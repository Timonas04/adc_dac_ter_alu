magic
tech sky130A
magscale 1 2
timestamp 1757960656
<< pwell >>
rect 2715 2465 2775 2541
rect 796 -1090 914 -12
rect 350 -4232 1606 -4142
rect 27757 -6782 28168 -6745
rect 27757 -6847 28061 -6782
<< psubdiff >>
rect 350 -4232 1606 -4142
<< locali >>
rect 350 -4232 1606 -4142
<< metal1 >>
rect 5577 3750 5773 3756
rect 975 3712 1034 3718
rect 443 1320 906 1713
rect 439 661 545 1161
rect 439 569 445 661
rect 537 569 545 661
rect 439 133 545 569
rect 801 128 911 1183
rect 434 -1054 540 -26
rect 796 -1090 914 -12
rect 431 -2279 549 -1212
rect 975 -1224 1034 3653
rect 2760 3284 2766 3369
rect 2851 3284 2984 3369
rect 5577 1982 5773 3614
rect 10640 3751 10855 3757
rect 7925 3352 7977 3358
rect 7925 3294 7977 3300
rect 10640 1801 10855 3620
rect 15643 3744 15851 3750
rect 12923 3352 12975 3358
rect 12923 3294 12975 3300
rect 15643 1908 15851 3618
rect 20651 3748 20843 3754
rect 25664 3750 25832 3760
rect 25664 3692 25678 3750
rect 17919 3352 17971 3358
rect 17913 3300 17919 3352
rect 17971 3300 17977 3352
rect 17919 3294 17971 3300
rect 20651 1954 20843 3626
rect 25814 3692 25832 3750
rect 30642 3750 30778 3756
rect 22919 3352 22971 3358
rect 22919 3294 22971 3300
rect 25678 2038 25814 3614
rect 27914 3352 27966 3358
rect 27914 3294 27966 3300
rect 30642 1920 30778 3614
rect 5665 -1119 5914 -1014
rect 5665 -1146 5968 -1119
rect 798 -1622 1034 -1224
rect 5704 -1251 5968 -1146
rect 975 -1623 1034 -1622
rect 807 -2057 1244 -1876
rect 807 -2189 1157 -2057
rect 1289 -2189 1394 -2057
rect 807 -2269 1244 -2189
rect 1262 -2410 1394 -2189
rect 440 -2819 877 -2426
rect 1710 -4168 1830 -4150
rect 1710 -4252 3990 -4168
rect 1710 -4342 1830 -4252
rect 1704 -4826 2102 -4708
rect 3906 -4890 3990 -4252
rect 5836 -4578 5968 -1251
rect 25652 -1279 25921 -1121
rect 21129 -2419 21417 -2261
rect 25763 -2377 25921 -1279
rect 21129 -2453 21287 -2419
rect 25763 -2541 25921 -2535
rect 21129 -2617 21287 -2611
rect 6328 -4228 9000 -4155
rect 5836 -4716 5968 -4710
rect 6592 -4810 6902 -4726
rect 6592 -4890 6676 -4810
rect 3906 -4974 6676 -4890
rect 8927 -4887 9000 -4228
rect 11208 -4240 14012 -4144
rect 16259 -4235 18997 -4148
rect 21269 -4235 24005 -4149
rect 26430 -4219 28991 -4165
rect 11549 -4805 12008 -4732
rect 11549 -4887 11622 -4805
rect 8927 -4960 11622 -4887
rect 13916 -4870 14012 -4240
rect 16466 -4812 17030 -4716
rect 16466 -4870 16562 -4812
rect 13916 -4966 16562 -4870
rect 18910 -4880 18997 -4235
rect 21446 -4812 22005 -4725
rect 21446 -4880 21533 -4812
rect 18910 -4967 21533 -4880
rect 23919 -4875 24005 -4235
rect 26465 -4815 26995 -4729
rect 28937 -4740 28991 -4219
rect 28937 -4794 29148 -4740
rect 26465 -4875 26551 -4815
rect 23919 -4961 26551 -4875
rect 28819 -4976 28977 -4970
rect 27466 -5029 27551 -5017
rect 24127 -5089 27551 -5029
rect 911 -5229 917 -5097
rect 1049 -5229 1055 -5097
rect 917 -5388 1049 -5229
rect 2232 -5247 5836 -5115
rect 5968 -5247 5974 -5115
rect 21123 -5334 21129 -5176
rect 21287 -5334 23868 -5176
rect 24127 -5199 24187 -5089
rect 25076 -5292 25763 -5134
rect 25921 -5292 25927 -5134
rect 25155 -5328 25252 -5292
rect 27466 -5454 27551 -5089
rect 28819 -5418 28977 -5134
rect 29094 -5335 29148 -4794
rect 29088 -5389 29094 -5335
rect 29148 -5389 29154 -5335
rect 1570 -6814 1675 -6711
rect 23965 -6814 24797 -6742
rect 28035 -6745 28217 -6743
rect 27757 -6814 28217 -6745
rect 28279 -6782 28300 -6738
rect 1570 -6884 28217 -6814
rect 1570 -6902 1675 -6884
<< via1 >>
rect 975 3653 1034 3712
rect 445 569 537 661
rect 5577 3614 5773 3750
rect 2766 3284 2851 3369
rect 10640 3620 10855 3751
rect 7925 3300 7977 3352
rect 15643 3618 15851 3744
rect 12923 3300 12975 3352
rect 20651 3626 20843 3748
rect 17919 3300 17971 3352
rect 25678 3614 25814 3750
rect 22919 3300 22971 3352
rect 30642 3614 30778 3750
rect 27914 3300 27966 3352
rect 1157 -2189 1289 -2057
rect 21129 -2611 21287 -2453
rect 25763 -2535 25921 -2377
rect 5836 -4710 5968 -4578
rect 917 -5229 1049 -5097
rect 5836 -5247 5968 -5115
rect 21129 -5334 21287 -5176
rect 25763 -5292 25921 -5134
rect 28819 -5134 28977 -4976
rect 29094 -5389 29148 -5335
<< metal2 >>
rect 10634 3750 10640 3751
rect 5571 3712 5577 3750
rect 969 3653 975 3712
rect 1034 3653 5577 3712
rect 5571 3614 5577 3653
rect 5773 3620 10640 3750
rect 10855 3750 10861 3751
rect 25666 3750 25888 3758
rect 10855 3748 25678 3750
rect 10855 3744 20651 3748
rect 10855 3620 15643 3744
rect 5773 3618 15643 3620
rect 15851 3626 20651 3744
rect 20843 3626 25678 3748
rect 15851 3618 25678 3626
rect 5773 3614 25678 3618
rect 25814 3614 30642 3750
rect 30778 3614 30784 3750
rect 3781 3409 28973 3536
rect 2766 3369 2851 3375
rect 1211 3284 2766 3369
rect 17919 3352 17971 3358
rect 7919 3351 7925 3352
rect 2851 3301 7925 3351
rect 7919 3300 7925 3301
rect 7977 3351 7983 3352
rect 12917 3351 12923 3352
rect 7977 3301 12923 3351
rect 7977 3300 7983 3301
rect 12917 3300 12923 3301
rect 12975 3351 12981 3352
rect 17913 3351 17919 3352
rect 12975 3301 17919 3351
rect 12975 3300 12981 3301
rect 17913 3300 17919 3301
rect 17971 3351 17977 3352
rect 22913 3351 22919 3352
rect 17971 3301 22919 3351
rect 17971 3300 17977 3301
rect 22913 3300 22919 3301
rect 22971 3351 22977 3352
rect 27908 3351 27914 3352
rect 22971 3301 27914 3351
rect 22971 3300 22977 3301
rect 27908 3300 27914 3301
rect 27966 3300 27972 3352
rect 17919 3294 17971 3300
rect 1211 661 1296 3284
rect 2766 3278 2851 3284
rect 439 569 445 661
rect 537 569 1299 661
rect 571 -5577 663 569
rect 26652 -640 26731 -333
rect 26043 -719 26731 -640
rect 1157 -2057 1289 -2051
rect 1157 -4981 1289 -2189
rect 21123 -2611 21129 -2453
rect 21287 -2611 21293 -2453
rect 25757 -2535 25763 -2377
rect 25921 -2535 25927 -2377
rect 5830 -4710 5836 -4578
rect 5968 -4710 5974 -4578
rect 917 -5097 1289 -4981
rect 1049 -5113 1289 -5097
rect 917 -5235 1049 -5229
rect 5836 -5115 5968 -4710
rect 5836 -5253 5968 -5247
rect 21129 -5176 21287 -2611
rect 25763 -4976 25921 -2535
rect 26043 -4670 26122 -719
rect 26043 -4758 26122 -4749
rect 25763 -5134 28819 -4976
rect 28977 -5134 28983 -4976
rect 25763 -5298 25921 -5292
rect 21129 -5340 21287 -5334
rect 24696 -5336 26122 -5330
rect 29094 -5335 29148 -5329
rect 24696 -5405 26048 -5336
rect 26117 -5405 26126 -5336
rect 28541 -5389 29094 -5335
rect 24696 -5409 26122 -5405
rect 571 -5669 1273 -5577
rect 24696 -5697 24775 -5409
rect 28541 -5734 28595 -5389
rect 29094 -5395 29148 -5389
<< via2 >>
rect 26043 -4749 26122 -4670
rect 26048 -5405 26117 -5336
<< metal3 >>
rect 26038 -4670 26127 -4665
rect 26038 -4749 26043 -4670
rect 26122 -4749 26127 -4670
rect 26038 -4754 26127 -4749
rect 26043 -5336 26122 -4754
rect 26043 -5405 26048 -5336
rect 26117 -5405 26122 -5336
rect 26043 -5410 26122 -5405
use anl_switch  anl_switch_0
timestamp 1757923025
transform 0 1 3602 -1 0 -3347
box 1756 -3202 3533 463
use anl_switch  anl_switch_1
timestamp 1757923025
transform 0 1 26402 -1 0 -3325
box 1756 -3202 3533 463
use anl_switch  anl_switch_2
timestamp 1757923025
transform 0 1 30202 -1 0 -3319
box 1756 -3202 3533 463
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_0
timestamp 1757903622
transform 0 1 987 -1 0 -4405
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_1
timestamp 1757903622
transform 1 0 857 0 1 -1147
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_2
timestamp 1757903622
transform 1 0 493 0 1 -1147
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_3
timestamp 1757903622
transform 1 0 857 0 1 49
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_4
timestamp 1757903622
transform 1 0 493 0 1 -2343
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_5
timestamp 1757903622
transform 1 0 857 0 1 -2343
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_6
timestamp 1757903622
transform 1 0 493 0 1 -3539
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_7
timestamp 1757903622
transform 1 0 857 0 1 -3539
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_8
timestamp 1757903622
transform 0 1 987 -1 0 -4769
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_9
timestamp 1757903622
transform 1 0 493 0 1 49
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_10
timestamp 1757903622
transform 1 0 493 0 1 1245
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_11
timestamp 1757903622
transform 1 0 857 0 1 1245
box -235 -651 235 651
use ter_dac_trit  ter_dac_trit_0
timestamp 1757960656
transform 0 1 -1028 -1 0 262
box -3396 2014 5266 6833
use ter_dac_trit  ter_dac_trit_1
timestamp 1757960656
transform 0 1 3986 -1 0 266
box -3396 2014 5266 6833
use ter_dac_trit  ter_dac_trit_2
timestamp 1757960656
transform 0 1 8986 -1 0 266
box -3396 2014 5266 6833
use ter_dac_trit  ter_dac_trit_3
timestamp 1757960656
transform 0 1 13986 -1 0 266
box -3396 2014 5266 6833
use ter_dac_trit  ter_dac_trit_4
timestamp 1757960656
transform 0 1 18986 -1 0 266
box -3396 2014 5266 6833
use ter_dac_trit  ter_dac_trit_5
timestamp 1757960656
transform 0 1 23986 -1 0 266
box -3396 2014 5266 6833
<< labels >>
rlabel space 22100 -6886 22738 -6809 1 a0
port 1 n
rlabel space 1528 -5299 1720 -5185 1 buffi_conn
port 2 n
rlabel space 28130 -5281 28322 -5158 1 DAC6_conn
port 19 n
rlabel space 24329 -5286 24515 -5163 1 buffo_conn
port 15 n
rlabel metal1 5597 2663 5763 3228 1 vdd
port 24 n
rlabel space 1139 -340 1242 209 1 vss
port 23 n
rlabel space 2060 -2635 2112 -2572 1 t0l
port 3 n
rlabel space 2936 -2635 2988 -2572 1 t0h
port 4 n
rlabel space 4119 -3784 4171 -3721 1 t0m
port 5 n
rlabel space 7596 -2629 7648 -2566 1 t1l
port 6 n
rlabel space 7948 -2633 8000 -2570 1 t1h
port 7 n
rlabel space 9134 -3775 9186 -3712 1 t1m
port 8 n
rlabel space 12599 -2633 12651 -2570 1 t2l
port 10 n
rlabel space 12950 -2632 13002 -2569 1 t2h
port 11 n
rlabel space 14145 -3774 14197 -3711 1 t2m
port 9 n
rlabel space 17600 -2630 17652 -2567 1 t3l
port 13 n
rlabel space 17949 -2633 18001 -2570 1 t3h
port 14 n
rlabel space 19144 -3767 19196 -3704 1 t3m
port 12 n
rlabel space 22597 -2629 22649 -2566 1 t4l
port 17 n
rlabel space 22950 -2629 23002 -2566 1 t4h
port 18 n
rlabel space 24132 -3774 24184 -3711 1 t4m
port 16 n
rlabel space 27073 -2628 27125 -2565 1 t5l
port 21 n
rlabel space 27950 -2631 28002 -2568 1 t5h
port 22 n
rlabel space 29139 -3769 29191 -3706 1 t5m
port 20 n
rlabel space 258 -6902 30819 3760 1 list
<< end >>
