MACRO r2r_dac
  CLASS BLOCK ;
  FOREIGN r2r_dac ;
  ORIGIN -14.505 113.075 ;
  SIZE 68.970 BY 14.235 ;
  PIN VDD
    ANTENNADIFFAREA 39.052799 ;
    PORT
      LAYER met1 ;
        RECT 42.560 -100.130 43.560 -99.130 ;
    END
  END VDD
  PIN B7
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 77.530 -108.625 78.530 -107.625 ;
    END
  END B7
  PIN B6
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 69.440 -108.585 70.440 -107.585 ;
    END
  END B6
  PIN B5
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 61.135 -108.615 62.135 -107.615 ;
    END
  END B5
  PIN B4
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 52.865 -108.600 53.865 -107.600 ;
    END
  END B4
  PIN B3
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 44.420 -108.560 45.420 -107.560 ;
    END
  END B3
  PIN B2
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 36.020 -108.720 37.020 -107.720 ;
    END
  END B2
  PIN B1
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 27.660 -108.605 28.660 -107.605 ;
    END
  END B1
  PIN B0
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met1 ;
        RECT 19.375 -108.600 20.375 -107.600 ;
    END
  END B0
  PIN OUT
    PORT
      LAYER met1 ;
        RECT 80.005 -106.990 81.005 -105.990 ;
    END
  END OUT
  PIN VSS
    ANTENNADIFFAREA 109.796898 ;
    PORT
      LAYER met1 ;
        RECT 42.730 -112.975 43.730 -111.975 ;
    END
  END VSS
  OBS
      LAYER pwell ;
        RECT 14.505 -112.365 18.675 -99.875 ;
      LAYER nwell ;
        RECT 18.795 -108.065 20.905 -99.875 ;
      LAYER pwell ;
        RECT 18.775 -112.360 20.885 -108.260 ;
        RECT 20.970 -112.350 26.960 -99.860 ;
      LAYER nwell ;
        RECT 27.090 -108.050 29.200 -99.860 ;
      LAYER pwell ;
        RECT 27.080 -112.360 29.190 -108.260 ;
        RECT 29.300 -112.360 35.290 -99.870 ;
      LAYER nwell ;
        RECT 35.405 -108.060 37.515 -99.870 ;
      LAYER pwell ;
        RECT 35.340 -112.360 37.450 -108.260 ;
        RECT 37.595 -112.370 43.585 -99.880 ;
      LAYER nwell ;
        RECT 43.785 -107.960 45.895 -99.770 ;
      LAYER pwell ;
        RECT 43.760 -112.340 45.870 -108.240 ;
        RECT 46.040 -112.355 52.030 -99.865 ;
      LAYER nwell ;
        RECT 52.175 -108.035 54.285 -99.845 ;
      LAYER pwell ;
        RECT 52.110 -112.360 54.220 -108.260 ;
        RECT 54.370 -112.355 60.360 -99.865 ;
      LAYER nwell ;
        RECT 60.505 -108.010 62.615 -99.820 ;
      LAYER pwell ;
        RECT 60.495 -112.365 62.605 -108.265 ;
        RECT 62.700 -112.355 68.690 -99.865 ;
      LAYER nwell ;
        RECT 68.800 -107.995 70.910 -99.805 ;
      LAYER pwell ;
        RECT 68.735 -112.355 70.845 -108.255 ;
        RECT 71.005 -112.360 76.995 -99.870 ;
      LAYER nwell ;
        RECT 77.100 -108.015 79.210 -99.825 ;
      LAYER pwell ;
        RECT 77.100 -112.355 79.210 -108.255 ;
        RECT 79.305 -112.350 83.475 -99.860 ;
      LAYER li1 ;
        RECT 19.200 -99.440 78.960 -98.990 ;
        RECT 19.200 -99.570 79.020 -99.440 ;
        RECT 18.980 -99.810 79.020 -99.570 ;
        RECT 18.980 -100.055 20.690 -99.810 ;
        RECT 27.270 -100.040 28.980 -99.810 ;
        RECT 14.685 -100.225 18.495 -100.055 ;
        RECT 14.685 -106.035 14.855 -100.225 ;
        RECT 15.335 -102.865 16.025 -100.705 ;
        RECT 15.335 -105.555 16.025 -103.395 ;
        RECT 16.505 -106.035 16.675 -100.225 ;
        RECT 17.155 -102.865 17.845 -100.705 ;
        RECT 17.155 -105.555 17.845 -103.395 ;
        RECT 18.325 -106.035 18.495 -100.225 ;
        RECT 14.685 -106.205 18.495 -106.035 ;
        RECT 14.685 -112.015 14.855 -106.205 ;
        RECT 15.335 -108.845 16.025 -106.685 ;
        RECT 15.335 -111.535 16.025 -109.375 ;
        RECT 16.505 -112.015 16.675 -106.205 ;
        RECT 17.155 -108.845 17.845 -106.685 ;
        RECT 17.155 -111.535 17.845 -109.375 ;
        RECT 18.325 -112.015 18.495 -106.205 ;
        RECT 18.975 -100.225 20.725 -100.055 ;
        RECT 18.975 -107.715 19.145 -100.225 ;
        RECT 19.685 -100.735 20.015 -100.565 ;
        RECT 19.545 -106.990 19.715 -100.950 ;
        RECT 19.985 -106.990 20.155 -100.950 ;
        RECT 19.685 -107.375 20.015 -107.205 ;
        RECT 20.555 -107.715 20.725 -100.225 ;
        RECT 18.975 -107.885 20.725 -107.715 ;
        RECT 21.150 -100.210 26.780 -100.040 ;
        RECT 21.150 -106.020 21.320 -100.210 ;
        RECT 21.800 -102.850 22.490 -100.690 ;
        RECT 21.800 -105.540 22.490 -103.380 ;
        RECT 22.970 -106.020 23.140 -100.210 ;
        RECT 23.620 -102.850 24.310 -100.690 ;
        RECT 23.620 -105.540 24.310 -103.380 ;
        RECT 24.790 -106.020 24.960 -100.210 ;
        RECT 25.440 -102.850 26.130 -100.690 ;
        RECT 25.440 -105.540 26.130 -103.380 ;
        RECT 26.610 -106.020 26.780 -100.210 ;
        RECT 21.150 -106.190 26.780 -106.020 ;
        RECT 18.955 -108.610 20.705 -108.440 ;
        RECT 18.955 -112.010 19.125 -108.610 ;
        RECT 19.665 -109.120 19.995 -108.950 ;
        RECT 19.525 -111.330 19.695 -109.290 ;
        RECT 19.965 -111.330 20.135 -109.290 ;
        RECT 19.665 -111.670 19.995 -111.500 ;
        RECT 20.535 -112.010 20.705 -108.610 ;
        RECT 18.955 -112.015 20.705 -112.010 ;
        RECT 21.150 -112.000 21.320 -106.190 ;
        RECT 21.800 -108.830 22.490 -106.670 ;
        RECT 21.800 -111.520 22.490 -109.360 ;
        RECT 22.970 -112.000 23.140 -106.190 ;
        RECT 23.620 -108.830 24.310 -106.670 ;
        RECT 23.620 -111.520 24.310 -109.360 ;
        RECT 24.790 -112.000 24.960 -106.190 ;
        RECT 25.440 -108.830 26.130 -106.670 ;
        RECT 25.440 -111.520 26.130 -109.360 ;
        RECT 26.610 -112.000 26.780 -106.190 ;
        RECT 27.270 -100.210 29.020 -100.040 ;
        RECT 27.270 -107.700 27.440 -100.210 ;
        RECT 27.980 -100.720 28.310 -100.550 ;
        RECT 27.840 -106.975 28.010 -100.935 ;
        RECT 28.280 -106.975 28.450 -100.935 ;
        RECT 27.980 -107.360 28.310 -107.190 ;
        RECT 28.850 -107.700 29.020 -100.210 ;
        RECT 27.270 -107.870 29.020 -107.700 ;
        RECT 29.480 -100.220 35.110 -100.050 ;
        RECT 29.480 -106.030 29.650 -100.220 ;
        RECT 30.130 -102.860 30.820 -100.700 ;
        RECT 30.130 -105.550 30.820 -103.390 ;
        RECT 31.300 -106.030 31.470 -100.220 ;
        RECT 31.950 -102.860 32.640 -100.700 ;
        RECT 31.950 -105.550 32.640 -103.390 ;
        RECT 33.120 -106.030 33.290 -100.220 ;
        RECT 33.770 -102.860 34.460 -100.700 ;
        RECT 33.770 -105.550 34.460 -103.390 ;
        RECT 34.940 -106.030 35.110 -100.220 ;
        RECT 35.410 -100.200 37.530 -99.810 ;
        RECT 43.920 -100.010 45.820 -99.810 ;
        RECT 35.410 -100.280 37.510 -100.200 ;
        RECT 37.775 -100.230 43.405 -100.060 ;
        RECT 29.480 -106.200 35.110 -106.030 ;
        RECT 21.150 -112.015 26.780 -112.000 ;
        RECT 27.260 -108.610 29.010 -108.440 ;
        RECT 27.260 -112.010 27.430 -108.610 ;
        RECT 27.970 -109.120 28.300 -108.950 ;
        RECT 27.830 -111.330 28.000 -109.290 ;
        RECT 28.270 -111.330 28.440 -109.290 ;
        RECT 27.970 -111.670 28.300 -111.500 ;
        RECT 28.840 -112.010 29.010 -108.610 ;
        RECT 27.260 -112.015 29.010 -112.010 ;
        RECT 29.480 -112.010 29.650 -106.200 ;
        RECT 30.130 -108.840 30.820 -106.680 ;
        RECT 30.130 -111.530 30.820 -109.370 ;
        RECT 31.300 -112.010 31.470 -106.200 ;
        RECT 31.950 -108.840 32.640 -106.680 ;
        RECT 31.950 -111.530 32.640 -109.370 ;
        RECT 33.120 -112.010 33.290 -106.200 ;
        RECT 33.770 -108.840 34.460 -106.680 ;
        RECT 33.770 -111.530 34.460 -109.370 ;
        RECT 34.940 -112.010 35.110 -106.200 ;
        RECT 35.585 -107.710 35.755 -100.280 ;
        RECT 36.295 -100.730 36.625 -100.560 ;
        RECT 36.155 -106.985 36.325 -100.945 ;
        RECT 36.595 -106.985 36.765 -100.945 ;
        RECT 36.295 -107.370 36.625 -107.200 ;
        RECT 37.165 -107.710 37.335 -100.280 ;
        RECT 35.585 -107.880 37.335 -107.710 ;
        RECT 37.775 -106.040 37.945 -100.230 ;
        RECT 38.425 -102.870 39.115 -100.710 ;
        RECT 38.425 -105.560 39.115 -103.400 ;
        RECT 39.595 -106.040 39.765 -100.230 ;
        RECT 40.245 -102.870 40.935 -100.710 ;
        RECT 40.245 -105.560 40.935 -103.400 ;
        RECT 41.415 -106.040 41.585 -100.230 ;
        RECT 42.065 -102.870 42.755 -100.710 ;
        RECT 42.065 -105.560 42.755 -103.400 ;
        RECT 43.235 -106.040 43.405 -100.230 ;
        RECT 37.775 -106.210 43.405 -106.040 ;
        RECT 29.480 -112.015 35.110 -112.010 ;
        RECT 35.520 -108.610 37.270 -108.440 ;
        RECT 35.520 -112.010 35.690 -108.610 ;
        RECT 36.230 -109.120 36.560 -108.950 ;
        RECT 36.090 -111.330 36.260 -109.290 ;
        RECT 36.530 -111.330 36.700 -109.290 ;
        RECT 36.230 -111.670 36.560 -111.500 ;
        RECT 37.100 -112.010 37.270 -108.610 ;
        RECT 35.520 -112.015 37.270 -112.010 ;
        RECT 37.775 -112.015 37.945 -106.210 ;
        RECT 38.425 -108.850 39.115 -106.690 ;
        RECT 38.425 -111.540 39.115 -109.380 ;
        RECT 39.595 -112.015 39.765 -106.210 ;
        RECT 40.245 -108.850 40.935 -106.690 ;
        RECT 40.245 -111.540 40.935 -109.380 ;
        RECT 41.415 -112.015 41.585 -106.210 ;
        RECT 42.065 -108.850 42.755 -106.690 ;
        RECT 42.065 -111.540 42.755 -109.380 ;
        RECT 43.235 -112.015 43.405 -106.210 ;
        RECT 43.965 -100.120 45.715 -100.010 ;
        RECT 52.360 -100.025 54.070 -99.810 ;
        RECT 60.690 -100.000 62.400 -99.810 ;
        RECT 68.980 -99.985 70.690 -99.810 ;
        RECT 43.965 -107.610 44.135 -100.120 ;
        RECT 44.675 -100.630 45.005 -100.460 ;
        RECT 44.535 -106.885 44.705 -100.845 ;
        RECT 44.975 -106.885 45.145 -100.845 ;
        RECT 44.675 -107.270 45.005 -107.100 ;
        RECT 45.545 -107.610 45.715 -100.120 ;
        RECT 43.965 -107.780 45.715 -107.610 ;
        RECT 46.220 -100.215 51.850 -100.045 ;
        RECT 46.220 -106.025 46.390 -100.215 ;
        RECT 46.870 -102.855 47.560 -100.695 ;
        RECT 46.870 -105.545 47.560 -103.385 ;
        RECT 48.040 -106.025 48.210 -100.215 ;
        RECT 48.690 -102.855 49.380 -100.695 ;
        RECT 48.690 -105.545 49.380 -103.385 ;
        RECT 49.860 -106.025 50.030 -100.215 ;
        RECT 50.510 -102.855 51.200 -100.695 ;
        RECT 50.510 -105.545 51.200 -103.385 ;
        RECT 51.680 -106.025 51.850 -100.215 ;
        RECT 46.220 -106.195 51.850 -106.025 ;
        RECT 43.940 -108.590 45.690 -108.420 ;
        RECT 43.940 -111.990 44.110 -108.590 ;
        RECT 44.650 -109.100 44.980 -108.930 ;
        RECT 44.510 -111.310 44.680 -109.270 ;
        RECT 44.950 -111.310 45.120 -109.270 ;
        RECT 44.650 -111.650 44.980 -111.480 ;
        RECT 45.520 -111.990 45.690 -108.590 ;
        RECT 43.940 -112.015 45.690 -111.990 ;
        RECT 46.220 -112.005 46.390 -106.195 ;
        RECT 46.870 -108.835 47.560 -106.675 ;
        RECT 46.870 -111.525 47.560 -109.365 ;
        RECT 48.040 -112.005 48.210 -106.195 ;
        RECT 48.690 -108.835 49.380 -106.675 ;
        RECT 48.690 -111.525 49.380 -109.365 ;
        RECT 49.860 -112.005 50.030 -106.195 ;
        RECT 50.510 -108.835 51.200 -106.675 ;
        RECT 50.510 -111.525 51.200 -109.365 ;
        RECT 51.680 -112.005 51.850 -106.195 ;
        RECT 52.355 -100.195 54.105 -100.025 ;
        RECT 52.355 -107.685 52.525 -100.195 ;
        RECT 53.065 -100.705 53.395 -100.535 ;
        RECT 52.925 -106.960 53.095 -100.920 ;
        RECT 53.365 -106.960 53.535 -100.920 ;
        RECT 53.065 -107.345 53.395 -107.175 ;
        RECT 53.935 -107.685 54.105 -100.195 ;
        RECT 52.355 -107.855 54.105 -107.685 ;
        RECT 54.550 -100.215 60.180 -100.045 ;
        RECT 54.550 -106.025 54.720 -100.215 ;
        RECT 55.200 -102.855 55.890 -100.695 ;
        RECT 55.200 -105.545 55.890 -103.385 ;
        RECT 56.370 -106.025 56.540 -100.215 ;
        RECT 57.020 -102.855 57.710 -100.695 ;
        RECT 57.020 -105.545 57.710 -103.385 ;
        RECT 58.190 -106.025 58.360 -100.215 ;
        RECT 58.840 -102.855 59.530 -100.695 ;
        RECT 58.840 -105.545 59.530 -103.385 ;
        RECT 60.010 -106.025 60.180 -100.215 ;
        RECT 54.550 -106.195 60.180 -106.025 ;
        RECT 46.220 -112.015 51.850 -112.005 ;
        RECT 52.290 -108.610 54.040 -108.440 ;
        RECT 52.290 -112.010 52.460 -108.610 ;
        RECT 53.000 -109.120 53.330 -108.950 ;
        RECT 52.860 -111.330 53.030 -109.290 ;
        RECT 53.300 -111.330 53.470 -109.290 ;
        RECT 53.000 -111.670 53.330 -111.500 ;
        RECT 53.870 -112.010 54.040 -108.610 ;
        RECT 52.290 -112.015 54.040 -112.010 ;
        RECT 54.550 -112.005 54.720 -106.195 ;
        RECT 55.200 -108.835 55.890 -106.675 ;
        RECT 55.200 -111.525 55.890 -109.365 ;
        RECT 56.370 -112.005 56.540 -106.195 ;
        RECT 57.020 -108.835 57.710 -106.675 ;
        RECT 57.020 -111.525 57.710 -109.365 ;
        RECT 58.190 -112.005 58.360 -106.195 ;
        RECT 58.840 -108.835 59.530 -106.675 ;
        RECT 58.840 -111.525 59.530 -109.365 ;
        RECT 60.010 -112.005 60.180 -106.195 ;
        RECT 60.685 -100.170 62.435 -100.000 ;
        RECT 60.685 -107.660 60.855 -100.170 ;
        RECT 61.395 -100.680 61.725 -100.510 ;
        RECT 61.255 -106.935 61.425 -100.895 ;
        RECT 61.695 -106.935 61.865 -100.895 ;
        RECT 61.395 -107.320 61.725 -107.150 ;
        RECT 62.265 -107.660 62.435 -100.170 ;
        RECT 60.685 -107.830 62.435 -107.660 ;
        RECT 62.880 -100.215 68.510 -100.045 ;
        RECT 62.880 -106.025 63.050 -100.215 ;
        RECT 63.530 -102.855 64.220 -100.695 ;
        RECT 63.530 -105.545 64.220 -103.385 ;
        RECT 64.700 -106.025 64.870 -100.215 ;
        RECT 65.350 -102.855 66.040 -100.695 ;
        RECT 65.350 -105.545 66.040 -103.385 ;
        RECT 66.520 -106.025 66.690 -100.215 ;
        RECT 67.170 -102.855 67.860 -100.695 ;
        RECT 67.170 -105.545 67.860 -103.385 ;
        RECT 68.340 -106.025 68.510 -100.215 ;
        RECT 62.880 -106.195 68.510 -106.025 ;
        RECT 54.550 -112.015 60.180 -112.005 ;
        RECT 60.675 -108.615 62.425 -108.445 ;
        RECT 60.675 -112.015 60.845 -108.615 ;
        RECT 61.385 -109.125 61.715 -108.955 ;
        RECT 61.245 -111.335 61.415 -109.295 ;
        RECT 61.685 -111.335 61.855 -109.295 ;
        RECT 61.385 -111.675 61.715 -111.505 ;
        RECT 62.255 -112.015 62.425 -108.615 ;
        RECT 62.880 -112.005 63.050 -106.195 ;
        RECT 63.530 -108.835 64.220 -106.675 ;
        RECT 63.530 -111.525 64.220 -109.365 ;
        RECT 64.700 -112.005 64.870 -106.195 ;
        RECT 65.350 -108.835 66.040 -106.675 ;
        RECT 65.350 -111.525 66.040 -109.365 ;
        RECT 66.520 -112.005 66.690 -106.195 ;
        RECT 67.170 -108.835 67.860 -106.675 ;
        RECT 67.170 -111.525 67.860 -109.365 ;
        RECT 68.340 -112.005 68.510 -106.195 ;
        RECT 68.980 -100.155 70.730 -99.985 ;
        RECT 77.310 -100.005 79.020 -99.810 ;
        RECT 68.980 -107.645 69.150 -100.155 ;
        RECT 69.690 -100.665 70.020 -100.495 ;
        RECT 69.550 -106.920 69.720 -100.880 ;
        RECT 69.990 -106.920 70.160 -100.880 ;
        RECT 69.690 -107.305 70.020 -107.135 ;
        RECT 70.560 -107.645 70.730 -100.155 ;
        RECT 68.980 -107.815 70.730 -107.645 ;
        RECT 71.185 -100.220 76.815 -100.050 ;
        RECT 71.185 -106.030 71.355 -100.220 ;
        RECT 71.835 -102.860 72.525 -100.700 ;
        RECT 71.835 -105.550 72.525 -103.390 ;
        RECT 73.005 -106.030 73.175 -100.220 ;
        RECT 73.655 -102.860 74.345 -100.700 ;
        RECT 73.655 -105.550 74.345 -103.390 ;
        RECT 74.825 -106.030 74.995 -100.220 ;
        RECT 75.475 -102.860 76.165 -100.700 ;
        RECT 75.475 -105.550 76.165 -103.390 ;
        RECT 76.645 -106.030 76.815 -100.220 ;
        RECT 71.185 -106.200 76.815 -106.030 ;
        RECT 62.880 -112.015 68.510 -112.005 ;
        RECT 68.915 -108.605 70.665 -108.435 ;
        RECT 68.915 -112.005 69.085 -108.605 ;
        RECT 69.625 -109.115 69.955 -108.945 ;
        RECT 69.485 -111.325 69.655 -109.285 ;
        RECT 69.925 -111.325 70.095 -109.285 ;
        RECT 69.625 -111.665 69.955 -111.495 ;
        RECT 70.495 -112.005 70.665 -108.605 ;
        RECT 68.915 -112.015 70.665 -112.005 ;
        RECT 71.185 -112.010 71.355 -106.200 ;
        RECT 71.835 -108.840 72.525 -106.680 ;
        RECT 71.835 -111.530 72.525 -109.370 ;
        RECT 73.005 -112.010 73.175 -106.200 ;
        RECT 73.655 -108.840 74.345 -106.680 ;
        RECT 73.655 -111.530 74.345 -109.370 ;
        RECT 74.825 -112.010 74.995 -106.200 ;
        RECT 75.475 -108.840 76.165 -106.680 ;
        RECT 75.475 -111.530 76.165 -109.370 ;
        RECT 76.645 -112.010 76.815 -106.200 ;
        RECT 77.280 -100.175 79.030 -100.005 ;
        RECT 77.280 -107.665 77.450 -100.175 ;
        RECT 77.990 -100.685 78.320 -100.515 ;
        RECT 77.850 -106.940 78.020 -100.900 ;
        RECT 78.290 -106.940 78.460 -100.900 ;
        RECT 77.990 -107.325 78.320 -107.155 ;
        RECT 78.860 -107.665 79.030 -100.175 ;
        RECT 77.280 -107.835 79.030 -107.665 ;
        RECT 79.485 -100.210 83.295 -100.040 ;
        RECT 79.485 -106.020 79.655 -100.210 ;
        RECT 80.135 -102.850 80.825 -100.690 ;
        RECT 80.135 -105.540 80.825 -103.380 ;
        RECT 81.305 -106.020 81.475 -100.210 ;
        RECT 81.955 -102.850 82.645 -100.690 ;
        RECT 81.955 -105.540 82.645 -103.380 ;
        RECT 83.125 -106.020 83.295 -100.210 ;
        RECT 79.485 -106.190 83.295 -106.020 ;
        RECT 71.185 -112.015 76.815 -112.010 ;
        RECT 77.280 -108.605 79.030 -108.435 ;
        RECT 77.280 -112.005 77.450 -108.605 ;
        RECT 77.990 -109.115 78.320 -108.945 ;
        RECT 77.850 -111.325 78.020 -109.285 ;
        RECT 78.290 -111.325 78.460 -109.285 ;
        RECT 77.990 -111.665 78.320 -111.495 ;
        RECT 78.860 -112.005 79.030 -108.605 ;
        RECT 77.280 -112.015 79.030 -112.005 ;
        RECT 79.485 -112.000 79.655 -106.190 ;
        RECT 80.135 -108.830 80.825 -106.670 ;
        RECT 80.135 -111.520 80.825 -109.360 ;
        RECT 81.305 -112.000 81.475 -106.190 ;
        RECT 81.955 -108.830 82.645 -106.670 ;
        RECT 81.955 -111.520 82.645 -109.360 ;
        RECT 83.125 -112.000 83.295 -106.190 ;
        RECT 79.485 -112.015 83.295 -112.000 ;
        RECT 14.685 -112.890 83.300 -112.015 ;
      LAYER met1 ;
        RECT 45.940 -98.845 46.580 -98.840 ;
        RECT 19.045 -98.850 46.580 -98.845 ;
        RECT 49.570 -98.845 50.300 -98.840 ;
        RECT 49.570 -98.850 79.150 -98.845 ;
        RECT 19.045 -99.130 79.150 -98.850 ;
        RECT 19.045 -99.385 42.560 -99.130 ;
        RECT 18.740 -100.130 42.560 -99.385 ;
        RECT 43.560 -100.085 79.150 -99.130 ;
        RECT 43.560 -100.130 44.390 -100.085 ;
        RECT 18.740 -100.250 44.390 -100.130 ;
        RECT 45.380 -100.250 79.150 -100.085 ;
        RECT 15.385 -100.785 15.975 -100.735 ;
        RECT 17.205 -100.785 17.795 -100.735 ;
        RECT 15.385 -102.740 17.795 -100.785 ;
        RECT 18.740 -101.015 19.200 -100.250 ;
        RECT 19.700 -100.765 20.015 -100.475 ;
        RECT 19.515 -101.015 19.745 -100.970 ;
        RECT 18.740 -101.685 19.745 -101.015 ;
        RECT 15.385 -102.840 15.975 -102.740 ;
        RECT 17.205 -102.840 17.795 -102.740 ;
        RECT 15.385 -103.745 15.975 -103.420 ;
        RECT 17.205 -103.725 17.795 -103.420 ;
        RECT 15.365 -108.765 15.990 -103.745 ;
        RECT 17.180 -108.745 17.805 -103.725 ;
        RECT 19.150 -106.890 19.745 -101.685 ;
        RECT 19.515 -106.970 19.745 -106.890 ;
        RECT 19.955 -101.030 20.185 -100.970 ;
        RECT 21.850 -101.015 22.440 -100.720 ;
        RECT 20.445 -101.030 22.440 -101.015 ;
        RECT 19.955 -102.800 22.440 -101.030 ;
        RECT 19.955 -104.410 20.860 -102.800 ;
        RECT 21.850 -102.825 22.440 -102.800 ;
        RECT 23.670 -100.815 24.260 -100.720 ;
        RECT 25.490 -100.815 26.080 -100.720 ;
        RECT 23.670 -102.600 26.080 -100.815 ;
        RECT 27.035 -101.015 27.495 -100.250 ;
        RECT 28.000 -100.740 28.315 -100.450 ;
        RECT 28.000 -100.750 28.290 -100.740 ;
        RECT 30.180 -100.930 30.770 -100.730 ;
        RECT 27.810 -101.015 28.040 -100.955 ;
        RECT 27.035 -101.845 28.040 -101.015 ;
        RECT 23.670 -102.825 24.260 -102.600 ;
        RECT 25.490 -102.825 26.080 -102.600 ;
        RECT 21.850 -103.585 22.440 -103.405 ;
        RECT 23.670 -103.585 24.260 -103.405 ;
        RECT 19.955 -106.865 20.985 -104.410 ;
        RECT 21.850 -105.370 24.260 -103.585 ;
        RECT 25.490 -103.735 26.080 -103.405 ;
        RECT 21.850 -105.510 22.440 -105.370 ;
        RECT 23.670 -105.510 24.260 -105.370 ;
        RECT 25.465 -105.510 26.080 -103.735 ;
        RECT 25.465 -106.700 25.995 -105.510 ;
        RECT 19.955 -106.970 20.185 -106.865 ;
        RECT 19.710 -107.175 20.040 -107.170 ;
        RECT 19.705 -107.405 20.040 -107.175 ;
        RECT 19.710 -107.430 20.040 -107.405 ;
        RECT 19.710 -107.600 19.970 -107.430 ;
        RECT 15.385 -108.820 15.975 -108.765 ;
        RECT 17.205 -108.820 17.795 -108.745 ;
        RECT 19.710 -108.920 20.040 -108.600 ;
        RECT 19.685 -109.135 20.040 -108.920 ;
        RECT 19.685 -109.150 19.975 -109.135 ;
        RECT 19.495 -109.370 19.725 -109.310 ;
        RECT 15.385 -109.490 15.975 -109.400 ;
        RECT 15.265 -112.015 15.990 -109.490 ;
        RECT 17.205 -109.500 17.795 -109.400 ;
        RECT 17.200 -111.595 17.795 -109.500 ;
        RECT 19.060 -110.155 19.725 -109.370 ;
        RECT 18.700 -111.240 19.725 -110.155 ;
        RECT 17.200 -112.015 17.795 -112.005 ;
        RECT 18.700 -112.015 19.160 -111.240 ;
        RECT 19.495 -111.310 19.725 -111.240 ;
        RECT 19.935 -109.380 20.165 -109.310 ;
        RECT 20.610 -109.380 20.985 -106.865 ;
        RECT 21.850 -106.880 22.440 -106.700 ;
        RECT 23.670 -106.880 24.260 -106.700 ;
        RECT 21.850 -108.665 24.260 -106.880 ;
        RECT 21.850 -108.805 22.440 -108.665 ;
        RECT 23.670 -108.805 24.260 -108.665 ;
        RECT 25.465 -108.680 26.080 -106.700 ;
        RECT 27.365 -106.890 28.040 -101.845 ;
        RECT 27.810 -106.955 28.040 -106.890 ;
        RECT 28.250 -101.010 28.480 -100.955 ;
        RECT 28.675 -101.010 30.770 -100.930 ;
        RECT 28.250 -102.715 30.770 -101.010 ;
        RECT 28.250 -104.295 29.195 -102.715 ;
        RECT 30.180 -102.835 30.770 -102.715 ;
        RECT 32.000 -100.980 32.590 -100.730 ;
        RECT 33.820 -100.980 34.410 -100.730 ;
        RECT 32.000 -102.765 34.410 -100.980 ;
        RECT 35.370 -101.035 35.830 -100.250 ;
        RECT 36.315 -100.765 36.630 -100.475 ;
        RECT 36.125 -101.035 36.355 -100.965 ;
        RECT 35.370 -101.835 36.355 -101.035 ;
        RECT 32.000 -102.835 32.590 -102.765 ;
        RECT 33.820 -102.835 34.410 -102.765 ;
        RECT 30.180 -103.670 30.770 -103.415 ;
        RECT 32.000 -103.670 32.590 -103.415 ;
        RECT 28.250 -106.845 29.375 -104.295 ;
        RECT 30.180 -105.455 32.590 -103.670 ;
        RECT 33.820 -103.745 34.410 -103.415 ;
        RECT 30.180 -105.520 30.770 -105.455 ;
        RECT 32.000 -105.520 32.590 -105.455 ;
        RECT 28.250 -106.955 28.480 -106.845 ;
        RECT 28.000 -107.190 28.290 -107.160 ;
        RECT 27.990 -107.605 28.320 -107.190 ;
        RECT 25.490 -108.805 26.080 -108.680 ;
        RECT 27.990 -109.155 28.320 -108.605 ;
        RECT 19.935 -111.200 21.010 -109.380 ;
        RECT 19.935 -111.310 20.165 -111.200 ;
        RECT 19.685 -111.755 20.000 -111.465 ;
        RECT 21.850 -111.490 22.440 -109.385 ;
        RECT 23.670 -109.600 24.260 -109.385 ;
        RECT 24.490 -109.600 25.085 -109.525 ;
        RECT 25.490 -109.600 26.080 -109.385 ;
        RECT 27.800 -109.400 28.030 -109.310 ;
        RECT 28.240 -109.390 28.470 -109.310 ;
        RECT 29.000 -109.390 29.375 -106.845 ;
        RECT 30.180 -106.840 30.770 -106.710 ;
        RECT 32.000 -106.840 32.590 -106.710 ;
        RECT 30.180 -108.625 32.590 -106.840 ;
        RECT 30.180 -108.815 30.770 -108.625 ;
        RECT 32.000 -108.815 32.590 -108.625 ;
        RECT 33.810 -108.765 34.435 -103.745 ;
        RECT 35.720 -106.910 36.355 -101.835 ;
        RECT 36.125 -106.965 36.355 -106.910 ;
        RECT 36.565 -100.985 36.795 -100.965 ;
        RECT 36.565 -101.005 37.490 -100.985 ;
        RECT 38.475 -101.005 39.065 -100.740 ;
        RECT 36.565 -102.820 39.065 -101.005 ;
        RECT 36.565 -104.420 37.490 -102.820 ;
        RECT 38.475 -102.845 39.065 -102.820 ;
        RECT 40.295 -100.925 40.885 -100.740 ;
        RECT 42.115 -100.925 42.705 -100.740 ;
        RECT 40.295 -102.740 42.705 -100.925 ;
        RECT 43.745 -100.895 44.205 -100.250 ;
        RECT 44.680 -100.640 44.995 -100.350 ;
        RECT 44.695 -100.660 44.985 -100.640 ;
        RECT 44.505 -100.895 44.735 -100.865 ;
        RECT 43.745 -101.455 44.735 -100.895 ;
        RECT 40.295 -102.845 40.885 -102.740 ;
        RECT 42.115 -102.845 42.705 -102.740 ;
        RECT 38.475 -103.565 39.065 -103.425 ;
        RECT 40.295 -103.565 40.885 -103.425 ;
        RECT 36.565 -106.820 37.565 -104.420 ;
        RECT 38.475 -105.380 40.885 -103.565 ;
        RECT 38.475 -105.530 39.065 -105.380 ;
        RECT 40.295 -105.530 40.885 -105.380 ;
        RECT 42.115 -103.705 42.705 -103.425 ;
        RECT 36.565 -106.965 36.795 -106.820 ;
        RECT 36.280 -107.400 36.605 -107.170 ;
        RECT 36.280 -107.720 36.540 -107.400 ;
        RECT 33.820 -108.815 34.410 -108.765 ;
        RECT 36.280 -108.920 36.540 -108.720 ;
        RECT 36.250 -109.150 36.540 -108.920 ;
        RECT 23.670 -111.385 26.080 -109.600 ;
        RECT 27.445 -110.005 28.045 -109.400 ;
        RECT 23.670 -111.490 24.260 -111.385 ;
        RECT 25.490 -111.490 26.080 -111.385 ;
        RECT 27.125 -111.270 28.045 -110.005 ;
        RECT 28.240 -111.080 29.375 -109.390 ;
        RECT 28.240 -111.210 29.290 -111.080 ;
        RECT 27.125 -112.015 27.585 -111.270 ;
        RECT 27.800 -111.310 28.030 -111.270 ;
        RECT 28.240 -111.310 28.470 -111.210 ;
        RECT 27.990 -111.745 28.305 -111.455 ;
        RECT 30.180 -111.500 30.770 -109.395 ;
        RECT 32.000 -109.660 32.590 -109.395 ;
        RECT 32.745 -109.660 33.335 -109.595 ;
        RECT 33.820 -109.660 34.410 -109.395 ;
        RECT 36.060 -109.410 36.290 -109.310 ;
        RECT 32.000 -111.445 34.410 -109.660 ;
        RECT 35.670 -109.995 36.290 -109.410 ;
        RECT 32.000 -111.500 32.590 -111.445 ;
        RECT 33.820 -111.500 34.410 -111.445 ;
        RECT 35.320 -111.280 36.290 -109.995 ;
        RECT 30.195 -111.525 30.740 -111.500 ;
        RECT 35.320 -112.015 35.780 -111.280 ;
        RECT 36.060 -111.310 36.290 -111.280 ;
        RECT 36.500 -109.405 36.730 -109.310 ;
        RECT 37.190 -109.405 37.565 -106.820 ;
        RECT 38.475 -106.870 39.065 -106.720 ;
        RECT 40.295 -106.870 40.885 -106.720 ;
        RECT 38.475 -108.685 40.885 -106.870 ;
        RECT 38.475 -108.825 39.065 -108.685 ;
        RECT 40.295 -108.825 40.885 -108.685 ;
        RECT 42.115 -108.725 42.740 -103.705 ;
        RECT 44.065 -106.770 44.735 -101.455 ;
        RECT 44.505 -106.865 44.735 -106.770 ;
        RECT 44.945 -100.935 45.175 -100.865 ;
        RECT 44.945 -100.985 45.845 -100.935 ;
        RECT 46.920 -100.985 47.510 -100.725 ;
        RECT 44.945 -102.800 47.510 -100.985 ;
        RECT 44.945 -104.370 45.845 -102.800 ;
        RECT 46.920 -102.830 47.510 -102.800 ;
        RECT 48.740 -100.865 49.330 -100.725 ;
        RECT 50.560 -100.865 51.150 -100.725 ;
        RECT 48.740 -102.680 51.150 -100.865 ;
        RECT 52.170 -100.985 52.630 -100.250 ;
        RECT 53.085 -100.725 53.400 -100.435 ;
        RECT 53.085 -100.735 53.375 -100.725 ;
        RECT 55.250 -100.925 55.840 -100.725 ;
        RECT 53.400 -100.940 55.840 -100.925 ;
        RECT 52.895 -100.985 53.125 -100.940 ;
        RECT 52.170 -101.475 53.125 -100.985 ;
        RECT 48.740 -102.830 49.330 -102.680 ;
        RECT 50.560 -102.830 51.150 -102.680 ;
        RECT 46.920 -103.665 47.510 -103.410 ;
        RECT 48.740 -103.665 49.330 -103.410 ;
        RECT 50.560 -103.480 51.150 -103.410 ;
        RECT 44.945 -106.770 45.970 -104.370 ;
        RECT 46.920 -105.480 49.330 -103.665 ;
        RECT 46.920 -105.515 47.510 -105.480 ;
        RECT 48.740 -105.515 49.330 -105.480 ;
        RECT 44.945 -106.865 45.175 -106.770 ;
        RECT 44.695 -107.300 44.985 -107.070 ;
        RECT 44.705 -107.560 44.955 -107.300 ;
        RECT 42.115 -108.825 42.705 -108.725 ;
        RECT 44.705 -108.900 44.955 -108.560 ;
        RECT 44.670 -109.130 44.960 -108.900 ;
        RECT 44.480 -109.370 44.710 -109.290 ;
        RECT 36.500 -111.225 37.585 -109.405 ;
        RECT 38.475 -109.555 39.065 -109.405 ;
        RECT 36.500 -111.310 36.730 -111.225 ;
        RECT 36.250 -111.490 36.540 -111.470 ;
        RECT 36.250 -111.700 36.605 -111.490 ;
        RECT 38.465 -111.510 39.065 -109.555 ;
        RECT 40.295 -109.650 40.885 -109.405 ;
        RECT 42.115 -109.650 42.705 -109.405 ;
        RECT 40.295 -111.465 42.705 -109.650 ;
        RECT 44.045 -109.855 44.710 -109.370 ;
        RECT 43.725 -109.905 44.710 -109.855 ;
        RECT 40.295 -111.510 40.885 -111.465 ;
        RECT 42.115 -111.510 42.705 -111.465 ;
        RECT 43.575 -111.240 44.710 -109.905 ;
        RECT 38.465 -111.545 39.010 -111.510 ;
        RECT 36.290 -111.780 36.605 -111.700 ;
        RECT 43.575 -111.975 44.185 -111.240 ;
        RECT 44.480 -111.290 44.710 -111.240 ;
        RECT 44.920 -109.380 45.150 -109.290 ;
        RECT 45.595 -109.380 45.970 -106.770 ;
        RECT 46.920 -106.970 47.510 -106.705 ;
        RECT 48.740 -106.970 49.330 -106.705 ;
        RECT 46.920 -108.785 49.330 -106.970 ;
        RECT 46.920 -108.810 47.510 -108.785 ;
        RECT 48.740 -108.810 49.330 -108.785 ;
        RECT 50.540 -108.800 51.160 -103.480 ;
        RECT 52.540 -106.860 53.125 -101.475 ;
        RECT 52.895 -106.940 53.125 -106.860 ;
        RECT 53.335 -102.740 55.840 -100.940 ;
        RECT 53.335 -104.435 54.225 -102.740 ;
        RECT 55.250 -102.830 55.840 -102.740 ;
        RECT 57.070 -100.885 57.660 -100.725 ;
        RECT 58.890 -100.885 59.480 -100.725 ;
        RECT 57.070 -102.700 59.480 -100.885 ;
        RECT 60.625 -100.935 61.085 -100.250 ;
        RECT 61.400 -100.690 61.715 -100.400 ;
        RECT 61.415 -100.710 61.705 -100.690 ;
        RECT 61.225 -100.935 61.455 -100.915 ;
        RECT 60.625 -101.755 61.455 -100.935 ;
        RECT 57.070 -102.830 57.660 -102.700 ;
        RECT 58.890 -102.830 59.480 -102.700 ;
        RECT 55.250 -103.625 55.840 -103.410 ;
        RECT 57.070 -103.625 57.660 -103.410 ;
        RECT 53.335 -106.870 54.450 -104.435 ;
        RECT 55.250 -105.440 57.660 -103.625 ;
        RECT 58.890 -103.705 59.480 -103.410 ;
        RECT 55.250 -105.515 55.840 -105.440 ;
        RECT 57.070 -105.515 57.660 -105.440 ;
        RECT 53.335 -106.940 53.565 -106.870 ;
        RECT 53.080 -107.145 53.330 -107.135 ;
        RECT 53.080 -107.375 53.375 -107.145 ;
        RECT 53.080 -107.600 53.330 -107.375 ;
        RECT 50.560 -108.810 51.150 -108.800 ;
        RECT 53.080 -108.920 53.330 -108.600 ;
        RECT 53.020 -109.120 53.330 -108.920 ;
        RECT 53.020 -109.150 53.310 -109.120 ;
        RECT 44.920 -111.200 45.970 -109.380 ;
        RECT 52.830 -109.390 53.060 -109.310 ;
        RECT 44.920 -111.290 45.150 -111.200 ;
        RECT 44.670 -111.465 44.960 -111.450 ;
        RECT 44.655 -111.755 44.970 -111.465 ;
        RECT 46.920 -111.510 47.510 -109.390 ;
        RECT 48.740 -109.630 49.330 -109.390 ;
        RECT 50.560 -109.630 51.150 -109.390 ;
        RECT 48.740 -111.445 51.150 -109.630 ;
        RECT 52.410 -109.845 53.060 -109.390 ;
        RECT 48.740 -111.495 49.330 -111.445 ;
        RECT 50.560 -111.495 51.150 -111.445 ;
        RECT 51.970 -111.290 53.060 -109.845 ;
        RECT 43.730 -112.015 44.185 -111.975 ;
        RECT 51.970 -112.015 52.430 -111.290 ;
        RECT 52.830 -111.310 53.060 -111.290 ;
        RECT 53.270 -109.430 53.500 -109.310 ;
        RECT 54.075 -109.430 54.450 -106.870 ;
        RECT 55.250 -106.890 55.840 -106.705 ;
        RECT 57.070 -106.890 57.660 -106.705 ;
        RECT 55.250 -108.705 57.660 -106.890 ;
        RECT 55.250 -108.810 55.840 -108.705 ;
        RECT 57.070 -108.810 57.660 -108.705 ;
        RECT 58.865 -108.725 59.490 -103.705 ;
        RECT 60.795 -106.810 61.455 -101.755 ;
        RECT 61.225 -106.915 61.455 -106.810 ;
        RECT 61.665 -101.000 61.895 -100.915 ;
        RECT 61.665 -101.005 62.585 -101.000 ;
        RECT 63.580 -101.005 64.170 -100.725 ;
        RECT 61.665 -102.820 64.170 -101.005 ;
        RECT 61.665 -104.410 62.585 -102.820 ;
        RECT 63.580 -102.830 64.170 -102.820 ;
        RECT 65.400 -100.905 65.990 -100.725 ;
        RECT 67.220 -100.905 67.810 -100.725 ;
        RECT 65.400 -102.720 67.810 -100.905 ;
        RECT 68.865 -100.975 69.325 -100.250 ;
        RECT 69.705 -100.715 70.020 -100.425 ;
        RECT 69.520 -100.975 69.750 -100.900 ;
        RECT 68.865 -101.705 69.750 -100.975 ;
        RECT 65.400 -102.830 65.990 -102.720 ;
        RECT 67.220 -102.830 67.810 -102.720 ;
        RECT 63.580 -103.665 64.170 -103.410 ;
        RECT 65.400 -103.665 65.990 -103.410 ;
        RECT 67.220 -103.665 67.810 -103.410 ;
        RECT 61.665 -106.835 62.780 -104.410 ;
        RECT 63.580 -105.480 66.000 -103.665 ;
        RECT 63.580 -105.515 64.170 -105.480 ;
        RECT 65.400 -105.515 65.990 -105.480 ;
        RECT 61.665 -106.915 61.895 -106.835 ;
        RECT 61.415 -107.350 61.705 -107.120 ;
        RECT 61.415 -107.615 61.665 -107.350 ;
        RECT 58.890 -108.810 59.480 -108.725 ;
        RECT 61.415 -108.925 61.665 -108.615 ;
        RECT 61.405 -109.155 61.695 -108.925 ;
        RECT 61.215 -109.370 61.445 -109.315 ;
        RECT 53.270 -111.220 54.450 -109.430 ;
        RECT 55.250 -109.405 55.840 -109.390 ;
        RECT 53.270 -111.250 54.335 -111.220 ;
        RECT 53.270 -111.310 53.500 -111.250 ;
        RECT 55.250 -111.425 55.845 -109.405 ;
        RECT 57.070 -109.610 57.660 -109.390 ;
        RECT 58.890 -109.610 59.480 -109.390 ;
        RECT 57.070 -111.425 59.480 -109.610 ;
        RECT 60.815 -109.835 61.445 -109.370 ;
        RECT 53.010 -111.745 53.325 -111.455 ;
        RECT 55.250 -111.495 55.840 -111.425 ;
        RECT 57.070 -111.495 57.660 -111.425 ;
        RECT 57.880 -111.510 58.470 -111.425 ;
        RECT 58.890 -111.495 59.480 -111.425 ;
        RECT 60.405 -111.270 61.445 -109.835 ;
        RECT 60.405 -112.015 60.865 -111.270 ;
        RECT 61.215 -111.315 61.445 -111.270 ;
        RECT 61.655 -109.440 61.885 -109.315 ;
        RECT 62.405 -109.440 62.780 -106.835 ;
        RECT 63.580 -106.910 64.170 -106.705 ;
        RECT 65.400 -106.910 65.990 -106.705 ;
        RECT 63.580 -108.725 65.990 -106.910 ;
        RECT 67.185 -108.685 67.810 -103.665 ;
        RECT 69.075 -106.850 69.750 -101.705 ;
        RECT 69.520 -106.900 69.750 -106.850 ;
        RECT 69.960 -101.005 70.190 -100.900 ;
        RECT 71.885 -101.005 72.475 -100.730 ;
        RECT 69.960 -102.820 72.475 -101.005 ;
        RECT 69.960 -104.310 70.865 -102.820 ;
        RECT 71.885 -102.835 72.475 -102.820 ;
        RECT 73.705 -100.905 74.295 -100.730 ;
        RECT 75.525 -100.905 76.115 -100.730 ;
        RECT 73.705 -102.720 76.115 -100.905 ;
        RECT 77.140 -100.975 77.600 -100.250 ;
        RECT 78.020 -100.485 78.335 -100.410 ;
        RECT 78.010 -100.700 78.335 -100.485 ;
        RECT 78.010 -100.715 78.300 -100.700 ;
        RECT 80.185 -100.905 80.775 -100.720 ;
        RECT 82.005 -100.905 82.595 -100.720 ;
        RECT 77.820 -100.975 78.050 -100.920 ;
        RECT 77.140 -101.935 78.050 -100.975 ;
        RECT 73.705 -102.835 74.295 -102.720 ;
        RECT 75.525 -102.835 76.115 -102.720 ;
        RECT 71.885 -103.665 72.475 -103.415 ;
        RECT 73.705 -103.665 74.295 -103.415 ;
        RECT 69.960 -106.860 71.000 -104.310 ;
        RECT 71.885 -105.480 74.295 -103.665 ;
        RECT 71.885 -105.520 72.475 -105.480 ;
        RECT 73.705 -105.520 74.295 -105.480 ;
        RECT 75.525 -103.685 76.115 -103.415 ;
        RECT 75.525 -105.520 76.175 -103.685 ;
        RECT 75.550 -106.710 76.175 -105.520 ;
        RECT 69.960 -106.900 70.190 -106.860 ;
        RECT 69.665 -107.585 70.010 -107.095 ;
        RECT 63.580 -108.810 64.170 -108.725 ;
        RECT 65.400 -108.810 65.990 -108.725 ;
        RECT 67.220 -108.810 67.810 -108.685 ;
        RECT 69.665 -108.915 70.010 -108.585 ;
        RECT 69.645 -109.130 70.010 -108.915 ;
        RECT 69.645 -109.145 69.935 -109.130 ;
        RECT 69.455 -109.380 69.685 -109.305 ;
        RECT 61.655 -111.195 62.780 -109.440 ;
        RECT 63.580 -109.485 64.170 -109.390 ;
        RECT 61.655 -111.260 62.695 -111.195 ;
        RECT 61.655 -111.315 61.885 -111.260 ;
        RECT 61.405 -111.490 61.695 -111.475 ;
        RECT 61.405 -111.705 61.745 -111.490 ;
        RECT 63.565 -111.495 64.170 -109.485 ;
        RECT 65.400 -109.610 65.990 -109.390 ;
        RECT 67.220 -109.610 67.810 -109.390 ;
        RECT 65.375 -111.425 67.810 -109.610 ;
        RECT 69.125 -109.875 69.685 -109.380 ;
        RECT 65.400 -111.495 65.990 -111.425 ;
        RECT 67.220 -111.495 67.810 -111.425 ;
        RECT 68.695 -111.280 69.685 -109.875 ;
        RECT 63.565 -111.515 64.110 -111.495 ;
        RECT 61.430 -111.780 61.745 -111.705 ;
        RECT 68.695 -112.015 69.155 -111.280 ;
        RECT 69.455 -111.305 69.685 -111.280 ;
        RECT 69.895 -109.405 70.125 -109.305 ;
        RECT 70.625 -109.405 71.000 -106.860 ;
        RECT 71.885 -106.910 72.475 -106.710 ;
        RECT 73.705 -106.910 74.295 -106.710 ;
        RECT 71.885 -108.725 74.295 -106.910 ;
        RECT 71.885 -108.815 72.475 -108.725 ;
        RECT 73.705 -108.815 74.295 -108.725 ;
        RECT 75.525 -108.705 76.175 -106.710 ;
        RECT 77.390 -106.850 78.050 -101.935 ;
        RECT 77.820 -106.920 78.050 -106.850 ;
        RECT 78.260 -100.940 78.490 -100.920 ;
        RECT 78.260 -103.525 79.045 -100.940 ;
        RECT 80.185 -102.720 82.595 -100.905 ;
        RECT 80.185 -102.825 80.775 -102.720 ;
        RECT 82.005 -102.825 82.595 -102.720 ;
        RECT 80.185 -103.525 80.775 -103.405 ;
        RECT 78.260 -105.340 80.775 -103.525 ;
        RECT 82.005 -103.645 82.595 -103.405 ;
        RECT 78.260 -106.105 79.045 -105.340 ;
        RECT 80.185 -105.510 80.775 -105.340 ;
        RECT 81.940 -105.510 82.595 -103.645 ;
        RECT 78.260 -106.840 79.085 -106.105 ;
        RECT 78.260 -106.920 78.490 -106.840 ;
        RECT 78.010 -107.180 78.300 -107.125 ;
        RECT 78.010 -107.190 78.525 -107.180 ;
        RECT 77.980 -107.625 78.525 -107.190 ;
        RECT 78.755 -107.420 79.085 -106.840 ;
        RECT 81.940 -106.700 82.565 -105.510 ;
        RECT 78.825 -108.420 79.085 -107.420 ;
        RECT 75.525 -108.815 76.115 -108.705 ;
        RECT 77.980 -109.090 78.525 -108.625 ;
        RECT 78.800 -108.715 79.085 -108.420 ;
        RECT 80.115 -108.675 80.830 -106.990 ;
        RECT 81.940 -108.665 82.595 -106.700 ;
        RECT 77.980 -109.100 78.455 -109.090 ;
        RECT 78.010 -109.115 78.455 -109.100 ;
        RECT 78.010 -109.145 78.300 -109.115 ;
        RECT 77.820 -109.350 78.050 -109.305 ;
        RECT 69.895 -111.095 71.000 -109.405 ;
        RECT 71.885 -109.505 72.475 -109.395 ;
        RECT 69.895 -111.225 70.960 -111.095 ;
        RECT 69.895 -111.305 70.125 -111.225 ;
        RECT 69.705 -111.465 70.020 -111.455 ;
        RECT 69.645 -111.695 70.020 -111.465 ;
        RECT 71.870 -111.500 72.475 -109.505 ;
        RECT 73.705 -109.550 74.295 -109.395 ;
        RECT 75.525 -109.550 76.115 -109.395 ;
        RECT 73.705 -111.365 76.115 -109.550 ;
        RECT 77.470 -109.785 78.050 -109.350 ;
        RECT 73.705 -111.500 74.295 -111.365 ;
        RECT 71.870 -111.525 72.415 -111.500 ;
        RECT 74.640 -111.515 75.185 -111.365 ;
        RECT 75.525 -111.500 76.115 -111.365 ;
        RECT 77.050 -111.250 78.050 -109.785 ;
        RECT 69.705 -111.745 70.020 -111.695 ;
        RECT 77.050 -112.015 77.510 -111.250 ;
        RECT 77.820 -111.305 78.050 -111.250 ;
        RECT 78.260 -109.365 78.490 -109.305 ;
        RECT 78.755 -109.365 79.085 -108.715 ;
        RECT 80.185 -108.710 80.790 -108.675 ;
        RECT 80.185 -108.805 80.775 -108.710 ;
        RECT 82.005 -108.805 82.595 -108.665 ;
        RECT 78.260 -110.860 79.085 -109.365 ;
        RECT 80.185 -109.570 80.775 -109.385 ;
        RECT 82.005 -109.570 82.595 -109.385 ;
        RECT 78.260 -111.245 78.860 -110.860 ;
        RECT 78.260 -111.305 78.490 -111.245 ;
        RECT 80.185 -111.385 82.595 -109.570 ;
        RECT 77.985 -111.755 78.300 -111.465 ;
        RECT 80.185 -111.490 80.775 -111.385 ;
        RECT 82.005 -111.490 82.595 -111.385 ;
        RECT 14.685 -112.495 42.730 -112.015 ;
        RECT 14.675 -112.975 42.730 -112.495 ;
        RECT 43.730 -112.495 83.300 -112.015 ;
        RECT 43.730 -112.975 83.305 -112.495 ;
        RECT 14.675 -113.075 83.305 -112.975 ;
      LAYER met2 ;
        RECT 21.820 -110.215 33.365 -109.625 ;
        RECT 80.245 -109.740 80.790 -107.740 ;
        RECT 38.410 -109.790 39.060 -109.770 ;
        RECT 38.410 -110.335 50.350 -109.790 ;
        RECT 38.410 -110.405 39.060 -110.335 ;
        RECT 55.270 -110.340 66.920 -109.795 ;
        RECT 71.840 -110.285 80.790 -109.740 ;
        RECT 24.490 -110.970 25.085 -110.530 ;
        RECT 17.170 -111.565 25.085 -110.970 ;
        RECT 30.150 -111.270 41.720 -110.680 ;
        RECT 46.890 -111.480 58.500 -110.890 ;
        RECT 63.535 -111.485 75.215 -110.940 ;
  END
END r2r_dac
END LIBRARY

