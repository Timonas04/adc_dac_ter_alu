MACRO digital
  CLASS BLOCK ;
  FOREIGN digital ;
  ORIGIN 0.000 0.000 ;
  SIZE 82.350 BY 93.070 ;
  PIN DAC6_conn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 27.240 82.350 27.840 ;
    END
  END DAC6_conn
  PIN DAC8_conn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 30.640 82.350 31.240 ;
    END
  END DAC8_conn
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 81.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 81.840 ;
    END
  END VPWR
  PIN a0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 54.440 82.350 55.040 ;
    END
  END a0
  PIN a0_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 92.570 29.350 93.070 ;
    END
  END a0_sel
  PIN aux1_conn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 34.040 82.350 34.640 ;
    END
  END aux1_conn
  PIN aux2_conn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 16.190 92.570 16.470 93.070 ;
    END
  END aux2_conn
  PIN buffi_conn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 0.090 92.570 0.370 93.070 ;
    END
  END buffi_conn
  PIN buffo_conn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 37.440 82.350 38.040 ;
    END
  END buffo_conn
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 81.850 51.040 82.350 51.640 ;
    END
  END clk
  PIN compr1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 92.570 10.030 93.070 ;
    END
  END compr1
  PIN compr2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 92.570 22.910 93.070 ;
    END
  END compr2
  PIN flash_adc_inp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 68.040 82.350 68.640 ;
    END
  END flash_adc_inp[0]
  PIN flash_adc_inp[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 92.570 61.550 93.070 ;
    END
  END flash_adc_inp[10]
  PIN flash_adc_inp[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 92.570 58.330 93.070 ;
    END
  END flash_adc_inp[11]
  PIN flash_adc_inp[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 92.570 55.110 93.070 ;
    END
  END flash_adc_inp[12]
  PIN flash_adc_inp[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.710 92.570 67.990 93.070 ;
    END
  END flash_adc_inp[13]
  PIN flash_adc_inp[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 92.570 71.210 93.070 ;
    END
  END flash_adc_inp[14]
  PIN flash_adc_inp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 81.850 91.840 82.350 92.440 ;
    END
  END flash_adc_inp[1]
  PIN flash_adc_inp[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 71.440 82.350 72.040 ;
    END
  END flash_adc_inp[2]
  PIN flash_adc_inp[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 88.440 82.350 89.040 ;
    END
  END flash_adc_inp[3]
  PIN flash_adc_inp[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 74.840 82.350 75.440 ;
    END
  END flash_adc_inp[4]
  PIN flash_adc_inp[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 81.850 85.040 82.350 85.640 ;
    END
  END flash_adc_inp[5]
  PIN flash_adc_inp[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 81.850 81.640 82.350 82.240 ;
    END
  END flash_adc_inp[6]
  PIN flash_adc_inp[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 92.570 77.650 93.070 ;
    END
  END flash_adc_inp[7]
  PIN flash_adc_inp[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 92.570 80.870 93.070 ;
    END
  END flash_adc_inp[8]
  PIN flash_adc_inp[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 92.570 64.770 93.070 ;
    END
  END flash_adc_inp[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 92.570 74.430 93.070 ;
    END
  END rst_n
  PIN tern_dac[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 0.500 21.040 ;
    END
  END tern_dac[0]
  PIN tern_dac[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 40.840 82.350 41.440 ;
    END
  END tern_dac[10]
  PIN tern_dac[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 44.240 82.350 44.840 ;
    END
  END tern_dac[11]
  PIN tern_dac[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 92.570 39.010 93.070 ;
    END
  END tern_dac[12]
  PIN tern_dac[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 92.570 6.810 93.070 ;
    END
  END tern_dac[13]
  PIN tern_dac[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 92.570 42.230 93.070 ;
    END
  END tern_dac[14]
  PIN tern_dac[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 92.570 19.690 93.070 ;
    END
  END tern_dac[15]
  PIN tern_dac[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 0.500 ;
    END
  END tern_dac[16]
  PIN tern_dac[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 81.850 13.640 82.350 14.240 ;
    END
  END tern_dac[17]
  PIN tern_dac[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 0.500 58.440 ;
    END
  END tern_dac[1]
  PIN tern_dac[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 0.500 61.840 ;
    END
  END tern_dac[2]
  PIN tern_dac[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 0.500 31.240 ;
    END
  END tern_dac[3]
  PIN tern_dac[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 0.500 ;
    END
  END tern_dac[4]
  PIN tern_dac[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 0.500 68.640 ;
    END
  END tern_dac[5]
  PIN tern_dac[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 0.500 82.240 ;
    END
  END tern_dac[6]
  PIN tern_dac[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 47.640 82.350 48.240 ;
    END
  END tern_dac[7]
  PIN tern_dac[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 0.500 72.040 ;
    END
  END tern_dac[8]
  PIN tern_dac[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 92.570 51.890 93.070 ;
    END
  END tern_dac[9]
  PIN ternff_conn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 57.840 82.350 58.440 ;
    END
  END ternff_conn
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 0.500 24.440 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 0.500 27.840 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 0.500 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 0.500 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 0.500 55.040 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 0.500 65.240 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 92.570 48.670 93.070 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 92.570 45.450 93.070 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3.310 92.570 3.590 93.070 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 92.570 13.250 93.070 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 0.500 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 0.500 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.500 48.240 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 23.840 82.350 24.440 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 81.850 17.040 82.350 17.640 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 81.850 20.440 82.350 21.040 ;
    END
  END uio_in[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 25.850 92.570 26.130 93.070 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 35.510 92.570 35.790 93.070 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 92.570 32.570 93.070 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 0.500 78.840 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 0.500 75.440 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 78.240 82.350 78.840 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 64.640 82.350 65.240 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 81.850 61.240 82.350 61.840 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 5.665 81.495 5.835 81.685 ;
        RECT 8.425 81.495 8.595 81.685 ;
        RECT 10.265 81.495 10.435 81.685 ;
        RECT 10.725 81.495 10.895 81.685 ;
        RECT 13.945 81.495 14.115 81.685 ;
        RECT 15.785 81.495 15.955 81.685 ;
        RECT 18.085 81.515 18.255 81.685 ;
        RECT 18.085 81.495 18.250 81.515 ;
        RECT 20.385 81.495 20.555 81.685 ;
        RECT 20.845 81.515 21.015 81.685 ;
        RECT 20.865 81.495 21.015 81.515 ;
        RECT 24.980 81.495 25.150 81.685 ;
        RECT 25.445 81.515 25.615 81.685 ;
        RECT 25.475 81.495 25.615 81.515 ;
        RECT 28.210 81.495 28.380 81.685 ;
        RECT 31.895 81.540 32.055 81.650 ;
        RECT 41.545 81.495 41.715 81.685 ;
        RECT 42.925 81.495 43.095 81.685 ;
        RECT 43.395 81.540 43.555 81.650 ;
        RECT 47.520 81.495 47.690 81.685 ;
        RECT 56.725 81.495 56.895 81.685 ;
        RECT 57.645 81.495 57.815 81.685 ;
        RECT 60.865 81.495 61.035 81.685 ;
        RECT 73.280 81.495 73.450 81.685 ;
        RECT 73.745 81.495 73.915 81.685 ;
        RECT 76.505 81.495 76.675 81.685 ;
        RECT 5.525 80.685 6.895 81.495 ;
        RECT 6.905 80.815 8.735 81.495 ;
        RECT 8.745 80.815 10.575 81.495 ;
        RECT 10.585 80.815 12.415 81.495 ;
        RECT 12.425 80.815 14.255 81.495 ;
        RECT 14.265 80.815 16.095 81.495 ;
        RECT 16.415 80.815 18.250 81.495 ;
        RECT 6.905 80.585 8.250 80.815 ;
        RECT 8.745 80.585 10.090 80.815 ;
        RECT 12.425 80.585 13.770 80.815 ;
        RECT 14.265 80.585 15.610 80.815 ;
        RECT 16.415 80.585 17.345 80.815 ;
        RECT 18.415 80.625 18.845 81.410 ;
        RECT 18.865 80.815 20.695 81.495 ;
        RECT 18.865 80.585 20.210 80.815 ;
        RECT 20.865 80.675 22.795 81.495 ;
        RECT 21.845 80.585 22.795 80.675 ;
        RECT 23.105 80.585 25.295 81.495 ;
        RECT 25.475 80.675 28.045 81.495 ;
        RECT 26.455 80.585 28.045 80.675 ;
        RECT 28.065 80.585 30.985 81.495 ;
        RECT 31.295 80.625 31.725 81.410 ;
        RECT 32.750 80.815 41.855 81.495 ;
        RECT 41.865 80.715 43.235 81.495 ;
        RECT 44.175 80.625 44.605 81.410 ;
        RECT 44.915 80.585 47.835 81.495 ;
        RECT 47.930 80.815 57.035 81.495 ;
        RECT 57.505 81.465 59.345 81.495 ;
        RECT 57.055 80.625 57.485 81.410 ;
        RECT 57.505 80.815 60.670 81.465 ;
        RECT 60.725 80.815 69.830 81.495 ;
        RECT 57.990 80.785 60.670 80.815 ;
        RECT 57.990 80.585 59.345 80.785 ;
        RECT 69.935 80.625 70.365 81.410 ;
        RECT 70.395 81.265 73.450 81.495 ;
        RECT 70.395 80.585 73.595 81.265 ;
        RECT 73.605 80.815 75.435 81.495 ;
        RECT 74.090 80.585 75.435 80.815 ;
        RECT 75.445 80.685 76.815 81.495 ;
      LAYER nwell ;
        RECT 5.330 77.465 77.010 80.295 ;
      LAYER pwell ;
        RECT 8.025 77.085 8.975 77.175 ;
        RECT 5.525 76.265 6.895 77.075 ;
        RECT 8.025 76.265 9.955 77.085 ;
        RECT 11.065 76.265 12.415 77.175 ;
        RECT 12.445 76.265 13.795 77.175 ;
        RECT 16.550 76.975 17.935 77.175 ;
        RECT 14.265 76.295 17.935 76.975 ;
        RECT 18.415 76.350 18.845 77.135 ;
        RECT 5.665 76.055 5.835 76.265 ;
        RECT 9.805 76.245 9.955 76.265 ;
        RECT 7.055 76.110 7.215 76.220 ;
        RECT 9.805 76.075 9.975 76.245 ;
        RECT 10.275 76.110 10.435 76.220 ;
        RECT 11.180 76.075 11.350 76.265 ;
        RECT 12.100 76.055 12.270 76.245 ;
        RECT 12.560 76.210 12.730 76.265 ;
        RECT 12.560 76.100 12.735 76.210 ;
        RECT 13.940 76.105 14.060 76.215 ;
        RECT 12.560 76.075 12.730 76.100 ;
        RECT 14.405 76.075 14.575 76.295 ;
        RECT 16.565 76.265 17.935 76.295 ;
        RECT 19.325 76.265 22.995 77.175 ;
        RECT 23.005 76.945 24.595 77.175 ;
        RECT 23.005 76.265 26.675 76.945 ;
        RECT 26.770 76.265 35.875 76.945 ;
        RECT 35.885 76.265 39.985 77.175 ;
        RECT 40.025 76.265 43.695 77.175 ;
        RECT 44.175 76.350 44.605 77.135 ;
        RECT 48.045 76.945 51.975 77.175 ;
        RECT 44.635 76.265 47.375 76.945 ;
        RECT 47.560 76.265 51.975 76.945 ;
        RECT 51.985 76.265 55.100 77.175 ;
        RECT 55.205 76.265 56.575 77.075 ;
        RECT 56.595 76.265 57.945 77.175 ;
        RECT 57.965 76.265 61.175 77.175 ;
        RECT 61.185 76.945 64.010 77.175 ;
        RECT 65.710 76.945 68.535 77.175 ;
        RECT 61.185 76.265 64.715 76.945 ;
        RECT 5.525 75.245 6.895 76.055 ;
        RECT 7.285 75.145 12.415 76.055 ;
        RECT 13.345 76.025 14.740 76.055 ;
        RECT 15.785 76.025 15.955 76.245 ;
        RECT 16.250 76.055 16.420 76.245 ;
        RECT 18.080 76.105 18.200 76.215 ;
        RECT 19.000 76.105 19.120 76.215 ;
        RECT 19.470 76.075 19.640 76.265 ;
        RECT 20.845 76.095 21.015 76.245 ;
        RECT 13.345 75.345 16.080 76.025 ;
        RECT 13.345 75.145 14.755 75.345 ;
        RECT 16.105 75.145 19.975 76.055 ;
        RECT 20.245 75.145 21.135 76.095 ;
        RECT 21.315 76.055 21.485 76.245 ;
        RECT 22.690 76.055 22.860 76.245 ;
        RECT 26.360 76.075 26.530 76.265 ;
        RECT 26.825 76.055 26.995 76.245 ;
        RECT 27.260 76.055 27.430 76.245 ;
        RECT 31.885 76.095 32.055 76.245 ;
        RECT 21.165 75.275 22.535 76.055 ;
        RECT 22.545 75.145 23.895 76.055 ;
        RECT 23.925 75.375 27.135 76.055 ;
        RECT 23.925 75.145 25.060 75.375 ;
        RECT 27.200 75.145 31.275 76.055 ;
        RECT 31.295 75.185 31.725 75.970 ;
        RECT 31.765 75.145 32.655 76.095 ;
        RECT 32.805 76.055 32.975 76.245 ;
        RECT 35.565 76.075 35.735 76.265 ;
        RECT 36.030 76.075 36.200 76.265 ;
        RECT 43.380 76.075 43.550 76.265 ;
        RECT 43.840 76.105 43.960 76.215 ;
        RECT 47.065 76.075 47.235 76.265 ;
        RECT 47.560 76.245 47.670 76.265 ;
        RECT 47.500 76.075 47.670 76.245 ;
        RECT 50.745 76.055 50.915 76.245 ;
        RECT 51.205 76.055 51.375 76.245 ;
        RECT 52.130 76.075 52.300 76.265 ;
        RECT 53.050 76.055 53.220 76.245 ;
        RECT 55.345 76.075 55.515 76.265 ;
        RECT 56.720 76.105 56.840 76.215 ;
        RECT 57.645 76.055 57.815 76.265 ;
        RECT 58.110 76.075 58.280 76.265 ;
        RECT 64.515 76.245 64.715 76.265 ;
        RECT 64.545 76.075 64.715 76.245 ;
        RECT 65.005 76.265 68.535 76.945 ;
        RECT 68.545 76.265 69.915 77.045 ;
        RECT 69.935 76.350 70.365 77.135 ;
        RECT 71.230 76.945 74.055 77.175 ;
        RECT 70.525 76.265 74.055 76.945 ;
        RECT 74.065 76.265 75.435 77.045 ;
        RECT 75.445 76.265 76.815 77.075 ;
        RECT 65.005 76.245 65.205 76.265 ;
        RECT 65.005 76.075 65.175 76.245 ;
        RECT 66.845 76.075 67.015 76.245 ;
        RECT 68.685 76.075 68.855 76.265 ;
        RECT 70.525 76.245 70.725 76.265 ;
        RECT 70.525 76.075 70.695 76.245 ;
        RECT 66.845 76.055 67.045 76.075 ;
        RECT 70.525 76.055 70.725 76.075 ;
        RECT 74.205 76.055 74.375 76.245 ;
        RECT 75.115 76.075 75.285 76.265 ;
        RECT 76.505 76.055 76.675 76.265 ;
        RECT 32.665 75.375 41.770 76.055 ;
        RECT 41.950 75.375 51.055 76.055 ;
        RECT 51.065 75.375 52.895 76.055 ;
        RECT 51.550 75.145 52.895 75.375 ;
        RECT 52.905 75.145 56.505 76.055 ;
        RECT 57.055 75.185 57.485 75.970 ;
        RECT 57.505 75.375 66.610 76.055 ;
        RECT 66.845 75.375 70.375 76.055 ;
        RECT 70.525 75.375 74.055 76.055 ;
        RECT 67.550 75.145 70.375 75.375 ;
        RECT 71.230 75.145 74.055 75.375 ;
        RECT 74.075 75.145 75.425 76.055 ;
        RECT 75.445 75.245 76.815 76.055 ;
      LAYER nwell ;
        RECT 5.330 72.025 77.010 74.855 ;
      LAYER pwell ;
        RECT 5.525 70.825 6.895 71.635 ;
        RECT 7.365 71.505 8.710 71.735 ;
        RECT 10.345 71.645 11.295 71.735 ;
        RECT 7.365 70.825 9.195 71.505 ;
        RECT 9.365 70.825 11.295 71.645 ;
        RECT 11.960 71.055 13.795 71.735 ;
        RECT 14.115 71.505 15.045 71.735 ;
        RECT 11.960 70.825 13.650 71.055 ;
        RECT 14.115 70.825 15.950 71.505 ;
        RECT 16.105 70.825 18.395 71.735 ;
        RECT 18.415 70.910 18.845 71.695 ;
        RECT 23.235 71.645 24.825 71.735 ;
        RECT 19.335 70.825 22.075 71.505 ;
        RECT 22.255 70.825 24.825 71.645 ;
        RECT 24.845 70.825 33.950 71.505 ;
        RECT 34.055 70.825 35.405 71.735 ;
        RECT 35.425 70.825 36.775 71.735 ;
        RECT 36.805 70.825 38.175 71.605 ;
        RECT 38.185 70.825 39.555 71.605 ;
        RECT 39.565 70.825 40.935 71.605 ;
        RECT 40.945 70.825 43.695 71.635 ;
        RECT 44.175 70.910 44.605 71.695 ;
        RECT 44.625 70.825 48.755 71.735 ;
        RECT 48.785 70.825 50.135 71.735 ;
        RECT 50.145 70.825 59.250 71.505 ;
        RECT 59.345 70.825 68.450 71.505 ;
        RECT 68.555 70.825 69.905 71.735 ;
        RECT 69.935 70.910 70.365 71.695 ;
        RECT 71.230 71.505 74.055 71.735 ;
        RECT 70.525 70.825 74.055 71.505 ;
        RECT 5.665 70.615 5.835 70.825 ;
        RECT 7.040 70.665 7.160 70.775 ;
        RECT 8.885 70.635 9.055 70.825 ;
        RECT 9.365 70.805 9.515 70.825 ;
        RECT 9.345 70.635 9.515 70.805 ;
        RECT 9.805 70.635 9.975 70.805 ;
        RECT 10.265 70.635 10.435 70.805 ;
        RECT 13.480 70.635 13.650 70.825 ;
        RECT 15.785 70.805 15.950 70.825 ;
        RECT 15.780 70.635 15.955 70.805 ;
        RECT 9.805 70.615 9.945 70.635 ;
        RECT 5.525 69.805 6.895 70.615 ;
        RECT 7.375 69.795 9.945 70.615 ;
        RECT 10.270 70.615 10.435 70.635 ;
        RECT 15.780 70.615 15.950 70.635 ;
        RECT 16.245 70.615 16.415 70.805 ;
        RECT 18.080 70.635 18.250 70.825 ;
        RECT 19.000 70.665 19.120 70.775 ;
        RECT 19.930 70.615 20.100 70.805 ;
        RECT 21.765 70.635 21.935 70.825 ;
        RECT 22.255 70.805 22.395 70.825 ;
        RECT 22.225 70.635 22.395 70.805 ;
        RECT 23.145 70.615 23.315 70.805 ;
        RECT 24.985 70.635 25.155 70.825 ;
        RECT 26.365 70.615 26.535 70.805 ;
        RECT 26.830 70.615 27.000 70.805 ;
        RECT 30.965 70.615 31.135 70.805 ;
        RECT 10.270 69.935 12.105 70.615 ;
        RECT 7.375 69.705 8.965 69.795 ;
        RECT 11.175 69.705 12.105 69.935 ;
        RECT 12.425 69.705 16.095 70.615 ;
        RECT 16.105 69.705 18.855 70.615 ;
        RECT 18.865 69.705 20.215 70.615 ;
        RECT 20.245 69.705 23.455 70.615 ;
        RECT 23.465 69.705 26.675 70.615 ;
        RECT 26.685 69.705 28.515 70.615 ;
        RECT 28.535 69.935 31.275 70.615 ;
        RECT 31.295 69.745 31.725 70.530 ;
        RECT 31.885 70.385 32.055 70.805 ;
        RECT 34.185 70.635 34.355 70.825 ;
        RECT 36.490 70.635 36.660 70.825 ;
        RECT 37.410 70.615 37.580 70.805 ;
        RECT 37.865 70.635 38.035 70.825 ;
        RECT 39.235 70.635 39.405 70.825 ;
        RECT 40.615 70.635 40.785 70.825 ;
        RECT 41.085 70.615 41.255 70.825 ;
        RECT 43.840 70.665 43.960 70.775 ;
        RECT 46.605 70.615 46.775 70.805 ;
        RECT 48.440 70.635 48.610 70.825 ;
        RECT 49.820 70.635 49.990 70.825 ;
        RECT 50.285 70.635 50.455 70.825 ;
        RECT 53.040 70.615 53.210 70.805 ;
        RECT 53.510 70.635 53.680 70.805 ;
        RECT 56.720 70.665 56.840 70.775 ;
        RECT 53.535 70.615 53.680 70.635 ;
        RECT 57.645 70.615 57.815 70.805 ;
        RECT 59.485 70.635 59.655 70.825 ;
        RECT 66.850 70.615 67.020 70.805 ;
        RECT 68.685 70.635 68.855 70.825 ;
        RECT 70.525 70.805 70.725 70.825 ;
        RECT 70.525 70.635 70.700 70.805 ;
        RECT 74.065 70.785 74.955 71.735 ;
        RECT 75.445 70.825 76.815 71.635 ;
        RECT 74.665 70.635 74.835 70.785 ;
        RECT 75.130 70.775 75.300 70.805 ;
        RECT 75.120 70.665 75.300 70.775 ;
        RECT 70.530 70.615 70.700 70.635 ;
        RECT 75.130 70.615 75.300 70.665 ;
        RECT 76.505 70.615 76.675 70.825 ;
        RECT 33.165 70.385 37.255 70.615 ;
        RECT 31.780 69.705 37.255 70.385 ;
        RECT 37.265 69.705 40.920 70.615 ;
        RECT 40.945 69.805 46.455 70.615 ;
        RECT 46.465 69.805 49.215 70.615 ;
        RECT 49.225 69.705 53.355 70.615 ;
        RECT 53.535 69.705 56.575 70.615 ;
        RECT 57.055 69.745 57.485 70.530 ;
        RECT 57.505 69.935 66.610 70.615 ;
        RECT 66.705 69.705 70.250 70.615 ;
        RECT 70.385 69.705 73.930 70.615 ;
        RECT 74.065 69.705 75.415 70.615 ;
        RECT 75.445 69.805 76.815 70.615 ;
      LAYER nwell ;
        RECT 5.330 66.585 77.010 69.415 ;
      LAYER pwell ;
        RECT 5.525 65.385 6.895 66.195 ;
        RECT 8.310 66.065 9.655 66.295 ;
        RECT 7.825 65.385 9.655 66.065 ;
        RECT 9.665 66.065 11.010 66.295 ;
        RECT 9.665 65.385 11.495 66.065 ;
        RECT 11.505 65.385 15.175 66.295 ;
        RECT 15.195 65.385 17.925 66.295 ;
        RECT 18.415 65.470 18.845 66.255 ;
        RECT 18.880 65.385 20.695 66.295 ;
        RECT 20.705 66.065 22.050 66.295 ;
        RECT 20.705 65.385 22.535 66.065 ;
        RECT 22.695 65.385 26.350 66.295 ;
        RECT 27.690 65.385 36.795 66.065 ;
        RECT 36.805 65.385 40.935 66.295 ;
        RECT 40.945 65.385 44.155 66.295 ;
        RECT 44.175 65.470 44.605 66.255 ;
        RECT 44.710 65.385 53.815 66.065 ;
        RECT 53.825 65.385 57.495 66.295 ;
        RECT 57.505 65.385 60.715 66.295 ;
        RECT 60.810 65.385 69.915 66.065 ;
        RECT 69.935 65.470 70.365 66.255 ;
        RECT 70.385 65.385 73.595 66.295 ;
        RECT 73.605 65.385 75.420 66.295 ;
        RECT 75.445 65.385 76.815 66.195 ;
        RECT 5.665 65.175 5.835 65.385 ;
        RECT 7.055 65.230 7.215 65.340 ;
        RECT 7.965 65.195 8.135 65.385 ;
        RECT 8.425 65.175 8.595 65.365 ;
        RECT 8.880 65.225 9.000 65.335 ;
        RECT 9.355 65.175 9.525 65.365 ;
        RECT 11.185 65.195 11.355 65.385 ;
        RECT 11.650 65.365 11.820 65.385 ;
        RECT 11.645 65.195 11.820 65.365 ;
        RECT 12.105 65.195 12.275 65.365 ;
        RECT 14.415 65.220 14.575 65.330 ;
        RECT 15.325 65.195 15.495 65.385 ;
        RECT 11.645 65.175 11.815 65.195 ;
        RECT 12.110 65.175 12.275 65.195 ;
        RECT 16.245 65.175 16.415 65.365 ;
        RECT 17.165 65.215 17.335 65.365 ;
        RECT 5.525 64.365 6.895 65.175 ;
        RECT 6.905 64.495 8.735 65.175 ;
        RECT 6.905 64.265 8.250 64.495 ;
        RECT 9.205 64.395 10.575 65.175 ;
        RECT 10.595 64.265 11.945 65.175 ;
        RECT 12.110 64.495 13.945 65.175 ;
        RECT 13.015 64.265 13.945 64.495 ;
        RECT 15.195 64.265 16.545 65.175 ;
        RECT 16.565 64.265 17.455 65.215 ;
        RECT 17.635 65.175 17.805 65.365 ;
        RECT 18.080 65.225 18.200 65.335 ;
        RECT 19.005 65.195 19.175 65.385 ;
        RECT 20.385 65.175 20.555 65.365 ;
        RECT 21.305 65.215 21.475 65.365 ;
        RECT 17.485 64.395 18.855 65.175 ;
        RECT 18.865 64.265 20.680 65.175 ;
        RECT 20.705 64.265 21.595 65.215 ;
        RECT 21.775 65.175 21.945 65.365 ;
        RECT 22.225 65.195 22.395 65.385 ;
        RECT 22.695 65.365 22.855 65.385 ;
        RECT 22.685 65.195 22.855 65.365 ;
        RECT 24.065 65.175 24.235 65.365 ;
        RECT 24.535 65.175 24.705 65.365 ;
        RECT 25.905 65.175 26.075 65.365 ;
        RECT 26.835 65.230 26.995 65.340 ;
        RECT 28.665 65.175 28.835 65.365 ;
        RECT 31.880 65.225 32.000 65.335 ;
        RECT 32.345 65.175 32.515 65.365 ;
        RECT 36.485 65.195 36.655 65.385 ;
        RECT 36.950 65.195 37.120 65.385 ;
        RECT 38.325 65.175 38.495 65.365 ;
        RECT 43.845 65.195 44.015 65.385 ;
        RECT 47.525 65.175 47.695 65.365 ;
        RECT 53.505 65.195 53.675 65.385 ;
        RECT 56.725 65.175 56.895 65.365 ;
        RECT 57.180 65.195 57.350 65.385 ;
        RECT 57.650 65.175 57.820 65.365 ;
        RECT 60.400 65.195 60.570 65.385 ;
        RECT 61.330 65.175 61.500 65.365 ;
        RECT 65.475 65.220 65.635 65.330 ;
        RECT 66.385 65.175 66.555 65.365 ;
        RECT 69.605 65.195 69.775 65.385 ;
        RECT 70.530 65.195 70.700 65.385 ;
        RECT 75.125 65.195 75.295 65.385 ;
        RECT 76.505 65.175 76.675 65.385 ;
        RECT 21.625 64.395 22.995 65.175 ;
        RECT 23.005 64.395 24.375 65.175 ;
        RECT 24.385 64.395 25.755 65.175 ;
        RECT 25.775 64.265 28.505 65.175 ;
        RECT 28.525 64.495 31.275 65.175 ;
        RECT 30.345 64.265 31.275 64.495 ;
        RECT 31.295 64.305 31.725 65.090 ;
        RECT 32.205 64.265 35.415 65.175 ;
        RECT 35.425 64.265 38.635 65.175 ;
        RECT 38.730 64.495 47.835 65.175 ;
        RECT 47.930 64.495 57.035 65.175 ;
        RECT 57.055 64.305 57.485 65.090 ;
        RECT 57.505 64.265 61.175 65.175 ;
        RECT 61.185 64.265 65.315 65.175 ;
        RECT 66.245 64.495 75.350 65.175 ;
        RECT 75.445 64.365 76.815 65.175 ;
      LAYER nwell ;
        RECT 5.330 61.145 77.010 63.975 ;
      LAYER pwell ;
        RECT 5.525 59.945 6.895 60.755 ;
        RECT 7.825 59.945 9.195 60.725 ;
        RECT 9.205 59.945 10.575 60.725 ;
        RECT 10.585 59.945 11.955 60.725 ;
        RECT 11.965 59.945 13.335 60.725 ;
        RECT 14.395 60.625 15.325 60.855 ;
        RECT 13.490 59.945 15.325 60.625 ;
        RECT 15.645 60.625 16.990 60.855 ;
        RECT 15.645 59.945 17.475 60.625 ;
        RECT 18.415 60.030 18.845 60.815 ;
        RECT 19.785 60.625 20.715 60.855 ;
        RECT 26.425 60.765 27.375 60.855 ;
        RECT 19.785 59.945 23.685 60.625 ;
        RECT 24.845 59.945 26.215 60.725 ;
        RECT 26.425 59.945 28.355 60.765 ;
        RECT 28.525 59.945 29.875 60.855 ;
        RECT 29.905 59.945 33.115 60.855 ;
        RECT 33.125 59.945 34.475 60.855 ;
        RECT 35.050 59.945 44.155 60.625 ;
        RECT 44.175 60.030 44.605 60.815 ;
        RECT 44.725 59.945 46.915 60.855 ;
        RECT 46.925 59.945 51.000 60.855 ;
        RECT 51.150 59.945 60.255 60.625 ;
        RECT 60.350 59.945 69.455 60.625 ;
        RECT 69.935 60.030 70.365 60.815 ;
        RECT 70.385 59.945 73.425 60.855 ;
        RECT 73.605 59.945 75.435 60.625 ;
        RECT 75.445 59.945 76.815 60.755 ;
        RECT 5.665 59.735 5.835 59.945 ;
        RECT 8.885 59.925 9.055 59.945 ;
        RECT 7.055 59.790 7.215 59.900 ;
        RECT 8.425 59.735 8.595 59.925 ;
        RECT 8.880 59.755 9.055 59.925 ;
        RECT 10.265 59.755 10.435 59.945 ;
        RECT 11.645 59.755 11.815 59.945 ;
        RECT 8.880 59.735 9.050 59.755 ;
        RECT 13.025 59.735 13.195 59.945 ;
        RECT 13.490 59.925 13.655 59.945 ;
        RECT 13.485 59.755 13.655 59.925 ;
        RECT 14.410 59.735 14.580 59.925 ;
        RECT 17.165 59.755 17.335 59.945 ;
        RECT 17.635 59.790 17.795 59.900 ;
        RECT 18.085 59.755 18.255 59.925 ;
        RECT 19.015 59.790 19.175 59.900 ;
        RECT 19.470 59.735 19.640 59.925 ;
        RECT 20.200 59.755 20.370 59.945 ;
        RECT 21.120 59.735 21.290 59.925 ;
        RECT 24.075 59.790 24.235 59.900 ;
        RECT 24.985 59.755 25.155 59.945 ;
        RECT 28.205 59.925 28.355 59.945 ;
        RECT 25.260 59.735 25.430 59.925 ;
        RECT 28.205 59.755 28.375 59.925 ;
        RECT 29.135 59.780 29.295 59.890 ;
        RECT 29.590 59.755 29.760 59.945 ;
        RECT 30.955 59.735 31.125 59.925 ;
        RECT 31.890 59.735 32.060 59.925 ;
        RECT 32.800 59.755 32.970 59.945 ;
        RECT 34.190 59.755 34.360 59.945 ;
        RECT 34.640 59.785 34.760 59.895 ;
        RECT 37.405 59.735 37.575 59.925 ;
        RECT 37.840 59.735 38.010 59.925 ;
        RECT 43.845 59.755 44.015 59.945 ;
        RECT 44.770 59.735 44.940 59.925 ;
        RECT 46.600 59.755 46.770 59.945 ;
        RECT 47.525 59.735 47.695 59.925 ;
        RECT 50.770 59.755 50.940 59.945 ;
        RECT 56.725 59.735 56.895 59.925 ;
        RECT 59.945 59.755 60.115 59.945 ;
        RECT 64.545 59.735 64.715 59.925 ;
        RECT 69.145 59.755 69.315 59.945 ;
        RECT 73.280 59.925 73.425 59.945 ;
        RECT 69.600 59.785 69.720 59.895 ;
        RECT 73.280 59.755 73.450 59.925 ;
        RECT 73.745 59.735 73.915 59.925 ;
        RECT 74.205 59.735 74.375 59.925 ;
        RECT 75.125 59.755 75.295 59.945 ;
        RECT 76.505 59.735 76.675 59.945 ;
        RECT 5.525 58.925 6.895 59.735 ;
        RECT 6.905 59.055 8.735 59.735 ;
        RECT 6.905 58.825 8.250 59.055 ;
        RECT 8.765 58.825 10.115 59.735 ;
        RECT 10.255 58.825 13.255 59.735 ;
        RECT 14.265 59.055 17.935 59.735 ;
        RECT 14.265 58.825 15.190 59.055 ;
        RECT 19.325 58.825 20.675 59.735 ;
        RECT 20.705 59.055 24.605 59.735 ;
        RECT 24.845 59.055 28.745 59.735 ;
        RECT 20.705 58.825 21.635 59.055 ;
        RECT 24.845 58.825 25.775 59.055 ;
        RECT 29.905 58.955 31.275 59.735 ;
        RECT 31.295 58.865 31.725 59.650 ;
        RECT 31.745 58.825 36.045 59.735 ;
        RECT 36.345 58.955 37.715 59.735 ;
        RECT 37.780 58.825 41.855 59.735 ;
        RECT 41.865 58.825 45.065 59.735 ;
        RECT 45.095 59.055 47.835 59.735 ;
        RECT 47.930 59.055 57.035 59.735 ;
        RECT 57.055 58.865 57.485 59.650 ;
        RECT 57.945 58.825 64.855 59.735 ;
        RECT 64.950 59.055 74.055 59.735 ;
        RECT 74.075 58.825 75.425 59.735 ;
        RECT 75.445 58.925 76.815 59.735 ;
      LAYER nwell ;
        RECT 5.330 55.705 77.010 58.535 ;
      LAYER pwell ;
        RECT 5.525 54.505 6.895 55.315 ;
        RECT 6.905 54.505 8.275 55.285 ;
        RECT 8.765 54.505 10.115 55.415 ;
        RECT 10.255 54.505 13.255 55.415 ;
        RECT 14.265 55.185 15.190 55.415 ;
        RECT 14.265 54.505 17.935 55.185 ;
        RECT 18.415 54.590 18.845 55.375 ;
        RECT 18.865 54.505 20.235 55.285 ;
        RECT 20.245 55.185 21.175 55.415 ;
        RECT 20.245 54.505 24.145 55.185 ;
        RECT 24.385 54.505 25.755 55.285 ;
        RECT 26.225 54.505 27.595 55.285 ;
        RECT 28.535 54.505 31.265 55.415 ;
        RECT 31.745 54.505 35.820 55.415 ;
        RECT 35.885 54.505 39.540 55.415 ;
        RECT 39.565 54.505 42.775 55.415 ;
        RECT 42.795 54.505 44.145 55.415 ;
        RECT 44.175 54.590 44.605 55.375 ;
        RECT 54.285 55.185 57.110 55.415 ;
        RECT 45.170 54.505 54.275 55.185 ;
        RECT 54.285 54.505 57.815 55.185 ;
        RECT 57.975 54.505 60.715 55.185 ;
        RECT 60.810 54.505 69.915 55.185 ;
        RECT 69.935 54.590 70.365 55.375 ;
        RECT 70.385 54.505 74.040 55.415 ;
        RECT 74.065 54.505 75.415 55.415 ;
        RECT 75.445 54.505 76.815 55.315 ;
        RECT 5.665 54.295 5.835 54.505 ;
        RECT 7.055 54.315 7.225 54.505 ;
        RECT 7.965 54.295 8.135 54.485 ;
        RECT 8.420 54.345 8.540 54.455 ;
        RECT 8.880 54.315 9.050 54.505 ;
        RECT 10.255 54.295 10.425 54.485 ;
        RECT 10.725 54.295 10.895 54.485 ;
        RECT 13.025 54.315 13.195 54.505 ;
        RECT 13.480 54.460 13.650 54.485 ;
        RECT 13.480 54.350 13.655 54.460 ;
        RECT 13.480 54.295 13.650 54.350 ;
        RECT 14.410 54.315 14.580 54.505 ;
        RECT 14.855 54.295 15.025 54.485 ;
        RECT 15.335 54.295 15.505 54.485 ;
        RECT 16.715 54.295 16.885 54.485 ;
        RECT 18.085 54.455 18.255 54.485 ;
        RECT 18.080 54.345 18.255 54.455 ;
        RECT 18.085 54.295 18.255 54.345 ;
        RECT 19.915 54.315 20.085 54.505 ;
        RECT 20.375 54.295 20.545 54.485 ;
        RECT 20.660 54.315 20.830 54.505 ;
        RECT 20.855 54.340 21.015 54.450 ;
        RECT 21.760 54.295 21.930 54.485 ;
        RECT 23.145 54.295 23.315 54.485 ;
        RECT 24.525 54.315 24.695 54.505 ;
        RECT 25.900 54.345 26.020 54.455 ;
        RECT 27.275 54.315 27.445 54.505 ;
        RECT 27.755 54.350 27.915 54.460 ;
        RECT 28.665 54.295 28.835 54.485 ;
        RECT 30.965 54.315 31.135 54.505 ;
        RECT 31.420 54.345 31.540 54.455 ;
        RECT 34.185 54.295 34.355 54.485 ;
        RECT 34.655 54.340 34.815 54.450 ;
        RECT 35.590 54.315 35.760 54.505 ;
        RECT 36.030 54.315 36.200 54.505 ;
        RECT 36.475 54.295 36.645 54.485 ;
        RECT 36.945 54.295 37.115 54.485 ;
        RECT 38.325 54.295 38.495 54.485 ;
        RECT 39.705 54.315 39.875 54.505 ;
        RECT 41.085 54.295 41.255 54.485 ;
        RECT 41.545 54.295 41.715 54.485 ;
        RECT 43.845 54.315 44.015 54.505 ;
        RECT 44.760 54.345 44.880 54.455 ;
        RECT 48.445 54.315 48.615 54.485 ;
        RECT 48.445 54.295 48.605 54.315 ;
        RECT 51.665 54.295 51.835 54.485 ;
        RECT 52.130 54.295 52.300 54.485 ;
        RECT 53.510 54.295 53.680 54.485 ;
        RECT 53.965 54.315 54.135 54.505 ;
        RECT 57.615 54.485 57.815 54.505 ;
        RECT 57.645 54.295 57.815 54.485 ;
        RECT 60.405 54.315 60.575 54.505 ;
        RECT 66.845 54.295 67.015 54.485 ;
        RECT 68.230 54.295 68.400 54.485 ;
        RECT 69.605 54.315 69.775 54.505 ;
        RECT 70.530 54.315 70.700 54.505 ;
        RECT 73.290 54.295 73.460 54.485 ;
        RECT 74.210 54.315 74.380 54.505 ;
        RECT 76.505 54.295 76.675 54.505 ;
        RECT 5.525 53.485 6.895 54.295 ;
        RECT 7.825 53.515 9.195 54.295 ;
        RECT 9.205 53.515 10.575 54.295 ;
        RECT 10.585 53.615 12.415 54.295 ;
        RECT 12.445 53.385 13.795 54.295 ;
        RECT 13.805 53.515 15.175 54.295 ;
        RECT 15.185 53.515 16.555 54.295 ;
        RECT 16.565 53.515 17.935 54.295 ;
        RECT 17.955 53.385 19.305 54.295 ;
        RECT 19.325 53.515 20.695 54.295 ;
        RECT 21.645 53.385 22.995 54.295 ;
        RECT 23.005 53.485 28.515 54.295 ;
        RECT 28.525 53.485 31.275 54.295 ;
        RECT 31.295 53.425 31.725 54.210 ;
        RECT 31.775 53.385 34.495 54.295 ;
        RECT 35.425 53.515 36.795 54.295 ;
        RECT 36.815 53.385 38.165 54.295 ;
        RECT 38.185 53.515 39.555 54.295 ;
        RECT 39.565 53.385 41.380 54.295 ;
        RECT 41.405 53.385 44.615 54.295 ;
        RECT 44.950 53.385 48.605 54.295 ;
        RECT 48.765 53.385 51.975 54.295 ;
        RECT 51.985 53.385 53.335 54.295 ;
        RECT 53.365 53.385 56.840 54.295 ;
        RECT 57.055 53.425 57.485 54.210 ;
        RECT 57.505 53.615 66.610 54.295 ;
        RECT 66.705 53.485 68.075 54.295 ;
        RECT 68.085 53.385 73.040 54.295 ;
        RECT 73.145 53.615 75.420 54.295 ;
        RECT 74.050 53.385 75.420 53.615 ;
        RECT 75.445 53.485 76.815 54.295 ;
      LAYER nwell ;
        RECT 5.330 50.265 77.010 53.095 ;
      LAYER pwell ;
        RECT 5.525 49.065 6.895 49.875 ;
        RECT 8.875 49.745 9.805 49.975 ;
        RECT 7.970 49.065 9.805 49.745 ;
        RECT 10.125 49.745 11.490 49.975 ;
        RECT 15.165 49.745 16.095 49.975 ;
        RECT 10.125 49.065 13.335 49.745 ;
        RECT 13.345 49.065 16.095 49.745 ;
        RECT 16.565 49.065 18.380 49.975 ;
        RECT 18.415 49.150 18.845 49.935 ;
        RECT 19.785 49.065 22.705 49.975 ;
        RECT 23.005 49.065 24.835 49.975 ;
        RECT 24.860 49.065 28.515 49.975 ;
        RECT 28.525 49.065 32.195 49.975 ;
        RECT 32.205 49.745 33.125 49.975 ;
        RECT 32.205 49.065 35.790 49.745 ;
        RECT 36.345 49.065 38.175 49.975 ;
        RECT 38.185 49.745 39.115 49.975 ;
        RECT 42.765 49.745 43.695 49.975 ;
        RECT 38.185 49.065 40.935 49.745 ;
        RECT 40.945 49.065 43.695 49.745 ;
        RECT 44.175 49.150 44.605 49.935 ;
        RECT 44.625 49.065 47.835 49.975 ;
        RECT 47.845 49.065 49.195 49.975 ;
        RECT 49.225 49.065 51.975 49.975 ;
        RECT 52.440 49.295 54.275 49.975 ;
        RECT 52.440 49.065 54.130 49.295 ;
        RECT 54.645 49.065 60.715 49.975 ;
        RECT 60.725 49.065 69.830 49.745 ;
        RECT 69.935 49.150 70.365 49.935 ;
        RECT 70.385 49.065 73.595 49.975 ;
        RECT 74.090 49.745 75.435 49.975 ;
        RECT 73.605 49.065 75.435 49.745 ;
        RECT 75.445 49.065 76.815 49.875 ;
        RECT 5.665 48.855 5.835 49.065 ;
        RECT 7.970 49.045 8.135 49.065 ;
        RECT 13.020 49.045 13.190 49.065 ;
        RECT 7.055 48.855 7.225 49.045 ;
        RECT 7.965 48.875 8.135 49.045 ;
        RECT 8.435 48.900 8.595 49.010 ;
        RECT 9.350 48.855 9.520 49.045 ;
        RECT 13.020 48.875 13.195 49.045 ;
        RECT 13.485 48.875 13.655 49.065 ;
        RECT 13.025 48.855 13.195 48.875 ;
        RECT 14.405 48.855 14.575 49.045 ;
        RECT 14.865 48.855 15.035 49.045 ;
        RECT 16.245 49.015 16.415 49.045 ;
        RECT 16.240 48.905 16.415 49.015 ;
        RECT 16.245 48.855 16.415 48.905 ;
        RECT 18.085 48.875 18.255 49.065 ;
        RECT 19.930 49.045 20.100 49.065 ;
        RECT 19.015 48.910 19.175 49.020 ;
        RECT 19.925 48.875 20.100 49.045 ;
        RECT 19.925 48.855 20.095 48.875 ;
        RECT 21.300 48.855 21.470 49.045 ;
        RECT 22.685 48.855 22.855 49.045 ;
        RECT 23.150 48.875 23.320 49.065 ;
        RECT 28.200 49.045 28.370 49.065 ;
        RECT 28.200 48.875 28.375 49.045 ;
        RECT 28.670 48.875 28.840 49.065 ;
        RECT 30.960 48.905 31.080 49.015 ;
        RECT 28.205 48.855 28.375 48.875 ;
        RECT 31.885 48.855 32.055 49.045 ;
        RECT 32.350 48.875 32.520 49.065 ;
        RECT 35.105 48.855 35.275 49.045 ;
        RECT 36.020 48.905 36.140 49.015 ;
        RECT 36.490 48.875 36.660 49.065 ;
        RECT 36.945 48.855 37.115 49.045 ;
        RECT 39.710 48.855 39.880 49.045 ;
        RECT 40.625 48.875 40.795 49.065 ;
        RECT 41.085 48.855 41.255 49.065 ;
        RECT 42.465 48.855 42.635 49.045 ;
        RECT 43.835 48.855 44.005 49.045 ;
        RECT 44.765 48.875 44.935 49.065 ;
        RECT 47.525 48.875 47.695 49.045 ;
        RECT 47.495 48.855 47.695 48.875 ;
        RECT 47.980 48.855 48.150 49.045 ;
        RECT 48.910 48.875 49.080 49.065 ;
        RECT 49.370 48.855 49.540 49.065 ;
        RECT 52.120 48.905 52.240 49.015 ;
        RECT 52.590 48.855 52.760 49.045 ;
        RECT 53.960 48.875 54.130 49.065 ;
        RECT 60.400 49.045 60.570 49.065 ;
        RECT 56.275 48.900 56.435 49.010 ;
        RECT 59.945 48.855 60.115 49.045 ;
        RECT 60.400 48.875 60.575 49.045 ;
        RECT 60.865 48.875 61.035 49.065 ;
        RECT 73.285 49.045 73.455 49.065 ;
        RECT 69.615 48.900 69.775 49.010 ;
        RECT 73.280 48.875 73.455 49.045 ;
        RECT 60.405 48.855 60.575 48.875 ;
        RECT 73.280 48.855 73.450 48.875 ;
        RECT 73.745 48.855 73.915 49.065 ;
        RECT 76.505 48.855 76.675 49.065 ;
        RECT 5.525 48.045 6.895 48.855 ;
        RECT 6.905 48.075 8.275 48.855 ;
        RECT 9.350 48.625 11.040 48.855 ;
        RECT 9.205 47.945 11.040 48.625 ;
        RECT 11.505 48.175 13.335 48.855 ;
        RECT 11.505 47.945 12.850 48.175 ;
        RECT 13.345 48.075 14.715 48.855 ;
        RECT 14.725 48.075 16.095 48.855 ;
        RECT 16.105 48.045 19.775 48.855 ;
        RECT 19.785 48.045 21.155 48.855 ;
        RECT 21.185 47.945 22.535 48.855 ;
        RECT 22.545 48.045 28.055 48.855 ;
        RECT 28.065 48.045 30.815 48.855 ;
        RECT 31.295 47.985 31.725 48.770 ;
        RECT 31.745 48.175 34.955 48.855 ;
        RECT 33.820 47.945 34.955 48.175 ;
        RECT 34.980 47.945 36.795 48.855 ;
        RECT 36.805 48.045 38.635 48.855 ;
        RECT 38.645 47.945 39.995 48.855 ;
        RECT 40.025 48.075 41.395 48.855 ;
        RECT 41.405 48.075 42.775 48.855 ;
        RECT 42.785 48.075 44.155 48.855 ;
        RECT 44.165 48.175 47.695 48.855 ;
        RECT 44.165 47.945 46.990 48.175 ;
        RECT 47.865 47.945 49.215 48.855 ;
        RECT 49.225 47.945 51.975 48.855 ;
        RECT 52.445 48.175 56.030 48.855 ;
        RECT 52.445 47.945 53.365 48.175 ;
        RECT 57.055 47.985 57.485 48.770 ;
        RECT 57.515 48.175 60.255 48.855 ;
        RECT 60.265 48.175 69.370 48.855 ;
        RECT 70.395 48.625 73.450 48.855 ;
        RECT 70.395 47.945 73.595 48.625 ;
        RECT 73.605 48.045 75.435 48.855 ;
        RECT 75.445 48.045 76.815 48.855 ;
      LAYER nwell ;
        RECT 5.330 44.825 77.010 47.655 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 7.825 43.625 11.035 44.535 ;
        RECT 11.045 43.625 16.555 44.435 ;
        RECT 16.565 43.625 18.395 44.435 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 18.875 43.625 21.605 44.535 ;
        RECT 21.625 43.625 25.295 44.435 ;
        RECT 25.765 43.625 27.115 44.535 ;
        RECT 27.145 43.625 32.655 44.435 ;
        RECT 32.665 43.625 38.175 44.435 ;
        RECT 38.185 43.625 39.555 44.435 ;
        RECT 39.565 43.625 41.380 44.535 ;
        RECT 41.880 43.625 43.695 44.535 ;
        RECT 44.175 43.710 44.605 44.495 ;
        RECT 45.085 43.625 46.455 44.405 ;
        RECT 46.465 43.625 47.835 44.405 ;
        RECT 47.845 43.625 49.215 44.405 ;
        RECT 49.225 43.625 52.435 44.535 ;
        RECT 52.455 43.625 53.805 44.535 ;
        RECT 53.835 43.625 55.185 44.535 ;
        RECT 55.285 43.625 57.495 44.535 ;
        RECT 57.770 43.625 60.705 44.535 ;
        RECT 60.810 43.625 69.915 44.305 ;
        RECT 69.935 43.710 70.365 44.495 ;
        RECT 70.385 43.855 73.585 44.535 ;
        RECT 70.530 43.625 73.585 43.855 ;
        RECT 73.605 43.625 75.435 44.535 ;
        RECT 75.445 43.625 76.815 44.435 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.415 7.215 43.605 ;
        RECT 7.965 43.435 8.135 43.625 ;
        RECT 8.880 43.465 9.000 43.575 ;
        RECT 9.620 43.415 9.790 43.605 ;
        RECT 11.185 43.435 11.355 43.625 ;
        RECT 13.485 43.415 13.655 43.605 ;
        RECT 16.705 43.435 16.875 43.625 ;
        RECT 17.625 43.415 17.795 43.605 ;
        RECT 19.925 43.435 20.095 43.605 ;
        RECT 21.305 43.435 21.475 43.625 ;
        RECT 21.765 43.435 21.935 43.625 ;
        RECT 19.925 43.415 20.090 43.435 ;
        RECT 23.145 43.415 23.315 43.605 ;
        RECT 23.600 43.465 23.720 43.575 ;
        RECT 24.340 43.415 24.510 43.605 ;
        RECT 25.440 43.465 25.560 43.575 ;
        RECT 26.830 43.435 27.000 43.625 ;
        RECT 27.285 43.435 27.455 43.625 ;
        RECT 28.205 43.415 28.375 43.605 ;
        RECT 30.960 43.465 31.080 43.575 ;
        RECT 32.805 43.435 32.975 43.625 ;
        RECT 33.265 43.415 33.435 43.605 ;
        RECT 33.720 43.465 33.840 43.575 ;
        RECT 34.185 43.415 34.355 43.605 ;
        RECT 36.945 43.415 37.115 43.605 ;
        RECT 38.325 43.435 38.495 43.625 ;
        RECT 39.705 43.415 39.875 43.605 ;
        RECT 41.085 43.435 41.255 43.625 ;
        RECT 41.540 43.570 41.660 43.575 ;
        RECT 41.540 43.465 41.715 43.570 ;
        RECT 41.555 43.460 41.715 43.465 ;
        RECT 42.005 43.435 42.175 43.625 ;
        RECT 42.465 43.415 42.635 43.605 ;
        RECT 43.840 43.465 43.960 43.575 ;
        RECT 44.305 43.415 44.475 43.605 ;
        RECT 44.760 43.465 44.880 43.575 ;
        RECT 45.235 43.435 45.405 43.625 ;
        RECT 46.140 43.465 46.260 43.575 ;
        RECT 46.615 43.435 46.785 43.625 ;
        RECT 48.895 43.435 49.065 43.625 ;
        RECT 52.125 43.605 52.295 43.625 ;
        RECT 49.825 43.435 49.995 43.605 ;
        RECT 50.280 43.465 50.400 43.575 ;
        RECT 49.795 43.415 49.995 43.435 ;
        RECT 50.745 43.415 50.915 43.605 ;
        RECT 52.125 43.435 52.305 43.605 ;
        RECT 53.505 43.435 53.675 43.625 ;
        RECT 53.965 43.435 54.135 43.625 ;
        RECT 52.135 43.415 52.305 43.435 ;
        RECT 56.720 43.415 56.890 43.605 ;
        RECT 57.180 43.435 57.350 43.625 ;
        RECT 57.770 43.605 57.815 43.625 ;
        RECT 57.645 43.435 57.815 43.605 ;
        RECT 58.570 43.415 58.740 43.605 ;
        RECT 64.085 43.415 64.255 43.605 ;
        RECT 64.545 43.415 64.715 43.605 ;
        RECT 66.385 43.415 66.555 43.605 ;
        RECT 69.605 43.435 69.775 43.625 ;
        RECT 70.530 43.435 70.700 43.625 ;
        RECT 75.120 43.435 75.290 43.625 ;
        RECT 76.505 43.415 76.675 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.905 42.605 8.735 43.415 ;
        RECT 9.205 42.735 13.105 43.415 ;
        RECT 9.205 42.505 10.135 42.735 ;
        RECT 13.345 42.605 16.095 43.415 ;
        RECT 16.105 42.505 17.920 43.415 ;
        RECT 18.255 42.735 20.090 43.415 ;
        RECT 18.255 42.505 19.185 42.735 ;
        RECT 20.245 42.505 23.455 43.415 ;
        RECT 23.925 42.735 27.825 43.415 ;
        RECT 23.925 42.505 24.855 42.735 ;
        RECT 28.065 42.605 30.815 43.415 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.745 42.505 33.560 43.415 ;
        RECT 34.055 42.505 36.785 43.415 ;
        RECT 36.805 42.605 39.555 43.415 ;
        RECT 39.580 42.505 41.395 43.415 ;
        RECT 42.340 42.505 44.155 43.415 ;
        RECT 44.165 42.605 45.995 43.415 ;
        RECT 46.465 42.735 49.995 43.415 ;
        RECT 46.465 42.505 49.290 42.735 ;
        RECT 50.605 42.635 51.975 43.415 ;
        RECT 51.985 42.635 53.355 43.415 ;
        RECT 53.380 42.505 57.035 43.415 ;
        RECT 57.055 42.545 57.485 43.330 ;
        RECT 58.425 42.505 60.635 43.415 ;
        RECT 60.865 42.505 64.315 43.415 ;
        RECT 64.405 42.735 66.235 43.415 ;
        RECT 66.245 42.735 75.350 43.415 ;
        RECT 64.890 42.505 66.235 42.735 ;
        RECT 75.445 42.605 76.815 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 77.010 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 6.905 38.185 8.735 38.995 ;
        RECT 8.745 38.865 9.675 39.095 ;
        RECT 8.745 38.185 12.645 38.865 ;
        RECT 12.885 38.185 14.715 38.995 ;
        RECT 15.185 38.185 17.000 39.095 ;
        RECT 17.025 38.185 18.395 38.995 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 19.175 38.865 20.105 39.095 ;
        RECT 19.175 38.185 21.010 38.865 ;
        RECT 21.165 38.185 22.980 39.095 ;
        RECT 23.925 38.865 24.855 39.095 ;
        RECT 23.925 38.185 27.825 38.865 ;
        RECT 28.075 38.185 29.425 39.095 ;
        RECT 29.445 38.185 30.795 39.095 ;
        RECT 30.825 38.185 32.195 38.995 ;
        RECT 32.220 38.185 34.035 39.095 ;
        RECT 34.045 38.185 35.875 38.995 ;
        RECT 36.345 38.185 37.695 39.095 ;
        RECT 37.725 38.185 43.235 38.995 ;
        RECT 44.175 38.270 44.605 39.055 ;
        RECT 44.625 38.895 45.570 39.095 ;
        RECT 46.905 38.895 47.835 39.095 ;
        RECT 44.625 38.415 47.835 38.895 ;
        RECT 44.625 38.215 47.695 38.415 ;
        RECT 44.625 38.185 45.570 38.215 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.045 37.975 7.215 38.185 ;
        RECT 9.160 37.995 9.330 38.185 ;
        RECT 10.080 37.975 10.250 38.165 ;
        RECT 13.025 37.995 13.195 38.185 ;
        RECT 14.220 37.975 14.390 38.165 ;
        RECT 14.860 38.025 14.980 38.135 ;
        RECT 16.705 37.995 16.875 38.185 ;
        RECT 17.165 37.995 17.335 38.185 ;
        RECT 20.845 38.165 21.010 38.185 ;
        RECT 18.085 37.975 18.255 38.165 ;
        RECT 20.845 37.995 21.015 38.165 ;
        RECT 22.685 37.995 22.855 38.185 ;
        RECT 23.155 38.030 23.315 38.140 ;
        RECT 23.605 37.975 23.775 38.165 ;
        RECT 24.340 37.995 24.510 38.185 ;
        RECT 28.205 37.995 28.375 38.185 ;
        RECT 29.125 37.975 29.295 38.165 ;
        RECT 30.510 37.995 30.680 38.185 ;
        RECT 30.965 38.135 31.135 38.185 ;
        RECT 30.960 38.025 31.135 38.135 ;
        RECT 30.965 37.995 31.135 38.025 ;
        RECT 31.885 37.975 32.055 38.165 ;
        RECT 32.345 37.995 32.515 38.185 ;
        RECT 33.265 37.975 33.435 38.165 ;
        RECT 34.185 37.995 34.355 38.185 ;
        RECT 35.110 37.975 35.280 38.165 ;
        RECT 36.020 38.025 36.140 38.135 ;
        RECT 37.410 37.995 37.580 38.185 ;
        RECT 37.865 37.995 38.035 38.185 ;
        RECT 38.785 37.975 38.955 38.165 ;
        RECT 40.630 37.975 40.800 38.165 ;
        RECT 43.395 38.030 43.555 38.140 ;
        RECT 47.060 37.975 47.230 38.165 ;
        RECT 47.525 37.995 47.695 38.215 ;
        RECT 47.845 38.185 51.515 38.995 ;
        RECT 51.985 38.185 55.195 39.095 ;
        RECT 56.595 39.005 58.185 39.095 ;
        RECT 55.205 38.185 56.575 38.995 ;
        RECT 56.595 38.185 59.165 39.005 ;
        RECT 59.425 38.185 62.425 39.095 ;
        RECT 62.575 38.185 65.510 39.095 ;
        RECT 65.795 38.185 67.145 39.095 ;
        RECT 67.175 38.185 69.915 38.865 ;
        RECT 69.935 38.270 70.365 39.055 ;
        RECT 70.395 38.415 73.595 39.095 ;
        RECT 70.395 38.185 73.450 38.415 ;
        RECT 73.605 38.185 75.435 38.995 ;
        RECT 75.445 38.185 76.815 38.995 ;
        RECT 47.985 37.995 48.155 38.185 ;
        RECT 47.530 37.975 47.695 37.995 ;
        RECT 50.750 37.975 50.920 38.165 ;
        RECT 51.205 37.975 51.375 38.165 ;
        RECT 51.660 38.025 51.780 38.135 ;
        RECT 52.115 37.995 52.285 38.185 ;
        RECT 52.595 37.975 52.765 38.165 ;
        RECT 53.975 37.975 54.145 38.165 ;
        RECT 55.345 37.975 55.515 38.185 ;
        RECT 59.025 38.165 59.165 38.185 ;
        RECT 59.485 38.165 59.655 38.185 ;
        RECT 65.465 38.165 65.510 38.185 ;
        RECT 59.025 37.975 59.195 38.165 ;
        RECT 59.485 37.995 59.660 38.165 ;
        RECT 59.490 37.975 59.660 37.995 ;
        RECT 61.785 37.975 61.955 38.165 ;
        RECT 65.465 37.995 65.635 38.165 ;
        RECT 66.385 37.975 66.555 38.165 ;
        RECT 66.845 37.995 67.015 38.185 ;
        RECT 69.605 37.995 69.775 38.185 ;
        RECT 73.280 37.995 73.450 38.185 ;
        RECT 73.745 37.995 73.915 38.185 ;
        RECT 76.505 37.975 76.675 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.905 37.165 9.655 37.975 ;
        RECT 9.665 37.295 13.565 37.975 ;
        RECT 13.805 37.295 17.705 37.975 ;
        RECT 9.665 37.065 10.595 37.295 ;
        RECT 13.805 37.065 14.735 37.295 ;
        RECT 17.945 37.165 23.455 37.975 ;
        RECT 23.465 37.165 28.975 37.975 ;
        RECT 28.985 37.165 30.815 37.975 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.755 37.065 33.105 37.975 ;
        RECT 33.125 37.165 34.955 37.975 ;
        RECT 34.965 37.295 38.635 37.975 ;
        RECT 34.965 37.065 35.890 37.295 ;
        RECT 38.645 37.165 40.475 37.975 ;
        RECT 40.485 37.065 43.405 37.975 ;
        RECT 43.900 37.065 47.375 37.975 ;
        RECT 47.530 37.295 49.365 37.975 ;
        RECT 48.435 37.065 49.365 37.295 ;
        RECT 49.685 37.065 51.035 37.975 ;
        RECT 51.065 37.165 52.435 37.975 ;
        RECT 52.445 37.195 53.815 37.975 ;
        RECT 53.825 37.195 55.195 37.975 ;
        RECT 55.220 37.065 57.035 37.975 ;
        RECT 57.055 37.105 57.485 37.890 ;
        RECT 57.505 37.065 59.320 37.975 ;
        RECT 59.345 37.065 61.535 37.975 ;
        RECT 61.725 37.065 65.175 37.975 ;
        RECT 66.245 37.295 75.350 37.975 ;
        RECT 75.445 37.165 76.815 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 77.010 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 32.745 8.735 33.555 ;
        RECT 8.745 32.745 11.955 33.655 ;
        RECT 11.965 32.745 17.475 33.555 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 18.875 32.745 20.225 33.655 ;
        RECT 20.245 32.745 21.615 33.555 ;
        RECT 21.625 33.425 22.555 33.655 ;
        RECT 21.625 32.745 25.525 33.425 ;
        RECT 25.765 32.745 27.115 33.655 ;
        RECT 27.145 32.745 30.815 33.555 ;
        RECT 30.825 32.745 34.035 33.655 ;
        RECT 34.045 32.745 39.555 33.555 ;
        RECT 39.565 32.745 43.235 33.555 ;
        RECT 44.175 32.830 44.605 33.615 ;
        RECT 44.625 33.455 45.570 33.655 ;
        RECT 46.905 33.455 47.835 33.655 ;
        RECT 44.625 32.975 47.835 33.455 ;
        RECT 44.625 32.775 47.695 32.975 ;
        RECT 44.625 32.745 45.570 32.775 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.045 32.555 7.215 32.745 ;
        RECT 8.425 32.535 8.595 32.725 ;
        RECT 8.885 32.535 9.055 32.725 ;
        RECT 11.645 32.535 11.815 32.745 ;
        RECT 12.105 32.535 12.275 32.745 ;
        RECT 15.795 32.580 15.955 32.690 ;
        RECT 16.700 32.535 16.870 32.725 ;
        RECT 17.635 32.590 17.795 32.700 ;
        RECT 19.925 32.555 20.095 32.745 ;
        RECT 20.385 32.555 20.555 32.745 ;
        RECT 20.845 32.535 21.015 32.725 ;
        RECT 21.580 32.535 21.750 32.725 ;
        RECT 22.040 32.555 22.210 32.745 ;
        RECT 25.445 32.555 25.615 32.725 ;
        RECT 26.830 32.555 27.000 32.745 ;
        RECT 27.285 32.555 27.455 32.745 ;
        RECT 27.740 32.585 27.860 32.695 ;
        RECT 28.205 32.555 28.375 32.725 ;
        RECT 30.515 32.580 30.675 32.690 ;
        RECT 30.955 32.555 31.125 32.745 ;
        RECT 34.185 32.555 34.355 32.745 ;
        RECT 35.565 32.555 35.735 32.725 ;
        RECT 25.465 32.535 25.615 32.555 ;
        RECT 28.210 32.535 28.375 32.555 ;
        RECT 35.565 32.535 35.725 32.555 ;
        RECT 39.240 32.535 39.410 32.725 ;
        RECT 39.705 32.535 39.875 32.745 ;
        RECT 43.395 32.590 43.555 32.700 ;
        RECT 45.225 32.535 45.395 32.725 ;
        RECT 45.685 32.535 45.855 32.725 ;
        RECT 47.525 32.555 47.695 32.775 ;
        RECT 48.765 32.745 53.155 33.655 ;
        RECT 47.995 32.590 48.155 32.700 ;
        RECT 48.910 32.555 49.080 32.745 ;
        RECT 49.375 32.580 49.535 32.690 ;
        RECT 52.585 32.535 52.755 32.725 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.905 31.855 8.735 32.535 ;
        RECT 8.745 31.855 10.575 32.535 ;
        RECT 6.905 31.625 8.250 31.855 ;
        RECT 10.585 31.755 11.955 32.535 ;
        RECT 11.965 31.725 15.635 32.535 ;
        RECT 16.585 31.625 17.935 32.535 ;
        RECT 17.945 31.625 21.155 32.535 ;
        RECT 21.165 31.855 25.065 32.535 ;
        RECT 21.165 31.625 22.095 31.855 ;
        RECT 25.465 31.715 27.395 32.535 ;
        RECT 28.210 31.855 30.045 32.535 ;
        RECT 26.445 31.625 27.395 31.715 ;
        RECT 29.115 31.625 30.045 31.855 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 32.070 31.625 35.725 32.535 ;
        RECT 35.885 31.625 39.555 32.535 ;
        RECT 39.565 31.725 42.315 32.535 ;
        RECT 42.755 31.625 45.535 32.535 ;
        RECT 45.545 31.725 49.215 32.535 ;
        RECT 50.155 31.625 52.885 32.535 ;
        RECT 53.050 32.505 53.220 32.725 ;
        RECT 53.825 32.705 54.715 33.655 ;
        RECT 54.745 32.745 56.095 33.655 ;
        RECT 56.125 33.425 57.470 33.655 ;
        RECT 58.450 33.425 59.795 33.655 ;
        RECT 61.635 33.425 62.555 33.655 ;
        RECT 64.820 33.455 65.775 33.655 ;
        RECT 56.125 32.745 57.955 33.425 ;
        RECT 57.965 32.745 59.795 33.425 ;
        RECT 60.265 32.745 62.555 33.425 ;
        RECT 63.495 32.775 65.775 33.455 ;
        RECT 53.500 32.585 53.620 32.695 ;
        RECT 54.425 32.555 54.595 32.705 ;
        RECT 54.890 32.555 55.060 32.745 ;
        RECT 55.805 32.535 55.975 32.725 ;
        RECT 57.645 32.535 57.815 32.745 ;
        RECT 58.105 32.555 58.275 32.745 ;
        RECT 59.940 32.585 60.060 32.695 ;
        RECT 60.405 32.555 60.575 32.745 ;
        RECT 62.705 32.535 62.875 32.725 ;
        RECT 63.165 32.535 63.335 32.725 ;
        RECT 63.620 32.555 63.790 32.775 ;
        RECT 64.820 32.745 65.775 32.775 ;
        RECT 65.785 32.745 67.155 33.525 ;
        RECT 67.175 32.745 69.915 33.425 ;
        RECT 69.935 32.830 70.365 33.615 ;
        RECT 70.385 32.745 71.755 33.525 ;
        RECT 71.845 32.745 75.430 33.655 ;
        RECT 75.445 32.745 76.815 33.555 ;
        RECT 65.465 32.535 65.635 32.725 ;
        RECT 65.935 32.555 66.105 32.745 ;
        RECT 69.605 32.535 69.775 32.745 ;
        RECT 70.075 32.580 70.235 32.690 ;
        RECT 70.535 32.555 70.705 32.745 ;
        RECT 75.120 32.535 75.290 32.745 ;
        RECT 76.505 32.535 76.675 32.745 ;
        RECT 54.710 32.505 55.655 32.535 ;
        RECT 52.905 31.825 55.655 32.505 ;
        RECT 54.710 31.625 55.655 31.825 ;
        RECT 55.665 31.725 57.035 32.535 ;
        RECT 57.055 31.665 57.485 32.450 ;
        RECT 57.505 31.625 60.715 32.535 ;
        RECT 60.725 31.855 63.015 32.535 ;
        RECT 63.025 31.855 65.315 32.535 ;
        RECT 60.725 31.625 61.645 31.855 ;
        RECT 64.395 31.625 65.315 31.855 ;
        RECT 65.325 31.725 67.155 32.535 ;
        RECT 67.165 31.855 69.915 32.535 ;
        RECT 70.845 31.855 75.435 32.535 ;
        RECT 67.165 31.625 68.095 31.855 ;
        RECT 73.610 31.625 74.950 31.855 ;
        RECT 75.445 31.725 76.815 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 77.010 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 7.825 27.305 9.655 28.215 ;
        RECT 11.510 27.985 12.875 28.215 ;
        RECT 9.665 27.305 12.875 27.985 ;
        RECT 12.885 27.305 14.715 28.215 ;
        RECT 14.725 27.305 18.395 28.115 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 20.475 28.125 22.065 28.215 ;
        RECT 19.495 27.305 22.065 28.125 ;
        RECT 22.085 27.985 23.430 28.215 ;
        RECT 22.085 27.305 23.915 27.985 ;
        RECT 23.925 27.305 29.435 28.115 ;
        RECT 29.445 27.305 33.115 28.115 ;
        RECT 33.125 27.305 35.875 28.215 ;
        RECT 35.885 27.305 39.095 28.215 ;
        RECT 40.950 27.985 42.315 28.215 ;
        RECT 39.105 27.305 42.315 27.985 ;
        RECT 42.325 27.305 44.155 28.115 ;
        RECT 44.175 27.390 44.605 28.175 ;
        RECT 44.625 27.305 50.135 28.115 ;
        RECT 51.080 27.305 52.895 28.215 ;
        RECT 52.905 27.305 58.415 28.115 ;
        RECT 58.425 27.305 60.255 28.115 ;
        RECT 61.635 27.985 62.555 28.215 ;
        RECT 60.265 27.305 62.555 27.985 ;
        RECT 62.565 27.305 63.935 28.115 ;
        RECT 63.965 27.305 65.315 28.215 ;
        RECT 66.660 28.015 67.615 28.215 ;
        RECT 65.335 27.335 67.615 28.015 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.020 27.260 7.190 27.285 ;
        RECT 7.020 27.150 7.215 27.260 ;
        RECT 7.020 27.115 7.190 27.150 ;
        RECT 7.970 27.115 8.140 27.305 ;
        RECT 9.810 27.115 9.980 27.305 ;
        RECT 14.400 27.285 14.570 27.305 ;
        RECT 13.945 27.115 14.115 27.285 ;
        RECT 14.400 27.115 14.575 27.285 ;
        RECT 14.865 27.115 15.035 27.305 ;
        RECT 19.495 27.285 19.635 27.305 ;
        RECT 7.080 27.095 7.190 27.115 ;
        RECT 13.945 27.095 14.085 27.115 ;
        RECT 14.405 27.095 14.575 27.115 ;
        RECT 16.250 27.095 16.420 27.285 ;
        RECT 19.000 27.145 19.120 27.255 ;
        RECT 19.465 27.115 19.635 27.285 ;
        RECT 22.225 27.095 22.395 27.285 ;
        RECT 22.695 27.140 22.855 27.250 ;
        RECT 23.605 27.115 23.775 27.305 ;
        RECT 24.065 27.115 24.235 27.305 ;
        RECT 26.825 27.095 26.995 27.285 ;
        RECT 27.285 27.095 27.455 27.285 ;
        RECT 29.585 27.115 29.755 27.305 ;
        RECT 30.960 27.145 31.080 27.255 ;
        RECT 33.265 27.115 33.435 27.305 ;
        RECT 34.655 27.095 34.825 27.285 ;
        RECT 35.105 27.095 35.275 27.285 ;
        RECT 37.865 27.095 38.035 27.285 ;
        RECT 38.785 27.115 38.955 27.305 ;
        RECT 39.250 27.115 39.420 27.305 ;
        RECT 40.620 27.095 40.790 27.285 ;
        RECT 41.085 27.095 41.255 27.285 ;
        RECT 42.465 27.115 42.635 27.305 ;
        RECT 44.765 27.095 44.935 27.305 ;
        RECT 47.985 27.095 48.155 27.285 ;
        RECT 49.820 27.145 49.940 27.255 ;
        RECT 50.295 27.150 50.455 27.260 ;
        RECT 51.205 27.095 51.375 27.305 ;
        RECT 51.665 27.095 51.835 27.285 ;
        RECT 53.045 27.115 53.215 27.305 ;
        RECT 58.565 27.115 58.735 27.305 ;
        RECT 59.945 27.095 60.115 27.285 ;
        RECT 60.405 27.115 60.575 27.305 ;
        RECT 62.705 27.115 62.875 27.305 ;
        RECT 63.165 27.115 63.335 27.285 ;
        RECT 63.165 27.095 63.315 27.115 ;
        RECT 63.625 27.095 63.795 27.285 ;
        RECT 65.000 27.115 65.170 27.305 ;
        RECT 65.460 27.115 65.630 27.335 ;
        RECT 66.660 27.305 67.615 27.335 ;
        RECT 67.705 27.305 69.915 28.215 ;
        RECT 69.935 27.390 70.365 28.175 ;
        RECT 70.385 27.305 71.755 28.085 ;
        RECT 71.765 28.015 73.175 28.215 ;
        RECT 71.765 27.335 74.500 28.015 ;
        RECT 71.765 27.305 73.160 27.335 ;
        RECT 69.600 27.285 69.770 27.305 ;
        RECT 66.380 27.145 66.500 27.255 ;
        RECT 67.755 27.095 67.925 27.285 ;
        RECT 69.600 27.115 69.775 27.285 ;
        RECT 69.605 27.095 69.775 27.115 ;
        RECT 70.075 27.095 70.245 27.285 ;
        RECT 70.535 27.115 70.705 27.305 ;
        RECT 71.440 27.145 71.560 27.255 ;
        RECT 73.285 27.095 73.455 27.285 ;
        RECT 74.205 27.115 74.375 27.335 ;
        RECT 75.445 27.305 76.815 28.115 ;
        RECT 74.675 27.150 74.835 27.260 ;
        RECT 75.125 27.095 75.295 27.285 ;
        RECT 76.505 27.095 76.675 27.305 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 7.080 26.415 11.495 27.095 ;
        RECT 7.565 26.185 11.495 26.415 ;
        RECT 11.515 26.275 14.085 27.095 ;
        RECT 14.265 26.285 16.095 27.095 ;
        RECT 16.105 26.415 20.695 27.095 ;
        RECT 20.705 26.415 22.535 27.095 ;
        RECT 11.515 26.185 13.105 26.275 ;
        RECT 16.590 26.185 17.930 26.415 ;
        RECT 20.705 26.185 22.050 26.415 ;
        RECT 23.605 26.185 27.055 27.095 ;
        RECT 27.145 26.285 30.815 27.095 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 31.745 26.185 34.955 27.095 ;
        RECT 34.975 26.185 37.705 27.095 ;
        RECT 37.725 26.285 39.555 27.095 ;
        RECT 39.585 26.185 40.935 27.095 ;
        RECT 40.945 26.285 44.615 27.095 ;
        RECT 44.625 26.185 47.835 27.095 ;
        RECT 47.845 26.285 49.675 27.095 ;
        RECT 50.155 26.185 51.505 27.095 ;
        RECT 51.525 26.285 57.035 27.095 ;
        RECT 57.055 26.225 57.485 27.010 ;
        RECT 57.515 26.185 60.245 27.095 ;
        RECT 61.385 26.275 63.315 27.095 ;
        RECT 63.485 26.285 66.235 27.095 ;
        RECT 66.705 26.315 68.075 27.095 ;
        RECT 68.085 26.415 69.915 27.095 ;
        RECT 61.385 26.185 62.335 26.275 ;
        RECT 68.085 26.185 69.430 26.415 ;
        RECT 69.925 26.315 71.295 27.095 ;
        RECT 71.765 26.415 73.595 27.095 ;
        RECT 73.605 26.415 75.435 27.095 ;
        RECT 71.765 26.185 73.110 26.415 ;
        RECT 75.445 26.285 76.815 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 77.010 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 6.905 22.545 8.250 22.775 ;
        RECT 11.485 22.545 12.415 22.775 ;
        RECT 6.905 21.865 8.735 22.545 ;
        RECT 9.665 21.865 12.415 22.545 ;
        RECT 12.425 21.865 15.175 22.675 ;
        RECT 15.185 22.575 16.115 22.775 ;
        RECT 17.445 22.575 18.395 22.775 ;
        RECT 15.185 22.095 18.395 22.575 ;
        RECT 15.330 21.895 18.395 22.095 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 21.605 22.545 22.535 22.775 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.055 21.700 7.215 21.810 ;
        RECT 7.965 21.655 8.135 21.845 ;
        RECT 8.425 21.675 8.595 21.865 ;
        RECT 8.895 21.710 9.055 21.820 ;
        RECT 9.805 21.675 9.975 21.865 ;
        RECT 10.265 21.655 10.435 21.845 ;
        RECT 10.725 21.655 10.895 21.845 ;
        RECT 12.565 21.675 12.735 21.865 ;
        RECT 14.400 21.705 14.520 21.815 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 7.835 20.745 9.185 21.655 ;
        RECT 9.205 20.875 10.575 21.655 ;
        RECT 10.585 20.845 14.255 21.655 ;
        RECT 14.870 21.625 15.040 21.845 ;
        RECT 15.330 21.675 15.500 21.895 ;
        RECT 17.460 21.865 18.395 21.895 ;
        RECT 18.865 21.865 22.535 22.545 ;
        RECT 23.005 21.865 27.125 22.775 ;
        RECT 29.470 22.545 30.815 22.775 ;
        RECT 27.145 21.865 28.975 22.545 ;
        RECT 28.985 21.865 30.815 22.545 ;
        RECT 31.025 22.685 31.975 22.775 ;
        RECT 31.025 21.865 32.955 22.685 ;
        RECT 33.125 22.095 34.960 22.775 ;
        RECT 18.085 21.655 18.255 21.845 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 21.765 21.655 21.935 21.845 ;
        RECT 22.680 21.705 22.800 21.815 ;
        RECT 23.145 21.655 23.315 21.865 ;
        RECT 24.985 21.675 25.155 21.865 ;
        RECT 26.820 21.655 26.990 21.845 ;
        RECT 27.285 21.655 27.455 21.845 ;
        RECT 28.665 21.675 28.835 21.865 ;
        RECT 29.125 21.675 29.295 21.865 ;
        RECT 32.805 21.845 32.955 21.865 ;
        RECT 33.270 21.865 34.960 22.095 ;
        RECT 35.425 21.865 37.255 22.675 ;
        RECT 37.725 21.865 41.395 22.775 ;
        RECT 41.405 22.545 42.750 22.775 ;
        RECT 41.405 21.865 43.235 22.545 ;
        RECT 44.175 21.950 44.605 22.735 ;
        RECT 44.625 21.865 46.455 22.675 ;
        RECT 46.965 22.545 48.340 22.775 ;
        RECT 50.130 22.545 51.510 22.775 ;
        RECT 52.010 22.545 55.620 22.775 ;
        RECT 46.965 22.095 51.510 22.545 ;
        RECT 30.960 21.705 31.080 21.815 ;
        RECT 31.885 21.655 32.055 21.845 ;
        RECT 32.805 21.675 32.975 21.845 ;
        RECT 33.270 21.675 33.440 21.865 ;
        RECT 35.565 21.675 35.735 21.865 ;
        RECT 37.400 21.705 37.520 21.815 ;
        RECT 37.865 21.655 38.035 21.865 ;
        RECT 42.925 21.675 43.095 21.865 ;
        RECT 43.385 21.675 43.555 21.845 ;
        RECT 43.385 21.655 43.550 21.675 ;
        RECT 43.850 21.655 44.020 21.845 ;
        RECT 44.765 21.675 44.935 21.865 ;
        RECT 45.225 21.655 45.395 21.845 ;
        RECT 46.600 21.705 46.720 21.815 ;
        RECT 47.070 21.675 47.240 22.095 ;
        RECT 48.350 21.865 51.510 22.095 ;
        RECT 51.525 21.865 55.620 22.545 ;
        RECT 55.665 21.865 57.035 22.675 ;
        RECT 57.060 21.865 58.875 22.775 ;
        RECT 58.885 21.865 64.395 22.675 ;
        RECT 64.405 21.865 69.915 22.675 ;
        RECT 69.935 21.950 70.365 22.735 ;
        RECT 70.385 21.865 71.755 22.645 ;
        RECT 72.685 21.865 74.055 22.645 ;
        RECT 74.065 21.865 75.435 22.645 ;
        RECT 75.445 21.865 76.815 22.675 ;
        RECT 48.455 21.700 48.615 21.810 ;
        RECT 49.360 21.655 49.530 21.845 ;
        RECT 51.670 21.655 51.840 21.865 ;
        RECT 52.125 21.655 52.295 21.845 ;
        RECT 54.880 21.705 55.000 21.815 ;
        RECT 55.805 21.675 55.975 21.865 ;
        RECT 56.725 21.655 56.895 21.845 ;
        RECT 57.185 21.675 57.355 21.865 ;
        RECT 59.025 21.675 59.195 21.865 ;
        RECT 59.945 21.655 60.115 21.845 ;
        RECT 60.405 21.655 60.575 21.845 ;
        RECT 64.545 21.675 64.715 21.865 ;
        RECT 65.925 21.655 66.095 21.845 ;
        RECT 71.445 21.655 71.615 21.865 ;
        RECT 71.915 21.710 72.075 21.820 ;
        RECT 73.735 21.675 73.905 21.865 ;
        RECT 74.215 21.675 74.385 21.865 ;
        RECT 75.120 21.705 75.240 21.815 ;
        RECT 76.505 21.655 76.675 21.865 ;
        RECT 17.000 21.625 17.935 21.655 ;
        RECT 14.870 21.425 17.935 21.625 ;
        RECT 14.725 20.945 17.935 21.425 ;
        RECT 14.725 20.745 15.655 20.945 ;
        RECT 16.985 20.745 17.935 20.945 ;
        RECT 17.945 20.845 21.615 21.655 ;
        RECT 21.625 20.845 22.995 21.655 ;
        RECT 23.020 20.745 24.835 21.655 ;
        RECT 25.785 20.745 27.135 21.655 ;
        RECT 27.145 20.845 30.815 21.655 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.845 37.255 21.655 ;
        RECT 37.725 20.745 41.395 21.655 ;
        RECT 41.715 20.975 43.550 21.655 ;
        RECT 41.715 20.745 42.645 20.975 ;
        RECT 43.705 20.745 45.055 21.655 ;
        RECT 45.085 20.745 48.295 21.655 ;
        RECT 49.245 20.745 50.595 21.655 ;
        RECT 50.605 20.745 51.955 21.655 ;
        RECT 51.985 20.845 54.735 21.655 ;
        RECT 55.205 20.745 57.020 21.655 ;
        RECT 57.055 20.785 57.485 21.570 ;
        RECT 57.515 20.745 60.245 21.655 ;
        RECT 60.265 20.845 65.775 21.655 ;
        RECT 65.785 20.845 71.295 21.655 ;
        RECT 71.305 20.845 74.975 21.655 ;
        RECT 75.445 20.845 76.815 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 77.010 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.905 16.425 12.415 17.235 ;
        RECT 12.425 16.425 17.935 17.235 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 18.865 16.425 22.535 17.235 ;
        RECT 23.635 16.425 27.135 17.335 ;
        RECT 27.145 16.425 28.975 17.335 ;
        RECT 28.985 16.425 32.655 17.235 ;
        RECT 33.135 16.655 36.335 17.335 ;
        RECT 33.135 16.425 36.190 16.655 ;
        RECT 36.345 16.425 41.855 17.235 ;
        RECT 41.865 16.425 43.695 17.235 ;
        RECT 44.175 16.510 44.605 17.295 ;
        RECT 45.580 17.105 46.955 17.335 ;
        RECT 48.725 17.105 49.675 17.335 ;
        RECT 45.580 16.655 49.675 17.105 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 7.045 16.215 7.215 16.425 ;
        RECT 12.565 16.215 12.735 16.425 ;
        RECT 18.085 16.375 18.255 16.405 ;
        RECT 18.080 16.265 18.255 16.375 ;
        RECT 18.085 16.215 18.255 16.265 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 23.635 16.405 23.770 16.425 ;
        RECT 22.670 16.380 22.840 16.405 ;
        RECT 21.775 16.260 21.935 16.370 ;
        RECT 22.670 16.270 22.855 16.380 ;
        RECT 22.670 16.215 22.840 16.270 ;
        RECT 23.600 16.235 23.770 16.405 ;
        RECT 26.360 16.215 26.530 16.405 ;
        RECT 28.660 16.235 28.830 16.425 ;
        RECT 29.125 16.235 29.295 16.425 ;
        RECT 29.580 16.215 29.750 16.405 ;
        RECT 30.970 16.215 31.140 16.405 ;
        RECT 31.885 16.215 32.055 16.405 ;
        RECT 32.800 16.265 32.920 16.375 ;
        RECT 33.725 16.215 33.895 16.405 ;
        RECT 35.105 16.215 35.275 16.405 ;
        RECT 36.020 16.235 36.190 16.425 ;
        RECT 36.485 16.235 36.655 16.425 ;
        RECT 40.625 16.215 40.795 16.405 ;
        RECT 42.005 16.235 42.175 16.425 ;
        RECT 43.840 16.265 43.960 16.375 ;
        RECT 44.775 16.270 44.935 16.380 ;
        RECT 45.685 16.235 45.855 16.655 ;
        RECT 46.965 16.425 49.675 16.655 ;
        RECT 50.180 17.105 53.790 17.335 ;
        RECT 50.180 16.425 54.275 17.105 ;
        RECT 54.285 16.425 59.795 17.235 ;
        RECT 59.805 16.425 65.315 17.235 ;
        RECT 65.325 16.425 68.995 17.235 ;
        RECT 69.935 16.510 70.365 17.295 ;
        RECT 70.385 16.425 73.135 17.235 ;
        RECT 73.605 16.425 75.435 17.105 ;
        RECT 75.445 16.425 76.815 17.235 ;
        RECT 46.145 16.215 46.315 16.405 ;
        RECT 49.820 16.265 49.940 16.375 ;
        RECT 51.665 16.215 51.835 16.405 ;
        RECT 53.960 16.235 54.130 16.425 ;
        RECT 54.425 16.235 54.595 16.425 ;
        RECT 57.645 16.215 57.815 16.405 ;
        RECT 59.945 16.235 60.115 16.425 ;
        RECT 63.165 16.215 63.335 16.405 ;
        RECT 65.465 16.235 65.635 16.425 ;
        RECT 68.685 16.215 68.855 16.405 ;
        RECT 69.155 16.270 69.315 16.380 ;
        RECT 70.525 16.235 70.695 16.425 ;
        RECT 73.280 16.265 73.400 16.375 ;
        RECT 75.125 16.235 75.295 16.425 ;
        RECT 76.505 16.215 76.675 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.405 12.415 16.215 ;
        RECT 12.425 15.405 17.935 16.215 ;
        RECT 17.945 15.405 21.615 16.215 ;
        RECT 22.555 15.305 26.215 16.215 ;
        RECT 26.245 15.305 27.595 16.215 ;
        RECT 27.620 15.535 29.895 16.215 ;
        RECT 27.620 15.305 28.990 15.535 ;
        RECT 29.905 15.305 31.255 16.215 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 31.745 15.535 33.575 16.215 ;
        RECT 33.585 15.435 34.955 16.215 ;
        RECT 34.965 15.405 40.475 16.215 ;
        RECT 40.485 15.405 45.995 16.215 ;
        RECT 46.005 15.405 51.515 16.215 ;
        RECT 51.525 15.405 57.035 16.215 ;
        RECT 57.055 15.345 57.485 16.130 ;
        RECT 57.505 15.405 63.015 16.215 ;
        RECT 63.025 15.405 68.535 16.215 ;
        RECT 68.545 15.405 74.055 16.215 ;
        RECT 75.445 15.405 76.815 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 77.010 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 12.415 11.795 ;
        RECT 14.725 10.985 18.395 11.795 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 25.965 11.805 26.915 11.895 ;
        RECT 18.865 10.985 22.535 11.795 ;
        RECT 23.005 10.985 24.375 11.765 ;
        RECT 24.385 10.985 25.755 11.795 ;
        RECT 25.965 10.985 27.895 11.805 ;
        RECT 28.550 11.665 29.895 11.895 ;
        RECT 28.065 10.985 29.895 11.665 ;
        RECT 29.905 10.985 31.275 11.765 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 32.665 10.985 34.495 11.665 ;
        RECT 34.505 10.985 35.875 11.795 ;
        RECT 36.370 11.665 37.715 11.895 ;
        RECT 35.885 10.985 37.715 11.665 ;
        RECT 37.725 10.985 43.235 11.795 ;
        RECT 44.175 11.070 44.605 11.855 ;
        RECT 44.625 10.985 50.135 11.795 ;
        RECT 50.145 10.985 55.655 11.795 ;
        RECT 55.665 10.985 57.035 11.795 ;
        RECT 57.055 11.070 57.485 11.855 ;
        RECT 57.505 10.985 63.015 11.795 ;
        RECT 63.025 10.985 68.535 11.795 ;
        RECT 68.545 10.985 69.915 11.795 ;
        RECT 69.935 11.070 70.365 11.855 ;
        RECT 70.385 10.985 74.055 11.795 ;
        RECT 74.065 10.985 75.435 11.795 ;
        RECT 75.445 10.985 76.815 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 12.575 10.830 12.735 10.940 ;
        RECT 14.405 10.795 14.575 10.965 ;
        RECT 14.865 10.795 15.035 10.985 ;
        RECT 19.005 10.795 19.175 10.985 ;
        RECT 22.680 10.825 22.800 10.935 ;
        RECT 23.145 10.795 23.315 10.985 ;
        RECT 24.525 10.795 24.695 10.985 ;
        RECT 27.745 10.965 27.895 10.985 ;
        RECT 27.745 10.795 27.915 10.965 ;
        RECT 28.205 10.795 28.375 10.985 ;
        RECT 30.055 10.795 30.225 10.985 ;
        RECT 31.895 10.830 32.055 10.940 ;
        RECT 32.805 10.795 32.975 10.985 ;
        RECT 34.645 10.795 34.815 10.985 ;
        RECT 36.025 10.795 36.195 10.985 ;
        RECT 37.865 10.795 38.035 10.985 ;
        RECT 43.395 10.830 43.555 10.940 ;
        RECT 44.765 10.795 44.935 10.985 ;
        RECT 50.285 10.795 50.455 10.985 ;
        RECT 55.805 10.795 55.975 10.985 ;
        RECT 57.645 10.795 57.815 10.985 ;
        RECT 63.165 10.795 63.335 10.985 ;
        RECT 68.685 10.795 68.855 10.985 ;
        RECT 70.525 10.795 70.695 10.985 ;
        RECT 74.205 10.795 74.375 10.985 ;
        RECT 76.505 10.795 76.675 10.985 ;
      LAYER li1 ;
        RECT 5.520 81.515 76.820 81.685 ;
        RECT 5.605 80.765 6.815 81.515 ;
        RECT 5.605 80.225 6.125 80.765 ;
        RECT 6.990 80.675 7.250 81.515 ;
        RECT 7.425 80.770 7.680 81.345 ;
        RECT 7.850 81.135 8.180 81.515 ;
        RECT 8.395 80.965 8.565 81.345 ;
        RECT 7.850 80.795 8.565 80.965 ;
        RECT 6.295 80.055 6.815 80.595 ;
        RECT 5.605 78.965 6.815 80.055 ;
        RECT 6.990 78.965 7.250 80.115 ;
        RECT 7.425 80.040 7.595 80.770 ;
        RECT 7.850 80.605 8.020 80.795 ;
        RECT 8.830 80.675 9.090 81.515 ;
        RECT 9.265 80.770 9.520 81.345 ;
        RECT 9.690 81.135 10.020 81.515 ;
        RECT 10.235 80.965 10.405 81.345 ;
        RECT 9.690 80.795 10.405 80.965 ;
        RECT 10.665 81.015 10.925 81.345 ;
        RECT 11.135 81.035 11.410 81.515 ;
        RECT 7.765 80.275 8.020 80.605 ;
        RECT 7.850 80.065 8.020 80.275 ;
        RECT 8.300 80.245 8.655 80.615 ;
        RECT 7.425 79.135 7.680 80.040 ;
        RECT 7.850 79.895 8.565 80.065 ;
        RECT 7.850 78.965 8.180 79.725 ;
        RECT 8.395 79.135 8.565 79.895 ;
        RECT 8.830 78.965 9.090 80.115 ;
        RECT 9.265 80.040 9.435 80.770 ;
        RECT 9.690 80.605 9.860 80.795 ;
        RECT 9.605 80.275 9.860 80.605 ;
        RECT 9.690 80.065 9.860 80.275 ;
        RECT 10.140 80.245 10.495 80.615 ;
        RECT 10.665 80.105 10.835 81.015 ;
        RECT 11.620 80.945 11.825 81.345 ;
        RECT 11.995 81.115 12.330 81.515 ;
        RECT 11.005 80.275 11.365 80.855 ;
        RECT 11.620 80.775 12.305 80.945 ;
        RECT 11.545 80.105 11.795 80.605 ;
        RECT 9.265 79.135 9.520 80.040 ;
        RECT 9.690 79.895 10.405 80.065 ;
        RECT 9.690 78.965 10.020 79.725 ;
        RECT 10.235 79.135 10.405 79.895 ;
        RECT 10.665 79.935 11.795 80.105 ;
        RECT 10.665 79.165 10.935 79.935 ;
        RECT 11.965 79.745 12.305 80.775 ;
        RECT 12.510 80.675 12.770 81.515 ;
        RECT 12.945 80.770 13.200 81.345 ;
        RECT 13.370 81.135 13.700 81.515 ;
        RECT 13.915 80.965 14.085 81.345 ;
        RECT 13.370 80.795 14.085 80.965 ;
        RECT 11.105 78.965 11.435 79.745 ;
        RECT 11.640 79.570 12.305 79.745 ;
        RECT 11.640 79.165 11.825 79.570 ;
        RECT 11.995 78.965 12.330 79.390 ;
        RECT 12.510 78.965 12.770 80.115 ;
        RECT 12.945 80.040 13.115 80.770 ;
        RECT 13.370 80.605 13.540 80.795 ;
        RECT 14.350 80.675 14.610 81.515 ;
        RECT 14.785 80.770 15.040 81.345 ;
        RECT 15.210 81.135 15.540 81.515 ;
        RECT 15.755 80.965 15.925 81.345 ;
        RECT 15.210 80.795 15.925 80.965 ;
        RECT 13.285 80.275 13.540 80.605 ;
        RECT 13.370 80.065 13.540 80.275 ;
        RECT 13.820 80.245 14.175 80.615 ;
        RECT 12.945 79.135 13.200 80.040 ;
        RECT 13.370 79.895 14.085 80.065 ;
        RECT 13.370 78.965 13.700 79.725 ;
        RECT 13.915 79.135 14.085 79.895 ;
        RECT 14.350 78.965 14.610 80.115 ;
        RECT 14.785 80.040 14.955 80.770 ;
        RECT 15.210 80.605 15.380 80.795 ;
        RECT 16.220 80.775 16.835 81.345 ;
        RECT 17.005 81.005 17.220 81.515 ;
        RECT 17.450 81.005 17.730 81.335 ;
        RECT 17.910 81.005 18.150 81.515 ;
        RECT 15.125 80.275 15.380 80.605 ;
        RECT 15.210 80.065 15.380 80.275 ;
        RECT 15.660 80.245 16.015 80.615 ;
        RECT 14.785 79.135 15.040 80.040 ;
        RECT 15.210 79.895 15.925 80.065 ;
        RECT 15.210 78.965 15.540 79.725 ;
        RECT 15.755 79.135 15.925 79.895 ;
        RECT 16.220 79.755 16.535 80.775 ;
        RECT 16.705 80.105 16.875 80.605 ;
        RECT 17.125 80.275 17.390 80.835 ;
        RECT 17.560 80.105 17.730 81.005 ;
        RECT 17.900 80.275 18.255 80.835 ;
        RECT 18.485 80.790 18.775 81.515 ;
        RECT 18.950 80.675 19.210 81.515 ;
        RECT 19.385 80.770 19.640 81.345 ;
        RECT 19.810 81.135 20.140 81.515 ;
        RECT 20.355 80.965 20.525 81.345 ;
        RECT 19.810 80.795 20.525 80.965 ;
        RECT 20.985 80.885 21.315 81.245 ;
        RECT 21.935 81.055 22.185 81.515 ;
        RECT 22.355 81.055 22.915 81.345 ;
        RECT 23.195 81.135 24.365 81.345 ;
        RECT 23.195 81.115 23.525 81.135 ;
        RECT 16.705 79.935 18.130 80.105 ;
        RECT 16.220 79.135 16.755 79.755 ;
        RECT 16.925 78.965 17.255 79.765 ;
        RECT 17.740 79.760 18.130 79.935 ;
        RECT 18.485 78.965 18.775 80.130 ;
        RECT 18.950 78.965 19.210 80.115 ;
        RECT 19.385 80.040 19.555 80.770 ;
        RECT 19.810 80.605 19.980 80.795 ;
        RECT 20.985 80.695 22.375 80.885 ;
        RECT 19.725 80.275 19.980 80.605 ;
        RECT 19.810 80.065 19.980 80.275 ;
        RECT 20.260 80.245 20.615 80.615 ;
        RECT 22.205 80.605 22.375 80.695 ;
        RECT 20.800 80.275 21.475 80.525 ;
        RECT 21.695 80.275 22.035 80.525 ;
        RECT 22.205 80.275 22.495 80.605 ;
        RECT 19.385 79.135 19.640 80.040 ;
        RECT 19.810 79.895 20.525 80.065 ;
        RECT 20.800 79.915 21.065 80.275 ;
        RECT 22.205 80.025 22.375 80.275 ;
        RECT 19.810 78.965 20.140 79.725 ;
        RECT 20.355 79.135 20.525 79.895 ;
        RECT 21.435 79.855 22.375 80.025 ;
        RECT 20.985 78.965 21.265 79.635 ;
        RECT 21.435 79.305 21.735 79.855 ;
        RECT 22.665 79.685 22.915 81.055 ;
        RECT 23.085 80.695 23.945 80.945 ;
        RECT 24.115 80.885 24.365 81.135 ;
        RECT 24.535 81.055 24.705 81.515 ;
        RECT 24.875 80.885 25.215 81.345 ;
        RECT 24.115 80.715 25.215 80.885 ;
        RECT 25.585 80.885 25.915 81.245 ;
        RECT 26.545 81.055 26.795 81.515 ;
        RECT 26.965 81.055 27.515 81.345 ;
        RECT 25.585 80.695 26.975 80.885 ;
        RECT 23.085 80.105 23.365 80.695 ;
        RECT 26.805 80.605 26.975 80.695 ;
        RECT 23.535 80.275 24.285 80.525 ;
        RECT 24.455 80.275 25.215 80.525 ;
        RECT 25.385 80.275 26.075 80.525 ;
        RECT 26.305 80.275 26.635 80.525 ;
        RECT 26.805 80.275 27.095 80.605 ;
        RECT 23.085 79.935 24.785 80.105 ;
        RECT 21.935 78.965 22.265 79.685 ;
        RECT 22.455 79.135 22.915 79.685 ;
        RECT 23.190 78.965 23.445 79.765 ;
        RECT 23.615 79.135 23.945 79.935 ;
        RECT 24.115 78.965 24.285 79.765 ;
        RECT 24.455 79.135 24.785 79.935 ;
        RECT 24.955 78.965 25.215 80.105 ;
        RECT 25.385 79.835 25.700 80.275 ;
        RECT 26.805 80.025 26.975 80.275 ;
        RECT 26.035 79.855 26.975 80.025 ;
        RECT 25.585 78.965 25.865 79.635 ;
        RECT 26.035 79.305 26.335 79.855 ;
        RECT 27.265 79.685 27.515 81.055 ;
        RECT 27.685 80.715 27.975 81.515 ;
        RECT 28.155 80.790 28.485 81.300 ;
        RECT 28.655 81.115 28.985 81.515 ;
        RECT 30.035 80.945 30.365 81.285 ;
        RECT 30.535 81.115 30.865 81.515 ;
        RECT 26.545 78.965 26.875 79.685 ;
        RECT 27.065 79.135 27.515 79.685 ;
        RECT 27.685 78.965 27.975 80.105 ;
        RECT 28.155 80.025 28.345 80.790 ;
        RECT 28.655 80.775 31.020 80.945 ;
        RECT 31.365 80.790 31.655 81.515 ;
        RECT 32.835 81.035 33.135 81.515 ;
        RECT 33.305 80.865 33.565 81.320 ;
        RECT 33.735 81.035 33.995 81.515 ;
        RECT 34.175 80.865 34.435 81.320 ;
        RECT 34.605 81.035 34.855 81.515 ;
        RECT 35.035 80.865 35.295 81.320 ;
        RECT 35.465 81.035 35.715 81.515 ;
        RECT 35.895 80.865 36.155 81.320 ;
        RECT 36.325 81.035 36.570 81.515 ;
        RECT 36.740 80.865 37.015 81.320 ;
        RECT 37.185 81.035 37.430 81.515 ;
        RECT 37.600 80.865 37.860 81.320 ;
        RECT 38.030 81.035 38.290 81.515 ;
        RECT 38.460 80.865 38.720 81.320 ;
        RECT 38.890 81.035 39.150 81.515 ;
        RECT 39.320 80.865 39.580 81.320 ;
        RECT 39.750 80.955 40.010 81.515 ;
        RECT 28.655 80.605 28.825 80.775 ;
        RECT 28.515 80.275 28.825 80.605 ;
        RECT 28.995 80.275 29.300 80.605 ;
        RECT 28.155 79.175 28.485 80.025 ;
        RECT 28.655 78.965 28.905 80.105 ;
        RECT 29.085 79.945 29.300 80.275 ;
        RECT 29.475 79.945 29.760 80.605 ;
        RECT 29.955 79.945 30.220 80.605 ;
        RECT 30.435 79.945 30.680 80.605 ;
        RECT 30.850 79.775 31.020 80.775 ;
        RECT 32.835 80.695 39.580 80.865 ;
        RECT 32.835 80.155 34.000 80.695 ;
        RECT 40.180 80.525 40.430 81.335 ;
        RECT 40.610 80.990 40.870 81.515 ;
        RECT 41.040 80.525 41.290 81.335 ;
        RECT 41.470 81.005 41.775 81.515 ;
        RECT 41.945 80.840 42.205 81.345 ;
        RECT 42.385 81.135 42.715 81.515 ;
        RECT 42.895 80.965 43.065 81.345 ;
        RECT 34.170 80.275 41.290 80.525 ;
        RECT 41.460 80.275 41.775 80.835 ;
        RECT 29.095 79.605 30.385 79.775 ;
        RECT 29.095 79.185 29.345 79.605 ;
        RECT 29.575 78.965 29.905 79.435 ;
        RECT 30.135 79.185 30.385 79.605 ;
        RECT 30.565 79.605 31.020 79.775 ;
        RECT 30.565 79.175 30.895 79.605 ;
        RECT 31.365 78.965 31.655 80.130 ;
        RECT 32.805 80.105 34.000 80.155 ;
        RECT 32.805 79.985 39.580 80.105 ;
        RECT 32.835 79.880 39.580 79.985 ;
        RECT 32.835 78.965 33.105 79.710 ;
        RECT 33.275 79.140 33.565 79.880 ;
        RECT 34.175 79.865 39.580 79.880 ;
        RECT 33.735 78.970 33.990 79.695 ;
        RECT 34.175 79.140 34.435 79.865 ;
        RECT 34.605 78.970 34.850 79.695 ;
        RECT 35.035 79.140 35.295 79.865 ;
        RECT 35.465 78.970 35.710 79.695 ;
        RECT 35.895 79.140 36.155 79.865 ;
        RECT 36.325 78.970 36.570 79.695 ;
        RECT 36.740 79.140 37.000 79.865 ;
        RECT 37.170 78.970 37.430 79.695 ;
        RECT 37.600 79.140 37.860 79.865 ;
        RECT 38.030 78.970 38.290 79.695 ;
        RECT 38.460 79.140 38.720 79.865 ;
        RECT 38.890 78.970 39.150 79.695 ;
        RECT 39.320 79.140 39.580 79.865 ;
        RECT 39.750 78.970 40.010 79.765 ;
        RECT 40.180 79.140 40.430 80.275 ;
        RECT 33.735 78.965 40.010 78.970 ;
        RECT 40.610 78.965 40.870 79.775 ;
        RECT 41.045 79.135 41.290 80.275 ;
        RECT 41.945 80.040 42.115 80.840 ;
        RECT 42.400 80.795 43.065 80.965 ;
        RECT 42.400 80.540 42.570 80.795 ;
        RECT 44.245 80.790 44.535 81.515 ;
        RECT 45.035 81.115 45.365 81.515 ;
        RECT 45.535 80.945 45.865 81.285 ;
        RECT 46.915 81.115 47.245 81.515 ;
        RECT 44.880 80.775 47.245 80.945 ;
        RECT 47.415 80.790 47.745 81.300 ;
        RECT 48.015 81.035 48.315 81.515 ;
        RECT 48.485 80.865 48.745 81.320 ;
        RECT 48.915 81.035 49.175 81.515 ;
        RECT 49.355 80.865 49.615 81.320 ;
        RECT 49.785 81.035 50.035 81.515 ;
        RECT 50.215 80.865 50.475 81.320 ;
        RECT 50.645 81.035 50.895 81.515 ;
        RECT 51.075 80.865 51.335 81.320 ;
        RECT 51.505 81.035 51.750 81.515 ;
        RECT 51.920 80.865 52.195 81.320 ;
        RECT 52.365 81.035 52.610 81.515 ;
        RECT 52.780 80.865 53.040 81.320 ;
        RECT 53.210 81.035 53.470 81.515 ;
        RECT 53.640 80.865 53.900 81.320 ;
        RECT 54.070 81.035 54.330 81.515 ;
        RECT 54.500 80.865 54.760 81.320 ;
        RECT 54.930 80.955 55.190 81.515 ;
        RECT 42.285 80.210 42.570 80.540 ;
        RECT 42.805 80.245 43.135 80.615 ;
        RECT 42.400 80.065 42.570 80.210 ;
        RECT 41.470 78.965 41.765 79.775 ;
        RECT 41.945 79.135 42.215 80.040 ;
        RECT 42.400 79.895 43.065 80.065 ;
        RECT 42.385 78.965 42.715 79.725 ;
        RECT 42.895 79.135 43.065 79.895 ;
        RECT 44.245 78.965 44.535 80.130 ;
        RECT 44.880 79.775 45.050 80.775 ;
        RECT 47.075 80.605 47.245 80.775 ;
        RECT 45.220 79.945 45.465 80.605 ;
        RECT 45.680 79.945 45.945 80.605 ;
        RECT 46.140 79.945 46.425 80.605 ;
        RECT 46.600 80.275 46.905 80.605 ;
        RECT 47.075 80.275 47.385 80.605 ;
        RECT 46.600 79.945 46.815 80.275 ;
        RECT 44.880 79.605 45.335 79.775 ;
        RECT 45.005 79.175 45.335 79.605 ;
        RECT 45.515 79.605 46.805 79.775 ;
        RECT 45.515 79.185 45.765 79.605 ;
        RECT 45.995 78.965 46.325 79.435 ;
        RECT 46.555 79.185 46.805 79.605 ;
        RECT 46.995 78.965 47.245 80.105 ;
        RECT 47.555 80.025 47.745 80.790 ;
        RECT 47.415 79.175 47.745 80.025 ;
        RECT 48.015 80.695 54.760 80.865 ;
        RECT 48.015 80.105 49.180 80.695 ;
        RECT 55.360 80.525 55.610 81.335 ;
        RECT 55.790 80.990 56.050 81.515 ;
        RECT 56.220 80.525 56.470 81.335 ;
        RECT 56.650 81.005 56.955 81.515 ;
        RECT 49.350 80.275 56.470 80.525 ;
        RECT 56.640 80.275 56.955 80.835 ;
        RECT 57.125 80.790 57.415 81.515 ;
        RECT 57.585 80.865 57.845 81.310 ;
        RECT 58.095 81.035 58.265 81.515 ;
        RECT 58.435 81.005 58.785 81.335 ;
        RECT 59.020 81.035 59.190 81.515 ;
        RECT 57.585 80.695 58.265 80.865 ;
        RECT 48.015 79.880 54.760 80.105 ;
        RECT 48.015 78.965 48.285 79.710 ;
        RECT 48.455 79.140 48.745 79.880 ;
        RECT 49.355 79.865 54.760 79.880 ;
        RECT 48.915 78.970 49.170 79.695 ;
        RECT 49.355 79.140 49.615 79.865 ;
        RECT 49.785 78.970 50.030 79.695 ;
        RECT 50.215 79.140 50.475 79.865 ;
        RECT 50.645 78.970 50.890 79.695 ;
        RECT 51.075 79.140 51.335 79.865 ;
        RECT 51.505 78.970 51.750 79.695 ;
        RECT 51.920 79.140 52.180 79.865 ;
        RECT 52.350 78.970 52.610 79.695 ;
        RECT 52.780 79.140 53.040 79.865 ;
        RECT 53.210 78.970 53.470 79.695 ;
        RECT 53.640 79.140 53.900 79.865 ;
        RECT 54.070 78.970 54.330 79.695 ;
        RECT 54.500 79.140 54.760 79.865 ;
        RECT 54.930 78.970 55.190 79.765 ;
        RECT 55.360 79.140 55.610 80.275 ;
        RECT 48.915 78.965 55.190 78.970 ;
        RECT 55.790 78.965 56.050 79.775 ;
        RECT 56.225 79.135 56.470 80.275 ;
        RECT 56.650 78.965 56.945 79.775 ;
        RECT 57.125 78.965 57.415 80.130 ;
        RECT 57.585 79.960 57.925 80.525 ;
        RECT 58.095 79.790 58.265 80.695 ;
        RECT 58.435 80.105 58.605 81.005 ;
        RECT 59.490 80.945 59.660 81.295 ;
        RECT 59.830 81.115 60.160 81.515 ;
        RECT 60.330 80.995 60.585 81.295 ;
        RECT 60.805 81.005 61.110 81.515 ;
        RECT 60.330 80.945 60.635 80.995 ;
        RECT 59.490 80.865 60.635 80.945 ;
        RECT 58.925 80.835 60.635 80.865 ;
        RECT 58.775 80.775 60.635 80.835 ;
        RECT 58.775 80.695 59.660 80.775 ;
        RECT 58.775 80.665 59.095 80.695 ;
        RECT 58.775 80.275 58.945 80.665 ;
        RECT 58.435 79.900 58.830 80.105 ;
        RECT 59.195 79.985 59.730 80.525 ;
        RECT 59.990 80.275 60.290 80.605 ;
        RECT 59.990 79.815 60.160 80.275 ;
        RECT 60.465 80.105 60.635 80.775 ;
        RECT 60.805 80.275 61.120 80.835 ;
        RECT 61.290 80.525 61.540 81.335 ;
        RECT 61.710 80.990 61.970 81.515 ;
        RECT 62.150 80.525 62.400 81.335 ;
        RECT 62.570 80.955 62.830 81.515 ;
        RECT 63.000 80.865 63.260 81.320 ;
        RECT 63.430 81.035 63.690 81.515 ;
        RECT 63.860 80.865 64.120 81.320 ;
        RECT 64.290 81.035 64.550 81.515 ;
        RECT 64.720 80.865 64.980 81.320 ;
        RECT 65.150 81.035 65.395 81.515 ;
        RECT 65.565 80.865 65.840 81.320 ;
        RECT 66.010 81.035 66.255 81.515 ;
        RECT 66.425 80.865 66.685 81.320 ;
        RECT 66.865 81.035 67.115 81.515 ;
        RECT 67.285 80.865 67.545 81.320 ;
        RECT 67.725 81.035 67.975 81.515 ;
        RECT 68.145 80.865 68.405 81.320 ;
        RECT 68.585 81.035 68.845 81.515 ;
        RECT 69.015 80.865 69.275 81.320 ;
        RECT 69.445 81.035 69.745 81.515 ;
        RECT 63.000 80.695 69.745 80.865 ;
        RECT 70.005 80.790 70.295 81.515 ;
        RECT 70.465 80.905 70.815 81.345 ;
        RECT 70.985 81.075 71.155 81.515 ;
        RECT 71.325 81.135 72.520 81.345 ;
        RECT 71.325 80.905 71.575 81.135 ;
        RECT 70.465 80.695 71.575 80.905 ;
        RECT 71.745 80.795 72.075 80.965 ;
        RECT 71.745 80.695 72.070 80.795 ;
        RECT 72.245 80.695 72.520 81.135 ;
        RECT 72.755 80.775 73.085 81.515 ;
        RECT 73.255 80.760 73.490 81.090 ;
        RECT 73.775 80.965 73.945 81.345 ;
        RECT 74.160 81.135 74.490 81.515 ;
        RECT 73.775 80.795 74.490 80.965 ;
        RECT 61.290 80.275 68.410 80.525 ;
        RECT 57.585 79.730 58.265 79.790 ;
        RECT 59.050 79.730 60.160 79.815 ;
        RECT 57.585 79.645 60.160 79.730 ;
        RECT 60.330 79.675 60.635 80.105 ;
        RECT 57.585 79.560 59.220 79.645 ;
        RECT 57.585 79.380 57.845 79.560 ;
        RECT 58.050 78.965 58.410 79.390 ;
        RECT 58.925 78.965 59.255 79.390 ;
        RECT 59.435 79.235 60.635 79.475 ;
        RECT 60.815 78.965 61.110 79.775 ;
        RECT 61.290 79.135 61.535 80.275 ;
        RECT 61.710 78.965 61.970 79.775 ;
        RECT 62.150 79.140 62.400 80.275 ;
        RECT 68.580 80.105 69.745 80.695 ;
        RECT 70.465 80.325 71.610 80.525 ;
        RECT 71.420 80.155 71.610 80.325 ;
        RECT 63.000 79.880 69.745 80.105 ;
        RECT 63.000 79.865 68.405 79.880 ;
        RECT 62.570 78.970 62.830 79.765 ;
        RECT 63.000 79.140 63.260 79.865 ;
        RECT 63.430 78.970 63.690 79.695 ;
        RECT 63.860 79.140 64.120 79.865 ;
        RECT 64.290 78.970 64.550 79.695 ;
        RECT 64.720 79.140 64.980 79.865 ;
        RECT 65.150 78.970 65.410 79.695 ;
        RECT 65.580 79.140 65.840 79.865 ;
        RECT 66.010 78.970 66.255 79.695 ;
        RECT 66.425 79.140 66.685 79.865 ;
        RECT 66.870 78.970 67.115 79.695 ;
        RECT 67.285 79.140 67.545 79.865 ;
        RECT 67.730 78.970 67.975 79.695 ;
        RECT 68.145 79.140 68.405 79.865 ;
        RECT 68.590 78.970 68.845 79.695 ;
        RECT 69.015 79.140 69.305 79.880 ;
        RECT 62.570 78.965 68.845 78.970 ;
        RECT 69.475 78.965 69.745 79.710 ;
        RECT 70.005 78.965 70.295 80.130 ;
        RECT 70.985 80.105 71.155 80.155 ;
        RECT 70.465 78.965 70.795 80.105 ;
        RECT 70.965 79.765 71.240 80.105 ;
        RECT 71.420 79.985 71.615 80.155 ;
        RECT 71.420 79.945 71.610 79.985 ;
        RECT 71.790 79.765 72.070 80.695 ;
        RECT 72.240 80.105 72.570 80.525 ;
        RECT 72.800 80.275 73.145 80.605 ;
        RECT 73.320 80.105 73.490 80.760 ;
        RECT 73.685 80.245 74.040 80.615 ;
        RECT 74.320 80.605 74.490 80.795 ;
        RECT 74.660 80.770 74.915 81.345 ;
        RECT 74.320 80.275 74.575 80.605 ;
        RECT 72.240 79.935 73.490 80.105 ;
        RECT 74.320 80.065 74.490 80.275 ;
        RECT 70.965 79.595 72.565 79.765 ;
        RECT 70.965 79.135 71.320 79.595 ;
        RECT 71.490 78.965 72.065 79.425 ;
        RECT 72.235 79.135 72.565 79.595 ;
        RECT 72.765 78.965 73.020 79.765 ;
        RECT 73.190 79.740 73.490 79.935 ;
        RECT 73.775 79.895 74.490 80.065 ;
        RECT 74.745 80.040 74.915 80.770 ;
        RECT 75.090 80.675 75.350 81.515 ;
        RECT 75.525 80.765 76.735 81.515 ;
        RECT 73.775 79.135 73.945 79.895 ;
        RECT 74.160 78.965 74.490 79.725 ;
        RECT 74.660 79.135 74.915 80.040 ;
        RECT 75.090 78.965 75.350 80.115 ;
        RECT 75.525 80.055 76.045 80.595 ;
        RECT 76.215 80.225 76.735 80.765 ;
        RECT 75.525 78.965 76.735 80.055 ;
        RECT 5.520 78.795 76.820 78.965 ;
        RECT 5.605 77.705 6.815 78.795 ;
        RECT 5.605 76.995 6.125 77.535 ;
        RECT 6.295 77.165 6.815 77.705 ;
        RECT 7.905 78.075 8.365 78.625 ;
        RECT 8.555 78.075 8.885 78.795 ;
        RECT 5.605 76.245 6.815 76.995 ;
        RECT 7.905 76.705 8.155 78.075 ;
        RECT 9.085 77.905 9.385 78.455 ;
        RECT 9.555 78.125 9.835 78.795 ;
        RECT 8.445 77.735 9.385 77.905 ;
        RECT 8.445 77.485 8.615 77.735 ;
        RECT 9.755 77.485 10.020 77.845 ;
        RECT 11.125 77.655 11.405 78.795 ;
        RECT 11.575 77.645 11.905 78.625 ;
        RECT 12.075 77.655 12.335 78.795 ;
        RECT 12.505 77.655 12.785 78.795 ;
        RECT 12.955 77.645 13.285 78.625 ;
        RECT 13.455 77.655 13.715 78.795 ;
        RECT 14.345 77.735 14.660 78.795 ;
        RECT 15.290 78.290 15.905 78.795 ;
        RECT 8.325 77.155 8.615 77.485 ;
        RECT 8.785 77.235 9.125 77.485 ;
        RECT 9.345 77.235 10.020 77.485 ;
        RECT 11.135 77.215 11.470 77.485 ;
        RECT 8.445 77.065 8.615 77.155 ;
        RECT 8.445 76.875 9.835 77.065 ;
        RECT 11.640 77.045 11.810 77.645 ;
        RECT 11.980 77.235 12.315 77.485 ;
        RECT 12.515 77.215 12.850 77.485 ;
        RECT 13.020 77.045 13.190 77.645 ;
        RECT 13.360 77.235 13.695 77.485 ;
        RECT 7.905 76.415 8.465 76.705 ;
        RECT 8.635 76.245 8.885 76.705 ;
        RECT 9.505 76.515 9.835 76.875 ;
        RECT 11.125 76.245 11.435 77.045 ;
        RECT 11.640 76.415 12.335 77.045 ;
        RECT 12.505 76.245 12.815 77.045 ;
        RECT 13.020 76.415 13.715 77.045 ;
        RECT 14.405 76.905 14.670 77.485 ;
        RECT 14.840 77.405 15.115 78.065 ;
        RECT 15.310 77.755 15.545 78.120 ;
        RECT 15.715 78.115 15.905 78.290 ;
        RECT 16.075 78.285 16.550 78.625 ;
        RECT 15.715 77.925 16.045 78.115 ;
        RECT 16.270 77.755 16.460 78.050 ;
        RECT 16.720 77.950 16.935 78.795 ;
        RECT 17.135 77.955 17.420 78.625 ;
        RECT 15.310 77.585 17.080 77.755 ;
        RECT 14.840 77.175 15.675 77.405 ;
        RECT 14.345 76.245 14.615 76.735 ;
        RECT 14.840 76.465 15.115 77.175 ;
        RECT 15.845 76.730 16.100 77.585 ;
        RECT 15.315 76.465 16.100 76.730 ;
        RECT 16.270 76.925 16.680 77.405 ;
        RECT 16.850 77.155 17.080 77.585 ;
        RECT 17.250 77.605 17.420 77.955 ;
        RECT 17.590 77.785 17.855 78.795 ;
        RECT 18.485 77.630 18.775 78.795 ;
        RECT 19.410 77.650 19.705 78.795 ;
        RECT 17.250 77.085 17.855 77.605 ;
        RECT 16.270 76.465 16.480 76.925 ;
        RECT 17.250 76.875 17.420 77.085 ;
        RECT 16.670 76.245 17.000 76.740 ;
        RECT 17.175 76.415 17.420 76.875 ;
        RECT 17.590 76.245 17.855 76.905 ;
        RECT 18.485 76.245 18.775 76.970 ;
        RECT 19.410 76.245 19.705 77.065 ;
        RECT 19.875 76.795 20.105 78.495 ;
        RECT 20.320 77.990 20.575 78.795 ;
        RECT 20.775 78.180 21.105 78.625 ;
        RECT 21.275 78.350 21.550 78.795 ;
        RECT 21.785 78.180 22.115 78.625 ;
        RECT 20.775 78.000 22.115 78.180 ;
        RECT 22.575 77.820 22.905 78.485 ;
        RECT 23.105 77.995 23.435 78.795 ;
        RECT 20.320 77.650 22.905 77.820 ;
        RECT 23.610 77.655 23.945 78.625 ;
        RECT 24.115 77.995 24.445 78.795 ;
        RECT 24.845 77.825 25.095 78.625 ;
        RECT 25.280 78.075 25.610 78.795 ;
        RECT 25.830 77.825 26.080 78.625 ;
        RECT 26.255 78.415 26.585 78.795 ;
        RECT 24.125 77.655 26.180 77.825 ;
        RECT 20.320 77.035 20.630 77.650 ;
        RECT 23.610 77.435 23.785 77.655 ;
        RECT 24.125 77.475 24.350 77.655 ;
        RECT 20.800 77.205 21.130 77.435 ;
        RECT 21.300 77.205 21.770 77.435 ;
        RECT 21.940 77.265 22.395 77.435 ;
        RECT 21.940 77.205 22.390 77.265 ;
        RECT 22.580 77.205 22.915 77.435 ;
        RECT 23.605 77.265 23.785 77.435 ;
        RECT 20.320 76.855 22.905 77.035 ;
        RECT 19.875 76.415 20.095 76.795 ;
        RECT 20.265 76.245 21.115 76.605 ;
        RECT 21.595 76.435 21.925 76.855 ;
        RECT 22.130 76.245 22.405 76.685 ;
        RECT 22.575 76.435 22.905 76.855 ;
        RECT 23.095 76.245 23.425 76.970 ;
        RECT 23.610 76.965 23.785 77.265 ;
        RECT 23.955 77.235 24.350 77.475 ;
        RECT 23.610 76.500 23.945 76.965 ;
        RECT 23.615 76.455 23.945 76.500 ;
        RECT 24.115 76.245 24.350 77.050 ;
        RECT 24.520 76.575 24.780 77.485 ;
        RECT 25.090 77.465 25.260 77.485 ;
        RECT 24.960 76.575 25.260 77.465 ;
        RECT 25.435 76.580 25.790 77.485 ;
        RECT 26.010 76.745 26.180 77.655 ;
        RECT 26.350 76.915 26.555 78.235 ;
        RECT 26.855 78.050 27.125 78.795 ;
        RECT 27.755 78.790 34.030 78.795 ;
        RECT 27.295 77.880 27.585 78.620 ;
        RECT 27.755 78.065 28.010 78.790 ;
        RECT 28.195 77.895 28.455 78.620 ;
        RECT 28.625 78.065 28.870 78.790 ;
        RECT 29.055 77.895 29.315 78.620 ;
        RECT 29.485 78.065 29.730 78.790 ;
        RECT 29.915 77.895 30.175 78.620 ;
        RECT 30.345 78.065 30.590 78.790 ;
        RECT 30.760 77.895 31.020 78.620 ;
        RECT 31.190 78.065 31.450 78.790 ;
        RECT 31.620 77.895 31.880 78.620 ;
        RECT 32.050 78.065 32.310 78.790 ;
        RECT 32.480 77.895 32.740 78.620 ;
        RECT 32.910 78.065 33.170 78.790 ;
        RECT 33.340 77.895 33.600 78.620 ;
        RECT 33.770 77.995 34.030 78.790 ;
        RECT 28.195 77.880 33.600 77.895 ;
        RECT 26.855 77.655 33.600 77.880 ;
        RECT 26.855 77.065 28.020 77.655 ;
        RECT 34.200 77.485 34.450 78.620 ;
        RECT 34.630 77.985 34.890 78.795 ;
        RECT 35.065 77.485 35.310 78.625 ;
        RECT 35.490 77.985 35.785 78.795 ;
        RECT 36.055 77.785 36.225 78.625 ;
        RECT 36.395 78.455 37.565 78.625 ;
        RECT 36.395 77.955 36.725 78.455 ;
        RECT 37.235 78.415 37.565 78.455 ;
        RECT 37.755 78.375 38.110 78.795 ;
        RECT 36.895 78.195 37.125 78.285 ;
        RECT 38.280 78.195 38.530 78.625 ;
        RECT 36.895 77.955 38.530 78.195 ;
        RECT 38.700 78.035 39.030 78.795 ;
        RECT 39.200 77.955 39.455 78.625 ;
        RECT 36.055 77.615 39.115 77.785 ;
        RECT 28.190 77.235 35.310 77.485 ;
        RECT 26.855 76.895 33.600 77.065 ;
        RECT 26.010 76.415 26.505 76.745 ;
        RECT 26.855 76.245 27.155 76.725 ;
        RECT 27.325 76.440 27.585 76.895 ;
        RECT 27.755 76.245 28.015 76.725 ;
        RECT 28.195 76.440 28.455 76.895 ;
        RECT 28.625 76.245 28.875 76.725 ;
        RECT 29.055 76.440 29.315 76.895 ;
        RECT 29.485 76.245 29.735 76.725 ;
        RECT 29.915 76.440 30.175 76.895 ;
        RECT 30.345 76.245 30.590 76.725 ;
        RECT 30.760 76.440 31.035 76.895 ;
        RECT 31.205 76.245 31.450 76.725 ;
        RECT 31.620 76.440 31.880 76.895 ;
        RECT 32.050 76.245 32.310 76.725 ;
        RECT 32.480 76.440 32.740 76.895 ;
        RECT 32.910 76.245 33.170 76.725 ;
        RECT 33.340 76.440 33.600 76.895 ;
        RECT 33.770 76.245 34.030 76.805 ;
        RECT 34.200 76.425 34.450 77.235 ;
        RECT 34.630 76.245 34.890 76.770 ;
        RECT 35.060 76.425 35.310 77.235 ;
        RECT 35.480 76.925 35.795 77.485 ;
        RECT 35.965 77.235 36.320 77.445 ;
        RECT 36.490 77.235 36.935 77.435 ;
        RECT 37.105 77.235 37.580 77.435 ;
        RECT 36.055 76.895 37.120 77.065 ;
        RECT 35.490 76.245 35.795 76.755 ;
        RECT 36.055 76.415 36.225 76.895 ;
        RECT 36.395 76.245 36.725 76.725 ;
        RECT 36.950 76.665 37.120 76.895 ;
        RECT 37.300 76.835 37.580 77.235 ;
        RECT 37.850 77.235 38.180 77.435 ;
        RECT 38.350 77.235 38.715 77.435 ;
        RECT 37.850 76.835 38.135 77.235 ;
        RECT 38.945 77.065 39.115 77.615 ;
        RECT 38.315 76.895 39.115 77.065 ;
        RECT 38.315 76.665 38.485 76.895 ;
        RECT 39.285 76.825 39.455 77.955 ;
        RECT 39.625 77.605 39.795 78.795 ;
        RECT 40.115 77.820 40.445 78.485 ;
        RECT 40.905 78.180 41.235 78.625 ;
        RECT 41.470 78.350 41.745 78.795 ;
        RECT 41.915 78.180 42.245 78.625 ;
        RECT 40.905 78.000 42.245 78.180 ;
        RECT 42.445 77.990 42.700 78.795 ;
        RECT 40.115 77.650 42.700 77.820 ;
        RECT 40.105 77.205 40.440 77.435 ;
        RECT 40.625 77.265 41.080 77.435 ;
        RECT 40.630 77.205 41.080 77.265 ;
        RECT 41.250 77.205 41.720 77.435 ;
        RECT 41.890 77.205 42.220 77.435 ;
        RECT 39.270 76.755 39.455 76.825 ;
        RECT 39.245 76.745 39.455 76.755 ;
        RECT 36.950 76.415 38.485 76.665 ;
        RECT 38.655 76.245 38.985 76.725 ;
        RECT 39.200 76.415 39.455 76.745 ;
        RECT 39.625 76.245 39.795 77.140 ;
        RECT 42.390 77.035 42.700 77.650 ;
        RECT 40.115 76.855 42.700 77.035 ;
        RECT 40.115 76.435 40.445 76.855 ;
        RECT 40.615 76.245 40.890 76.685 ;
        RECT 41.095 76.435 41.425 76.855 ;
        RECT 42.915 76.795 43.145 78.495 ;
        RECT 43.315 77.650 43.610 78.795 ;
        RECT 44.245 77.630 44.535 78.795 ;
        RECT 44.760 77.925 45.045 78.795 ;
        RECT 45.215 78.165 45.475 78.625 ;
        RECT 45.650 78.335 45.905 78.795 ;
        RECT 46.075 78.165 46.335 78.625 ;
        RECT 45.215 77.995 46.335 78.165 ;
        RECT 46.505 77.995 46.815 78.795 ;
        RECT 45.215 77.745 45.475 77.995 ;
        RECT 46.985 77.825 47.295 78.625 ;
        RECT 47.465 78.200 47.900 78.625 ;
        RECT 48.070 78.370 48.455 78.795 ;
        RECT 47.465 78.030 48.455 78.200 ;
        RECT 44.720 77.575 45.475 77.745 ;
        RECT 46.265 77.655 47.295 77.825 ;
        RECT 44.720 77.065 45.125 77.575 ;
        RECT 46.265 77.405 46.435 77.655 ;
        RECT 45.295 77.235 46.435 77.405 ;
        RECT 41.905 76.245 42.755 76.605 ;
        RECT 42.925 76.415 43.145 76.795 ;
        RECT 43.315 76.245 43.610 77.065 ;
        RECT 44.245 76.245 44.535 76.970 ;
        RECT 44.720 76.895 46.370 77.065 ;
        RECT 46.605 76.915 46.955 77.485 ;
        RECT 44.765 76.245 45.045 76.725 ;
        RECT 45.215 76.505 45.475 76.895 ;
        RECT 45.650 76.245 45.905 76.725 ;
        RECT 46.075 76.505 46.370 76.895 ;
        RECT 47.125 76.745 47.295 77.655 ;
        RECT 47.465 77.155 47.950 77.860 ;
        RECT 48.120 77.485 48.455 78.030 ;
        RECT 48.625 77.835 49.050 78.625 ;
        RECT 49.220 78.200 49.495 78.625 ;
        RECT 49.665 78.370 50.050 78.795 ;
        RECT 49.220 78.005 50.050 78.200 ;
        RECT 48.625 77.655 49.530 77.835 ;
        RECT 48.120 77.155 48.530 77.485 ;
        RECT 48.700 77.155 49.530 77.655 ;
        RECT 49.700 77.485 50.050 78.005 ;
        RECT 50.220 77.835 50.465 78.625 ;
        RECT 50.655 78.200 50.910 78.625 ;
        RECT 51.080 78.370 51.465 78.795 ;
        RECT 50.655 78.005 51.465 78.200 ;
        RECT 50.220 77.655 50.945 77.835 ;
        RECT 49.700 77.155 50.125 77.485 ;
        RECT 50.295 77.155 50.945 77.655 ;
        RECT 51.115 77.485 51.465 78.005 ;
        RECT 51.635 77.655 51.895 78.625 ;
        RECT 52.135 77.825 52.495 78.625 ;
        RECT 53.040 77.995 53.210 78.795 ;
        RECT 53.420 78.165 53.750 78.625 ;
        RECT 53.920 78.335 54.090 78.795 ;
        RECT 54.260 78.165 54.590 78.625 ;
        RECT 53.420 77.995 54.590 78.165 ;
        RECT 54.760 77.995 54.930 78.795 ;
        RECT 54.260 77.825 54.590 77.995 ;
        RECT 52.135 77.655 53.595 77.825 ;
        RECT 54.260 77.655 55.115 77.825 ;
        RECT 55.285 77.705 56.495 78.795 ;
        RECT 51.115 77.155 51.540 77.485 ;
        RECT 48.120 76.985 48.455 77.155 ;
        RECT 48.700 76.985 49.050 77.155 ;
        RECT 49.700 76.985 50.050 77.155 ;
        RECT 50.295 76.985 50.465 77.155 ;
        RECT 51.115 76.985 51.465 77.155 ;
        RECT 51.710 76.985 51.895 77.655 ;
        RECT 46.550 76.245 46.825 76.725 ;
        RECT 46.995 76.415 47.295 76.745 ;
        RECT 47.465 76.815 48.455 76.985 ;
        RECT 47.465 76.415 47.900 76.815 ;
        RECT 48.070 76.245 48.455 76.645 ;
        RECT 48.625 76.415 49.050 76.985 ;
        RECT 49.240 76.815 50.050 76.985 ;
        RECT 49.240 76.415 49.495 76.815 ;
        RECT 49.665 76.245 50.050 76.645 ;
        RECT 50.220 76.415 50.465 76.985 ;
        RECT 50.655 76.815 51.465 76.985 ;
        RECT 50.655 76.415 50.910 76.815 ;
        RECT 51.080 76.245 51.465 76.645 ;
        RECT 51.635 76.415 51.895 76.985 ;
        RECT 52.070 76.925 52.325 77.485 ;
        RECT 52.495 76.985 52.675 77.655 ;
        RECT 52.845 77.155 53.220 77.485 ;
        RECT 53.390 77.405 53.595 77.655 ;
        RECT 53.390 77.235 54.600 77.405 ;
        RECT 54.770 77.065 55.115 77.655 ;
        RECT 52.085 76.245 52.325 76.755 ;
        RECT 52.495 76.450 52.825 76.985 ;
        RECT 53.040 76.245 53.210 76.985 ;
        RECT 53.420 76.895 55.115 77.065 ;
        RECT 55.285 76.995 55.805 77.535 ;
        RECT 55.975 77.165 56.495 77.705 ;
        RECT 56.725 77.655 56.935 78.795 ;
        RECT 57.105 77.645 57.435 78.625 ;
        RECT 57.605 77.655 57.835 78.795 ;
        RECT 58.095 78.335 58.345 78.795 ;
        RECT 58.555 78.165 58.725 78.625 ;
        RECT 58.050 77.995 58.725 78.165 ;
        RECT 58.895 77.995 59.145 78.795 ;
        RECT 59.315 78.165 59.565 78.585 ;
        RECT 59.775 78.335 60.105 78.795 ;
        RECT 60.295 78.165 60.545 78.585 ;
        RECT 59.315 77.995 60.605 78.165 ;
        RECT 53.420 76.425 53.750 76.895 ;
        RECT 53.920 76.245 54.090 76.725 ;
        RECT 54.260 76.425 54.590 76.895 ;
        RECT 54.760 76.245 54.930 76.725 ;
        RECT 55.285 76.245 56.495 76.995 ;
        RECT 56.725 76.245 56.935 77.065 ;
        RECT 57.105 77.045 57.355 77.645 ;
        RECT 57.525 77.235 57.855 77.485 ;
        RECT 57.105 76.415 57.435 77.045 ;
        RECT 57.605 76.245 57.835 77.065 ;
        RECT 58.050 77.045 58.305 77.995 ;
        RECT 60.835 77.825 61.005 78.625 ;
        RECT 58.515 77.655 61.005 77.825 ;
        RECT 58.515 77.405 58.685 77.655 ;
        RECT 58.515 77.235 58.845 77.405 ;
        RECT 59.025 77.155 59.355 77.485 ;
        RECT 59.585 77.405 59.755 77.420 ;
        RECT 59.585 77.235 59.915 77.405 ;
        RECT 58.050 76.875 58.725 77.045 ;
        RECT 59.025 76.920 59.230 77.155 ;
        RECT 59.585 77.025 59.755 77.235 ;
        RECT 60.145 77.030 60.315 77.485 ;
        RECT 58.050 76.245 58.305 76.705 ;
        RECT 58.555 76.415 58.725 76.875 ;
        RECT 59.490 76.855 59.755 77.025 ;
        RECT 59.925 76.860 60.315 77.030 ;
        RECT 59.490 76.755 59.660 76.855 ;
        RECT 58.975 76.625 59.145 76.705 ;
        RECT 58.915 76.245 59.245 76.625 ;
        RECT 59.485 76.585 59.660 76.755 ;
        RECT 59.490 76.560 59.660 76.585 ;
        RECT 59.925 76.575 60.135 76.860 ;
        RECT 60.495 76.665 60.665 77.655 ;
        RECT 60.855 76.915 61.050 77.485 ;
        RECT 60.335 76.495 60.665 76.665 ;
        RECT 60.420 76.415 60.665 76.495 ;
        RECT 60.835 76.245 61.095 76.725 ;
        RECT 61.280 76.425 61.560 78.615 ;
        RECT 61.750 77.655 62.035 78.795 ;
        RECT 62.300 78.145 62.470 78.615 ;
        RECT 62.645 78.315 62.975 78.795 ;
        RECT 63.145 78.145 63.325 78.615 ;
        RECT 62.300 77.945 63.325 78.145 ;
        RECT 61.760 76.975 62.020 77.485 ;
        RECT 62.230 77.155 62.490 77.775 ;
        RECT 62.685 77.155 63.110 77.775 ;
        RECT 63.495 77.505 63.825 78.615 ;
        RECT 63.995 78.385 64.345 78.795 ;
        RECT 64.515 78.205 64.755 78.595 ;
        RECT 63.280 77.205 63.825 77.505 ;
        RECT 64.005 78.005 64.755 78.205 ;
        RECT 64.965 78.205 65.205 78.595 ;
        RECT 65.375 78.385 65.725 78.795 ;
        RECT 64.965 78.005 65.715 78.205 ;
        RECT 64.005 77.325 64.345 78.005 ;
        RECT 63.280 76.975 63.500 77.205 ;
        RECT 61.760 76.785 63.500 76.975 ;
        RECT 61.760 76.245 62.490 76.615 ;
        RECT 63.070 76.425 63.500 76.785 ;
        RECT 63.670 76.245 63.915 77.025 ;
        RECT 64.115 76.425 64.345 77.325 ;
        RECT 64.525 76.485 64.755 77.825 ;
        RECT 64.965 76.485 65.195 77.825 ;
        RECT 65.375 77.325 65.715 78.005 ;
        RECT 65.895 77.505 66.225 78.615 ;
        RECT 66.395 78.145 66.575 78.615 ;
        RECT 66.745 78.315 67.075 78.795 ;
        RECT 67.250 78.145 67.420 78.615 ;
        RECT 66.395 77.945 67.420 78.145 ;
        RECT 65.375 76.425 65.605 77.325 ;
        RECT 65.895 77.205 66.440 77.505 ;
        RECT 65.805 76.245 66.050 77.025 ;
        RECT 66.220 76.975 66.440 77.205 ;
        RECT 66.610 77.155 67.035 77.775 ;
        RECT 67.230 77.155 67.490 77.775 ;
        RECT 67.685 77.655 67.970 78.795 ;
        RECT 67.700 76.975 67.960 77.485 ;
        RECT 66.220 76.785 67.960 76.975 ;
        RECT 66.220 76.425 66.650 76.785 ;
        RECT 67.230 76.245 67.960 76.615 ;
        RECT 68.160 76.425 68.440 78.615 ;
        RECT 68.715 77.865 68.885 78.625 ;
        RECT 69.065 78.035 69.395 78.795 ;
        RECT 68.715 77.695 69.380 77.865 ;
        RECT 69.565 77.720 69.835 78.625 ;
        RECT 69.210 77.550 69.380 77.695 ;
        RECT 68.645 77.145 68.975 77.515 ;
        RECT 69.210 77.220 69.495 77.550 ;
        RECT 69.210 76.965 69.380 77.220 ;
        RECT 68.715 76.795 69.380 76.965 ;
        RECT 69.665 76.920 69.835 77.720 ;
        RECT 70.005 77.630 70.295 78.795 ;
        RECT 70.485 78.205 70.725 78.595 ;
        RECT 70.895 78.385 71.245 78.795 ;
        RECT 70.485 78.005 71.235 78.205 ;
        RECT 68.715 76.415 68.885 76.795 ;
        RECT 69.065 76.245 69.395 76.625 ;
        RECT 69.575 76.415 69.835 76.920 ;
        RECT 70.005 76.245 70.295 76.970 ;
        RECT 70.485 76.485 70.715 77.825 ;
        RECT 70.895 77.325 71.235 78.005 ;
        RECT 71.415 77.505 71.745 78.615 ;
        RECT 71.915 78.145 72.095 78.615 ;
        RECT 72.265 78.315 72.595 78.795 ;
        RECT 72.770 78.145 72.940 78.615 ;
        RECT 71.915 77.945 72.940 78.145 ;
        RECT 70.895 76.425 71.125 77.325 ;
        RECT 71.415 77.205 71.960 77.505 ;
        RECT 71.325 76.245 71.570 77.025 ;
        RECT 71.740 76.975 71.960 77.205 ;
        RECT 72.130 77.155 72.555 77.775 ;
        RECT 72.750 77.155 73.010 77.775 ;
        RECT 73.205 77.655 73.490 78.795 ;
        RECT 73.220 76.975 73.480 77.485 ;
        RECT 71.740 76.785 73.480 76.975 ;
        RECT 71.740 76.425 72.170 76.785 ;
        RECT 72.750 76.245 73.480 76.615 ;
        RECT 73.680 76.425 73.960 78.615 ;
        RECT 74.145 77.720 74.415 78.625 ;
        RECT 74.585 78.035 74.915 78.795 ;
        RECT 75.095 77.865 75.275 78.625 ;
        RECT 74.145 76.920 74.325 77.720 ;
        RECT 74.600 77.695 75.275 77.865 ;
        RECT 75.525 77.705 76.735 78.795 ;
        RECT 74.600 77.550 74.770 77.695 ;
        RECT 74.495 77.220 74.770 77.550 ;
        RECT 74.600 76.965 74.770 77.220 ;
        RECT 74.995 77.145 75.335 77.515 ;
        RECT 75.525 77.165 76.045 77.705 ;
        RECT 76.215 76.995 76.735 77.535 ;
        RECT 74.145 76.415 74.405 76.920 ;
        RECT 74.600 76.795 75.265 76.965 ;
        RECT 74.585 76.245 74.915 76.625 ;
        RECT 75.095 76.415 75.265 76.795 ;
        RECT 75.525 76.245 76.735 76.995 ;
        RECT 5.520 76.075 76.820 76.245 ;
        RECT 5.605 75.325 6.815 76.075 ;
        RECT 5.605 74.785 6.125 75.325 ;
        RECT 7.375 75.275 7.705 76.075 ;
        RECT 7.875 75.425 8.045 75.905 ;
        RECT 8.215 75.595 8.545 76.075 ;
        RECT 8.715 75.425 8.885 75.905 ;
        RECT 9.055 75.595 9.385 76.075 ;
        RECT 9.555 75.425 9.725 75.905 ;
        RECT 9.895 75.595 10.225 76.075 ;
        RECT 10.395 75.425 10.565 75.905 ;
        RECT 10.735 75.595 11.065 76.075 ;
        RECT 11.235 75.425 11.405 75.900 ;
        RECT 11.575 75.595 11.905 76.075 ;
        RECT 12.075 75.425 12.245 75.905 ;
        RECT 7.875 75.255 10.565 75.425 ;
        RECT 10.825 75.255 12.245 75.425 ;
        RECT 13.425 75.415 13.700 76.075 ;
        RECT 13.870 75.445 14.120 75.905 ;
        RECT 14.295 75.580 14.625 76.075 ;
        RECT 6.295 74.615 6.815 75.155 ;
        RECT 7.875 74.715 8.130 75.255 ;
        RECT 10.825 75.085 11.000 75.255 ;
        RECT 13.870 75.235 14.040 75.445 ;
        RECT 14.805 75.410 15.035 75.855 ;
        RECT 8.375 74.915 11.000 75.085 ;
        RECT 10.825 74.715 11.000 74.915 ;
        RECT 11.180 74.885 12.280 75.085 ;
        RECT 13.425 74.715 14.040 75.235 ;
        RECT 14.210 74.735 14.440 75.165 ;
        RECT 14.625 74.915 15.035 75.410 ;
        RECT 15.205 75.590 15.995 75.855 ;
        RECT 15.205 74.735 15.460 75.590 ;
        RECT 16.190 75.445 16.525 75.905 ;
        RECT 16.695 75.615 16.865 76.075 ;
        RECT 17.035 75.445 17.365 75.905 ;
        RECT 17.535 75.615 17.705 76.075 ;
        RECT 17.875 75.695 19.885 75.905 ;
        RECT 17.875 75.445 18.125 75.695 ;
        RECT 15.630 74.915 16.015 75.395 ;
        RECT 16.190 75.255 18.125 75.445 ;
        RECT 18.295 75.355 19.465 75.525 ;
        RECT 18.295 75.085 18.545 75.355 ;
        RECT 19.635 75.275 19.885 75.695 ;
        RECT 16.210 74.835 17.830 75.085 ;
        RECT 5.605 73.525 6.815 74.615 ;
        RECT 7.375 73.525 7.705 74.675 ;
        RECT 7.875 74.545 10.565 74.715 ;
        RECT 10.825 74.545 12.325 74.715 ;
        RECT 7.875 73.695 8.045 74.545 ;
        RECT 8.215 73.525 8.545 74.325 ;
        RECT 8.715 73.695 8.885 74.545 ;
        RECT 9.055 73.525 9.385 74.325 ;
        RECT 9.555 73.695 9.725 74.545 ;
        RECT 9.895 73.525 10.225 74.325 ;
        RECT 10.395 73.695 10.565 74.545 ;
        RECT 10.815 73.525 10.985 74.325 ;
        RECT 11.155 73.695 11.485 74.545 ;
        RECT 11.655 73.525 11.825 74.325 ;
        RECT 11.995 73.695 12.325 74.545 ;
        RECT 13.425 73.525 13.685 74.535 ;
        RECT 13.855 74.365 14.025 74.715 ;
        RECT 14.210 74.565 16.000 74.735 ;
        RECT 18.010 74.665 18.545 75.085 ;
        RECT 18.715 74.835 20.155 75.085 ;
        RECT 13.855 73.695 14.130 74.365 ;
        RECT 14.330 73.525 14.545 74.370 ;
        RECT 14.770 74.270 15.020 74.565 ;
        RECT 15.245 74.205 15.575 74.395 ;
        RECT 14.730 73.695 15.205 74.035 ;
        RECT 15.385 74.030 15.575 74.205 ;
        RECT 15.745 74.200 16.000 74.565 ;
        RECT 15.385 73.525 16.015 74.030 ;
        RECT 16.190 73.525 16.445 74.665 ;
        RECT 16.615 74.495 19.465 74.665 ;
        RECT 16.615 73.695 16.945 74.495 ;
        RECT 17.115 73.525 17.285 74.325 ;
        RECT 17.455 73.695 17.785 74.495 ;
        RECT 17.955 73.525 18.125 74.325 ;
        RECT 18.295 73.695 18.625 74.495 ;
        RECT 18.795 73.525 18.965 74.325 ;
        RECT 19.135 73.695 19.465 74.495 ;
        RECT 19.635 73.525 19.885 74.325 ;
        RECT 20.325 73.695 21.075 75.905 ;
        RECT 21.335 75.525 21.505 75.905 ;
        RECT 21.685 75.695 22.015 76.075 ;
        RECT 21.335 75.355 22.000 75.525 ;
        RECT 22.195 75.400 22.455 75.905 ;
        RECT 21.265 74.805 21.605 75.175 ;
        RECT 21.830 75.100 22.000 75.355 ;
        RECT 21.830 74.770 22.105 75.100 ;
        RECT 21.830 74.625 22.000 74.770 ;
        RECT 21.325 74.455 22.000 74.625 ;
        RECT 22.275 74.600 22.455 75.400 ;
        RECT 22.645 75.265 22.885 76.075 ;
        RECT 23.055 75.265 23.385 75.905 ;
        RECT 23.555 75.265 23.825 76.075 ;
        RECT 24.005 75.355 24.345 75.865 ;
        RECT 22.625 74.835 22.975 75.085 ;
        RECT 23.145 74.665 23.315 75.265 ;
        RECT 23.485 74.835 23.835 75.085 ;
        RECT 21.325 73.695 21.505 74.455 ;
        RECT 21.685 73.525 22.015 74.285 ;
        RECT 22.185 73.695 22.455 74.600 ;
        RECT 22.635 74.495 23.315 74.665 ;
        RECT 22.635 73.710 22.965 74.495 ;
        RECT 23.495 73.525 23.825 74.665 ;
        RECT 24.005 73.955 24.265 75.355 ;
        RECT 24.515 75.275 24.785 76.075 ;
        RECT 24.440 74.835 24.770 75.085 ;
        RECT 24.965 74.835 25.245 75.805 ;
        RECT 25.425 74.835 25.725 75.805 ;
        RECT 25.905 74.835 26.255 75.800 ;
        RECT 26.475 75.575 26.970 75.905 ;
        RECT 24.455 74.665 24.770 74.835 ;
        RECT 26.475 74.665 26.645 75.575 ;
        RECT 27.310 75.525 27.640 75.905 ;
        RECT 27.810 75.695 28.995 75.865 ;
        RECT 29.255 75.605 29.425 76.075 ;
        RECT 24.455 74.495 26.645 74.665 ;
        RECT 24.005 73.695 24.345 73.955 ;
        RECT 24.515 73.525 24.845 74.325 ;
        RECT 25.310 73.695 25.560 74.495 ;
        RECT 25.745 73.525 26.075 74.245 ;
        RECT 26.295 73.695 26.545 74.495 ;
        RECT 26.815 74.085 27.055 75.395 ;
        RECT 27.310 75.355 27.855 75.525 ;
        RECT 27.225 74.835 27.485 75.185 ;
        RECT 27.685 74.715 27.855 75.355 ;
        RECT 28.225 75.425 28.610 75.515 ;
        RECT 29.595 75.425 29.925 75.890 ;
        RECT 28.225 75.255 29.925 75.425 ;
        RECT 30.095 75.255 30.265 76.075 ;
        RECT 30.435 75.425 30.765 75.895 ;
        RECT 30.935 75.595 31.105 76.075 ;
        RECT 30.435 75.255 31.195 75.425 ;
        RECT 31.365 75.350 31.655 76.075 ;
        RECT 28.025 74.885 28.370 75.085 ;
        RECT 28.540 74.885 28.930 75.085 ;
        RECT 27.685 74.665 28.470 74.715 ;
        RECT 27.390 74.490 28.470 74.665 ;
        RECT 26.715 73.525 27.050 73.905 ;
        RECT 27.390 73.695 27.720 74.490 ;
        RECT 27.890 73.525 28.130 74.310 ;
        RECT 28.300 74.285 28.470 74.490 ;
        RECT 28.640 74.455 28.930 74.885 ;
        RECT 29.120 74.875 29.605 75.085 ;
        RECT 29.775 74.875 30.215 75.085 ;
        RECT 30.385 74.875 30.715 75.085 ;
        RECT 29.120 74.455 29.425 74.875 ;
        RECT 30.385 74.705 30.555 74.875 ;
        RECT 29.595 74.535 30.555 74.705 ;
        RECT 29.595 74.285 29.765 74.535 ;
        RECT 28.300 74.115 29.765 74.285 ;
        RECT 28.690 73.695 29.445 74.115 ;
        RECT 29.935 73.525 30.265 74.365 ;
        RECT 30.885 74.285 31.195 75.255 ;
        RECT 30.435 74.115 31.195 74.285 ;
        RECT 30.435 73.695 30.685 74.115 ;
        RECT 30.855 73.525 31.195 73.945 ;
        RECT 31.365 73.525 31.655 74.690 ;
        RECT 31.825 73.695 32.575 75.905 ;
        RECT 32.745 75.565 33.050 76.075 ;
        RECT 32.745 74.835 33.060 75.395 ;
        RECT 33.230 75.085 33.480 75.895 ;
        RECT 33.650 75.550 33.910 76.075 ;
        RECT 34.090 75.085 34.340 75.895 ;
        RECT 34.510 75.515 34.770 76.075 ;
        RECT 34.940 75.425 35.200 75.880 ;
        RECT 35.370 75.595 35.630 76.075 ;
        RECT 35.800 75.425 36.060 75.880 ;
        RECT 36.230 75.595 36.490 76.075 ;
        RECT 36.660 75.425 36.920 75.880 ;
        RECT 37.090 75.595 37.335 76.075 ;
        RECT 37.505 75.425 37.780 75.880 ;
        RECT 37.950 75.595 38.195 76.075 ;
        RECT 38.365 75.425 38.625 75.880 ;
        RECT 38.805 75.595 39.055 76.075 ;
        RECT 39.225 75.425 39.485 75.880 ;
        RECT 39.665 75.595 39.915 76.075 ;
        RECT 40.085 75.425 40.345 75.880 ;
        RECT 40.525 75.595 40.785 76.075 ;
        RECT 40.955 75.425 41.215 75.880 ;
        RECT 41.385 75.595 41.685 76.075 ;
        RECT 42.035 75.595 42.335 76.075 ;
        RECT 42.505 75.425 42.765 75.880 ;
        RECT 42.935 75.595 43.195 76.075 ;
        RECT 43.375 75.425 43.635 75.880 ;
        RECT 43.805 75.595 44.055 76.075 ;
        RECT 44.235 75.425 44.495 75.880 ;
        RECT 44.665 75.595 44.915 76.075 ;
        RECT 45.095 75.425 45.355 75.880 ;
        RECT 45.525 75.595 45.770 76.075 ;
        RECT 45.940 75.425 46.215 75.880 ;
        RECT 46.385 75.595 46.630 76.075 ;
        RECT 46.800 75.425 47.060 75.880 ;
        RECT 47.230 75.595 47.490 76.075 ;
        RECT 47.660 75.425 47.920 75.880 ;
        RECT 48.090 75.595 48.350 76.075 ;
        RECT 48.520 75.425 48.780 75.880 ;
        RECT 48.950 75.515 49.210 76.075 ;
        RECT 34.940 75.255 41.685 75.425 ;
        RECT 33.230 74.835 40.350 75.085 ;
        RECT 32.755 73.525 33.050 74.335 ;
        RECT 33.230 73.695 33.475 74.835 ;
        RECT 33.650 73.525 33.910 74.335 ;
        RECT 34.090 73.700 34.340 74.835 ;
        RECT 40.520 74.665 41.685 75.255 ;
        RECT 34.940 74.440 41.685 74.665 ;
        RECT 42.035 75.255 48.780 75.425 ;
        RECT 42.035 74.665 43.200 75.255 ;
        RECT 49.380 75.085 49.630 75.895 ;
        RECT 49.810 75.550 50.070 76.075 ;
        RECT 50.240 75.085 50.490 75.895 ;
        RECT 50.670 75.565 50.975 76.075 ;
        RECT 51.235 75.525 51.405 75.905 ;
        RECT 51.620 75.695 51.950 76.075 ;
        RECT 43.370 74.835 50.490 75.085 ;
        RECT 50.660 74.835 50.975 75.395 ;
        RECT 51.235 75.355 51.950 75.525 ;
        RECT 42.035 74.440 48.780 74.665 ;
        RECT 34.940 74.425 40.345 74.440 ;
        RECT 34.510 73.530 34.770 74.325 ;
        RECT 34.940 73.700 35.200 74.425 ;
        RECT 35.370 73.530 35.630 74.255 ;
        RECT 35.800 73.700 36.060 74.425 ;
        RECT 36.230 73.530 36.490 74.255 ;
        RECT 36.660 73.700 36.920 74.425 ;
        RECT 37.090 73.530 37.350 74.255 ;
        RECT 37.520 73.700 37.780 74.425 ;
        RECT 37.950 73.530 38.195 74.255 ;
        RECT 38.365 73.700 38.625 74.425 ;
        RECT 38.810 73.530 39.055 74.255 ;
        RECT 39.225 73.700 39.485 74.425 ;
        RECT 39.670 73.530 39.915 74.255 ;
        RECT 40.085 73.700 40.345 74.425 ;
        RECT 40.530 73.530 40.785 74.255 ;
        RECT 40.955 73.700 41.245 74.440 ;
        RECT 34.510 73.525 40.785 73.530 ;
        RECT 41.415 73.525 41.685 74.270 ;
        RECT 42.035 73.525 42.305 74.270 ;
        RECT 42.475 73.700 42.765 74.440 ;
        RECT 43.375 74.425 48.780 74.440 ;
        RECT 42.935 73.530 43.190 74.255 ;
        RECT 43.375 73.700 43.635 74.425 ;
        RECT 43.805 73.530 44.050 74.255 ;
        RECT 44.235 73.700 44.495 74.425 ;
        RECT 44.665 73.530 44.910 74.255 ;
        RECT 45.095 73.700 45.355 74.425 ;
        RECT 45.525 73.530 45.770 74.255 ;
        RECT 45.940 73.700 46.200 74.425 ;
        RECT 46.370 73.530 46.630 74.255 ;
        RECT 46.800 73.700 47.060 74.425 ;
        RECT 47.230 73.530 47.490 74.255 ;
        RECT 47.660 73.700 47.920 74.425 ;
        RECT 48.090 73.530 48.350 74.255 ;
        RECT 48.520 73.700 48.780 74.425 ;
        RECT 48.950 73.530 49.210 74.325 ;
        RECT 49.380 73.700 49.630 74.835 ;
        RECT 42.935 73.525 49.210 73.530 ;
        RECT 49.810 73.525 50.070 74.335 ;
        RECT 50.245 73.695 50.490 74.835 ;
        RECT 51.145 74.805 51.500 75.175 ;
        RECT 51.780 75.165 51.950 75.355 ;
        RECT 52.120 75.330 52.375 75.905 ;
        RECT 51.780 74.835 52.035 75.165 ;
        RECT 51.780 74.625 51.950 74.835 ;
        RECT 51.235 74.455 51.950 74.625 ;
        RECT 52.205 74.600 52.375 75.330 ;
        RECT 52.550 75.235 52.810 76.075 ;
        RECT 52.990 75.695 55.005 75.865 ;
        RECT 55.195 75.695 55.525 76.075 ;
        RECT 52.990 75.375 53.245 75.695 ;
        RECT 52.990 74.835 53.230 75.165 ;
        RECT 53.415 74.715 53.745 75.525 ;
        RECT 54.255 75.255 55.945 75.525 ;
        RECT 56.115 75.275 56.495 76.075 ;
        RECT 57.125 75.350 57.415 76.075 ;
        RECT 57.585 75.565 57.890 76.075 ;
        RECT 53.970 74.885 55.060 75.085 ;
        RECT 55.370 74.885 56.495 75.085 ;
        RECT 57.585 74.835 57.900 75.395 ;
        RECT 58.070 75.085 58.320 75.895 ;
        RECT 58.490 75.550 58.750 76.075 ;
        RECT 58.930 75.085 59.180 75.895 ;
        RECT 59.350 75.515 59.610 76.075 ;
        RECT 59.780 75.425 60.040 75.880 ;
        RECT 60.210 75.595 60.470 76.075 ;
        RECT 60.640 75.425 60.900 75.880 ;
        RECT 61.070 75.595 61.330 76.075 ;
        RECT 61.500 75.425 61.760 75.880 ;
        RECT 61.930 75.595 62.175 76.075 ;
        RECT 62.345 75.425 62.620 75.880 ;
        RECT 62.790 75.595 63.035 76.075 ;
        RECT 63.205 75.425 63.465 75.880 ;
        RECT 63.645 75.595 63.895 76.075 ;
        RECT 64.065 75.425 64.325 75.880 ;
        RECT 64.505 75.595 64.755 76.075 ;
        RECT 64.925 75.425 65.185 75.880 ;
        RECT 65.365 75.595 65.625 76.075 ;
        RECT 65.795 75.425 66.055 75.880 ;
        RECT 66.225 75.595 66.525 76.075 ;
        RECT 59.780 75.255 66.525 75.425 ;
        RECT 58.070 74.835 65.190 75.085 ;
        RECT 50.670 73.525 50.965 74.335 ;
        RECT 51.235 73.695 51.405 74.455 ;
        RECT 51.620 73.525 51.950 74.285 ;
        RECT 52.120 73.695 52.375 74.600 ;
        RECT 52.550 73.525 52.810 74.675 ;
        RECT 52.990 73.525 53.245 74.665 ;
        RECT 53.415 74.495 55.945 74.715 ;
        RECT 53.415 73.695 53.745 74.495 ;
        RECT 53.915 73.525 54.085 74.325 ;
        RECT 54.255 73.695 54.585 74.495 ;
        RECT 54.755 73.525 55.445 74.325 ;
        RECT 55.615 73.695 55.945 74.495 ;
        RECT 56.115 73.525 56.495 74.715 ;
        RECT 57.125 73.525 57.415 74.690 ;
        RECT 57.595 73.525 57.890 74.335 ;
        RECT 58.070 73.695 58.315 74.835 ;
        RECT 58.490 73.525 58.750 74.335 ;
        RECT 58.930 73.700 59.180 74.835 ;
        RECT 65.360 74.665 66.525 75.255 ;
        RECT 59.780 74.440 66.525 74.665 ;
        RECT 66.805 74.495 67.035 75.835 ;
        RECT 67.215 74.995 67.445 75.895 ;
        RECT 67.645 75.295 67.890 76.075 ;
        RECT 68.060 75.535 68.490 75.895 ;
        RECT 69.070 75.705 69.800 76.075 ;
        RECT 68.060 75.345 69.800 75.535 ;
        RECT 68.060 75.115 68.280 75.345 ;
        RECT 59.780 74.425 65.185 74.440 ;
        RECT 59.350 73.530 59.610 74.325 ;
        RECT 59.780 73.700 60.040 74.425 ;
        RECT 60.210 73.530 60.470 74.255 ;
        RECT 60.640 73.700 60.900 74.425 ;
        RECT 61.070 73.530 61.330 74.255 ;
        RECT 61.500 73.700 61.760 74.425 ;
        RECT 61.930 73.530 62.190 74.255 ;
        RECT 62.360 73.700 62.620 74.425 ;
        RECT 62.790 73.530 63.035 74.255 ;
        RECT 63.205 73.700 63.465 74.425 ;
        RECT 63.650 73.530 63.895 74.255 ;
        RECT 64.065 73.700 64.325 74.425 ;
        RECT 64.510 73.530 64.755 74.255 ;
        RECT 64.925 73.700 65.185 74.425 ;
        RECT 65.370 73.530 65.625 74.255 ;
        RECT 65.795 73.700 66.085 74.440 ;
        RECT 67.215 74.315 67.555 74.995 ;
        RECT 59.350 73.525 65.625 73.530 ;
        RECT 66.255 73.525 66.525 74.270 ;
        RECT 66.805 74.115 67.555 74.315 ;
        RECT 67.735 74.815 68.280 75.115 ;
        RECT 66.805 73.725 67.045 74.115 ;
        RECT 67.215 73.525 67.565 73.935 ;
        RECT 67.735 73.705 68.065 74.815 ;
        RECT 68.450 74.545 68.875 75.165 ;
        RECT 69.070 74.545 69.330 75.165 ;
        RECT 69.540 74.835 69.800 75.345 ;
        RECT 68.235 74.175 69.260 74.375 ;
        RECT 68.235 73.705 68.415 74.175 ;
        RECT 68.585 73.525 68.915 74.005 ;
        RECT 69.090 73.705 69.260 74.175 ;
        RECT 69.525 73.525 69.810 74.665 ;
        RECT 70.000 73.705 70.280 75.895 ;
        RECT 70.485 74.495 70.715 75.835 ;
        RECT 70.895 74.995 71.125 75.895 ;
        RECT 71.325 75.295 71.570 76.075 ;
        RECT 71.740 75.535 72.170 75.895 ;
        RECT 72.750 75.705 73.480 76.075 ;
        RECT 71.740 75.345 73.480 75.535 ;
        RECT 71.740 75.115 71.960 75.345 ;
        RECT 70.895 74.315 71.235 74.995 ;
        RECT 70.485 74.115 71.235 74.315 ;
        RECT 71.415 74.815 71.960 75.115 ;
        RECT 70.485 73.725 70.725 74.115 ;
        RECT 70.895 73.525 71.245 73.935 ;
        RECT 71.415 73.705 71.745 74.815 ;
        RECT 72.130 74.545 72.555 75.165 ;
        RECT 72.750 74.545 73.010 75.165 ;
        RECT 73.220 74.835 73.480 75.345 ;
        RECT 71.915 74.175 72.940 74.375 ;
        RECT 71.915 73.705 72.095 74.175 ;
        RECT 72.265 73.525 72.595 74.005 ;
        RECT 72.770 73.705 72.940 74.175 ;
        RECT 73.205 73.525 73.490 74.665 ;
        RECT 73.680 73.705 73.960 75.895 ;
        RECT 74.185 75.255 74.415 76.075 ;
        RECT 74.585 75.275 74.915 75.905 ;
        RECT 74.165 74.835 74.495 75.085 ;
        RECT 74.665 74.675 74.915 75.275 ;
        RECT 75.085 75.255 75.295 76.075 ;
        RECT 75.525 75.325 76.735 76.075 ;
        RECT 74.185 73.525 74.415 74.665 ;
        RECT 74.585 73.695 74.915 74.675 ;
        RECT 75.085 73.525 75.295 74.665 ;
        RECT 75.525 74.615 76.045 75.155 ;
        RECT 76.215 74.785 76.735 75.325 ;
        RECT 75.525 73.525 76.735 74.615 ;
        RECT 5.520 73.355 76.820 73.525 ;
        RECT 5.605 72.265 6.815 73.355 ;
        RECT 5.605 71.555 6.125 72.095 ;
        RECT 6.295 71.725 6.815 72.265 ;
        RECT 7.450 72.205 7.710 73.355 ;
        RECT 7.885 72.280 8.140 73.185 ;
        RECT 8.310 72.595 8.640 73.355 ;
        RECT 8.855 72.425 9.025 73.185 ;
        RECT 9.485 72.685 9.765 73.355 ;
        RECT 5.605 70.805 6.815 71.555 ;
        RECT 7.450 70.805 7.710 71.645 ;
        RECT 7.885 71.550 8.055 72.280 ;
        RECT 8.310 72.255 9.025 72.425 ;
        RECT 9.935 72.465 10.235 73.015 ;
        RECT 10.435 72.635 10.765 73.355 ;
        RECT 10.955 72.635 11.415 73.185 ;
        RECT 12.085 72.895 12.300 73.355 ;
        RECT 12.470 72.725 12.800 73.185 ;
        RECT 8.310 72.045 8.480 72.255 ;
        RECT 8.225 71.715 8.480 72.045 ;
        RECT 7.885 70.975 8.140 71.550 ;
        RECT 8.310 71.525 8.480 71.715 ;
        RECT 8.760 71.705 9.115 72.075 ;
        RECT 9.300 72.045 9.565 72.405 ;
        RECT 9.935 72.295 10.875 72.465 ;
        RECT 10.705 72.045 10.875 72.295 ;
        RECT 9.300 71.795 9.975 72.045 ;
        RECT 10.195 71.795 10.535 72.045 ;
        RECT 10.705 71.715 10.995 72.045 ;
        RECT 10.705 71.625 10.875 71.715 ;
        RECT 8.310 71.355 9.025 71.525 ;
        RECT 8.310 70.805 8.640 71.185 ;
        RECT 8.855 70.975 9.025 71.355 ;
        RECT 9.485 71.435 10.875 71.625 ;
        RECT 9.485 71.075 9.815 71.435 ;
        RECT 11.165 71.265 11.415 72.635 ;
        RECT 10.435 70.805 10.685 71.265 ;
        RECT 10.855 70.975 11.415 71.265 ;
        RECT 11.630 72.555 12.800 72.725 ;
        RECT 12.970 72.555 13.220 73.355 ;
        RECT 13.920 72.565 14.455 73.185 ;
        RECT 11.630 71.265 12.000 72.555 ;
        RECT 13.430 72.385 13.710 72.545 ;
        RECT 12.375 72.215 13.710 72.385 ;
        RECT 12.375 72.045 12.545 72.215 ;
        RECT 12.170 71.795 12.545 72.045 ;
        RECT 12.715 71.795 13.190 72.035 ;
        RECT 13.360 71.795 13.710 72.035 ;
        RECT 12.375 71.625 12.545 71.795 ;
        RECT 12.375 71.455 13.710 71.625 ;
        RECT 11.630 70.975 12.380 71.265 ;
        RECT 12.890 70.805 13.220 71.265 ;
        RECT 13.440 71.245 13.710 71.455 ;
        RECT 13.920 71.545 14.235 72.565 ;
        RECT 14.625 72.555 14.955 73.355 ;
        RECT 15.440 72.385 15.830 72.560 ;
        RECT 16.205 72.555 16.485 73.355 ;
        RECT 16.685 72.385 17.015 73.185 ;
        RECT 17.215 72.555 17.385 73.355 ;
        RECT 17.555 72.385 17.885 73.185 ;
        RECT 14.405 72.215 15.830 72.385 ;
        RECT 14.405 71.715 14.575 72.215 ;
        RECT 13.920 70.975 14.535 71.545 ;
        RECT 14.825 71.485 15.090 72.045 ;
        RECT 15.260 71.315 15.430 72.215 ;
        RECT 15.600 71.485 15.955 72.045 ;
        RECT 16.185 71.715 16.425 72.385 ;
        RECT 16.605 72.215 17.885 72.385 ;
        RECT 18.055 72.215 18.315 73.355 ;
        RECT 16.605 71.545 16.775 72.215 ;
        RECT 18.485 72.190 18.775 73.355 ;
        RECT 19.460 72.485 19.745 73.355 ;
        RECT 19.915 72.725 20.175 73.185 ;
        RECT 20.350 72.895 20.605 73.355 ;
        RECT 20.775 72.725 21.035 73.185 ;
        RECT 19.915 72.555 21.035 72.725 ;
        RECT 21.205 72.555 21.515 73.355 ;
        RECT 19.915 72.305 20.175 72.555 ;
        RECT 21.685 72.385 21.995 73.185 ;
        RECT 22.365 72.685 22.645 73.355 ;
        RECT 19.420 72.135 20.175 72.305 ;
        RECT 20.965 72.215 21.995 72.385 ;
        RECT 16.945 71.715 17.255 72.045 ;
        RECT 17.425 71.715 17.805 72.045 ;
        RECT 18.005 71.715 18.290 72.045 ;
        RECT 17.050 71.545 17.255 71.715 ;
        RECT 14.705 70.805 14.920 71.315 ;
        RECT 15.150 70.985 15.430 71.315 ;
        RECT 15.610 70.805 15.850 71.315 ;
        RECT 16.185 70.975 16.880 71.545 ;
        RECT 17.050 71.020 17.400 71.545 ;
        RECT 17.590 71.020 17.805 71.715 ;
        RECT 19.420 71.625 19.825 72.135 ;
        RECT 20.965 71.965 21.135 72.215 ;
        RECT 19.995 71.795 21.135 71.965 ;
        RECT 17.975 70.805 18.310 71.545 ;
        RECT 18.485 70.805 18.775 71.530 ;
        RECT 19.420 71.455 21.070 71.625 ;
        RECT 21.305 71.475 21.655 72.045 ;
        RECT 19.465 70.805 19.745 71.285 ;
        RECT 19.915 71.065 20.175 71.455 ;
        RECT 20.350 70.805 20.605 71.285 ;
        RECT 20.775 71.065 21.070 71.455 ;
        RECT 21.825 71.305 21.995 72.215 ;
        RECT 22.165 72.045 22.480 72.485 ;
        RECT 22.815 72.465 23.115 73.015 ;
        RECT 23.325 72.635 23.655 73.355 ;
        RECT 23.845 72.635 24.295 73.185 ;
        RECT 22.815 72.295 23.755 72.465 ;
        RECT 23.585 72.045 23.755 72.295 ;
        RECT 22.165 71.795 22.855 72.045 ;
        RECT 23.085 71.795 23.415 72.045 ;
        RECT 23.585 71.715 23.875 72.045 ;
        RECT 23.585 71.625 23.755 71.715 ;
        RECT 21.250 70.805 21.525 71.285 ;
        RECT 21.695 70.975 21.995 71.305 ;
        RECT 22.365 71.435 23.755 71.625 ;
        RECT 22.365 71.075 22.695 71.435 ;
        RECT 24.045 71.265 24.295 72.635 ;
        RECT 24.465 72.215 24.755 73.355 ;
        RECT 24.935 72.545 25.230 73.355 ;
        RECT 25.410 72.045 25.655 73.185 ;
        RECT 25.830 72.545 26.090 73.355 ;
        RECT 26.690 73.350 32.965 73.355 ;
        RECT 26.270 72.045 26.520 73.180 ;
        RECT 26.690 72.555 26.950 73.350 ;
        RECT 27.120 72.455 27.380 73.180 ;
        RECT 27.550 72.625 27.810 73.350 ;
        RECT 27.980 72.455 28.240 73.180 ;
        RECT 28.410 72.625 28.670 73.350 ;
        RECT 28.840 72.455 29.100 73.180 ;
        RECT 29.270 72.625 29.530 73.350 ;
        RECT 29.700 72.455 29.960 73.180 ;
        RECT 30.130 72.625 30.375 73.350 ;
        RECT 30.545 72.455 30.805 73.180 ;
        RECT 30.990 72.625 31.235 73.350 ;
        RECT 31.405 72.455 31.665 73.180 ;
        RECT 31.850 72.625 32.095 73.350 ;
        RECT 32.265 72.455 32.525 73.180 ;
        RECT 32.710 72.625 32.965 73.350 ;
        RECT 27.120 72.440 32.525 72.455 ;
        RECT 33.135 72.440 33.425 73.180 ;
        RECT 33.595 72.610 33.865 73.355 ;
        RECT 27.120 72.215 33.865 72.440 ;
        RECT 34.165 72.215 34.395 73.355 ;
        RECT 23.325 70.805 23.575 71.265 ;
        RECT 23.745 70.975 24.295 71.265 ;
        RECT 24.465 70.805 24.755 71.605 ;
        RECT 24.925 71.485 25.240 72.045 ;
        RECT 25.410 71.795 32.530 72.045 ;
        RECT 24.925 70.805 25.230 71.315 ;
        RECT 25.410 70.985 25.660 71.795 ;
        RECT 25.830 70.805 26.090 71.330 ;
        RECT 26.270 70.985 26.520 71.795 ;
        RECT 32.700 71.655 33.865 72.215 ;
        RECT 34.565 72.205 34.895 73.185 ;
        RECT 35.065 72.215 35.275 73.355 ;
        RECT 35.505 72.215 35.765 73.355 ;
        RECT 35.935 72.205 36.265 73.185 ;
        RECT 36.435 72.215 36.715 73.355 ;
        RECT 36.885 72.280 37.155 73.185 ;
        RECT 37.325 72.595 37.655 73.355 ;
        RECT 37.835 72.425 38.005 73.185 ;
        RECT 34.145 71.795 34.475 72.045 ;
        RECT 32.700 71.625 33.895 71.655 ;
        RECT 27.120 71.485 33.895 71.625 ;
        RECT 27.120 71.455 33.865 71.485 ;
        RECT 26.690 70.805 26.950 71.365 ;
        RECT 27.120 71.000 27.380 71.455 ;
        RECT 27.550 70.805 27.810 71.285 ;
        RECT 27.980 71.000 28.240 71.455 ;
        RECT 28.410 70.805 28.670 71.285 ;
        RECT 28.840 71.000 29.100 71.455 ;
        RECT 29.270 70.805 29.515 71.285 ;
        RECT 29.685 71.000 29.960 71.455 ;
        RECT 30.130 70.805 30.375 71.285 ;
        RECT 30.545 71.000 30.805 71.455 ;
        RECT 30.985 70.805 31.235 71.285 ;
        RECT 31.405 71.000 31.665 71.455 ;
        RECT 31.845 70.805 32.095 71.285 ;
        RECT 32.265 71.000 32.525 71.455 ;
        RECT 32.705 70.805 32.965 71.285 ;
        RECT 33.135 71.000 33.395 71.455 ;
        RECT 33.565 70.805 33.865 71.285 ;
        RECT 34.165 70.805 34.395 71.625 ;
        RECT 34.645 71.605 34.895 72.205 ;
        RECT 35.525 71.795 35.860 72.045 ;
        RECT 34.565 70.975 34.895 71.605 ;
        RECT 35.065 70.805 35.275 71.625 ;
        RECT 36.030 71.605 36.200 72.205 ;
        RECT 36.370 71.775 36.705 72.045 ;
        RECT 35.505 70.975 36.200 71.605 ;
        RECT 36.405 70.805 36.715 71.605 ;
        RECT 36.885 71.480 37.055 72.280 ;
        RECT 37.340 72.255 38.005 72.425 ;
        RECT 38.265 72.280 38.535 73.185 ;
        RECT 38.705 72.595 39.035 73.355 ;
        RECT 39.215 72.425 39.395 73.185 ;
        RECT 37.340 72.110 37.510 72.255 ;
        RECT 37.225 71.780 37.510 72.110 ;
        RECT 37.340 71.525 37.510 71.780 ;
        RECT 37.745 71.705 38.075 72.075 ;
        RECT 36.885 70.975 37.145 71.480 ;
        RECT 37.340 71.355 38.005 71.525 ;
        RECT 37.325 70.805 37.655 71.185 ;
        RECT 37.835 70.975 38.005 71.355 ;
        RECT 38.265 71.480 38.445 72.280 ;
        RECT 38.720 72.255 39.395 72.425 ;
        RECT 39.645 72.280 39.915 73.185 ;
        RECT 40.085 72.595 40.415 73.355 ;
        RECT 40.595 72.425 40.775 73.185 ;
        RECT 38.720 72.110 38.890 72.255 ;
        RECT 38.615 71.780 38.890 72.110 ;
        RECT 38.720 71.525 38.890 71.780 ;
        RECT 39.115 71.705 39.455 72.075 ;
        RECT 38.265 70.975 38.525 71.480 ;
        RECT 38.720 71.355 39.385 71.525 ;
        RECT 38.705 70.805 39.035 71.185 ;
        RECT 39.215 70.975 39.385 71.355 ;
        RECT 39.645 71.480 39.825 72.280 ;
        RECT 40.100 72.255 40.775 72.425 ;
        RECT 41.025 72.265 43.615 73.355 ;
        RECT 40.100 72.110 40.270 72.255 ;
        RECT 39.995 71.780 40.270 72.110 ;
        RECT 40.100 71.525 40.270 71.780 ;
        RECT 40.495 71.705 40.835 72.075 ;
        RECT 41.025 71.575 42.235 72.095 ;
        RECT 42.405 71.745 43.615 72.265 ;
        RECT 44.245 72.190 44.535 73.355 ;
        RECT 44.705 72.385 44.995 73.185 ;
        RECT 45.165 72.555 45.400 73.355 ;
        RECT 45.585 73.015 47.120 73.185 ;
        RECT 45.585 72.385 45.915 73.015 ;
        RECT 44.705 72.215 45.915 72.385 ;
        RECT 44.705 71.715 44.950 72.045 ;
        RECT 39.645 70.975 39.905 71.480 ;
        RECT 40.100 71.355 40.765 71.525 ;
        RECT 40.085 70.805 40.415 71.185 ;
        RECT 40.595 70.975 40.765 71.355 ;
        RECT 41.025 70.805 43.615 71.575 ;
        RECT 45.120 71.545 45.290 72.215 ;
        RECT 46.085 72.045 46.320 72.790 ;
        RECT 45.460 71.715 45.860 72.045 ;
        RECT 46.030 71.715 46.320 72.045 ;
        RECT 46.510 72.045 46.780 72.790 ;
        RECT 46.950 72.385 47.120 73.015 ;
        RECT 47.290 72.555 47.685 73.355 ;
        RECT 46.950 72.215 47.685 72.385 ;
        RECT 46.510 71.715 46.840 72.045 ;
        RECT 47.010 71.715 47.345 72.045 ;
        RECT 47.515 71.715 47.685 72.215 ;
        RECT 47.855 72.035 48.210 73.185 ;
        RECT 48.380 72.205 48.675 73.355 ;
        RECT 48.855 72.215 49.185 73.355 ;
        RECT 49.715 72.385 50.045 73.170 ;
        RECT 50.235 72.545 50.530 73.355 ;
        RECT 49.365 72.215 50.045 72.385 ;
        RECT 47.855 71.775 48.675 72.035 ;
        RECT 48.845 71.795 49.195 72.045 ;
        RECT 47.855 71.715 48.210 71.775 ;
        RECT 44.245 70.805 44.535 71.530 ;
        RECT 44.705 70.975 45.290 71.545 ;
        RECT 45.540 71.375 46.925 71.545 ;
        RECT 45.540 71.030 45.870 71.375 ;
        RECT 46.085 70.805 46.460 71.205 ;
        RECT 46.640 71.030 46.925 71.375 ;
        RECT 47.095 70.805 47.765 71.545 ;
        RECT 47.935 70.975 48.210 71.715 ;
        RECT 49.365 71.615 49.535 72.215 ;
        RECT 50.710 72.045 50.955 73.185 ;
        RECT 51.130 72.545 51.390 73.355 ;
        RECT 51.990 73.350 58.265 73.355 ;
        RECT 51.570 72.045 51.820 73.180 ;
        RECT 51.990 72.555 52.250 73.350 ;
        RECT 52.420 72.455 52.680 73.180 ;
        RECT 52.850 72.625 53.110 73.350 ;
        RECT 53.280 72.455 53.540 73.180 ;
        RECT 53.710 72.625 53.970 73.350 ;
        RECT 54.140 72.455 54.400 73.180 ;
        RECT 54.570 72.625 54.830 73.350 ;
        RECT 55.000 72.455 55.260 73.180 ;
        RECT 55.430 72.625 55.675 73.350 ;
        RECT 55.845 72.455 56.105 73.180 ;
        RECT 56.290 72.625 56.535 73.350 ;
        RECT 56.705 72.455 56.965 73.180 ;
        RECT 57.150 72.625 57.395 73.350 ;
        RECT 57.565 72.455 57.825 73.180 ;
        RECT 58.010 72.625 58.265 73.350 ;
        RECT 52.420 72.440 57.825 72.455 ;
        RECT 58.435 72.440 58.725 73.180 ;
        RECT 58.895 72.610 59.165 73.355 ;
        RECT 59.435 72.545 59.730 73.355 ;
        RECT 52.420 72.215 59.165 72.440 ;
        RECT 49.705 71.795 50.055 72.045 ;
        RECT 48.380 70.805 48.675 71.605 ;
        RECT 48.855 70.805 49.125 71.615 ;
        RECT 49.295 70.975 49.625 71.615 ;
        RECT 49.795 70.805 50.035 71.615 ;
        RECT 50.225 71.485 50.540 72.045 ;
        RECT 50.710 71.795 57.830 72.045 ;
        RECT 50.225 70.805 50.530 71.315 ;
        RECT 50.710 70.985 50.960 71.795 ;
        RECT 51.130 70.805 51.390 71.330 ;
        RECT 51.570 70.985 51.820 71.795 ;
        RECT 58.000 71.625 59.165 72.215 ;
        RECT 59.910 72.045 60.155 73.185 ;
        RECT 60.330 72.545 60.590 73.355 ;
        RECT 61.190 73.350 67.465 73.355 ;
        RECT 60.770 72.045 61.020 73.180 ;
        RECT 61.190 72.555 61.450 73.350 ;
        RECT 61.620 72.455 61.880 73.180 ;
        RECT 62.050 72.625 62.310 73.350 ;
        RECT 62.480 72.455 62.740 73.180 ;
        RECT 62.910 72.625 63.170 73.350 ;
        RECT 63.340 72.455 63.600 73.180 ;
        RECT 63.770 72.625 64.030 73.350 ;
        RECT 64.200 72.455 64.460 73.180 ;
        RECT 64.630 72.625 64.875 73.350 ;
        RECT 65.045 72.455 65.305 73.180 ;
        RECT 65.490 72.625 65.735 73.350 ;
        RECT 65.905 72.455 66.165 73.180 ;
        RECT 66.350 72.625 66.595 73.350 ;
        RECT 66.765 72.455 67.025 73.180 ;
        RECT 67.210 72.625 67.465 73.350 ;
        RECT 61.620 72.440 67.025 72.455 ;
        RECT 67.635 72.440 67.925 73.180 ;
        RECT 68.095 72.610 68.365 73.355 ;
        RECT 61.620 72.215 68.365 72.440 ;
        RECT 68.665 72.215 68.895 73.355 ;
        RECT 52.420 71.455 59.165 71.625 ;
        RECT 59.425 71.485 59.740 72.045 ;
        RECT 59.910 71.795 67.030 72.045 ;
        RECT 51.990 70.805 52.250 71.365 ;
        RECT 52.420 71.000 52.680 71.455 ;
        RECT 52.850 70.805 53.110 71.285 ;
        RECT 53.280 71.000 53.540 71.455 ;
        RECT 53.710 70.805 53.970 71.285 ;
        RECT 54.140 71.000 54.400 71.455 ;
        RECT 54.570 70.805 54.815 71.285 ;
        RECT 54.985 71.000 55.260 71.455 ;
        RECT 55.430 70.805 55.675 71.285 ;
        RECT 55.845 71.000 56.105 71.455 ;
        RECT 56.285 70.805 56.535 71.285 ;
        RECT 56.705 71.000 56.965 71.455 ;
        RECT 57.145 70.805 57.395 71.285 ;
        RECT 57.565 71.000 57.825 71.455 ;
        RECT 58.005 70.805 58.265 71.285 ;
        RECT 58.435 71.000 58.695 71.455 ;
        RECT 58.865 70.805 59.165 71.285 ;
        RECT 59.425 70.805 59.730 71.315 ;
        RECT 59.910 70.985 60.160 71.795 ;
        RECT 60.330 70.805 60.590 71.330 ;
        RECT 60.770 70.985 61.020 71.795 ;
        RECT 67.200 71.625 68.365 72.215 ;
        RECT 69.065 72.205 69.395 73.185 ;
        RECT 69.565 72.215 69.775 73.355 ;
        RECT 68.645 71.795 68.975 72.045 ;
        RECT 61.620 71.455 68.365 71.625 ;
        RECT 61.190 70.805 61.450 71.365 ;
        RECT 61.620 71.000 61.880 71.455 ;
        RECT 62.050 70.805 62.310 71.285 ;
        RECT 62.480 71.000 62.740 71.455 ;
        RECT 62.910 70.805 63.170 71.285 ;
        RECT 63.340 71.000 63.600 71.455 ;
        RECT 63.770 70.805 64.015 71.285 ;
        RECT 64.185 71.000 64.460 71.455 ;
        RECT 64.630 70.805 64.875 71.285 ;
        RECT 65.045 71.000 65.305 71.455 ;
        RECT 65.485 70.805 65.735 71.285 ;
        RECT 65.905 71.000 66.165 71.455 ;
        RECT 66.345 70.805 66.595 71.285 ;
        RECT 66.765 71.000 67.025 71.455 ;
        RECT 67.205 70.805 67.465 71.285 ;
        RECT 67.635 71.000 67.895 71.455 ;
        RECT 68.065 70.805 68.365 71.285 ;
        RECT 68.665 70.805 68.895 71.625 ;
        RECT 69.145 71.605 69.395 72.205 ;
        RECT 70.005 72.190 70.295 73.355 ;
        RECT 70.485 72.765 70.725 73.155 ;
        RECT 70.895 72.945 71.245 73.355 ;
        RECT 70.485 72.565 71.235 72.765 ;
        RECT 69.065 70.975 69.395 71.605 ;
        RECT 69.565 70.805 69.775 71.625 ;
        RECT 70.005 70.805 70.295 71.530 ;
        RECT 70.485 71.045 70.715 72.385 ;
        RECT 70.895 71.885 71.235 72.565 ;
        RECT 71.415 72.065 71.745 73.175 ;
        RECT 71.915 72.705 72.095 73.175 ;
        RECT 72.265 72.875 72.595 73.355 ;
        RECT 72.770 72.705 72.940 73.175 ;
        RECT 71.915 72.505 72.940 72.705 ;
        RECT 70.895 70.985 71.125 71.885 ;
        RECT 71.415 71.765 71.960 72.065 ;
        RECT 71.325 70.805 71.570 71.585 ;
        RECT 71.740 71.535 71.960 71.765 ;
        RECT 72.130 71.715 72.555 72.335 ;
        RECT 72.750 71.715 73.010 72.335 ;
        RECT 73.205 72.215 73.490 73.355 ;
        RECT 73.220 71.535 73.480 72.045 ;
        RECT 71.740 71.345 73.480 71.535 ;
        RECT 71.740 70.985 72.170 71.345 ;
        RECT 72.750 70.805 73.480 71.175 ;
        RECT 73.680 70.985 73.960 73.175 ;
        RECT 74.145 70.975 74.895 73.185 ;
        RECT 75.525 72.265 76.735 73.355 ;
        RECT 75.525 71.725 76.045 72.265 ;
        RECT 76.215 71.555 76.735 72.095 ;
        RECT 75.525 70.805 76.735 71.555 ;
        RECT 5.520 70.635 76.820 70.805 ;
        RECT 5.605 69.885 6.815 70.635 ;
        RECT 5.605 69.345 6.125 69.885 ;
        RECT 7.445 69.835 7.735 70.635 ;
        RECT 7.905 70.175 8.455 70.465 ;
        RECT 8.625 70.175 8.875 70.635 ;
        RECT 6.295 69.175 6.815 69.715 ;
        RECT 5.605 68.085 6.815 69.175 ;
        RECT 7.445 68.085 7.735 69.225 ;
        RECT 7.905 68.805 8.155 70.175 ;
        RECT 9.505 70.005 9.835 70.365 ;
        RECT 10.370 70.125 10.610 70.635 ;
        RECT 10.790 70.125 11.070 70.455 ;
        RECT 11.300 70.125 11.515 70.635 ;
        RECT 8.445 69.815 9.835 70.005 ;
        RECT 8.445 69.725 8.615 69.815 ;
        RECT 8.325 69.395 8.615 69.725 ;
        RECT 8.785 69.395 9.115 69.645 ;
        RECT 9.345 69.395 10.035 69.645 ;
        RECT 10.265 69.395 10.620 69.955 ;
        RECT 8.445 69.145 8.615 69.395 ;
        RECT 8.445 68.975 9.385 69.145 ;
        RECT 7.905 68.255 8.355 68.805 ;
        RECT 8.545 68.085 8.875 68.805 ;
        RECT 9.085 68.425 9.385 68.975 ;
        RECT 9.720 68.955 10.035 69.395 ;
        RECT 10.790 69.225 10.960 70.125 ;
        RECT 11.130 69.395 11.395 69.955 ;
        RECT 11.685 69.895 12.300 70.465 ;
        RECT 12.515 69.915 12.845 70.635 ;
        RECT 13.390 70.235 15.005 70.405 ;
        RECT 15.175 70.235 15.505 70.635 ;
        RECT 14.835 70.065 15.005 70.235 ;
        RECT 15.675 70.160 16.010 70.420 ;
        RECT 11.645 69.225 11.815 69.725 ;
        RECT 10.390 69.055 11.815 69.225 ;
        RECT 10.390 68.880 10.780 69.055 ;
        RECT 9.555 68.085 9.835 68.755 ;
        RECT 11.265 68.085 11.595 68.885 ;
        RECT 11.985 68.875 12.300 69.895 ;
        RECT 12.570 69.395 12.920 69.725 ;
        RECT 13.230 69.395 13.650 70.060 ;
        RECT 13.820 69.395 14.110 70.055 ;
        RECT 14.300 69.615 14.570 70.055 ;
        RECT 14.835 69.895 15.395 70.065 ;
        RECT 15.225 69.725 15.395 69.895 ;
        RECT 14.780 69.615 15.030 69.725 ;
        RECT 14.300 69.445 14.575 69.615 ;
        RECT 14.780 69.445 15.035 69.615 ;
        RECT 14.300 69.395 14.570 69.445 ;
        RECT 14.780 69.395 15.030 69.445 ;
        RECT 15.225 69.395 15.530 69.725 ;
        RECT 12.570 69.275 12.775 69.395 ;
        RECT 12.565 69.105 12.775 69.275 ;
        RECT 15.225 69.225 15.395 69.395 ;
        RECT 13.025 69.055 15.395 69.225 ;
        RECT 11.765 68.255 12.300 68.875 ;
        RECT 12.595 68.425 12.765 68.925 ;
        RECT 13.025 68.595 13.195 69.055 ;
        RECT 13.425 68.675 14.850 68.845 ;
        RECT 13.425 68.425 13.755 68.675 ;
        RECT 12.595 68.255 13.755 68.425 ;
        RECT 13.980 68.085 14.310 68.505 ;
        RECT 14.565 68.255 14.850 68.675 ;
        RECT 15.095 68.085 15.425 68.885 ;
        RECT 15.755 68.805 16.010 70.160 ;
        RECT 15.675 68.295 16.010 68.805 ;
        RECT 16.185 69.690 16.525 70.465 ;
        RECT 16.695 70.175 16.865 70.635 ;
        RECT 17.105 70.200 17.465 70.465 ;
        RECT 17.105 70.195 17.460 70.200 ;
        RECT 17.105 70.185 17.455 70.195 ;
        RECT 17.105 70.180 17.450 70.185 ;
        RECT 17.105 70.170 17.445 70.180 ;
        RECT 18.095 70.175 18.265 70.635 ;
        RECT 17.105 70.165 17.440 70.170 ;
        RECT 17.105 70.155 17.430 70.165 ;
        RECT 17.105 70.145 17.420 70.155 ;
        RECT 17.105 70.005 17.405 70.145 ;
        RECT 16.695 69.815 17.405 70.005 ;
        RECT 17.595 70.005 17.925 70.085 ;
        RECT 18.435 70.005 18.775 70.465 ;
        RECT 17.595 69.815 18.775 70.005 ;
        RECT 18.945 69.835 19.640 70.465 ;
        RECT 19.845 69.835 20.155 70.635 ;
        RECT 20.325 70.135 20.585 70.465 ;
        RECT 20.755 70.275 21.085 70.635 ;
        RECT 21.340 70.255 22.640 70.465 ;
        RECT 16.185 68.255 16.465 69.690 ;
        RECT 16.695 69.245 16.980 69.815 ;
        RECT 17.165 69.415 17.635 69.645 ;
        RECT 17.805 69.625 18.135 69.645 ;
        RECT 17.805 69.445 18.255 69.625 ;
        RECT 18.445 69.445 18.775 69.645 ;
        RECT 16.695 69.030 17.845 69.245 ;
        RECT 16.635 68.085 17.345 68.860 ;
        RECT 17.515 68.255 17.845 69.030 ;
        RECT 18.040 68.330 18.255 69.445 ;
        RECT 18.545 69.105 18.775 69.445 ;
        RECT 18.965 69.395 19.300 69.645 ;
        RECT 19.470 69.235 19.640 69.835 ;
        RECT 19.810 69.395 20.145 69.665 ;
        RECT 18.435 68.085 18.765 68.805 ;
        RECT 18.945 68.085 19.205 69.225 ;
        RECT 19.375 68.255 19.705 69.235 ;
        RECT 19.875 68.085 20.155 69.225 ;
        RECT 20.325 68.935 20.495 70.135 ;
        RECT 21.340 70.105 21.510 70.255 ;
        RECT 20.755 69.980 21.510 70.105 ;
        RECT 20.665 69.935 21.510 69.980 ;
        RECT 20.665 69.815 20.935 69.935 ;
        RECT 20.665 69.240 20.835 69.815 ;
        RECT 21.065 69.375 21.475 69.680 ;
        RECT 21.765 69.645 21.975 70.045 ;
        RECT 21.645 69.435 21.975 69.645 ;
        RECT 22.220 69.645 22.440 70.045 ;
        RECT 22.915 69.870 23.370 70.635 ;
        RECT 23.545 70.135 23.805 70.465 ;
        RECT 23.975 70.275 24.305 70.635 ;
        RECT 24.560 70.255 25.860 70.465 ;
        RECT 22.220 69.435 22.695 69.645 ;
        RECT 22.885 69.445 23.375 69.645 ;
        RECT 20.665 69.205 20.865 69.240 ;
        RECT 22.195 69.205 23.370 69.265 ;
        RECT 20.665 69.095 23.370 69.205 ;
        RECT 20.725 69.035 22.525 69.095 ;
        RECT 22.195 69.005 22.525 69.035 ;
        RECT 20.325 68.255 20.585 68.935 ;
        RECT 20.755 68.085 21.005 68.865 ;
        RECT 21.255 68.835 22.090 68.845 ;
        RECT 22.680 68.835 22.865 68.925 ;
        RECT 21.255 68.635 22.865 68.835 ;
        RECT 21.255 68.255 21.505 68.635 ;
        RECT 22.635 68.595 22.865 68.635 ;
        RECT 23.115 68.475 23.370 69.095 ;
        RECT 21.675 68.085 22.030 68.465 ;
        RECT 23.035 68.255 23.370 68.475 ;
        RECT 23.545 68.935 23.715 70.135 ;
        RECT 24.560 70.105 24.730 70.255 ;
        RECT 23.975 69.980 24.730 70.105 ;
        RECT 23.885 69.935 24.730 69.980 ;
        RECT 23.885 69.815 24.155 69.935 ;
        RECT 23.885 69.240 24.055 69.815 ;
        RECT 24.285 69.375 24.695 69.680 ;
        RECT 24.985 69.645 25.195 70.045 ;
        RECT 24.865 69.435 25.195 69.645 ;
        RECT 25.440 69.645 25.660 70.045 ;
        RECT 26.135 69.870 26.590 70.635 ;
        RECT 26.770 70.105 27.060 70.455 ;
        RECT 27.255 70.275 27.585 70.635 ;
        RECT 27.755 70.105 27.985 70.410 ;
        RECT 26.770 69.935 27.985 70.105 ;
        RECT 28.175 70.295 28.345 70.330 ;
        RECT 28.175 70.125 28.375 70.295 ;
        RECT 28.665 70.155 28.945 70.635 ;
        RECT 28.175 69.765 28.345 70.125 ;
        RECT 29.115 69.985 29.375 70.375 ;
        RECT 29.550 70.155 29.805 70.635 ;
        RECT 29.975 69.985 30.270 70.375 ;
        RECT 30.450 70.155 30.725 70.635 ;
        RECT 30.895 70.135 31.195 70.465 ;
        RECT 25.440 69.435 25.915 69.645 ;
        RECT 26.105 69.445 26.595 69.645 ;
        RECT 26.830 69.615 27.090 69.725 ;
        RECT 26.825 69.445 27.090 69.615 ;
        RECT 26.830 69.395 27.090 69.445 ;
        RECT 27.270 69.395 27.655 69.725 ;
        RECT 27.825 69.595 28.345 69.765 ;
        RECT 28.620 69.815 30.270 69.985 ;
        RECT 23.885 69.205 24.085 69.240 ;
        RECT 25.415 69.205 26.590 69.265 ;
        RECT 23.885 69.095 26.590 69.205 ;
        RECT 23.945 69.035 25.745 69.095 ;
        RECT 25.415 69.005 25.745 69.035 ;
        RECT 23.545 68.255 23.805 68.935 ;
        RECT 23.975 68.085 24.225 68.865 ;
        RECT 24.475 68.835 25.310 68.845 ;
        RECT 25.900 68.835 26.085 68.925 ;
        RECT 24.475 68.635 26.085 68.835 ;
        RECT 24.475 68.255 24.725 68.635 ;
        RECT 25.855 68.595 26.085 68.635 ;
        RECT 26.335 68.475 26.590 69.095 ;
        RECT 24.895 68.085 25.250 68.465 ;
        RECT 26.255 68.255 26.590 68.475 ;
        RECT 26.770 68.085 27.090 69.225 ;
        RECT 27.270 68.345 27.465 69.395 ;
        RECT 27.825 69.215 27.995 69.595 ;
        RECT 27.645 68.935 27.995 69.215 ;
        RECT 28.185 69.065 28.430 69.425 ;
        RECT 28.620 69.305 29.025 69.815 ;
        RECT 29.195 69.475 30.335 69.645 ;
        RECT 28.620 69.135 29.375 69.305 ;
        RECT 27.645 68.255 27.975 68.935 ;
        RECT 28.175 68.085 28.430 68.885 ;
        RECT 28.660 68.085 28.945 68.955 ;
        RECT 29.115 68.885 29.375 69.135 ;
        RECT 30.165 69.225 30.335 69.475 ;
        RECT 30.505 69.395 30.855 69.965 ;
        RECT 31.025 69.225 31.195 70.135 ;
        RECT 31.365 69.910 31.655 70.635 ;
        RECT 31.825 69.895 32.140 70.270 ;
        RECT 32.395 69.895 32.565 70.635 ;
        RECT 32.815 70.065 32.985 70.270 ;
        RECT 33.255 70.240 33.585 70.635 ;
        RECT 33.835 70.065 34.005 70.415 ;
        RECT 34.205 70.235 34.535 70.635 ;
        RECT 34.705 70.065 34.875 70.415 ;
        RECT 35.095 70.235 35.475 70.635 ;
        RECT 32.815 69.895 33.335 70.065 ;
        RECT 30.165 69.055 31.195 69.225 ;
        RECT 29.115 68.715 30.235 68.885 ;
        RECT 29.115 68.255 29.375 68.715 ;
        RECT 29.550 68.085 29.805 68.545 ;
        RECT 29.975 68.255 30.235 68.715 ;
        RECT 30.405 68.085 30.715 68.885 ;
        RECT 30.885 68.255 31.195 69.055 ;
        RECT 31.365 68.085 31.655 69.250 ;
        RECT 31.825 68.855 31.995 69.895 ;
        RECT 33.145 69.725 33.335 69.895 ;
        RECT 33.675 69.895 35.485 70.065 ;
        RECT 32.165 69.025 32.515 69.725 ;
        RECT 32.685 69.395 32.975 69.725 ;
        RECT 33.145 69.395 33.435 69.725 ;
        RECT 33.145 69.195 33.335 69.395 ;
        RECT 32.730 69.025 33.335 69.195 ;
        RECT 31.825 68.685 33.035 68.855 ;
        RECT 33.675 68.765 33.845 69.895 ;
        RECT 31.825 68.265 32.085 68.685 ;
        RECT 32.255 68.085 32.585 68.515 ;
        RECT 32.865 68.425 33.035 68.685 ;
        RECT 33.250 68.595 33.845 68.765 ;
        RECT 34.015 68.425 34.185 69.725 ;
        RECT 34.415 69.270 34.745 69.725 ;
        RECT 32.865 68.255 34.185 68.425 ;
        RECT 34.535 68.935 34.745 69.270 ;
        RECT 34.975 69.275 35.145 69.725 ;
        RECT 35.315 69.645 35.485 69.895 ;
        RECT 35.655 69.995 35.905 70.465 ;
        RECT 36.075 70.165 36.245 70.635 ;
        RECT 36.415 69.995 36.745 70.465 ;
        RECT 36.915 70.165 37.085 70.635 ;
        RECT 37.355 70.295 37.690 70.465 ;
        RECT 35.655 69.815 37.175 69.995 ;
        RECT 37.355 69.895 37.970 70.295 ;
        RECT 38.650 70.255 38.985 70.635 ;
        RECT 39.575 70.195 39.810 70.635 ;
        RECT 39.980 70.105 40.310 70.465 ;
        RECT 40.480 70.275 40.810 70.635 ;
        RECT 38.140 69.895 39.410 70.085 ;
        RECT 39.980 69.935 40.800 70.105 ;
        RECT 41.025 70.090 46.370 70.635 ;
        RECT 35.315 69.475 36.775 69.645 ;
        RECT 34.975 69.105 35.410 69.275 ;
        RECT 36.485 69.265 36.655 69.275 ;
        RECT 36.945 69.265 37.175 69.815 ;
        RECT 37.345 69.395 37.620 69.725 ;
        RECT 35.615 69.095 37.175 69.265 ;
        RECT 37.790 69.210 37.970 69.895 ;
        RECT 38.140 69.395 38.500 69.725 ;
        RECT 38.790 69.615 39.080 69.725 ;
        RECT 38.785 69.445 39.080 69.615 ;
        RECT 38.790 69.395 39.080 69.445 ;
        RECT 39.250 69.395 39.585 69.725 ;
        RECT 39.755 69.395 40.435 69.725 ;
        RECT 39.755 69.210 39.925 69.395 ;
        RECT 34.535 68.345 34.855 68.935 ;
        RECT 35.140 68.085 35.390 68.925 ;
        RECT 35.615 68.255 35.865 69.095 ;
        RECT 36.035 68.085 36.285 68.925 ;
        RECT 36.455 68.255 36.705 69.095 ;
        RECT 37.350 68.955 39.925 69.210 ;
        RECT 36.875 68.085 37.125 68.925 ;
        RECT 37.350 68.255 37.615 68.955 ;
        RECT 37.785 68.085 38.115 68.785 ;
        RECT 38.285 68.255 38.955 68.955 ;
        RECT 40.605 68.815 40.800 69.935 ;
        RECT 42.610 69.260 42.950 70.090 ;
        RECT 46.545 69.865 49.135 70.635 ;
        RECT 49.305 70.295 50.665 70.465 ;
        RECT 39.460 68.085 39.890 68.785 ;
        RECT 40.070 68.645 40.800 68.815 ;
        RECT 40.070 68.255 40.260 68.645 ;
        RECT 44.430 68.520 44.780 69.770 ;
        RECT 46.545 69.345 47.755 69.865 ;
        RECT 49.305 69.815 49.665 70.295 ;
        RECT 49.835 69.895 50.165 70.125 ;
        RECT 50.335 70.065 50.665 70.295 ;
        RECT 50.835 70.235 51.165 70.635 ;
        RECT 51.335 70.065 51.665 70.465 ;
        RECT 50.335 69.895 51.665 70.065 ;
        RECT 51.935 69.895 52.265 70.635 ;
        RECT 47.925 69.175 49.135 69.695 ;
        RECT 49.305 69.475 49.665 69.645 ;
        RECT 49.305 69.395 49.635 69.475 ;
        RECT 40.430 68.085 40.760 68.465 ;
        RECT 41.025 68.085 46.370 68.520 ;
        RECT 46.545 68.085 49.135 69.175 ;
        RECT 49.305 68.085 49.665 69.225 ;
        RECT 49.835 68.935 50.035 69.895 ;
        RECT 50.205 69.275 50.450 69.725 ;
        RECT 50.205 69.105 50.455 69.275 ;
        RECT 50.725 69.105 50.945 69.725 ;
        RECT 51.200 69.105 51.375 69.725 ;
        RECT 51.645 69.105 51.865 69.725 ;
        RECT 52.035 68.935 52.345 69.725 ;
        RECT 49.835 68.765 52.345 68.935 ;
        RECT 50.335 68.255 50.665 68.765 ;
        RECT 51.835 68.085 52.345 68.595 ;
        RECT 52.515 68.255 52.845 70.465 ;
        RECT 53.015 69.835 53.275 70.635 ;
        RECT 53.625 70.255 53.955 70.635 ;
        RECT 54.125 70.085 54.315 70.465 ;
        RECT 54.485 70.275 54.815 70.635 ;
        RECT 53.915 69.895 54.315 70.085 ;
        RECT 55.035 70.065 55.225 70.465 ;
        RECT 54.485 69.895 55.225 70.065 ;
        RECT 53.015 68.085 53.275 69.225 ;
        RECT 53.455 68.085 53.745 69.055 ;
        RECT 53.915 68.255 54.145 69.895 ;
        RECT 54.485 69.725 54.655 69.895 ;
        RECT 54.315 69.030 54.655 69.725 ;
        RECT 54.825 69.310 55.150 69.725 ;
        RECT 55.600 69.395 55.980 70.355 ;
        RECT 56.165 70.155 56.495 70.635 ;
        RECT 56.170 69.395 56.485 69.970 ;
        RECT 57.125 69.910 57.415 70.635 ;
        RECT 57.585 70.125 57.890 70.635 ;
        RECT 57.585 69.395 57.900 69.955 ;
        RECT 58.070 69.645 58.320 70.455 ;
        RECT 58.490 70.110 58.750 70.635 ;
        RECT 58.930 69.645 59.180 70.455 ;
        RECT 59.350 70.075 59.610 70.635 ;
        RECT 59.780 69.985 60.040 70.440 ;
        RECT 60.210 70.155 60.470 70.635 ;
        RECT 60.640 69.985 60.900 70.440 ;
        RECT 61.070 70.155 61.330 70.635 ;
        RECT 61.500 69.985 61.760 70.440 ;
        RECT 61.930 70.155 62.175 70.635 ;
        RECT 62.345 69.985 62.620 70.440 ;
        RECT 62.790 70.155 63.035 70.635 ;
        RECT 63.205 69.985 63.465 70.440 ;
        RECT 63.645 70.155 63.895 70.635 ;
        RECT 64.065 69.985 64.325 70.440 ;
        RECT 64.505 70.155 64.755 70.635 ;
        RECT 64.925 69.985 65.185 70.440 ;
        RECT 65.365 70.155 65.625 70.635 ;
        RECT 65.795 69.985 66.055 70.440 ;
        RECT 66.225 70.155 66.525 70.635 ;
        RECT 59.780 69.815 66.525 69.985 ;
        RECT 66.785 69.815 67.080 70.635 ;
        RECT 67.250 69.895 67.690 70.455 ;
        RECT 67.860 69.895 68.310 70.635 ;
        RECT 68.480 70.065 68.650 70.465 ;
        RECT 68.820 70.235 69.240 70.635 ;
        RECT 69.410 70.065 69.640 70.465 ;
        RECT 68.480 69.895 69.640 70.065 ;
        RECT 69.810 69.895 70.295 70.465 ;
        RECT 58.070 69.395 65.190 69.645 ;
        RECT 54.315 68.800 55.150 69.030 ;
        RECT 54.315 68.085 54.645 68.500 ;
        RECT 54.835 68.255 55.150 68.800 ;
        RECT 55.320 68.785 56.435 69.050 ;
        RECT 55.320 68.255 55.545 68.785 ;
        RECT 55.715 68.085 56.045 68.595 ;
        RECT 56.215 68.255 56.435 68.785 ;
        RECT 57.125 68.085 57.415 69.250 ;
        RECT 57.595 68.085 57.890 68.895 ;
        RECT 58.070 68.255 58.315 69.395 ;
        RECT 58.490 68.085 58.750 68.895 ;
        RECT 58.930 68.260 59.180 69.395 ;
        RECT 65.360 69.225 66.525 69.815 ;
        RECT 67.250 69.645 67.560 69.895 ;
        RECT 66.785 69.425 67.560 69.645 ;
        RECT 59.780 69.000 66.525 69.225 ;
        RECT 59.780 68.985 65.185 69.000 ;
        RECT 59.350 68.090 59.610 68.885 ;
        RECT 59.780 68.260 60.040 68.985 ;
        RECT 60.210 68.090 60.470 68.815 ;
        RECT 60.640 68.260 60.900 68.985 ;
        RECT 61.070 68.090 61.330 68.815 ;
        RECT 61.500 68.260 61.760 68.985 ;
        RECT 61.930 68.090 62.190 68.815 ;
        RECT 62.360 68.260 62.620 68.985 ;
        RECT 62.790 68.090 63.035 68.815 ;
        RECT 63.205 68.260 63.465 68.985 ;
        RECT 63.650 68.090 63.895 68.815 ;
        RECT 64.065 68.260 64.325 68.985 ;
        RECT 64.510 68.090 64.755 68.815 ;
        RECT 64.925 68.260 65.185 68.985 ;
        RECT 65.370 68.090 65.625 68.815 ;
        RECT 65.795 68.260 66.085 69.000 ;
        RECT 59.350 68.085 65.625 68.090 ;
        RECT 66.255 68.085 66.525 68.830 ;
        RECT 66.785 68.085 67.080 69.255 ;
        RECT 67.250 68.885 67.560 69.425 ;
        RECT 67.730 69.275 67.900 69.725 ;
        RECT 68.070 69.445 68.460 69.725 ;
        RECT 68.645 69.395 68.890 69.725 ;
        RECT 67.730 69.105 68.520 69.275 ;
        RECT 67.250 68.255 67.690 68.885 ;
        RECT 67.865 68.085 68.180 68.935 ;
        RECT 68.350 68.425 68.520 69.105 ;
        RECT 68.690 68.595 68.890 69.395 ;
        RECT 69.090 68.595 69.340 69.725 ;
        RECT 69.555 69.395 69.955 69.725 ;
        RECT 70.125 69.225 70.295 69.895 ;
        RECT 70.465 69.815 70.760 70.635 ;
        RECT 70.930 69.895 71.370 70.455 ;
        RECT 71.540 69.895 71.990 70.635 ;
        RECT 72.160 70.065 72.330 70.465 ;
        RECT 72.500 70.235 72.920 70.635 ;
        RECT 73.090 70.065 73.320 70.465 ;
        RECT 72.160 69.895 73.320 70.065 ;
        RECT 73.490 69.895 73.975 70.465 ;
        RECT 70.930 69.645 71.240 69.895 ;
        RECT 70.465 69.425 71.240 69.645 ;
        RECT 69.530 69.055 70.295 69.225 ;
        RECT 69.530 68.425 69.780 69.055 ;
        RECT 68.350 68.255 69.780 68.425 ;
        RECT 69.955 68.085 70.290 68.885 ;
        RECT 70.465 68.085 70.760 69.255 ;
        RECT 70.930 68.885 71.240 69.425 ;
        RECT 71.410 69.275 71.580 69.725 ;
        RECT 71.750 69.445 72.140 69.725 ;
        RECT 72.325 69.395 72.570 69.725 ;
        RECT 71.410 69.105 72.200 69.275 ;
        RECT 70.930 68.255 71.370 68.885 ;
        RECT 71.545 68.085 71.860 68.935 ;
        RECT 72.030 68.425 72.200 69.105 ;
        RECT 72.370 68.595 72.570 69.395 ;
        RECT 72.770 68.595 73.020 69.725 ;
        RECT 73.235 69.395 73.635 69.725 ;
        RECT 73.805 69.225 73.975 69.895 ;
        RECT 74.145 69.835 74.840 70.465 ;
        RECT 75.045 69.835 75.355 70.635 ;
        RECT 75.525 69.885 76.735 70.635 ;
        RECT 74.665 69.785 74.840 69.835 ;
        RECT 74.165 69.395 74.500 69.645 ;
        RECT 74.670 69.235 74.840 69.785 ;
        RECT 75.010 69.395 75.345 69.665 ;
        RECT 73.210 69.055 73.975 69.225 ;
        RECT 73.210 68.425 73.460 69.055 ;
        RECT 72.030 68.255 73.460 68.425 ;
        RECT 73.635 68.085 73.970 68.885 ;
        RECT 74.145 68.085 74.405 69.225 ;
        RECT 74.575 68.255 74.905 69.235 ;
        RECT 75.075 68.085 75.355 69.225 ;
        RECT 75.525 69.175 76.045 69.715 ;
        RECT 76.215 69.345 76.735 69.885 ;
        RECT 75.525 68.085 76.735 69.175 ;
        RECT 5.520 67.915 76.820 68.085 ;
        RECT 5.605 66.825 6.815 67.915 ;
        RECT 5.605 66.115 6.125 66.655 ;
        RECT 6.295 66.285 6.815 66.825 ;
        RECT 7.995 66.985 8.165 67.745 ;
        RECT 8.380 67.155 8.710 67.915 ;
        RECT 7.995 66.815 8.710 66.985 ;
        RECT 8.880 66.840 9.135 67.745 ;
        RECT 7.905 66.265 8.260 66.635 ;
        RECT 8.540 66.605 8.710 66.815 ;
        RECT 8.540 66.275 8.795 66.605 ;
        RECT 5.605 65.365 6.815 66.115 ;
        RECT 8.540 66.085 8.710 66.275 ;
        RECT 8.965 66.110 9.135 66.840 ;
        RECT 9.310 66.765 9.570 67.915 ;
        RECT 9.750 66.765 10.010 67.915 ;
        RECT 10.185 66.840 10.440 67.745 ;
        RECT 10.610 67.155 10.940 67.915 ;
        RECT 11.155 66.985 11.325 67.745 ;
        RECT 7.995 65.915 8.710 66.085 ;
        RECT 7.995 65.535 8.165 65.915 ;
        RECT 8.380 65.365 8.710 65.745 ;
        RECT 8.880 65.535 9.135 66.110 ;
        RECT 9.310 65.365 9.570 66.205 ;
        RECT 9.750 65.365 10.010 66.205 ;
        RECT 10.185 66.110 10.355 66.840 ;
        RECT 10.610 66.815 11.325 66.985 ;
        RECT 11.590 67.195 11.925 67.705 ;
        RECT 10.610 66.605 10.780 66.815 ;
        RECT 10.525 66.275 10.780 66.605 ;
        RECT 10.185 65.535 10.440 66.110 ;
        RECT 10.610 66.085 10.780 66.275 ;
        RECT 11.060 66.265 11.415 66.635 ;
        RECT 10.610 65.915 11.325 66.085 ;
        RECT 10.610 65.365 10.940 65.745 ;
        RECT 11.155 65.535 11.325 65.915 ;
        RECT 11.590 65.840 11.845 67.195 ;
        RECT 12.175 67.115 12.505 67.915 ;
        RECT 12.750 67.325 13.035 67.745 ;
        RECT 13.290 67.495 13.620 67.915 ;
        RECT 13.845 67.575 15.005 67.745 ;
        RECT 13.845 67.325 14.175 67.575 ;
        RECT 12.750 67.155 14.175 67.325 ;
        RECT 14.405 66.945 14.575 67.405 ;
        RECT 14.835 67.075 15.005 67.575 ;
        RECT 12.205 66.775 14.575 66.945 ;
        RECT 12.205 66.605 12.375 66.775 ;
        RECT 14.825 66.605 15.030 66.895 ;
        RECT 12.070 66.275 12.375 66.605 ;
        RECT 12.570 66.555 12.820 66.605 ;
        RECT 13.030 66.555 13.300 66.605 ;
        RECT 12.565 66.385 12.820 66.555 ;
        RECT 13.025 66.385 13.300 66.555 ;
        RECT 12.570 66.275 12.820 66.385 ;
        RECT 12.205 66.105 12.375 66.275 ;
        RECT 12.205 65.935 12.765 66.105 ;
        RECT 13.030 65.945 13.300 66.385 ;
        RECT 13.490 66.215 13.780 66.605 ;
        RECT 13.485 66.045 13.780 66.215 ;
        RECT 13.490 65.945 13.780 66.045 ;
        RECT 13.950 65.940 14.370 66.605 ;
        RECT 14.680 66.555 15.030 66.605 ;
        RECT 14.680 66.385 15.035 66.555 ;
        RECT 14.680 66.275 15.030 66.385 ;
        RECT 11.590 65.580 11.925 65.840 ;
        RECT 12.595 65.765 12.765 65.935 ;
        RECT 12.095 65.365 12.425 65.765 ;
        RECT 12.595 65.595 14.210 65.765 ;
        RECT 14.755 65.365 15.085 66.085 ;
        RECT 15.275 65.545 15.535 67.735 ;
        RECT 15.705 67.185 16.045 67.915 ;
        RECT 16.225 67.005 16.495 67.735 ;
        RECT 15.725 66.785 16.495 67.005 ;
        RECT 16.675 67.025 16.905 67.735 ;
        RECT 17.075 67.205 17.405 67.915 ;
        RECT 17.575 67.025 17.835 67.735 ;
        RECT 16.675 66.785 17.835 67.025 ;
        RECT 15.725 66.115 16.015 66.785 ;
        RECT 18.485 66.750 18.775 67.915 ;
        RECT 18.955 66.965 19.230 67.735 ;
        RECT 19.400 67.305 19.730 67.735 ;
        RECT 19.900 67.475 20.095 67.915 ;
        RECT 20.275 67.305 20.605 67.735 ;
        RECT 19.400 67.135 20.605 67.305 ;
        RECT 18.955 66.775 19.540 66.965 ;
        RECT 19.710 66.805 20.605 67.135 ;
        RECT 16.195 66.295 16.660 66.605 ;
        RECT 16.840 66.295 17.365 66.605 ;
        RECT 15.725 65.915 16.955 66.115 ;
        RECT 15.795 65.365 16.465 65.735 ;
        RECT 16.645 65.545 16.955 65.915 ;
        RECT 17.135 65.655 17.365 66.295 ;
        RECT 17.545 66.275 17.845 66.605 ;
        RECT 17.545 65.365 17.835 66.095 ;
        RECT 18.485 65.365 18.775 66.090 ;
        RECT 18.955 65.955 19.195 66.605 ;
        RECT 19.365 66.105 19.540 66.775 ;
        RECT 20.790 66.765 21.050 67.915 ;
        RECT 21.225 66.840 21.480 67.745 ;
        RECT 21.650 67.155 21.980 67.915 ;
        RECT 22.195 66.985 22.365 67.745 ;
        RECT 19.710 66.275 20.125 66.605 ;
        RECT 20.305 66.275 20.600 66.605 ;
        RECT 19.365 65.925 19.695 66.105 ;
        RECT 18.970 65.365 19.300 65.755 ;
        RECT 19.470 65.545 19.695 65.925 ;
        RECT 19.895 65.655 20.125 66.275 ;
        RECT 20.305 65.365 20.605 66.095 ;
        RECT 20.790 65.365 21.050 66.205 ;
        RECT 21.225 66.110 21.395 66.840 ;
        RECT 21.650 66.815 22.365 66.985 ;
        RECT 22.780 66.905 23.080 67.745 ;
        RECT 23.275 67.075 23.525 67.915 ;
        RECT 24.115 67.325 24.920 67.745 ;
        RECT 23.695 67.155 25.260 67.325 ;
        RECT 23.695 66.905 23.865 67.155 ;
        RECT 21.650 66.605 21.820 66.815 ;
        RECT 22.780 66.735 23.865 66.905 ;
        RECT 21.565 66.275 21.820 66.605 ;
        RECT 21.225 65.535 21.480 66.110 ;
        RECT 21.650 66.085 21.820 66.275 ;
        RECT 22.100 66.265 22.455 66.635 ;
        RECT 22.625 66.275 22.955 66.565 ;
        RECT 23.125 66.105 23.295 66.735 ;
        RECT 24.035 66.605 24.355 66.985 ;
        RECT 24.545 66.895 24.920 66.985 ;
        RECT 24.525 66.725 24.920 66.895 ;
        RECT 25.090 66.905 25.260 67.155 ;
        RECT 25.430 67.075 25.760 67.915 ;
        RECT 25.930 67.155 26.595 67.745 ;
        RECT 27.775 67.170 28.045 67.915 ;
        RECT 28.675 67.910 34.950 67.915 ;
        RECT 25.090 66.735 26.010 66.905 ;
        RECT 23.465 66.355 23.795 66.565 ;
        RECT 23.975 66.355 24.355 66.605 ;
        RECT 24.545 66.565 24.920 66.725 ;
        RECT 25.840 66.565 26.010 66.735 ;
        RECT 24.545 66.355 25.030 66.565 ;
        RECT 25.220 66.355 25.670 66.565 ;
        RECT 25.840 66.355 26.175 66.565 ;
        RECT 26.345 66.185 26.595 67.155 ;
        RECT 28.215 67.000 28.505 67.740 ;
        RECT 28.675 67.185 28.930 67.910 ;
        RECT 29.115 67.015 29.375 67.740 ;
        RECT 29.545 67.185 29.790 67.910 ;
        RECT 29.975 67.015 30.235 67.740 ;
        RECT 30.405 67.185 30.650 67.910 ;
        RECT 30.835 67.015 31.095 67.740 ;
        RECT 31.265 67.185 31.510 67.910 ;
        RECT 31.680 67.015 31.940 67.740 ;
        RECT 32.110 67.185 32.370 67.910 ;
        RECT 32.540 67.015 32.800 67.740 ;
        RECT 32.970 67.185 33.230 67.910 ;
        RECT 33.400 67.015 33.660 67.740 ;
        RECT 33.830 67.185 34.090 67.910 ;
        RECT 34.260 67.015 34.520 67.740 ;
        RECT 34.690 67.115 34.950 67.910 ;
        RECT 29.115 67.000 34.520 67.015 ;
        RECT 21.650 65.915 22.365 66.085 ;
        RECT 21.650 65.365 21.980 65.745 ;
        RECT 22.195 65.535 22.365 65.915 ;
        RECT 22.785 65.925 23.295 66.105 ;
        RECT 23.700 66.015 25.400 66.185 ;
        RECT 23.700 65.925 24.085 66.015 ;
        RECT 22.785 65.535 23.115 65.925 ;
        RECT 23.285 65.585 24.470 65.755 ;
        RECT 24.730 65.365 24.900 65.835 ;
        RECT 25.070 65.550 25.400 66.015 ;
        RECT 25.570 65.365 25.740 66.185 ;
        RECT 25.910 65.545 26.595 66.185 ;
        RECT 27.775 66.775 34.520 67.000 ;
        RECT 27.775 66.185 28.940 66.775 ;
        RECT 35.120 66.605 35.370 67.740 ;
        RECT 35.550 67.105 35.810 67.915 ;
        RECT 35.985 66.605 36.230 67.745 ;
        RECT 36.410 67.105 36.705 67.915 ;
        RECT 36.885 66.775 37.145 67.915 ;
        RECT 29.110 66.355 36.230 66.605 ;
        RECT 27.775 66.015 34.520 66.185 ;
        RECT 27.775 65.365 28.075 65.845 ;
        RECT 28.245 65.560 28.505 66.015 ;
        RECT 28.675 65.365 28.935 65.845 ;
        RECT 29.115 65.560 29.375 66.015 ;
        RECT 29.545 65.365 29.795 65.845 ;
        RECT 29.975 65.560 30.235 66.015 ;
        RECT 30.405 65.365 30.655 65.845 ;
        RECT 30.835 65.560 31.095 66.015 ;
        RECT 31.265 65.365 31.510 65.845 ;
        RECT 31.680 65.560 31.955 66.015 ;
        RECT 32.125 65.365 32.370 65.845 ;
        RECT 32.540 65.560 32.800 66.015 ;
        RECT 32.970 65.365 33.230 65.845 ;
        RECT 33.400 65.560 33.660 66.015 ;
        RECT 33.830 65.365 34.090 65.845 ;
        RECT 34.260 65.560 34.520 66.015 ;
        RECT 34.690 65.365 34.950 65.925 ;
        RECT 35.120 65.545 35.370 66.355 ;
        RECT 35.550 65.365 35.810 65.890 ;
        RECT 35.980 65.545 36.230 66.355 ;
        RECT 36.400 66.045 36.715 66.605 ;
        RECT 36.410 65.365 36.715 65.875 ;
        RECT 36.885 65.365 37.145 66.165 ;
        RECT 37.315 65.535 37.645 67.745 ;
        RECT 37.815 67.405 38.325 67.915 ;
        RECT 39.495 67.235 39.825 67.745 ;
        RECT 37.815 67.065 40.325 67.235 ;
        RECT 37.815 66.275 38.125 67.065 ;
        RECT 38.295 66.275 38.515 66.895 ;
        RECT 38.785 66.275 38.960 66.895 ;
        RECT 39.215 66.275 39.435 66.895 ;
        RECT 39.705 66.725 39.955 66.895 ;
        RECT 39.710 66.275 39.955 66.725 ;
        RECT 40.125 66.105 40.325 67.065 ;
        RECT 40.495 66.775 40.855 67.915 ;
        RECT 41.025 66.735 41.345 67.915 ;
        RECT 41.515 66.895 41.715 67.685 ;
        RECT 42.040 67.085 42.425 67.745 ;
        RECT 42.820 67.155 43.605 67.915 ;
        RECT 42.015 66.985 42.425 67.085 ;
        RECT 41.515 66.725 41.845 66.895 ;
        RECT 42.015 66.775 43.625 66.985 ;
        RECT 41.665 66.605 41.845 66.725 ;
        RECT 40.525 66.525 40.855 66.605 ;
        RECT 40.495 66.355 40.855 66.525 ;
        RECT 41.025 66.355 41.490 66.555 ;
        RECT 41.665 66.355 41.995 66.605 ;
        RECT 42.165 66.555 42.630 66.605 ;
        RECT 42.165 66.385 42.635 66.555 ;
        RECT 42.165 66.355 42.630 66.385 ;
        RECT 42.825 66.355 43.180 66.605 ;
        RECT 37.895 65.365 38.225 66.105 ;
        RECT 38.495 65.935 39.825 66.105 ;
        RECT 38.495 65.535 38.825 65.935 ;
        RECT 38.995 65.365 39.325 65.765 ;
        RECT 39.495 65.705 39.825 65.935 ;
        RECT 39.995 65.875 40.325 66.105 ;
        RECT 40.495 65.705 40.855 66.185 ;
        RECT 43.350 66.175 43.625 66.775 ;
        RECT 39.495 65.535 40.855 65.705 ;
        RECT 41.025 65.975 42.205 66.145 ;
        RECT 41.025 65.560 41.365 65.975 ;
        RECT 41.535 65.365 41.705 65.805 ;
        RECT 41.875 65.755 42.205 65.975 ;
        RECT 42.375 65.995 43.625 66.175 ;
        RECT 42.375 65.925 42.740 65.995 ;
        RECT 41.875 65.575 43.125 65.755 ;
        RECT 43.395 65.365 43.565 65.825 ;
        RECT 43.795 65.645 44.075 67.745 ;
        RECT 44.245 66.750 44.535 67.915 ;
        RECT 44.795 67.170 45.065 67.915 ;
        RECT 45.695 67.910 51.970 67.915 ;
        RECT 45.235 67.000 45.525 67.740 ;
        RECT 45.695 67.185 45.950 67.910 ;
        RECT 46.135 67.015 46.395 67.740 ;
        RECT 46.565 67.185 46.810 67.910 ;
        RECT 46.995 67.015 47.255 67.740 ;
        RECT 47.425 67.185 47.670 67.910 ;
        RECT 47.855 67.015 48.115 67.740 ;
        RECT 48.285 67.185 48.530 67.910 ;
        RECT 48.700 67.015 48.960 67.740 ;
        RECT 49.130 67.185 49.390 67.910 ;
        RECT 49.560 67.015 49.820 67.740 ;
        RECT 49.990 67.185 50.250 67.910 ;
        RECT 50.420 67.015 50.680 67.740 ;
        RECT 50.850 67.185 51.110 67.910 ;
        RECT 51.280 67.015 51.540 67.740 ;
        RECT 51.710 67.115 51.970 67.910 ;
        RECT 46.135 67.000 51.540 67.015 ;
        RECT 44.795 66.775 51.540 67.000 ;
        RECT 44.795 66.185 45.960 66.775 ;
        RECT 52.140 66.605 52.390 67.740 ;
        RECT 52.570 67.105 52.830 67.915 ;
        RECT 53.005 66.605 53.250 67.745 ;
        RECT 53.430 67.105 53.725 67.915 ;
        RECT 53.995 67.575 55.155 67.745 ;
        RECT 53.995 67.075 54.165 67.575 ;
        RECT 54.425 66.945 54.595 67.405 ;
        RECT 54.825 67.325 55.155 67.575 ;
        RECT 55.380 67.495 55.710 67.915 ;
        RECT 55.965 67.325 56.250 67.745 ;
        RECT 54.825 67.155 56.250 67.325 ;
        RECT 56.495 67.115 56.825 67.915 ;
        RECT 57.075 67.195 57.410 67.705 ;
        RECT 53.970 66.605 54.175 66.895 ;
        RECT 54.425 66.775 56.795 66.945 ;
        RECT 56.625 66.605 56.795 66.775 ;
        RECT 46.130 66.355 53.250 66.605 ;
        RECT 44.245 65.365 44.535 66.090 ;
        RECT 44.795 66.015 51.540 66.185 ;
        RECT 44.795 65.365 45.095 65.845 ;
        RECT 45.265 65.560 45.525 66.015 ;
        RECT 45.695 65.365 45.955 65.845 ;
        RECT 46.135 65.560 46.395 66.015 ;
        RECT 46.565 65.365 46.815 65.845 ;
        RECT 46.995 65.560 47.255 66.015 ;
        RECT 47.425 65.365 47.675 65.845 ;
        RECT 47.855 65.560 48.115 66.015 ;
        RECT 48.285 65.365 48.530 65.845 ;
        RECT 48.700 65.560 48.975 66.015 ;
        RECT 49.145 65.365 49.390 65.845 ;
        RECT 49.560 65.560 49.820 66.015 ;
        RECT 49.990 65.365 50.250 65.845 ;
        RECT 50.420 65.560 50.680 66.015 ;
        RECT 50.850 65.365 51.110 65.845 ;
        RECT 51.280 65.560 51.540 66.015 ;
        RECT 51.710 65.365 51.970 65.925 ;
        RECT 52.140 65.545 52.390 66.355 ;
        RECT 52.570 65.365 52.830 65.890 ;
        RECT 53.000 65.545 53.250 66.355 ;
        RECT 53.420 66.045 53.735 66.605 ;
        RECT 53.970 66.555 54.320 66.605 ;
        RECT 53.965 66.385 54.320 66.555 ;
        RECT 53.970 66.275 54.320 66.385 ;
        RECT 53.430 65.365 53.735 65.875 ;
        RECT 53.915 65.365 54.245 66.085 ;
        RECT 54.630 65.940 55.050 66.605 ;
        RECT 55.220 66.215 55.510 66.605 ;
        RECT 55.700 66.555 55.970 66.605 ;
        RECT 56.180 66.555 56.430 66.605 ;
        RECT 55.700 66.385 55.975 66.555 ;
        RECT 56.180 66.385 56.435 66.555 ;
        RECT 55.220 66.045 55.515 66.215 ;
        RECT 55.220 65.945 55.510 66.045 ;
        RECT 55.700 65.945 55.970 66.385 ;
        RECT 56.180 66.275 56.430 66.385 ;
        RECT 56.625 66.275 56.930 66.605 ;
        RECT 56.625 66.105 56.795 66.275 ;
        RECT 56.235 65.935 56.795 66.105 ;
        RECT 56.235 65.765 56.405 65.935 ;
        RECT 57.155 65.840 57.410 67.195 ;
        RECT 57.675 66.945 57.845 67.745 ;
        RECT 58.135 67.285 58.385 67.705 ;
        RECT 58.575 67.455 58.905 67.915 ;
        RECT 59.115 67.285 59.365 67.705 ;
        RECT 58.075 67.115 59.365 67.285 ;
        RECT 59.535 67.115 59.785 67.915 ;
        RECT 59.955 67.285 60.125 67.745 ;
        RECT 60.335 67.455 60.585 67.915 ;
        RECT 59.955 67.115 60.630 67.285 ;
        RECT 60.895 67.170 61.165 67.915 ;
        RECT 61.795 67.910 68.070 67.915 ;
        RECT 57.675 66.775 60.165 66.945 ;
        RECT 57.630 66.035 57.825 66.605 ;
        RECT 54.790 65.595 56.405 65.765 ;
        RECT 56.575 65.365 56.905 65.765 ;
        RECT 57.075 65.580 57.410 65.840 ;
        RECT 57.585 65.365 57.845 65.845 ;
        RECT 58.015 65.785 58.185 66.775 ;
        RECT 58.365 66.150 58.535 66.605 ;
        RECT 58.925 66.525 59.095 66.540 ;
        RECT 58.765 66.355 59.095 66.525 ;
        RECT 58.365 65.980 58.755 66.150 ;
        RECT 58.015 65.615 58.345 65.785 ;
        RECT 58.545 65.695 58.755 65.980 ;
        RECT 58.925 66.145 59.095 66.355 ;
        RECT 59.325 66.275 59.655 66.605 ;
        RECT 59.995 66.525 60.165 66.775 ;
        RECT 59.835 66.355 60.165 66.525 ;
        RECT 58.925 65.975 59.190 66.145 ;
        RECT 59.450 66.040 59.655 66.275 ;
        RECT 60.375 66.165 60.630 67.115 ;
        RECT 61.335 67.000 61.625 67.740 ;
        RECT 61.795 67.185 62.050 67.910 ;
        RECT 62.235 67.015 62.495 67.740 ;
        RECT 62.665 67.185 62.910 67.910 ;
        RECT 63.095 67.015 63.355 67.740 ;
        RECT 63.525 67.185 63.770 67.910 ;
        RECT 63.955 67.015 64.215 67.740 ;
        RECT 64.385 67.185 64.630 67.910 ;
        RECT 64.800 67.015 65.060 67.740 ;
        RECT 65.230 67.185 65.490 67.910 ;
        RECT 65.660 67.015 65.920 67.740 ;
        RECT 66.090 67.185 66.350 67.910 ;
        RECT 66.520 67.015 66.780 67.740 ;
        RECT 66.950 67.185 67.210 67.910 ;
        RECT 67.380 67.015 67.640 67.740 ;
        RECT 67.810 67.115 68.070 67.910 ;
        RECT 62.235 67.000 67.640 67.015 ;
        RECT 59.020 65.875 59.190 65.975 ;
        RECT 59.955 65.995 60.630 66.165 ;
        RECT 60.895 66.775 67.640 67.000 ;
        RECT 60.895 66.185 62.060 66.775 ;
        RECT 68.240 66.605 68.490 67.740 ;
        RECT 68.670 67.105 68.930 67.915 ;
        RECT 69.105 66.605 69.350 67.745 ;
        RECT 69.530 67.105 69.825 67.915 ;
        RECT 70.005 66.750 70.295 67.915 ;
        RECT 70.470 66.915 70.725 67.915 ;
        RECT 62.230 66.355 69.350 66.605 ;
        RECT 60.895 66.015 67.640 66.185 ;
        RECT 59.020 65.705 59.195 65.875 ;
        RECT 59.535 65.745 59.705 65.825 ;
        RECT 59.020 65.680 59.190 65.705 ;
        RECT 58.015 65.535 58.260 65.615 ;
        RECT 59.435 65.365 59.765 65.745 ;
        RECT 59.955 65.535 60.125 65.995 ;
        RECT 60.375 65.365 60.630 65.825 ;
        RECT 60.895 65.365 61.195 65.845 ;
        RECT 61.365 65.560 61.625 66.015 ;
        RECT 61.795 65.365 62.055 65.845 ;
        RECT 62.235 65.560 62.495 66.015 ;
        RECT 62.665 65.365 62.915 65.845 ;
        RECT 63.095 65.560 63.355 66.015 ;
        RECT 63.525 65.365 63.775 65.845 ;
        RECT 63.955 65.560 64.215 66.015 ;
        RECT 64.385 65.365 64.630 65.845 ;
        RECT 64.800 65.560 65.075 66.015 ;
        RECT 65.245 65.365 65.490 65.845 ;
        RECT 65.660 65.560 65.920 66.015 ;
        RECT 66.090 65.365 66.350 65.845 ;
        RECT 66.520 65.560 66.780 66.015 ;
        RECT 66.950 65.365 67.210 65.845 ;
        RECT 67.380 65.560 67.640 66.015 ;
        RECT 67.810 65.365 68.070 65.925 ;
        RECT 68.240 65.545 68.490 66.355 ;
        RECT 68.670 65.365 68.930 65.890 ;
        RECT 69.100 65.545 69.350 66.355 ;
        RECT 69.520 66.045 69.835 66.605 ;
        RECT 69.530 65.365 69.835 65.875 ;
        RECT 70.005 65.365 70.295 66.090 ;
        RECT 70.485 65.365 70.725 66.165 ;
        RECT 70.910 65.535 71.155 67.745 ;
        RECT 71.325 67.465 72.175 67.915 ;
        RECT 72.345 67.285 72.605 67.745 ;
        RECT 71.485 67.065 72.605 67.285 ;
        RECT 71.485 66.610 71.655 67.065 ;
        RECT 71.325 66.120 71.655 66.610 ;
        RECT 71.825 66.290 72.235 66.895 ;
        RECT 72.785 66.680 72.990 67.265 ;
        RECT 73.175 66.930 73.500 67.915 ;
        RECT 73.695 67.305 74.025 67.735 ;
        RECT 74.205 67.475 74.400 67.915 ;
        RECT 74.570 67.305 74.900 67.735 ;
        RECT 73.695 67.135 74.900 67.305 ;
        RECT 73.695 66.805 74.590 67.135 ;
        RECT 75.070 66.965 75.345 67.735 ;
        RECT 74.760 66.775 75.345 66.965 ;
        RECT 75.525 66.825 76.735 67.915 ;
        RECT 72.405 66.555 72.990 66.680 ;
        RECT 72.405 66.385 72.995 66.555 ;
        RECT 72.405 66.305 72.990 66.385 ;
        RECT 73.245 66.275 73.505 66.730 ;
        RECT 73.700 66.275 73.995 66.605 ;
        RECT 74.175 66.275 74.590 66.605 ;
        RECT 71.325 65.915 72.175 66.120 ;
        RECT 71.325 65.365 71.655 65.745 ;
        RECT 71.845 65.535 72.175 65.915 ;
        RECT 72.345 65.915 73.500 66.105 ;
        RECT 72.345 65.745 72.555 65.915 ;
        RECT 73.225 65.775 73.500 65.915 ;
        RECT 72.725 65.365 73.055 65.745 ;
        RECT 73.695 65.365 73.995 66.095 ;
        RECT 74.175 65.655 74.405 66.275 ;
        RECT 74.760 66.105 74.935 66.775 ;
        RECT 74.605 65.925 74.935 66.105 ;
        RECT 75.105 65.955 75.345 66.605 ;
        RECT 75.525 66.285 76.045 66.825 ;
        RECT 76.215 66.115 76.735 66.655 ;
        RECT 74.605 65.545 74.830 65.925 ;
        RECT 75.000 65.365 75.330 65.755 ;
        RECT 75.525 65.365 76.735 66.115 ;
        RECT 5.520 65.195 76.820 65.365 ;
        RECT 5.605 64.445 6.815 65.195 ;
        RECT 5.605 63.905 6.125 64.445 ;
        RECT 6.990 64.355 7.250 65.195 ;
        RECT 7.425 64.450 7.680 65.025 ;
        RECT 7.850 64.815 8.180 65.195 ;
        RECT 8.395 64.645 8.565 65.025 ;
        RECT 7.850 64.475 8.565 64.645 ;
        RECT 9.375 64.645 9.545 65.025 ;
        RECT 9.725 64.815 10.055 65.195 ;
        RECT 9.375 64.475 10.040 64.645 ;
        RECT 10.235 64.520 10.495 65.025 ;
        RECT 6.295 63.735 6.815 64.275 ;
        RECT 5.605 62.645 6.815 63.735 ;
        RECT 6.990 62.645 7.250 63.795 ;
        RECT 7.425 63.720 7.595 64.450 ;
        RECT 7.850 64.285 8.020 64.475 ;
        RECT 7.765 63.955 8.020 64.285 ;
        RECT 7.850 63.745 8.020 63.955 ;
        RECT 8.300 63.925 8.655 64.295 ;
        RECT 9.305 63.925 9.645 64.295 ;
        RECT 9.870 64.220 10.040 64.475 ;
        RECT 9.870 63.890 10.145 64.220 ;
        RECT 9.870 63.745 10.040 63.890 ;
        RECT 7.425 62.815 7.680 63.720 ;
        RECT 7.850 63.575 8.565 63.745 ;
        RECT 7.850 62.645 8.180 63.405 ;
        RECT 8.395 62.815 8.565 63.575 ;
        RECT 9.365 63.575 10.040 63.745 ;
        RECT 10.315 63.720 10.495 64.520 ;
        RECT 10.725 64.375 10.935 65.195 ;
        RECT 11.105 64.395 11.435 65.025 ;
        RECT 11.105 63.795 11.355 64.395 ;
        RECT 11.605 64.375 11.835 65.195 ;
        RECT 12.210 64.685 12.450 65.195 ;
        RECT 12.630 64.685 12.910 65.015 ;
        RECT 13.140 64.685 13.355 65.195 ;
        RECT 11.525 63.955 11.855 64.205 ;
        RECT 12.105 63.955 12.460 64.515 ;
        RECT 9.365 62.815 9.545 63.575 ;
        RECT 9.725 62.645 10.055 63.405 ;
        RECT 10.225 62.815 10.495 63.720 ;
        RECT 10.725 62.645 10.935 63.785 ;
        RECT 11.105 62.815 11.435 63.795 ;
        RECT 12.630 63.785 12.800 64.685 ;
        RECT 12.970 63.955 13.235 64.515 ;
        RECT 13.525 64.455 14.140 65.025 ;
        RECT 13.485 63.785 13.655 64.285 ;
        RECT 11.605 62.645 11.835 63.785 ;
        RECT 12.230 63.615 13.655 63.785 ;
        RECT 12.230 63.440 12.620 63.615 ;
        RECT 13.105 62.645 13.435 63.445 ;
        RECT 13.825 63.435 14.140 64.455 ;
        RECT 15.325 64.375 15.535 65.195 ;
        RECT 15.705 64.395 16.035 65.025 ;
        RECT 15.705 63.795 15.955 64.395 ;
        RECT 16.205 64.375 16.435 65.195 ;
        RECT 16.125 63.955 16.455 64.205 ;
        RECT 13.605 62.815 14.140 63.435 ;
        RECT 15.325 62.645 15.535 63.785 ;
        RECT 15.705 62.815 16.035 63.795 ;
        RECT 16.205 62.645 16.435 63.785 ;
        RECT 16.645 62.815 17.395 65.025 ;
        RECT 17.655 64.645 17.825 65.025 ;
        RECT 18.005 64.815 18.335 65.195 ;
        RECT 17.655 64.475 18.320 64.645 ;
        RECT 18.515 64.520 18.775 65.025 ;
        RECT 17.585 63.925 17.925 64.295 ;
        RECT 18.150 64.220 18.320 64.475 ;
        RECT 18.150 63.890 18.425 64.220 ;
        RECT 18.150 63.745 18.320 63.890 ;
        RECT 17.645 63.575 18.320 63.745 ;
        RECT 18.595 63.720 18.775 64.520 ;
        RECT 18.955 64.465 19.255 65.195 ;
        RECT 19.435 64.285 19.665 64.905 ;
        RECT 19.865 64.635 20.090 65.015 ;
        RECT 20.260 64.805 20.590 65.195 ;
        RECT 19.865 64.455 20.195 64.635 ;
        RECT 18.960 63.955 19.255 64.285 ;
        RECT 19.435 63.955 19.850 64.285 ;
        RECT 20.020 63.785 20.195 64.455 ;
        RECT 20.365 63.955 20.605 64.605 ;
        RECT 17.645 62.815 17.825 63.575 ;
        RECT 18.005 62.645 18.335 63.405 ;
        RECT 18.505 62.815 18.775 63.720 ;
        RECT 18.955 63.425 19.850 63.755 ;
        RECT 20.020 63.595 20.605 63.785 ;
        RECT 18.955 63.255 20.160 63.425 ;
        RECT 18.955 62.825 19.285 63.255 ;
        RECT 19.465 62.645 19.660 63.085 ;
        RECT 19.830 62.825 20.160 63.255 ;
        RECT 20.330 62.825 20.605 63.595 ;
        RECT 20.785 62.815 21.535 65.025 ;
        RECT 21.795 64.645 21.965 65.025 ;
        RECT 22.145 64.815 22.475 65.195 ;
        RECT 21.795 64.475 22.460 64.645 ;
        RECT 22.655 64.520 22.915 65.025 ;
        RECT 21.725 63.925 22.065 64.295 ;
        RECT 22.290 64.220 22.460 64.475 ;
        RECT 22.290 63.890 22.565 64.220 ;
        RECT 22.290 63.745 22.460 63.890 ;
        RECT 21.785 63.575 22.460 63.745 ;
        RECT 22.735 63.720 22.915 64.520 ;
        RECT 21.785 62.815 21.965 63.575 ;
        RECT 22.145 62.645 22.475 63.405 ;
        RECT 22.645 62.815 22.915 63.720 ;
        RECT 23.085 64.520 23.345 65.025 ;
        RECT 23.525 64.815 23.855 65.195 ;
        RECT 24.035 64.645 24.205 65.025 ;
        RECT 23.085 63.720 23.255 64.520 ;
        RECT 23.540 64.475 24.205 64.645 ;
        RECT 24.555 64.645 24.725 65.025 ;
        RECT 24.905 64.815 25.235 65.195 ;
        RECT 24.555 64.475 25.220 64.645 ;
        RECT 25.415 64.520 25.675 65.025 ;
        RECT 23.540 64.220 23.710 64.475 ;
        RECT 23.425 63.890 23.710 64.220 ;
        RECT 23.945 63.925 24.275 64.295 ;
        RECT 24.485 63.925 24.825 64.295 ;
        RECT 25.050 64.220 25.220 64.475 ;
        RECT 23.540 63.745 23.710 63.890 ;
        RECT 25.050 63.890 25.325 64.220 ;
        RECT 25.050 63.745 25.220 63.890 ;
        RECT 23.085 62.815 23.355 63.720 ;
        RECT 23.540 63.575 24.205 63.745 ;
        RECT 23.525 62.645 23.855 63.405 ;
        RECT 24.035 62.815 24.205 63.575 ;
        RECT 24.545 63.575 25.220 63.745 ;
        RECT 25.495 63.720 25.675 64.520 ;
        RECT 24.545 62.815 24.725 63.575 ;
        RECT 24.905 62.645 25.235 63.405 ;
        RECT 25.405 62.815 25.675 63.720 ;
        RECT 25.855 62.825 26.115 65.015 ;
        RECT 26.375 64.825 27.045 65.195 ;
        RECT 27.225 64.645 27.535 65.015 ;
        RECT 26.305 64.445 27.535 64.645 ;
        RECT 26.305 63.775 26.595 64.445 ;
        RECT 27.715 64.265 27.945 64.905 ;
        RECT 28.125 64.465 28.415 65.195 ;
        RECT 28.610 64.690 28.945 65.195 ;
        RECT 29.115 64.625 29.355 65.000 ;
        RECT 29.635 64.865 29.805 65.010 ;
        RECT 29.635 64.670 30.010 64.865 ;
        RECT 30.370 64.700 30.765 65.195 ;
        RECT 26.775 63.955 27.240 64.265 ;
        RECT 27.420 63.955 27.945 64.265 ;
        RECT 28.125 63.955 28.425 64.285 ;
        RECT 26.305 63.555 27.075 63.775 ;
        RECT 26.285 62.645 26.625 63.375 ;
        RECT 26.805 62.825 27.075 63.555 ;
        RECT 27.255 63.535 28.415 63.775 ;
        RECT 28.665 63.665 28.965 64.515 ;
        RECT 29.135 64.475 29.355 64.625 ;
        RECT 29.135 64.145 29.670 64.475 ;
        RECT 29.840 64.335 30.010 64.670 ;
        RECT 30.935 64.505 31.175 65.025 ;
        RECT 27.255 62.825 27.485 63.535 ;
        RECT 27.655 62.645 27.985 63.355 ;
        RECT 28.155 62.825 28.415 63.535 ;
        RECT 29.135 63.495 29.370 64.145 ;
        RECT 29.840 63.975 30.825 64.335 ;
        RECT 28.695 63.265 29.370 63.495 ;
        RECT 29.540 63.955 30.825 63.975 ;
        RECT 29.540 63.805 30.400 63.955 ;
        RECT 28.695 62.835 28.865 63.265 ;
        RECT 29.035 62.645 29.365 63.095 ;
        RECT 29.540 62.860 29.825 63.805 ;
        RECT 31.000 63.700 31.175 64.505 ;
        RECT 31.365 64.470 31.655 65.195 ;
        RECT 32.290 64.430 32.745 65.195 ;
        RECT 33.020 64.815 34.320 65.025 ;
        RECT 34.575 64.835 34.905 65.195 ;
        RECT 34.150 64.665 34.320 64.815 ;
        RECT 35.075 64.695 35.335 65.025 ;
        RECT 33.220 64.205 33.440 64.605 ;
        RECT 32.285 64.005 32.775 64.205 ;
        RECT 32.965 63.995 33.440 64.205 ;
        RECT 33.685 64.205 33.895 64.605 ;
        RECT 34.150 64.540 34.905 64.665 ;
        RECT 34.150 64.495 34.995 64.540 ;
        RECT 34.725 64.375 34.995 64.495 ;
        RECT 33.685 63.995 34.015 64.205 ;
        RECT 34.185 63.935 34.595 64.240 ;
        RECT 30.000 63.325 30.695 63.635 ;
        RECT 30.005 62.645 30.690 63.115 ;
        RECT 30.870 62.915 31.175 63.700 ;
        RECT 31.365 62.645 31.655 63.810 ;
        RECT 32.290 63.765 33.465 63.825 ;
        RECT 34.825 63.800 34.995 64.375 ;
        RECT 34.795 63.765 34.995 63.800 ;
        RECT 32.290 63.655 34.995 63.765 ;
        RECT 32.290 63.035 32.545 63.655 ;
        RECT 33.135 63.595 34.935 63.655 ;
        RECT 33.135 63.565 33.465 63.595 ;
        RECT 35.165 63.495 35.335 64.695 ;
        RECT 32.795 63.395 32.980 63.485 ;
        RECT 33.570 63.395 34.405 63.405 ;
        RECT 32.795 63.195 34.405 63.395 ;
        RECT 32.795 63.155 33.025 63.195 ;
        RECT 32.290 62.815 32.625 63.035 ;
        RECT 33.630 62.645 33.985 63.025 ;
        RECT 34.155 62.815 34.405 63.195 ;
        RECT 34.655 62.645 34.905 63.425 ;
        RECT 35.075 62.815 35.335 63.495 ;
        RECT 35.505 64.695 35.765 65.025 ;
        RECT 35.935 64.835 36.265 65.195 ;
        RECT 36.520 64.815 37.820 65.025 ;
        RECT 35.505 64.685 35.735 64.695 ;
        RECT 35.505 63.495 35.675 64.685 ;
        RECT 36.520 64.665 36.690 64.815 ;
        RECT 35.935 64.540 36.690 64.665 ;
        RECT 35.845 64.495 36.690 64.540 ;
        RECT 35.845 64.375 36.115 64.495 ;
        RECT 35.845 63.800 36.015 64.375 ;
        RECT 36.245 63.935 36.655 64.240 ;
        RECT 36.945 64.205 37.155 64.605 ;
        RECT 36.825 63.995 37.155 64.205 ;
        RECT 37.400 64.205 37.620 64.605 ;
        RECT 38.095 64.430 38.550 65.195 ;
        RECT 38.815 64.715 39.115 65.195 ;
        RECT 39.285 64.545 39.545 65.000 ;
        RECT 39.715 64.715 39.975 65.195 ;
        RECT 40.155 64.545 40.415 65.000 ;
        RECT 40.585 64.715 40.835 65.195 ;
        RECT 41.015 64.545 41.275 65.000 ;
        RECT 41.445 64.715 41.695 65.195 ;
        RECT 41.875 64.545 42.135 65.000 ;
        RECT 42.305 64.715 42.550 65.195 ;
        RECT 42.720 64.545 42.995 65.000 ;
        RECT 43.165 64.715 43.410 65.195 ;
        RECT 43.580 64.545 43.840 65.000 ;
        RECT 44.010 64.715 44.270 65.195 ;
        RECT 44.440 64.545 44.700 65.000 ;
        RECT 44.870 64.715 45.130 65.195 ;
        RECT 45.300 64.545 45.560 65.000 ;
        RECT 45.730 64.635 45.990 65.195 ;
        RECT 38.815 64.375 45.560 64.545 ;
        RECT 37.400 63.995 37.875 64.205 ;
        RECT 38.065 64.005 38.555 64.205 ;
        RECT 35.845 63.765 36.045 63.800 ;
        RECT 37.375 63.765 38.550 63.825 ;
        RECT 35.845 63.655 38.550 63.765 ;
        RECT 35.905 63.595 37.705 63.655 ;
        RECT 37.375 63.565 37.705 63.595 ;
        RECT 35.505 62.815 35.765 63.495 ;
        RECT 35.935 62.645 36.185 63.425 ;
        RECT 36.435 63.395 37.270 63.405 ;
        RECT 37.860 63.395 38.045 63.485 ;
        RECT 36.435 63.195 38.045 63.395 ;
        RECT 36.435 62.815 36.685 63.195 ;
        RECT 37.815 63.155 38.045 63.195 ;
        RECT 38.295 63.035 38.550 63.655 ;
        RECT 38.815 63.785 39.980 64.375 ;
        RECT 46.160 64.205 46.410 65.015 ;
        RECT 46.590 64.670 46.850 65.195 ;
        RECT 47.020 64.205 47.270 65.015 ;
        RECT 47.450 64.685 47.755 65.195 ;
        RECT 48.015 64.715 48.315 65.195 ;
        RECT 48.485 64.545 48.745 65.000 ;
        RECT 48.915 64.715 49.175 65.195 ;
        RECT 49.355 64.545 49.615 65.000 ;
        RECT 49.785 64.715 50.035 65.195 ;
        RECT 50.215 64.545 50.475 65.000 ;
        RECT 50.645 64.715 50.895 65.195 ;
        RECT 51.075 64.545 51.335 65.000 ;
        RECT 51.505 64.715 51.750 65.195 ;
        RECT 51.920 64.545 52.195 65.000 ;
        RECT 52.365 64.715 52.610 65.195 ;
        RECT 52.780 64.545 53.040 65.000 ;
        RECT 53.210 64.715 53.470 65.195 ;
        RECT 53.640 64.545 53.900 65.000 ;
        RECT 54.070 64.715 54.330 65.195 ;
        RECT 54.500 64.545 54.760 65.000 ;
        RECT 54.930 64.635 55.190 65.195 ;
        RECT 40.150 63.955 47.270 64.205 ;
        RECT 47.440 63.955 47.755 64.515 ;
        RECT 48.015 64.375 54.760 64.545 ;
        RECT 38.815 63.560 45.560 63.785 ;
        RECT 36.855 62.645 37.210 63.025 ;
        RECT 38.215 62.815 38.550 63.035 ;
        RECT 38.815 62.645 39.085 63.390 ;
        RECT 39.255 62.820 39.545 63.560 ;
        RECT 40.155 63.545 45.560 63.560 ;
        RECT 39.715 62.650 39.970 63.375 ;
        RECT 40.155 62.820 40.415 63.545 ;
        RECT 40.585 62.650 40.830 63.375 ;
        RECT 41.015 62.820 41.275 63.545 ;
        RECT 41.445 62.650 41.690 63.375 ;
        RECT 41.875 62.820 42.135 63.545 ;
        RECT 42.305 62.650 42.550 63.375 ;
        RECT 42.720 62.820 42.980 63.545 ;
        RECT 43.150 62.650 43.410 63.375 ;
        RECT 43.580 62.820 43.840 63.545 ;
        RECT 44.010 62.650 44.270 63.375 ;
        RECT 44.440 62.820 44.700 63.545 ;
        RECT 44.870 62.650 45.130 63.375 ;
        RECT 45.300 62.820 45.560 63.545 ;
        RECT 45.730 62.650 45.990 63.445 ;
        RECT 46.160 62.820 46.410 63.955 ;
        RECT 39.715 62.645 45.990 62.650 ;
        RECT 46.590 62.645 46.850 63.455 ;
        RECT 47.025 62.815 47.270 63.955 ;
        RECT 48.015 63.785 49.180 64.375 ;
        RECT 55.360 64.205 55.610 65.015 ;
        RECT 55.790 64.670 56.050 65.195 ;
        RECT 56.220 64.205 56.470 65.015 ;
        RECT 56.650 64.685 56.955 65.195 ;
        RECT 49.350 63.955 56.470 64.205 ;
        RECT 56.640 63.955 56.955 64.515 ;
        RECT 57.125 64.470 57.415 65.195 ;
        RECT 57.590 64.375 57.885 65.195 ;
        RECT 58.055 64.645 58.275 65.025 ;
        RECT 58.445 64.835 59.295 65.195 ;
        RECT 48.015 63.560 54.760 63.785 ;
        RECT 47.450 62.645 47.745 63.455 ;
        RECT 48.015 62.645 48.285 63.390 ;
        RECT 48.455 62.820 48.745 63.560 ;
        RECT 49.355 63.545 54.760 63.560 ;
        RECT 48.915 62.650 49.170 63.375 ;
        RECT 49.355 62.820 49.615 63.545 ;
        RECT 49.785 62.650 50.030 63.375 ;
        RECT 50.215 62.820 50.475 63.545 ;
        RECT 50.645 62.650 50.890 63.375 ;
        RECT 51.075 62.820 51.335 63.545 ;
        RECT 51.505 62.650 51.750 63.375 ;
        RECT 51.920 62.820 52.180 63.545 ;
        RECT 52.350 62.650 52.610 63.375 ;
        RECT 52.780 62.820 53.040 63.545 ;
        RECT 53.210 62.650 53.470 63.375 ;
        RECT 53.640 62.820 53.900 63.545 ;
        RECT 54.070 62.650 54.330 63.375 ;
        RECT 54.500 62.820 54.760 63.545 ;
        RECT 54.930 62.650 55.190 63.445 ;
        RECT 55.360 62.820 55.610 63.955 ;
        RECT 48.915 62.645 55.190 62.650 ;
        RECT 55.790 62.645 56.050 63.455 ;
        RECT 56.225 62.815 56.470 63.955 ;
        RECT 56.650 62.645 56.945 63.455 ;
        RECT 57.125 62.645 57.415 63.810 ;
        RECT 57.590 62.645 57.885 63.790 ;
        RECT 58.055 62.945 58.285 64.645 ;
        RECT 59.775 64.585 60.105 65.005 ;
        RECT 60.310 64.755 60.585 65.195 ;
        RECT 60.755 64.585 61.085 65.005 ;
        RECT 58.500 64.405 61.085 64.585 ;
        RECT 58.500 63.790 58.810 64.405 ;
        RECT 61.265 64.395 61.525 65.195 ;
        RECT 58.980 64.005 59.310 64.235 ;
        RECT 59.480 64.005 59.950 64.235 ;
        RECT 60.120 64.175 60.570 64.235 ;
        RECT 60.120 64.005 60.575 64.175 ;
        RECT 60.760 64.005 61.095 64.235 ;
        RECT 58.500 63.620 61.085 63.790 ;
        RECT 58.500 62.645 58.755 63.450 ;
        RECT 58.955 63.260 60.295 63.440 ;
        RECT 58.955 62.815 59.285 63.260 ;
        RECT 59.455 62.645 59.730 63.090 ;
        RECT 59.965 62.815 60.295 63.260 ;
        RECT 60.755 62.955 61.085 63.620 ;
        RECT 61.265 62.645 61.525 63.785 ;
        RECT 61.695 62.815 62.025 65.025 ;
        RECT 62.275 64.455 62.605 65.195 ;
        RECT 62.875 64.625 63.205 65.025 ;
        RECT 63.375 64.795 63.705 65.195 ;
        RECT 63.875 64.855 65.235 65.025 ;
        RECT 63.875 64.625 64.205 64.855 ;
        RECT 62.875 64.455 64.205 64.625 ;
        RECT 64.375 64.455 64.705 64.685 ;
        RECT 62.195 63.495 62.505 64.285 ;
        RECT 62.675 63.665 62.895 64.285 ;
        RECT 63.165 63.665 63.340 64.285 ;
        RECT 63.595 63.665 63.815 64.285 ;
        RECT 64.090 64.175 64.335 64.285 ;
        RECT 64.085 64.005 64.335 64.175 ;
        RECT 64.090 63.665 64.335 64.005 ;
        RECT 64.505 63.495 64.705 64.455 ;
        RECT 64.875 64.375 65.235 64.855 ;
        RECT 66.325 64.685 66.630 65.195 ;
        RECT 64.875 64.035 65.235 64.205 ;
        RECT 64.905 63.955 65.235 64.035 ;
        RECT 66.325 63.955 66.640 64.515 ;
        RECT 66.810 64.205 67.060 65.015 ;
        RECT 67.230 64.670 67.490 65.195 ;
        RECT 67.670 64.205 67.920 65.015 ;
        RECT 68.090 64.635 68.350 65.195 ;
        RECT 68.520 64.545 68.780 65.000 ;
        RECT 68.950 64.715 69.210 65.195 ;
        RECT 69.380 64.545 69.640 65.000 ;
        RECT 69.810 64.715 70.070 65.195 ;
        RECT 70.240 64.545 70.500 65.000 ;
        RECT 70.670 64.715 70.915 65.195 ;
        RECT 71.085 64.545 71.360 65.000 ;
        RECT 71.530 64.715 71.775 65.195 ;
        RECT 71.945 64.545 72.205 65.000 ;
        RECT 72.385 64.715 72.635 65.195 ;
        RECT 72.805 64.545 73.065 65.000 ;
        RECT 73.245 64.715 73.495 65.195 ;
        RECT 73.665 64.545 73.925 65.000 ;
        RECT 74.105 64.715 74.365 65.195 ;
        RECT 74.535 64.545 74.795 65.000 ;
        RECT 74.965 64.715 75.265 65.195 ;
        RECT 68.520 64.375 75.265 64.545 ;
        RECT 75.525 64.445 76.735 65.195 ;
        RECT 66.810 63.955 73.930 64.205 ;
        RECT 62.195 63.325 64.705 63.495 ;
        RECT 62.195 62.645 62.705 63.155 ;
        RECT 63.875 62.815 64.205 63.325 ;
        RECT 64.875 62.645 65.235 63.785 ;
        RECT 66.335 62.645 66.630 63.455 ;
        RECT 66.810 62.815 67.055 63.955 ;
        RECT 67.230 62.645 67.490 63.455 ;
        RECT 67.670 62.820 67.920 63.955 ;
        RECT 74.100 63.785 75.265 64.375 ;
        RECT 68.520 63.560 75.265 63.785 ;
        RECT 75.525 63.735 76.045 64.275 ;
        RECT 76.215 63.905 76.735 64.445 ;
        RECT 68.520 63.545 73.925 63.560 ;
        RECT 68.090 62.650 68.350 63.445 ;
        RECT 68.520 62.820 68.780 63.545 ;
        RECT 68.950 62.650 69.210 63.375 ;
        RECT 69.380 62.820 69.640 63.545 ;
        RECT 69.810 62.650 70.070 63.375 ;
        RECT 70.240 62.820 70.500 63.545 ;
        RECT 70.670 62.650 70.930 63.375 ;
        RECT 71.100 62.820 71.360 63.545 ;
        RECT 71.530 62.650 71.775 63.375 ;
        RECT 71.945 62.820 72.205 63.545 ;
        RECT 72.390 62.650 72.635 63.375 ;
        RECT 72.805 62.820 73.065 63.545 ;
        RECT 73.250 62.650 73.495 63.375 ;
        RECT 73.665 62.820 73.925 63.545 ;
        RECT 74.110 62.650 74.365 63.375 ;
        RECT 74.535 62.820 74.825 63.560 ;
        RECT 68.090 62.645 74.365 62.650 ;
        RECT 74.995 62.645 75.265 63.390 ;
        RECT 75.525 62.645 76.735 63.735 ;
        RECT 5.520 62.475 76.820 62.645 ;
        RECT 5.605 61.385 6.815 62.475 ;
        RECT 5.605 60.675 6.125 61.215 ;
        RECT 6.295 60.845 6.815 61.385 ;
        RECT 7.905 61.400 8.175 62.305 ;
        RECT 8.345 61.715 8.675 62.475 ;
        RECT 8.855 61.545 9.025 62.305 ;
        RECT 5.605 59.925 6.815 60.675 ;
        RECT 7.905 60.600 8.075 61.400 ;
        RECT 8.360 61.375 9.025 61.545 ;
        RECT 9.285 61.400 9.555 62.305 ;
        RECT 9.725 61.715 10.055 62.475 ;
        RECT 10.235 61.545 10.405 62.305 ;
        RECT 8.360 61.230 8.530 61.375 ;
        RECT 8.245 60.900 8.530 61.230 ;
        RECT 8.360 60.645 8.530 60.900 ;
        RECT 8.765 60.825 9.095 61.195 ;
        RECT 7.905 60.095 8.165 60.600 ;
        RECT 8.360 60.475 9.025 60.645 ;
        RECT 8.345 59.925 8.675 60.305 ;
        RECT 8.855 60.095 9.025 60.475 ;
        RECT 9.285 60.600 9.455 61.400 ;
        RECT 9.740 61.375 10.405 61.545 ;
        RECT 10.665 61.400 10.935 62.305 ;
        RECT 11.105 61.715 11.435 62.475 ;
        RECT 11.615 61.545 11.785 62.305 ;
        RECT 9.740 61.230 9.910 61.375 ;
        RECT 9.625 60.900 9.910 61.230 ;
        RECT 9.740 60.645 9.910 60.900 ;
        RECT 10.145 60.825 10.475 61.195 ;
        RECT 9.285 60.095 9.545 60.600 ;
        RECT 9.740 60.475 10.405 60.645 ;
        RECT 9.725 59.925 10.055 60.305 ;
        RECT 10.235 60.095 10.405 60.475 ;
        RECT 10.665 60.600 10.835 61.400 ;
        RECT 11.120 61.375 11.785 61.545 ;
        RECT 12.045 61.400 12.315 62.305 ;
        RECT 12.485 61.715 12.815 62.475 ;
        RECT 12.995 61.545 13.165 62.305 ;
        RECT 11.120 61.230 11.290 61.375 ;
        RECT 11.005 60.900 11.290 61.230 ;
        RECT 11.120 60.645 11.290 60.900 ;
        RECT 11.525 60.825 11.855 61.195 ;
        RECT 10.665 60.095 10.925 60.600 ;
        RECT 11.120 60.475 11.785 60.645 ;
        RECT 11.105 59.925 11.435 60.305 ;
        RECT 11.615 60.095 11.785 60.475 ;
        RECT 12.045 60.600 12.215 61.400 ;
        RECT 12.500 61.375 13.165 61.545 ;
        RECT 13.610 61.505 14.000 61.680 ;
        RECT 14.485 61.675 14.815 62.475 ;
        RECT 14.985 61.685 15.520 62.305 ;
        RECT 12.500 61.230 12.670 61.375 ;
        RECT 13.610 61.335 15.035 61.505 ;
        RECT 12.385 60.900 12.670 61.230 ;
        RECT 12.500 60.645 12.670 60.900 ;
        RECT 12.905 60.825 13.235 61.195 ;
        RECT 12.045 60.095 12.305 60.600 ;
        RECT 12.500 60.475 13.165 60.645 ;
        RECT 13.485 60.605 13.840 61.165 ;
        RECT 12.485 59.925 12.815 60.305 ;
        RECT 12.995 60.095 13.165 60.475 ;
        RECT 14.010 60.435 14.180 61.335 ;
        RECT 14.350 60.605 14.615 61.165 ;
        RECT 14.865 60.835 15.035 61.335 ;
        RECT 15.205 60.665 15.520 61.685 ;
        RECT 15.730 61.325 15.990 62.475 ;
        RECT 16.165 61.400 16.420 62.305 ;
        RECT 16.590 61.715 16.920 62.475 ;
        RECT 17.135 61.545 17.305 62.305 ;
        RECT 13.590 59.925 13.830 60.435 ;
        RECT 14.010 60.105 14.290 60.435 ;
        RECT 14.520 59.925 14.735 60.435 ;
        RECT 14.905 60.095 15.520 60.665 ;
        RECT 15.730 59.925 15.990 60.765 ;
        RECT 16.165 60.670 16.335 61.400 ;
        RECT 16.590 61.375 17.305 61.545 ;
        RECT 16.590 61.165 16.760 61.375 ;
        RECT 18.485 61.310 18.775 62.475 ;
        RECT 19.870 61.335 20.205 62.305 ;
        RECT 20.375 61.335 20.545 62.475 ;
        RECT 20.715 62.135 22.745 62.305 ;
        RECT 16.505 60.835 16.760 61.165 ;
        RECT 16.165 60.095 16.420 60.670 ;
        RECT 16.590 60.645 16.760 60.835 ;
        RECT 17.040 60.825 17.395 61.195 ;
        RECT 19.870 60.665 20.040 61.335 ;
        RECT 20.715 61.165 20.885 62.135 ;
        RECT 20.210 60.835 20.465 61.165 ;
        RECT 20.690 60.835 20.885 61.165 ;
        RECT 21.055 61.795 22.180 61.965 ;
        RECT 20.295 60.665 20.465 60.835 ;
        RECT 21.055 60.665 21.225 61.795 ;
        RECT 16.590 60.475 17.305 60.645 ;
        RECT 16.590 59.925 16.920 60.305 ;
        RECT 17.135 60.095 17.305 60.475 ;
        RECT 18.485 59.925 18.775 60.650 ;
        RECT 19.870 60.095 20.125 60.665 ;
        RECT 20.295 60.495 21.225 60.665 ;
        RECT 21.395 61.455 22.405 61.625 ;
        RECT 21.395 60.655 21.565 61.455 ;
        RECT 21.050 60.460 21.225 60.495 ;
        RECT 20.295 59.925 20.625 60.325 ;
        RECT 21.050 60.095 21.580 60.460 ;
        RECT 21.770 60.435 22.045 61.255 ;
        RECT 21.765 60.265 22.045 60.435 ;
        RECT 21.770 60.095 22.045 60.265 ;
        RECT 22.215 60.095 22.405 61.455 ;
        RECT 22.575 61.470 22.745 62.135 ;
        RECT 22.915 61.715 23.085 62.475 ;
        RECT 23.320 61.715 23.835 62.125 ;
        RECT 22.575 61.280 23.325 61.470 ;
        RECT 23.495 60.905 23.835 61.715 ;
        RECT 25.015 61.545 25.185 62.305 ;
        RECT 25.365 61.715 25.695 62.475 ;
        RECT 25.015 61.375 25.680 61.545 ;
        RECT 25.865 61.400 26.135 62.305 ;
        RECT 25.510 61.230 25.680 61.375 ;
        RECT 22.605 60.735 23.835 60.905 ;
        RECT 24.945 60.825 25.275 61.195 ;
        RECT 25.510 60.900 25.795 61.230 ;
        RECT 22.585 59.925 23.095 60.460 ;
        RECT 23.315 60.130 23.560 60.735 ;
        RECT 25.510 60.645 25.680 60.900 ;
        RECT 25.015 60.475 25.680 60.645 ;
        RECT 25.965 60.600 26.135 61.400 ;
        RECT 25.015 60.095 25.185 60.475 ;
        RECT 25.365 59.925 25.695 60.305 ;
        RECT 25.875 60.095 26.135 60.600 ;
        RECT 26.305 61.755 26.765 62.305 ;
        RECT 26.955 61.755 27.285 62.475 ;
        RECT 26.305 60.385 26.555 61.755 ;
        RECT 27.485 61.585 27.785 62.135 ;
        RECT 27.955 61.805 28.235 62.475 ;
        RECT 26.845 61.415 27.785 61.585 ;
        RECT 26.845 61.165 27.015 61.415 ;
        RECT 28.155 61.165 28.420 61.525 ;
        RECT 28.605 61.335 28.865 62.475 ;
        RECT 29.035 61.325 29.365 62.305 ;
        RECT 29.535 61.335 29.815 62.475 ;
        RECT 30.000 61.490 30.325 62.475 ;
        RECT 30.895 61.845 31.155 62.305 ;
        RECT 31.325 62.025 32.175 62.475 ;
        RECT 30.510 61.455 30.715 61.825 ;
        RECT 30.895 61.625 32.015 61.845 ;
        RECT 26.725 60.835 27.015 61.165 ;
        RECT 27.185 60.915 27.525 61.165 ;
        RECT 27.745 60.915 28.420 61.165 ;
        RECT 28.625 60.915 28.960 61.165 ;
        RECT 26.845 60.745 27.015 60.835 ;
        RECT 26.845 60.555 28.235 60.745 ;
        RECT 29.130 60.725 29.300 61.325 ;
        RECT 29.470 60.895 29.805 61.165 ;
        RECT 29.995 60.835 30.255 61.290 ;
        RECT 30.505 61.285 30.715 61.455 ;
        RECT 30.510 61.240 30.715 61.285 ;
        RECT 30.510 60.865 31.095 61.240 ;
        RECT 31.265 60.850 31.675 61.455 ;
        RECT 31.845 61.170 32.015 61.625 ;
        RECT 26.305 60.095 26.865 60.385 ;
        RECT 27.035 59.925 27.285 60.385 ;
        RECT 27.905 60.195 28.235 60.555 ;
        RECT 28.605 60.095 29.300 60.725 ;
        RECT 29.505 59.925 29.815 60.725 ;
        RECT 31.845 60.680 32.175 61.170 ;
        RECT 30.000 60.475 31.155 60.665 ;
        RECT 30.000 60.335 30.275 60.475 ;
        RECT 30.945 60.305 31.155 60.475 ;
        RECT 31.325 60.475 32.175 60.680 ;
        RECT 30.445 59.925 30.775 60.305 ;
        RECT 31.325 60.095 31.655 60.475 ;
        RECT 31.845 59.925 32.175 60.305 ;
        RECT 32.345 60.095 32.590 62.305 ;
        RECT 32.775 61.475 33.030 62.475 ;
        RECT 33.205 61.335 33.465 62.475 ;
        RECT 33.635 61.325 33.965 62.305 ;
        RECT 34.135 61.335 34.415 62.475 ;
        RECT 35.135 61.730 35.405 62.475 ;
        RECT 36.035 62.470 42.310 62.475 ;
        RECT 35.575 61.560 35.865 62.300 ;
        RECT 36.035 61.745 36.290 62.470 ;
        RECT 36.475 61.575 36.735 62.300 ;
        RECT 36.905 61.745 37.150 62.470 ;
        RECT 37.335 61.575 37.595 62.300 ;
        RECT 37.765 61.745 38.010 62.470 ;
        RECT 38.195 61.575 38.455 62.300 ;
        RECT 38.625 61.745 38.870 62.470 ;
        RECT 39.040 61.575 39.300 62.300 ;
        RECT 39.470 61.745 39.730 62.470 ;
        RECT 39.900 61.575 40.160 62.300 ;
        RECT 40.330 61.745 40.590 62.470 ;
        RECT 40.760 61.575 41.020 62.300 ;
        RECT 41.190 61.745 41.450 62.470 ;
        RECT 41.620 61.575 41.880 62.300 ;
        RECT 42.050 61.675 42.310 62.470 ;
        RECT 36.475 61.560 41.880 61.575 ;
        RECT 35.135 61.455 41.880 61.560 ;
        RECT 35.105 61.335 41.880 61.455 ;
        RECT 33.225 60.915 33.560 61.165 ;
        RECT 33.730 60.725 33.900 61.325 ;
        RECT 35.105 61.285 36.300 61.335 ;
        RECT 34.070 60.895 34.405 61.165 ;
        RECT 35.135 60.745 36.300 61.285 ;
        RECT 42.480 61.165 42.730 62.300 ;
        RECT 42.910 61.665 43.170 62.475 ;
        RECT 43.345 61.165 43.590 62.305 ;
        RECT 43.770 61.665 44.065 62.475 ;
        RECT 44.245 61.310 44.535 62.475 ;
        RECT 44.810 61.675 45.065 62.475 ;
        RECT 45.235 61.505 45.565 62.305 ;
        RECT 45.735 61.675 45.905 62.475 ;
        RECT 46.075 61.505 46.405 62.305 ;
        RECT 44.705 61.335 46.405 61.505 ;
        RECT 46.575 61.335 46.835 62.475 ;
        RECT 47.005 62.055 47.345 62.475 ;
        RECT 47.515 61.885 47.765 62.305 ;
        RECT 47.005 61.715 47.765 61.885 ;
        RECT 36.470 60.915 43.590 61.165 ;
        RECT 32.775 59.925 33.015 60.725 ;
        RECT 33.205 60.095 33.900 60.725 ;
        RECT 34.105 59.925 34.415 60.725 ;
        RECT 35.135 60.575 41.880 60.745 ;
        RECT 35.135 59.925 35.435 60.405 ;
        RECT 35.605 60.120 35.865 60.575 ;
        RECT 36.035 59.925 36.295 60.405 ;
        RECT 36.475 60.120 36.735 60.575 ;
        RECT 36.905 59.925 37.155 60.405 ;
        RECT 37.335 60.120 37.595 60.575 ;
        RECT 37.765 59.925 38.015 60.405 ;
        RECT 38.195 60.120 38.455 60.575 ;
        RECT 38.625 59.925 38.870 60.405 ;
        RECT 39.040 60.120 39.315 60.575 ;
        RECT 39.485 59.925 39.730 60.405 ;
        RECT 39.900 60.120 40.160 60.575 ;
        RECT 40.330 59.925 40.590 60.405 ;
        RECT 40.760 60.120 41.020 60.575 ;
        RECT 41.190 59.925 41.450 60.405 ;
        RECT 41.620 60.120 41.880 60.575 ;
        RECT 42.050 59.925 42.310 60.485 ;
        RECT 42.480 60.105 42.730 60.915 ;
        RECT 42.910 59.925 43.170 60.450 ;
        RECT 43.340 60.105 43.590 60.915 ;
        RECT 43.760 60.605 44.075 61.165 ;
        RECT 44.705 60.745 44.985 61.335 ;
        RECT 45.155 60.915 45.905 61.165 ;
        RECT 46.075 60.915 46.835 61.165 ;
        RECT 47.005 60.745 47.315 61.715 ;
        RECT 47.935 61.635 48.265 62.475 ;
        RECT 48.755 61.885 49.510 62.305 ;
        RECT 48.435 61.715 49.900 61.885 ;
        RECT 48.435 61.465 48.605 61.715 ;
        RECT 47.645 61.295 48.605 61.465 ;
        RECT 47.645 61.125 47.815 61.295 ;
        RECT 48.775 61.125 49.080 61.545 ;
        RECT 47.485 60.915 47.815 61.125 ;
        RECT 47.985 60.915 48.425 61.125 ;
        RECT 48.595 60.915 49.080 61.125 ;
        RECT 49.270 61.115 49.560 61.545 ;
        RECT 49.730 61.510 49.900 61.715 ;
        RECT 50.070 61.690 50.310 62.475 ;
        RECT 50.480 61.510 50.810 62.305 ;
        RECT 51.235 61.730 51.505 62.475 ;
        RECT 52.135 62.470 58.410 62.475 ;
        RECT 51.675 61.560 51.965 62.300 ;
        RECT 52.135 61.745 52.390 62.470 ;
        RECT 52.575 61.575 52.835 62.300 ;
        RECT 53.005 61.745 53.250 62.470 ;
        RECT 53.435 61.575 53.695 62.300 ;
        RECT 53.865 61.745 54.110 62.470 ;
        RECT 54.295 61.575 54.555 62.300 ;
        RECT 54.725 61.745 54.970 62.470 ;
        RECT 55.140 61.575 55.400 62.300 ;
        RECT 55.570 61.745 55.830 62.470 ;
        RECT 56.000 61.575 56.260 62.300 ;
        RECT 56.430 61.745 56.690 62.470 ;
        RECT 56.860 61.575 57.120 62.300 ;
        RECT 57.290 61.745 57.550 62.470 ;
        RECT 57.720 61.575 57.980 62.300 ;
        RECT 58.150 61.675 58.410 62.470 ;
        RECT 52.575 61.560 57.980 61.575 ;
        RECT 49.730 61.335 50.810 61.510 ;
        RECT 51.235 61.335 57.980 61.560 ;
        RECT 49.730 61.285 50.515 61.335 ;
        RECT 49.270 60.915 49.660 61.115 ;
        RECT 49.830 60.915 50.175 61.115 ;
        RECT 43.770 59.925 44.075 60.435 ;
        RECT 44.245 59.925 44.535 60.650 ;
        RECT 44.705 60.495 45.565 60.745 ;
        RECT 45.735 60.555 46.835 60.725 ;
        RECT 47.005 60.575 47.765 60.745 ;
        RECT 44.815 60.305 45.145 60.325 ;
        RECT 45.735 60.305 45.985 60.555 ;
        RECT 44.815 60.095 45.985 60.305 ;
        RECT 46.155 59.925 46.325 60.385 ;
        RECT 46.495 60.095 46.835 60.555 ;
        RECT 47.095 59.925 47.265 60.405 ;
        RECT 47.435 60.105 47.765 60.575 ;
        RECT 47.935 59.925 48.105 60.745 ;
        RECT 48.275 60.575 49.975 60.745 ;
        RECT 48.275 60.110 48.605 60.575 ;
        RECT 49.590 60.485 49.975 60.575 ;
        RECT 50.345 60.645 50.515 61.285 ;
        RECT 50.715 60.815 50.975 61.165 ;
        RECT 51.235 60.745 52.400 61.335 ;
        RECT 58.580 61.165 58.830 62.300 ;
        RECT 59.010 61.665 59.270 62.475 ;
        RECT 59.445 61.165 59.690 62.305 ;
        RECT 59.870 61.665 60.165 62.475 ;
        RECT 60.435 61.730 60.705 62.475 ;
        RECT 61.335 62.470 67.610 62.475 ;
        RECT 60.875 61.560 61.165 62.300 ;
        RECT 61.335 61.745 61.590 62.470 ;
        RECT 61.775 61.575 62.035 62.300 ;
        RECT 62.205 61.745 62.450 62.470 ;
        RECT 62.635 61.575 62.895 62.300 ;
        RECT 63.065 61.745 63.310 62.470 ;
        RECT 63.495 61.575 63.755 62.300 ;
        RECT 63.925 61.745 64.170 62.470 ;
        RECT 64.340 61.575 64.600 62.300 ;
        RECT 64.770 61.745 65.030 62.470 ;
        RECT 65.200 61.575 65.460 62.300 ;
        RECT 65.630 61.745 65.890 62.470 ;
        RECT 66.060 61.575 66.320 62.300 ;
        RECT 66.490 61.745 66.750 62.470 ;
        RECT 66.920 61.575 67.180 62.300 ;
        RECT 67.350 61.675 67.610 62.470 ;
        RECT 61.775 61.560 67.180 61.575 ;
        RECT 60.435 61.335 67.180 61.560 ;
        RECT 52.570 60.915 59.690 61.165 ;
        RECT 50.345 60.475 50.890 60.645 ;
        RECT 51.235 60.575 57.980 60.745 ;
        RECT 48.775 59.925 48.945 60.395 ;
        RECT 49.205 60.135 50.390 60.305 ;
        RECT 50.560 60.095 50.890 60.475 ;
        RECT 51.235 59.925 51.535 60.405 ;
        RECT 51.705 60.120 51.965 60.575 ;
        RECT 52.135 59.925 52.395 60.405 ;
        RECT 52.575 60.120 52.835 60.575 ;
        RECT 53.005 59.925 53.255 60.405 ;
        RECT 53.435 60.120 53.695 60.575 ;
        RECT 53.865 59.925 54.115 60.405 ;
        RECT 54.295 60.120 54.555 60.575 ;
        RECT 54.725 59.925 54.970 60.405 ;
        RECT 55.140 60.120 55.415 60.575 ;
        RECT 55.585 59.925 55.830 60.405 ;
        RECT 56.000 60.120 56.260 60.575 ;
        RECT 56.430 59.925 56.690 60.405 ;
        RECT 56.860 60.120 57.120 60.575 ;
        RECT 57.290 59.925 57.550 60.405 ;
        RECT 57.720 60.120 57.980 60.575 ;
        RECT 58.150 59.925 58.410 60.485 ;
        RECT 58.580 60.105 58.830 60.915 ;
        RECT 59.010 59.925 59.270 60.450 ;
        RECT 59.440 60.105 59.690 60.915 ;
        RECT 59.860 60.605 60.175 61.165 ;
        RECT 60.435 60.745 61.600 61.335 ;
        RECT 67.780 61.165 68.030 62.300 ;
        RECT 68.210 61.665 68.470 62.475 ;
        RECT 68.645 61.165 68.890 62.305 ;
        RECT 69.070 61.665 69.365 62.475 ;
        RECT 70.005 61.310 70.295 62.475 ;
        RECT 70.525 61.775 70.745 62.305 ;
        RECT 70.915 61.965 71.245 62.475 ;
        RECT 71.415 61.775 71.640 62.305 ;
        RECT 70.525 61.510 71.640 61.775 ;
        RECT 71.810 61.760 72.125 62.305 ;
        RECT 72.315 62.060 72.645 62.475 ;
        RECT 71.810 61.530 72.645 61.760 ;
        RECT 61.770 60.915 68.890 61.165 ;
        RECT 60.435 60.575 67.180 60.745 ;
        RECT 59.870 59.925 60.175 60.435 ;
        RECT 60.435 59.925 60.735 60.405 ;
        RECT 60.905 60.120 61.165 60.575 ;
        RECT 61.335 59.925 61.595 60.405 ;
        RECT 61.775 60.120 62.035 60.575 ;
        RECT 62.205 59.925 62.455 60.405 ;
        RECT 62.635 60.120 62.895 60.575 ;
        RECT 63.065 59.925 63.315 60.405 ;
        RECT 63.495 60.120 63.755 60.575 ;
        RECT 63.925 59.925 64.170 60.405 ;
        RECT 64.340 60.120 64.615 60.575 ;
        RECT 64.785 59.925 65.030 60.405 ;
        RECT 65.200 60.120 65.460 60.575 ;
        RECT 65.630 59.925 65.890 60.405 ;
        RECT 66.060 60.120 66.320 60.575 ;
        RECT 66.490 59.925 66.750 60.405 ;
        RECT 66.920 60.120 67.180 60.575 ;
        RECT 67.350 59.925 67.610 60.485 ;
        RECT 67.780 60.105 68.030 60.915 ;
        RECT 68.210 59.925 68.470 60.450 ;
        RECT 68.640 60.105 68.890 60.915 ;
        RECT 69.060 60.605 69.375 61.165 ;
        RECT 69.070 59.925 69.375 60.435 ;
        RECT 70.005 59.925 70.295 60.650 ;
        RECT 70.475 60.590 70.790 61.165 ;
        RECT 70.465 59.925 70.795 60.405 ;
        RECT 70.980 60.205 71.360 61.165 ;
        RECT 71.810 60.835 72.135 61.250 ;
        RECT 72.305 60.835 72.645 61.530 ;
        RECT 72.305 60.665 72.475 60.835 ;
        RECT 72.815 60.665 73.045 62.305 ;
        RECT 73.215 61.505 73.505 62.475 ;
        RECT 73.690 62.050 74.025 62.475 ;
        RECT 74.195 61.870 74.380 62.275 ;
        RECT 73.715 61.695 74.380 61.870 ;
        RECT 74.585 61.695 74.915 62.475 ;
        RECT 71.735 60.495 72.475 60.665 ;
        RECT 71.735 60.095 71.925 60.495 ;
        RECT 72.645 60.475 73.045 60.665 ;
        RECT 73.715 60.665 74.055 61.695 ;
        RECT 75.085 61.505 75.355 62.275 ;
        RECT 74.225 61.335 75.355 61.505 ;
        RECT 74.225 60.835 74.475 61.335 ;
        RECT 73.715 60.495 74.400 60.665 ;
        RECT 74.655 60.585 75.015 61.165 ;
        RECT 72.145 59.925 72.475 60.285 ;
        RECT 72.645 60.095 72.835 60.475 ;
        RECT 73.005 59.925 73.335 60.305 ;
        RECT 73.690 59.925 74.025 60.325 ;
        RECT 74.195 60.095 74.400 60.495 ;
        RECT 75.185 60.425 75.355 61.335 ;
        RECT 75.525 61.385 76.735 62.475 ;
        RECT 75.525 60.845 76.045 61.385 ;
        RECT 76.215 60.675 76.735 61.215 ;
        RECT 74.610 59.925 74.885 60.405 ;
        RECT 75.095 60.095 75.355 60.425 ;
        RECT 75.525 59.925 76.735 60.675 ;
        RECT 5.520 59.755 76.820 59.925 ;
        RECT 5.605 59.005 6.815 59.755 ;
        RECT 5.605 58.465 6.125 59.005 ;
        RECT 6.990 58.915 7.250 59.755 ;
        RECT 7.425 59.010 7.680 59.585 ;
        RECT 7.850 59.375 8.180 59.755 ;
        RECT 8.395 59.205 8.565 59.585 ;
        RECT 7.850 59.035 8.565 59.205 ;
        RECT 6.295 58.295 6.815 58.835 ;
        RECT 5.605 57.205 6.815 58.295 ;
        RECT 6.990 57.205 7.250 58.355 ;
        RECT 7.425 58.280 7.595 59.010 ;
        RECT 7.850 58.845 8.020 59.035 ;
        RECT 8.825 58.955 9.135 59.755 ;
        RECT 9.340 58.955 10.035 59.585 ;
        RECT 10.205 59.015 10.695 59.585 ;
        RECT 10.865 59.185 11.095 59.585 ;
        RECT 11.265 59.355 11.685 59.755 ;
        RECT 11.855 59.185 12.025 59.585 ;
        RECT 10.865 59.015 12.025 59.185 ;
        RECT 12.195 59.015 12.645 59.755 ;
        RECT 12.815 59.015 13.255 59.575 ;
        RECT 7.765 58.515 8.020 58.845 ;
        RECT 7.850 58.305 8.020 58.515 ;
        RECT 8.300 58.485 8.655 58.855 ;
        RECT 8.835 58.515 9.170 58.785 ;
        RECT 9.340 58.395 9.510 58.955 ;
        RECT 9.680 58.515 10.015 58.765 ;
        RECT 9.340 58.355 9.515 58.395 ;
        RECT 7.425 57.375 7.680 58.280 ;
        RECT 7.850 58.135 8.565 58.305 ;
        RECT 7.850 57.205 8.180 57.965 ;
        RECT 8.395 57.375 8.565 58.135 ;
        RECT 8.825 57.205 9.105 58.345 ;
        RECT 9.275 57.375 9.605 58.355 ;
        RECT 10.205 58.345 10.375 59.015 ;
        RECT 10.545 58.515 10.950 58.845 ;
        RECT 9.775 57.205 10.035 58.345 ;
        RECT 10.205 58.175 10.975 58.345 ;
        RECT 10.215 57.205 10.545 58.005 ;
        RECT 10.725 57.545 10.975 58.175 ;
        RECT 11.165 57.715 11.415 58.845 ;
        RECT 11.615 58.515 11.860 58.845 ;
        RECT 12.045 58.565 12.435 58.845 ;
        RECT 11.615 57.715 11.815 58.515 ;
        RECT 12.605 58.395 12.775 58.845 ;
        RECT 11.985 58.225 12.775 58.395 ;
        RECT 11.985 57.545 12.155 58.225 ;
        RECT 10.725 57.375 12.155 57.545 ;
        RECT 12.325 57.205 12.640 58.055 ;
        RECT 12.945 58.005 13.255 59.015 ;
        RECT 12.815 57.375 13.255 58.005 ;
        RECT 14.345 59.015 14.685 59.585 ;
        RECT 14.880 59.090 15.050 59.755 ;
        RECT 15.330 59.415 15.550 59.460 ;
        RECT 15.325 59.245 15.550 59.415 ;
        RECT 15.720 59.275 16.165 59.445 ;
        RECT 15.330 59.105 15.550 59.245 ;
        RECT 14.345 58.045 14.520 59.015 ;
        RECT 15.330 58.935 15.825 59.105 ;
        RECT 14.690 58.395 14.860 58.845 ;
        RECT 15.030 58.565 15.480 58.765 ;
        RECT 15.650 58.740 15.825 58.935 ;
        RECT 15.995 58.485 16.165 59.275 ;
        RECT 16.335 59.150 16.585 59.520 ;
        RECT 16.415 58.765 16.585 59.150 ;
        RECT 16.755 59.115 17.005 59.520 ;
        RECT 17.175 59.285 17.345 59.755 ;
        RECT 17.515 59.115 17.855 59.520 ;
        RECT 16.755 58.935 17.855 59.115 ;
        RECT 16.415 58.595 16.610 58.765 ;
        RECT 14.690 58.225 15.085 58.395 ;
        RECT 15.995 58.345 16.270 58.485 ;
        RECT 14.345 57.375 14.605 58.045 ;
        RECT 14.915 57.955 15.085 58.225 ;
        RECT 15.255 58.125 16.270 58.345 ;
        RECT 16.440 58.345 16.610 58.595 ;
        RECT 16.780 58.515 17.340 58.765 ;
        RECT 16.440 57.955 16.995 58.345 ;
        RECT 14.915 57.785 16.995 57.955 ;
        RECT 14.775 57.205 15.105 57.605 ;
        RECT 15.975 57.205 16.375 57.605 ;
        RECT 16.665 57.550 16.995 57.785 ;
        RECT 17.165 57.415 17.340 58.515 ;
        RECT 17.510 58.195 17.855 58.765 ;
        RECT 18.025 58.100 18.545 59.585 ;
        RECT 18.715 59.095 19.055 59.755 ;
        RECT 19.425 58.945 19.665 59.755 ;
        RECT 19.835 58.945 20.165 59.585 ;
        RECT 20.335 58.945 20.605 59.755 ;
        RECT 20.790 59.015 21.045 59.585 ;
        RECT 21.215 59.355 21.545 59.755 ;
        RECT 21.970 59.220 22.500 59.585 ;
        RECT 22.690 59.415 22.965 59.585 ;
        RECT 22.685 59.245 22.965 59.415 ;
        RECT 21.970 59.185 22.145 59.220 ;
        RECT 21.215 59.015 22.145 59.185 ;
        RECT 17.510 57.205 17.855 58.025 ;
        RECT 18.215 57.205 18.545 57.930 ;
        RECT 18.715 57.375 19.235 58.925 ;
        RECT 19.405 58.515 19.755 58.765 ;
        RECT 19.925 58.345 20.095 58.945 ;
        RECT 20.265 58.515 20.615 58.765 ;
        RECT 20.790 58.345 20.960 59.015 ;
        RECT 21.215 58.845 21.385 59.015 ;
        RECT 21.130 58.515 21.385 58.845 ;
        RECT 21.610 58.515 21.805 58.845 ;
        RECT 19.415 58.175 20.095 58.345 ;
        RECT 19.415 57.390 19.745 58.175 ;
        RECT 20.275 57.205 20.605 58.345 ;
        RECT 20.790 57.375 21.125 58.345 ;
        RECT 21.295 57.205 21.465 58.345 ;
        RECT 21.635 57.545 21.805 58.515 ;
        RECT 21.975 57.885 22.145 59.015 ;
        RECT 22.315 58.225 22.485 59.025 ;
        RECT 22.690 58.425 22.965 59.245 ;
        RECT 23.135 58.225 23.325 59.585 ;
        RECT 23.505 59.220 24.015 59.755 ;
        RECT 24.235 58.945 24.480 59.550 ;
        RECT 24.930 59.015 25.185 59.585 ;
        RECT 25.355 59.355 25.685 59.755 ;
        RECT 26.110 59.220 26.640 59.585 ;
        RECT 26.830 59.415 27.105 59.585 ;
        RECT 26.825 59.245 27.105 59.415 ;
        RECT 26.110 59.185 26.285 59.220 ;
        RECT 25.355 59.015 26.285 59.185 ;
        RECT 23.525 58.775 24.755 58.945 ;
        RECT 22.315 58.055 23.325 58.225 ;
        RECT 23.495 58.210 24.245 58.400 ;
        RECT 21.975 57.715 23.100 57.885 ;
        RECT 23.495 57.545 23.665 58.210 ;
        RECT 24.415 57.965 24.755 58.775 ;
        RECT 21.635 57.375 23.665 57.545 ;
        RECT 23.835 57.205 24.005 57.965 ;
        RECT 24.240 57.555 24.755 57.965 ;
        RECT 24.930 58.345 25.100 59.015 ;
        RECT 25.355 58.845 25.525 59.015 ;
        RECT 25.270 58.515 25.525 58.845 ;
        RECT 25.750 58.515 25.945 58.845 ;
        RECT 24.930 57.375 25.265 58.345 ;
        RECT 25.435 57.205 25.605 58.345 ;
        RECT 25.775 57.545 25.945 58.515 ;
        RECT 26.115 57.885 26.285 59.015 ;
        RECT 26.455 58.225 26.625 59.025 ;
        RECT 26.830 58.425 27.105 59.245 ;
        RECT 27.275 58.225 27.465 59.585 ;
        RECT 27.645 59.220 28.155 59.755 ;
        RECT 28.375 58.945 28.620 59.550 ;
        RECT 29.985 59.080 30.245 59.585 ;
        RECT 30.425 59.375 30.755 59.755 ;
        RECT 30.935 59.205 31.105 59.585 ;
        RECT 27.665 58.775 28.895 58.945 ;
        RECT 26.455 58.055 27.465 58.225 ;
        RECT 27.635 58.210 28.385 58.400 ;
        RECT 26.115 57.715 27.240 57.885 ;
        RECT 27.635 57.545 27.805 58.210 ;
        RECT 28.555 57.965 28.895 58.775 ;
        RECT 25.775 57.375 27.805 57.545 ;
        RECT 27.975 57.205 28.145 57.965 ;
        RECT 28.380 57.555 28.895 57.965 ;
        RECT 29.985 58.280 30.165 59.080 ;
        RECT 30.440 59.035 31.105 59.205 ;
        RECT 30.440 58.780 30.610 59.035 ;
        RECT 31.365 59.030 31.655 59.755 ;
        RECT 31.875 58.955 32.085 59.755 ;
        RECT 30.335 58.450 30.610 58.780 ;
        RECT 30.835 58.485 31.175 58.855 ;
        RECT 30.440 58.305 30.610 58.450 ;
        RECT 29.985 57.375 30.255 58.280 ;
        RECT 30.440 58.135 31.115 58.305 ;
        RECT 30.425 57.205 30.755 57.965 ;
        RECT 30.935 57.375 31.115 58.135 ;
        RECT 31.365 57.205 31.655 58.370 ;
        RECT 31.875 57.205 32.085 58.345 ;
        RECT 32.255 57.375 32.595 59.585 ;
        RECT 32.775 59.295 33.025 59.755 ;
        RECT 33.215 59.125 33.545 59.585 ;
        RECT 33.745 59.415 34.130 59.585 ;
        RECT 33.725 59.245 34.130 59.415 ;
        RECT 32.770 58.955 33.545 59.125 ;
        RECT 32.770 58.055 33.045 58.955 ;
        RECT 33.245 58.225 33.575 58.765 ;
        RECT 33.745 58.225 34.130 59.245 ;
        RECT 34.605 59.215 34.935 59.585 ;
        RECT 35.125 59.385 35.455 59.755 ;
        RECT 35.625 59.215 35.955 59.585 ;
        RECT 34.605 59.015 35.955 59.215 ;
        RECT 36.425 59.080 36.685 59.585 ;
        RECT 36.865 59.375 37.195 59.755 ;
        RECT 37.375 59.205 37.545 59.585 ;
        RECT 34.420 58.225 34.840 58.765 ;
        RECT 35.040 58.515 35.400 58.845 ;
        RECT 35.570 58.525 36.255 58.835 ;
        RECT 35.110 58.055 35.400 58.515 ;
        RECT 32.770 57.815 34.935 58.055 ;
        RECT 35.105 57.885 35.400 58.055 ;
        RECT 32.775 57.205 33.395 57.645 ;
        RECT 33.600 57.375 33.880 57.815 ;
        RECT 34.065 57.205 34.395 57.585 ;
        RECT 34.605 57.375 34.935 57.815 ;
        RECT 35.110 57.470 35.400 57.885 ;
        RECT 35.625 57.205 35.880 58.345 ;
        RECT 36.050 57.485 36.255 58.525 ;
        RECT 36.425 58.280 36.595 59.080 ;
        RECT 36.880 59.035 37.545 59.205 ;
        RECT 37.890 59.205 38.220 59.585 ;
        RECT 38.390 59.375 39.575 59.545 ;
        RECT 39.835 59.285 40.005 59.755 ;
        RECT 37.890 59.035 38.435 59.205 ;
        RECT 36.880 58.780 37.050 59.035 ;
        RECT 36.765 58.450 37.050 58.780 ;
        RECT 37.285 58.485 37.615 58.855 ;
        RECT 37.805 58.515 38.065 58.865 ;
        RECT 36.880 58.305 37.050 58.450 ;
        RECT 38.265 58.395 38.435 59.035 ;
        RECT 38.805 59.105 39.190 59.195 ;
        RECT 40.175 59.105 40.505 59.570 ;
        RECT 38.805 58.935 40.505 59.105 ;
        RECT 40.675 58.935 40.845 59.755 ;
        RECT 41.015 59.105 41.345 59.575 ;
        RECT 41.515 59.275 41.685 59.755 ;
        RECT 41.955 59.415 43.145 59.585 ;
        RECT 41.955 59.245 42.265 59.415 ;
        RECT 41.015 58.935 41.775 59.105 ;
        RECT 38.605 58.565 38.950 58.765 ;
        RECT 39.120 58.565 39.510 58.765 ;
        RECT 38.265 58.345 39.050 58.395 ;
        RECT 36.425 57.375 36.695 58.280 ;
        RECT 36.880 58.135 37.545 58.305 ;
        RECT 36.865 57.205 37.195 57.965 ;
        RECT 37.375 57.375 37.545 58.135 ;
        RECT 37.970 58.170 39.050 58.345 ;
        RECT 37.970 57.375 38.300 58.170 ;
        RECT 38.470 57.205 38.710 57.990 ;
        RECT 38.880 57.965 39.050 58.170 ;
        RECT 39.220 58.135 39.510 58.565 ;
        RECT 39.700 58.555 40.185 58.765 ;
        RECT 40.355 58.555 40.795 58.765 ;
        RECT 40.965 58.555 41.295 58.765 ;
        RECT 39.700 58.135 40.005 58.555 ;
        RECT 40.965 58.385 41.135 58.555 ;
        RECT 40.175 58.215 41.135 58.385 ;
        RECT 40.175 57.965 40.345 58.215 ;
        RECT 38.880 57.795 40.345 57.965 ;
        RECT 39.270 57.375 40.025 57.795 ;
        RECT 40.515 57.205 40.845 58.045 ;
        RECT 41.465 57.965 41.775 58.935 ;
        RECT 41.950 58.440 42.265 59.075 ;
        RECT 41.015 57.795 41.775 57.965 ;
        RECT 41.015 57.375 41.265 57.795 ;
        RECT 41.435 57.205 41.775 57.625 ;
        RECT 41.955 57.205 42.265 58.270 ;
        RECT 42.435 58.055 42.645 59.245 ;
        RECT 42.815 59.125 43.145 59.415 ;
        RECT 43.385 59.295 43.555 59.755 ;
        RECT 43.785 59.125 44.115 59.585 ;
        RECT 44.295 59.295 44.465 59.755 ;
        RECT 44.645 59.125 44.975 59.585 ;
        RECT 45.225 59.275 45.505 59.755 ;
        RECT 42.815 58.955 44.975 59.125 ;
        RECT 45.675 59.105 45.935 59.495 ;
        RECT 46.110 59.275 46.365 59.755 ;
        RECT 46.535 59.105 46.830 59.495 ;
        RECT 47.010 59.275 47.285 59.755 ;
        RECT 47.455 59.255 47.755 59.585 ;
        RECT 48.015 59.275 48.315 59.755 ;
        RECT 45.180 58.935 46.830 59.105 ;
        RECT 42.985 58.395 43.480 58.765 ;
        RECT 43.660 58.565 44.460 58.765 ;
        RECT 44.630 58.395 44.960 58.785 ;
        RECT 42.925 58.225 44.960 58.395 ;
        RECT 45.180 58.425 45.585 58.935 ;
        RECT 45.755 58.595 46.895 58.765 ;
        RECT 45.180 58.255 45.935 58.425 ;
        RECT 42.435 57.875 44.085 58.055 ;
        RECT 42.435 57.375 42.670 57.875 ;
        RECT 43.785 57.715 44.085 57.875 ;
        RECT 42.840 57.205 43.170 57.665 ;
        RECT 43.365 57.545 43.555 57.705 ;
        RECT 44.255 57.545 44.475 58.055 ;
        RECT 43.365 57.375 44.475 57.545 ;
        RECT 44.645 57.205 44.975 58.055 ;
        RECT 45.220 57.205 45.505 58.075 ;
        RECT 45.675 58.005 45.935 58.255 ;
        RECT 46.725 58.345 46.895 58.595 ;
        RECT 47.065 58.515 47.415 59.085 ;
        RECT 47.585 58.345 47.755 59.255 ;
        RECT 48.485 59.105 48.745 59.560 ;
        RECT 48.915 59.275 49.175 59.755 ;
        RECT 49.355 59.105 49.615 59.560 ;
        RECT 49.785 59.275 50.035 59.755 ;
        RECT 50.215 59.105 50.475 59.560 ;
        RECT 50.645 59.275 50.895 59.755 ;
        RECT 51.075 59.105 51.335 59.560 ;
        RECT 51.505 59.275 51.750 59.755 ;
        RECT 51.920 59.105 52.195 59.560 ;
        RECT 52.365 59.275 52.610 59.755 ;
        RECT 52.780 59.105 53.040 59.560 ;
        RECT 53.210 59.275 53.470 59.755 ;
        RECT 53.640 59.105 53.900 59.560 ;
        RECT 54.070 59.275 54.330 59.755 ;
        RECT 54.500 59.105 54.760 59.560 ;
        RECT 54.930 59.195 55.190 59.755 ;
        RECT 46.725 58.175 47.755 58.345 ;
        RECT 45.675 57.835 46.795 58.005 ;
        RECT 45.675 57.375 45.935 57.835 ;
        RECT 46.110 57.205 46.365 57.665 ;
        RECT 46.535 57.375 46.795 57.835 ;
        RECT 46.965 57.205 47.275 58.005 ;
        RECT 47.445 57.375 47.755 58.175 ;
        RECT 48.015 58.935 54.760 59.105 ;
        RECT 48.015 58.345 49.180 58.935 ;
        RECT 55.360 58.765 55.610 59.575 ;
        RECT 55.790 59.230 56.050 59.755 ;
        RECT 56.220 58.765 56.470 59.575 ;
        RECT 56.650 59.245 56.955 59.755 ;
        RECT 49.350 58.515 56.470 58.765 ;
        RECT 56.640 58.515 56.955 59.075 ;
        RECT 57.125 59.030 57.415 59.755 ;
        RECT 58.115 59.285 58.285 59.755 ;
        RECT 58.455 59.115 58.785 59.565 ;
        RECT 58.955 59.285 59.125 59.755 ;
        RECT 59.295 59.115 59.625 59.565 ;
        RECT 57.950 58.935 59.625 59.115 ;
        RECT 59.795 58.945 59.965 59.755 ;
        RECT 60.135 59.365 61.305 59.535 ;
        RECT 60.135 58.945 60.385 59.365 ;
        RECT 61.475 59.285 61.645 59.755 ;
        RECT 61.915 59.365 63.085 59.585 ;
        RECT 60.555 59.115 60.885 59.195 ;
        RECT 60.555 58.935 61.905 59.115 ;
        RECT 62.335 59.025 62.665 59.195 ;
        RECT 48.015 58.120 54.760 58.345 ;
        RECT 48.015 57.205 48.285 57.950 ;
        RECT 48.455 57.380 48.745 58.120 ;
        RECT 49.355 58.105 54.760 58.120 ;
        RECT 48.915 57.210 49.170 57.935 ;
        RECT 49.355 57.380 49.615 58.105 ;
        RECT 49.785 57.210 50.030 57.935 ;
        RECT 50.215 57.380 50.475 58.105 ;
        RECT 50.645 57.210 50.890 57.935 ;
        RECT 51.075 57.380 51.335 58.105 ;
        RECT 51.505 57.210 51.750 57.935 ;
        RECT 51.920 57.380 52.180 58.105 ;
        RECT 52.350 57.210 52.610 57.935 ;
        RECT 52.780 57.380 53.040 58.105 ;
        RECT 53.210 57.210 53.470 57.935 ;
        RECT 53.640 57.380 53.900 58.105 ;
        RECT 54.070 57.210 54.330 57.935 ;
        RECT 54.500 57.380 54.760 58.105 ;
        RECT 54.930 57.210 55.190 58.005 ;
        RECT 55.360 57.380 55.610 58.515 ;
        RECT 48.915 57.205 55.190 57.210 ;
        RECT 55.790 57.205 56.050 58.015 ;
        RECT 56.225 57.375 56.470 58.515 ;
        RECT 57.950 58.425 58.255 58.935 ;
        RECT 61.715 58.765 61.905 58.935 ;
        RECT 62.415 58.765 62.665 59.025 ;
        RECT 62.835 59.105 63.085 59.365 ;
        RECT 63.255 59.285 63.425 59.755 ;
        RECT 63.595 59.115 63.925 59.585 ;
        RECT 64.095 59.285 64.265 59.755 ;
        RECT 64.435 59.115 64.765 59.585 ;
        RECT 65.035 59.275 65.335 59.755 ;
        RECT 63.595 59.105 64.765 59.115 ;
        RECT 65.505 59.105 65.765 59.560 ;
        RECT 65.935 59.275 66.195 59.755 ;
        RECT 66.375 59.105 66.635 59.560 ;
        RECT 66.805 59.275 67.055 59.755 ;
        RECT 67.235 59.105 67.495 59.560 ;
        RECT 67.665 59.275 67.915 59.755 ;
        RECT 68.095 59.105 68.355 59.560 ;
        RECT 68.525 59.275 68.770 59.755 ;
        RECT 68.940 59.105 69.215 59.560 ;
        RECT 69.385 59.275 69.630 59.755 ;
        RECT 69.800 59.105 70.060 59.560 ;
        RECT 70.230 59.275 70.490 59.755 ;
        RECT 70.660 59.105 70.920 59.560 ;
        RECT 71.090 59.275 71.350 59.755 ;
        RECT 71.520 59.105 71.780 59.560 ;
        RECT 71.950 59.195 72.210 59.755 ;
        RECT 62.835 58.935 64.765 59.105 ;
        RECT 65.035 58.935 71.780 59.105 ;
        RECT 58.425 58.595 59.695 58.765 ;
        RECT 56.650 57.205 56.945 58.015 ;
        RECT 57.125 57.205 57.415 58.370 ;
        RECT 57.950 58.185 58.745 58.425 ;
        RECT 59.405 58.225 59.695 58.595 ;
        RECT 59.895 58.395 60.255 58.765 ;
        RECT 60.425 58.565 61.045 58.765 ;
        RECT 61.215 58.395 61.545 58.765 ;
        RECT 59.895 58.225 61.545 58.395 ;
        RECT 61.715 58.595 62.245 58.765 ;
        RECT 58.495 58.055 58.745 58.185 ;
        RECT 61.715 58.055 61.905 58.595 ;
        RECT 62.415 58.425 62.795 58.765 ;
        RECT 58.075 57.205 58.325 58.015 ;
        RECT 58.495 57.885 59.585 58.055 ;
        RECT 58.495 57.375 58.745 57.885 ;
        RECT 58.915 57.205 59.165 57.675 ;
        RECT 59.335 57.375 59.585 57.885 ;
        RECT 59.755 57.205 60.005 58.045 ;
        RECT 60.175 57.875 61.905 58.055 ;
        RECT 62.245 58.055 62.795 58.425 ;
        RECT 62.965 58.735 63.295 58.765 ;
        RECT 62.965 58.565 63.335 58.735 ;
        RECT 63.515 58.565 64.055 58.765 ;
        RECT 62.965 58.395 63.295 58.565 ;
        RECT 64.285 58.395 64.775 58.765 ;
        RECT 62.965 58.225 64.775 58.395 ;
        RECT 65.035 58.345 66.200 58.935 ;
        RECT 72.380 58.765 72.630 59.575 ;
        RECT 72.810 59.230 73.070 59.755 ;
        RECT 73.240 58.765 73.490 59.575 ;
        RECT 73.670 59.245 73.975 59.755 ;
        RECT 66.370 58.515 73.490 58.765 ;
        RECT 73.660 58.515 73.975 59.075 ;
        RECT 74.185 58.935 74.415 59.755 ;
        RECT 74.585 58.955 74.915 59.585 ;
        RECT 74.165 58.515 74.495 58.765 ;
        RECT 65.035 58.120 71.780 58.345 ;
        RECT 62.245 57.885 63.885 58.055 ;
        RECT 62.245 57.875 62.625 57.885 ;
        RECT 60.175 57.375 60.425 57.875 ;
        RECT 61.015 57.715 61.265 57.875 ;
        RECT 60.595 57.205 60.845 57.705 ;
        RECT 61.435 57.205 62.165 57.705 ;
        RECT 62.335 57.375 62.625 57.875 ;
        RECT 63.635 57.715 63.885 57.885 ;
        RECT 62.795 57.205 63.045 57.715 ;
        RECT 63.215 57.545 63.465 57.715 ;
        RECT 64.055 57.545 64.305 58.055 ;
        RECT 63.215 57.375 64.305 57.545 ;
        RECT 64.515 57.205 64.720 58.045 ;
        RECT 65.035 57.205 65.305 57.950 ;
        RECT 65.475 57.380 65.765 58.120 ;
        RECT 66.375 58.105 71.780 58.120 ;
        RECT 65.935 57.210 66.190 57.935 ;
        RECT 66.375 57.380 66.635 58.105 ;
        RECT 66.805 57.210 67.050 57.935 ;
        RECT 67.235 57.380 67.495 58.105 ;
        RECT 67.665 57.210 67.910 57.935 ;
        RECT 68.095 57.380 68.355 58.105 ;
        RECT 68.525 57.210 68.770 57.935 ;
        RECT 68.940 57.380 69.200 58.105 ;
        RECT 69.370 57.210 69.630 57.935 ;
        RECT 69.800 57.380 70.060 58.105 ;
        RECT 70.230 57.210 70.490 57.935 ;
        RECT 70.660 57.380 70.920 58.105 ;
        RECT 71.090 57.210 71.350 57.935 ;
        RECT 71.520 57.380 71.780 58.105 ;
        RECT 71.950 57.210 72.210 58.005 ;
        RECT 72.380 57.380 72.630 58.515 ;
        RECT 65.935 57.205 72.210 57.210 ;
        RECT 72.810 57.205 73.070 58.015 ;
        RECT 73.245 57.375 73.490 58.515 ;
        RECT 74.665 58.355 74.915 58.955 ;
        RECT 75.085 58.935 75.295 59.755 ;
        RECT 75.525 59.005 76.735 59.755 ;
        RECT 73.670 57.205 73.965 58.015 ;
        RECT 74.185 57.205 74.415 58.345 ;
        RECT 74.585 57.375 74.915 58.355 ;
        RECT 75.085 57.205 75.295 58.345 ;
        RECT 75.525 58.295 76.045 58.835 ;
        RECT 76.215 58.465 76.735 59.005 ;
        RECT 75.525 57.205 76.735 58.295 ;
        RECT 5.520 57.035 76.820 57.205 ;
        RECT 5.605 55.945 6.815 57.035 ;
        RECT 5.605 55.235 6.125 55.775 ;
        RECT 6.295 55.405 6.815 55.945 ;
        RECT 7.065 56.105 7.245 56.865 ;
        RECT 7.425 56.275 7.755 57.035 ;
        RECT 7.065 55.935 7.740 56.105 ;
        RECT 7.925 55.960 8.195 56.865 ;
        RECT 7.570 55.790 7.740 55.935 ;
        RECT 7.005 55.385 7.345 55.755 ;
        RECT 7.570 55.460 7.845 55.790 ;
        RECT 5.605 54.485 6.815 55.235 ;
        RECT 7.570 55.205 7.740 55.460 ;
        RECT 7.075 55.035 7.740 55.205 ;
        RECT 8.015 55.160 8.195 55.960 ;
        RECT 8.825 55.895 9.105 57.035 ;
        RECT 9.275 55.885 9.605 56.865 ;
        RECT 9.775 55.895 10.035 57.035 ;
        RECT 10.215 56.235 10.545 57.035 ;
        RECT 10.725 56.695 12.155 56.865 ;
        RECT 10.725 56.065 10.975 56.695 ;
        RECT 10.205 55.895 10.975 56.065 ;
        RECT 8.835 55.455 9.170 55.725 ;
        RECT 9.340 55.335 9.510 55.885 ;
        RECT 9.680 55.475 10.015 55.725 ;
        RECT 9.340 55.285 9.515 55.335 ;
        RECT 7.075 54.655 7.245 55.035 ;
        RECT 7.425 54.485 7.755 54.865 ;
        RECT 7.935 54.655 8.195 55.160 ;
        RECT 8.825 54.485 9.135 55.285 ;
        RECT 9.340 54.655 10.035 55.285 ;
        RECT 10.205 55.225 10.375 55.895 ;
        RECT 10.545 55.395 10.950 55.725 ;
        RECT 11.165 55.395 11.415 56.525 ;
        RECT 11.615 55.725 11.815 56.525 ;
        RECT 11.985 56.015 12.155 56.695 ;
        RECT 12.325 56.185 12.640 57.035 ;
        RECT 12.815 56.235 13.255 56.865 ;
        RECT 11.985 55.845 12.775 56.015 ;
        RECT 11.615 55.395 11.860 55.725 ;
        RECT 12.045 55.395 12.435 55.675 ;
        RECT 12.605 55.395 12.775 55.845 ;
        RECT 12.945 55.225 13.255 56.235 ;
        RECT 10.205 54.655 10.695 55.225 ;
        RECT 10.865 55.055 12.025 55.225 ;
        RECT 10.865 54.655 11.095 55.055 ;
        RECT 11.265 54.485 11.685 54.885 ;
        RECT 11.855 54.655 12.025 55.055 ;
        RECT 12.195 54.485 12.645 55.225 ;
        RECT 12.815 54.665 13.255 55.225 ;
        RECT 14.345 56.195 14.605 56.865 ;
        RECT 14.775 56.635 15.105 57.035 ;
        RECT 15.975 56.635 16.375 57.035 ;
        RECT 16.665 56.455 16.995 56.690 ;
        RECT 14.915 56.285 16.995 56.455 ;
        RECT 14.345 55.225 14.520 56.195 ;
        RECT 14.915 56.015 15.085 56.285 ;
        RECT 14.690 55.845 15.085 56.015 ;
        RECT 15.255 55.895 16.270 56.115 ;
        RECT 14.690 55.395 14.860 55.845 ;
        RECT 15.995 55.755 16.270 55.895 ;
        RECT 16.440 55.895 16.995 56.285 ;
        RECT 15.030 55.475 15.480 55.675 ;
        RECT 15.650 55.305 15.825 55.500 ;
        RECT 14.345 54.655 14.685 55.225 ;
        RECT 14.880 54.485 15.050 55.150 ;
        RECT 15.330 55.135 15.825 55.305 ;
        RECT 15.330 54.995 15.550 55.135 ;
        RECT 15.325 54.825 15.550 54.995 ;
        RECT 15.995 54.965 16.165 55.755 ;
        RECT 16.440 55.645 16.610 55.895 ;
        RECT 17.165 55.725 17.340 56.825 ;
        RECT 17.510 56.215 17.855 57.035 ;
        RECT 16.415 55.475 16.610 55.645 ;
        RECT 16.780 55.475 17.340 55.725 ;
        RECT 17.510 55.475 17.855 56.045 ;
        RECT 18.485 55.870 18.775 57.035 ;
        RECT 18.945 55.960 19.215 56.865 ;
        RECT 19.385 56.275 19.715 57.035 ;
        RECT 19.895 56.105 20.075 56.865 ;
        RECT 16.415 55.090 16.585 55.475 ;
        RECT 15.330 54.780 15.550 54.825 ;
        RECT 15.720 54.795 16.165 54.965 ;
        RECT 16.335 54.720 16.585 55.090 ;
        RECT 16.755 55.125 17.855 55.305 ;
        RECT 16.755 54.720 17.005 55.125 ;
        RECT 17.175 54.485 17.345 54.955 ;
        RECT 17.515 54.720 17.855 55.125 ;
        RECT 18.485 54.485 18.775 55.210 ;
        RECT 18.945 55.160 19.125 55.960 ;
        RECT 19.400 55.935 20.075 56.105 ;
        RECT 19.400 55.790 19.570 55.935 ;
        RECT 19.295 55.460 19.570 55.790 ;
        RECT 20.330 55.895 20.665 56.865 ;
        RECT 20.835 55.895 21.005 57.035 ;
        RECT 21.175 56.695 23.205 56.865 ;
        RECT 19.400 55.205 19.570 55.460 ;
        RECT 19.795 55.385 20.135 55.755 ;
        RECT 20.330 55.225 20.500 55.895 ;
        RECT 21.175 55.725 21.345 56.695 ;
        RECT 20.670 55.395 20.925 55.725 ;
        RECT 21.150 55.395 21.345 55.725 ;
        RECT 21.515 56.355 22.640 56.525 ;
        RECT 20.755 55.225 20.925 55.395 ;
        RECT 21.515 55.225 21.685 56.355 ;
        RECT 18.945 54.655 19.205 55.160 ;
        RECT 19.400 55.035 20.065 55.205 ;
        RECT 19.385 54.485 19.715 54.865 ;
        RECT 19.895 54.655 20.065 55.035 ;
        RECT 20.330 54.655 20.585 55.225 ;
        RECT 20.755 55.055 21.685 55.225 ;
        RECT 21.855 56.015 22.865 56.185 ;
        RECT 21.855 55.215 22.025 56.015 ;
        RECT 22.230 55.335 22.505 55.815 ;
        RECT 22.225 55.165 22.505 55.335 ;
        RECT 21.510 55.020 21.685 55.055 ;
        RECT 20.755 54.485 21.085 54.885 ;
        RECT 21.510 54.655 22.040 55.020 ;
        RECT 22.230 54.655 22.505 55.165 ;
        RECT 22.675 54.655 22.865 56.015 ;
        RECT 23.035 56.030 23.205 56.695 ;
        RECT 23.375 56.275 23.545 57.035 ;
        RECT 23.780 56.275 24.295 56.685 ;
        RECT 23.035 55.840 23.785 56.030 ;
        RECT 23.955 55.465 24.295 56.275 ;
        RECT 24.555 56.105 24.725 56.865 ;
        RECT 24.905 56.275 25.235 57.035 ;
        RECT 24.555 55.935 25.220 56.105 ;
        RECT 25.405 55.960 25.675 56.865 ;
        RECT 25.050 55.790 25.220 55.935 ;
        RECT 23.065 55.295 24.295 55.465 ;
        RECT 24.485 55.385 24.815 55.755 ;
        RECT 25.050 55.460 25.335 55.790 ;
        RECT 23.045 54.485 23.555 55.020 ;
        RECT 23.775 54.690 24.020 55.295 ;
        RECT 25.050 55.205 25.220 55.460 ;
        RECT 24.555 55.035 25.220 55.205 ;
        RECT 25.505 55.160 25.675 55.960 ;
        RECT 24.555 54.655 24.725 55.035 ;
        RECT 24.905 54.485 25.235 54.865 ;
        RECT 25.415 54.655 25.675 55.160 ;
        RECT 26.305 55.960 26.575 56.865 ;
        RECT 26.745 56.275 27.075 57.035 ;
        RECT 27.255 56.105 27.435 56.865 ;
        RECT 26.305 55.160 26.485 55.960 ;
        RECT 26.760 55.935 27.435 56.105 ;
        RECT 28.625 56.145 28.885 56.855 ;
        RECT 29.055 56.325 29.385 57.035 ;
        RECT 29.555 56.145 29.785 56.855 ;
        RECT 26.760 55.790 26.930 55.935 ;
        RECT 28.625 55.905 29.785 56.145 ;
        RECT 29.965 56.125 30.235 56.855 ;
        RECT 30.415 56.305 30.755 57.035 ;
        RECT 29.965 55.905 30.735 56.125 ;
        RECT 26.655 55.460 26.930 55.790 ;
        RECT 26.760 55.205 26.930 55.460 ;
        RECT 27.155 55.385 27.495 55.755 ;
        RECT 28.615 55.395 28.915 55.725 ;
        RECT 29.095 55.415 29.620 55.725 ;
        RECT 29.800 55.415 30.265 55.725 ;
        RECT 26.305 54.655 26.565 55.160 ;
        RECT 26.760 55.035 27.425 55.205 ;
        RECT 26.745 54.485 27.075 54.865 ;
        RECT 27.255 54.655 27.425 55.035 ;
        RECT 28.625 54.485 28.915 55.215 ;
        RECT 29.095 54.775 29.325 55.415 ;
        RECT 30.445 55.235 30.735 55.905 ;
        RECT 29.505 55.035 30.735 55.235 ;
        RECT 29.505 54.665 29.815 55.035 ;
        RECT 29.995 54.485 30.665 54.855 ;
        RECT 30.925 54.665 31.185 56.855 ;
        RECT 31.825 56.615 32.165 57.035 ;
        RECT 32.335 56.445 32.585 56.865 ;
        RECT 31.825 56.275 32.585 56.445 ;
        RECT 31.825 55.305 32.135 56.275 ;
        RECT 32.755 56.195 33.085 57.035 ;
        RECT 33.575 56.445 34.330 56.865 ;
        RECT 33.255 56.275 34.720 56.445 ;
        RECT 33.255 56.025 33.425 56.275 ;
        RECT 32.465 55.855 33.425 56.025 ;
        RECT 32.465 55.685 32.635 55.855 ;
        RECT 33.595 55.685 33.900 56.105 ;
        RECT 32.305 55.475 32.635 55.685 ;
        RECT 32.805 55.475 33.245 55.685 ;
        RECT 33.415 55.475 33.900 55.685 ;
        RECT 34.090 55.675 34.380 56.105 ;
        RECT 34.550 56.070 34.720 56.275 ;
        RECT 34.890 56.250 35.130 57.035 ;
        RECT 35.300 56.070 35.630 56.865 ;
        RECT 34.550 55.895 35.630 56.070 ;
        RECT 35.970 56.165 36.235 56.865 ;
        RECT 36.405 56.335 36.735 57.035 ;
        RECT 36.905 56.165 37.575 56.865 ;
        RECT 38.080 56.335 38.510 57.035 ;
        RECT 38.690 56.475 38.880 56.865 ;
        RECT 39.050 56.655 39.380 57.035 ;
        RECT 38.690 56.305 39.420 56.475 ;
        RECT 35.970 55.910 38.545 56.165 ;
        RECT 34.550 55.845 35.335 55.895 ;
        RECT 34.090 55.475 34.480 55.675 ;
        RECT 34.650 55.475 34.995 55.675 ;
        RECT 31.825 55.135 32.585 55.305 ;
        RECT 31.915 54.485 32.085 54.965 ;
        RECT 32.255 54.665 32.585 55.135 ;
        RECT 32.755 54.485 32.925 55.305 ;
        RECT 33.095 55.135 34.795 55.305 ;
        RECT 33.095 54.670 33.425 55.135 ;
        RECT 34.410 55.045 34.795 55.135 ;
        RECT 35.165 55.205 35.335 55.845 ;
        RECT 35.535 55.375 35.795 55.725 ;
        RECT 35.965 55.395 36.240 55.725 ;
        RECT 36.410 55.225 36.590 55.910 ;
        RECT 38.375 55.725 38.545 55.910 ;
        RECT 36.760 55.395 37.120 55.725 ;
        RECT 37.410 55.675 37.700 55.725 ;
        RECT 37.405 55.505 37.700 55.675 ;
        RECT 37.410 55.395 37.700 55.505 ;
        RECT 37.870 55.395 38.205 55.725 ;
        RECT 38.375 55.395 39.055 55.725 ;
        RECT 35.165 55.035 35.710 55.205 ;
        RECT 33.595 54.485 33.765 54.955 ;
        RECT 34.025 54.695 35.210 54.865 ;
        RECT 35.380 54.655 35.710 55.035 ;
        RECT 35.975 54.825 36.590 55.225 ;
        RECT 36.760 55.035 38.030 55.225 ;
        RECT 39.225 55.185 39.420 56.305 ;
        RECT 38.600 55.015 39.420 55.185 ;
        RECT 35.975 54.655 36.310 54.825 ;
        RECT 37.270 54.485 37.605 54.865 ;
        RECT 38.195 54.485 38.430 54.925 ;
        RECT 38.600 54.655 38.930 55.015 ;
        RECT 39.100 54.485 39.430 54.845 ;
        RECT 39.645 54.765 39.925 56.865 ;
        RECT 40.115 56.275 40.900 57.035 ;
        RECT 41.295 56.205 41.680 56.865 ;
        RECT 41.295 56.105 41.705 56.205 ;
        RECT 40.095 55.895 41.705 56.105 ;
        RECT 42.005 56.015 42.205 56.805 ;
        RECT 40.095 55.295 40.370 55.895 ;
        RECT 41.875 55.845 42.205 56.015 ;
        RECT 42.375 55.855 42.695 57.035 ;
        RECT 42.925 55.895 43.135 57.035 ;
        RECT 43.305 55.885 43.635 56.865 ;
        RECT 43.805 55.895 44.035 57.035 ;
        RECT 41.875 55.725 42.055 55.845 ;
        RECT 40.540 55.475 40.895 55.725 ;
        RECT 41.090 55.675 41.555 55.725 ;
        RECT 41.085 55.505 41.555 55.675 ;
        RECT 41.090 55.475 41.555 55.505 ;
        RECT 41.725 55.475 42.055 55.725 ;
        RECT 42.230 55.475 42.695 55.675 ;
        RECT 40.095 55.115 41.345 55.295 ;
        RECT 40.980 55.045 41.345 55.115 ;
        RECT 41.515 55.095 42.695 55.265 ;
        RECT 40.155 54.485 40.325 54.945 ;
        RECT 41.515 54.875 41.845 55.095 ;
        RECT 40.595 54.695 41.845 54.875 ;
        RECT 42.015 54.485 42.185 54.925 ;
        RECT 42.355 54.680 42.695 55.095 ;
        RECT 42.925 54.485 43.135 55.305 ;
        RECT 43.305 55.285 43.555 55.885 ;
        RECT 44.245 55.870 44.535 57.035 ;
        RECT 45.255 56.290 45.525 57.035 ;
        RECT 46.155 57.030 52.430 57.035 ;
        RECT 45.695 56.120 45.985 56.860 ;
        RECT 46.155 56.305 46.410 57.030 ;
        RECT 46.595 56.135 46.855 56.860 ;
        RECT 47.025 56.305 47.270 57.030 ;
        RECT 47.455 56.135 47.715 56.860 ;
        RECT 47.885 56.305 48.130 57.030 ;
        RECT 48.315 56.135 48.575 56.860 ;
        RECT 48.745 56.305 48.990 57.030 ;
        RECT 49.160 56.135 49.420 56.860 ;
        RECT 49.590 56.305 49.850 57.030 ;
        RECT 50.020 56.135 50.280 56.860 ;
        RECT 50.450 56.305 50.710 57.030 ;
        RECT 50.880 56.135 51.140 56.860 ;
        RECT 51.310 56.305 51.570 57.030 ;
        RECT 51.740 56.135 52.000 56.860 ;
        RECT 52.170 56.235 52.430 57.030 ;
        RECT 46.595 56.120 52.000 56.135 ;
        RECT 45.255 55.895 52.000 56.120 ;
        RECT 43.725 55.475 44.055 55.725 ;
        RECT 45.255 55.305 46.420 55.895 ;
        RECT 52.600 55.725 52.850 56.860 ;
        RECT 53.030 56.225 53.290 57.035 ;
        RECT 53.465 55.725 53.710 56.865 ;
        RECT 53.890 56.225 54.185 57.035 ;
        RECT 46.590 55.475 53.710 55.725 ;
        RECT 43.305 54.655 43.635 55.285 ;
        RECT 43.805 54.485 44.035 55.305 ;
        RECT 44.245 54.485 44.535 55.210 ;
        RECT 45.255 55.135 52.000 55.305 ;
        RECT 45.255 54.485 45.555 54.965 ;
        RECT 45.725 54.680 45.985 55.135 ;
        RECT 46.155 54.485 46.415 54.965 ;
        RECT 46.595 54.680 46.855 55.135 ;
        RECT 47.025 54.485 47.275 54.965 ;
        RECT 47.455 54.680 47.715 55.135 ;
        RECT 47.885 54.485 48.135 54.965 ;
        RECT 48.315 54.680 48.575 55.135 ;
        RECT 48.745 54.485 48.990 54.965 ;
        RECT 49.160 54.680 49.435 55.135 ;
        RECT 49.605 54.485 49.850 54.965 ;
        RECT 50.020 54.680 50.280 55.135 ;
        RECT 50.450 54.485 50.710 54.965 ;
        RECT 50.880 54.680 51.140 55.135 ;
        RECT 51.310 54.485 51.570 54.965 ;
        RECT 51.740 54.680 52.000 55.135 ;
        RECT 52.170 54.485 52.430 55.045 ;
        RECT 52.600 54.665 52.850 55.475 ;
        RECT 53.030 54.485 53.290 55.010 ;
        RECT 53.460 54.665 53.710 55.475 ;
        RECT 53.880 55.165 54.195 55.725 ;
        RECT 53.890 54.485 54.195 54.995 ;
        RECT 54.380 54.665 54.660 56.855 ;
        RECT 54.850 55.895 55.135 57.035 ;
        RECT 55.400 56.385 55.570 56.855 ;
        RECT 55.745 56.555 56.075 57.035 ;
        RECT 56.245 56.385 56.425 56.855 ;
        RECT 55.400 56.185 56.425 56.385 ;
        RECT 54.860 55.215 55.120 55.725 ;
        RECT 55.330 55.395 55.590 56.015 ;
        RECT 55.785 55.395 56.210 56.015 ;
        RECT 56.595 55.745 56.925 56.855 ;
        RECT 57.095 56.625 57.445 57.035 ;
        RECT 57.615 56.445 57.855 56.835 ;
        RECT 56.380 55.445 56.925 55.745 ;
        RECT 57.105 56.245 57.855 56.445 ;
        RECT 57.105 55.565 57.445 56.245 ;
        RECT 58.100 56.165 58.385 57.035 ;
        RECT 58.555 56.405 58.815 56.865 ;
        RECT 58.990 56.575 59.245 57.035 ;
        RECT 59.415 56.405 59.675 56.865 ;
        RECT 58.555 56.235 59.675 56.405 ;
        RECT 59.845 56.235 60.155 57.035 ;
        RECT 56.380 55.215 56.600 55.445 ;
        RECT 54.860 55.025 56.600 55.215 ;
        RECT 54.860 54.485 55.590 54.855 ;
        RECT 56.170 54.665 56.600 55.025 ;
        RECT 56.770 54.485 57.015 55.265 ;
        RECT 57.215 54.665 57.445 55.565 ;
        RECT 57.625 54.725 57.855 56.065 ;
        RECT 58.555 55.985 58.815 56.235 ;
        RECT 60.325 56.065 60.635 56.865 ;
        RECT 60.895 56.290 61.165 57.035 ;
        RECT 61.795 57.030 68.070 57.035 ;
        RECT 61.335 56.120 61.625 56.860 ;
        RECT 61.795 56.305 62.050 57.030 ;
        RECT 62.235 56.135 62.495 56.860 ;
        RECT 62.665 56.305 62.910 57.030 ;
        RECT 63.095 56.135 63.355 56.860 ;
        RECT 63.525 56.305 63.770 57.030 ;
        RECT 63.955 56.135 64.215 56.860 ;
        RECT 64.385 56.305 64.630 57.030 ;
        RECT 64.800 56.135 65.060 56.860 ;
        RECT 65.230 56.305 65.490 57.030 ;
        RECT 65.660 56.135 65.920 56.860 ;
        RECT 66.090 56.305 66.350 57.030 ;
        RECT 66.520 56.135 66.780 56.860 ;
        RECT 66.950 56.305 67.210 57.030 ;
        RECT 67.380 56.135 67.640 56.860 ;
        RECT 67.810 56.235 68.070 57.030 ;
        RECT 62.235 56.120 67.640 56.135 ;
        RECT 58.060 55.815 58.815 55.985 ;
        RECT 59.605 55.895 60.635 56.065 ;
        RECT 58.060 55.305 58.465 55.815 ;
        RECT 59.605 55.645 59.775 55.895 ;
        RECT 58.635 55.475 59.775 55.645 ;
        RECT 58.060 55.135 59.710 55.305 ;
        RECT 59.945 55.155 60.295 55.725 ;
        RECT 58.105 54.485 58.385 54.965 ;
        RECT 58.555 54.745 58.815 55.135 ;
        RECT 58.990 54.485 59.245 54.965 ;
        RECT 59.415 54.745 59.710 55.135 ;
        RECT 60.465 54.985 60.635 55.895 ;
        RECT 60.895 55.895 67.640 56.120 ;
        RECT 60.895 55.305 62.060 55.895 ;
        RECT 68.240 55.725 68.490 56.860 ;
        RECT 68.670 56.225 68.930 57.035 ;
        RECT 69.105 55.725 69.350 56.865 ;
        RECT 69.530 56.225 69.825 57.035 ;
        RECT 70.005 55.870 70.295 57.035 ;
        RECT 70.470 56.165 70.735 56.865 ;
        RECT 70.905 56.335 71.235 57.035 ;
        RECT 71.405 56.165 72.075 56.865 ;
        RECT 72.580 56.335 73.010 57.035 ;
        RECT 73.190 56.475 73.380 56.865 ;
        RECT 73.550 56.655 73.880 57.035 ;
        RECT 73.190 56.305 73.920 56.475 ;
        RECT 70.470 55.910 73.045 56.165 ;
        RECT 62.230 55.475 69.350 55.725 ;
        RECT 60.895 55.135 67.640 55.305 ;
        RECT 59.890 54.485 60.165 54.965 ;
        RECT 60.335 54.655 60.635 54.985 ;
        RECT 60.895 54.485 61.195 54.965 ;
        RECT 61.365 54.680 61.625 55.135 ;
        RECT 61.795 54.485 62.055 54.965 ;
        RECT 62.235 54.680 62.495 55.135 ;
        RECT 62.665 54.485 62.915 54.965 ;
        RECT 63.095 54.680 63.355 55.135 ;
        RECT 63.525 54.485 63.775 54.965 ;
        RECT 63.955 54.680 64.215 55.135 ;
        RECT 64.385 54.485 64.630 54.965 ;
        RECT 64.800 54.680 65.075 55.135 ;
        RECT 65.245 54.485 65.490 54.965 ;
        RECT 65.660 54.680 65.920 55.135 ;
        RECT 66.090 54.485 66.350 54.965 ;
        RECT 66.520 54.680 66.780 55.135 ;
        RECT 66.950 54.485 67.210 54.965 ;
        RECT 67.380 54.680 67.640 55.135 ;
        RECT 67.810 54.485 68.070 55.045 ;
        RECT 68.240 54.665 68.490 55.475 ;
        RECT 68.670 54.485 68.930 55.010 ;
        RECT 69.100 54.665 69.350 55.475 ;
        RECT 69.520 55.165 69.835 55.725 ;
        RECT 70.465 55.395 70.740 55.725 ;
        RECT 70.910 55.225 71.090 55.910 ;
        RECT 72.875 55.725 73.045 55.910 ;
        RECT 71.260 55.395 71.620 55.725 ;
        RECT 71.910 55.675 72.200 55.725 ;
        RECT 71.905 55.505 72.200 55.675 ;
        RECT 71.910 55.395 72.200 55.505 ;
        RECT 72.370 55.395 72.705 55.725 ;
        RECT 72.875 55.395 73.555 55.725 ;
        RECT 69.530 54.485 69.835 54.995 ;
        RECT 70.005 54.485 70.295 55.210 ;
        RECT 70.475 54.825 71.090 55.225 ;
        RECT 71.260 55.035 72.530 55.225 ;
        RECT 73.725 55.185 73.920 56.305 ;
        RECT 74.155 56.065 74.485 56.850 ;
        RECT 74.155 55.895 74.835 56.065 ;
        RECT 75.015 55.895 75.345 57.035 ;
        RECT 75.525 55.945 76.735 57.035 ;
        RECT 74.145 55.475 74.495 55.725 ;
        RECT 74.665 55.295 74.835 55.895 ;
        RECT 75.005 55.475 75.355 55.725 ;
        RECT 75.525 55.405 76.045 55.945 ;
        RECT 73.100 55.015 73.920 55.185 ;
        RECT 70.475 54.655 70.810 54.825 ;
        RECT 71.770 54.485 72.105 54.865 ;
        RECT 72.695 54.485 72.930 54.925 ;
        RECT 73.100 54.655 73.430 55.015 ;
        RECT 73.600 54.485 73.930 54.845 ;
        RECT 74.165 54.485 74.405 55.295 ;
        RECT 74.575 54.655 74.905 55.295 ;
        RECT 75.075 54.485 75.345 55.295 ;
        RECT 76.215 55.235 76.735 55.775 ;
        RECT 75.525 54.485 76.735 55.235 ;
        RECT 5.520 54.315 76.820 54.485 ;
        RECT 5.605 53.565 6.815 54.315 ;
        RECT 7.995 53.765 8.165 54.145 ;
        RECT 8.345 53.935 8.675 54.315 ;
        RECT 7.995 53.595 8.660 53.765 ;
        RECT 8.855 53.640 9.115 54.145 ;
        RECT 5.605 53.025 6.125 53.565 ;
        RECT 6.295 52.855 6.815 53.395 ;
        RECT 7.925 53.045 8.255 53.415 ;
        RECT 8.490 53.340 8.660 53.595 ;
        RECT 8.490 53.010 8.775 53.340 ;
        RECT 8.490 52.865 8.660 53.010 ;
        RECT 5.605 51.765 6.815 52.855 ;
        RECT 7.995 52.695 8.660 52.865 ;
        RECT 8.945 52.840 9.115 53.640 ;
        RECT 7.995 51.935 8.165 52.695 ;
        RECT 8.345 51.765 8.675 52.525 ;
        RECT 8.845 51.935 9.115 52.840 ;
        RECT 9.285 53.640 9.545 54.145 ;
        RECT 9.725 53.935 10.055 54.315 ;
        RECT 10.235 53.765 10.405 54.145 ;
        RECT 9.285 52.840 9.465 53.640 ;
        RECT 9.740 53.595 10.405 53.765 ;
        RECT 10.665 53.815 10.925 54.145 ;
        RECT 11.135 53.835 11.410 54.315 ;
        RECT 9.740 53.340 9.910 53.595 ;
        RECT 9.635 53.010 9.910 53.340 ;
        RECT 10.135 53.045 10.475 53.415 ;
        RECT 9.740 52.865 9.910 53.010 ;
        RECT 10.665 52.905 10.835 53.815 ;
        RECT 11.620 53.745 11.825 54.145 ;
        RECT 11.995 53.915 12.330 54.315 ;
        RECT 11.005 53.075 11.365 53.655 ;
        RECT 11.620 53.575 12.305 53.745 ;
        RECT 11.545 52.905 11.795 53.405 ;
        RECT 9.285 51.935 9.555 52.840 ;
        RECT 9.740 52.695 10.415 52.865 ;
        RECT 9.725 51.765 10.055 52.525 ;
        RECT 10.235 51.935 10.415 52.695 ;
        RECT 10.665 52.735 11.795 52.905 ;
        RECT 10.665 51.965 10.935 52.735 ;
        RECT 11.965 52.545 12.305 53.575 ;
        RECT 12.515 53.505 12.785 54.315 ;
        RECT 12.955 53.505 13.285 54.145 ;
        RECT 13.455 53.505 13.695 54.315 ;
        RECT 13.885 53.640 14.145 54.145 ;
        RECT 14.325 53.935 14.655 54.315 ;
        RECT 14.835 53.765 15.005 54.145 ;
        RECT 12.505 53.075 12.855 53.325 ;
        RECT 13.025 52.905 13.195 53.505 ;
        RECT 13.365 53.075 13.715 53.325 ;
        RECT 11.105 51.765 11.435 52.545 ;
        RECT 11.640 52.370 12.305 52.545 ;
        RECT 11.640 51.965 11.825 52.370 ;
        RECT 11.995 51.765 12.330 52.190 ;
        RECT 12.515 51.765 12.845 52.905 ;
        RECT 13.025 52.735 13.705 52.905 ;
        RECT 13.375 51.950 13.705 52.735 ;
        RECT 13.885 52.840 14.065 53.640 ;
        RECT 14.340 53.595 15.005 53.765 ;
        RECT 15.355 53.765 15.525 54.145 ;
        RECT 15.705 53.935 16.035 54.315 ;
        RECT 15.355 53.595 16.020 53.765 ;
        RECT 16.215 53.640 16.475 54.145 ;
        RECT 14.340 53.340 14.510 53.595 ;
        RECT 14.235 53.010 14.510 53.340 ;
        RECT 14.735 53.045 15.075 53.415 ;
        RECT 15.285 53.045 15.625 53.415 ;
        RECT 15.850 53.340 16.020 53.595 ;
        RECT 14.340 52.865 14.510 53.010 ;
        RECT 15.850 53.010 16.125 53.340 ;
        RECT 15.850 52.865 16.020 53.010 ;
        RECT 13.885 51.935 14.155 52.840 ;
        RECT 14.340 52.695 15.015 52.865 ;
        RECT 14.325 51.765 14.655 52.525 ;
        RECT 14.835 51.935 15.015 52.695 ;
        RECT 15.345 52.695 16.020 52.865 ;
        RECT 16.295 52.840 16.475 53.640 ;
        RECT 16.735 53.765 16.905 54.145 ;
        RECT 17.085 53.935 17.415 54.315 ;
        RECT 16.735 53.595 17.400 53.765 ;
        RECT 17.595 53.640 17.855 54.145 ;
        RECT 16.665 53.045 17.005 53.415 ;
        RECT 17.230 53.340 17.400 53.595 ;
        RECT 17.230 53.010 17.505 53.340 ;
        RECT 17.230 52.865 17.400 53.010 ;
        RECT 15.345 51.935 15.525 52.695 ;
        RECT 15.705 51.765 16.035 52.525 ;
        RECT 16.205 51.935 16.475 52.840 ;
        RECT 16.725 52.695 17.400 52.865 ;
        RECT 17.675 52.840 17.855 53.640 ;
        RECT 18.065 53.495 18.295 54.315 ;
        RECT 18.465 53.515 18.795 54.145 ;
        RECT 18.045 53.075 18.375 53.325 ;
        RECT 18.545 52.915 18.795 53.515 ;
        RECT 18.965 53.495 19.175 54.315 ;
        RECT 19.405 53.640 19.665 54.145 ;
        RECT 19.845 53.935 20.175 54.315 ;
        RECT 20.355 53.765 20.525 54.145 ;
        RECT 16.725 51.935 16.905 52.695 ;
        RECT 17.085 51.765 17.415 52.525 ;
        RECT 17.585 51.935 17.855 52.840 ;
        RECT 18.065 51.765 18.295 52.905 ;
        RECT 18.465 51.935 18.795 52.915 ;
        RECT 18.965 51.765 19.175 52.905 ;
        RECT 19.405 52.840 19.585 53.640 ;
        RECT 19.860 53.595 20.525 53.765 ;
        RECT 19.860 53.340 20.030 53.595 ;
        RECT 21.705 53.515 22.015 54.315 ;
        RECT 22.220 53.515 22.915 54.145 ;
        RECT 23.085 53.770 28.430 54.315 ;
        RECT 19.755 53.010 20.030 53.340 ;
        RECT 20.255 53.045 20.595 53.415 ;
        RECT 21.715 53.075 22.050 53.345 ;
        RECT 19.860 52.865 20.030 53.010 ;
        RECT 22.220 52.915 22.390 53.515 ;
        RECT 22.560 53.075 22.895 53.325 ;
        RECT 24.670 52.940 25.010 53.770 ;
        RECT 28.605 53.545 31.195 54.315 ;
        RECT 31.365 53.590 31.655 54.315 ;
        RECT 31.825 53.555 32.535 54.145 ;
        RECT 33.045 53.785 33.375 54.145 ;
        RECT 33.575 53.955 33.905 54.315 ;
        RECT 34.075 53.785 34.405 54.145 ;
        RECT 33.045 53.575 34.405 53.785 ;
        RECT 35.505 53.640 35.765 54.145 ;
        RECT 35.945 53.935 36.275 54.315 ;
        RECT 36.455 53.765 36.625 54.145 ;
        RECT 19.405 51.935 19.675 52.840 ;
        RECT 19.860 52.695 20.535 52.865 ;
        RECT 19.845 51.765 20.175 52.525 ;
        RECT 20.355 51.935 20.535 52.695 ;
        RECT 21.705 51.765 21.985 52.905 ;
        RECT 22.155 51.935 22.485 52.915 ;
        RECT 22.655 51.765 22.915 52.905 ;
        RECT 26.490 52.200 26.840 53.450 ;
        RECT 28.605 53.025 29.815 53.545 ;
        RECT 29.985 52.855 31.195 53.375 ;
        RECT 23.085 51.765 28.430 52.200 ;
        RECT 28.605 51.765 31.195 52.855 ;
        RECT 31.365 51.765 31.655 52.930 ;
        RECT 31.825 52.585 32.030 53.555 ;
        RECT 32.200 52.785 32.530 53.325 ;
        RECT 32.705 53.075 33.200 53.405 ;
        RECT 33.520 53.075 33.895 53.405 ;
        RECT 34.105 53.075 34.415 53.405 ;
        RECT 32.705 52.785 33.030 53.075 ;
        RECT 33.225 52.585 33.555 52.805 ;
        RECT 31.825 52.355 33.555 52.585 ;
        RECT 31.825 51.935 32.525 52.355 ;
        RECT 32.725 51.765 33.055 52.125 ;
        RECT 33.225 51.955 33.555 52.355 ;
        RECT 33.725 52.105 33.895 53.075 ;
        RECT 35.505 52.840 35.685 53.640 ;
        RECT 35.960 53.595 36.625 53.765 ;
        RECT 35.960 53.340 36.130 53.595 ;
        RECT 36.925 53.495 37.155 54.315 ;
        RECT 37.325 53.515 37.655 54.145 ;
        RECT 35.855 53.010 36.130 53.340 ;
        RECT 36.355 53.045 36.695 53.415 ;
        RECT 36.905 53.075 37.235 53.325 ;
        RECT 35.960 52.865 36.130 53.010 ;
        RECT 37.405 52.915 37.655 53.515 ;
        RECT 37.825 53.495 38.035 54.315 ;
        RECT 38.355 53.765 38.525 54.145 ;
        RECT 38.705 53.935 39.035 54.315 ;
        RECT 38.355 53.595 39.020 53.765 ;
        RECT 39.215 53.640 39.475 54.145 ;
        RECT 38.285 53.045 38.615 53.415 ;
        RECT 38.850 53.340 39.020 53.595 ;
        RECT 34.075 51.765 34.405 52.825 ;
        RECT 35.505 51.935 35.775 52.840 ;
        RECT 35.960 52.695 36.635 52.865 ;
        RECT 35.945 51.765 36.275 52.525 ;
        RECT 36.455 51.935 36.635 52.695 ;
        RECT 36.925 51.765 37.155 52.905 ;
        RECT 37.325 51.935 37.655 52.915 ;
        RECT 38.850 53.010 39.135 53.340 ;
        RECT 37.825 51.765 38.035 52.905 ;
        RECT 38.850 52.865 39.020 53.010 ;
        RECT 38.355 52.695 39.020 52.865 ;
        RECT 39.305 52.840 39.475 53.640 ;
        RECT 39.655 53.585 39.955 54.315 ;
        RECT 40.135 53.405 40.365 54.025 ;
        RECT 40.565 53.755 40.790 54.135 ;
        RECT 40.960 53.925 41.290 54.315 ;
        RECT 40.565 53.575 40.895 53.755 ;
        RECT 39.660 53.075 39.955 53.405 ;
        RECT 40.135 53.075 40.550 53.405 ;
        RECT 40.720 52.905 40.895 53.575 ;
        RECT 41.065 53.075 41.305 53.725 ;
        RECT 41.490 53.550 41.945 54.315 ;
        RECT 42.220 53.935 43.520 54.145 ;
        RECT 43.775 53.955 44.105 54.315 ;
        RECT 43.350 53.785 43.520 53.935 ;
        RECT 44.275 53.815 44.535 54.145 ;
        RECT 42.420 53.325 42.640 53.725 ;
        RECT 41.485 53.125 41.975 53.325 ;
        RECT 42.165 53.115 42.640 53.325 ;
        RECT 42.885 53.325 43.095 53.725 ;
        RECT 43.350 53.660 44.105 53.785 ;
        RECT 43.350 53.615 44.195 53.660 ;
        RECT 43.925 53.495 44.195 53.615 ;
        RECT 42.885 53.115 43.215 53.325 ;
        RECT 43.385 53.055 43.795 53.360 ;
        RECT 38.355 51.935 38.525 52.695 ;
        RECT 38.705 51.765 39.035 52.525 ;
        RECT 39.205 51.935 39.475 52.840 ;
        RECT 39.655 52.545 40.550 52.875 ;
        RECT 40.720 52.715 41.305 52.905 ;
        RECT 39.655 52.375 40.860 52.545 ;
        RECT 39.655 51.945 39.985 52.375 ;
        RECT 40.165 51.765 40.360 52.205 ;
        RECT 40.530 51.945 40.860 52.375 ;
        RECT 41.030 51.945 41.305 52.715 ;
        RECT 41.490 52.885 42.665 52.945 ;
        RECT 44.025 52.920 44.195 53.495 ;
        RECT 43.995 52.885 44.195 52.920 ;
        RECT 41.490 52.775 44.195 52.885 ;
        RECT 41.490 52.155 41.745 52.775 ;
        RECT 42.335 52.715 44.135 52.775 ;
        RECT 42.335 52.685 42.665 52.715 ;
        RECT 44.365 52.615 44.535 53.815 ;
        RECT 41.995 52.515 42.180 52.605 ;
        RECT 42.770 52.515 43.605 52.525 ;
        RECT 41.995 52.315 43.605 52.515 ;
        RECT 41.995 52.275 42.225 52.315 ;
        RECT 41.490 51.935 41.825 52.155 ;
        RECT 42.830 51.765 43.185 52.145 ;
        RECT 43.355 51.935 43.605 52.315 ;
        RECT 43.855 51.765 44.105 52.545 ;
        RECT 44.275 51.935 44.535 52.615 ;
        RECT 44.705 53.495 45.390 54.135 ;
        RECT 45.560 53.495 45.730 54.315 ;
        RECT 45.900 53.665 46.230 54.130 ;
        RECT 46.400 53.845 46.570 54.315 ;
        RECT 46.830 53.925 48.015 54.095 ;
        RECT 48.185 53.755 48.515 54.145 ;
        RECT 47.215 53.665 47.600 53.755 ;
        RECT 45.900 53.495 47.600 53.665 ;
        RECT 48.005 53.575 48.515 53.755 ;
        RECT 48.845 53.815 49.105 54.145 ;
        RECT 49.275 53.955 49.605 54.315 ;
        RECT 49.860 53.935 51.160 54.145 ;
        RECT 44.705 52.525 44.955 53.495 ;
        RECT 45.125 53.115 45.460 53.325 ;
        RECT 45.630 53.115 46.080 53.325 ;
        RECT 46.270 53.295 46.755 53.325 ;
        RECT 46.270 53.125 46.775 53.295 ;
        RECT 46.270 53.115 46.755 53.125 ;
        RECT 45.290 52.945 45.460 53.115 ;
        RECT 45.290 52.775 46.210 52.945 ;
        RECT 44.705 51.935 45.370 52.525 ;
        RECT 45.540 51.765 45.870 52.605 ;
        RECT 46.040 52.525 46.210 52.775 ;
        RECT 46.380 52.695 46.755 53.115 ;
        RECT 46.945 53.075 47.325 53.325 ;
        RECT 47.505 53.115 47.835 53.325 ;
        RECT 46.945 52.695 47.265 53.075 ;
        RECT 48.005 52.945 48.175 53.575 ;
        RECT 48.345 53.115 48.675 53.405 ;
        RECT 47.435 52.775 48.520 52.945 ;
        RECT 47.435 52.525 47.605 52.775 ;
        RECT 46.040 52.355 47.605 52.525 ;
        RECT 46.380 51.935 47.185 52.355 ;
        RECT 47.775 51.765 48.025 52.605 ;
        RECT 48.220 51.935 48.520 52.775 ;
        RECT 48.845 52.615 49.015 53.815 ;
        RECT 49.860 53.785 50.030 53.935 ;
        RECT 49.275 53.660 50.030 53.785 ;
        RECT 49.185 53.615 50.030 53.660 ;
        RECT 49.185 53.495 49.455 53.615 ;
        RECT 49.185 52.920 49.355 53.495 ;
        RECT 49.585 53.055 49.995 53.360 ;
        RECT 50.285 53.325 50.495 53.725 ;
        RECT 50.165 53.115 50.495 53.325 ;
        RECT 50.740 53.325 50.960 53.725 ;
        RECT 51.435 53.550 51.890 54.315 ;
        RECT 52.085 53.505 52.325 54.315 ;
        RECT 52.495 53.505 52.825 54.145 ;
        RECT 52.995 53.505 53.265 54.315 ;
        RECT 53.445 53.515 53.785 54.145 ;
        RECT 53.955 53.515 54.205 54.315 ;
        RECT 54.395 53.665 54.725 54.145 ;
        RECT 54.895 53.855 55.120 54.315 ;
        RECT 55.290 53.665 55.620 54.145 ;
        RECT 50.740 53.115 51.215 53.325 ;
        RECT 51.405 53.125 51.895 53.325 ;
        RECT 52.065 53.075 52.415 53.325 ;
        RECT 49.185 52.885 49.385 52.920 ;
        RECT 50.715 52.885 51.890 52.945 ;
        RECT 52.585 52.905 52.755 53.505 ;
        RECT 52.925 53.075 53.275 53.325 ;
        RECT 53.445 52.905 53.620 53.515 ;
        RECT 54.395 53.495 55.620 53.665 ;
        RECT 56.250 53.535 56.750 54.145 ;
        RECT 57.125 53.590 57.415 54.315 ;
        RECT 57.585 53.805 57.890 54.315 ;
        RECT 53.790 53.155 54.485 53.325 ;
        RECT 54.315 52.905 54.485 53.155 ;
        RECT 54.660 53.125 55.080 53.325 ;
        RECT 55.250 53.125 55.580 53.325 ;
        RECT 55.750 53.125 56.080 53.325 ;
        RECT 56.250 52.905 56.420 53.535 ;
        RECT 56.605 53.075 56.955 53.325 ;
        RECT 57.585 53.075 57.900 53.635 ;
        RECT 58.070 53.325 58.320 54.135 ;
        RECT 58.490 53.790 58.750 54.315 ;
        RECT 58.930 53.325 59.180 54.135 ;
        RECT 59.350 53.755 59.610 54.315 ;
        RECT 59.780 53.665 60.040 54.120 ;
        RECT 60.210 53.835 60.470 54.315 ;
        RECT 60.640 53.665 60.900 54.120 ;
        RECT 61.070 53.835 61.330 54.315 ;
        RECT 61.500 53.665 61.760 54.120 ;
        RECT 61.930 53.835 62.175 54.315 ;
        RECT 62.345 53.665 62.620 54.120 ;
        RECT 62.790 53.835 63.035 54.315 ;
        RECT 63.205 53.665 63.465 54.120 ;
        RECT 63.645 53.835 63.895 54.315 ;
        RECT 64.065 53.665 64.325 54.120 ;
        RECT 64.505 53.835 64.755 54.315 ;
        RECT 64.925 53.665 65.185 54.120 ;
        RECT 65.365 53.835 65.625 54.315 ;
        RECT 65.795 53.665 66.055 54.120 ;
        RECT 66.225 53.835 66.525 54.315 ;
        RECT 59.780 53.495 66.525 53.665 ;
        RECT 58.070 53.075 65.190 53.325 ;
        RECT 49.185 52.775 51.890 52.885 ;
        RECT 49.245 52.715 51.045 52.775 ;
        RECT 50.715 52.685 51.045 52.715 ;
        RECT 48.845 51.935 49.105 52.615 ;
        RECT 49.275 51.765 49.525 52.545 ;
        RECT 49.775 52.515 50.610 52.525 ;
        RECT 51.200 52.515 51.385 52.605 ;
        RECT 49.775 52.315 51.385 52.515 ;
        RECT 49.775 51.935 50.025 52.315 ;
        RECT 51.155 52.275 51.385 52.315 ;
        RECT 51.635 52.155 51.890 52.775 ;
        RECT 50.195 51.765 50.550 52.145 ;
        RECT 51.555 51.935 51.890 52.155 ;
        RECT 52.075 52.735 52.755 52.905 ;
        RECT 52.075 51.950 52.405 52.735 ;
        RECT 52.935 51.765 53.265 52.905 ;
        RECT 53.445 51.935 53.785 52.905 ;
        RECT 53.955 51.765 54.125 52.905 ;
        RECT 54.315 52.735 56.750 52.905 ;
        RECT 54.395 51.765 54.645 52.565 ;
        RECT 55.290 51.935 55.620 52.735 ;
        RECT 55.920 51.765 56.250 52.565 ;
        RECT 56.420 51.935 56.750 52.735 ;
        RECT 57.125 51.765 57.415 52.930 ;
        RECT 57.595 51.765 57.890 52.575 ;
        RECT 58.070 51.935 58.315 53.075 ;
        RECT 58.490 51.765 58.750 52.575 ;
        RECT 58.930 51.940 59.180 53.075 ;
        RECT 65.360 52.955 66.525 53.495 ;
        RECT 66.785 53.565 67.995 54.315 ;
        RECT 68.170 53.685 68.505 54.145 ;
        RECT 68.675 53.855 68.870 54.315 ;
        RECT 69.115 53.935 71.140 54.145 ;
        RECT 66.785 53.025 67.305 53.565 ;
        RECT 68.170 53.495 68.860 53.685 ;
        RECT 69.115 53.495 69.365 53.935 ;
        RECT 69.535 53.495 70.720 53.765 ;
        RECT 70.890 53.685 71.140 53.935 ;
        RECT 71.310 53.855 71.480 54.315 ;
        RECT 71.650 53.685 71.980 54.145 ;
        RECT 72.150 53.855 72.390 54.315 ;
        RECT 72.600 53.685 72.930 54.145 ;
        RECT 73.245 53.805 73.485 54.315 ;
        RECT 73.655 53.805 73.945 54.145 ;
        RECT 74.175 53.805 74.490 54.315 ;
        RECT 70.890 53.495 72.930 53.685 ;
        RECT 65.360 52.905 66.555 52.955 ;
        RECT 59.780 52.785 66.555 52.905 ;
        RECT 67.475 52.855 67.995 53.395 ;
        RECT 68.690 53.325 68.860 53.495 ;
        RECT 68.190 53.125 68.520 53.325 ;
        RECT 68.690 53.125 70.285 53.325 ;
        RECT 68.690 52.955 68.860 53.125 ;
        RECT 70.455 52.955 70.720 53.495 ;
        RECT 73.285 53.465 73.485 53.635 ;
        RECT 71.235 53.125 73.020 53.325 ;
        RECT 73.290 53.075 73.485 53.465 ;
        RECT 59.780 52.680 66.525 52.785 ;
        RECT 59.780 52.665 65.185 52.680 ;
        RECT 59.350 51.770 59.610 52.565 ;
        RECT 59.780 51.940 60.040 52.665 ;
        RECT 60.210 51.770 60.470 52.495 ;
        RECT 60.640 51.940 60.900 52.665 ;
        RECT 61.070 51.770 61.330 52.495 ;
        RECT 61.500 51.940 61.760 52.665 ;
        RECT 61.930 51.770 62.190 52.495 ;
        RECT 62.360 51.940 62.620 52.665 ;
        RECT 62.790 51.770 63.035 52.495 ;
        RECT 63.205 51.940 63.465 52.665 ;
        RECT 63.650 51.770 63.895 52.495 ;
        RECT 64.065 51.940 64.325 52.665 ;
        RECT 64.510 51.770 64.755 52.495 ;
        RECT 64.925 51.940 65.185 52.665 ;
        RECT 65.370 51.770 65.625 52.495 ;
        RECT 65.795 51.940 66.085 52.680 ;
        RECT 59.350 51.765 65.625 51.770 ;
        RECT 66.255 51.765 66.525 52.510 ;
        RECT 66.785 51.765 67.995 52.855 ;
        RECT 68.170 52.735 68.860 52.955 ;
        RECT 68.170 51.935 68.505 52.735 ;
        RECT 69.050 52.565 69.365 52.955 ;
        RECT 68.675 51.765 69.365 52.565 ;
        RECT 69.535 52.735 72.400 52.955 ;
        RECT 73.655 52.905 73.835 53.805 ;
        RECT 74.660 53.745 74.830 54.015 ;
        RECT 75.000 53.915 75.330 54.315 ;
        RECT 74.005 53.075 74.415 53.635 ;
        RECT 74.660 53.575 75.355 53.745 ;
        RECT 74.585 52.905 74.755 53.405 ;
        RECT 69.535 51.935 69.865 52.735 ;
        RECT 70.035 51.765 70.205 52.565 ;
        RECT 70.375 51.935 70.720 52.735 ;
        RECT 70.890 51.765 71.060 52.565 ;
        RECT 71.230 51.935 71.560 52.735 ;
        RECT 71.730 51.765 71.900 52.565 ;
        RECT 72.070 51.935 72.400 52.735 ;
        RECT 72.600 51.765 72.930 52.905 ;
        RECT 73.295 52.735 74.755 52.905 ;
        RECT 73.295 52.560 73.655 52.735 ;
        RECT 74.925 52.565 75.355 53.575 ;
        RECT 75.525 53.565 76.735 54.315 ;
        RECT 74.240 51.765 74.410 52.565 ;
        RECT 74.580 52.395 75.355 52.565 ;
        RECT 75.525 52.855 76.045 53.395 ;
        RECT 76.215 53.025 76.735 53.565 ;
        RECT 74.580 51.935 74.910 52.395 ;
        RECT 75.080 51.765 75.250 52.225 ;
        RECT 75.525 51.765 76.735 52.855 ;
        RECT 5.520 51.595 76.820 51.765 ;
        RECT 5.605 50.505 6.815 51.595 ;
        RECT 5.605 49.795 6.125 50.335 ;
        RECT 6.295 49.965 6.815 50.505 ;
        RECT 8.090 50.625 8.480 50.800 ;
        RECT 8.965 50.795 9.295 51.595 ;
        RECT 9.465 50.805 10.000 51.425 ;
        RECT 8.090 50.455 9.515 50.625 ;
        RECT 5.605 49.045 6.815 49.795 ;
        RECT 7.965 49.725 8.320 50.285 ;
        RECT 8.490 49.555 8.660 50.455 ;
        RECT 8.830 49.725 9.095 50.285 ;
        RECT 9.345 49.955 9.515 50.455 ;
        RECT 9.685 49.785 10.000 50.805 ;
        RECT 10.205 50.640 10.475 51.595 ;
        RECT 8.070 49.045 8.310 49.555 ;
        RECT 8.490 49.225 8.770 49.555 ;
        RECT 9.000 49.045 9.215 49.555 ;
        RECT 9.385 49.215 10.000 49.785 ;
        RECT 10.660 50.540 10.965 51.325 ;
        RECT 11.145 51.125 11.830 51.595 ;
        RECT 11.140 50.605 11.835 50.915 ;
        RECT 10.660 49.735 10.835 50.540 ;
        RECT 12.010 50.435 12.295 51.380 ;
        RECT 12.495 51.145 12.825 51.595 ;
        RECT 12.995 50.975 13.165 51.405 ;
        RECT 11.435 50.285 12.295 50.435 ;
        RECT 11.005 50.265 12.295 50.285 ;
        RECT 12.485 50.745 13.165 50.975 ;
        RECT 13.515 50.975 13.685 51.405 ;
        RECT 13.855 51.145 14.185 51.595 ;
        RECT 13.515 50.745 14.190 50.975 ;
        RECT 11.005 49.905 11.995 50.265 ;
        RECT 12.485 50.095 12.720 50.745 ;
        RECT 10.205 49.045 10.475 49.680 ;
        RECT 10.660 49.215 10.895 49.735 ;
        RECT 11.825 49.570 11.995 49.905 ;
        RECT 12.165 49.765 12.720 50.095 ;
        RECT 12.505 49.615 12.720 49.765 ;
        RECT 12.890 49.895 13.190 50.575 ;
        RECT 12.890 49.725 13.195 49.895 ;
        RECT 13.485 49.725 13.785 50.575 ;
        RECT 13.955 50.095 14.190 50.745 ;
        RECT 14.360 50.435 14.645 51.380 ;
        RECT 14.825 51.125 15.510 51.595 ;
        RECT 14.820 50.605 15.515 50.915 ;
        RECT 15.690 50.540 15.995 51.325 ;
        RECT 14.360 50.285 15.220 50.435 ;
        RECT 14.360 50.265 15.645 50.285 ;
        RECT 13.955 49.765 14.490 50.095 ;
        RECT 14.660 49.905 15.645 50.265 ;
        RECT 13.955 49.615 14.175 49.765 ;
        RECT 11.065 49.045 11.465 49.540 ;
        RECT 11.825 49.375 12.225 49.570 ;
        RECT 12.055 49.230 12.225 49.375 ;
        RECT 12.505 49.240 12.745 49.615 ;
        RECT 12.915 49.045 13.245 49.550 ;
        RECT 13.430 49.045 13.765 49.550 ;
        RECT 13.935 49.240 14.175 49.615 ;
        RECT 14.660 49.570 14.830 49.905 ;
        RECT 15.820 49.735 15.995 50.540 ;
        RECT 16.655 50.985 16.985 51.415 ;
        RECT 17.165 51.155 17.360 51.595 ;
        RECT 17.530 50.985 17.860 51.415 ;
        RECT 16.655 50.815 17.860 50.985 ;
        RECT 16.655 50.485 17.550 50.815 ;
        RECT 18.030 50.645 18.305 51.415 ;
        RECT 17.720 50.455 18.305 50.645 ;
        RECT 16.660 49.955 16.955 50.285 ;
        RECT 17.135 49.955 17.550 50.285 ;
        RECT 14.455 49.375 14.830 49.570 ;
        RECT 14.455 49.230 14.625 49.375 ;
        RECT 15.190 49.045 15.585 49.540 ;
        RECT 15.755 49.215 15.995 49.735 ;
        RECT 16.655 49.045 16.955 49.775 ;
        RECT 17.135 49.335 17.365 49.955 ;
        RECT 17.720 49.785 17.895 50.455 ;
        RECT 18.485 50.430 18.775 51.595 ;
        RECT 19.875 50.535 20.205 51.385 ;
        RECT 19.875 50.405 20.095 50.535 ;
        RECT 20.375 50.455 20.625 51.595 ;
        RECT 20.815 50.955 21.065 51.375 ;
        RECT 21.295 51.125 21.625 51.595 ;
        RECT 21.855 50.955 22.105 51.375 ;
        RECT 20.815 50.785 22.105 50.955 ;
        RECT 22.285 50.955 22.615 51.385 ;
        RECT 22.285 50.785 22.740 50.955 ;
        RECT 17.565 49.605 17.895 49.785 ;
        RECT 18.065 49.635 18.305 50.285 ;
        RECT 19.875 49.770 20.065 50.405 ;
        RECT 20.805 50.285 21.020 50.615 ;
        RECT 20.235 49.955 20.545 50.285 ;
        RECT 20.715 49.955 21.020 50.285 ;
        RECT 21.195 49.955 21.480 50.615 ;
        RECT 21.675 49.955 21.940 50.615 ;
        RECT 22.155 49.955 22.400 50.615 ;
        RECT 20.375 49.785 20.545 49.955 ;
        RECT 22.570 49.785 22.740 50.785 ;
        RECT 23.090 50.455 23.410 51.595 ;
        RECT 23.590 50.285 23.785 51.335 ;
        RECT 23.965 50.745 24.295 51.425 ;
        RECT 24.495 50.795 24.750 51.595 ;
        RECT 24.945 50.755 25.200 51.425 ;
        RECT 25.370 50.835 25.700 51.595 ;
        RECT 25.870 50.995 26.120 51.425 ;
        RECT 26.290 51.175 26.645 51.595 ;
        RECT 26.835 51.255 28.005 51.425 ;
        RECT 26.835 51.215 27.165 51.255 ;
        RECT 27.275 50.995 27.505 51.085 ;
        RECT 25.870 50.755 27.505 50.995 ;
        RECT 27.675 50.755 28.005 51.255 ;
        RECT 24.945 50.745 25.155 50.755 ;
        RECT 23.965 50.465 24.315 50.745 ;
        RECT 23.150 50.235 23.410 50.285 ;
        RECT 23.145 50.065 23.410 50.235 ;
        RECT 23.150 49.955 23.410 50.065 ;
        RECT 23.590 49.955 23.975 50.285 ;
        RECT 24.145 50.085 24.315 50.465 ;
        RECT 24.505 50.255 24.750 50.615 ;
        RECT 24.145 49.915 24.665 50.085 ;
        RECT 17.565 49.225 17.790 49.605 ;
        RECT 17.960 49.045 18.290 49.435 ;
        RECT 18.485 49.045 18.775 49.770 ;
        RECT 19.875 49.260 20.205 49.770 ;
        RECT 20.375 49.615 22.740 49.785 ;
        RECT 20.375 49.045 20.705 49.445 ;
        RECT 21.755 49.275 22.085 49.615 ;
        RECT 23.090 49.575 24.305 49.745 ;
        RECT 22.255 49.045 22.585 49.445 ;
        RECT 23.090 49.225 23.380 49.575 ;
        RECT 23.575 49.045 23.905 49.405 ;
        RECT 24.075 49.270 24.305 49.575 ;
        RECT 24.495 49.350 24.665 49.915 ;
        RECT 24.945 49.625 25.115 50.745 ;
        RECT 28.175 50.585 28.345 51.425 ;
        RECT 25.285 50.415 28.345 50.585 ;
        RECT 28.610 50.875 28.945 51.385 ;
        RECT 25.285 49.865 25.455 50.415 ;
        RECT 25.685 50.035 26.050 50.235 ;
        RECT 26.220 50.035 26.550 50.235 ;
        RECT 25.285 49.695 26.085 49.865 ;
        RECT 24.945 49.545 25.130 49.625 ;
        RECT 24.945 49.215 25.200 49.545 ;
        RECT 25.415 49.045 25.745 49.525 ;
        RECT 25.915 49.465 26.085 49.695 ;
        RECT 26.265 49.635 26.550 50.035 ;
        RECT 26.820 50.035 27.295 50.235 ;
        RECT 27.465 50.035 27.910 50.235 ;
        RECT 28.080 50.035 28.430 50.245 ;
        RECT 26.820 49.635 27.100 50.035 ;
        RECT 27.280 49.695 28.345 49.865 ;
        RECT 27.280 49.465 27.450 49.695 ;
        RECT 25.915 49.215 27.450 49.465 ;
        RECT 27.675 49.045 28.005 49.525 ;
        RECT 28.175 49.215 28.345 49.695 ;
        RECT 28.610 49.520 28.865 50.875 ;
        RECT 29.195 50.795 29.525 51.595 ;
        RECT 29.770 51.005 30.055 51.425 ;
        RECT 30.310 51.175 30.640 51.595 ;
        RECT 30.865 51.255 32.025 51.425 ;
        RECT 30.865 51.005 31.195 51.255 ;
        RECT 29.770 50.835 31.195 51.005 ;
        RECT 31.425 50.625 31.595 51.085 ;
        RECT 31.855 50.755 32.025 51.255 ;
        RECT 29.225 50.455 31.595 50.625 ;
        RECT 29.225 50.285 29.395 50.455 ;
        RECT 31.845 50.405 32.055 50.575 ;
        RECT 32.285 50.485 32.545 51.425 ;
        RECT 32.715 51.195 33.045 51.595 ;
        RECT 34.190 51.330 34.445 51.425 ;
        RECT 33.305 51.160 34.445 51.330 ;
        RECT 34.615 51.215 34.945 51.385 ;
        RECT 33.305 50.935 33.475 51.160 ;
        RECT 32.715 50.765 33.475 50.935 ;
        RECT 34.190 51.025 34.445 51.160 ;
        RECT 31.845 50.285 32.050 50.405 ;
        RECT 29.090 49.955 29.395 50.285 ;
        RECT 29.590 50.235 29.840 50.285 ;
        RECT 29.585 50.065 29.840 50.235 ;
        RECT 29.590 49.955 29.840 50.065 ;
        RECT 29.225 49.785 29.395 49.955 ;
        RECT 30.050 49.895 30.320 50.285 ;
        RECT 30.510 49.895 30.800 50.285 ;
        RECT 29.225 49.615 29.785 49.785 ;
        RECT 30.045 49.725 30.320 49.895 ;
        RECT 30.505 49.725 30.800 49.895 ;
        RECT 30.050 49.625 30.320 49.725 ;
        RECT 30.510 49.625 30.800 49.725 ;
        RECT 30.970 49.620 31.390 50.285 ;
        RECT 31.700 49.955 32.050 50.285 ;
        RECT 32.285 49.770 32.460 50.485 ;
        RECT 32.715 50.285 32.885 50.765 ;
        RECT 33.740 50.675 33.910 50.865 ;
        RECT 34.190 50.855 34.600 51.025 ;
        RECT 32.630 49.955 32.885 50.285 ;
        RECT 33.110 49.955 33.440 50.575 ;
        RECT 33.740 50.505 34.260 50.675 ;
        RECT 33.610 49.955 33.900 50.335 ;
        RECT 34.090 49.785 34.260 50.505 ;
        RECT 28.610 49.260 28.945 49.520 ;
        RECT 29.615 49.445 29.785 49.615 ;
        RECT 29.115 49.045 29.445 49.445 ;
        RECT 29.615 49.275 31.230 49.445 ;
        RECT 31.775 49.045 32.105 49.765 ;
        RECT 32.285 49.215 32.545 49.770 ;
        RECT 33.380 49.615 34.260 49.785 ;
        RECT 34.430 49.830 34.600 50.855 ;
        RECT 34.775 50.965 34.945 51.215 ;
        RECT 35.115 51.135 35.365 51.595 ;
        RECT 35.535 50.965 35.715 51.425 ;
        RECT 34.775 50.795 35.715 50.965 ;
        RECT 34.800 50.315 35.280 50.615 ;
        RECT 34.430 49.660 34.780 49.830 ;
        RECT 35.020 49.725 35.280 50.315 ;
        RECT 35.480 49.725 35.740 50.615 ;
        RECT 36.430 50.455 36.750 51.595 ;
        RECT 36.930 50.285 37.125 51.335 ;
        RECT 37.305 50.745 37.635 51.425 ;
        RECT 37.835 50.795 38.090 51.595 ;
        RECT 37.305 50.465 37.655 50.745 ;
        RECT 36.490 50.235 36.750 50.285 ;
        RECT 36.485 50.065 36.750 50.235 ;
        RECT 36.490 49.955 36.750 50.065 ;
        RECT 36.930 49.955 37.315 50.285 ;
        RECT 37.485 50.085 37.655 50.465 ;
        RECT 37.845 50.255 38.090 50.615 ;
        RECT 38.285 50.540 38.590 51.325 ;
        RECT 38.770 51.125 39.455 51.595 ;
        RECT 38.765 50.605 39.460 50.915 ;
        RECT 38.285 50.405 38.495 50.540 ;
        RECT 39.635 50.435 39.920 51.380 ;
        RECT 40.095 51.145 40.425 51.595 ;
        RECT 40.595 50.975 40.765 51.405 ;
        RECT 37.485 49.915 38.005 50.085 ;
        RECT 32.715 49.045 33.145 49.490 ;
        RECT 33.380 49.215 33.550 49.615 ;
        RECT 33.720 49.045 34.440 49.445 ;
        RECT 34.610 49.215 34.780 49.660 ;
        RECT 36.430 49.575 37.645 49.745 ;
        RECT 35.355 49.045 35.755 49.555 ;
        RECT 36.430 49.225 36.720 49.575 ;
        RECT 36.915 49.045 37.245 49.405 ;
        RECT 37.415 49.270 37.645 49.575 ;
        RECT 37.835 49.555 38.005 49.915 ;
        RECT 38.285 49.735 38.460 50.405 ;
        RECT 39.060 50.285 39.920 50.435 ;
        RECT 38.635 50.265 39.920 50.285 ;
        RECT 40.090 50.745 40.765 50.975 ;
        RECT 41.115 50.975 41.285 51.405 ;
        RECT 41.455 51.145 41.785 51.595 ;
        RECT 41.115 50.745 41.790 50.975 ;
        RECT 38.635 49.905 39.620 50.265 ;
        RECT 40.090 50.095 40.325 50.745 ;
        RECT 37.835 49.385 38.035 49.555 ;
        RECT 37.835 49.350 38.005 49.385 ;
        RECT 38.285 49.215 38.525 49.735 ;
        RECT 39.450 49.570 39.620 49.905 ;
        RECT 39.790 49.765 40.325 50.095 ;
        RECT 40.105 49.615 40.325 49.765 ;
        RECT 40.495 49.725 40.795 50.575 ;
        RECT 41.085 49.725 41.385 50.575 ;
        RECT 41.555 50.095 41.790 50.745 ;
        RECT 41.960 50.435 42.245 51.380 ;
        RECT 42.425 51.125 43.110 51.595 ;
        RECT 42.420 50.605 43.115 50.915 ;
        RECT 43.290 50.540 43.595 51.325 ;
        RECT 41.960 50.285 42.820 50.435 ;
        RECT 41.960 50.265 43.245 50.285 ;
        RECT 41.555 49.765 42.090 50.095 ;
        RECT 42.260 49.905 43.245 50.265 ;
        RECT 41.555 49.615 41.775 49.765 ;
        RECT 38.695 49.045 39.090 49.540 ;
        RECT 39.450 49.375 39.825 49.570 ;
        RECT 39.655 49.230 39.825 49.375 ;
        RECT 40.105 49.240 40.345 49.615 ;
        RECT 40.515 49.045 40.850 49.550 ;
        RECT 41.030 49.045 41.365 49.550 ;
        RECT 41.535 49.240 41.775 49.615 ;
        RECT 42.260 49.570 42.430 49.905 ;
        RECT 43.420 49.735 43.595 50.540 ;
        RECT 44.245 50.430 44.535 51.595 ;
        RECT 44.710 51.205 45.045 51.425 ;
        RECT 46.050 51.215 46.405 51.595 ;
        RECT 44.710 50.585 44.965 51.205 ;
        RECT 45.215 51.045 45.445 51.085 ;
        RECT 46.575 51.045 46.825 51.425 ;
        RECT 45.215 50.845 46.825 51.045 ;
        RECT 45.215 50.755 45.400 50.845 ;
        RECT 45.990 50.835 46.825 50.845 ;
        RECT 47.075 50.815 47.325 51.595 ;
        RECT 47.495 50.745 47.755 51.425 ;
        RECT 45.555 50.645 45.885 50.675 ;
        RECT 45.555 50.585 47.355 50.645 ;
        RECT 44.710 50.475 47.415 50.585 ;
        RECT 44.710 50.415 45.885 50.475 ;
        RECT 47.215 50.440 47.415 50.475 ;
        RECT 44.705 50.035 45.195 50.235 ;
        RECT 45.385 50.035 45.860 50.245 ;
        RECT 42.055 49.375 42.430 49.570 ;
        RECT 42.055 49.230 42.225 49.375 ;
        RECT 42.790 49.045 43.185 49.540 ;
        RECT 43.355 49.215 43.595 49.735 ;
        RECT 44.245 49.045 44.535 49.770 ;
        RECT 44.710 49.045 45.165 49.810 ;
        RECT 45.640 49.635 45.860 50.035 ;
        RECT 46.105 50.035 46.435 50.245 ;
        RECT 46.105 49.635 46.315 50.035 ;
        RECT 46.605 50.000 47.015 50.305 ;
        RECT 47.245 49.865 47.415 50.440 ;
        RECT 47.145 49.745 47.415 49.865 ;
        RECT 46.570 49.700 47.415 49.745 ;
        RECT 46.570 49.575 47.325 49.700 ;
        RECT 46.570 49.425 46.740 49.575 ;
        RECT 47.585 49.555 47.755 50.745 ;
        RECT 47.925 50.455 48.185 51.595 ;
        RECT 48.355 50.445 48.685 51.425 ;
        RECT 48.855 50.455 49.135 51.595 ;
        RECT 49.315 51.255 50.485 51.425 ;
        RECT 49.315 50.585 49.645 51.255 ;
        RECT 50.155 51.215 50.485 51.255 ;
        RECT 50.655 51.215 51.030 51.595 ;
        RECT 49.815 51.045 50.045 51.085 ;
        RECT 49.815 50.995 50.430 51.045 ;
        RECT 51.175 50.995 51.345 51.125 ;
        RECT 49.815 50.795 51.345 50.995 ;
        RECT 51.580 50.815 51.845 51.595 ;
        RECT 52.565 51.135 52.780 51.595 ;
        RECT 52.950 50.965 53.280 51.425 ;
        RECT 52.110 50.795 53.280 50.965 ;
        RECT 53.450 50.795 53.700 51.595 ;
        RECT 54.815 50.795 54.985 51.595 ;
        RECT 49.815 50.755 50.695 50.795 ;
        RECT 50.835 50.585 51.895 50.625 ;
        RECT 49.315 50.455 51.895 50.585 ;
        RECT 47.945 50.035 48.280 50.285 ;
        RECT 48.450 49.845 48.620 50.445 ;
        RECT 49.315 50.405 51.060 50.455 ;
        RECT 48.790 50.015 49.125 50.285 ;
        RECT 47.525 49.545 47.755 49.555 ;
        RECT 45.440 49.215 46.740 49.425 ;
        RECT 46.995 49.045 47.325 49.405 ;
        RECT 47.495 49.215 47.755 49.545 ;
        RECT 47.925 49.215 48.620 49.845 ;
        RECT 48.825 49.045 49.135 49.845 ;
        RECT 49.345 49.725 49.795 50.235 ;
        RECT 49.985 50.035 50.460 50.235 ;
        RECT 50.210 49.635 50.460 50.035 ;
        RECT 50.710 50.035 51.060 50.235 ;
        RECT 50.710 49.635 50.920 50.035 ;
        RECT 51.230 49.955 51.555 50.285 ;
        RECT 51.725 49.785 51.895 50.455 ;
        RECT 51.165 49.615 51.895 49.785 ;
        RECT 49.315 49.045 49.765 49.555 ;
        RECT 51.165 49.465 51.345 49.615 ;
        RECT 50.040 49.215 51.345 49.465 ;
        RECT 52.110 49.505 52.480 50.795 ;
        RECT 53.910 50.625 54.190 50.785 ;
        RECT 52.855 50.455 54.190 50.625 ;
        RECT 55.155 50.575 55.485 51.425 ;
        RECT 55.655 50.795 55.825 51.595 ;
        RECT 55.995 50.575 56.325 51.425 ;
        RECT 56.495 50.795 56.665 51.595 ;
        RECT 56.835 50.575 57.165 51.425 ;
        RECT 57.335 50.795 57.505 51.595 ;
        RECT 57.675 50.575 58.005 51.425 ;
        RECT 58.175 50.745 58.345 51.595 ;
        RECT 58.515 50.575 58.845 51.425 ;
        RECT 59.015 50.745 59.185 51.595 ;
        RECT 59.355 50.575 59.685 51.425 ;
        RECT 52.855 50.285 53.025 50.455 ;
        RECT 52.650 50.035 53.025 50.285 ;
        RECT 54.365 50.405 58.005 50.575 ;
        RECT 58.175 50.405 59.685 50.575 ;
        RECT 59.875 50.505 60.205 51.425 ;
        RECT 53.195 50.035 53.670 50.275 ;
        RECT 53.840 50.035 54.190 50.275 ;
        RECT 52.855 49.865 53.025 50.035 ;
        RECT 54.365 49.865 54.750 50.405 ;
        RECT 58.175 50.235 58.345 50.405 ;
        RECT 59.875 50.235 60.045 50.505 ;
        RECT 60.375 50.405 60.545 51.595 ;
        RECT 60.815 50.785 61.110 51.595 ;
        RECT 61.290 50.285 61.535 51.425 ;
        RECT 61.710 50.785 61.970 51.595 ;
        RECT 62.570 51.590 68.845 51.595 ;
        RECT 62.150 50.285 62.400 51.420 ;
        RECT 62.570 50.795 62.830 51.590 ;
        RECT 63.000 50.695 63.260 51.420 ;
        RECT 63.430 50.865 63.690 51.590 ;
        RECT 63.860 50.695 64.120 51.420 ;
        RECT 64.290 50.865 64.550 51.590 ;
        RECT 64.720 50.695 64.980 51.420 ;
        RECT 65.150 50.865 65.410 51.590 ;
        RECT 65.580 50.695 65.840 51.420 ;
        RECT 66.010 50.865 66.255 51.590 ;
        RECT 66.425 50.695 66.685 51.420 ;
        RECT 66.870 50.865 67.115 51.590 ;
        RECT 67.285 50.695 67.545 51.420 ;
        RECT 67.730 50.865 67.975 51.590 ;
        RECT 68.145 50.695 68.405 51.420 ;
        RECT 68.590 50.865 68.845 51.590 ;
        RECT 63.000 50.680 68.405 50.695 ;
        RECT 69.015 50.680 69.305 51.420 ;
        RECT 69.475 50.850 69.745 51.595 ;
        RECT 63.000 50.455 69.745 50.680 ;
        RECT 54.960 50.035 58.345 50.235 ;
        RECT 58.515 50.035 60.045 50.235 ;
        RECT 60.215 50.035 60.635 50.235 ;
        RECT 58.175 49.865 58.345 50.035 ;
        RECT 59.875 49.865 60.045 50.035 ;
        RECT 52.855 49.695 54.190 49.865 ;
        RECT 54.365 49.695 58.005 49.865 ;
        RECT 58.175 49.695 59.685 49.865 ;
        RECT 51.525 49.045 51.855 49.445 ;
        RECT 52.110 49.215 52.860 49.505 ;
        RECT 53.370 49.045 53.700 49.505 ;
        RECT 53.920 49.485 54.190 49.695 ;
        RECT 54.815 49.045 54.985 49.525 ;
        RECT 55.155 49.220 55.485 49.695 ;
        RECT 55.655 49.045 55.825 49.525 ;
        RECT 55.995 49.220 56.325 49.695 ;
        RECT 56.495 49.045 56.665 49.525 ;
        RECT 56.835 49.220 57.165 49.695 ;
        RECT 57.335 49.045 57.505 49.525 ;
        RECT 57.675 49.220 58.005 49.695 ;
        RECT 58.175 49.045 58.345 49.525 ;
        RECT 58.515 49.220 58.845 49.695 ;
        RECT 59.015 49.045 59.185 49.525 ;
        RECT 59.355 49.220 59.685 49.695 ;
        RECT 59.875 49.220 60.205 49.865 ;
        RECT 60.375 49.045 60.545 49.865 ;
        RECT 60.805 49.725 61.120 50.285 ;
        RECT 61.290 50.035 68.410 50.285 ;
        RECT 60.805 49.045 61.110 49.555 ;
        RECT 61.290 49.225 61.540 50.035 ;
        RECT 61.710 49.045 61.970 49.570 ;
        RECT 62.150 49.225 62.400 50.035 ;
        RECT 68.580 49.865 69.745 50.455 ;
        RECT 70.005 50.430 70.295 51.595 ;
        RECT 70.465 50.745 70.725 51.425 ;
        RECT 70.895 50.815 71.145 51.595 ;
        RECT 71.395 51.045 71.645 51.425 ;
        RECT 71.815 51.215 72.170 51.595 ;
        RECT 73.175 51.205 73.510 51.425 ;
        RECT 72.775 51.045 73.005 51.085 ;
        RECT 71.395 50.845 73.005 51.045 ;
        RECT 71.395 50.835 72.230 50.845 ;
        RECT 72.820 50.755 73.005 50.845 ;
        RECT 63.000 49.695 69.745 49.865 ;
        RECT 62.570 49.045 62.830 49.605 ;
        RECT 63.000 49.240 63.260 49.695 ;
        RECT 63.430 49.045 63.690 49.525 ;
        RECT 63.860 49.240 64.120 49.695 ;
        RECT 64.290 49.045 64.550 49.525 ;
        RECT 64.720 49.240 64.980 49.695 ;
        RECT 65.150 49.045 65.395 49.525 ;
        RECT 65.565 49.240 65.840 49.695 ;
        RECT 66.010 49.045 66.255 49.525 ;
        RECT 66.425 49.240 66.685 49.695 ;
        RECT 66.865 49.045 67.115 49.525 ;
        RECT 67.285 49.240 67.545 49.695 ;
        RECT 67.725 49.045 67.975 49.525 ;
        RECT 68.145 49.240 68.405 49.695 ;
        RECT 68.585 49.045 68.845 49.525 ;
        RECT 69.015 49.240 69.275 49.695 ;
        RECT 69.445 49.045 69.745 49.525 ;
        RECT 70.005 49.045 70.295 49.770 ;
        RECT 70.465 49.555 70.635 50.745 ;
        RECT 72.335 50.645 72.665 50.675 ;
        RECT 70.865 50.585 72.665 50.645 ;
        RECT 73.255 50.585 73.510 51.205 ;
        RECT 70.805 50.475 73.510 50.585 ;
        RECT 73.775 50.665 73.945 51.425 ;
        RECT 74.160 50.835 74.490 51.595 ;
        RECT 73.775 50.495 74.490 50.665 ;
        RECT 74.660 50.520 74.915 51.425 ;
        RECT 70.805 50.440 71.005 50.475 ;
        RECT 70.805 49.865 70.975 50.440 ;
        RECT 72.335 50.415 73.510 50.475 ;
        RECT 71.205 50.000 71.615 50.305 ;
        RECT 71.785 50.035 72.115 50.245 ;
        RECT 70.805 49.745 71.075 49.865 ;
        RECT 70.805 49.700 71.650 49.745 ;
        RECT 70.895 49.575 71.650 49.700 ;
        RECT 71.905 49.635 72.115 50.035 ;
        RECT 72.360 50.035 72.835 50.245 ;
        RECT 73.025 50.035 73.515 50.235 ;
        RECT 72.360 49.635 72.580 50.035 ;
        RECT 73.685 49.945 74.040 50.315 ;
        RECT 74.320 50.285 74.490 50.495 ;
        RECT 74.320 49.955 74.575 50.285 ;
        RECT 70.465 49.545 70.695 49.555 ;
        RECT 70.465 49.215 70.725 49.545 ;
        RECT 71.480 49.425 71.650 49.575 ;
        RECT 70.895 49.045 71.225 49.405 ;
        RECT 71.480 49.215 72.780 49.425 ;
        RECT 73.055 49.045 73.510 49.810 ;
        RECT 74.320 49.765 74.490 49.955 ;
        RECT 74.745 49.790 74.915 50.520 ;
        RECT 75.090 50.445 75.350 51.595 ;
        RECT 75.525 50.505 76.735 51.595 ;
        RECT 75.525 49.965 76.045 50.505 ;
        RECT 73.775 49.595 74.490 49.765 ;
        RECT 73.775 49.215 73.945 49.595 ;
        RECT 74.160 49.045 74.490 49.425 ;
        RECT 74.660 49.215 74.915 49.790 ;
        RECT 75.090 49.045 75.350 49.885 ;
        RECT 76.215 49.795 76.735 50.335 ;
        RECT 75.525 49.045 76.735 49.795 ;
        RECT 5.520 48.875 76.820 49.045 ;
        RECT 5.605 48.125 6.815 48.875 ;
        RECT 7.075 48.325 7.245 48.705 ;
        RECT 7.425 48.495 7.755 48.875 ;
        RECT 7.075 48.155 7.740 48.325 ;
        RECT 7.935 48.200 8.195 48.705 ;
        RECT 5.605 47.585 6.125 48.125 ;
        RECT 6.295 47.415 6.815 47.955 ;
        RECT 7.005 47.605 7.345 47.975 ;
        RECT 7.570 47.900 7.740 48.155 ;
        RECT 7.570 47.570 7.845 47.900 ;
        RECT 7.570 47.425 7.740 47.570 ;
        RECT 5.605 46.325 6.815 47.415 ;
        RECT 7.065 47.255 7.740 47.425 ;
        RECT 8.015 47.400 8.195 48.200 ;
        RECT 9.290 48.225 9.560 48.435 ;
        RECT 9.780 48.415 10.110 48.875 ;
        RECT 10.620 48.415 11.370 48.705 ;
        RECT 9.290 48.055 10.625 48.225 ;
        RECT 10.455 47.885 10.625 48.055 ;
        RECT 9.290 47.645 9.640 47.885 ;
        RECT 9.810 47.645 10.285 47.885 ;
        RECT 10.455 47.635 10.830 47.885 ;
        RECT 10.455 47.465 10.625 47.635 ;
        RECT 7.065 46.495 7.245 47.255 ;
        RECT 7.425 46.325 7.755 47.085 ;
        RECT 7.925 46.495 8.195 47.400 ;
        RECT 9.290 47.295 10.625 47.465 ;
        RECT 9.290 47.135 9.570 47.295 ;
        RECT 11.000 47.125 11.370 48.415 ;
        RECT 11.590 48.035 11.850 48.875 ;
        RECT 12.025 48.130 12.280 48.705 ;
        RECT 12.450 48.495 12.780 48.875 ;
        RECT 12.995 48.325 13.165 48.705 ;
        RECT 12.450 48.155 13.165 48.325 ;
        RECT 13.425 48.200 13.685 48.705 ;
        RECT 13.865 48.495 14.195 48.875 ;
        RECT 14.375 48.325 14.545 48.705 ;
        RECT 9.780 46.325 10.030 47.125 ;
        RECT 10.200 46.955 11.370 47.125 ;
        RECT 10.200 46.495 10.530 46.955 ;
        RECT 10.700 46.325 10.915 46.785 ;
        RECT 11.590 46.325 11.850 47.475 ;
        RECT 12.025 47.400 12.195 48.130 ;
        RECT 12.450 47.965 12.620 48.155 ;
        RECT 12.365 47.635 12.620 47.965 ;
        RECT 12.450 47.425 12.620 47.635 ;
        RECT 12.900 47.605 13.255 47.975 ;
        RECT 12.025 46.495 12.280 47.400 ;
        RECT 12.450 47.255 13.165 47.425 ;
        RECT 12.450 46.325 12.780 47.085 ;
        RECT 12.995 46.495 13.165 47.255 ;
        RECT 13.425 47.400 13.595 48.200 ;
        RECT 13.880 48.155 14.545 48.325 ;
        RECT 14.895 48.325 15.065 48.705 ;
        RECT 15.245 48.495 15.575 48.875 ;
        RECT 14.895 48.155 15.560 48.325 ;
        RECT 15.755 48.200 16.015 48.705 ;
        RECT 13.880 47.900 14.050 48.155 ;
        RECT 13.765 47.570 14.050 47.900 ;
        RECT 14.285 47.605 14.615 47.975 ;
        RECT 14.825 47.605 15.155 47.975 ;
        RECT 15.390 47.900 15.560 48.155 ;
        RECT 13.880 47.425 14.050 47.570 ;
        RECT 15.390 47.570 15.675 47.900 ;
        RECT 15.390 47.425 15.560 47.570 ;
        RECT 13.425 46.495 13.695 47.400 ;
        RECT 13.880 47.255 14.545 47.425 ;
        RECT 13.865 46.325 14.195 47.085 ;
        RECT 14.375 46.495 14.545 47.255 ;
        RECT 14.895 47.255 15.560 47.425 ;
        RECT 15.845 47.400 16.015 48.200 ;
        RECT 16.185 48.105 19.695 48.875 ;
        RECT 19.865 48.125 21.075 48.875 ;
        RECT 16.185 47.585 17.835 48.105 ;
        RECT 18.005 47.415 19.695 47.935 ;
        RECT 19.865 47.585 20.385 48.125 ;
        RECT 21.245 48.075 21.555 48.875 ;
        RECT 21.760 48.075 22.455 48.705 ;
        RECT 22.625 48.330 27.970 48.875 ;
        RECT 20.555 47.415 21.075 47.955 ;
        RECT 21.255 47.635 21.590 47.905 ;
        RECT 21.760 47.475 21.930 48.075 ;
        RECT 22.100 47.635 22.435 47.885 ;
        RECT 24.210 47.500 24.550 48.330 ;
        RECT 28.145 48.105 30.735 48.875 ;
        RECT 31.365 48.150 31.655 48.875 ;
        RECT 31.910 48.375 32.405 48.705 ;
        RECT 14.895 46.495 15.065 47.255 ;
        RECT 15.245 46.325 15.575 47.085 ;
        RECT 15.745 46.495 16.015 47.400 ;
        RECT 16.185 46.325 19.695 47.415 ;
        RECT 19.865 46.325 21.075 47.415 ;
        RECT 21.245 46.325 21.525 47.465 ;
        RECT 21.695 46.495 22.025 47.475 ;
        RECT 22.195 46.325 22.455 47.465 ;
        RECT 26.030 46.760 26.380 48.010 ;
        RECT 28.145 47.585 29.355 48.105 ;
        RECT 29.525 47.415 30.735 47.935 ;
        RECT 22.625 46.325 27.970 46.760 ;
        RECT 28.145 46.325 30.735 47.415 ;
        RECT 31.365 46.325 31.655 47.490 ;
        RECT 31.825 46.885 32.065 48.195 ;
        RECT 32.235 47.465 32.405 48.375 ;
        RECT 32.625 47.635 32.975 48.600 ;
        RECT 33.155 47.635 33.455 48.605 ;
        RECT 33.635 47.635 33.915 48.605 ;
        RECT 34.095 48.075 34.365 48.875 ;
        RECT 34.535 48.155 34.875 48.665 ;
        RECT 35.070 48.485 35.400 48.875 ;
        RECT 35.570 48.315 35.795 48.695 ;
        RECT 34.110 47.635 34.440 47.885 ;
        RECT 34.110 47.465 34.425 47.635 ;
        RECT 32.235 47.295 34.425 47.465 ;
        RECT 31.830 46.325 32.165 46.705 ;
        RECT 32.335 46.495 32.585 47.295 ;
        RECT 32.805 46.325 33.135 47.045 ;
        RECT 33.320 46.495 33.570 47.295 ;
        RECT 34.035 46.325 34.365 47.125 ;
        RECT 34.615 46.755 34.875 48.155 ;
        RECT 35.055 47.635 35.295 48.285 ;
        RECT 35.465 48.135 35.795 48.315 ;
        RECT 35.465 47.465 35.640 48.135 ;
        RECT 35.995 47.965 36.225 48.585 ;
        RECT 36.405 48.145 36.705 48.875 ;
        RECT 36.885 48.105 38.555 48.875 ;
        RECT 35.810 47.635 36.225 47.965 ;
        RECT 36.405 47.635 36.700 47.965 ;
        RECT 36.885 47.585 37.635 48.105 ;
        RECT 38.725 48.075 39.420 48.705 ;
        RECT 39.625 48.075 39.935 48.875 ;
        RECT 40.105 48.200 40.365 48.705 ;
        RECT 40.545 48.495 40.875 48.875 ;
        RECT 41.055 48.325 41.225 48.705 ;
        RECT 39.245 48.025 39.420 48.075 ;
        RECT 34.535 46.495 34.875 46.755 ;
        RECT 35.055 47.275 35.640 47.465 ;
        RECT 35.055 46.505 35.330 47.275 ;
        RECT 35.810 47.105 36.705 47.435 ;
        RECT 37.805 47.415 38.555 47.935 ;
        RECT 38.745 47.635 39.080 47.885 ;
        RECT 39.250 47.475 39.420 48.025 ;
        RECT 39.590 47.635 39.925 47.905 ;
        RECT 35.500 46.935 36.705 47.105 ;
        RECT 35.500 46.505 35.830 46.935 ;
        RECT 36.000 46.325 36.195 46.765 ;
        RECT 36.375 46.505 36.705 46.935 ;
        RECT 36.885 46.325 38.555 47.415 ;
        RECT 38.725 46.325 38.985 47.465 ;
        RECT 39.155 46.495 39.485 47.475 ;
        RECT 39.655 46.325 39.935 47.465 ;
        RECT 40.105 47.400 40.275 48.200 ;
        RECT 40.560 48.155 41.225 48.325 ;
        RECT 41.485 48.200 41.745 48.705 ;
        RECT 41.925 48.495 42.255 48.875 ;
        RECT 42.435 48.325 42.605 48.705 ;
        RECT 40.560 47.900 40.730 48.155 ;
        RECT 40.445 47.570 40.730 47.900 ;
        RECT 40.965 47.605 41.295 47.975 ;
        RECT 40.560 47.425 40.730 47.570 ;
        RECT 40.105 46.495 40.375 47.400 ;
        RECT 40.560 47.255 41.225 47.425 ;
        RECT 40.545 46.325 40.875 47.085 ;
        RECT 41.055 46.495 41.225 47.255 ;
        RECT 41.485 47.400 41.655 48.200 ;
        RECT 41.940 48.155 42.605 48.325 ;
        RECT 42.865 48.200 43.125 48.705 ;
        RECT 43.305 48.495 43.635 48.875 ;
        RECT 43.815 48.325 43.985 48.705 ;
        RECT 41.940 47.900 42.110 48.155 ;
        RECT 41.825 47.570 42.110 47.900 ;
        RECT 42.345 47.605 42.675 47.975 ;
        RECT 41.940 47.425 42.110 47.570 ;
        RECT 41.485 46.495 41.755 47.400 ;
        RECT 41.940 47.255 42.605 47.425 ;
        RECT 41.925 46.325 42.255 47.085 ;
        RECT 42.435 46.495 42.605 47.255 ;
        RECT 42.865 47.400 43.045 48.200 ;
        RECT 43.320 48.155 43.985 48.325 ;
        RECT 43.320 47.900 43.490 48.155 ;
        RECT 43.215 47.570 43.490 47.900 ;
        RECT 43.715 47.605 44.055 47.975 ;
        RECT 43.320 47.425 43.490 47.570 ;
        RECT 42.865 46.495 43.135 47.400 ;
        RECT 43.320 47.255 43.995 47.425 ;
        RECT 43.305 46.325 43.635 47.085 ;
        RECT 43.815 46.495 43.995 47.255 ;
        RECT 44.260 46.505 44.540 48.695 ;
        RECT 44.740 48.505 45.470 48.875 ;
        RECT 46.050 48.335 46.480 48.695 ;
        RECT 44.740 48.145 46.480 48.335 ;
        RECT 44.740 47.635 45.000 48.145 ;
        RECT 44.730 46.325 45.015 47.465 ;
        RECT 45.210 47.345 45.470 47.965 ;
        RECT 45.665 47.345 46.090 47.965 ;
        RECT 46.260 47.915 46.480 48.145 ;
        RECT 46.650 48.095 46.895 48.875 ;
        RECT 46.260 47.615 46.805 47.915 ;
        RECT 47.095 47.795 47.325 48.695 ;
        RECT 45.280 46.975 46.305 47.175 ;
        RECT 45.280 46.505 45.450 46.975 ;
        RECT 45.625 46.325 45.955 46.805 ;
        RECT 46.125 46.505 46.305 46.975 ;
        RECT 46.475 46.505 46.805 47.615 ;
        RECT 46.985 47.115 47.325 47.795 ;
        RECT 47.505 47.295 47.735 48.635 ;
        RECT 47.925 48.075 48.235 48.875 ;
        RECT 48.440 48.075 49.135 48.705 ;
        RECT 49.315 48.365 49.765 48.875 ;
        RECT 50.040 48.455 51.345 48.705 ;
        RECT 51.525 48.475 51.855 48.875 ;
        RECT 51.165 48.305 51.345 48.455 ;
        RECT 47.935 47.635 48.270 47.905 ;
        RECT 48.440 47.475 48.610 48.075 ;
        RECT 48.780 47.635 49.115 47.885 ;
        RECT 49.345 47.685 49.795 48.195 ;
        RECT 50.210 47.885 50.460 48.285 ;
        RECT 49.985 47.685 50.460 47.885 ;
        RECT 50.710 47.885 50.920 48.285 ;
        RECT 51.165 48.135 51.895 48.305 ;
        RECT 50.710 47.685 51.060 47.885 ;
        RECT 51.230 47.635 51.555 47.965 ;
        RECT 46.985 46.915 47.735 47.115 ;
        RECT 46.975 46.325 47.325 46.735 ;
        RECT 47.495 46.525 47.735 46.915 ;
        RECT 47.925 46.325 48.205 47.465 ;
        RECT 48.375 46.495 48.705 47.475 ;
        RECT 49.315 47.465 51.060 47.515 ;
        RECT 51.725 47.465 51.895 48.135 ;
        RECT 48.875 46.325 49.135 47.465 ;
        RECT 49.315 47.335 51.895 47.465 ;
        RECT 49.315 46.665 49.645 47.335 ;
        RECT 50.835 47.295 51.895 47.335 ;
        RECT 52.525 48.150 52.785 48.705 ;
        RECT 52.955 48.430 53.385 48.875 ;
        RECT 53.620 48.305 53.790 48.705 ;
        RECT 53.960 48.475 54.680 48.875 ;
        RECT 52.525 47.435 52.700 48.150 ;
        RECT 53.620 48.135 54.500 48.305 ;
        RECT 54.850 48.260 55.020 48.705 ;
        RECT 55.595 48.365 55.995 48.875 ;
        RECT 52.870 47.635 53.125 47.965 ;
        RECT 49.815 47.125 50.695 47.165 ;
        RECT 49.815 46.925 51.345 47.125 ;
        RECT 49.815 46.875 50.430 46.925 ;
        RECT 49.815 46.835 50.045 46.875 ;
        RECT 51.175 46.795 51.345 46.925 ;
        RECT 50.155 46.665 50.485 46.705 ;
        RECT 49.315 46.495 50.485 46.665 ;
        RECT 50.655 46.325 51.030 46.705 ;
        RECT 51.580 46.325 51.845 47.105 ;
        RECT 52.525 46.495 52.785 47.435 ;
        RECT 52.955 47.155 53.125 47.635 ;
        RECT 53.350 47.345 53.680 47.965 ;
        RECT 53.850 47.585 54.140 47.965 ;
        RECT 54.330 47.415 54.500 48.135 ;
        RECT 53.980 47.245 54.500 47.415 ;
        RECT 54.670 48.090 55.020 48.260 ;
        RECT 52.955 46.985 53.715 47.155 ;
        RECT 53.980 47.055 54.150 47.245 ;
        RECT 54.670 47.065 54.840 48.090 ;
        RECT 55.260 47.605 55.520 48.195 ;
        RECT 55.040 47.305 55.520 47.605 ;
        RECT 55.720 47.305 55.980 48.195 ;
        RECT 57.125 48.150 57.415 48.875 ;
        RECT 57.645 48.395 57.925 48.875 ;
        RECT 58.095 48.225 58.355 48.615 ;
        RECT 58.530 48.395 58.785 48.875 ;
        RECT 58.955 48.225 59.250 48.615 ;
        RECT 59.430 48.395 59.705 48.875 ;
        RECT 59.875 48.375 60.175 48.705 ;
        RECT 57.600 48.055 59.250 48.225 ;
        RECT 57.600 47.545 58.005 48.055 ;
        RECT 58.175 47.715 59.315 47.885 ;
        RECT 53.545 46.760 53.715 46.985 ;
        RECT 54.430 46.895 54.840 47.065 ;
        RECT 55.015 46.955 55.955 47.125 ;
        RECT 54.430 46.760 54.685 46.895 ;
        RECT 52.955 46.325 53.285 46.725 ;
        RECT 53.545 46.590 54.685 46.760 ;
        RECT 55.015 46.705 55.185 46.955 ;
        RECT 54.430 46.495 54.685 46.590 ;
        RECT 54.855 46.535 55.185 46.705 ;
        RECT 55.355 46.325 55.605 46.785 ;
        RECT 55.775 46.495 55.955 46.955 ;
        RECT 57.125 46.325 57.415 47.490 ;
        RECT 57.600 47.375 58.355 47.545 ;
        RECT 57.640 46.325 57.925 47.195 ;
        RECT 58.095 47.125 58.355 47.375 ;
        RECT 59.145 47.465 59.315 47.715 ;
        RECT 59.485 47.635 59.835 48.205 ;
        RECT 60.005 47.465 60.175 48.375 ;
        RECT 60.345 48.365 60.650 48.875 ;
        RECT 60.345 47.635 60.660 48.195 ;
        RECT 60.830 47.885 61.080 48.695 ;
        RECT 61.250 48.350 61.510 48.875 ;
        RECT 61.690 47.885 61.940 48.695 ;
        RECT 62.110 48.315 62.370 48.875 ;
        RECT 62.540 48.225 62.800 48.680 ;
        RECT 62.970 48.395 63.230 48.875 ;
        RECT 63.400 48.225 63.660 48.680 ;
        RECT 63.830 48.395 64.090 48.875 ;
        RECT 64.260 48.225 64.520 48.680 ;
        RECT 64.690 48.395 64.935 48.875 ;
        RECT 65.105 48.225 65.380 48.680 ;
        RECT 65.550 48.395 65.795 48.875 ;
        RECT 65.965 48.225 66.225 48.680 ;
        RECT 66.405 48.395 66.655 48.875 ;
        RECT 66.825 48.225 67.085 48.680 ;
        RECT 67.265 48.395 67.515 48.875 ;
        RECT 67.685 48.225 67.945 48.680 ;
        RECT 68.125 48.395 68.385 48.875 ;
        RECT 68.555 48.225 68.815 48.680 ;
        RECT 68.985 48.395 69.285 48.875 ;
        RECT 70.465 48.265 70.815 48.705 ;
        RECT 70.985 48.435 71.155 48.875 ;
        RECT 71.325 48.495 72.520 48.705 ;
        RECT 71.325 48.265 71.575 48.495 ;
        RECT 62.540 48.055 69.285 48.225 ;
        RECT 70.465 48.055 71.575 48.265 ;
        RECT 71.745 48.155 72.075 48.325 ;
        RECT 71.745 48.055 72.070 48.155 ;
        RECT 72.245 48.055 72.520 48.495 ;
        RECT 72.755 48.135 73.085 48.875 ;
        RECT 73.255 48.120 73.490 48.450 ;
        RECT 60.830 47.635 67.950 47.885 ;
        RECT 59.145 47.295 60.175 47.465 ;
        RECT 58.095 46.955 59.215 47.125 ;
        RECT 58.095 46.495 58.355 46.955 ;
        RECT 58.530 46.325 58.785 46.785 ;
        RECT 58.955 46.495 59.215 46.955 ;
        RECT 59.385 46.325 59.695 47.125 ;
        RECT 59.865 46.495 60.175 47.295 ;
        RECT 60.355 46.325 60.650 47.135 ;
        RECT 60.830 46.495 61.075 47.635 ;
        RECT 61.250 46.325 61.510 47.135 ;
        RECT 61.690 46.500 61.940 47.635 ;
        RECT 68.120 47.465 69.285 48.055 ;
        RECT 70.465 47.685 71.610 47.885 ;
        RECT 70.985 47.465 71.155 47.515 ;
        RECT 62.540 47.240 69.285 47.465 ;
        RECT 62.540 47.225 67.945 47.240 ;
        RECT 62.110 46.330 62.370 47.125 ;
        RECT 62.540 46.500 62.800 47.225 ;
        RECT 62.970 46.330 63.230 47.055 ;
        RECT 63.400 46.500 63.660 47.225 ;
        RECT 63.830 46.330 64.090 47.055 ;
        RECT 64.260 46.500 64.520 47.225 ;
        RECT 64.690 46.330 64.950 47.055 ;
        RECT 65.120 46.500 65.380 47.225 ;
        RECT 65.550 46.330 65.795 47.055 ;
        RECT 65.965 46.500 66.225 47.225 ;
        RECT 66.410 46.330 66.655 47.055 ;
        RECT 66.825 46.500 67.085 47.225 ;
        RECT 67.270 46.330 67.515 47.055 ;
        RECT 67.685 46.500 67.945 47.225 ;
        RECT 68.130 46.330 68.385 47.055 ;
        RECT 68.555 46.500 68.845 47.240 ;
        RECT 62.110 46.325 68.385 46.330 ;
        RECT 69.015 46.325 69.285 47.070 ;
        RECT 70.465 46.325 70.795 47.465 ;
        RECT 70.965 47.125 71.240 47.465 ;
        RECT 71.420 47.305 71.610 47.685 ;
        RECT 71.790 47.125 72.070 48.055 ;
        RECT 72.240 47.465 72.570 47.885 ;
        RECT 72.800 47.635 73.145 47.965 ;
        RECT 73.320 47.465 73.490 48.120 ;
        RECT 73.685 48.105 75.355 48.875 ;
        RECT 75.525 48.125 76.735 48.875 ;
        RECT 73.685 47.585 74.435 48.105 ;
        RECT 72.240 47.295 73.490 47.465 ;
        RECT 74.605 47.415 75.355 47.935 ;
        RECT 70.965 46.955 72.565 47.125 ;
        RECT 70.965 46.495 71.320 46.955 ;
        RECT 71.490 46.325 72.065 46.785 ;
        RECT 72.235 46.495 72.565 46.955 ;
        RECT 72.765 46.325 73.020 47.125 ;
        RECT 73.190 47.100 73.490 47.295 ;
        RECT 73.685 46.325 75.355 47.415 ;
        RECT 75.525 47.415 76.045 47.955 ;
        RECT 76.215 47.585 76.735 48.125 ;
        RECT 75.525 46.325 76.735 47.415 ;
        RECT 5.520 46.155 76.820 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 7.905 43.885 8.185 45.985 ;
        RECT 8.375 45.395 9.160 46.155 ;
        RECT 9.555 45.325 9.940 45.985 ;
        RECT 9.555 45.225 9.965 45.325 ;
        RECT 8.355 45.015 9.965 45.225 ;
        RECT 10.265 45.135 10.465 45.925 ;
        RECT 8.355 44.415 8.630 45.015 ;
        RECT 10.135 44.965 10.465 45.135 ;
        RECT 10.635 44.975 10.955 46.155 ;
        RECT 11.125 45.720 16.470 46.155 ;
        RECT 10.135 44.845 10.315 44.965 ;
        RECT 8.800 44.595 9.155 44.845 ;
        RECT 9.350 44.795 9.815 44.845 ;
        RECT 9.345 44.625 9.815 44.795 ;
        RECT 9.350 44.595 9.815 44.625 ;
        RECT 9.985 44.595 10.315 44.845 ;
        RECT 10.490 44.595 10.955 44.795 ;
        RECT 8.355 44.235 9.605 44.415 ;
        RECT 9.240 44.165 9.605 44.235 ;
        RECT 9.775 44.215 10.955 44.385 ;
        RECT 8.415 43.605 8.585 44.065 ;
        RECT 9.775 43.995 10.105 44.215 ;
        RECT 8.855 43.815 10.105 43.995 ;
        RECT 10.275 43.605 10.445 44.045 ;
        RECT 10.615 43.800 10.955 44.215 ;
        RECT 12.710 44.150 13.050 44.980 ;
        RECT 14.530 44.470 14.880 45.720 ;
        RECT 16.645 45.065 18.315 46.155 ;
        RECT 16.645 44.375 17.395 44.895 ;
        RECT 17.565 44.545 18.315 45.065 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 18.965 45.265 19.225 45.975 ;
        RECT 19.395 45.445 19.725 46.155 ;
        RECT 19.895 45.265 20.125 45.975 ;
        RECT 18.965 45.025 20.125 45.265 ;
        RECT 20.305 45.245 20.575 45.975 ;
        RECT 20.755 45.425 21.095 46.155 ;
        RECT 20.305 45.025 21.075 45.245 ;
        RECT 18.955 44.515 19.255 44.845 ;
        RECT 19.435 44.535 19.960 44.845 ;
        RECT 20.140 44.535 20.605 44.845 ;
        RECT 11.125 43.605 16.470 44.150 ;
        RECT 16.645 43.605 18.315 44.375 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 18.965 43.605 19.255 44.335 ;
        RECT 19.435 43.895 19.665 44.535 ;
        RECT 20.785 44.355 21.075 45.025 ;
        RECT 19.845 44.155 21.075 44.355 ;
        RECT 19.845 43.785 20.155 44.155 ;
        RECT 20.335 43.605 21.005 43.975 ;
        RECT 21.265 43.785 21.525 45.975 ;
        RECT 21.705 45.065 25.215 46.155 ;
        RECT 21.705 44.375 23.355 44.895 ;
        RECT 23.525 44.545 25.215 45.065 ;
        RECT 25.845 45.015 26.105 46.155 ;
        RECT 26.275 45.005 26.605 45.985 ;
        RECT 26.775 45.015 27.055 46.155 ;
        RECT 27.225 45.720 32.570 46.155 ;
        RECT 32.745 45.720 38.090 46.155 ;
        RECT 26.365 44.965 26.540 45.005 ;
        RECT 25.865 44.595 26.200 44.845 ;
        RECT 26.370 44.405 26.540 44.965 ;
        RECT 26.710 44.575 27.045 44.845 ;
        RECT 21.705 43.605 25.215 44.375 ;
        RECT 25.845 43.775 26.540 44.405 ;
        RECT 26.745 43.605 27.055 44.405 ;
        RECT 28.810 44.150 29.150 44.980 ;
        RECT 30.630 44.470 30.980 45.720 ;
        RECT 34.330 44.150 34.670 44.980 ;
        RECT 36.150 44.470 36.500 45.720 ;
        RECT 38.265 45.065 39.475 46.155 ;
        RECT 38.265 44.355 38.785 44.895 ;
        RECT 38.955 44.525 39.475 45.065 ;
        RECT 39.655 45.545 39.985 45.975 ;
        RECT 40.165 45.715 40.360 46.155 ;
        RECT 40.530 45.545 40.860 45.975 ;
        RECT 39.655 45.375 40.860 45.545 ;
        RECT 39.655 45.045 40.550 45.375 ;
        RECT 41.030 45.205 41.305 45.975 ;
        RECT 40.720 45.015 41.305 45.205 ;
        RECT 41.955 45.205 42.230 45.975 ;
        RECT 42.400 45.545 42.730 45.975 ;
        RECT 42.900 45.715 43.095 46.155 ;
        RECT 43.275 45.545 43.605 45.975 ;
        RECT 42.400 45.375 43.605 45.545 ;
        RECT 41.955 45.015 42.540 45.205 ;
        RECT 42.710 45.045 43.605 45.375 ;
        RECT 39.660 44.515 39.955 44.845 ;
        RECT 40.135 44.515 40.550 44.845 ;
        RECT 27.225 43.605 32.570 44.150 ;
        RECT 32.745 43.605 38.090 44.150 ;
        RECT 38.265 43.605 39.475 44.355 ;
        RECT 39.655 43.605 39.955 44.335 ;
        RECT 40.135 43.895 40.365 44.515 ;
        RECT 40.720 44.345 40.895 45.015 ;
        RECT 40.565 44.165 40.895 44.345 ;
        RECT 41.065 44.195 41.305 44.845 ;
        RECT 41.955 44.195 42.195 44.845 ;
        RECT 42.365 44.345 42.540 45.015 ;
        RECT 44.245 44.990 44.535 46.155 ;
        RECT 45.245 45.225 45.425 45.985 ;
        RECT 45.605 45.395 45.935 46.155 ;
        RECT 45.245 45.055 45.920 45.225 ;
        RECT 46.105 45.080 46.375 45.985 ;
        RECT 45.750 44.910 45.920 45.055 ;
        RECT 42.710 44.515 43.125 44.845 ;
        RECT 43.305 44.515 43.600 44.845 ;
        RECT 42.365 44.165 42.695 44.345 ;
        RECT 40.565 43.785 40.790 44.165 ;
        RECT 40.960 43.605 41.290 43.995 ;
        RECT 41.970 43.605 42.300 43.995 ;
        RECT 42.470 43.785 42.695 44.165 ;
        RECT 42.895 43.895 43.125 44.515 ;
        RECT 45.185 44.505 45.525 44.875 ;
        RECT 45.750 44.580 46.025 44.910 ;
        RECT 43.305 43.605 43.605 44.335 ;
        RECT 44.245 43.605 44.535 44.330 ;
        RECT 45.750 44.325 45.920 44.580 ;
        RECT 45.255 44.155 45.920 44.325 ;
        RECT 46.195 44.280 46.375 45.080 ;
        RECT 46.625 45.225 46.805 45.985 ;
        RECT 46.985 45.395 47.315 46.155 ;
        RECT 46.625 45.055 47.300 45.225 ;
        RECT 47.485 45.080 47.755 45.985 ;
        RECT 47.130 44.910 47.300 45.055 ;
        RECT 46.565 44.505 46.905 44.875 ;
        RECT 47.130 44.580 47.405 44.910 ;
        RECT 47.130 44.325 47.300 44.580 ;
        RECT 45.255 43.775 45.425 44.155 ;
        RECT 45.605 43.605 45.935 43.985 ;
        RECT 46.115 43.775 46.375 44.280 ;
        RECT 46.635 44.155 47.300 44.325 ;
        RECT 47.575 44.280 47.755 45.080 ;
        RECT 46.635 43.775 46.805 44.155 ;
        RECT 46.985 43.605 47.315 43.985 ;
        RECT 47.495 43.775 47.755 44.280 ;
        RECT 47.925 45.080 48.195 45.985 ;
        RECT 48.365 45.395 48.695 46.155 ;
        RECT 48.875 45.225 49.055 45.985 ;
        RECT 47.925 44.280 48.105 45.080 ;
        RECT 48.380 45.055 49.055 45.225 ;
        RECT 49.305 45.305 49.565 45.985 ;
        RECT 49.735 45.375 49.985 46.155 ;
        RECT 50.235 45.605 50.485 45.985 ;
        RECT 50.655 45.775 51.010 46.155 ;
        RECT 52.015 45.765 52.350 45.985 ;
        RECT 51.615 45.605 51.845 45.645 ;
        RECT 50.235 45.405 51.845 45.605 ;
        RECT 50.235 45.395 51.070 45.405 ;
        RECT 51.660 45.315 51.845 45.405 ;
        RECT 48.380 44.910 48.550 45.055 ;
        RECT 48.275 44.580 48.550 44.910 ;
        RECT 48.380 44.325 48.550 44.580 ;
        RECT 48.775 44.505 49.115 44.875 ;
        RECT 47.925 43.775 48.185 44.280 ;
        RECT 48.380 44.155 49.045 44.325 ;
        RECT 48.365 43.605 48.695 43.985 ;
        RECT 48.875 43.775 49.045 44.155 ;
        RECT 49.305 44.105 49.475 45.305 ;
        RECT 51.175 45.205 51.505 45.235 ;
        RECT 49.705 45.145 51.505 45.205 ;
        RECT 52.095 45.145 52.350 45.765 ;
        RECT 49.645 45.035 52.350 45.145 ;
        RECT 49.645 45.000 49.845 45.035 ;
        RECT 49.645 44.425 49.815 45.000 ;
        RECT 51.175 44.975 52.350 45.035 ;
        RECT 52.585 45.015 52.795 46.155 ;
        RECT 52.965 45.005 53.295 45.985 ;
        RECT 53.465 45.015 53.695 46.155 ;
        RECT 53.945 45.015 54.175 46.155 ;
        RECT 54.345 45.005 54.675 45.985 ;
        RECT 54.845 45.015 55.055 46.155 ;
        RECT 55.325 45.815 56.465 45.985 ;
        RECT 55.325 45.355 55.625 45.815 ;
        RECT 55.795 45.185 56.125 45.645 ;
        RECT 55.365 45.135 56.125 45.185 ;
        RECT 50.045 44.560 50.455 44.865 ;
        RECT 50.625 44.595 50.955 44.805 ;
        RECT 49.645 44.305 49.915 44.425 ;
        RECT 49.645 44.260 50.490 44.305 ;
        RECT 49.735 44.135 50.490 44.260 ;
        RECT 50.745 44.195 50.955 44.595 ;
        RECT 51.200 44.595 51.675 44.805 ;
        RECT 51.865 44.595 52.355 44.795 ;
        RECT 51.200 44.195 51.420 44.595 ;
        RECT 49.305 43.775 49.565 44.105 ;
        RECT 50.320 43.985 50.490 44.135 ;
        RECT 49.735 43.605 50.065 43.965 ;
        RECT 50.320 43.775 51.620 43.985 ;
        RECT 51.895 43.605 52.350 44.370 ;
        RECT 52.585 43.605 52.795 44.425 ;
        RECT 52.965 44.405 53.215 45.005 ;
        RECT 53.385 44.595 53.715 44.845 ;
        RECT 53.925 44.595 54.255 44.845 ;
        RECT 52.965 43.775 53.295 44.405 ;
        RECT 53.465 43.605 53.695 44.425 ;
        RECT 53.945 43.605 54.175 44.425 ;
        RECT 54.425 44.405 54.675 45.005 ;
        RECT 55.345 44.965 56.125 45.135 ;
        RECT 56.295 45.185 56.465 45.815 ;
        RECT 56.635 45.355 56.965 46.155 ;
        RECT 57.135 45.185 57.410 45.985 ;
        RECT 57.790 45.715 58.120 46.155 ;
        RECT 58.290 45.545 58.525 45.985 ;
        RECT 58.710 45.775 59.040 46.155 ;
        RECT 59.250 45.545 59.595 45.985 ;
        RECT 56.295 44.975 57.410 45.185 ;
        RECT 57.585 45.305 59.595 45.545 ;
        RECT 55.365 44.425 55.580 44.965 ;
        RECT 55.750 44.595 56.520 44.795 ;
        RECT 56.690 44.595 57.410 44.795 ;
        RECT 54.345 43.775 54.675 44.405 ;
        RECT 54.845 43.605 55.055 44.425 ;
        RECT 55.365 44.255 56.965 44.425 ;
        RECT 55.795 44.245 56.965 44.255 ;
        RECT 55.335 43.605 55.625 44.075 ;
        RECT 55.795 43.775 56.125 44.245 ;
        RECT 56.295 43.605 56.465 44.075 ;
        RECT 56.635 43.775 56.965 44.245 ;
        RECT 57.135 43.605 57.410 44.425 ;
        RECT 57.585 44.405 57.815 45.305 ;
        RECT 59.770 45.135 60.115 45.890 ;
        RECT 60.285 45.315 60.615 46.155 ;
        RECT 60.895 45.410 61.165 46.155 ;
        RECT 61.795 46.150 68.070 46.155 ;
        RECT 61.335 45.240 61.625 45.980 ;
        RECT 61.795 45.425 62.050 46.150 ;
        RECT 62.235 45.255 62.495 45.980 ;
        RECT 62.665 45.425 62.910 46.150 ;
        RECT 63.095 45.255 63.355 45.980 ;
        RECT 63.525 45.425 63.770 46.150 ;
        RECT 63.955 45.255 64.215 45.980 ;
        RECT 64.385 45.425 64.630 46.150 ;
        RECT 64.800 45.255 65.060 45.980 ;
        RECT 65.230 45.425 65.490 46.150 ;
        RECT 65.660 45.255 65.920 45.980 ;
        RECT 66.090 45.425 66.350 46.150 ;
        RECT 66.520 45.255 66.780 45.980 ;
        RECT 66.950 45.425 67.210 46.150 ;
        RECT 67.380 45.255 67.640 45.980 ;
        RECT 67.810 45.355 68.070 46.150 ;
        RECT 62.235 45.240 67.640 45.255 ;
        RECT 57.985 44.595 58.315 45.135 ;
        RECT 57.585 43.775 58.190 44.405 ;
        RECT 58.525 43.775 58.855 45.135 ;
        RECT 59.025 44.515 59.315 45.135 ;
        RECT 59.485 44.515 60.115 45.135 ;
        RECT 60.285 44.525 60.615 45.135 ;
        RECT 60.895 45.015 67.640 45.240 ;
        RECT 60.895 44.425 62.060 45.015 ;
        RECT 68.240 44.845 68.490 45.980 ;
        RECT 68.670 45.345 68.930 46.155 ;
        RECT 69.105 44.845 69.350 45.985 ;
        RECT 69.530 45.345 69.825 46.155 ;
        RECT 70.005 44.990 70.295 46.155 ;
        RECT 70.490 45.185 70.790 45.380 ;
        RECT 70.960 45.355 71.215 46.155 ;
        RECT 71.415 45.525 71.745 45.985 ;
        RECT 71.915 45.695 72.490 46.155 ;
        RECT 72.660 45.525 73.015 45.985 ;
        RECT 71.415 45.355 73.015 45.525 ;
        RECT 70.490 45.015 71.740 45.185 ;
        RECT 62.230 44.595 69.350 44.845 ;
        RECT 59.250 44.145 60.615 44.345 ;
        RECT 60.895 44.255 67.640 44.425 ;
        RECT 59.250 43.775 59.595 44.145 ;
        RECT 59.785 43.605 60.115 43.975 ;
        RECT 60.285 43.775 60.615 44.145 ;
        RECT 60.895 43.605 61.195 44.085 ;
        RECT 61.365 43.800 61.625 44.255 ;
        RECT 61.795 43.605 62.055 44.085 ;
        RECT 62.235 43.800 62.495 44.255 ;
        RECT 62.665 43.605 62.915 44.085 ;
        RECT 63.095 43.800 63.355 44.255 ;
        RECT 63.525 43.605 63.775 44.085 ;
        RECT 63.955 43.800 64.215 44.255 ;
        RECT 64.385 43.605 64.630 44.085 ;
        RECT 64.800 43.800 65.075 44.255 ;
        RECT 65.245 43.605 65.490 44.085 ;
        RECT 65.660 43.800 65.920 44.255 ;
        RECT 66.090 43.605 66.350 44.085 ;
        RECT 66.520 43.800 66.780 44.255 ;
        RECT 66.950 43.605 67.210 44.085 ;
        RECT 67.380 43.800 67.640 44.255 ;
        RECT 67.810 43.605 68.070 44.165 ;
        RECT 68.240 43.785 68.490 44.595 ;
        RECT 68.670 43.605 68.930 44.130 ;
        RECT 69.100 43.785 69.350 44.595 ;
        RECT 69.520 44.285 69.835 44.845 ;
        RECT 70.490 44.360 70.660 45.015 ;
        RECT 70.835 44.515 71.180 44.845 ;
        RECT 71.410 44.595 71.740 45.015 ;
        RECT 71.910 44.425 72.190 45.355 ;
        RECT 72.370 44.795 72.560 45.175 ;
        RECT 72.740 45.015 73.015 45.355 ;
        RECT 73.185 45.015 73.515 46.155 ;
        RECT 73.690 45.355 73.945 46.155 ;
        RECT 74.145 45.305 74.475 45.985 ;
        RECT 73.690 44.815 73.935 45.175 ;
        RECT 74.125 45.025 74.475 45.305 ;
        RECT 72.370 44.595 73.515 44.795 ;
        RECT 74.125 44.645 74.295 45.025 ;
        RECT 74.655 44.845 74.850 45.895 ;
        RECT 75.030 45.015 75.350 46.155 ;
        RECT 75.525 45.065 76.735 46.155 ;
        RECT 73.775 44.475 74.295 44.645 ;
        RECT 74.465 44.515 74.850 44.845 ;
        RECT 75.030 44.795 75.290 44.845 ;
        RECT 75.030 44.625 75.295 44.795 ;
        RECT 75.030 44.515 75.290 44.625 ;
        RECT 75.525 44.525 76.045 45.065 ;
        RECT 69.530 43.605 69.835 44.115 ;
        RECT 70.005 43.605 70.295 44.330 ;
        RECT 70.490 44.030 70.725 44.360 ;
        RECT 70.895 43.605 71.225 44.345 ;
        RECT 71.460 43.985 71.735 44.425 ;
        RECT 71.910 44.325 72.235 44.425 ;
        RECT 71.905 44.155 72.235 44.325 ;
        RECT 72.405 44.215 73.515 44.425 ;
        RECT 72.405 43.985 72.655 44.215 ;
        RECT 71.460 43.775 72.655 43.985 ;
        RECT 72.825 43.605 72.995 44.045 ;
        RECT 73.165 43.775 73.515 44.215 ;
        RECT 73.775 43.910 73.945 44.475 ;
        RECT 76.215 44.355 76.735 44.895 ;
        RECT 74.135 44.135 75.350 44.305 ;
        RECT 74.135 43.830 74.365 44.135 ;
        RECT 74.535 43.605 74.865 43.965 ;
        RECT 75.060 43.785 75.350 44.135 ;
        RECT 75.525 43.605 76.735 44.355 ;
        RECT 5.520 43.435 76.820 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.985 42.665 8.655 43.435 ;
        RECT 9.290 42.695 9.545 43.265 ;
        RECT 9.715 43.035 10.045 43.435 ;
        RECT 10.470 42.900 11.000 43.265 ;
        RECT 11.190 43.095 11.465 43.265 ;
        RECT 11.185 42.925 11.465 43.095 ;
        RECT 10.470 42.865 10.645 42.900 ;
        RECT 9.715 42.695 10.645 42.865 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 6.985 42.145 7.735 42.665 ;
        RECT 7.905 41.975 8.655 42.495 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 6.985 40.885 8.655 41.975 ;
        RECT 9.290 42.025 9.460 42.695 ;
        RECT 9.715 42.525 9.885 42.695 ;
        RECT 9.630 42.195 9.885 42.525 ;
        RECT 10.110 42.195 10.305 42.525 ;
        RECT 9.290 41.055 9.625 42.025 ;
        RECT 9.795 40.885 9.965 42.025 ;
        RECT 10.135 41.225 10.305 42.195 ;
        RECT 10.475 41.565 10.645 42.695 ;
        RECT 10.815 41.905 10.985 42.705 ;
        RECT 11.190 42.105 11.465 42.925 ;
        RECT 11.635 41.905 11.825 43.265 ;
        RECT 12.005 42.900 12.515 43.435 ;
        RECT 12.735 42.625 12.980 43.230 ;
        RECT 13.425 42.665 16.015 43.435 ;
        RECT 16.195 42.705 16.495 43.435 ;
        RECT 12.025 42.455 13.255 42.625 ;
        RECT 10.815 41.735 11.825 41.905 ;
        RECT 11.995 41.890 12.745 42.080 ;
        RECT 10.475 41.395 11.600 41.565 ;
        RECT 11.995 41.225 12.165 41.890 ;
        RECT 12.915 41.645 13.255 42.455 ;
        RECT 13.425 42.145 14.635 42.665 ;
        RECT 16.675 42.525 16.905 43.145 ;
        RECT 17.105 42.875 17.330 43.255 ;
        RECT 17.500 43.045 17.830 43.435 ;
        RECT 17.105 42.695 17.435 42.875 ;
        RECT 14.805 41.975 16.015 42.495 ;
        RECT 16.200 42.195 16.495 42.525 ;
        RECT 16.675 42.195 17.090 42.525 ;
        RECT 17.260 42.025 17.435 42.695 ;
        RECT 17.605 42.195 17.845 42.845 ;
        RECT 18.060 42.695 18.675 43.265 ;
        RECT 18.845 42.925 19.060 43.435 ;
        RECT 19.290 42.925 19.570 43.255 ;
        RECT 19.750 42.925 19.990 43.435 ;
        RECT 10.135 41.055 12.165 41.225 ;
        RECT 12.335 40.885 12.505 41.645 ;
        RECT 12.740 41.235 13.255 41.645 ;
        RECT 13.425 40.885 16.015 41.975 ;
        RECT 16.195 41.665 17.090 41.995 ;
        RECT 17.260 41.835 17.845 42.025 ;
        RECT 16.195 41.495 17.400 41.665 ;
        RECT 16.195 41.065 16.525 41.495 ;
        RECT 16.705 40.885 16.900 41.325 ;
        RECT 17.070 41.065 17.400 41.495 ;
        RECT 17.570 41.065 17.845 41.835 ;
        RECT 18.060 41.675 18.375 42.695 ;
        RECT 18.545 42.025 18.715 42.525 ;
        RECT 18.965 42.195 19.230 42.755 ;
        RECT 19.400 42.025 19.570 42.925 ;
        RECT 20.325 42.825 20.665 43.240 ;
        RECT 20.835 42.995 21.005 43.435 ;
        RECT 21.175 43.045 22.425 43.225 ;
        RECT 21.175 42.825 21.505 43.045 ;
        RECT 22.695 42.975 22.865 43.435 ;
        RECT 19.740 42.195 20.095 42.755 ;
        RECT 20.325 42.655 21.505 42.825 ;
        RECT 21.675 42.805 22.040 42.875 ;
        RECT 21.675 42.625 22.925 42.805 ;
        RECT 20.325 42.245 20.790 42.445 ;
        RECT 20.965 42.195 21.295 42.445 ;
        RECT 21.465 42.415 21.930 42.445 ;
        RECT 21.465 42.245 21.935 42.415 ;
        RECT 21.465 42.195 21.930 42.245 ;
        RECT 22.125 42.195 22.480 42.445 ;
        RECT 20.965 42.075 21.145 42.195 ;
        RECT 18.545 41.855 19.970 42.025 ;
        RECT 18.060 41.055 18.595 41.675 ;
        RECT 18.765 40.885 19.095 41.685 ;
        RECT 19.580 41.680 19.970 41.855 ;
        RECT 20.325 40.885 20.645 42.065 ;
        RECT 20.815 41.905 21.145 42.075 ;
        RECT 22.650 42.025 22.925 42.625 ;
        RECT 20.815 41.115 21.015 41.905 ;
        RECT 21.315 41.815 22.925 42.025 ;
        RECT 21.315 41.715 21.725 41.815 ;
        RECT 21.340 41.055 21.725 41.715 ;
        RECT 22.120 40.885 22.905 41.645 ;
        RECT 23.095 41.055 23.375 43.155 ;
        RECT 24.010 42.695 24.265 43.265 ;
        RECT 24.435 43.035 24.765 43.435 ;
        RECT 25.190 42.900 25.720 43.265 ;
        RECT 25.190 42.865 25.365 42.900 ;
        RECT 24.435 42.695 25.365 42.865 ;
        RECT 24.010 42.025 24.180 42.695 ;
        RECT 24.435 42.525 24.605 42.695 ;
        RECT 24.350 42.195 24.605 42.525 ;
        RECT 24.830 42.195 25.025 42.525 ;
        RECT 24.010 41.055 24.345 42.025 ;
        RECT 24.515 40.885 24.685 42.025 ;
        RECT 24.855 41.225 25.025 42.195 ;
        RECT 25.195 41.565 25.365 42.695 ;
        RECT 25.535 41.905 25.705 42.705 ;
        RECT 25.910 42.415 26.185 43.265 ;
        RECT 25.905 42.245 26.185 42.415 ;
        RECT 25.910 42.105 26.185 42.245 ;
        RECT 26.355 41.905 26.545 43.265 ;
        RECT 26.725 42.900 27.235 43.435 ;
        RECT 27.455 42.625 27.700 43.230 ;
        RECT 28.145 42.665 30.735 43.435 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 31.835 42.705 32.135 43.435 ;
        RECT 26.745 42.455 27.975 42.625 ;
        RECT 25.535 41.735 26.545 41.905 ;
        RECT 26.715 41.890 27.465 42.080 ;
        RECT 25.195 41.395 26.320 41.565 ;
        RECT 26.715 41.225 26.885 41.890 ;
        RECT 27.635 41.645 27.975 42.455 ;
        RECT 28.145 42.145 29.355 42.665 ;
        RECT 32.315 42.525 32.545 43.145 ;
        RECT 32.745 42.875 32.970 43.255 ;
        RECT 33.140 43.045 33.470 43.435 ;
        RECT 32.745 42.695 33.075 42.875 ;
        RECT 29.525 41.975 30.735 42.495 ;
        RECT 31.840 42.195 32.135 42.525 ;
        RECT 32.315 42.195 32.730 42.525 ;
        RECT 24.855 41.055 26.885 41.225 ;
        RECT 27.055 40.885 27.225 41.645 ;
        RECT 27.460 41.235 27.975 41.645 ;
        RECT 28.145 40.885 30.735 41.975 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 32.900 42.025 33.075 42.695 ;
        RECT 33.245 42.195 33.485 42.845 ;
        RECT 31.835 41.665 32.730 41.995 ;
        RECT 32.900 41.835 33.485 42.025 ;
        RECT 31.835 41.495 33.040 41.665 ;
        RECT 31.835 41.065 32.165 41.495 ;
        RECT 32.345 40.885 32.540 41.325 ;
        RECT 32.710 41.065 33.040 41.495 ;
        RECT 33.210 41.065 33.485 41.835 ;
        RECT 34.135 41.065 34.395 43.255 ;
        RECT 34.655 43.065 35.325 43.435 ;
        RECT 35.505 42.885 35.815 43.255 ;
        RECT 34.585 42.685 35.815 42.885 ;
        RECT 34.585 42.015 34.875 42.685 ;
        RECT 35.995 42.505 36.225 43.145 ;
        RECT 36.405 42.705 36.695 43.435 ;
        RECT 36.885 42.665 39.475 43.435 ;
        RECT 39.670 43.045 40.000 43.435 ;
        RECT 40.170 42.875 40.395 43.255 ;
        RECT 35.055 42.195 35.520 42.505 ;
        RECT 35.700 42.195 36.225 42.505 ;
        RECT 36.405 42.195 36.705 42.525 ;
        RECT 36.885 42.145 38.095 42.665 ;
        RECT 34.585 41.795 35.355 42.015 ;
        RECT 34.565 40.885 34.905 41.615 ;
        RECT 35.085 41.065 35.355 41.795 ;
        RECT 35.535 41.775 36.695 42.015 ;
        RECT 38.265 41.975 39.475 42.495 ;
        RECT 39.655 42.195 39.895 42.845 ;
        RECT 40.065 42.695 40.395 42.875 ;
        RECT 40.065 42.025 40.240 42.695 ;
        RECT 40.595 42.525 40.825 43.145 ;
        RECT 41.005 42.705 41.305 43.435 ;
        RECT 42.430 43.045 42.760 43.435 ;
        RECT 42.930 42.875 43.155 43.255 ;
        RECT 40.410 42.195 40.825 42.525 ;
        RECT 41.005 42.195 41.300 42.525 ;
        RECT 42.415 42.195 42.655 42.845 ;
        RECT 42.825 42.695 43.155 42.875 ;
        RECT 42.825 42.025 43.000 42.695 ;
        RECT 43.355 42.525 43.585 43.145 ;
        RECT 43.765 42.705 44.065 43.435 ;
        RECT 44.245 42.665 45.915 43.435 ;
        RECT 43.170 42.195 43.585 42.525 ;
        RECT 43.765 42.195 44.060 42.525 ;
        RECT 44.245 42.145 44.995 42.665 ;
        RECT 35.535 41.065 35.765 41.775 ;
        RECT 35.935 40.885 36.265 41.595 ;
        RECT 36.435 41.065 36.695 41.775 ;
        RECT 36.885 40.885 39.475 41.975 ;
        RECT 39.655 41.835 40.240 42.025 ;
        RECT 39.655 41.065 39.930 41.835 ;
        RECT 40.410 41.665 41.305 41.995 ;
        RECT 40.100 41.495 41.305 41.665 ;
        RECT 40.100 41.065 40.430 41.495 ;
        RECT 40.600 40.885 40.795 41.325 ;
        RECT 40.975 41.065 41.305 41.495 ;
        RECT 42.415 41.835 43.000 42.025 ;
        RECT 42.415 41.065 42.690 41.835 ;
        RECT 43.170 41.665 44.065 41.995 ;
        RECT 45.165 41.975 45.915 42.495 ;
        RECT 42.860 41.495 44.065 41.665 ;
        RECT 42.860 41.065 43.190 41.495 ;
        RECT 43.360 40.885 43.555 41.325 ;
        RECT 43.735 41.065 44.065 41.495 ;
        RECT 44.245 40.885 45.915 41.975 ;
        RECT 46.560 41.065 46.840 43.255 ;
        RECT 47.040 43.065 47.770 43.435 ;
        RECT 48.350 42.895 48.780 43.255 ;
        RECT 47.040 42.705 48.780 42.895 ;
        RECT 47.040 42.195 47.300 42.705 ;
        RECT 47.030 40.885 47.315 42.025 ;
        RECT 47.510 41.905 47.770 42.525 ;
        RECT 47.965 41.905 48.390 42.525 ;
        RECT 48.560 42.475 48.780 42.705 ;
        RECT 48.950 42.655 49.195 43.435 ;
        RECT 48.560 42.175 49.105 42.475 ;
        RECT 49.395 42.355 49.625 43.255 ;
        RECT 47.580 41.535 48.605 41.735 ;
        RECT 47.580 41.065 47.750 41.535 ;
        RECT 47.925 40.885 48.255 41.365 ;
        RECT 48.425 41.065 48.605 41.535 ;
        RECT 48.775 41.065 49.105 42.175 ;
        RECT 49.285 41.675 49.625 42.355 ;
        RECT 49.805 41.855 50.035 43.195 ;
        RECT 50.775 42.885 50.945 43.265 ;
        RECT 51.125 43.055 51.455 43.435 ;
        RECT 50.775 42.715 51.440 42.885 ;
        RECT 51.635 42.760 51.895 43.265 ;
        RECT 50.705 42.165 51.035 42.535 ;
        RECT 51.270 42.460 51.440 42.715 ;
        RECT 51.270 42.130 51.555 42.460 ;
        RECT 51.270 41.985 51.440 42.130 ;
        RECT 50.775 41.815 51.440 41.985 ;
        RECT 51.725 41.960 51.895 42.760 ;
        RECT 52.155 42.885 52.325 43.265 ;
        RECT 52.505 43.055 52.835 43.435 ;
        RECT 52.155 42.715 52.820 42.885 ;
        RECT 53.015 42.760 53.275 43.265 ;
        RECT 52.085 42.165 52.425 42.535 ;
        RECT 52.650 42.460 52.820 42.715 ;
        RECT 52.650 42.130 52.925 42.460 ;
        RECT 52.650 41.985 52.820 42.130 ;
        RECT 49.285 41.475 50.035 41.675 ;
        RECT 49.275 40.885 49.625 41.295 ;
        RECT 49.795 41.085 50.035 41.475 ;
        RECT 50.775 41.055 50.945 41.815 ;
        RECT 51.125 40.885 51.455 41.645 ;
        RECT 51.625 41.055 51.895 41.960 ;
        RECT 52.145 41.815 52.820 41.985 ;
        RECT 53.095 41.960 53.275 42.760 ;
        RECT 52.145 41.055 52.325 41.815 ;
        RECT 52.505 40.885 52.835 41.645 ;
        RECT 53.005 41.055 53.275 41.960 ;
        RECT 53.465 42.935 53.720 43.265 ;
        RECT 53.935 42.955 54.265 43.435 ;
        RECT 54.435 43.015 55.970 43.265 ;
        RECT 53.465 42.855 53.650 42.935 ;
        RECT 53.465 41.725 53.635 42.855 ;
        RECT 54.435 42.785 54.605 43.015 ;
        RECT 53.805 42.615 54.605 42.785 ;
        RECT 53.805 42.065 53.975 42.615 ;
        RECT 54.785 42.445 55.070 42.845 ;
        RECT 54.205 42.415 54.570 42.445 ;
        RECT 54.195 42.245 54.570 42.415 ;
        RECT 54.740 42.245 55.070 42.445 ;
        RECT 55.340 42.445 55.620 42.845 ;
        RECT 55.800 42.785 55.970 43.015 ;
        RECT 56.195 42.955 56.525 43.435 ;
        RECT 56.695 42.785 56.865 43.265 ;
        RECT 55.800 42.615 56.865 42.785 ;
        RECT 57.125 42.710 57.415 43.435 ;
        RECT 58.510 42.615 58.785 43.435 ;
        RECT 58.955 42.795 59.285 43.265 ;
        RECT 59.455 42.965 59.625 43.435 ;
        RECT 59.795 42.795 60.125 43.265 ;
        RECT 60.295 42.965 60.585 43.435 ;
        RECT 58.955 42.785 60.125 42.795 ;
        RECT 60.960 42.785 61.290 43.250 ;
        RECT 61.460 42.965 61.630 43.435 ;
        RECT 61.800 42.785 62.130 43.265 ;
        RECT 58.955 42.615 60.555 42.785 ;
        RECT 60.960 42.615 62.130 42.785 ;
        RECT 55.340 42.245 55.815 42.445 ;
        RECT 55.985 42.245 56.430 42.445 ;
        RECT 56.600 42.235 56.950 42.445 ;
        RECT 58.510 42.245 59.230 42.445 ;
        RECT 59.400 42.245 60.170 42.445 ;
        RECT 60.340 42.075 60.555 42.615 ;
        RECT 60.805 42.235 61.450 42.445 ;
        RECT 61.620 42.235 62.190 42.445 ;
        RECT 53.805 41.895 56.865 42.065 ;
        RECT 53.465 41.055 53.720 41.725 ;
        RECT 53.890 40.885 54.220 41.645 ;
        RECT 54.390 41.485 56.025 41.725 ;
        RECT 54.390 41.055 54.640 41.485 ;
        RECT 55.795 41.395 56.025 41.485 ;
        RECT 54.810 40.885 55.165 41.305 ;
        RECT 55.355 41.225 55.685 41.265 ;
        RECT 56.195 41.225 56.525 41.725 ;
        RECT 55.355 41.055 56.525 41.225 ;
        RECT 56.695 41.055 56.865 41.895 ;
        RECT 57.125 40.885 57.415 42.050 ;
        RECT 58.510 41.855 59.625 42.065 ;
        RECT 58.510 41.055 58.785 41.855 ;
        RECT 58.955 40.885 59.285 41.685 ;
        RECT 59.455 41.225 59.625 41.855 ;
        RECT 59.795 41.905 60.575 42.075 ;
        RECT 62.360 42.065 62.530 43.265 ;
        RECT 63.070 42.865 63.240 43.070 ;
        RECT 59.795 41.855 60.555 41.905 ;
        RECT 59.795 41.395 60.125 41.855 ;
        RECT 60.295 41.225 60.595 41.685 ;
        RECT 59.455 41.055 60.595 41.225 ;
        RECT 61.020 40.885 61.350 41.985 ;
        RECT 61.825 41.655 62.530 42.065 ;
        RECT 62.700 42.695 63.240 42.865 ;
        RECT 63.520 42.695 63.690 43.435 ;
        RECT 63.955 42.695 64.315 43.070 ;
        RECT 64.575 42.885 64.745 43.265 ;
        RECT 64.960 43.055 65.290 43.435 ;
        RECT 64.575 42.715 65.290 42.885 ;
        RECT 62.700 41.995 62.870 42.695 ;
        RECT 63.040 42.195 63.370 42.525 ;
        RECT 63.540 42.195 63.890 42.525 ;
        RECT 62.700 41.825 63.325 41.995 ;
        RECT 63.540 41.655 63.805 42.195 ;
        RECT 64.060 42.040 64.315 42.695 ;
        RECT 64.485 42.165 64.840 42.535 ;
        RECT 65.120 42.525 65.290 42.715 ;
        RECT 65.460 42.690 65.715 43.265 ;
        RECT 65.120 42.195 65.375 42.525 ;
        RECT 61.825 41.485 63.805 41.655 ;
        RECT 61.825 41.055 62.150 41.485 ;
        RECT 62.320 40.885 62.650 41.305 ;
        RECT 63.395 40.885 63.805 41.315 ;
        RECT 63.975 41.055 64.315 42.040 ;
        RECT 65.120 41.985 65.290 42.195 ;
        RECT 64.575 41.815 65.290 41.985 ;
        RECT 65.545 41.960 65.715 42.690 ;
        RECT 65.890 42.595 66.150 43.435 ;
        RECT 66.325 42.925 66.630 43.435 ;
        RECT 66.325 42.195 66.640 42.755 ;
        RECT 66.810 42.445 67.060 43.255 ;
        RECT 67.230 42.910 67.490 43.435 ;
        RECT 67.670 42.445 67.920 43.255 ;
        RECT 68.090 42.875 68.350 43.435 ;
        RECT 68.520 42.785 68.780 43.240 ;
        RECT 68.950 42.955 69.210 43.435 ;
        RECT 69.380 42.785 69.640 43.240 ;
        RECT 69.810 42.955 70.070 43.435 ;
        RECT 70.240 42.785 70.500 43.240 ;
        RECT 70.670 42.955 70.915 43.435 ;
        RECT 71.085 42.785 71.360 43.240 ;
        RECT 71.530 42.955 71.775 43.435 ;
        RECT 71.945 42.785 72.205 43.240 ;
        RECT 72.385 42.955 72.635 43.435 ;
        RECT 72.805 42.785 73.065 43.240 ;
        RECT 73.245 42.955 73.495 43.435 ;
        RECT 73.665 42.785 73.925 43.240 ;
        RECT 74.105 42.955 74.365 43.435 ;
        RECT 74.535 42.785 74.795 43.240 ;
        RECT 74.965 42.955 75.265 43.435 ;
        RECT 68.520 42.615 75.265 42.785 ;
        RECT 75.525 42.685 76.735 43.435 ;
        RECT 66.810 42.195 73.930 42.445 ;
        RECT 64.575 41.055 64.745 41.815 ;
        RECT 64.960 40.885 65.290 41.645 ;
        RECT 65.460 41.055 65.715 41.960 ;
        RECT 65.890 40.885 66.150 42.035 ;
        RECT 66.335 40.885 66.630 41.695 ;
        RECT 66.810 41.055 67.055 42.195 ;
        RECT 67.230 40.885 67.490 41.695 ;
        RECT 67.670 41.060 67.920 42.195 ;
        RECT 74.100 42.025 75.265 42.615 ;
        RECT 68.520 41.800 75.265 42.025 ;
        RECT 75.525 41.975 76.045 42.515 ;
        RECT 76.215 42.145 76.735 42.685 ;
        RECT 68.520 41.785 73.925 41.800 ;
        RECT 68.090 40.890 68.350 41.685 ;
        RECT 68.520 41.060 68.780 41.785 ;
        RECT 68.950 40.890 69.210 41.615 ;
        RECT 69.380 41.060 69.640 41.785 ;
        RECT 69.810 40.890 70.070 41.615 ;
        RECT 70.240 41.060 70.500 41.785 ;
        RECT 70.670 40.890 70.930 41.615 ;
        RECT 71.100 41.060 71.360 41.785 ;
        RECT 71.530 40.890 71.775 41.615 ;
        RECT 71.945 41.060 72.205 41.785 ;
        RECT 72.390 40.890 72.635 41.615 ;
        RECT 72.805 41.060 73.065 41.785 ;
        RECT 73.250 40.890 73.495 41.615 ;
        RECT 73.665 41.060 73.925 41.785 ;
        RECT 74.110 40.890 74.365 41.615 ;
        RECT 74.535 41.060 74.825 41.800 ;
        RECT 68.090 40.885 74.365 40.890 ;
        RECT 74.995 40.885 75.265 41.630 ;
        RECT 75.525 40.885 76.735 41.975 ;
        RECT 5.520 40.715 76.820 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 6.985 39.625 8.655 40.715 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 6.985 38.935 7.735 39.455 ;
        RECT 7.905 39.105 8.655 39.625 ;
        RECT 8.830 39.575 9.165 40.545 ;
        RECT 9.335 39.575 9.505 40.715 ;
        RECT 9.675 40.375 11.705 40.545 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 6.985 38.165 8.655 38.935 ;
        RECT 8.830 38.905 9.000 39.575 ;
        RECT 9.675 39.405 9.845 40.375 ;
        RECT 9.170 39.075 9.425 39.405 ;
        RECT 9.650 39.075 9.845 39.405 ;
        RECT 10.015 40.035 11.140 40.205 ;
        RECT 9.255 38.905 9.425 39.075 ;
        RECT 10.015 38.905 10.185 40.035 ;
        RECT 8.830 38.335 9.085 38.905 ;
        RECT 9.255 38.735 10.185 38.905 ;
        RECT 10.355 39.695 11.365 39.865 ;
        RECT 10.355 38.895 10.525 39.695 ;
        RECT 10.010 38.700 10.185 38.735 ;
        RECT 9.255 38.165 9.585 38.565 ;
        RECT 10.010 38.335 10.540 38.700 ;
        RECT 10.730 38.675 11.005 39.495 ;
        RECT 10.725 38.505 11.005 38.675 ;
        RECT 10.730 38.335 11.005 38.505 ;
        RECT 11.175 38.335 11.365 39.695 ;
        RECT 11.535 39.710 11.705 40.375 ;
        RECT 11.875 39.955 12.045 40.715 ;
        RECT 12.280 39.955 12.795 40.365 ;
        RECT 11.535 39.520 12.285 39.710 ;
        RECT 12.455 39.145 12.795 39.955 ;
        RECT 12.965 39.625 14.635 40.715 ;
        RECT 11.565 38.975 12.795 39.145 ;
        RECT 11.545 38.165 12.055 38.700 ;
        RECT 12.275 38.370 12.520 38.975 ;
        RECT 12.965 38.935 13.715 39.455 ;
        RECT 13.885 39.105 14.635 39.625 ;
        RECT 15.275 40.105 15.605 40.535 ;
        RECT 15.785 40.275 15.980 40.715 ;
        RECT 16.150 40.105 16.480 40.535 ;
        RECT 15.275 39.935 16.480 40.105 ;
        RECT 15.275 39.605 16.170 39.935 ;
        RECT 16.650 39.765 16.925 40.535 ;
        RECT 16.340 39.575 16.925 39.765 ;
        RECT 17.105 39.625 18.315 40.715 ;
        RECT 15.280 39.075 15.575 39.405 ;
        RECT 15.755 39.075 16.170 39.405 ;
        RECT 12.965 38.165 14.635 38.935 ;
        RECT 15.275 38.165 15.575 38.895 ;
        RECT 15.755 38.455 15.985 39.075 ;
        RECT 16.340 38.905 16.515 39.575 ;
        RECT 16.185 38.725 16.515 38.905 ;
        RECT 16.685 38.755 16.925 39.405 ;
        RECT 17.105 38.915 17.625 39.455 ;
        RECT 17.795 39.085 18.315 39.625 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.980 39.925 19.515 40.545 ;
        RECT 16.185 38.345 16.410 38.725 ;
        RECT 16.580 38.165 16.910 38.555 ;
        RECT 17.105 38.165 18.315 38.915 ;
        RECT 18.980 38.905 19.295 39.925 ;
        RECT 19.685 39.915 20.015 40.715 ;
        RECT 21.255 40.105 21.585 40.535 ;
        RECT 21.765 40.275 21.960 40.715 ;
        RECT 22.130 40.105 22.460 40.535 ;
        RECT 21.255 39.935 22.460 40.105 ;
        RECT 20.500 39.745 20.890 39.920 ;
        RECT 19.465 39.575 20.890 39.745 ;
        RECT 21.255 39.605 22.150 39.935 ;
        RECT 22.630 39.765 22.905 40.535 ;
        RECT 22.320 39.575 22.905 39.765 ;
        RECT 24.010 39.575 24.345 40.545 ;
        RECT 24.515 39.575 24.685 40.715 ;
        RECT 24.855 40.375 26.885 40.545 ;
        RECT 19.465 39.075 19.635 39.575 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 18.980 38.335 19.595 38.905 ;
        RECT 19.885 38.845 20.150 39.405 ;
        RECT 20.320 38.675 20.490 39.575 ;
        RECT 20.660 38.845 21.015 39.405 ;
        RECT 21.260 39.075 21.555 39.405 ;
        RECT 21.735 39.075 22.150 39.405 ;
        RECT 19.765 38.165 19.980 38.675 ;
        RECT 20.210 38.345 20.490 38.675 ;
        RECT 20.670 38.165 20.910 38.675 ;
        RECT 21.255 38.165 21.555 38.895 ;
        RECT 21.735 38.455 21.965 39.075 ;
        RECT 22.320 38.905 22.495 39.575 ;
        RECT 22.165 38.725 22.495 38.905 ;
        RECT 22.665 38.755 22.905 39.405 ;
        RECT 24.010 38.905 24.180 39.575 ;
        RECT 24.855 39.405 25.025 40.375 ;
        RECT 24.350 39.075 24.605 39.405 ;
        RECT 24.830 39.075 25.025 39.405 ;
        RECT 25.195 40.035 26.320 40.205 ;
        RECT 24.435 38.905 24.605 39.075 ;
        RECT 25.195 38.905 25.365 40.035 ;
        RECT 22.165 38.345 22.390 38.725 ;
        RECT 22.560 38.165 22.890 38.555 ;
        RECT 24.010 38.335 24.265 38.905 ;
        RECT 24.435 38.735 25.365 38.905 ;
        RECT 25.535 39.695 26.545 39.865 ;
        RECT 25.535 38.895 25.705 39.695 ;
        RECT 25.190 38.700 25.365 38.735 ;
        RECT 24.435 38.165 24.765 38.565 ;
        RECT 25.190 38.335 25.720 38.700 ;
        RECT 25.910 38.675 26.185 39.495 ;
        RECT 25.905 38.505 26.185 38.675 ;
        RECT 25.910 38.335 26.185 38.505 ;
        RECT 26.355 38.335 26.545 39.695 ;
        RECT 26.715 39.710 26.885 40.375 ;
        RECT 27.055 39.955 27.225 40.715 ;
        RECT 27.460 39.955 27.975 40.365 ;
        RECT 26.715 39.520 27.465 39.710 ;
        RECT 27.635 39.145 27.975 39.955 ;
        RECT 28.185 39.575 28.415 40.715 ;
        RECT 28.585 39.565 28.915 40.545 ;
        RECT 29.085 39.575 29.295 40.715 ;
        RECT 29.525 39.575 29.785 40.715 ;
        RECT 29.955 39.565 30.285 40.545 ;
        RECT 30.455 39.575 30.735 40.715 ;
        RECT 30.905 39.625 32.115 40.715 ;
        RECT 28.165 39.155 28.495 39.405 ;
        RECT 26.745 38.975 27.975 39.145 ;
        RECT 26.725 38.165 27.235 38.700 ;
        RECT 27.455 38.370 27.700 38.975 ;
        RECT 28.185 38.165 28.415 38.985 ;
        RECT 28.665 38.965 28.915 39.565 ;
        RECT 30.045 39.525 30.220 39.565 ;
        RECT 29.545 39.155 29.880 39.405 ;
        RECT 28.585 38.335 28.915 38.965 ;
        RECT 29.085 38.165 29.295 38.985 ;
        RECT 30.050 38.965 30.220 39.525 ;
        RECT 30.390 39.135 30.725 39.405 ;
        RECT 29.525 38.335 30.220 38.965 ;
        RECT 30.425 38.165 30.735 38.965 ;
        RECT 30.905 38.915 31.425 39.455 ;
        RECT 31.595 39.085 32.115 39.625 ;
        RECT 32.295 39.765 32.570 40.535 ;
        RECT 32.740 40.105 33.070 40.535 ;
        RECT 33.240 40.275 33.435 40.715 ;
        RECT 33.615 40.105 33.945 40.535 ;
        RECT 32.740 39.935 33.945 40.105 ;
        RECT 32.295 39.575 32.880 39.765 ;
        RECT 33.050 39.605 33.945 39.935 ;
        RECT 34.125 39.625 35.795 40.715 ;
        RECT 30.905 38.165 32.115 38.915 ;
        RECT 32.295 38.755 32.535 39.405 ;
        RECT 32.705 38.905 32.880 39.575 ;
        RECT 33.050 39.075 33.465 39.405 ;
        RECT 33.645 39.075 33.940 39.405 ;
        RECT 32.705 38.725 33.035 38.905 ;
        RECT 32.310 38.165 32.640 38.555 ;
        RECT 32.810 38.345 33.035 38.725 ;
        RECT 33.235 38.455 33.465 39.075 ;
        RECT 34.125 38.935 34.875 39.455 ;
        RECT 35.045 39.105 35.795 39.625 ;
        RECT 36.425 39.575 36.685 40.715 ;
        RECT 36.855 39.565 37.185 40.545 ;
        RECT 37.355 39.575 37.635 40.715 ;
        RECT 37.805 40.280 43.150 40.715 ;
        RECT 36.445 39.155 36.780 39.405 ;
        RECT 36.950 38.965 37.120 39.565 ;
        RECT 37.290 39.135 37.625 39.405 ;
        RECT 33.645 38.165 33.945 38.895 ;
        RECT 34.125 38.165 35.795 38.935 ;
        RECT 36.425 38.335 37.120 38.965 ;
        RECT 37.325 38.165 37.635 38.965 ;
        RECT 39.390 38.710 39.730 39.540 ;
        RECT 41.210 39.030 41.560 40.280 ;
        RECT 44.245 39.550 44.535 40.715 ;
        RECT 44.705 39.575 44.980 40.545 ;
        RECT 45.190 39.915 45.470 40.715 ;
        RECT 45.640 40.205 47.255 40.535 ;
        RECT 45.640 39.865 46.815 40.035 ;
        RECT 45.640 39.745 45.810 39.865 ;
        RECT 45.150 39.575 45.810 39.745 ;
        RECT 37.805 38.165 43.150 38.710 ;
        RECT 44.245 38.165 44.535 38.890 ;
        RECT 44.705 38.840 44.875 39.575 ;
        RECT 45.150 39.405 45.320 39.575 ;
        RECT 46.070 39.405 46.315 39.695 ;
        RECT 46.485 39.575 46.815 39.865 ;
        RECT 47.075 39.405 47.245 39.965 ;
        RECT 47.495 39.575 47.755 40.715 ;
        RECT 47.925 39.625 51.435 40.715 ;
        RECT 45.045 39.075 45.320 39.405 ;
        RECT 45.490 39.075 46.315 39.405 ;
        RECT 46.530 39.075 47.245 39.405 ;
        RECT 47.415 39.155 47.750 39.405 ;
        RECT 45.150 38.905 45.320 39.075 ;
        RECT 46.995 38.985 47.245 39.075 ;
        RECT 44.705 38.495 44.980 38.840 ;
        RECT 45.150 38.735 46.815 38.905 ;
        RECT 45.170 38.165 45.545 38.565 ;
        RECT 45.715 38.385 45.885 38.735 ;
        RECT 46.055 38.165 46.385 38.565 ;
        RECT 46.555 38.335 46.815 38.735 ;
        RECT 46.995 38.565 47.325 38.985 ;
        RECT 47.495 38.165 47.755 38.985 ;
        RECT 47.925 38.935 49.575 39.455 ;
        RECT 49.745 39.105 51.435 39.625 ;
        RECT 52.070 39.765 52.335 40.535 ;
        RECT 52.505 39.995 52.835 40.715 ;
        RECT 53.025 40.175 53.285 40.535 ;
        RECT 53.455 40.345 53.785 40.715 ;
        RECT 53.955 40.175 54.215 40.535 ;
        RECT 53.025 39.945 54.215 40.175 ;
        RECT 54.785 39.765 55.075 40.535 ;
        RECT 47.925 38.165 51.435 38.935 ;
        RECT 52.070 38.345 52.405 39.765 ;
        RECT 52.580 39.585 55.075 39.765 ;
        RECT 55.285 39.625 56.495 40.715 ;
        RECT 52.580 38.895 52.805 39.585 ;
        RECT 53.005 39.075 53.285 39.405 ;
        RECT 53.465 39.075 54.040 39.405 ;
        RECT 54.220 39.075 54.655 39.405 ;
        RECT 54.835 39.075 55.105 39.405 ;
        RECT 55.285 38.915 55.805 39.455 ;
        RECT 55.975 39.085 56.495 39.625 ;
        RECT 56.665 39.575 56.955 40.715 ;
        RECT 57.125 39.995 57.575 40.545 ;
        RECT 57.765 39.995 58.095 40.715 ;
        RECT 52.580 38.705 55.065 38.895 ;
        RECT 52.585 38.165 53.330 38.535 ;
        RECT 53.895 38.345 54.150 38.705 ;
        RECT 54.330 38.165 54.660 38.535 ;
        RECT 54.840 38.345 55.065 38.705 ;
        RECT 55.285 38.165 56.495 38.915 ;
        RECT 56.665 38.165 56.955 38.965 ;
        RECT 57.125 38.625 57.375 39.995 ;
        RECT 58.305 39.825 58.605 40.375 ;
        RECT 58.775 40.045 59.055 40.715 ;
        RECT 59.425 39.915 59.865 40.545 ;
        RECT 57.665 39.655 58.605 39.825 ;
        RECT 57.665 39.405 57.835 39.655 ;
        RECT 58.940 39.405 59.255 39.845 ;
        RECT 57.545 39.075 57.835 39.405 ;
        RECT 58.005 39.155 58.335 39.405 ;
        RECT 58.565 39.155 59.255 39.405 ;
        RECT 57.665 38.985 57.835 39.075 ;
        RECT 57.665 38.795 59.055 38.985 ;
        RECT 57.125 38.335 57.675 38.625 ;
        RECT 57.845 38.165 58.095 38.625 ;
        RECT 58.725 38.435 59.055 38.795 ;
        RECT 59.425 38.905 59.735 39.915 ;
        RECT 60.040 39.865 60.355 40.715 ;
        RECT 60.525 40.375 61.955 40.545 ;
        RECT 60.525 39.695 60.695 40.375 ;
        RECT 59.905 39.525 60.695 39.695 ;
        RECT 59.905 39.075 60.075 39.525 ;
        RECT 60.865 39.405 61.065 40.205 ;
        RECT 60.245 39.075 60.635 39.355 ;
        RECT 60.820 39.075 61.065 39.405 ;
        RECT 61.265 39.075 61.515 40.205 ;
        RECT 61.705 39.745 61.955 40.375 ;
        RECT 62.135 39.915 62.465 40.715 ;
        RECT 62.665 39.875 62.995 40.715 ;
        RECT 61.705 39.575 62.475 39.745 ;
        RECT 63.165 39.695 63.510 40.450 ;
        RECT 63.685 40.105 64.030 40.545 ;
        RECT 64.240 40.335 64.570 40.715 ;
        RECT 64.755 40.105 64.990 40.545 ;
        RECT 65.160 40.275 65.490 40.715 ;
        RECT 63.685 39.865 65.695 40.105 ;
        RECT 61.730 39.075 62.135 39.405 ;
        RECT 62.305 38.905 62.475 39.575 ;
        RECT 62.665 39.085 62.995 39.695 ;
        RECT 63.165 39.075 63.795 39.695 ;
        RECT 63.965 39.075 64.255 39.695 ;
        RECT 59.425 38.345 59.865 38.905 ;
        RECT 60.035 38.165 60.485 38.905 ;
        RECT 60.655 38.735 61.815 38.905 ;
        RECT 60.655 38.335 60.825 38.735 ;
        RECT 60.995 38.165 61.415 38.565 ;
        RECT 61.585 38.335 61.815 38.735 ;
        RECT 61.985 38.335 62.475 38.905 ;
        RECT 62.665 38.705 64.030 38.905 ;
        RECT 62.665 38.335 62.995 38.705 ;
        RECT 63.165 38.165 63.495 38.535 ;
        RECT 63.685 38.335 64.030 38.705 ;
        RECT 64.425 38.335 64.755 39.695 ;
        RECT 64.965 39.155 65.295 39.695 ;
        RECT 65.465 38.965 65.695 39.865 ;
        RECT 65.925 39.575 66.135 40.715 ;
        RECT 66.305 39.565 66.635 40.545 ;
        RECT 66.805 39.575 67.035 40.715 ;
        RECT 67.300 39.845 67.585 40.715 ;
        RECT 67.755 40.085 68.015 40.545 ;
        RECT 68.190 40.255 68.445 40.715 ;
        RECT 68.615 40.085 68.875 40.545 ;
        RECT 67.755 39.915 68.875 40.085 ;
        RECT 69.045 39.915 69.355 40.715 ;
        RECT 67.755 39.665 68.015 39.915 ;
        RECT 69.525 39.745 69.835 40.545 ;
        RECT 65.090 38.335 65.695 38.965 ;
        RECT 65.925 38.165 66.135 38.985 ;
        RECT 66.305 38.965 66.555 39.565 ;
        RECT 67.260 39.495 68.015 39.665 ;
        RECT 68.805 39.575 69.835 39.745 ;
        RECT 66.725 39.155 67.055 39.405 ;
        RECT 67.260 38.985 67.665 39.495 ;
        RECT 68.805 39.325 68.975 39.575 ;
        RECT 67.835 39.155 68.975 39.325 ;
        RECT 66.305 38.335 66.635 38.965 ;
        RECT 66.805 38.165 67.035 38.985 ;
        RECT 67.260 38.815 68.910 38.985 ;
        RECT 69.145 38.835 69.495 39.405 ;
        RECT 67.305 38.165 67.585 38.645 ;
        RECT 67.755 38.425 68.015 38.815 ;
        RECT 68.190 38.165 68.445 38.645 ;
        RECT 68.615 38.425 68.910 38.815 ;
        RECT 69.665 38.665 69.835 39.575 ;
        RECT 70.005 39.550 70.295 40.715 ;
        RECT 70.465 39.575 70.795 40.715 ;
        RECT 70.965 40.085 71.320 40.545 ;
        RECT 71.490 40.255 72.065 40.715 ;
        RECT 72.235 40.085 72.565 40.545 ;
        RECT 70.965 39.915 72.565 40.085 ;
        RECT 72.765 39.915 73.020 40.715 ;
        RECT 70.965 39.575 71.240 39.915 ;
        RECT 71.420 39.355 71.610 39.735 ;
        RECT 70.465 39.185 71.615 39.355 ;
        RECT 70.465 39.155 71.610 39.185 ;
        RECT 71.790 38.985 72.070 39.915 ;
        RECT 73.190 39.745 73.490 39.940 ;
        RECT 72.240 39.575 73.490 39.745 ;
        RECT 73.685 39.625 75.355 40.715 ;
        RECT 72.240 39.155 72.570 39.575 ;
        RECT 72.800 39.075 73.145 39.405 ;
        RECT 69.090 38.165 69.365 38.645 ;
        RECT 69.535 38.335 69.835 38.665 ;
        RECT 70.005 38.165 70.295 38.890 ;
        RECT 70.465 38.775 71.575 38.985 ;
        RECT 70.465 38.335 70.815 38.775 ;
        RECT 70.985 38.165 71.155 38.605 ;
        RECT 71.325 38.545 71.575 38.775 ;
        RECT 71.745 38.885 72.070 38.985 ;
        RECT 71.745 38.715 72.075 38.885 ;
        RECT 72.245 38.545 72.520 38.985 ;
        RECT 73.320 38.920 73.490 39.575 ;
        RECT 71.325 38.335 72.520 38.545 ;
        RECT 72.755 38.165 73.085 38.905 ;
        RECT 73.255 38.590 73.490 38.920 ;
        RECT 73.685 38.935 74.435 39.455 ;
        RECT 74.605 39.105 75.355 39.625 ;
        RECT 75.525 39.625 76.735 40.715 ;
        RECT 75.525 39.085 76.045 39.625 ;
        RECT 73.685 38.165 75.355 38.935 ;
        RECT 76.215 38.915 76.735 39.455 ;
        RECT 75.525 38.165 76.735 38.915 ;
        RECT 5.520 37.995 76.820 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 6.985 37.225 9.575 37.995 ;
        RECT 9.750 37.255 10.005 37.825 ;
        RECT 10.175 37.595 10.505 37.995 ;
        RECT 10.930 37.460 11.460 37.825 ;
        RECT 10.930 37.425 11.105 37.460 ;
        RECT 10.175 37.255 11.105 37.425 ;
        RECT 11.650 37.315 11.925 37.825 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 6.985 36.705 8.195 37.225 ;
        RECT 8.365 36.535 9.575 37.055 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 6.985 35.445 9.575 36.535 ;
        RECT 9.750 36.585 9.920 37.255 ;
        RECT 10.175 37.085 10.345 37.255 ;
        RECT 10.090 36.755 10.345 37.085 ;
        RECT 10.570 36.755 10.765 37.085 ;
        RECT 9.750 35.615 10.085 36.585 ;
        RECT 10.255 35.445 10.425 36.585 ;
        RECT 10.595 35.785 10.765 36.755 ;
        RECT 10.935 36.125 11.105 37.255 ;
        RECT 11.275 36.465 11.445 37.265 ;
        RECT 11.645 37.145 11.925 37.315 ;
        RECT 11.650 36.665 11.925 37.145 ;
        RECT 12.095 36.465 12.285 37.825 ;
        RECT 12.465 37.460 12.975 37.995 ;
        RECT 13.195 37.185 13.440 37.790 ;
        RECT 13.890 37.255 14.145 37.825 ;
        RECT 14.315 37.595 14.645 37.995 ;
        RECT 15.070 37.460 15.600 37.825 ;
        RECT 15.790 37.655 16.065 37.825 ;
        RECT 15.785 37.485 16.065 37.655 ;
        RECT 15.070 37.425 15.245 37.460 ;
        RECT 14.315 37.255 15.245 37.425 ;
        RECT 12.485 37.015 13.715 37.185 ;
        RECT 11.275 36.295 12.285 36.465 ;
        RECT 12.455 36.450 13.205 36.640 ;
        RECT 10.935 35.955 12.060 36.125 ;
        RECT 12.455 35.785 12.625 36.450 ;
        RECT 13.375 36.205 13.715 37.015 ;
        RECT 10.595 35.615 12.625 35.785 ;
        RECT 12.795 35.445 12.965 36.205 ;
        RECT 13.200 35.795 13.715 36.205 ;
        RECT 13.890 36.585 14.060 37.255 ;
        RECT 14.315 37.085 14.485 37.255 ;
        RECT 14.230 36.755 14.485 37.085 ;
        RECT 14.710 36.755 14.905 37.085 ;
        RECT 13.890 35.615 14.225 36.585 ;
        RECT 14.395 35.445 14.565 36.585 ;
        RECT 14.735 35.785 14.905 36.755 ;
        RECT 15.075 36.125 15.245 37.255 ;
        RECT 15.415 36.465 15.585 37.265 ;
        RECT 15.790 36.665 16.065 37.485 ;
        RECT 16.235 36.465 16.425 37.825 ;
        RECT 16.605 37.460 17.115 37.995 ;
        RECT 17.335 37.185 17.580 37.790 ;
        RECT 18.025 37.450 23.370 37.995 ;
        RECT 23.545 37.450 28.890 37.995 ;
        RECT 16.625 37.015 17.855 37.185 ;
        RECT 15.415 36.295 16.425 36.465 ;
        RECT 16.595 36.450 17.345 36.640 ;
        RECT 15.075 35.955 16.200 36.125 ;
        RECT 16.595 35.785 16.765 36.450 ;
        RECT 17.515 36.205 17.855 37.015 ;
        RECT 19.610 36.620 19.950 37.450 ;
        RECT 14.735 35.615 16.765 35.785 ;
        RECT 16.935 35.445 17.105 36.205 ;
        RECT 17.340 35.795 17.855 36.205 ;
        RECT 21.430 35.880 21.780 37.130 ;
        RECT 25.130 36.620 25.470 37.450 ;
        RECT 29.065 37.225 30.735 37.995 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 26.950 35.880 27.300 37.130 ;
        RECT 29.065 36.705 29.815 37.225 ;
        RECT 31.865 37.175 32.095 37.995 ;
        RECT 32.265 37.195 32.595 37.825 ;
        RECT 29.985 36.535 30.735 37.055 ;
        RECT 31.845 36.755 32.175 37.005 ;
        RECT 18.025 35.445 23.370 35.880 ;
        RECT 23.545 35.445 28.890 35.880 ;
        RECT 29.065 35.445 30.735 36.535 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 32.345 36.595 32.595 37.195 ;
        RECT 32.765 37.175 32.975 37.995 ;
        RECT 33.205 37.225 34.875 37.995 ;
        RECT 35.045 37.255 35.385 37.825 ;
        RECT 35.580 37.330 35.750 37.995 ;
        RECT 36.030 37.655 36.250 37.700 ;
        RECT 36.025 37.485 36.250 37.655 ;
        RECT 36.420 37.515 36.865 37.685 ;
        RECT 36.030 37.345 36.250 37.485 ;
        RECT 33.205 36.705 33.955 37.225 ;
        RECT 31.865 35.445 32.095 36.585 ;
        RECT 32.265 35.615 32.595 36.595 ;
        RECT 32.765 35.445 32.975 36.585 ;
        RECT 34.125 36.535 34.875 37.055 ;
        RECT 33.205 35.445 34.875 36.535 ;
        RECT 35.045 36.285 35.220 37.255 ;
        RECT 36.030 37.175 36.525 37.345 ;
        RECT 35.390 36.635 35.560 37.085 ;
        RECT 35.730 36.805 36.180 37.005 ;
        RECT 36.350 36.980 36.525 37.175 ;
        RECT 36.695 36.725 36.865 37.515 ;
        RECT 37.035 37.390 37.285 37.760 ;
        RECT 37.115 37.005 37.285 37.390 ;
        RECT 37.455 37.355 37.705 37.760 ;
        RECT 37.875 37.525 38.045 37.995 ;
        RECT 38.215 37.355 38.555 37.760 ;
        RECT 37.455 37.175 38.555 37.355 ;
        RECT 38.725 37.225 40.395 37.995 ;
        RECT 40.575 37.270 40.905 37.780 ;
        RECT 41.075 37.595 41.405 37.995 ;
        RECT 42.455 37.425 42.785 37.765 ;
        RECT 42.955 37.595 43.285 37.995 ;
        RECT 37.115 36.835 37.310 37.005 ;
        RECT 35.390 36.465 35.785 36.635 ;
        RECT 36.695 36.585 36.970 36.725 ;
        RECT 35.045 35.615 35.305 36.285 ;
        RECT 35.615 36.195 35.785 36.465 ;
        RECT 35.955 36.365 36.970 36.585 ;
        RECT 37.140 36.585 37.310 36.835 ;
        RECT 37.480 36.755 38.040 37.005 ;
        RECT 37.140 36.195 37.695 36.585 ;
        RECT 35.615 36.025 37.695 36.195 ;
        RECT 35.475 35.445 35.805 35.845 ;
        RECT 36.675 35.445 37.075 35.845 ;
        RECT 37.365 35.790 37.695 36.025 ;
        RECT 37.865 35.655 38.040 36.755 ;
        RECT 38.210 36.435 38.555 37.005 ;
        RECT 38.725 36.705 39.475 37.225 ;
        RECT 39.645 36.535 40.395 37.055 ;
        RECT 38.210 35.445 38.555 36.265 ;
        RECT 38.725 35.445 40.395 36.535 ;
        RECT 40.575 36.505 40.765 37.270 ;
        RECT 41.075 37.255 43.440 37.425 ;
        RECT 41.075 37.085 41.245 37.255 ;
        RECT 40.935 36.755 41.245 37.085 ;
        RECT 41.415 36.755 41.720 37.085 ;
        RECT 40.575 35.655 40.905 36.505 ;
        RECT 41.075 35.445 41.325 36.585 ;
        RECT 41.505 36.425 41.720 36.755 ;
        RECT 41.895 36.425 42.180 37.085 ;
        RECT 42.375 36.425 42.640 37.085 ;
        RECT 42.855 36.425 43.100 37.085 ;
        RECT 43.270 36.255 43.440 37.255 ;
        RECT 43.990 37.215 44.490 37.825 ;
        RECT 43.785 36.755 44.135 37.005 ;
        RECT 44.320 36.585 44.490 37.215 ;
        RECT 45.120 37.345 45.450 37.825 ;
        RECT 45.620 37.535 45.845 37.995 ;
        RECT 46.015 37.345 46.345 37.825 ;
        RECT 45.120 37.175 46.345 37.345 ;
        RECT 46.535 37.195 46.785 37.995 ;
        RECT 46.955 37.195 47.295 37.825 ;
        RECT 47.630 37.485 47.870 37.995 ;
        RECT 48.050 37.485 48.330 37.815 ;
        RECT 48.560 37.485 48.775 37.995 ;
        RECT 44.660 36.805 44.990 37.005 ;
        RECT 45.160 36.805 45.490 37.005 ;
        RECT 45.660 36.805 46.080 37.005 ;
        RECT 46.255 36.835 46.950 37.005 ;
        RECT 46.255 36.585 46.425 36.835 ;
        RECT 47.120 36.585 47.295 37.195 ;
        RECT 47.525 36.755 47.880 37.315 ;
        RECT 48.050 36.585 48.220 37.485 ;
        RECT 48.390 36.755 48.655 37.315 ;
        RECT 48.945 37.255 49.560 37.825 ;
        RECT 48.905 36.585 49.075 37.085 ;
        RECT 41.515 36.085 42.805 36.255 ;
        RECT 41.515 35.665 41.765 36.085 ;
        RECT 41.995 35.445 42.325 35.915 ;
        RECT 42.555 35.665 42.805 36.085 ;
        RECT 42.985 36.085 43.440 36.255 ;
        RECT 43.990 36.415 46.425 36.585 ;
        RECT 42.985 35.655 43.315 36.085 ;
        RECT 43.990 35.615 44.320 36.415 ;
        RECT 44.490 35.445 44.820 36.245 ;
        RECT 45.120 35.615 45.450 36.415 ;
        RECT 46.095 35.445 46.345 36.245 ;
        RECT 46.615 35.445 46.785 36.585 ;
        RECT 46.955 35.615 47.295 36.585 ;
        RECT 47.650 36.415 49.075 36.585 ;
        RECT 47.650 36.240 48.040 36.415 ;
        RECT 48.525 35.445 48.855 36.245 ;
        RECT 49.245 36.235 49.560 37.255 ;
        RECT 49.765 37.195 50.460 37.825 ;
        RECT 50.665 37.195 50.975 37.995 ;
        RECT 51.145 37.245 52.355 37.995 ;
        RECT 52.615 37.445 52.785 37.825 ;
        RECT 52.965 37.615 53.295 37.995 ;
        RECT 52.615 37.275 53.280 37.445 ;
        RECT 53.475 37.320 53.735 37.825 ;
        RECT 49.785 36.755 50.120 37.005 ;
        RECT 50.290 36.635 50.460 37.195 ;
        RECT 50.630 36.755 50.965 37.025 ;
        RECT 51.145 36.705 51.665 37.245 ;
        RECT 50.285 36.595 50.460 36.635 ;
        RECT 49.025 35.615 49.560 36.235 ;
        RECT 49.765 35.445 50.025 36.585 ;
        RECT 50.195 35.615 50.525 36.595 ;
        RECT 50.695 35.445 50.975 36.585 ;
        RECT 51.835 36.535 52.355 37.075 ;
        RECT 52.545 36.725 52.885 37.095 ;
        RECT 53.110 37.020 53.280 37.275 ;
        RECT 53.110 36.690 53.385 37.020 ;
        RECT 53.110 36.545 53.280 36.690 ;
        RECT 51.145 35.445 52.355 36.535 ;
        RECT 52.605 36.375 53.280 36.545 ;
        RECT 53.555 36.520 53.735 37.320 ;
        RECT 53.995 37.445 54.165 37.825 ;
        RECT 54.345 37.615 54.675 37.995 ;
        RECT 53.995 37.275 54.660 37.445 ;
        RECT 54.855 37.320 55.115 37.825 ;
        RECT 55.310 37.605 55.640 37.995 ;
        RECT 55.810 37.435 56.035 37.815 ;
        RECT 53.925 36.725 54.265 37.095 ;
        RECT 54.490 37.020 54.660 37.275 ;
        RECT 54.490 36.690 54.765 37.020 ;
        RECT 54.490 36.545 54.660 36.690 ;
        RECT 52.605 35.615 52.785 36.375 ;
        RECT 52.965 35.445 53.295 36.205 ;
        RECT 53.465 35.615 53.735 36.520 ;
        RECT 53.985 36.375 54.660 36.545 ;
        RECT 54.935 36.520 55.115 37.320 ;
        RECT 55.295 36.755 55.535 37.405 ;
        RECT 55.705 37.255 56.035 37.435 ;
        RECT 55.705 36.585 55.880 37.255 ;
        RECT 56.235 37.085 56.465 37.705 ;
        RECT 56.645 37.265 56.945 37.995 ;
        RECT 57.125 37.270 57.415 37.995 ;
        RECT 57.595 37.265 57.895 37.995 ;
        RECT 58.075 37.085 58.305 37.705 ;
        RECT 58.505 37.435 58.730 37.815 ;
        RECT 58.900 37.605 59.230 37.995 ;
        RECT 58.505 37.255 58.835 37.435 ;
        RECT 56.050 36.755 56.465 37.085 ;
        RECT 56.645 36.755 56.940 37.085 ;
        RECT 57.600 36.755 57.895 37.085 ;
        RECT 58.075 36.755 58.490 37.085 ;
        RECT 53.985 35.615 54.165 36.375 ;
        RECT 54.345 35.445 54.675 36.205 ;
        RECT 54.845 35.615 55.115 36.520 ;
        RECT 55.295 36.395 55.880 36.585 ;
        RECT 55.295 35.625 55.570 36.395 ;
        RECT 56.050 36.225 56.945 36.555 ;
        RECT 55.740 36.055 56.945 36.225 ;
        RECT 55.740 35.625 56.070 36.055 ;
        RECT 56.240 35.445 56.435 35.885 ;
        RECT 56.615 35.625 56.945 36.055 ;
        RECT 57.125 35.445 57.415 36.610 ;
        RECT 58.660 36.585 58.835 37.255 ;
        RECT 59.005 36.755 59.245 37.405 ;
        RECT 59.425 37.365 59.765 37.825 ;
        RECT 59.935 37.535 60.105 37.995 ;
        RECT 60.275 37.615 61.445 37.825 ;
        RECT 60.275 37.365 60.525 37.615 ;
        RECT 61.115 37.595 61.445 37.615 ;
        RECT 59.425 37.195 60.525 37.365 ;
        RECT 60.695 37.175 61.555 37.425 ;
        RECT 59.425 36.755 60.185 37.005 ;
        RECT 60.355 36.755 61.105 37.005 ;
        RECT 61.275 36.585 61.555 37.175 ;
        RECT 57.595 36.225 58.490 36.555 ;
        RECT 58.660 36.395 59.245 36.585 ;
        RECT 57.595 36.055 58.800 36.225 ;
        RECT 57.595 35.625 57.925 36.055 ;
        RECT 58.105 35.445 58.300 35.885 ;
        RECT 58.470 35.625 58.800 36.055 ;
        RECT 58.970 35.625 59.245 36.395 ;
        RECT 59.425 35.445 59.685 36.585 ;
        RECT 59.855 36.415 61.555 36.585 ;
        RECT 61.725 37.255 62.085 37.630 ;
        RECT 62.350 37.255 62.520 37.995 ;
        RECT 62.800 37.425 62.970 37.630 ;
        RECT 62.800 37.255 63.340 37.425 ;
        RECT 61.725 36.600 61.980 37.255 ;
        RECT 62.150 36.755 62.500 37.085 ;
        RECT 62.670 36.755 63.000 37.085 ;
        RECT 59.855 35.615 60.185 36.415 ;
        RECT 60.355 35.445 60.525 36.245 ;
        RECT 60.695 35.615 61.025 36.415 ;
        RECT 61.195 35.445 61.450 36.245 ;
        RECT 61.725 35.615 62.065 36.600 ;
        RECT 62.235 36.215 62.500 36.755 ;
        RECT 63.170 36.555 63.340 37.255 ;
        RECT 62.715 36.385 63.340 36.555 ;
        RECT 63.510 36.625 63.680 37.825 ;
        RECT 63.910 37.345 64.240 37.825 ;
        RECT 64.410 37.525 64.580 37.995 ;
        RECT 64.750 37.345 65.080 37.810 ;
        RECT 66.325 37.485 66.630 37.995 ;
        RECT 63.910 37.175 65.080 37.345 ;
        RECT 63.850 36.795 64.420 37.005 ;
        RECT 64.590 36.795 65.235 37.005 ;
        RECT 66.325 36.755 66.640 37.315 ;
        RECT 66.810 37.005 67.060 37.815 ;
        RECT 67.230 37.470 67.490 37.995 ;
        RECT 67.670 37.005 67.920 37.815 ;
        RECT 68.090 37.435 68.350 37.995 ;
        RECT 68.520 37.345 68.780 37.800 ;
        RECT 68.950 37.515 69.210 37.995 ;
        RECT 69.380 37.345 69.640 37.800 ;
        RECT 69.810 37.515 70.070 37.995 ;
        RECT 70.240 37.345 70.500 37.800 ;
        RECT 70.670 37.515 70.915 37.995 ;
        RECT 71.085 37.345 71.360 37.800 ;
        RECT 71.530 37.515 71.775 37.995 ;
        RECT 71.945 37.345 72.205 37.800 ;
        RECT 72.385 37.515 72.635 37.995 ;
        RECT 72.805 37.345 73.065 37.800 ;
        RECT 73.245 37.515 73.495 37.995 ;
        RECT 73.665 37.345 73.925 37.800 ;
        RECT 74.105 37.515 74.365 37.995 ;
        RECT 74.535 37.345 74.795 37.800 ;
        RECT 74.965 37.515 75.265 37.995 ;
        RECT 68.520 37.175 75.265 37.345 ;
        RECT 75.525 37.245 76.735 37.995 ;
        RECT 66.810 36.755 73.930 37.005 ;
        RECT 63.510 36.215 64.215 36.625 ;
        RECT 62.235 36.045 64.215 36.215 ;
        RECT 62.235 35.445 62.645 35.875 ;
        RECT 63.390 35.445 63.720 35.865 ;
        RECT 63.890 35.615 64.215 36.045 ;
        RECT 64.690 35.445 65.020 36.545 ;
        RECT 66.335 35.445 66.630 36.255 ;
        RECT 66.810 35.615 67.055 36.755 ;
        RECT 67.230 35.445 67.490 36.255 ;
        RECT 67.670 35.620 67.920 36.755 ;
        RECT 74.100 36.585 75.265 37.175 ;
        RECT 68.520 36.360 75.265 36.585 ;
        RECT 75.525 36.535 76.045 37.075 ;
        RECT 76.215 36.705 76.735 37.245 ;
        RECT 68.520 36.345 73.925 36.360 ;
        RECT 68.090 35.450 68.350 36.245 ;
        RECT 68.520 35.620 68.780 36.345 ;
        RECT 68.950 35.450 69.210 36.175 ;
        RECT 69.380 35.620 69.640 36.345 ;
        RECT 69.810 35.450 70.070 36.175 ;
        RECT 70.240 35.620 70.500 36.345 ;
        RECT 70.670 35.450 70.930 36.175 ;
        RECT 71.100 35.620 71.360 36.345 ;
        RECT 71.530 35.450 71.775 36.175 ;
        RECT 71.945 35.620 72.205 36.345 ;
        RECT 72.390 35.450 72.635 36.175 ;
        RECT 72.805 35.620 73.065 36.345 ;
        RECT 73.250 35.450 73.495 36.175 ;
        RECT 73.665 35.620 73.925 36.345 ;
        RECT 74.110 35.450 74.365 36.175 ;
        RECT 74.535 35.620 74.825 36.360 ;
        RECT 68.090 35.445 74.365 35.450 ;
        RECT 74.995 35.445 75.265 36.190 ;
        RECT 75.525 35.445 76.735 36.535 ;
        RECT 5.520 35.275 76.820 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 6.985 34.185 8.655 35.275 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 6.985 33.495 7.735 34.015 ;
        RECT 7.905 33.665 8.655 34.185 ;
        RECT 8.825 34.095 9.145 35.275 ;
        RECT 9.315 34.255 9.515 35.045 ;
        RECT 9.840 34.445 10.225 35.105 ;
        RECT 10.620 34.515 11.405 35.275 ;
        RECT 9.815 34.345 10.225 34.445 ;
        RECT 9.315 34.085 9.645 34.255 ;
        RECT 9.815 34.135 11.425 34.345 ;
        RECT 9.465 33.965 9.645 34.085 ;
        RECT 8.825 33.715 9.290 33.915 ;
        RECT 9.465 33.715 9.795 33.965 ;
        RECT 9.965 33.915 10.430 33.965 ;
        RECT 9.965 33.745 10.435 33.915 ;
        RECT 9.965 33.715 10.430 33.745 ;
        RECT 10.625 33.715 10.980 33.965 ;
        RECT 11.150 33.535 11.425 34.135 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 6.985 32.725 8.655 33.495 ;
        RECT 8.825 33.335 10.005 33.505 ;
        RECT 8.825 32.920 9.165 33.335 ;
        RECT 9.335 32.725 9.505 33.165 ;
        RECT 9.675 33.115 10.005 33.335 ;
        RECT 10.175 33.355 11.425 33.535 ;
        RECT 10.175 33.285 10.540 33.355 ;
        RECT 9.675 32.935 10.925 33.115 ;
        RECT 11.195 32.725 11.365 33.185 ;
        RECT 11.595 33.005 11.875 35.105 ;
        RECT 12.045 34.840 17.390 35.275 ;
        RECT 13.630 33.270 13.970 34.100 ;
        RECT 15.450 33.590 15.800 34.840 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 19.005 34.135 19.215 35.275 ;
        RECT 19.385 34.125 19.715 35.105 ;
        RECT 19.885 34.135 20.115 35.275 ;
        RECT 20.325 34.185 21.535 35.275 ;
        RECT 12.045 32.725 17.390 33.270 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 19.005 32.725 19.215 33.545 ;
        RECT 19.385 33.525 19.635 34.125 ;
        RECT 19.805 33.715 20.135 33.965 ;
        RECT 19.385 32.895 19.715 33.525 ;
        RECT 19.885 32.725 20.115 33.545 ;
        RECT 20.325 33.475 20.845 34.015 ;
        RECT 21.015 33.645 21.535 34.185 ;
        RECT 21.710 34.135 22.045 35.105 ;
        RECT 22.215 34.135 22.385 35.275 ;
        RECT 22.555 34.935 24.585 35.105 ;
        RECT 20.325 32.725 21.535 33.475 ;
        RECT 21.710 33.465 21.880 34.135 ;
        RECT 22.555 33.965 22.725 34.935 ;
        RECT 22.050 33.635 22.305 33.965 ;
        RECT 22.530 33.635 22.725 33.965 ;
        RECT 22.895 34.595 24.020 34.765 ;
        RECT 22.135 33.465 22.305 33.635 ;
        RECT 22.895 33.465 23.065 34.595 ;
        RECT 21.710 32.895 21.965 33.465 ;
        RECT 22.135 33.295 23.065 33.465 ;
        RECT 23.235 34.255 24.245 34.425 ;
        RECT 23.235 33.455 23.405 34.255 ;
        RECT 22.890 33.260 23.065 33.295 ;
        RECT 22.135 32.725 22.465 33.125 ;
        RECT 22.890 32.895 23.420 33.260 ;
        RECT 23.610 33.235 23.885 34.055 ;
        RECT 23.605 33.065 23.885 33.235 ;
        RECT 23.610 32.895 23.885 33.065 ;
        RECT 24.055 32.895 24.245 34.255 ;
        RECT 24.415 34.270 24.585 34.935 ;
        RECT 24.755 34.515 24.925 35.275 ;
        RECT 25.160 34.515 25.675 34.925 ;
        RECT 24.415 34.080 25.165 34.270 ;
        RECT 25.335 33.705 25.675 34.515 ;
        RECT 25.845 34.135 26.105 35.275 ;
        RECT 26.275 34.125 26.605 35.105 ;
        RECT 26.775 34.135 27.055 35.275 ;
        RECT 27.225 34.185 30.735 35.275 ;
        RECT 25.865 33.715 26.200 33.965 ;
        RECT 24.445 33.535 25.675 33.705 ;
        RECT 24.425 32.725 24.935 33.260 ;
        RECT 25.155 32.930 25.400 33.535 ;
        RECT 26.370 33.525 26.540 34.125 ;
        RECT 26.710 33.695 27.045 33.965 ;
        RECT 25.845 32.895 26.540 33.525 ;
        RECT 26.745 32.725 27.055 33.525 ;
        RECT 27.225 33.495 28.875 34.015 ;
        RECT 29.045 33.665 30.735 34.185 ;
        RECT 30.910 34.325 31.175 35.095 ;
        RECT 31.345 34.555 31.675 35.275 ;
        RECT 31.865 34.735 32.125 35.095 ;
        RECT 32.295 34.905 32.625 35.275 ;
        RECT 32.795 34.735 33.055 35.095 ;
        RECT 31.865 34.505 33.055 34.735 ;
        RECT 33.625 34.325 33.915 35.095 ;
        RECT 34.125 34.840 39.470 35.275 ;
        RECT 27.225 32.725 30.735 33.495 ;
        RECT 30.910 32.905 31.245 34.325 ;
        RECT 31.420 34.145 33.915 34.325 ;
        RECT 31.420 33.455 31.645 34.145 ;
        RECT 31.845 33.635 32.125 33.965 ;
        RECT 32.305 33.635 32.880 33.965 ;
        RECT 33.060 33.635 33.495 33.965 ;
        RECT 33.675 33.635 33.945 33.965 ;
        RECT 31.420 33.265 33.905 33.455 ;
        RECT 35.710 33.270 36.050 34.100 ;
        RECT 37.530 33.590 37.880 34.840 ;
        RECT 39.645 34.185 43.155 35.275 ;
        RECT 39.645 33.495 41.295 34.015 ;
        RECT 41.465 33.665 43.155 34.185 ;
        RECT 44.245 34.110 44.535 35.275 ;
        RECT 44.705 34.135 44.980 35.105 ;
        RECT 45.190 34.475 45.470 35.275 ;
        RECT 45.640 34.765 47.255 35.095 ;
        RECT 45.640 34.425 46.815 34.595 ;
        RECT 45.640 34.305 45.810 34.425 ;
        RECT 45.150 34.135 45.810 34.305 ;
        RECT 31.425 32.725 32.170 33.095 ;
        RECT 32.735 32.905 32.990 33.265 ;
        RECT 33.170 32.725 33.500 33.095 ;
        RECT 33.680 32.905 33.905 33.265 ;
        RECT 34.125 32.725 39.470 33.270 ;
        RECT 39.645 32.725 43.155 33.495 ;
        RECT 44.245 32.725 44.535 33.450 ;
        RECT 44.705 33.400 44.875 34.135 ;
        RECT 45.150 33.965 45.320 34.135 ;
        RECT 46.070 33.965 46.315 34.255 ;
        RECT 46.485 34.135 46.815 34.425 ;
        RECT 47.075 33.965 47.245 34.525 ;
        RECT 47.495 34.135 47.755 35.275 ;
        RECT 48.855 34.295 49.105 35.105 ;
        RECT 49.275 34.935 51.385 35.105 ;
        RECT 49.275 34.465 49.525 34.935 ;
        RECT 49.695 34.295 50.025 34.765 ;
        RECT 50.195 34.465 50.365 34.935 ;
        RECT 50.535 34.295 50.920 34.765 ;
        RECT 48.855 34.125 50.920 34.295 ;
        RECT 51.135 34.295 51.385 34.935 ;
        RECT 51.555 34.465 51.725 35.275 ;
        RECT 51.895 34.295 52.225 35.105 ;
        RECT 52.395 34.465 52.565 35.275 ;
        RECT 52.735 34.295 53.065 35.105 ;
        RECT 51.135 34.125 53.065 34.295 ;
        RECT 45.045 33.635 45.320 33.965 ;
        RECT 45.490 33.635 46.315 33.965 ;
        RECT 46.530 33.635 47.245 33.965 ;
        RECT 47.415 33.715 47.750 33.965 ;
        RECT 48.905 33.745 49.540 33.915 ;
        RECT 49.825 33.745 50.460 33.915 ;
        RECT 48.910 33.715 49.540 33.745 ;
        RECT 49.830 33.715 50.460 33.745 ;
        RECT 45.150 33.465 45.320 33.635 ;
        RECT 46.995 33.545 47.245 33.635 ;
        RECT 44.705 33.055 44.980 33.400 ;
        RECT 45.150 33.295 46.815 33.465 ;
        RECT 45.170 32.725 45.545 33.125 ;
        RECT 45.715 32.945 45.885 33.295 ;
        RECT 46.055 32.725 46.385 33.125 ;
        RECT 46.555 32.895 46.815 33.295 ;
        RECT 46.995 33.125 47.325 33.545 ;
        RECT 47.495 32.725 47.755 33.545 ;
        RECT 48.855 33.320 49.945 33.490 ;
        RECT 50.630 33.485 50.920 34.125 ;
        RECT 51.205 33.715 51.860 33.915 ;
        RECT 52.125 33.745 53.260 33.915 ;
        RECT 52.150 33.715 53.260 33.745 ;
        RECT 48.855 32.895 49.105 33.320 ;
        RECT 49.275 32.725 49.605 33.150 ;
        RECT 49.775 33.145 49.945 33.320 ;
        RECT 50.115 33.315 51.805 33.485 ;
        RECT 51.975 33.320 53.135 33.490 ;
        RECT 51.975 33.145 52.145 33.320 ;
        RECT 49.775 32.895 50.865 33.145 ;
        RECT 51.055 32.895 52.145 33.145 ;
        RECT 52.315 32.725 52.645 33.150 ;
        RECT 52.815 32.895 53.135 33.320 ;
        RECT 53.905 32.895 54.655 35.105 ;
        RECT 54.835 34.305 55.165 35.090 ;
        RECT 54.835 34.135 55.515 34.305 ;
        RECT 55.695 34.135 56.025 35.275 ;
        RECT 54.825 33.715 55.175 33.965 ;
        RECT 55.345 33.535 55.515 34.135 ;
        RECT 56.210 34.125 56.470 35.275 ;
        RECT 56.645 34.200 56.900 35.105 ;
        RECT 57.070 34.515 57.400 35.275 ;
        RECT 57.615 34.345 57.785 35.105 ;
        RECT 55.685 33.715 56.035 33.965 ;
        RECT 54.845 32.725 55.085 33.535 ;
        RECT 55.255 32.895 55.585 33.535 ;
        RECT 55.755 32.725 56.025 33.535 ;
        RECT 56.210 32.725 56.470 33.565 ;
        RECT 56.645 33.470 56.815 34.200 ;
        RECT 57.070 34.175 57.785 34.345 ;
        RECT 58.135 34.345 58.305 35.105 ;
        RECT 58.520 34.515 58.850 35.275 ;
        RECT 58.135 34.175 58.850 34.345 ;
        RECT 59.020 34.200 59.275 35.105 ;
        RECT 57.070 33.965 57.240 34.175 ;
        RECT 56.985 33.635 57.240 33.965 ;
        RECT 56.645 32.895 56.900 33.470 ;
        RECT 57.070 33.445 57.240 33.635 ;
        RECT 57.520 33.625 57.875 33.995 ;
        RECT 58.045 33.625 58.400 33.995 ;
        RECT 58.680 33.965 58.850 34.175 ;
        RECT 58.680 33.635 58.935 33.965 ;
        RECT 58.680 33.445 58.850 33.635 ;
        RECT 59.105 33.470 59.275 34.200 ;
        RECT 59.450 34.125 59.710 35.275 ;
        RECT 60.345 34.720 60.950 35.275 ;
        RECT 61.125 34.765 61.605 35.105 ;
        RECT 61.775 34.730 62.030 35.275 ;
        RECT 60.345 34.620 60.960 34.720 ;
        RECT 60.775 34.595 60.960 34.620 ;
        RECT 60.345 34.000 60.605 34.450 ;
        RECT 60.775 34.350 61.105 34.595 ;
        RECT 61.275 34.275 62.030 34.525 ;
        RECT 62.200 34.405 62.475 35.105 ;
        RECT 63.565 34.765 64.755 35.055 ;
        RECT 61.260 34.240 62.030 34.275 ;
        RECT 61.245 34.230 62.030 34.240 ;
        RECT 61.240 34.215 62.135 34.230 ;
        RECT 61.220 34.200 62.135 34.215 ;
        RECT 61.200 34.190 62.135 34.200 ;
        RECT 61.175 34.180 62.135 34.190 ;
        RECT 61.105 34.150 62.135 34.180 ;
        RECT 61.085 34.120 62.135 34.150 ;
        RECT 61.065 34.090 62.135 34.120 ;
        RECT 61.035 34.065 62.135 34.090 ;
        RECT 61.000 34.030 62.135 34.065 ;
        RECT 60.970 34.025 62.135 34.030 ;
        RECT 60.970 34.020 61.360 34.025 ;
        RECT 60.970 34.010 61.335 34.020 ;
        RECT 60.970 34.005 61.320 34.010 ;
        RECT 60.970 34.000 61.305 34.005 ;
        RECT 60.345 33.995 61.305 34.000 ;
        RECT 60.345 33.985 61.295 33.995 ;
        RECT 60.345 33.980 61.285 33.985 ;
        RECT 60.345 33.970 61.275 33.980 ;
        RECT 60.345 33.960 61.270 33.970 ;
        RECT 60.345 33.955 61.265 33.960 ;
        RECT 60.345 33.940 61.255 33.955 ;
        RECT 60.345 33.925 61.250 33.940 ;
        RECT 60.345 33.900 61.240 33.925 ;
        RECT 60.345 33.830 61.235 33.900 ;
        RECT 57.070 33.275 57.785 33.445 ;
        RECT 57.070 32.725 57.400 33.105 ;
        RECT 57.615 32.895 57.785 33.275 ;
        RECT 58.135 33.275 58.850 33.445 ;
        RECT 58.135 32.895 58.305 33.275 ;
        RECT 58.520 32.725 58.850 33.105 ;
        RECT 59.020 32.895 59.275 33.470 ;
        RECT 59.450 32.725 59.710 33.565 ;
        RECT 60.345 33.275 60.895 33.660 ;
        RECT 61.065 33.105 61.235 33.830 ;
        RECT 60.345 32.935 61.235 33.105 ;
        RECT 61.405 33.430 61.735 33.855 ;
        RECT 61.905 33.630 62.135 34.025 ;
        RECT 61.405 32.945 61.625 33.430 ;
        RECT 62.305 33.375 62.475 34.405 ;
        RECT 63.585 34.425 64.755 34.595 ;
        RECT 64.925 34.475 65.205 35.275 ;
        RECT 63.585 34.135 63.910 34.425 ;
        RECT 64.585 34.305 64.755 34.425 ;
        RECT 64.080 33.965 64.275 34.255 ;
        RECT 64.585 34.135 65.245 34.305 ;
        RECT 65.415 34.135 65.690 35.105 ;
        RECT 65.945 34.345 66.125 35.105 ;
        RECT 66.305 34.515 66.635 35.275 ;
        RECT 65.945 34.175 66.620 34.345 ;
        RECT 66.805 34.200 67.075 35.105 ;
        RECT 67.300 34.405 67.585 35.275 ;
        RECT 67.755 34.645 68.015 35.105 ;
        RECT 68.190 34.815 68.445 35.275 ;
        RECT 68.615 34.645 68.875 35.105 ;
        RECT 67.755 34.475 68.875 34.645 ;
        RECT 69.045 34.475 69.355 35.275 ;
        RECT 67.755 34.225 68.015 34.475 ;
        RECT 69.525 34.305 69.835 35.105 ;
        RECT 65.075 33.965 65.245 34.135 ;
        RECT 63.565 33.635 63.910 33.965 ;
        RECT 64.080 33.635 64.905 33.965 ;
        RECT 65.075 33.635 65.350 33.965 ;
        RECT 65.075 33.465 65.245 33.635 ;
        RECT 61.795 32.725 62.045 33.265 ;
        RECT 62.215 32.895 62.475 33.375 ;
        RECT 63.580 33.295 65.245 33.465 ;
        RECT 65.520 33.400 65.690 34.135 ;
        RECT 66.450 34.030 66.620 34.175 ;
        RECT 65.885 33.625 66.225 33.995 ;
        RECT 66.450 33.700 66.725 34.030 ;
        RECT 66.450 33.445 66.620 33.700 ;
        RECT 63.580 32.945 63.835 33.295 ;
        RECT 64.005 32.725 64.335 33.125 ;
        RECT 64.505 32.945 64.675 33.295 ;
        RECT 64.845 32.725 65.225 33.125 ;
        RECT 65.415 33.055 65.690 33.400 ;
        RECT 65.955 33.275 66.620 33.445 ;
        RECT 66.895 33.400 67.075 34.200 ;
        RECT 65.955 32.895 66.125 33.275 ;
        RECT 66.305 32.725 66.635 33.105 ;
        RECT 66.815 32.895 67.075 33.400 ;
        RECT 67.260 34.055 68.015 34.225 ;
        RECT 68.805 34.135 69.835 34.305 ;
        RECT 67.260 33.545 67.665 34.055 ;
        RECT 68.805 33.885 68.975 34.135 ;
        RECT 67.835 33.715 68.975 33.885 ;
        RECT 67.260 33.375 68.910 33.545 ;
        RECT 69.145 33.395 69.495 33.965 ;
        RECT 67.305 32.725 67.585 33.205 ;
        RECT 67.755 32.985 68.015 33.375 ;
        RECT 68.190 32.725 68.445 33.205 ;
        RECT 68.615 32.985 68.910 33.375 ;
        RECT 69.665 33.225 69.835 34.135 ;
        RECT 70.005 34.110 70.295 35.275 ;
        RECT 70.545 34.345 70.725 35.105 ;
        RECT 70.905 34.515 71.235 35.275 ;
        RECT 70.545 34.175 71.220 34.345 ;
        RECT 71.405 34.200 71.675 35.105 ;
        RECT 71.975 34.935 74.025 35.105 ;
        RECT 71.975 34.435 72.225 34.935 ;
        RECT 72.395 34.265 72.605 34.765 ;
        RECT 72.815 34.435 73.025 34.935 ;
        RECT 73.355 34.265 73.605 34.765 ;
        RECT 73.775 34.435 74.025 34.935 ;
        RECT 74.195 34.265 74.445 35.105 ;
        RECT 74.615 34.435 74.865 35.275 ;
        RECT 75.035 34.265 75.290 35.105 ;
        RECT 71.050 34.030 71.220 34.175 ;
        RECT 70.485 33.625 70.825 33.995 ;
        RECT 71.050 33.700 71.325 34.030 ;
        RECT 69.090 32.725 69.365 33.205 ;
        RECT 69.535 32.895 69.835 33.225 ;
        RECT 70.005 32.725 70.295 33.450 ;
        RECT 71.050 33.445 71.220 33.700 ;
        RECT 70.555 33.275 71.220 33.445 ;
        RECT 71.495 33.400 71.675 34.200 ;
        RECT 70.555 32.895 70.725 33.275 ;
        RECT 70.905 32.725 71.235 33.105 ;
        RECT 71.415 32.895 71.675 33.400 ;
        RECT 71.845 34.095 72.605 34.265 ;
        RECT 71.845 33.545 72.305 34.095 ;
        RECT 72.800 33.925 73.065 34.265 ;
        RECT 73.355 34.095 75.290 34.265 ;
        RECT 75.525 34.185 76.735 35.275 ;
        RECT 72.475 33.715 73.065 33.925 ;
        RECT 73.255 33.715 74.305 33.925 ;
        RECT 74.475 33.715 75.305 33.925 ;
        RECT 75.525 33.645 76.045 34.185 ;
        RECT 71.845 33.365 74.905 33.545 ;
        RECT 71.895 32.725 72.185 33.195 ;
        RECT 72.355 32.895 72.685 33.365 ;
        RECT 72.855 32.725 73.565 33.195 ;
        RECT 73.735 32.895 74.065 33.365 ;
        RECT 74.235 32.725 74.405 33.195 ;
        RECT 74.575 32.895 74.905 33.365 ;
        RECT 75.075 32.725 75.350 33.545 ;
        RECT 76.215 33.475 76.735 34.015 ;
        RECT 75.525 32.725 76.735 33.475 ;
        RECT 5.520 32.555 76.820 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.990 31.715 7.250 32.555 ;
        RECT 7.425 31.810 7.680 32.385 ;
        RECT 7.850 32.175 8.180 32.555 ;
        RECT 8.395 32.005 8.565 32.385 ;
        RECT 7.850 31.835 8.565 32.005 ;
        RECT 8.825 32.055 9.085 32.385 ;
        RECT 9.295 32.075 9.570 32.555 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 6.990 30.005 7.250 31.155 ;
        RECT 7.425 31.080 7.595 31.810 ;
        RECT 7.850 31.645 8.020 31.835 ;
        RECT 7.765 31.315 8.020 31.645 ;
        RECT 7.850 31.105 8.020 31.315 ;
        RECT 8.300 31.285 8.655 31.655 ;
        RECT 8.825 31.145 8.995 32.055 ;
        RECT 9.780 31.985 9.985 32.385 ;
        RECT 10.155 32.155 10.490 32.555 ;
        RECT 9.165 31.315 9.525 31.895 ;
        RECT 9.780 31.815 10.465 31.985 ;
        RECT 9.705 31.145 9.955 31.645 ;
        RECT 7.425 30.175 7.680 31.080 ;
        RECT 7.850 30.935 8.565 31.105 ;
        RECT 7.850 30.005 8.180 30.765 ;
        RECT 8.395 30.175 8.565 30.935 ;
        RECT 8.825 30.975 9.955 31.145 ;
        RECT 8.825 30.205 9.095 30.975 ;
        RECT 10.125 30.785 10.465 31.815 ;
        RECT 9.265 30.005 9.595 30.785 ;
        RECT 9.800 30.610 10.465 30.785 ;
        RECT 10.665 31.880 10.925 32.385 ;
        RECT 11.105 32.175 11.435 32.555 ;
        RECT 11.615 32.005 11.785 32.385 ;
        RECT 10.665 31.080 10.835 31.880 ;
        RECT 11.120 31.835 11.785 32.005 ;
        RECT 11.120 31.580 11.290 31.835 ;
        RECT 12.045 31.785 15.555 32.555 ;
        RECT 11.005 31.250 11.290 31.580 ;
        RECT 11.525 31.285 11.855 31.655 ;
        RECT 12.045 31.265 13.695 31.785 ;
        RECT 16.645 31.755 16.955 32.555 ;
        RECT 17.160 31.755 17.855 32.385 ;
        RECT 18.025 31.945 18.365 32.360 ;
        RECT 18.535 32.115 18.705 32.555 ;
        RECT 18.875 32.165 20.125 32.345 ;
        RECT 18.875 31.945 19.205 32.165 ;
        RECT 20.395 32.095 20.565 32.555 ;
        RECT 18.025 31.775 19.205 31.945 ;
        RECT 19.375 31.925 19.740 31.995 ;
        RECT 17.160 31.705 17.335 31.755 ;
        RECT 19.375 31.745 20.625 31.925 ;
        RECT 11.120 31.105 11.290 31.250 ;
        RECT 9.800 30.205 9.985 30.610 ;
        RECT 10.155 30.005 10.490 30.430 ;
        RECT 10.665 30.175 10.935 31.080 ;
        RECT 11.120 30.935 11.785 31.105 ;
        RECT 13.865 31.095 15.555 31.615 ;
        RECT 16.655 31.315 16.990 31.585 ;
        RECT 17.160 31.155 17.330 31.705 ;
        RECT 17.500 31.315 17.835 31.565 ;
        RECT 18.025 31.365 18.490 31.565 ;
        RECT 18.665 31.315 18.995 31.565 ;
        RECT 19.165 31.535 19.630 31.565 ;
        RECT 19.165 31.365 19.635 31.535 ;
        RECT 19.165 31.315 19.630 31.365 ;
        RECT 19.825 31.315 20.180 31.565 ;
        RECT 18.665 31.195 18.845 31.315 ;
        RECT 11.105 30.005 11.435 30.765 ;
        RECT 11.615 30.175 11.785 30.935 ;
        RECT 12.045 30.005 15.555 31.095 ;
        RECT 16.645 30.005 16.925 31.145 ;
        RECT 17.095 30.175 17.425 31.155 ;
        RECT 17.595 30.005 17.855 31.145 ;
        RECT 18.025 30.005 18.345 31.185 ;
        RECT 18.515 31.025 18.845 31.195 ;
        RECT 20.350 31.145 20.625 31.745 ;
        RECT 18.515 30.235 18.715 31.025 ;
        RECT 19.015 30.935 20.625 31.145 ;
        RECT 19.015 30.835 19.425 30.935 ;
        RECT 19.040 30.175 19.425 30.835 ;
        RECT 19.820 30.005 20.605 30.765 ;
        RECT 20.795 30.175 21.075 32.275 ;
        RECT 21.250 31.815 21.505 32.385 ;
        RECT 21.675 32.155 22.005 32.555 ;
        RECT 22.430 32.020 22.960 32.385 ;
        RECT 22.430 31.985 22.605 32.020 ;
        RECT 21.675 31.815 22.605 31.985 ;
        RECT 21.250 31.145 21.420 31.815 ;
        RECT 21.675 31.645 21.845 31.815 ;
        RECT 21.590 31.315 21.845 31.645 ;
        RECT 22.070 31.315 22.265 31.645 ;
        RECT 21.250 30.175 21.585 31.145 ;
        RECT 21.755 30.005 21.925 31.145 ;
        RECT 22.095 30.345 22.265 31.315 ;
        RECT 22.435 30.685 22.605 31.815 ;
        RECT 22.775 31.025 22.945 31.825 ;
        RECT 23.150 31.535 23.425 32.385 ;
        RECT 23.145 31.365 23.425 31.535 ;
        RECT 23.150 31.225 23.425 31.365 ;
        RECT 23.595 31.025 23.785 32.385 ;
        RECT 23.965 32.020 24.475 32.555 ;
        RECT 24.695 31.745 24.940 32.350 ;
        RECT 25.585 31.925 25.915 32.285 ;
        RECT 26.535 32.095 26.785 32.555 ;
        RECT 26.955 32.095 27.515 32.385 ;
        RECT 23.985 31.575 25.215 31.745 ;
        RECT 25.585 31.735 26.975 31.925 ;
        RECT 22.775 30.855 23.785 31.025 ;
        RECT 23.955 31.010 24.705 31.200 ;
        RECT 22.435 30.515 23.560 30.685 ;
        RECT 23.955 30.345 24.125 31.010 ;
        RECT 24.875 30.765 25.215 31.575 ;
        RECT 26.805 31.645 26.975 31.735 ;
        RECT 25.400 31.315 26.075 31.565 ;
        RECT 26.295 31.315 26.635 31.565 ;
        RECT 26.805 31.315 27.095 31.645 ;
        RECT 25.400 30.955 25.665 31.315 ;
        RECT 26.805 31.065 26.975 31.315 ;
        RECT 22.095 30.175 24.125 30.345 ;
        RECT 24.295 30.005 24.465 30.765 ;
        RECT 24.700 30.355 25.215 30.765 ;
        RECT 26.035 30.895 26.975 31.065 ;
        RECT 25.585 30.005 25.865 30.675 ;
        RECT 26.035 30.345 26.335 30.895 ;
        RECT 27.265 30.725 27.515 32.095 ;
        RECT 28.310 32.045 28.550 32.555 ;
        RECT 28.730 32.045 29.010 32.375 ;
        RECT 29.240 32.045 29.455 32.555 ;
        RECT 28.205 31.315 28.560 31.875 ;
        RECT 28.730 31.145 28.900 32.045 ;
        RECT 29.070 31.315 29.335 31.875 ;
        RECT 29.625 31.815 30.240 32.385 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 29.585 31.145 29.755 31.645 ;
        RECT 28.330 30.975 29.755 31.145 ;
        RECT 28.330 30.800 28.720 30.975 ;
        RECT 26.535 30.005 26.865 30.725 ;
        RECT 27.055 30.175 27.515 30.725 ;
        RECT 29.205 30.005 29.535 30.805 ;
        RECT 29.925 30.795 30.240 31.815 ;
        RECT 31.825 31.735 32.510 32.375 ;
        RECT 32.680 31.735 32.850 32.555 ;
        RECT 33.020 31.905 33.350 32.370 ;
        RECT 33.520 32.085 33.690 32.555 ;
        RECT 33.950 32.165 35.135 32.335 ;
        RECT 35.305 31.995 35.635 32.385 ;
        RECT 34.335 31.905 34.720 31.995 ;
        RECT 33.020 31.735 34.720 31.905 ;
        RECT 35.125 31.815 35.635 31.995 ;
        RECT 35.975 31.835 36.305 32.555 ;
        RECT 36.850 32.155 38.465 32.325 ;
        RECT 38.635 32.155 38.965 32.555 ;
        RECT 38.295 31.985 38.465 32.155 ;
        RECT 39.135 32.080 39.470 32.340 ;
        RECT 29.705 30.175 30.240 30.795 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 31.825 30.765 32.075 31.735 ;
        RECT 32.245 31.355 32.580 31.565 ;
        RECT 32.750 31.355 33.200 31.565 ;
        RECT 33.390 31.355 33.875 31.565 ;
        RECT 32.410 31.185 32.580 31.355 ;
        RECT 33.500 31.195 33.875 31.355 ;
        RECT 34.065 31.315 34.445 31.565 ;
        RECT 34.625 31.355 34.955 31.565 ;
        RECT 32.410 31.015 33.330 31.185 ;
        RECT 31.825 30.175 32.490 30.765 ;
        RECT 32.660 30.005 32.990 30.845 ;
        RECT 33.160 30.765 33.330 31.015 ;
        RECT 33.500 31.025 33.895 31.195 ;
        RECT 33.500 30.935 33.875 31.025 ;
        RECT 34.065 30.935 34.385 31.315 ;
        RECT 35.125 31.185 35.295 31.815 ;
        RECT 35.465 31.355 35.795 31.645 ;
        RECT 36.030 31.535 36.380 31.645 ;
        RECT 36.025 31.365 36.380 31.535 ;
        RECT 36.030 31.315 36.380 31.365 ;
        RECT 36.690 31.315 37.110 31.980 ;
        RECT 37.280 31.535 37.570 31.975 ;
        RECT 37.760 31.535 38.030 31.975 ;
        RECT 38.295 31.815 38.855 31.985 ;
        RECT 38.685 31.645 38.855 31.815 ;
        RECT 38.240 31.535 38.490 31.645 ;
        RECT 37.280 31.365 37.575 31.535 ;
        RECT 37.760 31.365 38.035 31.535 ;
        RECT 38.240 31.365 38.495 31.535 ;
        RECT 37.280 31.315 37.570 31.365 ;
        RECT 37.760 31.315 38.030 31.365 ;
        RECT 38.240 31.315 38.490 31.365 ;
        RECT 38.685 31.315 38.990 31.645 ;
        RECT 34.555 31.015 35.640 31.185 ;
        RECT 36.030 31.025 36.235 31.315 ;
        RECT 38.685 31.145 38.855 31.315 ;
        RECT 34.555 30.765 34.725 31.015 ;
        RECT 33.160 30.595 34.725 30.765 ;
        RECT 33.500 30.175 34.305 30.595 ;
        RECT 34.895 30.005 35.145 30.845 ;
        RECT 35.340 30.175 35.640 31.015 ;
        RECT 36.485 30.975 38.855 31.145 ;
        RECT 36.055 30.345 36.225 30.845 ;
        RECT 36.485 30.515 36.655 30.975 ;
        RECT 36.885 30.595 38.310 30.765 ;
        RECT 36.885 30.345 37.215 30.595 ;
        RECT 36.055 30.175 37.215 30.345 ;
        RECT 37.440 30.005 37.770 30.425 ;
        RECT 38.025 30.175 38.310 30.595 ;
        RECT 38.555 30.005 38.885 30.805 ;
        RECT 39.215 30.725 39.470 32.080 ;
        RECT 39.645 31.785 42.235 32.555 ;
        RECT 42.845 31.835 43.185 32.555 ;
        RECT 39.645 31.265 40.855 31.785 ;
        RECT 43.375 31.645 43.575 32.225 ;
        RECT 43.835 31.875 44.135 32.295 ;
        RECT 44.375 32.215 44.625 32.345 ;
        RECT 44.305 32.045 44.625 32.215 ;
        RECT 45.115 32.175 45.445 32.555 ;
        RECT 41.025 31.095 42.235 31.615 ;
        RECT 42.790 31.315 43.205 31.625 ;
        RECT 43.375 31.315 43.735 31.645 ;
        RECT 43.945 31.565 44.135 31.875 ;
        RECT 44.375 32.005 44.625 32.045 ;
        RECT 44.375 31.835 45.025 32.005 ;
        RECT 43.945 31.385 44.310 31.565 ;
        RECT 44.515 31.215 44.685 31.645 ;
        RECT 39.135 30.215 39.470 30.725 ;
        RECT 39.645 30.005 42.235 31.095 ;
        RECT 42.845 30.005 43.185 31.145 ;
        RECT 44.285 31.025 44.685 31.215 ;
        RECT 43.355 30.855 43.525 30.895 ;
        RECT 44.855 30.855 45.025 31.835 ;
        RECT 45.625 31.785 49.135 32.555 ;
        RECT 50.245 31.825 50.535 32.555 ;
        RECT 45.195 31.315 45.455 31.645 ;
        RECT 45.625 31.265 47.275 31.785 ;
        RECT 47.445 31.095 49.135 31.615 ;
        RECT 50.235 31.315 50.535 31.645 ;
        RECT 50.715 31.625 50.945 32.265 ;
        RECT 51.125 32.005 51.435 32.375 ;
        RECT 51.615 32.185 52.285 32.555 ;
        RECT 51.125 31.805 52.355 32.005 ;
        RECT 50.715 31.315 51.240 31.625 ;
        RECT 51.420 31.315 51.885 31.625 ;
        RECT 52.065 31.135 52.355 31.805 ;
        RECT 43.355 30.685 44.445 30.855 ;
        RECT 43.355 30.175 43.525 30.685 ;
        RECT 43.735 30.005 43.985 30.505 ;
        RECT 44.195 30.385 44.445 30.685 ;
        RECT 44.675 30.555 45.025 30.855 ;
        RECT 45.195 30.385 45.455 30.805 ;
        RECT 44.195 30.175 45.455 30.385 ;
        RECT 45.625 30.005 49.135 31.095 ;
        RECT 50.245 30.895 51.405 31.135 ;
        RECT 50.245 30.185 50.505 30.895 ;
        RECT 50.675 30.005 51.005 30.715 ;
        RECT 51.175 30.185 51.405 30.895 ;
        RECT 51.585 30.915 52.355 31.135 ;
        RECT 51.585 30.185 51.855 30.915 ;
        RECT 52.035 30.005 52.375 30.735 ;
        RECT 52.545 30.185 52.805 32.375 ;
        RECT 52.995 32.055 53.325 32.555 ;
        RECT 53.525 31.985 53.695 32.335 ;
        RECT 53.895 32.155 54.225 32.555 ;
        RECT 54.395 31.985 54.565 32.335 ;
        RECT 54.735 32.155 55.115 32.555 ;
        RECT 52.990 31.315 53.340 31.885 ;
        RECT 53.525 31.815 55.135 31.985 ;
        RECT 55.305 31.880 55.575 32.225 ;
        RECT 54.965 31.645 55.135 31.815 ;
        RECT 52.990 30.855 53.310 31.145 ;
        RECT 53.510 31.025 54.220 31.645 ;
        RECT 54.390 31.315 54.795 31.645 ;
        RECT 54.965 31.315 55.235 31.645 ;
        RECT 54.965 31.145 55.135 31.315 ;
        RECT 55.405 31.145 55.575 31.880 ;
        RECT 55.745 31.805 56.955 32.555 ;
        RECT 57.125 31.830 57.415 32.555 ;
        RECT 55.745 31.265 56.265 31.805 ;
        RECT 54.410 30.975 55.135 31.145 ;
        RECT 54.410 30.855 54.580 30.975 ;
        RECT 52.990 30.685 54.580 30.855 ;
        RECT 52.990 30.225 54.645 30.515 ;
        RECT 54.815 30.005 55.095 30.805 ;
        RECT 55.305 30.175 55.575 31.145 ;
        RECT 56.435 31.095 56.955 31.635 ;
        RECT 55.745 30.005 56.955 31.095 ;
        RECT 57.125 30.005 57.415 31.170 ;
        RECT 57.585 30.175 57.865 32.275 ;
        RECT 58.095 32.095 58.265 32.555 ;
        RECT 58.535 32.165 59.785 32.345 ;
        RECT 58.920 31.925 59.285 31.995 ;
        RECT 58.035 31.745 59.285 31.925 ;
        RECT 59.455 31.945 59.785 32.165 ;
        RECT 59.955 32.115 60.125 32.555 ;
        RECT 60.295 31.945 60.635 32.360 ;
        RECT 59.455 31.775 60.635 31.945 ;
        RECT 60.805 31.905 61.065 32.385 ;
        RECT 61.235 32.015 61.485 32.555 ;
        RECT 58.035 31.145 58.310 31.745 ;
        RECT 58.480 31.315 58.835 31.565 ;
        RECT 59.030 31.535 59.495 31.565 ;
        RECT 59.025 31.365 59.495 31.535 ;
        RECT 59.030 31.315 59.495 31.365 ;
        RECT 59.665 31.315 59.995 31.565 ;
        RECT 60.170 31.365 60.635 31.565 ;
        RECT 59.815 31.195 59.995 31.315 ;
        RECT 58.035 30.935 59.645 31.145 ;
        RECT 59.815 31.025 60.145 31.195 ;
        RECT 59.235 30.835 59.645 30.935 ;
        RECT 58.055 30.005 58.840 30.765 ;
        RECT 59.235 30.175 59.620 30.835 ;
        RECT 59.945 30.235 60.145 31.025 ;
        RECT 60.315 30.005 60.635 31.185 ;
        RECT 60.805 30.875 60.975 31.905 ;
        RECT 61.655 31.875 61.875 32.335 ;
        RECT 61.625 31.850 61.875 31.875 ;
        RECT 61.145 31.255 61.375 31.650 ;
        RECT 61.545 31.425 61.875 31.850 ;
        RECT 62.045 32.175 62.935 32.345 ;
        RECT 63.105 32.175 63.995 32.345 ;
        RECT 62.045 31.450 62.215 32.175 ;
        RECT 62.385 31.620 62.935 32.005 ;
        RECT 63.105 31.620 63.655 32.005 ;
        RECT 63.825 31.450 63.995 32.175 ;
        RECT 62.045 31.380 62.935 31.450 ;
        RECT 62.040 31.355 62.935 31.380 ;
        RECT 62.030 31.340 62.935 31.355 ;
        RECT 62.025 31.325 62.935 31.340 ;
        RECT 62.015 31.320 62.935 31.325 ;
        RECT 62.010 31.310 62.935 31.320 ;
        RECT 62.005 31.300 62.935 31.310 ;
        RECT 61.995 31.295 62.935 31.300 ;
        RECT 61.985 31.285 62.935 31.295 ;
        RECT 61.975 31.280 62.935 31.285 ;
        RECT 61.975 31.275 62.310 31.280 ;
        RECT 61.960 31.270 62.310 31.275 ;
        RECT 61.945 31.260 62.310 31.270 ;
        RECT 61.920 31.255 62.310 31.260 ;
        RECT 61.145 31.250 62.310 31.255 ;
        RECT 61.145 31.215 62.280 31.250 ;
        RECT 61.145 31.190 62.245 31.215 ;
        RECT 61.145 31.160 62.215 31.190 ;
        RECT 61.145 31.130 62.195 31.160 ;
        RECT 61.145 31.100 62.175 31.130 ;
        RECT 61.145 31.090 62.105 31.100 ;
        RECT 61.145 31.080 62.080 31.090 ;
        RECT 61.145 31.065 62.060 31.080 ;
        RECT 61.145 31.050 62.040 31.065 ;
        RECT 61.250 31.040 62.035 31.050 ;
        RECT 61.250 31.005 62.020 31.040 ;
        RECT 60.805 30.175 61.080 30.875 ;
        RECT 61.250 30.755 62.005 31.005 ;
        RECT 62.175 30.685 62.505 30.930 ;
        RECT 62.675 30.830 62.935 31.280 ;
        RECT 63.105 31.380 63.995 31.450 ;
        RECT 64.165 31.875 64.385 32.335 ;
        RECT 64.555 32.015 64.805 32.555 ;
        RECT 64.975 31.905 65.235 32.385 ;
        RECT 64.165 31.850 64.415 31.875 ;
        RECT 64.165 31.425 64.495 31.850 ;
        RECT 63.105 31.355 64.000 31.380 ;
        RECT 63.105 31.340 64.010 31.355 ;
        RECT 63.105 31.325 64.015 31.340 ;
        RECT 63.105 31.320 64.025 31.325 ;
        RECT 63.105 31.310 64.030 31.320 ;
        RECT 63.105 31.300 64.035 31.310 ;
        RECT 63.105 31.295 64.045 31.300 ;
        RECT 63.105 31.285 64.055 31.295 ;
        RECT 63.105 31.280 64.065 31.285 ;
        RECT 63.105 30.830 63.365 31.280 ;
        RECT 63.730 31.275 64.065 31.280 ;
        RECT 63.730 31.270 64.080 31.275 ;
        RECT 63.730 31.260 64.095 31.270 ;
        RECT 63.730 31.255 64.120 31.260 ;
        RECT 64.665 31.255 64.895 31.650 ;
        RECT 63.730 31.250 64.895 31.255 ;
        RECT 63.760 31.215 64.895 31.250 ;
        RECT 63.795 31.190 64.895 31.215 ;
        RECT 63.825 31.160 64.895 31.190 ;
        RECT 63.845 31.130 64.895 31.160 ;
        RECT 63.865 31.100 64.895 31.130 ;
        RECT 63.935 31.090 64.895 31.100 ;
        RECT 63.960 31.080 64.895 31.090 ;
        RECT 63.980 31.065 64.895 31.080 ;
        RECT 64.000 31.050 64.895 31.065 ;
        RECT 64.005 31.040 64.790 31.050 ;
        RECT 64.020 31.005 64.790 31.040 ;
        RECT 62.320 30.660 62.505 30.685 ;
        RECT 63.535 30.685 63.865 30.930 ;
        RECT 64.035 30.755 64.790 31.005 ;
        RECT 65.065 30.875 65.235 31.905 ;
        RECT 65.405 31.785 67.075 32.555 ;
        RECT 67.265 31.865 67.505 32.385 ;
        RECT 67.675 32.060 68.070 32.555 ;
        RECT 68.635 32.225 68.805 32.370 ;
        RECT 68.430 32.030 68.805 32.225 ;
        RECT 65.405 31.265 66.155 31.785 ;
        RECT 66.325 31.095 67.075 31.615 ;
        RECT 63.535 30.660 63.720 30.685 ;
        RECT 62.320 30.560 62.935 30.660 ;
        RECT 61.250 30.005 61.505 30.550 ;
        RECT 61.675 30.175 62.155 30.515 ;
        RECT 62.330 30.005 62.935 30.560 ;
        RECT 63.105 30.560 63.720 30.660 ;
        RECT 63.105 30.005 63.710 30.560 ;
        RECT 63.885 30.175 64.365 30.515 ;
        RECT 64.535 30.005 64.790 30.550 ;
        RECT 64.960 30.175 65.235 30.875 ;
        RECT 65.405 30.005 67.075 31.095 ;
        RECT 67.265 31.060 67.440 31.865 ;
        RECT 68.430 31.695 68.600 32.030 ;
        RECT 69.085 31.985 69.325 32.360 ;
        RECT 69.495 32.050 69.830 32.555 ;
        RECT 70.925 32.055 71.185 32.385 ;
        RECT 71.355 32.055 71.605 32.555 ;
        RECT 69.085 31.835 69.305 31.985 ;
        RECT 67.615 31.335 68.600 31.695 ;
        RECT 68.770 31.505 69.305 31.835 ;
        RECT 67.615 31.315 68.900 31.335 ;
        RECT 68.040 31.165 68.900 31.315 ;
        RECT 67.265 30.275 67.570 31.060 ;
        RECT 67.745 30.685 68.440 30.995 ;
        RECT 67.750 30.005 68.435 30.475 ;
        RECT 68.615 30.220 68.900 31.165 ;
        RECT 69.070 30.855 69.305 31.505 ;
        RECT 69.475 31.025 69.775 31.875 ;
        RECT 69.070 30.625 69.745 30.855 ;
        RECT 69.075 30.005 69.405 30.455 ;
        RECT 69.575 30.195 69.745 30.625 ;
        RECT 70.925 30.725 71.095 32.055 ;
        RECT 71.265 31.335 71.615 31.875 ;
        RECT 71.785 31.235 72.090 32.215 ;
        RECT 72.265 31.535 72.530 32.220 ;
        RECT 73.260 32.005 73.430 32.385 ;
        RECT 73.700 32.175 74.030 32.555 ;
        RECT 73.035 31.835 74.025 32.005 ;
        RECT 72.265 31.365 72.535 31.535 ;
        RECT 72.695 31.065 72.865 31.240 ;
        RECT 71.685 30.895 72.865 31.065 ;
        RECT 71.685 30.725 71.855 30.895 ;
        RECT 73.035 30.725 73.205 31.835 ;
        RECT 73.375 31.315 73.685 31.645 ;
        RECT 73.855 31.315 74.025 31.835 ;
        RECT 70.925 30.555 71.855 30.725 ;
        RECT 72.025 30.555 73.205 30.725 ;
        RECT 73.515 30.755 73.685 31.315 ;
        RECT 74.200 31.095 74.425 32.385 ;
        RECT 74.595 32.175 74.925 32.555 ;
        RECT 75.095 32.005 75.265 32.385 ;
        RECT 74.770 31.835 75.265 32.005 ;
        RECT 74.120 30.925 74.450 31.095 ;
        RECT 74.770 30.755 74.940 31.835 ;
        RECT 75.525 31.805 76.735 32.555 ;
        RECT 75.110 31.535 75.290 31.645 ;
        RECT 75.110 31.365 75.295 31.535 ;
        RECT 75.110 31.005 75.290 31.365 ;
        RECT 75.525 31.095 76.045 31.635 ;
        RECT 76.215 31.265 76.735 31.805 ;
        RECT 73.515 30.585 75.265 30.755 ;
        RECT 70.925 30.175 71.185 30.555 ;
        RECT 71.355 30.005 71.685 30.385 ;
        RECT 72.025 30.175 72.195 30.555 ;
        RECT 72.365 30.005 72.705 30.385 ;
        RECT 72.875 30.175 73.045 30.555 ;
        RECT 73.280 30.005 73.950 30.385 ;
        RECT 74.595 30.005 74.925 30.385 ;
        RECT 75.095 30.175 75.265 30.585 ;
        RECT 75.525 30.005 76.735 31.095 ;
        RECT 5.520 29.835 76.820 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 7.910 28.695 8.230 29.835 ;
        RECT 8.410 28.525 8.605 29.575 ;
        RECT 8.785 28.985 9.115 29.665 ;
        RECT 9.315 29.035 9.570 29.835 ;
        RECT 9.835 29.215 10.005 29.645 ;
        RECT 10.175 29.385 10.505 29.835 ;
        RECT 9.835 28.985 10.515 29.215 ;
        RECT 8.785 28.705 9.135 28.985 ;
        RECT 7.970 28.475 8.230 28.525 ;
        RECT 7.965 28.305 8.230 28.475 ;
        RECT 7.970 28.195 8.230 28.305 ;
        RECT 8.410 28.195 8.795 28.525 ;
        RECT 8.965 28.325 9.135 28.705 ;
        RECT 9.325 28.495 9.570 28.855 ;
        RECT 9.810 28.475 10.110 28.815 ;
        RECT 8.965 28.155 9.485 28.325 ;
        RECT 9.805 28.305 10.110 28.475 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 7.910 27.815 9.125 27.985 ;
        RECT 7.910 27.465 8.200 27.815 ;
        RECT 8.395 27.285 8.725 27.645 ;
        RECT 8.895 27.510 9.125 27.815 ;
        RECT 9.315 27.590 9.485 28.155 ;
        RECT 9.810 27.965 10.110 28.305 ;
        RECT 10.280 28.335 10.515 28.985 ;
        RECT 10.705 28.675 10.990 29.620 ;
        RECT 11.170 29.365 11.855 29.835 ;
        RECT 11.165 28.845 11.860 29.155 ;
        RECT 12.035 28.780 12.340 29.565 ;
        RECT 12.525 28.880 12.795 29.835 ;
        RECT 12.970 29.035 13.225 29.835 ;
        RECT 13.425 28.985 13.755 29.665 ;
        RECT 10.705 28.525 11.565 28.675 ;
        RECT 10.705 28.505 11.995 28.525 ;
        RECT 10.280 28.005 10.835 28.335 ;
        RECT 11.005 28.145 11.995 28.505 ;
        RECT 10.280 27.855 10.495 28.005 ;
        RECT 9.755 27.285 10.085 27.790 ;
        RECT 10.255 27.480 10.495 27.855 ;
        RECT 11.005 27.810 11.175 28.145 ;
        RECT 12.165 27.975 12.340 28.780 ;
        RECT 12.970 28.495 13.215 28.855 ;
        RECT 13.405 28.705 13.755 28.985 ;
        RECT 13.405 28.325 13.575 28.705 ;
        RECT 13.935 28.525 14.130 29.575 ;
        RECT 14.310 28.695 14.630 29.835 ;
        RECT 14.805 28.745 18.315 29.835 ;
        RECT 10.775 27.615 11.175 27.810 ;
        RECT 10.775 27.470 10.945 27.615 ;
        RECT 11.535 27.285 11.935 27.780 ;
        RECT 12.105 27.455 12.340 27.975 ;
        RECT 13.055 28.155 13.575 28.325 ;
        RECT 13.745 28.195 14.130 28.525 ;
        RECT 14.310 28.475 14.570 28.525 ;
        RECT 14.310 28.305 14.575 28.475 ;
        RECT 14.310 28.195 14.570 28.305 ;
        RECT 12.525 27.285 12.795 27.920 ;
        RECT 13.055 27.590 13.225 28.155 ;
        RECT 14.805 28.055 16.455 28.575 ;
        RECT 16.625 28.225 18.315 28.745 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 19.605 29.165 19.885 29.835 ;
        RECT 19.405 28.525 19.720 28.965 ;
        RECT 20.055 28.945 20.355 29.495 ;
        RECT 20.565 29.115 20.895 29.835 ;
        RECT 21.085 29.115 21.535 29.665 ;
        RECT 20.055 28.775 20.995 28.945 ;
        RECT 20.825 28.525 20.995 28.775 ;
        RECT 19.405 28.275 20.095 28.525 ;
        RECT 20.325 28.275 20.655 28.525 ;
        RECT 20.825 28.195 21.115 28.525 ;
        RECT 20.825 28.105 20.995 28.195 ;
        RECT 13.415 27.815 14.630 27.985 ;
        RECT 13.415 27.510 13.645 27.815 ;
        RECT 13.815 27.285 14.145 27.645 ;
        RECT 14.340 27.465 14.630 27.815 ;
        RECT 14.805 27.285 18.315 28.055 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 19.605 27.915 20.995 28.105 ;
        RECT 19.605 27.555 19.935 27.915 ;
        RECT 21.285 27.745 21.535 29.115 ;
        RECT 21.705 28.695 21.995 29.835 ;
        RECT 22.170 28.685 22.430 29.835 ;
        RECT 22.605 28.760 22.860 29.665 ;
        RECT 23.030 29.075 23.360 29.835 ;
        RECT 23.575 28.905 23.745 29.665 ;
        RECT 24.005 29.400 29.350 29.835 ;
        RECT 20.565 27.285 20.815 27.745 ;
        RECT 20.985 27.455 21.535 27.745 ;
        RECT 21.705 27.285 21.995 28.085 ;
        RECT 22.170 27.285 22.430 28.125 ;
        RECT 22.605 28.030 22.775 28.760 ;
        RECT 23.030 28.735 23.745 28.905 ;
        RECT 23.030 28.525 23.200 28.735 ;
        RECT 22.945 28.195 23.200 28.525 ;
        RECT 22.605 27.455 22.860 28.030 ;
        RECT 23.030 28.005 23.200 28.195 ;
        RECT 23.480 28.185 23.835 28.555 ;
        RECT 23.030 27.835 23.745 28.005 ;
        RECT 23.030 27.285 23.360 27.665 ;
        RECT 23.575 27.455 23.745 27.835 ;
        RECT 25.590 27.830 25.930 28.660 ;
        RECT 27.410 28.150 27.760 29.400 ;
        RECT 29.525 28.745 33.035 29.835 ;
        RECT 29.525 28.055 31.175 28.575 ;
        RECT 31.345 28.225 33.035 28.745 ;
        RECT 33.205 28.230 33.485 29.665 ;
        RECT 33.655 29.060 34.365 29.835 ;
        RECT 34.535 28.890 34.865 29.665 ;
        RECT 33.715 28.675 34.865 28.890 ;
        RECT 24.005 27.285 29.350 27.830 ;
        RECT 29.525 27.285 33.035 28.055 ;
        RECT 33.205 27.455 33.545 28.230 ;
        RECT 33.715 28.105 34.000 28.675 ;
        RECT 34.185 28.275 34.655 28.505 ;
        RECT 35.060 28.475 35.275 29.590 ;
        RECT 35.455 29.115 35.785 29.835 ;
        RECT 35.965 28.985 36.225 29.665 ;
        RECT 36.395 29.055 36.645 29.835 ;
        RECT 36.895 29.285 37.145 29.665 ;
        RECT 37.315 29.455 37.670 29.835 ;
        RECT 38.675 29.445 39.010 29.665 ;
        RECT 38.275 29.285 38.505 29.325 ;
        RECT 36.895 29.085 38.505 29.285 ;
        RECT 36.895 29.075 37.730 29.085 ;
        RECT 38.320 28.995 38.505 29.085 ;
        RECT 35.565 28.475 35.795 28.815 ;
        RECT 34.825 28.295 35.275 28.475 ;
        RECT 34.825 28.275 35.155 28.295 ;
        RECT 35.465 28.275 35.795 28.475 ;
        RECT 33.715 27.915 34.425 28.105 ;
        RECT 34.125 27.775 34.425 27.915 ;
        RECT 34.615 27.915 35.795 28.105 ;
        RECT 34.615 27.835 34.945 27.915 ;
        RECT 34.125 27.765 34.440 27.775 ;
        RECT 34.125 27.755 34.450 27.765 ;
        RECT 34.125 27.750 34.460 27.755 ;
        RECT 33.715 27.285 33.885 27.745 ;
        RECT 34.125 27.740 34.465 27.750 ;
        RECT 34.125 27.735 34.470 27.740 ;
        RECT 34.125 27.725 34.475 27.735 ;
        RECT 34.125 27.720 34.480 27.725 ;
        RECT 34.125 27.455 34.485 27.720 ;
        RECT 35.115 27.285 35.285 27.745 ;
        RECT 35.455 27.455 35.795 27.915 ;
        RECT 35.965 27.785 36.135 28.985 ;
        RECT 37.835 28.885 38.165 28.915 ;
        RECT 36.365 28.825 38.165 28.885 ;
        RECT 38.755 28.825 39.010 29.445 ;
        RECT 39.275 29.215 39.445 29.645 ;
        RECT 39.615 29.385 39.945 29.835 ;
        RECT 39.275 28.985 39.955 29.215 ;
        RECT 36.305 28.715 39.010 28.825 ;
        RECT 36.305 28.680 36.505 28.715 ;
        RECT 36.305 28.105 36.475 28.680 ;
        RECT 37.835 28.655 39.010 28.715 ;
        RECT 36.705 28.240 37.115 28.545 ;
        RECT 37.285 28.275 37.615 28.485 ;
        RECT 36.305 27.985 36.575 28.105 ;
        RECT 36.305 27.940 37.150 27.985 ;
        RECT 36.395 27.815 37.150 27.940 ;
        RECT 37.405 27.875 37.615 28.275 ;
        RECT 37.860 28.275 38.335 28.485 ;
        RECT 38.525 28.275 39.015 28.475 ;
        RECT 37.860 27.875 38.080 28.275 ;
        RECT 39.250 28.135 39.550 28.815 ;
        RECT 35.965 27.455 36.225 27.785 ;
        RECT 36.980 27.665 37.150 27.815 ;
        RECT 36.395 27.285 36.725 27.645 ;
        RECT 36.980 27.455 38.280 27.665 ;
        RECT 38.555 27.285 39.010 28.050 ;
        RECT 39.245 27.965 39.550 28.135 ;
        RECT 39.720 28.335 39.955 28.985 ;
        RECT 40.145 28.675 40.430 29.620 ;
        RECT 40.610 29.365 41.295 29.835 ;
        RECT 40.605 28.845 41.300 29.155 ;
        RECT 41.475 28.780 41.780 29.565 ;
        RECT 41.965 28.880 42.235 29.835 ;
        RECT 40.145 28.525 41.005 28.675 ;
        RECT 40.145 28.505 41.435 28.525 ;
        RECT 39.720 28.005 40.275 28.335 ;
        RECT 40.445 28.145 41.435 28.505 ;
        RECT 39.720 27.855 39.935 28.005 ;
        RECT 39.195 27.285 39.525 27.790 ;
        RECT 39.695 27.480 39.935 27.855 ;
        RECT 40.445 27.810 40.615 28.145 ;
        RECT 41.605 27.975 41.780 28.780 ;
        RECT 42.405 28.745 44.075 29.835 ;
        RECT 40.215 27.615 40.615 27.810 ;
        RECT 40.215 27.470 40.385 27.615 ;
        RECT 40.975 27.285 41.375 27.780 ;
        RECT 41.545 27.455 41.780 27.975 ;
        RECT 42.405 28.055 43.155 28.575 ;
        RECT 43.325 28.225 44.075 28.745 ;
        RECT 44.245 28.670 44.535 29.835 ;
        RECT 44.705 29.400 50.050 29.835 ;
        RECT 41.965 27.285 42.235 27.920 ;
        RECT 42.405 27.285 44.075 28.055 ;
        RECT 44.245 27.285 44.535 28.010 ;
        RECT 46.290 27.830 46.630 28.660 ;
        RECT 48.110 28.150 48.460 29.400 ;
        RECT 51.155 28.885 51.430 29.655 ;
        RECT 51.600 29.225 51.930 29.655 ;
        RECT 52.100 29.395 52.295 29.835 ;
        RECT 52.475 29.225 52.805 29.655 ;
        RECT 52.985 29.400 58.330 29.835 ;
        RECT 51.600 29.055 52.805 29.225 ;
        RECT 51.155 28.695 51.740 28.885 ;
        RECT 51.910 28.725 52.805 29.055 ;
        RECT 51.155 27.875 51.395 28.525 ;
        RECT 51.565 28.025 51.740 28.695 ;
        RECT 51.910 28.195 52.325 28.525 ;
        RECT 52.505 28.195 52.800 28.525 ;
        RECT 51.565 27.845 51.895 28.025 ;
        RECT 44.705 27.285 50.050 27.830 ;
        RECT 51.170 27.285 51.500 27.675 ;
        RECT 51.670 27.465 51.895 27.845 ;
        RECT 52.095 27.575 52.325 28.195 ;
        RECT 52.505 27.285 52.805 28.015 ;
        RECT 54.570 27.830 54.910 28.660 ;
        RECT 56.390 28.150 56.740 29.400 ;
        RECT 58.505 28.745 60.175 29.835 ;
        RECT 60.345 29.280 60.950 29.835 ;
        RECT 61.125 29.325 61.605 29.665 ;
        RECT 61.775 29.290 62.030 29.835 ;
        RECT 60.345 29.180 60.960 29.280 ;
        RECT 60.775 29.155 60.960 29.180 ;
        RECT 58.505 28.055 59.255 28.575 ;
        RECT 59.425 28.225 60.175 28.745 ;
        RECT 60.345 28.560 60.605 29.010 ;
        RECT 60.775 28.910 61.105 29.155 ;
        RECT 61.275 28.835 62.030 29.085 ;
        RECT 62.200 28.965 62.475 29.665 ;
        RECT 61.260 28.800 62.030 28.835 ;
        RECT 61.245 28.790 62.030 28.800 ;
        RECT 61.240 28.775 62.135 28.790 ;
        RECT 61.220 28.760 62.135 28.775 ;
        RECT 61.200 28.750 62.135 28.760 ;
        RECT 61.175 28.740 62.135 28.750 ;
        RECT 61.105 28.710 62.135 28.740 ;
        RECT 61.085 28.680 62.135 28.710 ;
        RECT 61.065 28.650 62.135 28.680 ;
        RECT 61.035 28.625 62.135 28.650 ;
        RECT 61.000 28.590 62.135 28.625 ;
        RECT 60.970 28.585 62.135 28.590 ;
        RECT 60.970 28.580 61.360 28.585 ;
        RECT 60.970 28.570 61.335 28.580 ;
        RECT 60.970 28.565 61.320 28.570 ;
        RECT 60.970 28.560 61.305 28.565 ;
        RECT 60.345 28.555 61.305 28.560 ;
        RECT 60.345 28.545 61.295 28.555 ;
        RECT 60.345 28.540 61.285 28.545 ;
        RECT 60.345 28.530 61.275 28.540 ;
        RECT 60.345 28.520 61.270 28.530 ;
        RECT 60.345 28.515 61.265 28.520 ;
        RECT 60.345 28.500 61.255 28.515 ;
        RECT 60.345 28.485 61.250 28.500 ;
        RECT 60.345 28.460 61.240 28.485 ;
        RECT 60.345 28.390 61.235 28.460 ;
        RECT 52.985 27.285 58.330 27.830 ;
        RECT 58.505 27.285 60.175 28.055 ;
        RECT 60.345 27.835 60.895 28.220 ;
        RECT 61.065 27.665 61.235 28.390 ;
        RECT 60.345 27.495 61.235 27.665 ;
        RECT 61.405 27.990 61.735 28.415 ;
        RECT 61.905 28.190 62.135 28.585 ;
        RECT 61.405 27.505 61.625 27.990 ;
        RECT 62.305 27.935 62.475 28.965 ;
        RECT 62.645 28.745 63.855 29.835 ;
        RECT 61.795 27.285 62.045 27.825 ;
        RECT 62.215 27.455 62.475 27.935 ;
        RECT 62.645 28.035 63.165 28.575 ;
        RECT 63.335 28.205 63.855 28.745 ;
        RECT 64.035 28.695 64.365 29.835 ;
        RECT 64.895 28.865 65.225 29.650 ;
        RECT 65.405 29.325 66.595 29.615 ;
        RECT 64.545 28.695 65.225 28.865 ;
        RECT 65.425 28.985 66.595 29.155 ;
        RECT 66.765 29.035 67.045 29.835 ;
        RECT 65.425 28.695 65.750 28.985 ;
        RECT 66.425 28.865 66.595 28.985 ;
        RECT 64.025 28.275 64.375 28.525 ;
        RECT 64.545 28.095 64.715 28.695 ;
        RECT 65.920 28.525 66.115 28.815 ;
        RECT 66.425 28.695 67.085 28.865 ;
        RECT 67.255 28.695 67.530 29.665 ;
        RECT 67.745 29.495 68.885 29.665 ;
        RECT 67.745 29.035 68.045 29.495 ;
        RECT 68.215 28.865 68.545 29.325 ;
        RECT 67.785 28.815 68.545 28.865 ;
        RECT 66.915 28.525 67.085 28.695 ;
        RECT 64.885 28.275 65.235 28.525 ;
        RECT 65.405 28.195 65.750 28.525 ;
        RECT 65.920 28.195 66.745 28.525 ;
        RECT 66.915 28.195 67.190 28.525 ;
        RECT 62.645 27.285 63.855 28.035 ;
        RECT 64.035 27.285 64.305 28.095 ;
        RECT 64.475 27.455 64.805 28.095 ;
        RECT 64.975 27.285 65.215 28.095 ;
        RECT 66.915 28.025 67.085 28.195 ;
        RECT 65.420 27.855 67.085 28.025 ;
        RECT 67.360 27.960 67.530 28.695 ;
        RECT 67.765 28.645 68.545 28.815 ;
        RECT 68.715 28.865 68.885 29.495 ;
        RECT 69.055 29.035 69.385 29.835 ;
        RECT 69.555 28.865 69.830 29.665 ;
        RECT 68.715 28.655 69.830 28.865 ;
        RECT 70.005 28.670 70.295 29.835 ;
        RECT 70.545 28.905 70.725 29.665 ;
        RECT 70.905 29.075 71.235 29.835 ;
        RECT 70.545 28.735 71.220 28.905 ;
        RECT 71.405 28.760 71.675 29.665 ;
        RECT 71.845 28.825 72.105 29.835 ;
        RECT 72.275 28.995 72.550 29.665 ;
        RECT 65.420 27.505 65.675 27.855 ;
        RECT 65.845 27.285 66.175 27.685 ;
        RECT 66.345 27.505 66.515 27.855 ;
        RECT 66.685 27.285 67.065 27.685 ;
        RECT 67.255 27.615 67.530 27.960 ;
        RECT 67.785 28.105 68.000 28.645 ;
        RECT 71.050 28.590 71.220 28.735 ;
        RECT 68.170 28.275 68.940 28.475 ;
        RECT 69.110 28.275 69.830 28.475 ;
        RECT 70.485 28.185 70.825 28.555 ;
        RECT 71.050 28.260 71.325 28.590 ;
        RECT 67.785 27.935 69.385 28.105 ;
        RECT 68.215 27.925 69.385 27.935 ;
        RECT 67.755 27.285 68.045 27.755 ;
        RECT 68.215 27.455 68.545 27.925 ;
        RECT 68.715 27.285 68.885 27.755 ;
        RECT 69.055 27.455 69.385 27.925 ;
        RECT 69.555 27.285 69.830 28.105 ;
        RECT 70.005 27.285 70.295 28.010 ;
        RECT 71.050 28.005 71.220 28.260 ;
        RECT 70.555 27.835 71.220 28.005 ;
        RECT 71.495 27.960 71.675 28.760 ;
        RECT 72.275 28.645 72.445 28.995 ;
        RECT 72.750 28.990 72.965 29.835 ;
        RECT 73.150 29.325 73.625 29.665 ;
        RECT 73.805 29.330 74.435 29.835 ;
        RECT 73.805 29.155 73.995 29.330 ;
        RECT 73.190 28.795 73.440 29.090 ;
        RECT 73.665 28.965 73.995 29.155 ;
        RECT 74.165 28.795 74.420 29.160 ;
        RECT 71.845 28.125 72.460 28.645 ;
        RECT 72.630 28.625 74.420 28.795 ;
        RECT 75.525 28.745 76.735 29.835 ;
        RECT 72.630 28.195 72.860 28.625 ;
        RECT 70.555 27.455 70.725 27.835 ;
        RECT 70.905 27.285 71.235 27.665 ;
        RECT 71.415 27.455 71.675 27.960 ;
        RECT 71.845 27.285 72.120 27.945 ;
        RECT 72.290 27.915 72.460 28.125 ;
        RECT 73.045 27.950 73.455 28.445 ;
        RECT 72.290 27.455 72.540 27.915 ;
        RECT 72.715 27.285 73.045 27.780 ;
        RECT 73.225 27.505 73.455 27.950 ;
        RECT 73.625 27.770 73.880 28.625 ;
        RECT 74.050 27.965 74.435 28.445 ;
        RECT 75.525 28.205 76.045 28.745 ;
        RECT 76.215 28.035 76.735 28.575 ;
        RECT 73.625 27.505 74.415 27.770 ;
        RECT 75.525 27.285 76.735 28.035 ;
        RECT 5.520 27.115 76.820 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 6.985 26.545 7.420 26.945 ;
        RECT 7.590 26.715 7.975 27.115 ;
        RECT 6.985 26.375 7.975 26.545 ;
        RECT 8.145 26.375 8.570 26.945 ;
        RECT 8.760 26.545 9.015 26.945 ;
        RECT 9.185 26.715 9.570 27.115 ;
        RECT 8.760 26.375 9.570 26.545 ;
        RECT 9.740 26.375 9.985 26.945 ;
        RECT 10.175 26.545 10.430 26.945 ;
        RECT 10.600 26.715 10.985 27.115 ;
        RECT 10.175 26.375 10.985 26.545 ;
        RECT 11.155 26.375 11.415 26.945 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 7.640 26.205 7.975 26.375 ;
        RECT 8.220 26.205 8.570 26.375 ;
        RECT 9.220 26.205 9.570 26.375 ;
        RECT 9.815 26.205 9.985 26.375 ;
        RECT 10.635 26.205 10.985 26.375 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 6.985 25.500 7.470 26.205 ;
        RECT 7.640 25.875 8.050 26.205 ;
        RECT 7.640 25.330 7.975 25.875 ;
        RECT 8.220 25.705 9.050 26.205 ;
        RECT 6.985 25.160 7.975 25.330 ;
        RECT 8.145 25.525 9.050 25.705 ;
        RECT 9.220 25.875 9.645 26.205 ;
        RECT 6.985 24.735 7.420 25.160 ;
        RECT 7.590 24.565 7.975 24.990 ;
        RECT 8.145 24.735 8.570 25.525 ;
        RECT 9.220 25.355 9.570 25.875 ;
        RECT 9.815 25.705 10.465 26.205 ;
        RECT 8.740 25.160 9.570 25.355 ;
        RECT 9.740 25.525 10.465 25.705 ;
        RECT 10.635 25.875 11.060 26.205 ;
        RECT 8.740 24.735 9.015 25.160 ;
        RECT 9.185 24.565 9.570 24.990 ;
        RECT 9.740 24.735 9.985 25.525 ;
        RECT 10.635 25.355 10.985 25.875 ;
        RECT 11.230 25.705 11.415 26.375 ;
        RECT 11.585 26.315 11.875 27.115 ;
        RECT 12.045 26.655 12.595 26.945 ;
        RECT 12.765 26.655 13.015 27.115 ;
        RECT 10.175 25.160 10.985 25.355 ;
        RECT 10.175 24.735 10.430 25.160 ;
        RECT 10.600 24.565 10.985 24.990 ;
        RECT 11.155 24.735 11.415 25.705 ;
        RECT 11.585 24.565 11.875 25.705 ;
        RECT 12.045 25.285 12.295 26.655 ;
        RECT 13.645 26.485 13.975 26.845 ;
        RECT 12.585 26.295 13.975 26.485 ;
        RECT 14.345 26.345 16.015 27.115 ;
        RECT 16.275 26.565 16.445 26.945 ;
        RECT 16.615 26.735 16.945 27.115 ;
        RECT 16.275 26.395 16.770 26.565 ;
        RECT 12.585 26.205 12.755 26.295 ;
        RECT 12.465 25.875 12.755 26.205 ;
        RECT 12.925 25.875 13.255 26.125 ;
        RECT 13.485 25.875 14.175 26.125 ;
        RECT 12.585 25.625 12.755 25.875 ;
        RECT 12.585 25.455 13.525 25.625 ;
        RECT 12.045 24.735 12.495 25.285 ;
        RECT 12.685 24.565 13.015 25.285 ;
        RECT 13.225 24.905 13.525 25.455 ;
        RECT 13.860 25.435 14.175 25.875 ;
        RECT 14.345 25.825 15.095 26.345 ;
        RECT 15.265 25.655 16.015 26.175 ;
        RECT 16.250 25.755 16.430 26.205 ;
        RECT 13.695 24.565 13.975 25.235 ;
        RECT 14.345 24.565 16.015 25.655 ;
        RECT 16.245 25.585 16.430 25.755 ;
        RECT 16.250 25.565 16.430 25.585 ;
        RECT 16.600 25.315 16.770 26.395 ;
        RECT 17.115 25.655 17.340 26.945 ;
        RECT 17.510 26.735 17.840 27.115 ;
        RECT 18.110 26.565 18.280 26.945 ;
        RECT 17.515 26.395 18.505 26.565 ;
        RECT 17.515 25.875 17.685 26.395 ;
        RECT 17.855 25.875 18.165 26.205 ;
        RECT 17.090 25.485 17.420 25.655 ;
        RECT 17.855 25.315 18.025 25.875 ;
        RECT 16.275 25.145 18.025 25.315 ;
        RECT 18.335 25.285 18.505 26.395 ;
        RECT 19.010 26.095 19.275 26.780 ;
        RECT 19.005 25.925 19.275 26.095 ;
        RECT 18.675 25.625 18.845 25.800 ;
        RECT 19.450 25.795 19.755 26.775 ;
        RECT 19.935 26.615 20.185 27.115 ;
        RECT 20.355 26.615 20.615 26.945 ;
        RECT 19.925 25.895 20.275 26.435 ;
        RECT 18.675 25.455 19.855 25.625 ;
        RECT 19.685 25.285 19.855 25.455 ;
        RECT 20.445 25.285 20.615 26.615 ;
        RECT 20.790 26.275 21.050 27.115 ;
        RECT 21.225 26.370 21.480 26.945 ;
        RECT 21.650 26.735 21.980 27.115 ;
        RECT 22.195 26.565 22.365 26.945 ;
        RECT 21.650 26.395 22.365 26.565 ;
        RECT 23.700 26.465 24.030 26.930 ;
        RECT 24.200 26.645 24.370 27.115 ;
        RECT 24.540 26.465 24.870 26.945 ;
        RECT 16.275 24.735 16.445 25.145 ;
        RECT 18.335 25.115 19.515 25.285 ;
        RECT 19.685 25.115 20.615 25.285 ;
        RECT 16.615 24.565 16.945 24.945 ;
        RECT 17.590 24.565 18.260 24.945 ;
        RECT 18.495 24.735 18.665 25.115 ;
        RECT 18.835 24.565 19.175 24.945 ;
        RECT 19.345 24.735 19.515 25.115 ;
        RECT 19.855 24.565 20.185 24.945 ;
        RECT 20.355 24.735 20.615 25.115 ;
        RECT 20.790 24.565 21.050 25.715 ;
        RECT 21.225 25.640 21.395 26.370 ;
        RECT 21.650 26.205 21.820 26.395 ;
        RECT 23.700 26.295 24.870 26.465 ;
        RECT 21.565 25.875 21.820 26.205 ;
        RECT 21.650 25.665 21.820 25.875 ;
        RECT 22.100 25.845 22.455 26.215 ;
        RECT 23.545 25.915 24.190 26.125 ;
        RECT 24.360 25.915 24.930 26.125 ;
        RECT 25.100 25.745 25.270 26.945 ;
        RECT 25.810 26.545 25.980 26.750 ;
        RECT 21.225 24.735 21.480 25.640 ;
        RECT 21.650 25.495 22.365 25.665 ;
        RECT 21.650 24.565 21.980 25.325 ;
        RECT 22.195 24.735 22.365 25.495 ;
        RECT 23.760 24.565 24.090 25.665 ;
        RECT 24.565 25.335 25.270 25.745 ;
        RECT 25.440 26.375 25.980 26.545 ;
        RECT 26.260 26.375 26.430 27.115 ;
        RECT 26.695 26.375 27.055 26.750 ;
        RECT 25.440 25.675 25.610 26.375 ;
        RECT 25.780 25.875 26.110 26.205 ;
        RECT 26.280 25.875 26.630 26.205 ;
        RECT 25.440 25.505 26.065 25.675 ;
        RECT 26.280 25.335 26.545 25.875 ;
        RECT 26.800 25.720 27.055 26.375 ;
        RECT 27.225 26.345 30.735 27.115 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 31.875 26.575 32.100 26.935 ;
        RECT 32.280 26.745 32.610 27.115 ;
        RECT 32.790 26.575 33.045 26.935 ;
        RECT 33.610 26.745 34.355 27.115 ;
        RECT 31.875 26.385 34.360 26.575 ;
        RECT 27.225 25.825 28.875 26.345 ;
        RECT 24.565 25.165 26.545 25.335 ;
        RECT 24.565 24.735 24.890 25.165 ;
        RECT 25.060 24.565 25.390 24.985 ;
        RECT 26.135 24.565 26.545 24.995 ;
        RECT 26.715 24.735 27.055 25.720 ;
        RECT 29.045 25.655 30.735 26.175 ;
        RECT 31.835 25.875 32.105 26.205 ;
        RECT 32.285 25.875 32.720 26.205 ;
        RECT 32.900 25.875 33.475 26.205 ;
        RECT 33.655 25.875 33.935 26.205 ;
        RECT 27.225 24.565 30.735 25.655 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 34.135 25.695 34.360 26.385 ;
        RECT 31.865 25.515 34.360 25.695 ;
        RECT 34.535 25.515 34.870 26.935 ;
        RECT 31.865 24.745 32.155 25.515 ;
        RECT 32.725 25.105 33.915 25.335 ;
        RECT 32.725 24.745 32.985 25.105 ;
        RECT 33.155 24.565 33.485 24.935 ;
        RECT 33.655 24.745 33.915 25.105 ;
        RECT 34.105 24.565 34.435 25.285 ;
        RECT 34.605 24.745 34.870 25.515 ;
        RECT 35.055 24.745 35.315 26.935 ;
        RECT 35.575 26.745 36.245 27.115 ;
        RECT 36.425 26.565 36.735 26.935 ;
        RECT 35.505 26.365 36.735 26.565 ;
        RECT 35.505 25.695 35.795 26.365 ;
        RECT 36.915 26.185 37.145 26.825 ;
        RECT 37.325 26.385 37.615 27.115 ;
        RECT 37.805 26.345 39.475 27.115 ;
        RECT 35.975 25.875 36.440 26.185 ;
        RECT 36.620 25.875 37.145 26.185 ;
        RECT 37.325 25.875 37.625 26.205 ;
        RECT 37.805 25.825 38.555 26.345 ;
        RECT 39.655 26.305 39.925 27.115 ;
        RECT 40.095 26.305 40.425 26.945 ;
        RECT 40.595 26.305 40.835 27.115 ;
        RECT 41.025 26.345 44.535 27.115 ;
        RECT 35.505 25.475 36.275 25.695 ;
        RECT 35.485 24.565 35.825 25.295 ;
        RECT 36.005 24.745 36.275 25.475 ;
        RECT 36.455 25.455 37.615 25.695 ;
        RECT 38.725 25.655 39.475 26.175 ;
        RECT 39.645 25.875 39.995 26.125 ;
        RECT 40.165 25.705 40.335 26.305 ;
        RECT 40.505 25.875 40.855 26.125 ;
        RECT 41.025 25.825 42.675 26.345 ;
        RECT 36.455 24.745 36.685 25.455 ;
        RECT 36.855 24.565 37.185 25.275 ;
        RECT 37.355 24.745 37.615 25.455 ;
        RECT 37.805 24.565 39.475 25.655 ;
        RECT 39.655 24.565 39.985 25.705 ;
        RECT 40.165 25.535 40.845 25.705 ;
        RECT 42.845 25.655 44.535 26.175 ;
        RECT 40.515 24.750 40.845 25.535 ;
        RECT 41.025 24.565 44.535 25.655 ;
        RECT 44.705 24.735 44.985 26.835 ;
        RECT 45.215 26.655 45.385 27.115 ;
        RECT 45.655 26.725 46.905 26.905 ;
        RECT 46.040 26.485 46.405 26.555 ;
        RECT 45.155 26.305 46.405 26.485 ;
        RECT 46.575 26.505 46.905 26.725 ;
        RECT 47.075 26.675 47.245 27.115 ;
        RECT 47.415 26.505 47.755 26.920 ;
        RECT 46.575 26.335 47.755 26.505 ;
        RECT 47.925 26.345 49.595 27.115 ;
        RECT 45.155 25.705 45.430 26.305 ;
        RECT 45.600 25.875 45.955 26.125 ;
        RECT 46.150 26.095 46.615 26.125 ;
        RECT 46.145 25.925 46.615 26.095 ;
        RECT 46.150 25.875 46.615 25.925 ;
        RECT 46.785 25.875 47.115 26.125 ;
        RECT 47.290 25.925 47.755 26.125 ;
        RECT 46.935 25.755 47.115 25.875 ;
        RECT 47.925 25.825 48.675 26.345 ;
        RECT 50.285 26.295 50.495 27.115 ;
        RECT 50.665 26.315 50.995 26.945 ;
        RECT 45.155 25.495 46.765 25.705 ;
        RECT 46.935 25.585 47.265 25.755 ;
        RECT 46.355 25.395 46.765 25.495 ;
        RECT 45.175 24.565 45.960 25.325 ;
        RECT 46.355 24.735 46.740 25.395 ;
        RECT 47.065 24.795 47.265 25.585 ;
        RECT 47.435 24.565 47.755 25.745 ;
        RECT 48.845 25.655 49.595 26.175 ;
        RECT 50.665 25.715 50.915 26.315 ;
        RECT 51.165 26.295 51.395 27.115 ;
        RECT 51.605 26.570 56.950 27.115 ;
        RECT 51.085 25.875 51.415 26.125 ;
        RECT 53.190 25.740 53.530 26.570 ;
        RECT 57.125 26.390 57.415 27.115 ;
        RECT 57.605 26.385 57.895 27.115 ;
        RECT 47.925 24.565 49.595 25.655 ;
        RECT 50.285 24.565 50.495 25.705 ;
        RECT 50.665 24.735 50.995 25.715 ;
        RECT 51.165 24.565 51.395 25.705 ;
        RECT 55.010 25.000 55.360 26.250 ;
        RECT 57.595 25.875 57.895 26.205 ;
        RECT 58.075 26.185 58.305 26.825 ;
        RECT 58.485 26.565 58.795 26.935 ;
        RECT 58.975 26.745 59.645 27.115 ;
        RECT 58.485 26.365 59.715 26.565 ;
        RECT 58.075 25.875 58.600 26.185 ;
        RECT 58.780 25.875 59.245 26.185 ;
        RECT 51.605 24.565 56.950 25.000 ;
        RECT 57.125 24.565 57.415 25.730 ;
        RECT 59.425 25.695 59.715 26.365 ;
        RECT 57.605 25.455 58.765 25.695 ;
        RECT 57.605 24.745 57.865 25.455 ;
        RECT 58.035 24.565 58.365 25.275 ;
        RECT 58.535 24.745 58.765 25.455 ;
        RECT 58.945 25.475 59.715 25.695 ;
        RECT 58.945 24.745 59.215 25.475 ;
        RECT 59.395 24.565 59.735 25.295 ;
        RECT 59.905 24.745 60.165 26.935 ;
        RECT 61.265 26.655 61.825 26.945 ;
        RECT 61.995 26.655 62.245 27.115 ;
        RECT 61.265 25.285 61.515 26.655 ;
        RECT 62.865 26.485 63.195 26.845 ;
        RECT 61.805 26.295 63.195 26.485 ;
        RECT 63.565 26.345 66.155 27.115 ;
        RECT 66.785 26.440 67.045 26.945 ;
        RECT 67.225 26.735 67.555 27.115 ;
        RECT 67.735 26.565 67.905 26.945 ;
        RECT 61.805 26.205 61.975 26.295 ;
        RECT 61.685 25.875 61.975 26.205 ;
        RECT 62.145 25.875 62.485 26.125 ;
        RECT 62.705 25.875 63.380 26.125 ;
        RECT 61.805 25.625 61.975 25.875 ;
        RECT 61.805 25.455 62.745 25.625 ;
        RECT 63.115 25.515 63.380 25.875 ;
        RECT 63.565 25.825 64.775 26.345 ;
        RECT 64.945 25.655 66.155 26.175 ;
        RECT 61.265 24.735 61.725 25.285 ;
        RECT 61.915 24.565 62.245 25.285 ;
        RECT 62.445 24.905 62.745 25.455 ;
        RECT 62.915 24.565 63.195 25.235 ;
        RECT 63.565 24.565 66.155 25.655 ;
        RECT 66.785 25.640 66.965 26.440 ;
        RECT 67.240 26.395 67.905 26.565 ;
        RECT 67.240 26.140 67.410 26.395 ;
        RECT 68.170 26.275 68.430 27.115 ;
        RECT 68.605 26.370 68.860 26.945 ;
        RECT 69.030 26.735 69.360 27.115 ;
        RECT 69.575 26.565 69.745 26.945 ;
        RECT 69.030 26.395 69.745 26.565 ;
        RECT 70.095 26.565 70.265 26.945 ;
        RECT 70.445 26.735 70.775 27.115 ;
        RECT 70.095 26.395 70.760 26.565 ;
        RECT 70.955 26.440 71.215 26.945 ;
        RECT 67.135 25.810 67.410 26.140 ;
        RECT 67.635 25.845 67.975 26.215 ;
        RECT 67.240 25.665 67.410 25.810 ;
        RECT 66.785 24.735 67.055 25.640 ;
        RECT 67.240 25.495 67.915 25.665 ;
        RECT 67.225 24.565 67.555 25.325 ;
        RECT 67.735 24.735 67.915 25.495 ;
        RECT 68.170 24.565 68.430 25.715 ;
        RECT 68.605 25.640 68.775 26.370 ;
        RECT 69.030 26.205 69.200 26.395 ;
        RECT 68.945 25.875 69.200 26.205 ;
        RECT 69.030 25.665 69.200 25.875 ;
        RECT 69.480 25.845 69.835 26.215 ;
        RECT 70.025 25.845 70.365 26.215 ;
        RECT 70.590 26.140 70.760 26.395 ;
        RECT 70.590 25.810 70.865 26.140 ;
        RECT 70.590 25.665 70.760 25.810 ;
        RECT 68.605 24.735 68.860 25.640 ;
        RECT 69.030 25.495 69.745 25.665 ;
        RECT 69.030 24.565 69.360 25.325 ;
        RECT 69.575 24.735 69.745 25.495 ;
        RECT 70.085 25.495 70.760 25.665 ;
        RECT 71.035 25.640 71.215 26.440 ;
        RECT 71.850 26.275 72.110 27.115 ;
        RECT 72.285 26.370 72.540 26.945 ;
        RECT 72.710 26.735 73.040 27.115 ;
        RECT 73.255 26.565 73.425 26.945 ;
        RECT 73.690 26.715 74.025 27.115 ;
        RECT 72.710 26.395 73.425 26.565 ;
        RECT 74.195 26.545 74.400 26.945 ;
        RECT 74.610 26.635 74.885 27.115 ;
        RECT 75.095 26.615 75.355 26.945 ;
        RECT 70.085 24.735 70.265 25.495 ;
        RECT 70.445 24.565 70.775 25.325 ;
        RECT 70.945 24.735 71.215 25.640 ;
        RECT 71.850 24.565 72.110 25.715 ;
        RECT 72.285 25.640 72.455 26.370 ;
        RECT 72.710 26.205 72.880 26.395 ;
        RECT 73.715 26.375 74.400 26.545 ;
        RECT 72.625 25.875 72.880 26.205 ;
        RECT 72.710 25.665 72.880 25.875 ;
        RECT 73.160 25.845 73.515 26.215 ;
        RECT 72.285 24.735 72.540 25.640 ;
        RECT 72.710 25.495 73.425 25.665 ;
        RECT 72.710 24.565 73.040 25.325 ;
        RECT 73.255 24.735 73.425 25.495 ;
        RECT 73.715 25.345 74.055 26.375 ;
        RECT 74.225 25.705 74.475 26.205 ;
        RECT 74.655 25.875 75.015 26.455 ;
        RECT 75.185 25.705 75.355 26.615 ;
        RECT 75.525 26.365 76.735 27.115 ;
        RECT 74.225 25.535 75.355 25.705 ;
        RECT 73.715 25.170 74.380 25.345 ;
        RECT 73.690 24.565 74.025 24.990 ;
        RECT 74.195 24.765 74.380 25.170 ;
        RECT 74.585 24.565 74.915 25.345 ;
        RECT 75.085 24.765 75.355 25.535 ;
        RECT 75.525 25.655 76.045 26.195 ;
        RECT 76.215 25.825 76.735 26.365 ;
        RECT 75.525 24.565 76.735 25.655 ;
        RECT 5.520 24.395 76.820 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 6.990 23.245 7.250 24.395 ;
        RECT 7.425 23.320 7.680 24.225 ;
        RECT 7.850 23.635 8.180 24.395 ;
        RECT 8.395 23.465 8.565 24.225 ;
        RECT 9.835 23.775 10.005 24.205 ;
        RECT 10.175 23.945 10.505 24.395 ;
        RECT 9.835 23.545 10.510 23.775 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 6.990 21.845 7.250 22.685 ;
        RECT 7.425 22.590 7.595 23.320 ;
        RECT 7.850 23.295 8.565 23.465 ;
        RECT 7.850 23.085 8.020 23.295 ;
        RECT 7.765 22.755 8.020 23.085 ;
        RECT 7.425 22.015 7.680 22.590 ;
        RECT 7.850 22.565 8.020 22.755 ;
        RECT 8.300 22.745 8.655 23.115 ;
        RECT 7.850 22.395 8.565 22.565 ;
        RECT 9.805 22.525 10.105 23.375 ;
        RECT 10.275 22.895 10.510 23.545 ;
        RECT 10.680 23.235 10.965 24.180 ;
        RECT 11.145 23.925 11.830 24.395 ;
        RECT 11.140 23.405 11.835 23.715 ;
        RECT 12.010 23.340 12.315 24.125 ;
        RECT 10.680 23.085 11.540 23.235 ;
        RECT 10.680 23.065 11.965 23.085 ;
        RECT 10.275 22.565 10.810 22.895 ;
        RECT 10.980 22.705 11.965 23.065 ;
        RECT 10.275 22.415 10.495 22.565 ;
        RECT 7.850 21.845 8.180 22.225 ;
        RECT 8.395 22.015 8.565 22.395 ;
        RECT 9.750 21.845 10.085 22.350 ;
        RECT 10.255 22.040 10.495 22.415 ;
        RECT 10.980 22.370 11.150 22.705 ;
        RECT 12.140 22.535 12.315 23.340 ;
        RECT 12.505 23.305 15.095 24.395 ;
        RECT 15.265 23.885 15.525 24.395 ;
        RECT 10.775 22.175 11.150 22.370 ;
        RECT 10.775 22.030 10.945 22.175 ;
        RECT 11.510 21.845 11.905 22.340 ;
        RECT 12.075 22.015 12.315 22.535 ;
        RECT 12.505 22.615 13.715 23.135 ;
        RECT 13.885 22.785 15.095 23.305 ;
        RECT 15.265 22.835 15.605 23.715 ;
        RECT 15.775 23.005 15.945 24.225 ;
        RECT 16.185 23.890 16.800 24.395 ;
        RECT 16.185 23.355 16.435 23.720 ;
        RECT 16.605 23.715 16.800 23.890 ;
        RECT 16.970 23.885 17.445 24.225 ;
        RECT 17.615 23.850 17.830 24.395 ;
        RECT 16.605 23.525 16.935 23.715 ;
        RECT 17.155 23.355 17.870 23.650 ;
        RECT 18.040 23.525 18.315 24.225 ;
        RECT 16.185 23.185 17.975 23.355 ;
        RECT 15.775 22.755 16.570 23.005 ;
        RECT 15.775 22.665 16.025 22.755 ;
        RECT 12.505 21.845 15.095 22.615 ;
        RECT 15.265 21.845 15.525 22.665 ;
        RECT 15.695 22.245 16.025 22.665 ;
        RECT 16.740 22.330 16.995 23.185 ;
        RECT 16.205 22.065 16.995 22.330 ;
        RECT 17.165 22.485 17.575 23.005 ;
        RECT 17.745 22.755 17.975 23.185 ;
        RECT 18.145 22.495 18.315 23.525 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 19.030 23.775 19.205 24.225 ;
        RECT 19.375 23.955 19.705 24.395 ;
        RECT 20.010 23.805 20.180 24.225 ;
        RECT 20.415 23.985 21.085 24.395 ;
        RECT 21.300 23.805 21.470 24.225 ;
        RECT 21.670 23.985 22.000 24.395 ;
        RECT 19.030 23.605 19.660 23.775 ;
        RECT 18.945 22.755 19.310 23.435 ;
        RECT 19.490 23.085 19.660 23.605 ;
        RECT 20.010 23.635 22.025 23.805 ;
        RECT 19.490 22.755 19.840 23.085 ;
        RECT 19.490 22.585 19.660 22.755 ;
        RECT 17.165 22.065 17.365 22.485 ;
        RECT 17.555 21.845 17.885 22.305 ;
        RECT 18.055 22.015 18.315 22.495 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 19.030 22.415 19.660 22.585 ;
        RECT 19.030 22.015 19.205 22.415 ;
        RECT 20.010 22.345 20.180 23.635 ;
        RECT 19.375 21.845 19.705 22.225 ;
        RECT 19.950 22.015 20.180 22.345 ;
        RECT 20.380 22.180 20.660 23.455 ;
        RECT 20.885 22.355 21.155 23.455 ;
        RECT 21.345 22.425 21.685 23.455 ;
        RECT 21.855 23.085 22.025 23.635 ;
        RECT 22.195 23.255 22.455 24.225 ;
        RECT 21.855 22.755 22.115 23.085 ;
        RECT 22.285 22.565 22.455 23.255 ;
        RECT 20.845 22.185 21.155 22.355 ;
        RECT 20.885 22.180 21.155 22.185 ;
        RECT 21.615 21.845 21.945 22.225 ;
        RECT 22.115 22.100 22.455 22.565 ;
        RECT 23.135 23.380 23.390 24.220 ;
        RECT 23.565 23.575 23.895 24.395 ;
        RECT 24.135 23.405 24.345 24.220 ;
        RECT 22.115 22.055 22.450 22.100 ;
        RECT 23.135 22.015 23.465 23.380 ;
        RECT 23.695 23.225 24.345 23.405 ;
        RECT 23.695 22.585 23.915 23.225 ;
        RECT 24.515 23.050 24.720 24.225 ;
        RECT 24.290 22.810 24.720 23.050 ;
        RECT 24.890 22.810 25.220 24.225 ;
        RECT 25.400 22.755 25.680 24.225 ;
        RECT 25.860 23.425 26.145 24.220 ;
        RECT 26.325 23.595 26.540 24.395 ;
        RECT 26.720 23.425 26.990 24.220 ;
        RECT 27.230 23.970 27.565 24.395 ;
        RECT 27.735 23.790 27.920 24.195 ;
        RECT 25.860 23.255 26.990 23.425 ;
        RECT 27.255 23.615 27.920 23.790 ;
        RECT 28.125 23.615 28.455 24.395 ;
        RECT 25.905 22.755 26.290 23.085 ;
        RECT 26.510 22.785 27.010 23.050 ;
        RECT 25.985 22.605 26.290 22.755 ;
        RECT 23.695 22.415 25.805 22.585 ;
        RECT 23.695 22.410 24.915 22.415 ;
        RECT 23.635 21.845 24.310 22.230 ;
        RECT 24.585 22.020 24.915 22.410 ;
        RECT 25.085 21.845 25.430 22.245 ;
        RECT 25.600 22.020 25.805 22.415 ;
        RECT 25.985 22.045 26.540 22.605 ;
        RECT 27.255 22.585 27.595 23.615 ;
        RECT 28.625 23.425 28.895 24.195 ;
        RECT 27.765 23.255 28.895 23.425 ;
        RECT 29.155 23.465 29.325 24.225 ;
        RECT 29.540 23.635 29.870 24.395 ;
        RECT 29.155 23.295 29.870 23.465 ;
        RECT 30.040 23.320 30.295 24.225 ;
        RECT 27.765 22.755 28.015 23.255 ;
        RECT 26.715 21.845 26.955 22.520 ;
        RECT 27.255 22.415 27.940 22.585 ;
        RECT 28.195 22.505 28.555 23.085 ;
        RECT 27.230 21.845 27.565 22.245 ;
        RECT 27.735 22.015 27.940 22.415 ;
        RECT 28.725 22.345 28.895 23.255 ;
        RECT 29.065 22.745 29.420 23.115 ;
        RECT 29.700 23.085 29.870 23.295 ;
        RECT 29.700 22.755 29.955 23.085 ;
        RECT 29.700 22.565 29.870 22.755 ;
        RECT 30.125 22.590 30.295 23.320 ;
        RECT 30.470 23.245 30.730 24.395 ;
        RECT 30.905 23.675 31.365 24.225 ;
        RECT 31.555 23.675 31.885 24.395 ;
        RECT 28.150 21.845 28.425 22.325 ;
        RECT 28.635 22.015 28.895 22.345 ;
        RECT 29.155 22.395 29.870 22.565 ;
        RECT 29.155 22.015 29.325 22.395 ;
        RECT 29.540 21.845 29.870 22.225 ;
        RECT 30.040 22.015 30.295 22.590 ;
        RECT 30.470 21.845 30.730 22.685 ;
        RECT 30.905 22.305 31.155 23.675 ;
        RECT 32.085 23.505 32.385 24.055 ;
        RECT 32.555 23.725 32.835 24.395 ;
        RECT 33.700 23.595 33.950 24.395 ;
        RECT 34.120 23.765 34.450 24.225 ;
        RECT 34.620 23.935 34.835 24.395 ;
        RECT 34.120 23.595 35.290 23.765 ;
        RECT 31.445 23.335 32.385 23.505 ;
        RECT 31.445 23.085 31.615 23.335 ;
        RECT 32.755 23.085 33.020 23.445 ;
        RECT 33.210 23.425 33.490 23.585 ;
        RECT 33.210 23.255 34.545 23.425 ;
        RECT 31.325 22.755 31.615 23.085 ;
        RECT 31.785 22.835 32.125 23.085 ;
        RECT 32.345 22.835 33.020 23.085 ;
        RECT 34.375 23.085 34.545 23.255 ;
        RECT 33.210 22.835 33.560 23.075 ;
        RECT 33.730 22.835 34.205 23.075 ;
        RECT 34.375 22.835 34.750 23.085 ;
        RECT 31.445 22.665 31.615 22.755 ;
        RECT 34.375 22.665 34.545 22.835 ;
        RECT 31.445 22.475 32.835 22.665 ;
        RECT 30.905 22.015 31.465 22.305 ;
        RECT 31.635 21.845 31.885 22.305 ;
        RECT 32.505 22.115 32.835 22.475 ;
        RECT 33.210 22.495 34.545 22.665 ;
        RECT 33.210 22.285 33.480 22.495 ;
        RECT 34.920 22.305 35.290 23.595 ;
        RECT 35.505 23.305 37.175 24.395 ;
        RECT 33.700 21.845 34.030 22.305 ;
        RECT 34.540 22.015 35.290 22.305 ;
        RECT 35.505 22.615 36.255 23.135 ;
        RECT 36.425 22.785 37.175 23.305 ;
        RECT 37.805 23.545 38.145 24.185 ;
        RECT 38.315 23.935 38.560 24.395 ;
        RECT 38.735 23.765 38.985 24.225 ;
        RECT 39.175 24.015 39.845 24.395 ;
        RECT 40.045 23.765 40.295 24.225 ;
        RECT 38.735 23.595 40.295 23.765 ;
        RECT 35.505 21.845 37.175 22.615 ;
        RECT 37.805 22.430 37.975 23.545 ;
        RECT 41.055 23.425 41.225 24.225 ;
        RECT 38.285 23.255 41.225 23.425 ;
        RECT 38.285 23.085 38.455 23.255 ;
        RECT 41.490 23.245 41.750 24.395 ;
        RECT 41.925 23.320 42.180 24.225 ;
        RECT 42.350 23.635 42.680 24.395 ;
        RECT 42.895 23.465 43.065 24.225 ;
        RECT 38.145 22.755 38.455 23.085 ;
        RECT 38.625 22.755 38.960 23.085 ;
        RECT 38.285 22.585 38.455 22.755 ;
        RECT 37.805 22.015 38.115 22.430 ;
        RECT 38.285 22.415 38.980 22.585 ;
        RECT 39.230 22.510 39.425 23.085 ;
        RECT 39.685 22.755 40.030 23.085 ;
        RECT 40.340 22.755 40.815 23.085 ;
        RECT 41.070 22.755 41.255 23.085 ;
        RECT 39.685 22.525 39.875 22.755 ;
        RECT 38.310 21.845 38.640 22.225 ;
        RECT 38.810 22.185 38.980 22.415 ;
        RECT 40.045 22.415 41.225 22.585 ;
        RECT 40.045 22.185 40.215 22.415 ;
        RECT 38.810 22.015 40.215 22.185 ;
        RECT 40.485 21.845 40.815 22.245 ;
        RECT 41.055 22.015 41.225 22.415 ;
        RECT 41.490 21.845 41.750 22.685 ;
        RECT 41.925 22.590 42.095 23.320 ;
        RECT 42.350 23.295 43.065 23.465 ;
        RECT 42.350 23.085 42.520 23.295 ;
        RECT 44.245 23.230 44.535 24.395 ;
        RECT 44.705 23.305 46.375 24.395 ;
        RECT 42.265 22.755 42.520 23.085 ;
        RECT 41.925 22.015 42.180 22.590 ;
        RECT 42.350 22.565 42.520 22.755 ;
        RECT 42.800 22.745 43.155 23.115 ;
        RECT 44.705 22.615 45.455 23.135 ;
        RECT 45.625 22.785 46.375 23.305 ;
        RECT 47.005 23.795 47.265 24.215 ;
        RECT 47.435 23.965 47.765 24.395 ;
        RECT 48.455 23.965 49.200 24.135 ;
        RECT 47.005 23.625 48.860 23.795 ;
        RECT 42.350 22.395 43.065 22.565 ;
        RECT 42.350 21.845 42.680 22.225 ;
        RECT 42.895 22.015 43.065 22.395 ;
        RECT 44.245 21.845 44.535 22.570 ;
        RECT 44.705 21.845 46.375 22.615 ;
        RECT 47.005 22.585 47.180 23.625 ;
        RECT 47.350 22.755 47.700 23.455 ;
        RECT 47.915 23.285 48.520 23.455 ;
        RECT 47.870 22.755 48.160 23.085 ;
        RECT 48.330 23.005 48.520 23.285 ;
        RECT 48.690 23.345 48.860 23.625 ;
        RECT 49.030 23.715 49.200 23.965 ;
        RECT 49.425 23.885 50.065 24.215 ;
        RECT 49.030 23.545 50.065 23.715 ;
        RECT 50.235 23.595 50.515 24.395 ;
        RECT 49.895 23.425 50.065 23.545 ;
        RECT 48.690 23.175 49.340 23.345 ;
        RECT 49.895 23.255 50.555 23.425 ;
        RECT 50.725 23.255 51.000 24.225 ;
        RECT 48.330 22.835 48.775 23.005 ;
        RECT 48.330 22.585 48.520 22.835 ;
        RECT 49.170 22.755 49.340 23.175 ;
        RECT 50.385 23.085 50.555 23.255 ;
        RECT 49.560 22.755 50.215 23.085 ;
        RECT 50.385 22.755 50.660 23.085 ;
        RECT 50.385 22.585 50.555 22.755 ;
        RECT 47.005 22.210 47.325 22.585 ;
        RECT 47.580 21.845 47.750 22.585 ;
        RECT 48.000 22.415 48.520 22.585 ;
        RECT 48.945 22.415 50.555 22.585 ;
        RECT 50.830 22.520 51.000 23.255 ;
        RECT 51.170 23.200 51.340 24.395 ;
        RECT 51.610 23.825 51.930 24.225 ;
        RECT 51.610 23.375 51.780 23.825 ;
        RECT 52.100 23.595 52.410 24.395 ;
        RECT 52.580 23.765 52.910 24.225 ;
        RECT 53.080 23.935 53.250 24.395 ;
        RECT 53.420 23.765 53.750 24.225 ;
        RECT 53.920 23.935 54.170 24.395 ;
        RECT 54.360 23.935 54.610 24.395 ;
        RECT 52.580 23.715 53.750 23.765 ;
        RECT 54.780 23.765 55.030 24.225 ;
        RECT 55.280 23.935 55.570 24.395 ;
        RECT 54.780 23.715 55.570 23.765 ;
        RECT 52.580 23.545 55.570 23.715 ;
        RECT 55.370 23.375 55.570 23.545 ;
        RECT 51.610 23.205 55.170 23.375 ;
        RECT 55.345 23.205 55.570 23.375 ;
        RECT 55.745 23.305 56.955 24.395 ;
        RECT 48.000 22.210 48.170 22.415 ;
        RECT 48.415 21.845 48.770 22.245 ;
        RECT 48.945 22.065 49.115 22.415 ;
        RECT 49.315 21.845 49.645 22.245 ;
        RECT 49.815 22.065 49.985 22.415 ;
        RECT 50.155 21.845 50.535 22.245 ;
        RECT 50.725 22.175 51.000 22.520 ;
        RECT 51.170 21.845 51.340 22.785 ;
        RECT 51.610 22.415 51.780 23.205 ;
        RECT 51.950 22.835 52.300 23.035 ;
        RECT 52.580 22.835 53.260 23.035 ;
        RECT 53.470 22.835 54.660 23.035 ;
        RECT 54.840 22.835 55.170 23.205 ;
        RECT 55.370 22.665 55.570 23.205 ;
        RECT 51.610 22.015 51.930 22.415 ;
        RECT 52.100 21.845 52.410 22.665 ;
        RECT 52.580 22.475 54.270 22.665 ;
        RECT 52.580 22.015 52.910 22.475 ;
        RECT 53.520 22.395 54.270 22.475 ;
        RECT 53.080 21.845 53.330 22.305 ;
        RECT 54.440 22.225 54.610 22.665 ;
        RECT 54.780 22.395 55.570 22.665 ;
        RECT 55.745 22.595 56.265 23.135 ;
        RECT 56.435 22.765 56.955 23.305 ;
        RECT 57.135 23.445 57.410 24.215 ;
        RECT 57.580 23.785 57.910 24.215 ;
        RECT 58.080 23.955 58.275 24.395 ;
        RECT 58.455 23.785 58.785 24.215 ;
        RECT 58.965 23.960 64.310 24.395 ;
        RECT 64.485 23.960 69.830 24.395 ;
        RECT 57.580 23.615 58.785 23.785 ;
        RECT 57.135 23.255 57.720 23.445 ;
        RECT 57.890 23.285 58.785 23.615 ;
        RECT 53.520 22.015 55.570 22.225 ;
        RECT 55.745 21.845 56.955 22.595 ;
        RECT 57.135 22.435 57.375 23.085 ;
        RECT 57.545 22.585 57.720 23.255 ;
        RECT 57.890 22.755 58.305 23.085 ;
        RECT 58.485 22.755 58.780 23.085 ;
        RECT 57.545 22.405 57.875 22.585 ;
        RECT 57.150 21.845 57.480 22.235 ;
        RECT 57.650 22.025 57.875 22.405 ;
        RECT 58.075 22.135 58.305 22.755 ;
        RECT 58.485 21.845 58.785 22.575 ;
        RECT 60.550 22.390 60.890 23.220 ;
        RECT 62.370 22.710 62.720 23.960 ;
        RECT 66.070 22.390 66.410 23.220 ;
        RECT 67.890 22.710 68.240 23.960 ;
        RECT 70.005 23.230 70.295 24.395 ;
        RECT 70.465 23.320 70.735 24.225 ;
        RECT 70.905 23.635 71.235 24.395 ;
        RECT 71.415 23.465 71.585 24.225 ;
        RECT 58.965 21.845 64.310 22.390 ;
        RECT 64.485 21.845 69.830 22.390 ;
        RECT 70.005 21.845 70.295 22.570 ;
        RECT 70.465 22.520 70.635 23.320 ;
        RECT 70.920 23.295 71.585 23.465 ;
        RECT 72.765 23.320 73.035 24.225 ;
        RECT 73.205 23.635 73.535 24.395 ;
        RECT 73.715 23.465 73.895 24.225 ;
        RECT 70.920 23.150 71.090 23.295 ;
        RECT 70.805 22.820 71.090 23.150 ;
        RECT 70.920 22.565 71.090 22.820 ;
        RECT 71.325 22.745 71.655 23.115 ;
        RECT 70.465 22.015 70.725 22.520 ;
        RECT 70.920 22.395 71.585 22.565 ;
        RECT 70.905 21.845 71.235 22.225 ;
        RECT 71.415 22.015 71.585 22.395 ;
        RECT 72.765 22.520 72.945 23.320 ;
        RECT 73.220 23.295 73.895 23.465 ;
        RECT 74.225 23.465 74.405 24.225 ;
        RECT 74.585 23.635 74.915 24.395 ;
        RECT 74.225 23.295 74.900 23.465 ;
        RECT 75.085 23.320 75.355 24.225 ;
        RECT 73.220 23.150 73.390 23.295 ;
        RECT 73.115 22.820 73.390 23.150 ;
        RECT 74.730 23.150 74.900 23.295 ;
        RECT 73.220 22.565 73.390 22.820 ;
        RECT 73.615 22.745 73.955 23.115 ;
        RECT 74.165 22.745 74.505 23.115 ;
        RECT 74.730 22.820 75.005 23.150 ;
        RECT 74.730 22.565 74.900 22.820 ;
        RECT 72.765 22.015 73.025 22.520 ;
        RECT 73.220 22.395 73.885 22.565 ;
        RECT 73.205 21.845 73.535 22.225 ;
        RECT 73.715 22.015 73.885 22.395 ;
        RECT 74.235 22.395 74.900 22.565 ;
        RECT 75.175 22.520 75.355 23.320 ;
        RECT 75.525 23.305 76.735 24.395 ;
        RECT 75.525 22.765 76.045 23.305 ;
        RECT 76.215 22.595 76.735 23.135 ;
        RECT 74.235 22.015 74.405 22.395 ;
        RECT 74.585 21.845 74.915 22.225 ;
        RECT 75.095 22.015 75.355 22.520 ;
        RECT 75.525 21.845 76.735 22.595 ;
        RECT 5.520 21.675 76.820 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 7.945 20.855 8.175 21.675 ;
        RECT 8.345 20.875 8.675 21.505 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 7.925 20.435 8.255 20.685 ;
        RECT 8.425 20.275 8.675 20.875 ;
        RECT 8.845 20.855 9.055 21.675 ;
        RECT 9.285 21.000 9.545 21.505 ;
        RECT 9.725 21.295 10.055 21.675 ;
        RECT 10.235 21.125 10.405 21.505 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 7.945 19.125 8.175 20.265 ;
        RECT 8.345 19.295 8.675 20.275 ;
        RECT 8.845 19.125 9.055 20.265 ;
        RECT 9.285 20.200 9.455 21.000 ;
        RECT 9.740 20.955 10.405 21.125 ;
        RECT 9.740 20.700 9.910 20.955 ;
        RECT 10.665 20.905 14.175 21.675 ;
        RECT 9.625 20.370 9.910 20.700 ;
        RECT 10.145 20.405 10.475 20.775 ;
        RECT 10.665 20.385 12.315 20.905 ;
        RECT 14.805 20.855 15.065 21.675 ;
        RECT 15.235 20.855 15.565 21.275 ;
        RECT 15.745 21.190 16.535 21.455 ;
        RECT 15.315 20.765 15.565 20.855 ;
        RECT 9.740 20.225 9.910 20.370 ;
        RECT 9.285 19.295 9.555 20.200 ;
        RECT 9.740 20.055 10.405 20.225 ;
        RECT 12.485 20.215 14.175 20.735 ;
        RECT 9.725 19.125 10.055 19.885 ;
        RECT 10.235 19.295 10.405 20.055 ;
        RECT 10.665 19.125 14.175 20.215 ;
        RECT 14.805 19.805 15.145 20.685 ;
        RECT 15.315 20.515 16.110 20.765 ;
        RECT 14.805 19.125 15.065 19.635 ;
        RECT 15.315 19.295 15.485 20.515 ;
        RECT 16.280 20.335 16.535 21.190 ;
        RECT 16.705 21.035 16.905 21.455 ;
        RECT 17.095 21.215 17.425 21.675 ;
        RECT 16.705 20.515 17.115 21.035 ;
        RECT 17.595 21.025 17.855 21.505 ;
        RECT 17.285 20.335 17.515 20.765 ;
        RECT 15.725 20.165 17.515 20.335 ;
        RECT 15.725 19.800 15.975 20.165 ;
        RECT 16.145 19.805 16.475 19.995 ;
        RECT 16.695 19.870 17.410 20.165 ;
        RECT 17.685 19.995 17.855 21.025 ;
        RECT 18.025 20.905 21.535 21.675 ;
        RECT 21.705 20.925 22.915 21.675 ;
        RECT 23.110 21.285 23.440 21.675 ;
        RECT 23.610 21.115 23.835 21.495 ;
        RECT 18.025 20.385 19.675 20.905 ;
        RECT 19.845 20.215 21.535 20.735 ;
        RECT 21.705 20.385 22.225 20.925 ;
        RECT 22.395 20.215 22.915 20.755 ;
        RECT 23.095 20.435 23.335 21.085 ;
        RECT 23.505 20.935 23.835 21.115 ;
        RECT 23.505 20.265 23.680 20.935 ;
        RECT 24.035 20.765 24.265 21.385 ;
        RECT 24.445 20.945 24.745 21.675 ;
        RECT 25.855 20.865 26.125 21.675 ;
        RECT 26.295 20.865 26.625 21.505 ;
        RECT 26.795 20.865 27.035 21.675 ;
        RECT 27.225 20.905 30.735 21.675 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 31.825 21.130 37.170 21.675 ;
        RECT 23.850 20.435 24.265 20.765 ;
        RECT 24.445 20.435 24.740 20.765 ;
        RECT 25.845 20.435 26.195 20.685 ;
        RECT 26.365 20.265 26.535 20.865 ;
        RECT 26.705 20.435 27.055 20.685 ;
        RECT 27.225 20.385 28.875 20.905 ;
        RECT 16.145 19.630 16.340 19.805 ;
        RECT 15.725 19.125 16.340 19.630 ;
        RECT 16.510 19.295 16.985 19.635 ;
        RECT 17.155 19.125 17.370 19.670 ;
        RECT 17.580 19.295 17.855 19.995 ;
        RECT 18.025 19.125 21.535 20.215 ;
        RECT 21.705 19.125 22.915 20.215 ;
        RECT 23.095 20.075 23.680 20.265 ;
        RECT 23.095 19.305 23.370 20.075 ;
        RECT 23.850 19.905 24.745 20.235 ;
        RECT 23.540 19.735 24.745 19.905 ;
        RECT 23.540 19.305 23.870 19.735 ;
        RECT 24.040 19.125 24.235 19.565 ;
        RECT 24.415 19.305 24.745 19.735 ;
        RECT 25.855 19.125 26.185 20.265 ;
        RECT 26.365 20.095 27.045 20.265 ;
        RECT 29.045 20.215 30.735 20.735 ;
        RECT 33.410 20.300 33.750 21.130 ;
        RECT 37.805 21.090 38.115 21.505 ;
        RECT 38.310 21.295 38.640 21.675 ;
        RECT 38.810 21.335 40.215 21.505 ;
        RECT 38.810 21.105 38.980 21.335 ;
        RECT 26.715 19.310 27.045 20.095 ;
        RECT 27.225 19.125 30.735 20.215 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 35.230 19.560 35.580 20.810 ;
        RECT 37.805 19.975 37.975 21.090 ;
        RECT 38.285 20.935 38.980 21.105 ;
        RECT 40.045 21.105 40.215 21.335 ;
        RECT 40.485 21.275 40.815 21.675 ;
        RECT 41.055 21.105 41.225 21.505 ;
        RECT 38.285 20.765 38.455 20.935 ;
        RECT 38.145 20.435 38.455 20.765 ;
        RECT 38.625 20.435 38.960 20.765 ;
        RECT 39.230 20.435 39.425 21.010 ;
        RECT 39.685 20.765 39.875 20.995 ;
        RECT 40.045 20.935 41.225 21.105 ;
        RECT 41.520 20.935 42.135 21.505 ;
        RECT 42.305 21.165 42.520 21.675 ;
        RECT 42.750 21.165 43.030 21.495 ;
        RECT 43.210 21.165 43.450 21.675 ;
        RECT 39.685 20.435 40.030 20.765 ;
        RECT 40.340 20.435 40.815 20.765 ;
        RECT 41.070 20.435 41.255 20.765 ;
        RECT 38.285 20.265 38.455 20.435 ;
        RECT 38.285 20.095 41.225 20.265 ;
        RECT 31.825 19.125 37.170 19.560 ;
        RECT 37.805 19.335 38.145 19.975 ;
        RECT 38.735 19.755 40.295 19.925 ;
        RECT 38.315 19.125 38.560 19.585 ;
        RECT 38.735 19.295 38.985 19.755 ;
        RECT 39.175 19.125 39.845 19.505 ;
        RECT 40.045 19.295 40.295 19.755 ;
        RECT 41.055 19.295 41.225 20.095 ;
        RECT 41.520 19.915 41.835 20.935 ;
        RECT 42.005 20.265 42.175 20.765 ;
        RECT 42.425 20.435 42.690 20.995 ;
        RECT 42.860 20.265 43.030 21.165 ;
        RECT 43.200 20.435 43.555 20.995 ;
        RECT 43.805 20.865 44.045 21.675 ;
        RECT 44.215 20.865 44.545 21.505 ;
        RECT 44.715 20.865 44.985 21.675 ;
        RECT 43.785 20.435 44.135 20.685 ;
        RECT 44.305 20.265 44.475 20.865 ;
        RECT 44.645 20.435 44.995 20.685 ;
        RECT 42.005 20.095 43.430 20.265 ;
        RECT 41.520 19.295 42.055 19.915 ;
        RECT 42.225 19.125 42.555 19.925 ;
        RECT 43.040 19.920 43.430 20.095 ;
        RECT 43.795 20.095 44.475 20.265 ;
        RECT 43.795 19.310 44.125 20.095 ;
        RECT 44.655 19.125 44.985 20.265 ;
        RECT 45.165 19.295 45.445 21.395 ;
        RECT 45.675 21.215 45.845 21.675 ;
        RECT 46.115 21.285 47.365 21.465 ;
        RECT 46.500 21.045 46.865 21.115 ;
        RECT 45.615 20.865 46.865 21.045 ;
        RECT 47.035 21.065 47.365 21.285 ;
        RECT 47.535 21.235 47.705 21.675 ;
        RECT 47.875 21.065 48.215 21.480 ;
        RECT 47.035 20.895 48.215 21.065 ;
        RECT 49.305 20.875 49.615 21.675 ;
        RECT 49.820 20.875 50.515 21.505 ;
        RECT 50.685 20.875 51.380 21.505 ;
        RECT 51.585 20.875 51.895 21.675 ;
        RECT 52.065 20.905 54.655 21.675 ;
        RECT 55.295 20.945 55.595 21.675 ;
        RECT 45.615 20.265 45.890 20.865 ;
        RECT 46.060 20.435 46.415 20.685 ;
        RECT 46.610 20.655 47.075 20.685 ;
        RECT 46.605 20.485 47.075 20.655 ;
        RECT 46.610 20.435 47.075 20.485 ;
        RECT 47.245 20.435 47.575 20.685 ;
        RECT 47.750 20.485 48.215 20.685 ;
        RECT 49.315 20.435 49.650 20.705 ;
        RECT 47.395 20.315 47.575 20.435 ;
        RECT 45.615 20.055 47.225 20.265 ;
        RECT 47.395 20.145 47.725 20.315 ;
        RECT 46.815 19.955 47.225 20.055 ;
        RECT 45.635 19.125 46.420 19.885 ;
        RECT 46.815 19.295 47.200 19.955 ;
        RECT 47.525 19.355 47.725 20.145 ;
        RECT 47.895 19.125 48.215 20.305 ;
        RECT 49.820 20.275 49.990 20.875 ;
        RECT 50.160 20.435 50.495 20.685 ;
        RECT 50.705 20.435 51.040 20.685 ;
        RECT 51.210 20.275 51.380 20.875 ;
        RECT 51.550 20.435 51.885 20.705 ;
        RECT 52.065 20.385 53.275 20.905 ;
        RECT 55.775 20.765 56.005 21.385 ;
        RECT 56.205 21.115 56.430 21.495 ;
        RECT 56.600 21.285 56.930 21.675 ;
        RECT 56.205 20.935 56.535 21.115 ;
        RECT 49.305 19.125 49.585 20.265 ;
        RECT 49.755 19.295 50.085 20.275 ;
        RECT 50.255 19.125 50.515 20.265 ;
        RECT 50.685 19.125 50.945 20.265 ;
        RECT 51.115 19.295 51.445 20.275 ;
        RECT 51.615 19.125 51.895 20.265 ;
        RECT 53.445 20.215 54.655 20.735 ;
        RECT 55.300 20.435 55.595 20.765 ;
        RECT 55.775 20.435 56.190 20.765 ;
        RECT 56.360 20.265 56.535 20.935 ;
        RECT 56.705 20.435 56.945 21.085 ;
        RECT 57.125 20.950 57.415 21.675 ;
        RECT 57.605 20.945 57.895 21.675 ;
        RECT 57.595 20.435 57.895 20.765 ;
        RECT 58.075 20.745 58.305 21.385 ;
        RECT 58.485 21.125 58.795 21.495 ;
        RECT 58.975 21.305 59.645 21.675 ;
        RECT 58.485 20.925 59.715 21.125 ;
        RECT 58.075 20.435 58.600 20.745 ;
        RECT 58.780 20.435 59.245 20.745 ;
        RECT 52.065 19.125 54.655 20.215 ;
        RECT 55.295 19.905 56.190 20.235 ;
        RECT 56.360 20.075 56.945 20.265 ;
        RECT 55.295 19.735 56.500 19.905 ;
        RECT 55.295 19.305 55.625 19.735 ;
        RECT 55.805 19.125 56.000 19.565 ;
        RECT 56.170 19.305 56.500 19.735 ;
        RECT 56.670 19.305 56.945 20.075 ;
        RECT 57.125 19.125 57.415 20.290 ;
        RECT 59.425 20.255 59.715 20.925 ;
        RECT 57.605 20.015 58.765 20.255 ;
        RECT 57.605 19.305 57.865 20.015 ;
        RECT 58.035 19.125 58.365 19.835 ;
        RECT 58.535 19.305 58.765 20.015 ;
        RECT 58.945 20.035 59.715 20.255 ;
        RECT 58.945 19.305 59.215 20.035 ;
        RECT 59.395 19.125 59.735 19.855 ;
        RECT 59.905 19.305 60.165 21.495 ;
        RECT 60.345 21.130 65.690 21.675 ;
        RECT 65.865 21.130 71.210 21.675 ;
        RECT 61.930 20.300 62.270 21.130 ;
        RECT 63.750 19.560 64.100 20.810 ;
        RECT 67.450 20.300 67.790 21.130 ;
        RECT 71.385 20.905 74.895 21.675 ;
        RECT 75.525 20.925 76.735 21.675 ;
        RECT 69.270 19.560 69.620 20.810 ;
        RECT 71.385 20.385 73.035 20.905 ;
        RECT 73.205 20.215 74.895 20.735 ;
        RECT 60.345 19.125 65.690 19.560 ;
        RECT 65.865 19.125 71.210 19.560 ;
        RECT 71.385 19.125 74.895 20.215 ;
        RECT 75.525 20.215 76.045 20.755 ;
        RECT 76.215 20.385 76.735 20.925 ;
        RECT 75.525 19.125 76.735 20.215 ;
        RECT 5.520 18.955 76.820 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 6.985 18.520 12.330 18.955 ;
        RECT 12.505 18.520 17.850 18.955 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 8.570 16.950 8.910 17.780 ;
        RECT 10.390 17.270 10.740 18.520 ;
        RECT 14.090 16.950 14.430 17.780 ;
        RECT 15.910 17.270 16.260 18.520 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.945 17.865 22.455 18.955 ;
        RECT 18.945 17.175 20.595 17.695 ;
        RECT 20.765 17.345 22.455 17.865 ;
        RECT 23.545 17.815 23.930 18.775 ;
        RECT 24.145 18.155 24.435 18.955 ;
        RECT 24.605 18.615 25.970 18.785 ;
        RECT 24.605 17.985 24.775 18.615 ;
        RECT 24.100 17.815 24.775 17.985 ;
        RECT 6.985 16.405 12.330 16.950 ;
        RECT 12.505 16.405 17.850 16.950 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 18.945 16.405 22.455 17.175 ;
        RECT 23.545 17.145 23.720 17.815 ;
        RECT 24.100 17.645 24.270 17.815 ;
        RECT 24.945 17.645 25.270 18.445 ;
        RECT 25.640 18.405 25.970 18.615 ;
        RECT 25.640 18.155 26.595 18.405 ;
        RECT 23.905 17.395 24.270 17.645 ;
        RECT 24.465 17.395 24.715 17.645 ;
        RECT 23.905 17.315 24.095 17.395 ;
        RECT 24.465 17.315 24.635 17.395 ;
        RECT 24.925 17.315 25.270 17.645 ;
        RECT 25.440 17.315 25.715 17.980 ;
        RECT 25.900 17.315 26.255 17.980 ;
        RECT 26.425 17.145 26.595 18.155 ;
        RECT 26.765 17.815 27.055 18.955 ;
        RECT 27.230 18.155 27.485 18.955 ;
        RECT 27.685 18.105 28.015 18.785 ;
        RECT 26.780 17.315 27.055 17.645 ;
        RECT 27.230 17.615 27.475 17.975 ;
        RECT 27.665 17.825 28.015 18.105 ;
        RECT 27.665 17.445 27.835 17.825 ;
        RECT 28.195 17.645 28.390 18.695 ;
        RECT 28.570 17.815 28.890 18.955 ;
        RECT 29.065 17.865 32.575 18.955 ;
        RECT 27.315 17.275 27.835 17.445 ;
        RECT 28.005 17.315 28.390 17.645 ;
        RECT 28.570 17.595 28.830 17.645 ;
        RECT 28.570 17.425 28.835 17.595 ;
        RECT 28.570 17.315 28.830 17.425 ;
        RECT 27.315 17.255 27.485 17.275 ;
        RECT 23.545 16.575 24.055 17.145 ;
        RECT 24.600 16.975 26.000 17.145 ;
        RECT 24.225 16.405 24.395 16.965 ;
        RECT 24.600 16.575 24.930 16.975 ;
        RECT 25.105 16.405 25.435 16.805 ;
        RECT 25.670 16.785 26.000 16.975 ;
        RECT 26.170 16.955 26.595 17.145 ;
        RECT 27.285 17.085 27.485 17.255 ;
        RECT 29.065 17.175 30.715 17.695 ;
        RECT 30.885 17.345 32.575 17.865 ;
        RECT 33.205 17.815 33.535 18.955 ;
        RECT 33.705 18.325 34.060 18.785 ;
        RECT 34.230 18.495 34.805 18.955 ;
        RECT 34.975 18.325 35.305 18.785 ;
        RECT 33.705 18.155 35.305 18.325 ;
        RECT 35.505 18.155 35.760 18.955 ;
        RECT 36.425 18.520 41.770 18.955 ;
        RECT 33.705 17.815 33.980 18.155 ;
        RECT 34.160 17.595 34.350 17.975 ;
        RECT 33.205 17.395 34.350 17.595 ;
        RECT 34.530 17.225 34.810 18.155 ;
        RECT 35.930 17.985 36.230 18.180 ;
        RECT 34.980 17.815 36.230 17.985 ;
        RECT 34.980 17.395 35.310 17.815 ;
        RECT 35.540 17.315 35.885 17.645 ;
        RECT 26.765 16.785 27.055 17.055 ;
        RECT 25.670 16.575 27.055 16.785 ;
        RECT 27.315 16.710 27.485 17.085 ;
        RECT 27.675 16.935 28.890 17.105 ;
        RECT 27.675 16.630 27.905 16.935 ;
        RECT 28.075 16.405 28.405 16.765 ;
        RECT 28.600 16.585 28.890 16.935 ;
        RECT 29.065 16.405 32.575 17.175 ;
        RECT 33.205 17.015 34.315 17.225 ;
        RECT 33.205 16.575 33.555 17.015 ;
        RECT 33.725 16.405 33.895 16.845 ;
        RECT 34.065 16.785 34.315 17.015 ;
        RECT 34.485 17.125 34.810 17.225 ;
        RECT 34.485 16.955 34.815 17.125 ;
        RECT 34.985 16.785 35.260 17.225 ;
        RECT 36.060 17.160 36.230 17.815 ;
        RECT 34.065 16.575 35.260 16.785 ;
        RECT 35.495 16.405 35.825 17.145 ;
        RECT 35.995 16.830 36.230 17.160 ;
        RECT 38.010 16.950 38.350 17.780 ;
        RECT 39.830 17.270 40.180 18.520 ;
        RECT 41.945 17.865 43.615 18.955 ;
        RECT 41.945 17.175 42.695 17.695 ;
        RECT 42.865 17.345 43.615 17.865 ;
        RECT 44.245 17.790 44.535 18.955 ;
        RECT 45.625 18.355 45.885 18.775 ;
        RECT 46.055 18.525 46.385 18.955 ;
        RECT 47.050 18.525 47.795 18.695 ;
        RECT 45.625 18.185 47.455 18.355 ;
        RECT 36.425 16.405 41.770 16.950 ;
        RECT 41.945 16.405 43.615 17.175 ;
        RECT 45.625 17.145 45.795 18.185 ;
        RECT 45.965 17.315 46.315 18.015 ;
        RECT 46.530 17.845 47.115 18.015 ;
        RECT 46.485 17.315 46.775 17.645 ;
        RECT 46.945 17.565 47.115 17.845 ;
        RECT 47.285 17.905 47.455 18.185 ;
        RECT 47.625 18.275 47.795 18.525 ;
        RECT 48.020 18.445 48.660 18.775 ;
        RECT 47.625 18.105 48.660 18.275 ;
        RECT 48.830 18.155 49.110 18.955 ;
        RECT 48.490 17.985 48.660 18.105 ;
        RECT 47.285 17.735 47.935 17.905 ;
        RECT 48.490 17.815 49.150 17.985 ;
        RECT 49.320 17.815 49.595 18.785 ;
        RECT 50.230 18.495 50.520 18.955 ;
        RECT 50.770 18.325 51.020 18.785 ;
        RECT 51.190 18.495 51.440 18.955 ;
        RECT 51.630 18.495 51.880 18.955 ;
        RECT 46.945 17.395 47.370 17.565 ;
        RECT 46.945 17.145 47.115 17.395 ;
        RECT 47.765 17.315 47.935 17.735 ;
        RECT 48.980 17.645 49.150 17.815 ;
        RECT 48.155 17.315 48.810 17.645 ;
        RECT 48.980 17.315 49.255 17.645 ;
        RECT 48.980 17.145 49.150 17.315 ;
        RECT 44.245 16.405 44.535 17.130 ;
        RECT 45.625 16.770 45.940 17.145 ;
        RECT 46.195 16.405 46.365 17.145 ;
        RECT 46.615 16.975 47.115 17.145 ;
        RECT 47.555 16.975 49.150 17.145 ;
        RECT 49.425 17.080 49.595 17.815 ;
        RECT 46.615 16.770 46.785 16.975 ;
        RECT 47.010 16.405 47.385 16.805 ;
        RECT 47.555 16.625 47.725 16.975 ;
        RECT 47.910 16.405 48.240 16.805 ;
        RECT 48.410 16.625 48.580 16.975 ;
        RECT 48.750 16.405 49.130 16.805 ;
        RECT 49.320 16.735 49.595 17.080 ;
        RECT 50.230 18.275 51.020 18.325 ;
        RECT 52.050 18.325 52.380 18.785 ;
        RECT 52.550 18.495 52.720 18.955 ;
        RECT 52.890 18.325 53.220 18.785 ;
        RECT 52.050 18.275 53.220 18.325 ;
        RECT 50.230 18.105 53.220 18.275 ;
        RECT 53.390 18.155 53.700 18.955 ;
        RECT 53.870 18.385 54.190 18.785 ;
        RECT 54.365 18.520 59.710 18.955 ;
        RECT 59.885 18.520 65.230 18.955 ;
        RECT 50.230 17.225 50.430 18.105 ;
        RECT 54.020 17.935 54.190 18.385 ;
        RECT 50.630 17.765 54.190 17.935 ;
        RECT 50.630 17.395 50.960 17.765 ;
        RECT 51.140 17.395 52.330 17.595 ;
        RECT 52.540 17.395 53.220 17.595 ;
        RECT 53.500 17.395 53.850 17.595 ;
        RECT 50.230 16.955 51.020 17.225 ;
        RECT 51.190 16.785 51.360 17.225 ;
        RECT 51.530 17.035 53.220 17.225 ;
        RECT 51.530 16.955 52.280 17.035 ;
        RECT 50.230 16.575 52.280 16.785 ;
        RECT 52.470 16.405 52.720 16.865 ;
        RECT 52.890 16.575 53.220 17.035 ;
        RECT 53.390 16.405 53.700 17.225 ;
        RECT 54.020 16.975 54.190 17.765 ;
        RECT 53.870 16.575 54.190 16.975 ;
        RECT 55.950 16.950 56.290 17.780 ;
        RECT 57.770 17.270 58.120 18.520 ;
        RECT 61.470 16.950 61.810 17.780 ;
        RECT 63.290 17.270 63.640 18.520 ;
        RECT 65.405 17.865 68.915 18.955 ;
        RECT 65.405 17.175 67.055 17.695 ;
        RECT 67.225 17.345 68.915 17.865 ;
        RECT 70.005 17.790 70.295 18.955 ;
        RECT 70.465 17.865 73.055 18.955 ;
        RECT 73.690 18.530 74.025 18.955 ;
        RECT 74.195 18.350 74.380 18.755 ;
        RECT 70.465 17.175 71.675 17.695 ;
        RECT 71.845 17.345 73.055 17.865 ;
        RECT 73.715 18.175 74.380 18.350 ;
        RECT 74.585 18.175 74.915 18.955 ;
        RECT 54.365 16.405 59.710 16.950 ;
        RECT 59.885 16.405 65.230 16.950 ;
        RECT 65.405 16.405 68.915 17.175 ;
        RECT 70.005 16.405 70.295 17.130 ;
        RECT 70.465 16.405 73.055 17.175 ;
        RECT 73.715 17.145 74.055 18.175 ;
        RECT 75.085 17.985 75.355 18.755 ;
        RECT 74.225 17.815 75.355 17.985 ;
        RECT 74.225 17.315 74.475 17.815 ;
        RECT 73.715 16.975 74.400 17.145 ;
        RECT 74.655 17.065 75.015 17.645 ;
        RECT 73.690 16.405 74.025 16.805 ;
        RECT 74.195 16.575 74.400 16.975 ;
        RECT 75.185 16.905 75.355 17.815 ;
        RECT 75.525 17.865 76.735 18.955 ;
        RECT 75.525 17.325 76.045 17.865 ;
        RECT 76.215 17.155 76.735 17.695 ;
        RECT 74.610 16.405 74.885 16.885 ;
        RECT 75.095 16.575 75.355 16.905 ;
        RECT 75.525 16.405 76.735 17.155 ;
        RECT 5.520 16.235 76.820 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 6.985 15.690 12.330 16.235 ;
        RECT 12.505 15.690 17.850 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 8.570 14.860 8.910 15.690 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 10.390 14.120 10.740 15.370 ;
        RECT 14.090 14.860 14.430 15.690 ;
        RECT 18.025 15.465 21.535 16.235 ;
        RECT 15.910 14.120 16.260 15.370 ;
        RECT 18.025 14.945 19.675 15.465 ;
        RECT 22.725 15.435 22.895 16.235 ;
        RECT 19.845 14.775 21.535 15.295 ;
        RECT 6.985 13.685 12.330 14.120 ;
        RECT 12.505 13.685 17.850 14.120 ;
        RECT 18.025 13.685 21.535 14.775 ;
        RECT 22.655 13.685 22.905 14.875 ;
        RECT 23.130 13.855 23.345 15.955 ;
        RECT 23.565 15.775 23.745 16.235 ;
        RECT 24.005 15.845 25.270 16.025 ;
        RECT 24.390 15.605 24.755 15.675 ;
        RECT 23.515 15.425 24.755 15.605 ;
        RECT 24.930 15.625 25.270 15.845 ;
        RECT 25.455 15.795 25.625 16.235 ;
        RECT 25.795 15.625 26.130 16.040 ;
        RECT 24.930 15.495 26.130 15.625 ;
        RECT 25.100 15.455 26.130 15.495 ;
        RECT 26.305 15.435 26.615 16.235 ;
        RECT 26.820 15.435 27.515 16.065 ;
        RECT 27.710 15.835 28.040 16.235 ;
        RECT 28.210 15.665 28.380 15.935 ;
        RECT 28.550 15.725 28.865 16.235 ;
        RECT 29.095 15.725 29.385 16.065 ;
        RECT 29.555 15.725 29.795 16.235 ;
        RECT 27.685 15.495 28.380 15.665 ;
        RECT 23.515 14.825 23.795 15.425 ;
        RECT 26.820 15.385 26.995 15.435 ;
        RECT 23.975 14.995 24.330 15.245 ;
        RECT 24.500 14.995 24.965 15.245 ;
        RECT 25.135 14.995 25.465 15.245 ;
        RECT 25.635 15.045 26.130 15.245 ;
        RECT 25.285 14.875 25.465 14.995 ;
        RECT 23.515 14.615 25.115 14.825 ;
        RECT 25.285 14.705 25.640 14.875 ;
        RECT 25.810 14.705 26.130 15.045 ;
        RECT 26.315 14.995 26.650 15.265 ;
        RECT 26.820 14.835 26.990 15.385 ;
        RECT 27.160 14.995 27.495 15.245 ;
        RECT 23.535 13.685 24.335 14.445 ;
        RECT 24.730 13.855 25.115 14.615 ;
        RECT 25.440 13.915 25.640 14.705 ;
        RECT 25.810 13.685 26.130 14.525 ;
        RECT 26.305 13.685 26.585 14.825 ;
        RECT 26.755 13.855 27.085 14.835 ;
        RECT 27.255 13.685 27.515 14.825 ;
        RECT 27.685 14.485 28.115 15.495 ;
        RECT 28.285 14.825 28.455 15.325 ;
        RECT 28.625 14.995 29.035 15.555 ;
        RECT 29.205 14.825 29.385 15.725 ;
        RECT 29.555 15.215 29.750 15.555 ;
        RECT 29.985 15.435 30.680 16.065 ;
        RECT 30.885 15.435 31.195 16.235 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.735 32.085 16.065 ;
        RECT 32.295 15.755 32.570 16.235 ;
        RECT 30.505 15.385 30.680 15.435 ;
        RECT 29.555 15.045 29.755 15.215 ;
        RECT 29.555 14.995 29.750 15.045 ;
        RECT 30.005 14.995 30.340 15.245 ;
        RECT 30.510 14.835 30.680 15.385 ;
        RECT 30.850 14.995 31.185 15.265 ;
        RECT 28.285 14.655 29.745 14.825 ;
        RECT 27.685 14.315 28.460 14.485 ;
        RECT 27.790 13.685 27.960 14.145 ;
        RECT 28.130 13.855 28.460 14.315 ;
        RECT 28.630 13.685 28.800 14.485 ;
        RECT 29.385 14.480 29.745 14.655 ;
        RECT 29.985 13.685 30.245 14.825 ;
        RECT 30.415 13.855 30.745 14.835 ;
        RECT 30.915 13.685 31.195 14.825 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 31.825 14.825 31.995 15.735 ;
        RECT 32.780 15.665 32.985 16.065 ;
        RECT 33.155 15.835 33.490 16.235 ;
        RECT 33.755 15.685 33.925 16.065 ;
        RECT 34.105 15.855 34.435 16.235 ;
        RECT 32.165 14.995 32.525 15.575 ;
        RECT 32.780 15.495 33.465 15.665 ;
        RECT 33.755 15.515 34.420 15.685 ;
        RECT 34.615 15.560 34.875 16.065 ;
        RECT 35.045 15.690 40.390 16.235 ;
        RECT 40.565 15.690 45.910 16.235 ;
        RECT 46.085 15.690 51.430 16.235 ;
        RECT 51.605 15.690 56.950 16.235 ;
        RECT 32.705 14.825 32.955 15.325 ;
        RECT 31.825 14.655 32.955 14.825 ;
        RECT 31.825 13.885 32.095 14.655 ;
        RECT 33.125 14.465 33.465 15.495 ;
        RECT 33.685 14.965 34.015 15.335 ;
        RECT 34.250 15.260 34.420 15.515 ;
        RECT 34.250 14.930 34.535 15.260 ;
        RECT 34.250 14.785 34.420 14.930 ;
        RECT 32.265 13.685 32.595 14.465 ;
        RECT 32.800 14.290 33.465 14.465 ;
        RECT 33.755 14.615 34.420 14.785 ;
        RECT 34.705 14.760 34.875 15.560 ;
        RECT 36.630 14.860 36.970 15.690 ;
        RECT 32.800 13.885 32.985 14.290 ;
        RECT 33.155 13.685 33.490 14.110 ;
        RECT 33.755 13.855 33.925 14.615 ;
        RECT 34.105 13.685 34.435 14.445 ;
        RECT 34.605 13.855 34.875 14.760 ;
        RECT 38.450 14.120 38.800 15.370 ;
        RECT 42.150 14.860 42.490 15.690 ;
        RECT 43.970 14.120 44.320 15.370 ;
        RECT 47.670 14.860 48.010 15.690 ;
        RECT 49.490 14.120 49.840 15.370 ;
        RECT 53.190 14.860 53.530 15.690 ;
        RECT 57.125 15.510 57.415 16.235 ;
        RECT 57.585 15.690 62.930 16.235 ;
        RECT 63.105 15.690 68.450 16.235 ;
        RECT 68.625 15.690 73.970 16.235 ;
        RECT 55.010 14.120 55.360 15.370 ;
        RECT 59.170 14.860 59.510 15.690 ;
        RECT 35.045 13.685 40.390 14.120 ;
        RECT 40.565 13.685 45.910 14.120 ;
        RECT 46.085 13.685 51.430 14.120 ;
        RECT 51.605 13.685 56.950 14.120 ;
        RECT 57.125 13.685 57.415 14.850 ;
        RECT 60.990 14.120 61.340 15.370 ;
        RECT 64.690 14.860 65.030 15.690 ;
        RECT 66.510 14.120 66.860 15.370 ;
        RECT 70.210 14.860 70.550 15.690 ;
        RECT 74.325 15.575 74.665 16.235 ;
        RECT 72.030 14.120 72.380 15.370 ;
        RECT 57.585 13.685 62.930 14.120 ;
        RECT 63.105 13.685 68.450 14.120 ;
        RECT 68.625 13.685 73.970 14.120 ;
        RECT 74.145 13.855 74.665 15.405 ;
        RECT 74.835 14.580 75.355 16.065 ;
        RECT 75.525 15.485 76.735 16.235 ;
        RECT 75.525 14.775 76.045 15.315 ;
        RECT 76.215 14.945 76.735 15.485 ;
        RECT 74.835 13.685 75.165 14.410 ;
        RECT 75.525 13.685 76.735 14.775 ;
        RECT 5.520 13.515 76.820 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 6.985 13.080 12.330 13.515 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 8.570 11.510 8.910 12.340 ;
        RECT 10.390 11.830 10.740 13.080 ;
        RECT 13.425 11.795 13.945 13.345 ;
        RECT 14.115 12.790 14.445 13.515 ;
        RECT 6.985 10.965 12.330 11.510 ;
        RECT 13.605 10.965 13.945 11.625 ;
        RECT 14.115 11.135 14.635 12.620 ;
        RECT 14.805 12.425 18.315 13.515 ;
        RECT 14.805 11.735 16.455 12.255 ;
        RECT 16.625 11.905 18.315 12.425 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 18.945 12.425 22.455 13.515 ;
        RECT 18.945 11.735 20.595 12.255 ;
        RECT 20.765 11.905 22.455 12.425 ;
        RECT 23.175 12.585 23.345 13.345 ;
        RECT 23.525 12.755 23.855 13.515 ;
        RECT 23.175 12.415 23.840 12.585 ;
        RECT 24.025 12.440 24.295 13.345 ;
        RECT 23.670 12.270 23.840 12.415 ;
        RECT 23.105 11.865 23.435 12.235 ;
        RECT 23.670 11.940 23.955 12.270 ;
        RECT 14.805 10.965 18.315 11.735 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 18.945 10.965 22.455 11.735 ;
        RECT 23.670 11.685 23.840 11.940 ;
        RECT 23.175 11.515 23.840 11.685 ;
        RECT 24.125 11.640 24.295 12.440 ;
        RECT 24.465 12.425 25.675 13.515 ;
        RECT 23.175 11.135 23.345 11.515 ;
        RECT 23.525 10.965 23.855 11.345 ;
        RECT 24.035 11.135 24.295 11.640 ;
        RECT 24.465 11.715 24.985 12.255 ;
        RECT 25.155 11.885 25.675 12.425 ;
        RECT 25.845 12.795 26.305 13.345 ;
        RECT 26.495 12.795 26.825 13.515 ;
        RECT 24.465 10.965 25.675 11.715 ;
        RECT 25.845 11.425 26.095 12.795 ;
        RECT 27.025 12.625 27.325 13.175 ;
        RECT 27.495 12.845 27.775 13.515 ;
        RECT 26.385 12.455 27.325 12.625 ;
        RECT 28.235 12.585 28.405 13.345 ;
        RECT 28.620 12.755 28.950 13.515 ;
        RECT 26.385 12.205 26.555 12.455 ;
        RECT 27.695 12.205 27.960 12.565 ;
        RECT 28.235 12.415 28.950 12.585 ;
        RECT 29.120 12.440 29.375 13.345 ;
        RECT 26.265 11.875 26.555 12.205 ;
        RECT 26.725 11.955 27.065 12.205 ;
        RECT 27.285 11.955 27.960 12.205 ;
        RECT 26.385 11.785 26.555 11.875 ;
        RECT 28.145 11.865 28.500 12.235 ;
        RECT 28.780 12.205 28.950 12.415 ;
        RECT 28.780 11.875 29.035 12.205 ;
        RECT 26.385 11.595 27.775 11.785 ;
        RECT 28.780 11.685 28.950 11.875 ;
        RECT 29.205 11.710 29.375 12.440 ;
        RECT 29.550 12.365 29.810 13.515 ;
        RECT 30.065 12.585 30.245 13.345 ;
        RECT 30.425 12.755 30.755 13.515 ;
        RECT 30.065 12.415 30.740 12.585 ;
        RECT 30.925 12.440 31.195 13.345 ;
        RECT 30.570 12.270 30.740 12.415 ;
        RECT 30.005 11.865 30.345 12.235 ;
        RECT 30.570 11.940 30.845 12.270 ;
        RECT 25.845 11.135 26.405 11.425 ;
        RECT 26.575 10.965 26.825 11.425 ;
        RECT 27.445 11.235 27.775 11.595 ;
        RECT 28.235 11.515 28.950 11.685 ;
        RECT 28.235 11.135 28.405 11.515 ;
        RECT 28.620 10.965 28.950 11.345 ;
        RECT 29.120 11.135 29.375 11.710 ;
        RECT 29.550 10.965 29.810 11.805 ;
        RECT 30.570 11.685 30.740 11.940 ;
        RECT 30.075 11.515 30.740 11.685 ;
        RECT 31.015 11.640 31.195 12.440 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 32.745 12.545 33.015 13.315 ;
        RECT 33.185 12.735 33.515 13.515 ;
        RECT 33.720 12.910 33.905 13.315 ;
        RECT 34.075 13.090 34.410 13.515 ;
        RECT 33.720 12.735 34.385 12.910 ;
        RECT 32.745 12.375 33.875 12.545 ;
        RECT 30.075 11.135 30.245 11.515 ;
        RECT 30.425 10.965 30.755 11.345 ;
        RECT 30.935 11.135 31.195 11.640 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 32.745 11.465 32.915 12.375 ;
        RECT 33.085 11.625 33.445 12.205 ;
        RECT 33.625 11.875 33.875 12.375 ;
        RECT 34.045 11.705 34.385 12.735 ;
        RECT 34.585 12.425 35.795 13.515 ;
        RECT 33.700 11.535 34.385 11.705 ;
        RECT 34.585 11.715 35.105 12.255 ;
        RECT 35.275 11.885 35.795 12.425 ;
        RECT 36.055 12.585 36.225 13.345 ;
        RECT 36.440 12.755 36.770 13.515 ;
        RECT 36.055 12.415 36.770 12.585 ;
        RECT 36.940 12.440 37.195 13.345 ;
        RECT 35.965 11.865 36.320 12.235 ;
        RECT 36.600 12.205 36.770 12.415 ;
        RECT 36.600 11.875 36.855 12.205 ;
        RECT 32.745 11.135 33.005 11.465 ;
        RECT 33.215 10.965 33.490 11.445 ;
        RECT 33.700 11.135 33.905 11.535 ;
        RECT 34.075 10.965 34.410 11.365 ;
        RECT 34.585 10.965 35.795 11.715 ;
        RECT 36.600 11.685 36.770 11.875 ;
        RECT 37.025 11.710 37.195 12.440 ;
        RECT 37.370 12.365 37.630 13.515 ;
        RECT 37.805 13.080 43.150 13.515 ;
        RECT 36.055 11.515 36.770 11.685 ;
        RECT 36.055 11.135 36.225 11.515 ;
        RECT 36.440 10.965 36.770 11.345 ;
        RECT 36.940 11.135 37.195 11.710 ;
        RECT 37.370 10.965 37.630 11.805 ;
        RECT 39.390 11.510 39.730 12.340 ;
        RECT 41.210 11.830 41.560 13.080 ;
        RECT 44.245 12.350 44.535 13.515 ;
        RECT 44.705 13.080 50.050 13.515 ;
        RECT 50.225 13.080 55.570 13.515 ;
        RECT 37.805 10.965 43.150 11.510 ;
        RECT 44.245 10.965 44.535 11.690 ;
        RECT 46.290 11.510 46.630 12.340 ;
        RECT 48.110 11.830 48.460 13.080 ;
        RECT 51.810 11.510 52.150 12.340 ;
        RECT 53.630 11.830 53.980 13.080 ;
        RECT 55.745 12.425 56.955 13.515 ;
        RECT 55.745 11.715 56.265 12.255 ;
        RECT 56.435 11.885 56.955 12.425 ;
        RECT 57.125 12.350 57.415 13.515 ;
        RECT 57.585 13.080 62.930 13.515 ;
        RECT 63.105 13.080 68.450 13.515 ;
        RECT 44.705 10.965 50.050 11.510 ;
        RECT 50.225 10.965 55.570 11.510 ;
        RECT 55.745 10.965 56.955 11.715 ;
        RECT 57.125 10.965 57.415 11.690 ;
        RECT 59.170 11.510 59.510 12.340 ;
        RECT 60.990 11.830 61.340 13.080 ;
        RECT 64.690 11.510 65.030 12.340 ;
        RECT 66.510 11.830 66.860 13.080 ;
        RECT 68.625 12.425 69.835 13.515 ;
        RECT 68.625 11.715 69.145 12.255 ;
        RECT 69.315 11.885 69.835 12.425 ;
        RECT 70.005 12.350 70.295 13.515 ;
        RECT 70.465 12.425 73.975 13.515 ;
        RECT 74.145 12.425 75.355 13.515 ;
        RECT 70.465 11.735 72.115 12.255 ;
        RECT 72.285 11.905 73.975 12.425 ;
        RECT 57.585 10.965 62.930 11.510 ;
        RECT 63.105 10.965 68.450 11.510 ;
        RECT 68.625 10.965 69.835 11.715 ;
        RECT 70.005 10.965 70.295 11.690 ;
        RECT 70.465 10.965 73.975 11.735 ;
        RECT 74.145 11.715 74.665 12.255 ;
        RECT 74.835 11.885 75.355 12.425 ;
        RECT 75.525 12.425 76.735 13.515 ;
        RECT 75.525 11.885 76.045 12.425 ;
        RECT 76.215 11.715 76.735 12.255 ;
        RECT 74.145 10.965 75.355 11.715 ;
        RECT 75.525 10.965 76.735 11.715 ;
        RECT 5.520 10.795 76.820 10.965 ;
      LAYER met1 ;
        RECT 11.110 92.720 11.430 92.780 ;
        RECT 73.670 92.720 73.990 92.780 ;
        RECT 11.110 92.580 73.990 92.720 ;
        RECT 11.110 92.520 11.430 92.580 ;
        RECT 73.670 92.520 73.990 92.580 ;
        RECT 10.190 91.020 10.510 91.080 ;
        RECT 32.270 91.020 32.590 91.080 ;
        RECT 10.190 90.880 32.590 91.020 ;
        RECT 10.190 90.820 10.510 90.880 ;
        RECT 32.270 90.820 32.590 90.880 ;
        RECT 4.210 87.620 4.530 87.680 ;
        RECT 9.730 87.620 10.050 87.680 ;
        RECT 4.210 87.480 10.050 87.620 ;
        RECT 4.210 87.420 4.530 87.480 ;
        RECT 9.730 87.420 10.050 87.480 ;
        RECT 23.990 84.900 24.310 84.960 ;
        RECT 69.530 84.900 69.850 84.960 ;
        RECT 23.990 84.760 69.850 84.900 ;
        RECT 23.990 84.700 24.310 84.760 ;
        RECT 69.530 84.700 69.850 84.760 ;
        RECT 12.030 84.220 12.350 84.280 ;
        RECT 41.010 84.220 41.330 84.280 ;
        RECT 12.030 84.080 41.330 84.220 ;
        RECT 12.030 84.020 12.350 84.080 ;
        RECT 41.010 84.020 41.330 84.080 ;
        RECT 23.070 83.880 23.390 83.940 ;
        RECT 56.650 83.880 56.970 83.940 ;
        RECT 23.070 83.740 56.970 83.880 ;
        RECT 23.070 83.680 23.390 83.740 ;
        RECT 56.650 83.680 56.970 83.740 ;
        RECT 19.850 83.540 20.170 83.600 ;
        RECT 41.930 83.540 42.250 83.600 ;
        RECT 19.850 83.400 42.250 83.540 ;
        RECT 19.850 83.340 20.170 83.400 ;
        RECT 41.930 83.340 42.250 83.400 ;
        RECT 26.290 83.200 26.610 83.260 ;
        RECT 26.290 83.060 62.170 83.200 ;
        RECT 26.290 83.000 26.610 83.060 ;
        RECT 62.030 82.920 62.170 83.060 ;
        RECT 22.610 82.860 22.930 82.920 ;
        RECT 48.830 82.860 49.150 82.920 ;
        RECT 22.610 82.720 49.150 82.860 ;
        RECT 62.030 82.720 62.490 82.920 ;
        RECT 22.610 82.660 22.930 82.720 ;
        RECT 48.830 82.660 49.150 82.720 ;
        RECT 62.170 82.660 62.490 82.720 ;
        RECT 18.010 82.520 18.330 82.580 ;
        RECT 21.690 82.520 22.010 82.580 ;
        RECT 34.570 82.520 34.890 82.580 ;
        RECT 18.010 82.380 34.890 82.520 ;
        RECT 18.010 82.320 18.330 82.380 ;
        RECT 21.690 82.320 22.010 82.380 ;
        RECT 34.570 82.320 34.890 82.380 ;
        RECT 41.010 82.520 41.330 82.580 ;
        RECT 59.870 82.520 60.190 82.580 ;
        RECT 41.010 82.380 60.190 82.520 ;
        RECT 41.010 82.320 41.330 82.380 ;
        RECT 59.870 82.320 60.190 82.380 ;
        RECT 16.630 82.180 16.950 82.240 ;
        RECT 37.330 82.180 37.650 82.240 ;
        RECT 16.630 82.040 37.650 82.180 ;
        RECT 16.630 81.980 16.950 82.040 ;
        RECT 37.330 81.980 37.650 82.040 ;
        RECT 43.310 82.180 43.630 82.240 ;
        RECT 70.910 82.180 71.230 82.240 ;
        RECT 43.310 82.040 71.230 82.180 ;
        RECT 43.310 81.980 43.630 82.040 ;
        RECT 70.910 81.980 71.230 82.040 ;
        RECT 5.520 81.360 76.820 81.840 ;
        RECT 6.510 81.160 6.830 81.220 ;
        RECT 7.445 81.160 7.735 81.205 ;
        RECT 6.510 81.020 7.735 81.160 ;
        RECT 6.510 80.960 6.830 81.020 ;
        RECT 7.445 80.975 7.735 81.020 ;
        RECT 12.965 81.160 13.255 81.205 ;
        RECT 20.310 81.160 20.630 81.220 ;
        RECT 22.150 81.160 22.470 81.220 ;
        RECT 36.410 81.160 36.730 81.220 ;
        RECT 54.350 81.160 54.670 81.220 ;
        RECT 12.965 81.020 20.630 81.160 ;
        RECT 12.965 80.975 13.255 81.020 ;
        RECT 20.310 80.960 20.630 81.020 ;
        RECT 20.860 81.020 22.470 81.160 ;
        RECT 11.110 80.620 11.430 80.880 ;
        RECT 12.030 80.620 12.350 80.880 ;
        RECT 20.860 80.820 21.000 81.020 ;
        RECT 22.150 80.960 22.470 81.020 ;
        RECT 22.700 81.020 36.730 81.160 ;
        RECT 22.700 80.820 22.840 81.020 ;
        RECT 36.410 80.960 36.730 81.020 ;
        RECT 42.940 81.020 54.670 81.160 ;
        RECT 13.960 80.680 21.000 80.820 ;
        RECT 21.320 80.680 22.840 80.820 ;
        RECT 23.085 80.820 23.375 80.865 ;
        RECT 31.350 80.820 31.670 80.880 ;
        RECT 23.085 80.680 31.670 80.820 ;
        RECT 5.130 80.480 5.450 80.540 ;
        RECT 8.365 80.480 8.655 80.525 ;
        RECT 5.130 80.340 8.655 80.480 ;
        RECT 5.130 80.280 5.450 80.340 ;
        RECT 8.365 80.295 8.655 80.340 ;
        RECT 10.205 80.480 10.495 80.525 ;
        RECT 11.570 80.480 11.890 80.540 ;
        RECT 13.960 80.525 14.100 80.680 ;
        RECT 10.205 80.340 11.890 80.480 ;
        RECT 10.205 80.295 10.495 80.340 ;
        RECT 11.570 80.280 11.890 80.340 ;
        RECT 13.885 80.295 14.175 80.525 ;
        RECT 15.710 80.280 16.030 80.540 ;
        RECT 16.185 80.480 16.475 80.525 ;
        RECT 16.630 80.480 16.950 80.540 ;
        RECT 16.185 80.340 16.950 80.480 ;
        RECT 16.185 80.295 16.475 80.340 ;
        RECT 16.630 80.280 16.950 80.340 ;
        RECT 17.090 80.280 17.410 80.540 ;
        RECT 18.010 80.280 18.330 80.540 ;
        RECT 20.385 80.480 20.675 80.525 ;
        RECT 21.320 80.480 21.460 80.680 ;
        RECT 23.085 80.635 23.375 80.680 ;
        RECT 31.350 80.620 31.670 80.680 ;
        RECT 20.385 80.340 21.460 80.480 ;
        RECT 20.385 80.295 20.675 80.340 ;
        RECT 21.690 80.280 22.010 80.540 ;
        RECT 22.610 80.480 22.930 80.540 ;
        RECT 23.545 80.480 23.835 80.525 ;
        RECT 22.610 80.340 23.835 80.480 ;
        RECT 22.610 80.280 22.930 80.340 ;
        RECT 23.545 80.295 23.835 80.340 ;
        RECT 24.910 80.280 25.230 80.540 ;
        RECT 26.290 80.280 26.610 80.540 ;
        RECT 28.130 80.480 28.450 80.540 ;
        RECT 29.985 80.480 30.275 80.525 ;
        RECT 33.190 80.480 33.510 80.540 ;
        RECT 28.130 80.340 33.510 80.480 ;
        RECT 28.130 80.280 28.450 80.340 ;
        RECT 29.985 80.295 30.275 80.340 ;
        RECT 33.190 80.280 33.510 80.340 ;
        RECT 41.470 80.280 41.790 80.540 ;
        RECT 42.940 80.525 43.080 81.020 ;
        RECT 54.350 80.960 54.670 81.020 ;
        RECT 54.810 81.160 55.130 81.220 ;
        RECT 58.505 81.160 58.795 81.205 ;
        RECT 54.810 81.020 58.795 81.160 ;
        RECT 54.810 80.960 55.130 81.020 ;
        RECT 58.505 80.975 58.795 81.020 ;
        RECT 74.605 80.975 74.895 81.205 ;
        RECT 51.590 80.820 51.910 80.880 ;
        RECT 74.680 80.820 74.820 80.975 ;
        RECT 51.590 80.680 74.820 80.820 ;
        RECT 51.590 80.620 51.910 80.680 ;
        RECT 42.865 80.295 43.155 80.525 ;
        RECT 44.690 80.480 45.010 80.540 ;
        RECT 45.625 80.480 45.915 80.525 ;
        RECT 44.690 80.340 45.915 80.480 ;
        RECT 44.690 80.280 45.010 80.340 ;
        RECT 45.625 80.295 45.915 80.340 ;
        RECT 56.665 80.480 56.955 80.525 ;
        RECT 56.665 80.340 60.100 80.480 ;
        RECT 56.665 80.295 56.955 80.340 ;
        RECT 9.730 80.140 10.050 80.200 ;
        RECT 20.785 80.140 21.075 80.185 ;
        RECT 21.230 80.140 21.550 80.200 ;
        RECT 9.730 80.000 20.600 80.140 ;
        RECT 9.730 79.940 10.050 80.000 ;
        RECT 6.050 79.800 6.370 79.860 ;
        RECT 9.285 79.800 9.575 79.845 ;
        RECT 6.050 79.660 9.575 79.800 ;
        RECT 6.050 79.600 6.370 79.660 ;
        RECT 9.285 79.615 9.575 79.660 ;
        RECT 14.790 79.600 15.110 79.860 ;
        RECT 19.405 79.800 19.695 79.845 ;
        RECT 19.850 79.800 20.170 79.860 ;
        RECT 19.405 79.660 20.170 79.800 ;
        RECT 20.460 79.800 20.600 80.000 ;
        RECT 20.785 80.000 21.550 80.140 ;
        RECT 20.785 79.955 21.075 80.000 ;
        RECT 21.230 79.940 21.550 80.000 ;
        RECT 22.150 80.140 22.470 80.200 ;
        RECT 24.450 80.140 24.770 80.200 ;
        RECT 22.150 80.000 24.770 80.140 ;
        RECT 22.150 79.940 22.470 80.000 ;
        RECT 24.450 79.940 24.770 80.000 ;
        RECT 25.385 79.955 25.675 80.185 ;
        RECT 25.460 79.800 25.600 79.955 ;
        RECT 29.050 79.940 29.370 80.200 ;
        RECT 29.510 79.940 29.830 80.200 ;
        RECT 30.430 79.940 30.750 80.200 ;
        RECT 30.890 80.140 31.210 80.200 ;
        RECT 32.745 80.140 33.035 80.185 ;
        RECT 30.890 80.000 33.035 80.140 ;
        RECT 30.890 79.940 31.210 80.000 ;
        RECT 32.745 79.955 33.035 80.000 ;
        RECT 45.150 79.940 45.470 80.200 ;
        RECT 46.070 79.940 46.390 80.200 ;
        RECT 46.545 79.955 46.835 80.185 ;
        RECT 57.585 80.140 57.875 80.185 ;
        RECT 58.030 80.140 58.350 80.200 ;
        RECT 59.195 80.140 59.485 80.185 ;
        RECT 57.585 80.000 58.350 80.140 ;
        RECT 57.585 79.955 57.875 80.000 ;
        RECT 26.750 79.800 27.070 79.860 ;
        RECT 20.460 79.660 27.070 79.800 ;
        RECT 19.405 79.615 19.695 79.660 ;
        RECT 19.850 79.600 20.170 79.660 ;
        RECT 26.750 79.600 27.070 79.660 ;
        RECT 27.225 79.800 27.515 79.845 ;
        RECT 38.710 79.800 39.030 79.860 ;
        RECT 46.620 79.800 46.760 79.955 ;
        RECT 58.030 79.940 58.350 80.000 ;
        RECT 58.580 80.000 59.485 80.140 ;
        RECT 59.960 80.140 60.100 80.340 ;
        RECT 60.790 80.280 61.110 80.540 ;
        RECT 71.830 80.480 72.150 80.540 ;
        RECT 72.765 80.480 73.055 80.525 ;
        RECT 71.830 80.340 73.055 80.480 ;
        RECT 71.830 80.280 72.150 80.340 ;
        RECT 72.765 80.295 73.055 80.340 ;
        RECT 73.670 80.280 73.990 80.540 ;
        RECT 66.770 80.140 67.090 80.200 ;
        RECT 59.960 80.000 67.090 80.140 ;
        RECT 27.225 79.660 39.030 79.800 ;
        RECT 27.225 79.615 27.515 79.660 ;
        RECT 38.710 79.600 39.030 79.660 ;
        RECT 41.560 79.660 46.760 79.800 ;
        RECT 47.465 79.800 47.755 79.845 ;
        RECT 53.430 79.800 53.750 79.860 ;
        RECT 47.465 79.660 53.750 79.800 ;
        RECT 17.090 79.460 17.410 79.520 ;
        RECT 21.230 79.460 21.550 79.520 ;
        RECT 17.090 79.320 21.550 79.460 ;
        RECT 17.090 79.260 17.410 79.320 ;
        RECT 21.230 79.260 21.550 79.320 ;
        RECT 22.625 79.460 22.915 79.505 ;
        RECT 27.670 79.460 27.990 79.520 ;
        RECT 22.625 79.320 27.990 79.460 ;
        RECT 22.625 79.275 22.915 79.320 ;
        RECT 27.670 79.260 27.990 79.320 ;
        RECT 28.145 79.460 28.435 79.505 ;
        RECT 41.560 79.460 41.700 79.660 ;
        RECT 47.465 79.615 47.755 79.660 ;
        RECT 53.430 79.600 53.750 79.660 ;
        RECT 53.890 79.800 54.210 79.860 ;
        RECT 58.580 79.800 58.720 80.000 ;
        RECT 59.195 79.955 59.485 80.000 ;
        RECT 66.770 79.940 67.090 80.000 ;
        RECT 70.910 79.940 71.230 80.200 ;
        RECT 71.385 80.140 71.675 80.185 ;
        RECT 73.210 80.140 73.530 80.200 ;
        RECT 71.385 80.000 73.530 80.140 ;
        RECT 71.385 79.955 71.675 80.000 ;
        RECT 73.210 79.940 73.530 80.000 ;
        RECT 59.870 79.800 60.190 79.860 ;
        RECT 71.830 79.800 72.150 79.860 ;
        RECT 53.890 79.660 58.720 79.800 ;
        RECT 59.500 79.660 72.150 79.800 ;
        RECT 53.890 79.600 54.210 79.660 ;
        RECT 28.145 79.320 41.700 79.460 ;
        RECT 28.145 79.275 28.435 79.320 ;
        RECT 41.930 79.260 42.250 79.520 ;
        RECT 50.225 79.460 50.515 79.505 ;
        RECT 58.950 79.460 59.270 79.520 ;
        RECT 59.500 79.505 59.640 79.660 ;
        RECT 59.870 79.600 60.190 79.660 ;
        RECT 71.830 79.600 72.150 79.660 ;
        RECT 50.225 79.320 59.270 79.460 ;
        RECT 50.225 79.275 50.515 79.320 ;
        RECT 58.950 79.260 59.270 79.320 ;
        RECT 59.425 79.275 59.715 79.505 ;
        RECT 66.770 79.460 67.090 79.520 ;
        RECT 67.245 79.460 67.535 79.505 ;
        RECT 66.770 79.320 67.535 79.460 ;
        RECT 66.770 79.260 67.090 79.320 ;
        RECT 67.245 79.275 67.535 79.320 ;
        RECT 5.520 78.640 76.820 79.120 ;
        RECT 16.185 78.440 16.475 78.485 ;
        RECT 17.550 78.440 17.870 78.500 ;
        RECT 27.210 78.440 27.530 78.500 ;
        RECT 16.185 78.300 17.870 78.440 ;
        RECT 16.185 78.255 16.475 78.300 ;
        RECT 17.550 78.240 17.870 78.300 ;
        RECT 20.400 78.300 27.530 78.440 ;
        RECT 11.585 78.100 11.875 78.145 ;
        RECT 20.400 78.100 20.540 78.300 ;
        RECT 27.210 78.240 27.530 78.300 ;
        RECT 27.670 78.440 27.990 78.500 ;
        RECT 34.110 78.440 34.430 78.500 ;
        RECT 27.670 78.300 34.430 78.440 ;
        RECT 27.670 78.240 27.990 78.300 ;
        RECT 34.110 78.240 34.430 78.300 ;
        RECT 41.930 78.440 42.250 78.500 ;
        RECT 64.930 78.440 65.250 78.500 ;
        RECT 41.930 78.300 65.250 78.440 ;
        RECT 41.930 78.240 42.250 78.300 ;
        RECT 64.930 78.240 65.250 78.300 ;
        RECT 69.545 78.440 69.835 78.485 ;
        RECT 73.670 78.440 73.990 78.500 ;
        RECT 69.545 78.300 73.990 78.440 ;
        RECT 69.545 78.255 69.835 78.300 ;
        RECT 73.670 78.240 73.990 78.300 ;
        RECT 45.610 78.100 45.930 78.160 ;
        RECT 11.585 77.960 20.540 78.100 ;
        RECT 20.860 77.960 41.700 78.100 ;
        RECT 11.585 77.915 11.875 77.960 ;
        RECT 9.270 77.760 9.590 77.820 ;
        RECT 9.745 77.760 10.035 77.805 ;
        RECT 17.090 77.760 17.410 77.820 ;
        RECT 9.270 77.620 17.410 77.760 ;
        RECT 9.270 77.560 9.590 77.620 ;
        RECT 9.745 77.575 10.035 77.620 ;
        RECT 17.090 77.560 17.410 77.620 ;
        RECT 8.825 77.420 9.115 77.465 ;
        RECT 8.825 77.280 9.960 77.420 ;
        RECT 8.825 77.235 9.115 77.280 ;
        RECT 9.820 77.140 9.960 77.280 ;
        RECT 11.110 77.220 11.430 77.480 ;
        RECT 12.030 77.220 12.350 77.480 ;
        RECT 12.505 77.420 12.795 77.465 ;
        RECT 12.950 77.420 13.270 77.480 ;
        RECT 12.505 77.280 13.270 77.420 ;
        RECT 12.505 77.235 12.795 77.280 ;
        RECT 12.950 77.220 13.270 77.280 ;
        RECT 13.410 77.220 13.730 77.480 ;
        RECT 17.565 77.420 17.855 77.465 ;
        RECT 19.390 77.420 19.710 77.480 ;
        RECT 20.860 77.465 21.000 77.960 ;
        RECT 21.690 77.760 22.010 77.820 ;
        RECT 23.990 77.760 24.310 77.820 ;
        RECT 33.650 77.760 33.970 77.820 ;
        RECT 41.010 77.760 41.330 77.820 ;
        RECT 21.690 77.620 24.310 77.760 ;
        RECT 21.690 77.560 22.010 77.620 ;
        RECT 23.990 77.560 24.310 77.620 ;
        RECT 24.540 77.620 33.970 77.760 ;
        RECT 20.785 77.420 21.075 77.465 ;
        RECT 17.565 77.280 19.710 77.420 ;
        RECT 17.565 77.235 17.855 77.280 ;
        RECT 19.390 77.220 19.710 77.280 ;
        RECT 19.940 77.280 21.075 77.420 ;
        RECT 9.730 76.880 10.050 77.140 ;
        RECT 14.330 76.880 14.650 77.140 ;
        RECT 14.790 77.080 15.110 77.140 ;
        RECT 16.415 77.080 16.705 77.125 ;
        RECT 19.940 77.080 20.080 77.280 ;
        RECT 20.785 77.235 21.075 77.280 ;
        RECT 21.230 77.220 21.550 77.480 ;
        RECT 22.150 77.220 22.470 77.480 ;
        RECT 24.540 77.465 24.680 77.620 ;
        RECT 33.650 77.560 33.970 77.620 ;
        RECT 35.580 77.620 41.330 77.760 ;
        RECT 22.625 77.420 22.915 77.465 ;
        RECT 23.545 77.420 23.835 77.465 ;
        RECT 22.625 77.280 23.835 77.420 ;
        RECT 22.625 77.235 22.915 77.280 ;
        RECT 23.545 77.235 23.835 77.280 ;
        RECT 24.465 77.235 24.755 77.465 ;
        RECT 25.385 77.420 25.675 77.465 ;
        RECT 30.890 77.420 31.210 77.480 ;
        RECT 35.580 77.465 35.720 77.620 ;
        RECT 41.010 77.560 41.330 77.620 ;
        RECT 25.385 77.280 31.210 77.420 ;
        RECT 25.385 77.235 25.675 77.280 ;
        RECT 14.790 76.940 20.080 77.080 ;
        RECT 20.310 77.080 20.630 77.140 ;
        RECT 25.460 77.080 25.600 77.235 ;
        RECT 30.890 77.220 31.210 77.280 ;
        RECT 35.505 77.235 35.795 77.465 ;
        RECT 35.950 77.220 36.270 77.480 ;
        RECT 36.430 77.235 36.720 77.465 ;
        RECT 38.290 77.420 38.580 77.465 ;
        RECT 38.290 77.280 38.940 77.420 ;
        RECT 38.290 77.235 38.580 77.280 ;
        RECT 20.310 76.940 25.600 77.080 ;
        RECT 25.830 77.080 26.150 77.140 ;
        RECT 26.305 77.080 26.595 77.125 ;
        RECT 27.670 77.080 27.990 77.140 ;
        RECT 35.030 77.080 35.350 77.140 ;
        RECT 25.830 76.940 27.990 77.080 ;
        RECT 14.790 76.880 15.110 76.940 ;
        RECT 16.415 76.895 16.705 76.940 ;
        RECT 20.310 76.880 20.630 76.940 ;
        RECT 25.830 76.880 26.150 76.940 ;
        RECT 26.305 76.895 26.595 76.940 ;
        RECT 27.670 76.880 27.990 76.940 ;
        RECT 28.200 76.940 35.350 77.080 ;
        RECT 7.890 76.540 8.210 76.800 ;
        RECT 12.490 76.740 12.810 76.800 ;
        RECT 12.965 76.740 13.255 76.785 ;
        RECT 12.490 76.600 13.255 76.740 ;
        RECT 12.490 76.540 12.810 76.600 ;
        RECT 12.965 76.555 13.255 76.600 ;
        RECT 19.850 76.540 20.170 76.800 ;
        RECT 20.770 76.740 21.090 76.800 ;
        RECT 24.925 76.740 25.215 76.785 ;
        RECT 28.200 76.740 28.340 76.940 ;
        RECT 35.030 76.880 35.350 76.940 ;
        RECT 20.770 76.600 28.340 76.740 ;
        RECT 29.065 76.740 29.355 76.785 ;
        RECT 29.970 76.740 30.290 76.800 ;
        RECT 29.065 76.600 30.290 76.740 ;
        RECT 20.770 76.540 21.090 76.600 ;
        RECT 24.925 76.555 25.215 76.600 ;
        RECT 29.065 76.555 29.355 76.600 ;
        RECT 29.970 76.540 30.290 76.600 ;
        RECT 30.890 76.740 31.210 76.800 ;
        RECT 36.500 76.740 36.640 77.235 ;
        RECT 36.870 77.080 37.190 77.140 ;
        RECT 37.345 77.080 37.635 77.125 ;
        RECT 36.870 76.940 37.635 77.080 ;
        RECT 36.870 76.880 37.190 76.940 ;
        RECT 37.345 76.895 37.635 76.940 ;
        RECT 37.790 76.880 38.110 77.140 ;
        RECT 38.800 77.080 38.940 77.280 ;
        RECT 40.090 77.220 40.410 77.480 ;
        RECT 40.550 77.220 40.870 77.480 ;
        RECT 41.560 77.465 41.700 77.960 ;
        RECT 45.610 77.960 75.280 78.100 ;
        RECT 45.610 77.900 45.930 77.960 ;
        RECT 47.465 77.760 47.755 77.805 ;
        RECT 47.910 77.760 48.230 77.820 ;
        RECT 61.265 77.760 61.555 77.805 ;
        RECT 47.465 77.620 48.230 77.760 ;
        RECT 47.465 77.575 47.755 77.620 ;
        RECT 47.910 77.560 48.230 77.620 ;
        RECT 48.460 77.620 61.555 77.760 ;
        RECT 41.485 77.235 41.775 77.465 ;
        RECT 41.945 77.420 42.235 77.465 ;
        RECT 48.460 77.420 48.600 77.620 ;
        RECT 61.265 77.575 61.555 77.620 ;
        RECT 62.185 77.760 62.475 77.805 ;
        RECT 68.165 77.760 68.455 77.805 ;
        RECT 62.185 77.620 68.455 77.760 ;
        RECT 62.185 77.575 62.475 77.620 ;
        RECT 68.165 77.575 68.455 77.620 ;
        RECT 70.450 77.560 70.770 77.820 ;
        RECT 41.945 77.280 48.600 77.420 ;
        RECT 48.830 77.420 49.150 77.480 ;
        RECT 51.590 77.420 51.910 77.480 ;
        RECT 48.830 77.280 51.910 77.420 ;
        RECT 41.945 77.235 42.235 77.280 ;
        RECT 41.560 77.080 41.700 77.235 ;
        RECT 48.830 77.220 49.150 77.280 ;
        RECT 51.590 77.220 51.910 77.280 ;
        RECT 52.985 77.420 53.275 77.465 ;
        RECT 54.350 77.420 54.670 77.480 ;
        RECT 52.985 77.280 54.670 77.420 ;
        RECT 52.985 77.235 53.275 77.280 ;
        RECT 54.350 77.220 54.670 77.280 ;
        RECT 55.270 77.420 55.590 77.480 ;
        RECT 57.545 77.430 57.835 77.475 ;
        RECT 57.200 77.420 57.835 77.430 ;
        RECT 55.270 77.290 57.835 77.420 ;
        RECT 55.270 77.280 57.340 77.290 ;
        RECT 55.270 77.220 55.590 77.280 ;
        RECT 57.545 77.245 57.835 77.290 ;
        RECT 58.950 77.220 59.270 77.480 ;
        RECT 59.410 77.420 59.730 77.480 ;
        RECT 60.805 77.420 61.095 77.465 ;
        RECT 59.410 77.280 61.095 77.420 ;
        RECT 59.410 77.220 59.730 77.280 ;
        RECT 60.805 77.235 61.095 77.280 ;
        RECT 62.645 77.420 62.935 77.465 ;
        RECT 64.010 77.420 64.330 77.480 ;
        RECT 62.645 77.280 64.330 77.420 ;
        RECT 62.645 77.235 62.935 77.280 ;
        RECT 64.010 77.220 64.330 77.280 ;
        RECT 64.485 77.420 64.775 77.465 ;
        RECT 66.310 77.420 66.630 77.480 ;
        RECT 66.785 77.420 67.075 77.465 ;
        RECT 64.485 77.280 66.080 77.420 ;
        RECT 64.485 77.235 64.775 77.280 ;
        RECT 46.545 77.080 46.835 77.125 ;
        RECT 51.130 77.080 51.450 77.140 ;
        RECT 52.065 77.080 52.355 77.125 ;
        RECT 38.800 76.940 42.160 77.080 ;
        RECT 42.020 76.800 42.160 76.940 ;
        RECT 46.545 76.940 52.355 77.080 ;
        RECT 46.545 76.895 46.835 76.940 ;
        RECT 51.130 76.880 51.450 76.940 ;
        RECT 52.065 76.895 52.355 76.940 ;
        RECT 56.190 77.080 56.510 77.140 ;
        RECT 58.045 77.080 58.335 77.125 ;
        RECT 64.560 77.080 64.700 77.235 ;
        RECT 56.190 76.940 58.335 77.080 ;
        RECT 56.190 76.880 56.510 76.940 ;
        RECT 58.045 76.895 58.335 76.940 ;
        RECT 61.340 76.940 64.700 77.080 ;
        RECT 30.890 76.600 36.640 76.740 ;
        RECT 30.890 76.540 31.210 76.600 ;
        RECT 39.170 76.540 39.490 76.800 ;
        RECT 41.930 76.540 42.250 76.800 ;
        RECT 42.850 76.540 43.170 76.800 ;
        RECT 52.510 76.740 52.830 76.800 ;
        RECT 53.445 76.740 53.735 76.785 ;
        RECT 52.510 76.600 53.735 76.740 ;
        RECT 52.510 76.540 52.830 76.600 ;
        RECT 53.445 76.555 53.735 76.600 ;
        RECT 55.730 76.740 56.050 76.800 ;
        RECT 57.125 76.740 57.415 76.785 ;
        RECT 58.490 76.740 58.810 76.800 ;
        RECT 55.730 76.600 58.810 76.740 ;
        RECT 55.730 76.540 56.050 76.600 ;
        RECT 57.125 76.555 57.415 76.600 ;
        RECT 58.490 76.540 58.810 76.600 ;
        RECT 58.950 76.740 59.270 76.800 ;
        RECT 59.425 76.740 59.715 76.785 ;
        RECT 58.950 76.600 59.715 76.740 ;
        RECT 58.950 76.540 59.270 76.600 ;
        RECT 59.425 76.555 59.715 76.600 ;
        RECT 59.885 76.740 60.175 76.785 ;
        RECT 61.340 76.740 61.480 76.940 ;
        RECT 64.930 76.880 65.250 77.140 ;
        RECT 65.940 77.080 66.080 77.280 ;
        RECT 66.310 77.280 67.075 77.420 ;
        RECT 66.310 77.220 66.630 77.280 ;
        RECT 66.785 77.235 67.075 77.280 ;
        RECT 67.230 77.220 67.550 77.480 ;
        RECT 68.625 77.235 68.915 77.465 ;
        RECT 67.690 77.080 68.010 77.140 ;
        RECT 65.940 76.940 68.010 77.080 ;
        RECT 67.690 76.880 68.010 76.940 ;
        RECT 59.885 76.600 61.480 76.740 ;
        RECT 61.710 76.740 62.030 76.800 ;
        RECT 68.700 76.740 68.840 77.235 ;
        RECT 72.290 77.220 72.610 77.480 ;
        RECT 72.750 77.220 73.070 77.480 ;
        RECT 75.140 77.465 75.280 77.960 ;
        RECT 75.065 77.235 75.355 77.465 ;
        RECT 61.710 76.600 68.840 76.740 ;
        RECT 70.910 76.740 71.230 76.800 ;
        RECT 73.685 76.740 73.975 76.785 ;
        RECT 70.910 76.600 73.975 76.740 ;
        RECT 59.885 76.555 60.175 76.600 ;
        RECT 61.710 76.540 62.030 76.600 ;
        RECT 70.910 76.540 71.230 76.600 ;
        RECT 73.685 76.555 73.975 76.600 ;
        RECT 74.130 76.540 74.450 76.800 ;
        RECT 5.520 75.920 76.820 76.400 ;
        RECT 14.790 75.520 15.110 75.780 ;
        RECT 20.785 75.720 21.075 75.765 ;
        RECT 21.230 75.720 21.550 75.780 ;
        RECT 22.610 75.720 22.930 75.780 ;
        RECT 20.785 75.580 22.930 75.720 ;
        RECT 20.785 75.535 21.075 75.580 ;
        RECT 21.230 75.520 21.550 75.580 ;
        RECT 22.610 75.520 22.930 75.580 ;
        RECT 23.070 75.520 23.390 75.780 ;
        RECT 24.910 75.520 25.230 75.780 ;
        RECT 25.830 75.720 26.150 75.780 ;
        RECT 31.825 75.720 32.115 75.765 ;
        RECT 25.830 75.580 32.115 75.720 ;
        RECT 25.830 75.520 26.150 75.580 ;
        RECT 31.825 75.535 32.115 75.580 ;
        RECT 34.110 75.720 34.430 75.780 ;
        RECT 37.790 75.720 38.110 75.780 ;
        RECT 34.110 75.580 38.110 75.720 ;
        RECT 14.330 75.380 14.650 75.440 ;
        RECT 15.725 75.380 16.015 75.425 ;
        RECT 14.330 75.240 16.015 75.380 ;
        RECT 14.330 75.180 14.650 75.240 ;
        RECT 15.725 75.195 16.015 75.240 ;
        RECT 18.100 75.240 30.660 75.380 ;
        RECT 12.045 75.040 12.335 75.085 ;
        RECT 15.250 75.040 15.570 75.100 ;
        RECT 18.100 75.085 18.240 75.240 ;
        RECT 12.045 74.900 15.570 75.040 ;
        RECT 12.045 74.855 12.335 74.900 ;
        RECT 15.250 74.840 15.570 74.900 ;
        RECT 17.565 74.855 17.855 75.085 ;
        RECT 18.025 74.855 18.315 75.085 ;
        RECT 19.865 75.040 20.155 75.085 ;
        RECT 20.310 75.040 20.630 75.100 ;
        RECT 19.865 74.900 20.630 75.040 ;
        RECT 19.865 74.855 20.155 74.900 ;
        RECT 10.190 74.500 10.510 74.760 ;
        RECT 17.640 74.700 17.780 74.855 ;
        RECT 20.310 74.840 20.630 74.900 ;
        RECT 21.230 74.840 21.550 75.100 ;
        RECT 21.690 75.040 22.010 75.100 ;
        RECT 22.625 75.040 22.915 75.085 ;
        RECT 21.690 74.900 22.915 75.040 ;
        RECT 21.690 74.840 22.010 74.900 ;
        RECT 22.625 74.855 22.915 74.900 ;
        RECT 23.545 74.855 23.835 75.085 ;
        RECT 25.385 75.040 25.675 75.085 ;
        RECT 27.225 75.040 27.515 75.085 ;
        RECT 27.670 75.040 27.990 75.100 ;
        RECT 25.385 74.900 26.980 75.040 ;
        RECT 25.385 74.855 25.675 74.900 ;
        RECT 23.620 74.700 23.760 74.855 ;
        RECT 24.005 74.700 24.295 74.745 ;
        RECT 17.640 74.560 21.000 74.700 ;
        RECT 23.620 74.560 24.295 74.700 ;
        RECT 26.840 74.700 26.980 74.900 ;
        RECT 27.225 74.900 27.990 75.040 ;
        RECT 27.225 74.855 27.515 74.900 ;
        RECT 27.670 74.840 27.990 74.900 ;
        RECT 28.140 75.040 28.430 75.085 ;
        RECT 28.140 74.900 29.740 75.040 ;
        RECT 28.140 74.855 28.430 74.900 ;
        RECT 26.840 74.560 27.440 74.700 ;
        RECT 13.870 73.820 14.190 74.080 ;
        RECT 14.805 74.020 15.095 74.065 ;
        RECT 18.010 74.020 18.330 74.080 ;
        RECT 14.805 73.880 18.330 74.020 ;
        RECT 20.860 74.020 21.000 74.560 ;
        RECT 24.005 74.515 24.295 74.560 ;
        RECT 22.165 74.360 22.455 74.405 ;
        RECT 23.530 74.360 23.850 74.420 ;
        RECT 22.165 74.220 23.850 74.360 ;
        RECT 22.165 74.175 22.455 74.220 ;
        RECT 23.530 74.160 23.850 74.220 ;
        RECT 26.290 74.360 26.610 74.420 ;
        RECT 26.765 74.360 27.055 74.405 ;
        RECT 26.290 74.220 27.055 74.360 ;
        RECT 26.290 74.160 26.610 74.220 ;
        RECT 26.765 74.175 27.055 74.220 ;
        RECT 24.910 74.020 25.230 74.080 ;
        RECT 20.860 73.880 25.230 74.020 ;
        RECT 27.300 74.020 27.440 74.560 ;
        RECT 28.590 74.500 28.910 74.760 ;
        RECT 29.065 74.515 29.355 74.745 ;
        RECT 29.600 74.700 29.740 74.900 ;
        RECT 29.970 74.840 30.290 75.100 ;
        RECT 30.520 75.040 30.660 75.240 ;
        RECT 30.890 75.180 31.210 75.440 ;
        RECT 31.900 75.380 32.040 75.535 ;
        RECT 34.110 75.520 34.430 75.580 ;
        RECT 37.790 75.520 38.110 75.580 ;
        RECT 41.470 75.720 41.790 75.780 ;
        RECT 44.245 75.720 44.535 75.765 ;
        RECT 41.470 75.580 44.535 75.720 ;
        RECT 41.470 75.520 41.790 75.580 ;
        RECT 44.245 75.535 44.535 75.580 ;
        RECT 45.150 75.720 45.470 75.780 ;
        RECT 67.230 75.720 67.550 75.780 ;
        RECT 70.005 75.720 70.295 75.765 ;
        RECT 45.150 75.580 60.100 75.720 ;
        RECT 43.770 75.380 44.090 75.440 ;
        RECT 31.900 75.240 44.090 75.380 ;
        RECT 44.320 75.380 44.460 75.535 ;
        RECT 45.150 75.520 45.470 75.580 ;
        RECT 57.585 75.380 57.875 75.425 ;
        RECT 44.320 75.240 57.875 75.380 ;
        RECT 59.960 75.380 60.100 75.580 ;
        RECT 67.230 75.580 70.295 75.720 ;
        RECT 67.230 75.520 67.550 75.580 ;
        RECT 70.005 75.535 70.295 75.580 ;
        RECT 72.750 75.720 73.070 75.780 ;
        RECT 73.685 75.720 73.975 75.765 ;
        RECT 72.750 75.580 73.975 75.720 ;
        RECT 72.750 75.520 73.070 75.580 ;
        RECT 73.685 75.535 73.975 75.580 ;
        RECT 60.790 75.380 61.110 75.440 ;
        RECT 59.960 75.240 61.110 75.380 ;
        RECT 43.770 75.180 44.090 75.240 ;
        RECT 57.585 75.195 57.875 75.240 ;
        RECT 60.790 75.180 61.110 75.240 ;
        RECT 62.630 75.380 62.950 75.440 ;
        RECT 70.465 75.380 70.755 75.425 ;
        RECT 62.630 75.240 70.755 75.380 ;
        RECT 62.630 75.180 62.950 75.240 ;
        RECT 70.465 75.195 70.755 75.240 ;
        RECT 32.745 75.040 33.035 75.085 ;
        RECT 30.520 74.900 33.035 75.040 ;
        RECT 32.745 74.855 33.035 74.900 ;
        RECT 33.190 75.040 33.510 75.100 ;
        RECT 48.830 75.040 49.150 75.100 ;
        RECT 33.190 74.900 49.150 75.040 ;
        RECT 33.190 74.840 33.510 74.900 ;
        RECT 48.830 74.840 49.150 74.900 ;
        RECT 50.670 74.840 50.990 75.100 ;
        RECT 51.145 74.855 51.435 75.085 ;
        RECT 34.110 74.700 34.430 74.760 ;
        RECT 29.600 74.560 34.430 74.700 ;
        RECT 27.670 74.360 27.990 74.420 ;
        RECT 29.140 74.360 29.280 74.515 ;
        RECT 34.110 74.500 34.430 74.560 ;
        RECT 41.010 74.500 41.330 74.760 ;
        RECT 49.290 74.700 49.610 74.760 ;
        RECT 41.560 74.560 49.610 74.700 ;
        RECT 27.670 74.220 29.280 74.360 ;
        RECT 30.430 74.360 30.750 74.420 ;
        RECT 41.560 74.360 41.700 74.560 ;
        RECT 49.290 74.500 49.610 74.560 ;
        RECT 49.750 74.700 50.070 74.760 ;
        RECT 51.250 74.700 51.390 74.855 ;
        RECT 52.970 74.840 53.290 75.100 ;
        RECT 54.810 74.840 55.130 75.100 ;
        RECT 56.190 74.840 56.510 75.100 ;
        RECT 58.490 75.040 58.810 75.100 ;
        RECT 61.710 75.040 62.030 75.100 ;
        RECT 58.490 74.900 62.030 75.040 ;
        RECT 58.490 74.840 58.810 74.900 ;
        RECT 61.710 74.840 62.030 74.900 ;
        RECT 69.085 75.040 69.375 75.085 ;
        RECT 70.910 75.040 71.230 75.100 ;
        RECT 69.085 74.900 71.230 75.040 ;
        RECT 69.085 74.855 69.375 74.900 ;
        RECT 70.910 74.840 71.230 74.900 ;
        RECT 71.830 75.040 72.150 75.100 ;
        RECT 74.145 75.040 74.435 75.085 ;
        RECT 74.590 75.040 74.910 75.100 ;
        RECT 71.830 74.900 74.910 75.040 ;
        RECT 71.830 74.840 72.150 74.900 ;
        RECT 74.145 74.855 74.435 74.900 ;
        RECT 74.590 74.840 74.910 74.900 ;
        RECT 49.750 74.560 51.390 74.700 ;
        RECT 58.950 74.700 59.270 74.760 ;
        RECT 64.470 74.700 64.790 74.760 ;
        RECT 58.950 74.560 64.790 74.700 ;
        RECT 49.750 74.500 50.070 74.560 ;
        RECT 58.950 74.500 59.270 74.560 ;
        RECT 64.470 74.500 64.790 74.560 ;
        RECT 66.785 74.700 67.075 74.745 ;
        RECT 67.230 74.700 67.550 74.760 ;
        RECT 66.785 74.560 67.550 74.700 ;
        RECT 66.785 74.515 67.075 74.560 ;
        RECT 67.230 74.500 67.550 74.560 ;
        RECT 68.625 74.515 68.915 74.745 ;
        RECT 30.430 74.220 41.700 74.360 ;
        RECT 46.990 74.360 47.310 74.420 ;
        RECT 53.445 74.360 53.735 74.405 ;
        RECT 46.990 74.220 53.735 74.360 ;
        RECT 27.670 74.160 27.990 74.220 ;
        RECT 30.430 74.160 30.750 74.220 ;
        RECT 46.990 74.160 47.310 74.220 ;
        RECT 53.445 74.175 53.735 74.220 ;
        RECT 55.270 74.360 55.590 74.420 ;
        RECT 68.700 74.360 68.840 74.515 ;
        RECT 72.290 74.500 72.610 74.760 ;
        RECT 72.765 74.700 73.055 74.745 ;
        RECT 73.670 74.700 73.990 74.760 ;
        RECT 72.765 74.560 73.990 74.700 ;
        RECT 72.765 74.515 73.055 74.560 ;
        RECT 73.670 74.500 73.990 74.560 ;
        RECT 55.270 74.220 68.840 74.360 ;
        RECT 55.270 74.160 55.590 74.220 ;
        RECT 28.130 74.020 28.450 74.080 ;
        RECT 29.510 74.020 29.830 74.080 ;
        RECT 27.300 73.880 29.830 74.020 ;
        RECT 14.805 73.835 15.095 73.880 ;
        RECT 18.010 73.820 18.330 73.880 ;
        RECT 24.910 73.820 25.230 73.880 ;
        RECT 28.130 73.820 28.450 73.880 ;
        RECT 29.510 73.820 29.830 73.880 ;
        RECT 30.890 74.020 31.210 74.080 ;
        RECT 52.065 74.020 52.355 74.065 ;
        RECT 53.890 74.020 54.210 74.080 ;
        RECT 30.890 73.880 54.210 74.020 ;
        RECT 30.890 73.820 31.210 73.880 ;
        RECT 52.065 73.835 52.355 73.880 ;
        RECT 53.890 73.820 54.210 73.880 ;
        RECT 58.490 74.020 58.810 74.080 ;
        RECT 64.025 74.020 64.315 74.065 ;
        RECT 58.490 73.880 64.315 74.020 ;
        RECT 58.490 73.820 58.810 73.880 ;
        RECT 64.025 73.835 64.315 73.880 ;
        RECT 69.530 74.020 69.850 74.080 ;
        RECT 74.605 74.020 74.895 74.065 ;
        RECT 69.530 73.880 74.895 74.020 ;
        RECT 69.530 73.820 69.850 73.880 ;
        RECT 74.605 73.835 74.895 73.880 ;
        RECT 5.520 73.200 76.820 73.680 ;
        RECT 12.505 73.000 12.795 73.045 ;
        RECT 27.670 73.000 27.990 73.060 ;
        RECT 12.505 72.860 27.990 73.000 ;
        RECT 12.505 72.815 12.795 72.860 ;
        RECT 27.670 72.800 27.990 72.860 ;
        RECT 35.490 73.000 35.810 73.060 ;
        RECT 38.265 73.000 38.555 73.045 ;
        RECT 35.490 72.860 38.555 73.000 ;
        RECT 35.490 72.800 35.810 72.860 ;
        RECT 38.265 72.815 38.555 72.860 ;
        RECT 44.690 73.000 45.010 73.060 ;
        RECT 55.270 73.000 55.590 73.060 ;
        RECT 44.690 72.860 55.590 73.000 ;
        RECT 44.690 72.800 45.010 72.860 ;
        RECT 55.270 72.800 55.590 72.860 ;
        RECT 73.670 72.800 73.990 73.060 ;
        RECT 16.645 72.660 16.935 72.705 ;
        RECT 25.830 72.660 26.150 72.720 ;
        RECT 15.340 72.520 16.935 72.660 ;
        RECT 15.340 72.380 15.480 72.520 ;
        RECT 16.645 72.475 16.935 72.520 ;
        RECT 17.640 72.520 26.150 72.660 ;
        RECT 7.430 72.320 7.750 72.380 ;
        RECT 9.285 72.320 9.575 72.365 ;
        RECT 7.430 72.180 9.575 72.320 ;
        RECT 7.430 72.120 7.750 72.180 ;
        RECT 9.285 72.135 9.575 72.180 ;
        RECT 11.125 72.320 11.415 72.365 ;
        RECT 11.125 72.180 15.020 72.320 ;
        RECT 11.125 72.135 11.415 72.180 ;
        RECT 8.810 71.780 9.130 72.040 ;
        RECT 10.205 71.980 10.495 72.025 ;
        RECT 10.650 71.980 10.970 72.040 ;
        RECT 12.950 71.980 13.270 72.040 ;
        RECT 14.880 72.025 15.020 72.180 ;
        RECT 15.250 72.120 15.570 72.380 ;
        RECT 15.710 72.320 16.030 72.380 ;
        RECT 16.185 72.320 16.475 72.365 ;
        RECT 15.710 72.180 16.475 72.320 ;
        RECT 15.710 72.120 16.030 72.180 ;
        RECT 16.185 72.135 16.475 72.180 ;
        RECT 17.090 72.025 17.410 72.040 ;
        RECT 17.640 72.025 17.780 72.520 ;
        RECT 25.830 72.460 26.150 72.520 ;
        RECT 26.750 72.660 27.070 72.720 ;
        RECT 34.110 72.660 34.430 72.720 ;
        RECT 35.965 72.660 36.255 72.705 ;
        RECT 65.865 72.660 66.155 72.705 ;
        RECT 26.750 72.520 31.120 72.660 ;
        RECT 26.750 72.460 27.070 72.520 ;
        RECT 28.590 72.320 28.910 72.380 ;
        RECT 21.320 72.180 28.910 72.320 ;
        RECT 21.320 72.025 21.460 72.180 ;
        RECT 28.590 72.120 28.910 72.180 ;
        RECT 10.205 71.840 10.970 71.980 ;
        RECT 12.755 71.840 13.270 71.980 ;
        RECT 10.205 71.795 10.495 71.840 ;
        RECT 10.650 71.780 10.970 71.840 ;
        RECT 12.950 71.780 13.270 71.840 ;
        RECT 13.425 71.980 13.715 72.025 ;
        RECT 13.425 71.840 14.100 71.980 ;
        RECT 13.425 71.795 13.715 71.840 ;
        RECT 3.750 71.300 4.070 71.360 ;
        RECT 13.960 71.345 14.100 71.840 ;
        RECT 14.805 71.795 15.095 72.025 ;
        RECT 17.005 71.795 17.410 72.025 ;
        RECT 17.565 71.795 17.855 72.025 ;
        RECT 18.025 71.980 18.315 72.025 ;
        RECT 18.025 71.840 21.000 71.980 ;
        RECT 18.025 71.795 18.315 71.840 ;
        RECT 14.880 71.640 15.020 71.795 ;
        RECT 17.090 71.780 17.410 71.795 ;
        RECT 15.250 71.640 15.570 71.700 ;
        RECT 14.880 71.500 15.570 71.640 ;
        RECT 15.250 71.440 15.570 71.500 ;
        RECT 15.725 71.640 16.015 71.685 ;
        RECT 20.860 71.640 21.000 71.840 ;
        RECT 21.245 71.795 21.535 72.025 ;
        RECT 21.690 71.980 22.010 72.040 ;
        RECT 22.165 71.980 22.455 72.025 ;
        RECT 21.690 71.840 22.455 71.980 ;
        RECT 21.690 71.780 22.010 71.840 ;
        RECT 22.165 71.795 22.455 71.840 ;
        RECT 23.070 71.780 23.390 72.040 ;
        RECT 23.530 71.780 23.850 72.040 ;
        RECT 24.910 71.980 25.230 72.040 ;
        RECT 30.430 71.980 30.750 72.040 ;
        RECT 24.910 71.840 30.750 71.980 ;
        RECT 30.980 71.980 31.120 72.520 ;
        RECT 34.110 72.520 36.255 72.660 ;
        RECT 34.110 72.460 34.430 72.520 ;
        RECT 35.965 72.475 36.255 72.520 ;
        RECT 46.620 72.520 66.155 72.660 ;
        RECT 32.270 72.320 32.590 72.380 ;
        RECT 33.650 72.320 33.970 72.380 ;
        RECT 46.085 72.320 46.375 72.365 ;
        RECT 32.270 72.180 36.640 72.320 ;
        RECT 32.270 72.120 32.590 72.180 ;
        RECT 33.650 72.120 33.970 72.180 ;
        RECT 34.125 71.980 34.415 72.025 ;
        RECT 30.980 71.840 34.415 71.980 ;
        RECT 24.910 71.780 25.230 71.840 ;
        RECT 30.430 71.780 30.750 71.840 ;
        RECT 34.125 71.795 34.415 71.840 ;
        RECT 35.030 71.980 35.350 72.040 ;
        RECT 36.500 72.025 36.640 72.180 ;
        RECT 36.960 72.180 46.375 72.320 ;
        RECT 35.505 71.980 35.795 72.025 ;
        RECT 35.030 71.840 35.795 71.980 ;
        RECT 35.030 71.780 35.350 71.840 ;
        RECT 35.505 71.795 35.795 71.840 ;
        RECT 36.425 71.795 36.715 72.025 ;
        RECT 23.620 71.640 23.760 71.780 ;
        RECT 15.725 71.500 20.600 71.640 ;
        RECT 20.860 71.500 23.760 71.640 ;
        RECT 25.830 71.640 26.150 71.700 ;
        RECT 26.750 71.640 27.070 71.700 ;
        RECT 25.830 71.500 27.070 71.640 ;
        RECT 15.725 71.455 16.015 71.500 ;
        RECT 7.905 71.300 8.195 71.345 ;
        RECT 3.750 71.160 8.195 71.300 ;
        RECT 3.750 71.100 4.070 71.160 ;
        RECT 7.905 71.115 8.195 71.160 ;
        RECT 13.885 71.300 14.175 71.345 ;
        RECT 16.630 71.300 16.950 71.360 ;
        RECT 13.885 71.160 16.950 71.300 ;
        RECT 20.460 71.300 20.600 71.500 ;
        RECT 25.830 71.440 26.150 71.500 ;
        RECT 26.750 71.440 27.070 71.500 ;
        RECT 28.130 71.640 28.450 71.700 ;
        RECT 33.650 71.640 33.970 71.700 ;
        RECT 36.960 71.640 37.100 72.180 ;
        RECT 46.085 72.135 46.375 72.180 ;
        RECT 46.620 72.040 46.760 72.520 ;
        RECT 65.865 72.475 66.155 72.520 ;
        RECT 48.370 72.320 48.690 72.380 ;
        RECT 69.085 72.320 69.375 72.365 ;
        RECT 48.370 72.180 69.375 72.320 ;
        RECT 48.370 72.120 48.690 72.180 ;
        RECT 69.085 72.135 69.375 72.180 ;
        RECT 37.330 71.980 37.650 72.040 ;
        RECT 37.805 71.980 38.095 72.025 ;
        RECT 37.330 71.840 38.095 71.980 ;
        RECT 37.330 71.780 37.650 71.840 ;
        RECT 37.805 71.795 38.095 71.840 ;
        RECT 38.710 71.980 39.030 72.040 ;
        RECT 39.185 71.980 39.475 72.025 ;
        RECT 38.710 71.840 39.475 71.980 ;
        RECT 38.710 71.780 39.030 71.840 ;
        RECT 39.185 71.795 39.475 71.840 ;
        RECT 39.630 71.980 39.950 72.040 ;
        RECT 40.565 71.980 40.855 72.025 ;
        RECT 39.630 71.840 40.855 71.980 ;
        RECT 39.630 71.780 39.950 71.840 ;
        RECT 40.565 71.795 40.855 71.840 ;
        RECT 44.230 71.980 44.550 72.040 ;
        RECT 44.705 71.980 44.995 72.025 ;
        RECT 45.150 71.980 45.470 72.040 ;
        RECT 44.230 71.840 45.470 71.980 ;
        RECT 44.230 71.780 44.550 71.840 ;
        RECT 44.705 71.795 44.995 71.840 ;
        RECT 45.150 71.780 45.470 71.840 ;
        RECT 45.610 71.780 45.930 72.040 ;
        RECT 46.530 71.780 46.850 72.040 ;
        RECT 47.005 71.980 47.295 72.025 ;
        RECT 47.450 71.980 47.770 72.040 ;
        RECT 47.005 71.840 47.770 71.980 ;
        RECT 47.005 71.795 47.295 71.840 ;
        RECT 47.450 71.780 47.770 71.840 ;
        RECT 48.830 71.780 49.150 72.040 ;
        RECT 49.765 71.980 50.055 72.025 ;
        RECT 52.050 71.980 52.370 72.040 ;
        RECT 49.765 71.840 52.370 71.980 ;
        RECT 49.765 71.795 50.055 71.840 ;
        RECT 52.050 71.780 52.370 71.840 ;
        RECT 58.030 71.980 58.350 72.040 ;
        RECT 68.625 71.980 68.915 72.025 ;
        RECT 58.030 71.840 68.915 71.980 ;
        RECT 58.030 71.780 58.350 71.840 ;
        RECT 68.625 71.795 68.915 71.840 ;
        RECT 72.290 71.780 72.610 72.040 ;
        RECT 72.765 71.980 73.055 72.025 ;
        RECT 75.050 71.980 75.370 72.040 ;
        RECT 72.765 71.840 75.370 71.980 ;
        RECT 72.765 71.795 73.055 71.840 ;
        RECT 75.050 71.780 75.370 71.840 ;
        RECT 28.130 71.500 33.970 71.640 ;
        RECT 28.130 71.440 28.450 71.500 ;
        RECT 33.650 71.440 33.970 71.500 ;
        RECT 34.200 71.500 37.100 71.640 ;
        RECT 41.010 71.640 41.330 71.700 ;
        RECT 50.225 71.640 50.515 71.685 ;
        RECT 41.010 71.500 50.515 71.640 ;
        RECT 23.530 71.300 23.850 71.360 ;
        RECT 20.460 71.160 23.850 71.300 ;
        RECT 13.885 71.115 14.175 71.160 ;
        RECT 16.630 71.100 16.950 71.160 ;
        RECT 23.530 71.100 23.850 71.160 ;
        RECT 24.005 71.300 24.295 71.345 ;
        RECT 27.210 71.300 27.530 71.360 ;
        RECT 24.005 71.160 27.530 71.300 ;
        RECT 24.005 71.115 24.295 71.160 ;
        RECT 27.210 71.100 27.530 71.160 ;
        RECT 28.590 71.300 28.910 71.360 ;
        RECT 34.200 71.300 34.340 71.500 ;
        RECT 41.010 71.440 41.330 71.500 ;
        RECT 50.225 71.455 50.515 71.500 ;
        RECT 52.510 71.640 52.830 71.700 ;
        RECT 59.425 71.640 59.715 71.685 ;
        RECT 52.510 71.500 59.715 71.640 ;
        RECT 52.510 71.440 52.830 71.500 ;
        RECT 59.425 71.455 59.715 71.500 ;
        RECT 68.150 71.640 68.470 71.700 ;
        RECT 71.830 71.640 72.150 71.700 ;
        RECT 68.150 71.500 72.150 71.640 ;
        RECT 68.150 71.440 68.470 71.500 ;
        RECT 71.830 71.440 72.150 71.500 ;
        RECT 28.590 71.160 34.340 71.300 ;
        RECT 34.570 71.300 34.890 71.360 ;
        RECT 35.490 71.300 35.810 71.360 ;
        RECT 34.570 71.160 35.810 71.300 ;
        RECT 28.590 71.100 28.910 71.160 ;
        RECT 34.570 71.100 34.890 71.160 ;
        RECT 35.490 71.100 35.810 71.160 ;
        RECT 36.410 71.300 36.730 71.360 ;
        RECT 36.885 71.300 37.175 71.345 ;
        RECT 36.410 71.160 37.175 71.300 ;
        RECT 36.410 71.100 36.730 71.160 ;
        RECT 36.885 71.115 37.175 71.160 ;
        RECT 38.250 71.300 38.570 71.360 ;
        RECT 39.645 71.300 39.935 71.345 ;
        RECT 38.250 71.160 39.935 71.300 ;
        RECT 38.250 71.100 38.570 71.160 ;
        RECT 39.645 71.115 39.935 71.160 ;
        RECT 47.910 71.100 48.230 71.360 ;
        RECT 49.290 71.100 49.610 71.360 ;
        RECT 51.130 71.300 51.450 71.360 ;
        RECT 56.665 71.300 56.955 71.345 ;
        RECT 51.130 71.160 56.955 71.300 ;
        RECT 51.130 71.100 51.450 71.160 ;
        RECT 56.665 71.115 56.955 71.160 ;
        RECT 58.950 71.300 59.270 71.360 ;
        RECT 70.465 71.300 70.755 71.345 ;
        RECT 74.145 71.300 74.435 71.345 ;
        RECT 58.950 71.160 74.435 71.300 ;
        RECT 58.950 71.100 59.270 71.160 ;
        RECT 70.465 71.115 70.755 71.160 ;
        RECT 74.145 71.115 74.435 71.160 ;
        RECT 5.520 70.480 76.820 70.960 ;
        RECT 16.630 70.280 16.950 70.340 ;
        RECT 28.145 70.280 28.435 70.325 ;
        RECT 28.590 70.280 28.910 70.340 ;
        RECT 46.530 70.280 46.850 70.340 ;
        RECT 62.170 70.280 62.490 70.340 ;
        RECT 64.025 70.280 64.315 70.325 ;
        RECT 74.130 70.280 74.450 70.340 ;
        RECT 14.420 70.140 15.465 70.280 ;
        RECT 7.430 69.940 7.750 70.000 ;
        RECT 11.125 69.940 11.415 69.985 ;
        RECT 13.760 69.940 14.050 69.985 ;
        RECT 14.420 69.940 14.560 70.140 ;
        RECT 7.430 69.800 11.415 69.940 ;
        RECT 7.430 69.740 7.750 69.800 ;
        RECT 11.125 69.755 11.415 69.800 ;
        RECT 11.660 69.800 14.560 69.940 ;
        RECT 8.825 69.600 9.115 69.645 ;
        RECT 10.190 69.600 10.510 69.660 ;
        RECT 11.660 69.600 11.800 69.800 ;
        RECT 13.760 69.755 14.050 69.800 ;
        RECT 8.825 69.460 10.510 69.600 ;
        RECT 8.825 69.415 9.115 69.460 ;
        RECT 10.190 69.400 10.510 69.460 ;
        RECT 10.740 69.460 11.800 69.600 ;
        RECT 12.950 69.645 13.270 69.660 ;
        RECT 9.270 69.260 9.590 69.320 ;
        RECT 9.745 69.260 10.035 69.305 ;
        RECT 9.270 69.120 10.035 69.260 ;
        RECT 9.270 69.060 9.590 69.120 ;
        RECT 9.745 69.075 10.035 69.120 ;
        RECT 10.740 68.920 10.880 69.460 ;
        RECT 12.950 69.415 13.485 69.645 ;
        RECT 14.345 69.415 14.635 69.645 ;
        RECT 12.950 69.400 13.270 69.415 ;
        RECT 12.030 69.260 12.350 69.320 ;
        RECT 12.505 69.260 12.795 69.305 ;
        RECT 14.420 69.260 14.560 69.415 ;
        RECT 14.790 69.400 15.110 69.660 ;
        RECT 15.325 69.600 15.465 70.140 ;
        RECT 16.630 70.140 25.600 70.280 ;
        RECT 16.630 70.080 16.950 70.140 ;
        RECT 21.705 69.940 21.995 69.985 ;
        RECT 22.610 69.940 22.930 70.000 ;
        RECT 24.925 69.940 25.215 69.985 ;
        RECT 21.705 69.800 25.215 69.940 ;
        RECT 25.460 69.940 25.600 70.140 ;
        RECT 28.145 70.140 28.910 70.280 ;
        RECT 28.145 70.095 28.435 70.140 ;
        RECT 28.590 70.080 28.910 70.140 ;
        RECT 30.060 70.140 46.850 70.280 ;
        RECT 30.060 69.940 30.200 70.140 ;
        RECT 46.530 70.080 46.850 70.140 ;
        RECT 47.080 70.140 55.960 70.280 ;
        RECT 30.445 69.940 30.735 69.985 ;
        RECT 25.460 69.800 28.820 69.940 ;
        RECT 30.060 69.800 30.735 69.940 ;
        RECT 21.705 69.755 21.995 69.800 ;
        RECT 22.610 69.740 22.930 69.800 ;
        RECT 24.925 69.755 25.215 69.800 ;
        RECT 17.105 69.600 17.395 69.645 ;
        RECT 18.945 69.600 19.235 69.645 ;
        RECT 15.325 69.460 17.395 69.600 ;
        RECT 17.105 69.415 17.395 69.460 ;
        RECT 18.100 69.460 19.235 69.600 ;
        RECT 12.030 69.120 12.795 69.260 ;
        RECT 12.030 69.060 12.350 69.120 ;
        RECT 12.505 69.075 12.795 69.120 ;
        RECT 13.040 69.120 14.560 69.260 ;
        RECT 16.630 69.260 16.950 69.320 ;
        RECT 18.100 69.260 18.240 69.460 ;
        RECT 18.945 69.415 19.235 69.460 ;
        RECT 19.865 69.600 20.155 69.645 ;
        RECT 20.310 69.600 20.630 69.660 ;
        RECT 19.865 69.460 20.630 69.600 ;
        RECT 19.865 69.415 20.155 69.460 ;
        RECT 20.310 69.400 20.630 69.460 ;
        RECT 21.230 69.400 21.550 69.660 ;
        RECT 22.150 69.400 22.470 69.660 ;
        RECT 23.085 69.600 23.375 69.645 ;
        RECT 24.465 69.600 24.755 69.645 ;
        RECT 25.370 69.600 25.690 69.660 ;
        RECT 23.085 69.460 24.755 69.600 ;
        RECT 23.085 69.415 23.375 69.460 ;
        RECT 24.465 69.415 24.755 69.460 ;
        RECT 25.000 69.460 25.690 69.600 ;
        RECT 16.630 69.120 18.240 69.260 ;
        RECT 18.470 69.260 18.790 69.320 ;
        RECT 23.160 69.260 23.300 69.415 ;
        RECT 18.470 69.120 23.300 69.260 ;
        RECT 7.980 68.780 10.880 68.920 ;
        RECT 11.570 68.920 11.890 68.980 ;
        RECT 13.040 68.920 13.180 69.120 ;
        RECT 16.630 69.060 16.950 69.120 ;
        RECT 18.470 69.060 18.790 69.120 ;
        RECT 11.570 68.780 13.180 68.920 ;
        RECT 13.410 68.920 13.730 68.980 ;
        RECT 16.185 68.920 16.475 68.965 ;
        RECT 13.410 68.780 16.475 68.920 ;
        RECT 2.830 68.580 3.150 68.640 ;
        RECT 7.980 68.625 8.120 68.780 ;
        RECT 11.570 68.720 11.890 68.780 ;
        RECT 13.410 68.720 13.730 68.780 ;
        RECT 16.185 68.735 16.475 68.780 ;
        RECT 18.010 68.920 18.330 68.980 ;
        RECT 18.010 68.780 20.080 68.920 ;
        RECT 18.010 68.720 18.330 68.780 ;
        RECT 7.905 68.580 8.195 68.625 ;
        RECT 2.830 68.440 8.195 68.580 ;
        RECT 2.830 68.380 3.150 68.440 ;
        RECT 7.905 68.395 8.195 68.440 ;
        RECT 12.045 68.580 12.335 68.625 ;
        RECT 12.490 68.580 12.810 68.640 ;
        RECT 12.045 68.440 12.810 68.580 ;
        RECT 12.045 68.395 12.335 68.440 ;
        RECT 12.490 68.380 12.810 68.440 ;
        RECT 15.710 68.380 16.030 68.640 ;
        RECT 17.090 68.580 17.410 68.640 ;
        RECT 19.405 68.580 19.695 68.625 ;
        RECT 17.090 68.440 19.695 68.580 ;
        RECT 19.940 68.580 20.080 68.780 ;
        RECT 20.310 68.720 20.630 68.980 ;
        RECT 21.230 68.920 21.550 68.980 ;
        RECT 25.000 68.920 25.140 69.460 ;
        RECT 25.370 69.400 25.690 69.460 ;
        RECT 26.290 69.400 26.610 69.660 ;
        RECT 26.765 69.600 27.055 69.645 ;
        RECT 26.765 69.460 27.900 69.600 ;
        RECT 26.765 69.415 27.055 69.460 ;
        RECT 27.760 69.320 27.900 69.460 ;
        RECT 27.670 69.060 27.990 69.320 ;
        RECT 28.130 69.060 28.450 69.320 ;
        RECT 28.680 69.260 28.820 69.800 ;
        RECT 30.445 69.755 30.735 69.800 ;
        RECT 30.980 69.800 40.320 69.940 ;
        RECT 29.050 69.600 29.370 69.660 ;
        RECT 30.980 69.600 31.120 69.800 ;
        RECT 29.050 69.460 31.120 69.600 ;
        RECT 32.745 69.600 33.035 69.645 ;
        RECT 34.570 69.600 34.890 69.660 ;
        RECT 37.345 69.600 37.635 69.645 ;
        RECT 32.745 69.460 33.420 69.600 ;
        RECT 29.050 69.400 29.370 69.460 ;
        RECT 32.745 69.415 33.035 69.460 ;
        RECT 32.270 69.305 32.590 69.320 ;
        RECT 28.680 69.120 32.040 69.260 ;
        RECT 27.225 68.920 27.515 68.965 ;
        RECT 31.900 68.920 32.040 69.120 ;
        RECT 32.195 69.075 32.590 69.305 ;
        RECT 32.270 69.060 32.590 69.075 ;
        RECT 33.280 68.920 33.420 69.460 ;
        RECT 34.570 69.460 37.635 69.600 ;
        RECT 34.570 69.400 34.890 69.460 ;
        RECT 37.345 69.415 37.635 69.460 ;
        RECT 34.110 69.260 34.430 69.320 ;
        RECT 35.045 69.260 35.335 69.305 ;
        RECT 34.110 69.120 35.335 69.260 ;
        RECT 34.110 69.060 34.430 69.120 ;
        RECT 35.045 69.075 35.335 69.120 ;
        RECT 36.410 69.060 36.730 69.320 ;
        RECT 37.420 69.260 37.560 69.415 ;
        RECT 38.250 69.400 38.570 69.660 ;
        RECT 38.710 69.400 39.030 69.660 ;
        RECT 39.170 69.600 39.490 69.660 ;
        RECT 40.180 69.600 40.320 69.800 ;
        RECT 40.550 69.740 40.870 70.000 ;
        RECT 47.080 69.940 47.220 70.140 ;
        RECT 55.820 69.985 55.960 70.140 ;
        RECT 62.170 70.140 64.315 70.280 ;
        RECT 62.170 70.080 62.490 70.140 ;
        RECT 64.025 70.095 64.315 70.140 ;
        RECT 68.240 70.140 74.450 70.280 ;
        RECT 53.905 69.940 54.195 69.985 ;
        RECT 41.330 69.800 47.220 69.940 ;
        RECT 47.540 69.800 54.195 69.940 ;
        RECT 41.330 69.600 41.470 69.800 ;
        RECT 39.170 69.460 39.685 69.600 ;
        RECT 40.180 69.460 41.470 69.600 ;
        RECT 46.530 69.590 46.850 69.660 ;
        RECT 47.540 69.590 47.680 69.800 ;
        RECT 53.905 69.755 54.195 69.800 ;
        RECT 55.745 69.940 56.035 69.985 ;
        RECT 68.240 69.940 68.380 70.140 ;
        RECT 74.130 70.080 74.450 70.140 ;
        RECT 74.605 69.940 74.895 69.985 ;
        RECT 55.745 69.800 68.380 69.940 ;
        RECT 68.700 69.800 74.895 69.940 ;
        RECT 55.745 69.755 56.035 69.800 ;
        RECT 39.170 69.400 39.490 69.460 ;
        RECT 46.530 69.450 47.680 69.590 ;
        RECT 48.370 69.600 48.690 69.660 ;
        RECT 49.305 69.600 49.595 69.645 ;
        RECT 50.300 69.600 51.360 69.630 ;
        RECT 51.605 69.600 51.895 69.645 ;
        RECT 48.370 69.460 49.595 69.600 ;
        RECT 46.530 69.400 46.850 69.450 ;
        RECT 48.370 69.400 48.690 69.460 ;
        RECT 49.305 69.415 49.595 69.460 ;
        RECT 49.840 69.490 51.895 69.600 ;
        RECT 49.840 69.460 50.440 69.490 ;
        RECT 51.220 69.460 51.895 69.490 ;
        RECT 44.230 69.260 44.550 69.320 ;
        RECT 37.420 69.120 44.550 69.260 ;
        RECT 44.230 69.060 44.550 69.120 ;
        RECT 45.610 69.260 45.930 69.320 ;
        RECT 49.840 69.260 49.980 69.460 ;
        RECT 51.605 69.415 51.895 69.460 ;
        RECT 52.525 69.600 52.815 69.645 ;
        RECT 54.825 69.600 55.115 69.645 ;
        RECT 52.525 69.460 55.115 69.600 ;
        RECT 52.525 69.415 52.815 69.460 ;
        RECT 54.825 69.415 55.115 69.460 ;
        RECT 56.190 69.400 56.510 69.660 ;
        RECT 57.570 69.400 57.890 69.660 ;
        RECT 68.150 69.400 68.470 69.660 ;
        RECT 68.700 69.645 68.840 69.800 ;
        RECT 68.625 69.415 68.915 69.645 ;
        RECT 69.070 69.400 69.390 69.660 ;
        RECT 69.545 69.600 69.835 69.645 ;
        RECT 69.990 69.600 70.310 69.660 ;
        RECT 69.545 69.460 70.310 69.600 ;
        RECT 69.545 69.415 69.835 69.460 ;
        RECT 69.990 69.400 70.310 69.460 ;
        RECT 71.830 69.400 72.150 69.660 ;
        RECT 72.380 69.645 72.520 69.800 ;
        RECT 74.605 69.755 74.895 69.800 ;
        RECT 72.305 69.415 72.595 69.645 ;
        RECT 73.225 69.415 73.515 69.645 ;
        RECT 73.670 69.600 73.990 69.660 ;
        RECT 74.145 69.600 74.435 69.645 ;
        RECT 73.670 69.460 74.435 69.600 ;
        RECT 45.610 69.120 49.980 69.260 ;
        RECT 45.610 69.060 45.930 69.120 ;
        RECT 50.210 69.060 50.530 69.320 ;
        RECT 50.685 69.075 50.975 69.305 ;
        RECT 21.230 68.780 25.140 68.920 ;
        RECT 25.895 68.780 31.580 68.920 ;
        RECT 31.900 68.780 33.420 68.920 ;
        RECT 34.570 68.920 34.890 68.980 ;
        RECT 38.710 68.920 39.030 68.980 ;
        RECT 47.450 68.920 47.770 68.980 ;
        RECT 34.570 68.780 39.030 68.920 ;
        RECT 21.230 68.720 21.550 68.780 ;
        RECT 21.320 68.580 21.460 68.720 ;
        RECT 19.940 68.440 21.460 68.580 ;
        RECT 17.090 68.380 17.410 68.440 ;
        RECT 19.405 68.395 19.695 68.440 ;
        RECT 23.530 68.380 23.850 68.640 ;
        RECT 24.450 68.580 24.770 68.640 ;
        RECT 25.895 68.580 26.035 68.780 ;
        RECT 27.225 68.735 27.515 68.780 ;
        RECT 31.440 68.640 31.580 68.780 ;
        RECT 34.570 68.720 34.890 68.780 ;
        RECT 38.710 68.720 39.030 68.780 ;
        RECT 39.260 68.780 47.770 68.920 ;
        RECT 24.450 68.440 26.035 68.580 ;
        RECT 26.290 68.580 26.610 68.640 ;
        RECT 30.890 68.580 31.210 68.640 ;
        RECT 26.290 68.440 31.210 68.580 ;
        RECT 24.450 68.380 24.770 68.440 ;
        RECT 26.290 68.380 26.610 68.440 ;
        RECT 30.890 68.380 31.210 68.440 ;
        RECT 31.350 68.380 31.670 68.640 ;
        RECT 32.730 68.580 33.050 68.640 ;
        RECT 39.260 68.580 39.400 68.780 ;
        RECT 47.450 68.720 47.770 68.780 ;
        RECT 48.370 68.920 48.690 68.980 ;
        RECT 50.820 68.920 50.960 69.075 ;
        RECT 51.130 69.060 51.450 69.320 ;
        RECT 56.650 69.260 56.970 69.320 ;
        RECT 70.080 69.260 70.220 69.400 ;
        RECT 73.300 69.260 73.440 69.415 ;
        RECT 73.670 69.400 73.990 69.460 ;
        RECT 74.145 69.415 74.435 69.460 ;
        RECT 75.065 69.600 75.355 69.645 ;
        RECT 75.510 69.600 75.830 69.660 ;
        RECT 75.065 69.460 75.830 69.600 ;
        RECT 75.065 69.415 75.355 69.460 ;
        RECT 75.510 69.400 75.830 69.460 ;
        RECT 56.650 69.120 69.760 69.260 ;
        RECT 70.080 69.120 73.440 69.260 ;
        RECT 56.650 69.060 56.970 69.120 ;
        RECT 48.370 68.780 50.960 68.920 ;
        RECT 59.870 68.920 60.190 68.980 ;
        RECT 67.245 68.920 67.535 68.965 ;
        RECT 59.870 68.780 67.535 68.920 ;
        RECT 69.620 68.920 69.760 69.120 ;
        RECT 72.765 68.920 73.055 68.965 ;
        RECT 69.620 68.780 73.055 68.920 ;
        RECT 48.370 68.720 48.690 68.780 ;
        RECT 59.870 68.720 60.190 68.780 ;
        RECT 67.245 68.735 67.535 68.780 ;
        RECT 72.765 68.735 73.055 68.780 ;
        RECT 32.730 68.440 39.400 68.580 ;
        RECT 41.470 68.580 41.790 68.640 ;
        RECT 63.090 68.580 63.410 68.640 ;
        RECT 41.470 68.440 63.410 68.580 ;
        RECT 32.730 68.380 33.050 68.440 ;
        RECT 41.470 68.380 41.790 68.440 ;
        RECT 63.090 68.380 63.410 68.440 ;
        RECT 70.910 68.380 71.230 68.640 ;
        RECT 5.520 67.760 76.820 68.240 ;
        RECT 5.590 67.560 5.910 67.620 ;
        RECT 10.205 67.560 10.495 67.605 ;
        RECT 5.590 67.420 10.495 67.560 ;
        RECT 5.590 67.360 5.910 67.420 ;
        RECT 10.205 67.375 10.495 67.420 ;
        RECT 10.650 67.560 10.970 67.620 ;
        RECT 17.090 67.560 17.410 67.620 ;
        RECT 10.650 67.420 17.410 67.560 ;
        RECT 10.650 67.360 10.970 67.420 ;
        RECT 17.090 67.360 17.410 67.420 ;
        RECT 22.150 67.560 22.470 67.620 ;
        RECT 29.985 67.560 30.275 67.605 ;
        RECT 34.570 67.560 34.890 67.620 ;
        RECT 22.150 67.420 29.740 67.560 ;
        RECT 22.150 67.360 22.470 67.420 ;
        RECT 8.825 67.220 9.115 67.265 ;
        RECT 9.270 67.220 9.590 67.280 ;
        RECT 8.825 67.080 9.590 67.220 ;
        RECT 8.825 67.035 9.115 67.080 ;
        RECT 9.270 67.020 9.590 67.080 ;
        RECT 11.570 67.220 11.890 67.280 ;
        RECT 18.010 67.220 18.330 67.280 ;
        RECT 11.570 67.080 18.330 67.220 ;
        RECT 11.570 67.020 11.890 67.080 ;
        RECT 9.360 66.880 9.500 67.020 ;
        RECT 10.650 66.880 10.970 66.940 ;
        RECT 9.360 66.740 10.970 66.880 ;
        RECT 10.650 66.680 10.970 66.740 ;
        RECT 7.430 66.540 7.750 66.600 ;
        RECT 7.905 66.540 8.195 66.585 ;
        RECT 7.430 66.400 8.195 66.540 ;
        RECT 7.430 66.340 7.750 66.400 ;
        RECT 7.905 66.355 8.195 66.400 ;
        RECT 11.110 66.340 11.430 66.600 ;
        RECT 12.490 66.340 12.810 66.600 ;
        RECT 13.040 66.585 13.180 67.080 ;
        RECT 18.010 67.020 18.330 67.080 ;
        RECT 18.930 67.020 19.250 67.280 ;
        RECT 23.530 67.020 23.850 67.280 ;
        RECT 26.750 67.220 27.070 67.280 ;
        RECT 29.050 67.220 29.370 67.280 ;
        RECT 24.080 67.080 29.370 67.220 ;
        RECT 29.600 67.220 29.740 67.420 ;
        RECT 29.985 67.420 34.890 67.560 ;
        RECT 29.985 67.375 30.275 67.420 ;
        RECT 34.570 67.360 34.890 67.420 ;
        RECT 37.345 67.560 37.635 67.605 ;
        RECT 38.250 67.560 38.570 67.620 ;
        RECT 37.345 67.420 38.570 67.560 ;
        RECT 37.345 67.375 37.635 67.420 ;
        RECT 38.250 67.360 38.570 67.420 ;
        RECT 40.090 67.360 40.410 67.620 ;
        RECT 41.470 67.360 41.790 67.620 ;
        RECT 45.150 67.560 45.470 67.620 ;
        RECT 47.005 67.560 47.295 67.605 ;
        RECT 57.570 67.560 57.890 67.620 ;
        RECT 45.150 67.420 57.890 67.560 ;
        RECT 45.150 67.360 45.470 67.420 ;
        RECT 47.005 67.375 47.295 67.420 ;
        RECT 57.570 67.360 57.890 67.420 ;
        RECT 67.690 67.560 68.010 67.620 ;
        RECT 73.670 67.560 73.990 67.620 ;
        RECT 67.690 67.420 73.990 67.560 ;
        RECT 67.690 67.360 68.010 67.420 ;
        RECT 73.670 67.360 73.990 67.420 ;
        RECT 33.190 67.220 33.510 67.280 ;
        RECT 29.600 67.080 33.510 67.220 ;
        RECT 13.410 66.880 13.730 66.940 ;
        RECT 20.770 66.880 21.090 66.940 ;
        RECT 23.620 66.880 23.760 67.020 ;
        RECT 24.080 66.925 24.220 67.080 ;
        RECT 26.750 67.020 27.070 67.080 ;
        RECT 29.050 67.020 29.370 67.080 ;
        RECT 33.190 67.020 33.510 67.080 ;
        RECT 33.650 67.220 33.970 67.280 ;
        RECT 33.650 67.080 39.860 67.220 ;
        RECT 33.650 67.020 33.970 67.080 ;
        RECT 13.410 66.740 14.230 66.880 ;
        RECT 13.410 66.680 13.730 66.740 ;
        RECT 14.090 66.585 14.230 66.740 ;
        RECT 17.640 66.740 23.760 66.880 ;
        RECT 12.965 66.355 13.255 66.585 ;
        RECT 14.015 66.355 14.305 66.585 ;
        RECT 14.790 66.340 15.110 66.600 ;
        RECT 15.710 66.540 16.030 66.600 ;
        RECT 17.640 66.585 17.780 66.740 ;
        RECT 20.770 66.680 21.090 66.740 ;
        RECT 24.005 66.695 24.295 66.925 ;
        RECT 24.465 66.880 24.755 66.925 ;
        RECT 28.590 66.880 28.910 66.940 ;
        RECT 24.465 66.740 28.910 66.880 ;
        RECT 24.465 66.695 24.755 66.740 ;
        RECT 28.590 66.680 28.910 66.740 ;
        RECT 29.970 66.880 30.290 66.940 ;
        RECT 39.720 66.925 39.860 67.080 ;
        RECT 38.725 66.880 39.015 66.925 ;
        RECT 29.970 66.740 39.015 66.880 ;
        RECT 29.970 66.680 30.290 66.740 ;
        RECT 38.725 66.695 39.015 66.740 ;
        RECT 39.645 66.695 39.935 66.925 ;
        RECT 40.180 66.600 40.320 67.360 ;
        RECT 51.130 67.220 51.450 67.280 ;
        RECT 53.890 67.220 54.210 67.280 ;
        RECT 51.130 67.080 54.210 67.220 ;
        RECT 51.130 67.020 51.450 67.080 ;
        RECT 53.890 67.020 54.210 67.080 ;
        RECT 56.190 67.220 56.510 67.280 ;
        RECT 57.125 67.220 57.415 67.265 ;
        RECT 59.410 67.220 59.730 67.280 ;
        RECT 75.065 67.220 75.355 67.265 ;
        RECT 56.190 67.080 59.730 67.220 ;
        RECT 56.190 67.020 56.510 67.080 ;
        RECT 57.125 67.035 57.415 67.080 ;
        RECT 59.410 67.020 59.730 67.080 ;
        RECT 59.960 67.080 75.355 67.220 ;
        RECT 53.430 66.880 53.750 66.940 ;
        RECT 59.960 66.880 60.100 67.080 ;
        RECT 75.065 67.035 75.355 67.080 ;
        RECT 40.640 66.740 53.750 66.880 ;
        RECT 40.640 66.600 40.780 66.740 ;
        RECT 53.430 66.680 53.750 66.740 ;
        RECT 59.500 66.740 60.100 66.880 ;
        RECT 60.790 66.880 61.110 66.940 ;
        RECT 70.925 66.880 71.215 66.925 ;
        RECT 60.790 66.740 71.215 66.880 ;
        RECT 16.185 66.540 16.475 66.585 ;
        RECT 15.710 66.400 16.475 66.540 ;
        RECT 15.710 66.340 16.030 66.400 ;
        RECT 16.185 66.355 16.475 66.400 ;
        RECT 17.565 66.355 17.855 66.585 ;
        RECT 20.310 66.340 20.630 66.600 ;
        RECT 22.150 66.340 22.470 66.600 ;
        RECT 22.610 66.340 22.930 66.600 ;
        RECT 23.545 66.345 23.835 66.575 ;
        RECT 25.385 66.355 25.675 66.585 ;
        RECT 25.830 66.540 26.150 66.600 ;
        RECT 26.305 66.540 26.595 66.585 ;
        RECT 25.830 66.400 26.595 66.540 ;
        RECT 12.030 66.200 12.350 66.260 ;
        RECT 13.425 66.200 13.715 66.245 ;
        RECT 17.105 66.200 17.395 66.245 ;
        RECT 12.030 66.060 17.395 66.200 ;
        RECT 12.030 66.000 12.350 66.060 ;
        RECT 13.425 66.015 13.715 66.060 ;
        RECT 17.105 66.015 17.395 66.060 ;
        RECT 18.945 66.200 19.235 66.245 ;
        RECT 23.070 66.200 23.390 66.260 ;
        RECT 23.620 66.200 23.760 66.345 ;
        RECT 18.945 66.060 21.880 66.200 ;
        RECT 18.945 66.015 19.235 66.060 ;
        RECT 11.570 65.660 11.890 65.920 ;
        RECT 15.250 65.660 15.570 65.920 ;
        RECT 17.180 65.860 17.320 66.015 ;
        RECT 20.400 65.920 20.540 66.060 ;
        RECT 19.850 65.860 20.170 65.920 ;
        RECT 17.180 65.720 20.170 65.860 ;
        RECT 19.850 65.660 20.170 65.720 ;
        RECT 20.310 65.660 20.630 65.920 ;
        RECT 21.230 65.660 21.550 65.920 ;
        RECT 21.740 65.860 21.880 66.060 ;
        RECT 23.070 66.060 23.760 66.200 ;
        RECT 23.070 66.000 23.390 66.060 ;
        RECT 24.910 65.860 25.230 65.920 ;
        RECT 21.740 65.720 25.230 65.860 ;
        RECT 25.460 65.860 25.600 66.355 ;
        RECT 25.830 66.340 26.150 66.400 ;
        RECT 26.305 66.355 26.595 66.400 ;
        RECT 31.350 66.540 31.670 66.600 ;
        RECT 31.350 66.400 38.075 66.540 ;
        RECT 31.350 66.340 31.670 66.400 ;
        RECT 28.130 66.200 28.450 66.260 ;
        RECT 30.890 66.200 31.210 66.260 ;
        RECT 28.130 66.060 31.210 66.200 ;
        RECT 28.130 66.000 28.450 66.060 ;
        RECT 30.890 66.000 31.210 66.060 ;
        RECT 36.410 66.000 36.730 66.260 ;
        RECT 37.935 66.200 38.075 66.400 ;
        RECT 38.250 66.340 38.570 66.600 ;
        RECT 39.185 66.355 39.475 66.585 ;
        RECT 39.260 66.200 39.400 66.355 ;
        RECT 40.090 66.340 40.410 66.600 ;
        RECT 40.550 66.340 40.870 66.600 ;
        RECT 41.010 66.340 41.330 66.600 ;
        RECT 41.470 66.540 41.790 66.600 ;
        RECT 42.405 66.540 42.695 66.585 ;
        RECT 41.470 66.400 42.695 66.540 ;
        RECT 41.470 66.340 41.790 66.400 ;
        RECT 42.405 66.355 42.695 66.400 ;
        RECT 42.865 66.540 43.155 66.585 ;
        RECT 43.310 66.540 43.630 66.600 ;
        RECT 42.865 66.400 43.630 66.540 ;
        RECT 42.865 66.355 43.155 66.400 ;
        RECT 43.310 66.340 43.630 66.400 ;
        RECT 53.890 66.340 54.210 66.600 ;
        RECT 54.350 66.585 54.670 66.600 ;
        RECT 54.350 66.355 54.885 66.585 ;
        RECT 54.350 66.340 54.670 66.355 ;
        RECT 55.730 66.340 56.050 66.600 ;
        RECT 56.190 66.340 56.510 66.600 ;
        RECT 57.585 66.540 57.875 66.585 ;
        RECT 58.950 66.540 59.270 66.600 ;
        RECT 57.585 66.400 59.270 66.540 ;
        RECT 57.585 66.355 57.875 66.400 ;
        RECT 58.950 66.340 59.270 66.400 ;
        RECT 43.785 66.200 44.075 66.245 ;
        RECT 37.935 66.060 44.075 66.200 ;
        RECT 43.785 66.015 44.075 66.060 ;
        RECT 44.230 66.200 44.550 66.260 ;
        RECT 52.510 66.200 52.830 66.260 ;
        RECT 44.230 66.060 52.830 66.200 ;
        RECT 25.830 65.860 26.150 65.920 ;
        RECT 25.460 65.720 26.150 65.860 ;
        RECT 24.910 65.660 25.230 65.720 ;
        RECT 25.830 65.660 26.150 65.720 ;
        RECT 34.570 65.860 34.890 65.920 ;
        RECT 38.250 65.860 38.570 65.920 ;
        RECT 34.570 65.720 38.570 65.860 ;
        RECT 43.860 65.860 44.000 66.015 ;
        RECT 44.230 66.000 44.550 66.060 ;
        RECT 52.510 66.000 52.830 66.060 ;
        RECT 53.430 66.000 53.750 66.260 ;
        RECT 55.285 66.015 55.575 66.245 ;
        RECT 57.110 66.200 57.430 66.260 ;
        RECT 58.490 66.245 58.810 66.260 ;
        RECT 59.500 66.245 59.640 66.740 ;
        RECT 60.790 66.680 61.110 66.740 ;
        RECT 70.925 66.695 71.215 66.740 ;
        RECT 71.830 66.340 72.150 66.600 ;
        RECT 72.750 66.340 73.070 66.600 ;
        RECT 73.225 66.355 73.515 66.585 ;
        RECT 73.685 66.355 73.975 66.585 ;
        RECT 58.305 66.200 58.810 66.245 ;
        RECT 57.110 66.060 58.810 66.200 ;
        RECT 48.370 65.860 48.690 65.920 ;
        RECT 43.860 65.720 48.690 65.860 ;
        RECT 34.570 65.660 34.890 65.720 ;
        RECT 38.250 65.660 38.570 65.720 ;
        RECT 48.370 65.660 48.690 65.720 ;
        RECT 51.590 65.860 51.910 65.920 ;
        RECT 55.360 65.860 55.500 66.015 ;
        RECT 57.110 66.000 57.430 66.060 ;
        RECT 58.305 66.015 58.810 66.060 ;
        RECT 59.425 66.015 59.715 66.245 ;
        RECT 60.345 66.200 60.635 66.245 ;
        RECT 61.710 66.200 62.030 66.260 ;
        RECT 66.310 66.200 66.630 66.260 ;
        RECT 69.545 66.200 69.835 66.245 ;
        RECT 60.345 66.060 62.030 66.200 ;
        RECT 60.345 66.015 60.635 66.060 ;
        RECT 58.490 66.000 58.810 66.015 ;
        RECT 61.710 66.000 62.030 66.060 ;
        RECT 62.720 66.060 66.080 66.200 ;
        RECT 51.590 65.720 55.500 65.860 ;
        RECT 51.590 65.660 51.910 65.720 ;
        RECT 58.950 65.660 59.270 65.920 ;
        RECT 59.870 65.860 60.190 65.920 ;
        RECT 62.720 65.860 62.860 66.060 ;
        RECT 59.870 65.720 62.860 65.860 ;
        RECT 63.105 65.860 63.395 65.905 ;
        RECT 64.010 65.860 64.330 65.920 ;
        RECT 63.105 65.720 64.330 65.860 ;
        RECT 65.940 65.860 66.080 66.060 ;
        RECT 66.310 66.060 69.835 66.200 ;
        RECT 66.310 66.000 66.630 66.060 ;
        RECT 69.545 66.015 69.835 66.060 ;
        RECT 70.450 66.200 70.770 66.260 ;
        RECT 73.300 66.200 73.440 66.355 ;
        RECT 70.450 66.060 73.440 66.200 ;
        RECT 70.450 66.000 70.770 66.060 ;
        RECT 73.760 65.860 73.900 66.355 ;
        RECT 74.130 66.340 74.450 66.600 ;
        RECT 74.590 66.540 74.910 66.600 ;
        RECT 75.065 66.540 75.355 66.585 ;
        RECT 74.590 66.400 75.355 66.540 ;
        RECT 74.590 66.340 74.910 66.400 ;
        RECT 75.065 66.355 75.355 66.400 ;
        RECT 65.940 65.720 73.900 65.860 ;
        RECT 59.870 65.660 60.190 65.720 ;
        RECT 63.105 65.675 63.395 65.720 ;
        RECT 64.010 65.660 64.330 65.720 ;
        RECT 5.520 65.040 76.820 65.520 ;
        RECT 13.885 64.840 14.175 64.885 ;
        RECT 14.790 64.840 15.110 64.900 ;
        RECT 13.885 64.700 15.110 64.840 ;
        RECT 13.885 64.655 14.175 64.700 ;
        RECT 14.790 64.640 15.110 64.700 ;
        RECT 15.725 64.840 16.015 64.885 ;
        RECT 17.550 64.840 17.870 64.900 ;
        RECT 15.725 64.700 17.870 64.840 ;
        RECT 15.725 64.655 16.015 64.700 ;
        RECT 17.550 64.640 17.870 64.700 ;
        RECT 18.485 64.840 18.775 64.885 ;
        RECT 21.245 64.840 21.535 64.885 ;
        RECT 22.150 64.840 22.470 64.900 ;
        RECT 25.370 64.840 25.690 64.900 ;
        RECT 18.485 64.700 21.000 64.840 ;
        RECT 18.485 64.655 18.775 64.700 ;
        RECT 4.670 64.500 4.990 64.560 ;
        RECT 11.125 64.500 11.415 64.545 ;
        RECT 13.410 64.500 13.730 64.560 ;
        RECT 4.670 64.360 9.500 64.500 ;
        RECT 4.670 64.300 4.990 64.360 ;
        RECT 8.350 63.960 8.670 64.220 ;
        RECT 9.360 64.205 9.500 64.360 ;
        RECT 11.125 64.360 13.730 64.500 ;
        RECT 11.125 64.315 11.415 64.360 ;
        RECT 13.410 64.300 13.730 64.360 ;
        RECT 19.405 64.500 19.695 64.545 ;
        RECT 19.850 64.500 20.170 64.560 ;
        RECT 19.405 64.360 20.170 64.500 ;
        RECT 19.405 64.315 19.695 64.360 ;
        RECT 19.850 64.300 20.170 64.360 ;
        RECT 20.310 64.300 20.630 64.560 ;
        RECT 20.860 64.500 21.000 64.700 ;
        RECT 21.245 64.700 25.690 64.840 ;
        RECT 21.245 64.655 21.535 64.700 ;
        RECT 22.150 64.640 22.470 64.700 ;
        RECT 25.370 64.640 25.690 64.700 ;
        RECT 25.845 64.840 26.135 64.885 ;
        RECT 30.430 64.840 30.750 64.900 ;
        RECT 34.110 64.840 34.430 64.900 ;
        RECT 35.505 64.840 35.795 64.885 ;
        RECT 25.845 64.700 30.750 64.840 ;
        RECT 25.845 64.655 26.135 64.700 ;
        RECT 30.430 64.640 30.750 64.700 ;
        RECT 33.280 64.700 35.795 64.840 ;
        RECT 33.280 64.545 33.420 64.700 ;
        RECT 34.110 64.640 34.430 64.700 ;
        RECT 35.505 64.655 35.795 64.700 ;
        RECT 36.410 64.840 36.730 64.900 ;
        RECT 40.550 64.840 40.870 64.900 ;
        RECT 36.410 64.700 40.870 64.840 ;
        RECT 36.410 64.640 36.730 64.700 ;
        RECT 40.550 64.640 40.870 64.700 ;
        RECT 41.025 64.840 41.315 64.885 ;
        RECT 41.930 64.840 42.250 64.900 ;
        RECT 62.170 64.840 62.490 64.900 ;
        RECT 41.025 64.700 42.250 64.840 ;
        RECT 41.025 64.655 41.315 64.700 ;
        RECT 41.930 64.640 42.250 64.700 ;
        RECT 59.500 64.700 62.490 64.840 ;
        RECT 20.860 64.360 27.900 64.500 ;
        RECT 9.285 63.975 9.575 64.205 ;
        RECT 11.585 63.975 11.875 64.205 ;
        RECT 12.045 64.160 12.335 64.205 ;
        RECT 12.490 64.160 12.810 64.220 ;
        RECT 12.045 64.020 12.810 64.160 ;
        RECT 12.045 63.975 12.335 64.020 ;
        RECT 5.130 63.820 5.450 63.880 ;
        RECT 11.660 63.820 11.800 63.975 ;
        RECT 12.490 63.960 12.810 64.020 ;
        RECT 12.965 63.975 13.255 64.205 ;
        RECT 16.185 64.160 16.475 64.205 ;
        RECT 16.630 64.160 16.950 64.220 ;
        RECT 16.185 64.020 16.950 64.160 ;
        RECT 16.185 63.975 16.475 64.020 ;
        RECT 13.040 63.820 13.180 63.975 ;
        RECT 16.630 63.960 16.950 64.020 ;
        RECT 17.105 64.160 17.395 64.205 ;
        RECT 17.565 64.160 17.855 64.205 ;
        RECT 18.470 64.160 18.790 64.220 ;
        RECT 17.105 64.020 18.790 64.160 ;
        RECT 17.105 63.975 17.395 64.020 ;
        RECT 17.565 63.975 17.855 64.020 ;
        RECT 18.470 63.960 18.790 64.020 ;
        RECT 18.945 64.160 19.235 64.205 ;
        RECT 20.770 64.160 21.090 64.220 ;
        RECT 18.945 64.020 21.090 64.160 ;
        RECT 18.945 63.975 19.235 64.020 ;
        RECT 20.770 63.960 21.090 64.020 ;
        RECT 21.665 64.160 21.955 64.205 ;
        RECT 22.150 64.160 22.470 64.220 ;
        RECT 21.665 64.020 22.470 64.160 ;
        RECT 21.665 63.975 21.955 64.020 ;
        RECT 22.150 63.960 22.470 64.020 ;
        RECT 23.530 64.160 23.850 64.220 ;
        RECT 24.005 64.160 24.295 64.205 ;
        RECT 23.530 64.020 24.295 64.160 ;
        RECT 23.530 63.960 23.850 64.020 ;
        RECT 24.005 63.975 24.295 64.020 ;
        RECT 24.450 63.960 24.770 64.220 ;
        RECT 27.760 64.205 27.900 64.360 ;
        RECT 33.205 64.315 33.495 64.545 ;
        RECT 33.665 64.500 33.955 64.545 ;
        RECT 34.570 64.500 34.890 64.560 ;
        RECT 33.665 64.360 34.890 64.500 ;
        RECT 33.665 64.315 33.955 64.360 ;
        RECT 34.570 64.300 34.890 64.360 ;
        RECT 36.870 64.300 37.190 64.560 ;
        RECT 37.330 64.500 37.650 64.560 ;
        RECT 41.470 64.500 41.790 64.560 ;
        RECT 37.330 64.360 41.790 64.500 ;
        RECT 37.330 64.300 37.650 64.360 ;
        RECT 41.470 64.300 41.790 64.360 ;
        RECT 44.230 64.500 44.550 64.560 ;
        RECT 51.590 64.500 51.910 64.560 ;
        RECT 44.230 64.360 51.910 64.500 ;
        RECT 44.230 64.300 44.550 64.360 ;
        RECT 51.590 64.300 51.910 64.360 ;
        RECT 53.890 64.500 54.210 64.560 ;
        RECT 57.110 64.500 57.430 64.560 ;
        RECT 53.890 64.360 57.430 64.500 ;
        RECT 53.890 64.300 54.210 64.360 ;
        RECT 57.110 64.300 57.430 64.360 ;
        RECT 26.765 63.975 27.055 64.205 ;
        RECT 27.685 63.975 27.975 64.205 ;
        RECT 5.130 63.680 13.180 63.820 ;
        RECT 13.410 63.820 13.730 63.880 ;
        RECT 26.840 63.820 26.980 63.975 ;
        RECT 13.410 63.680 26.980 63.820 ;
        RECT 27.760 63.820 27.900 63.975 ;
        RECT 28.130 63.960 28.450 64.220 ;
        RECT 28.590 64.160 28.910 64.220 ;
        RECT 30.430 64.160 30.750 64.220 ;
        RECT 28.590 64.020 30.750 64.160 ;
        RECT 28.590 63.960 28.910 64.020 ;
        RECT 30.430 63.960 30.750 64.020 ;
        RECT 32.270 63.960 32.590 64.220 ;
        RECT 32.730 64.160 33.050 64.220 ;
        RECT 34.125 64.160 34.415 64.205 ;
        RECT 32.730 64.020 34.415 64.160 ;
        RECT 32.730 63.960 33.050 64.020 ;
        RECT 34.125 63.975 34.415 64.020 ;
        RECT 36.425 64.160 36.715 64.205 ;
        RECT 36.425 64.020 37.560 64.160 ;
        RECT 36.425 63.975 36.715 64.020 ;
        RECT 33.190 63.820 33.510 63.880 ;
        RECT 27.760 63.680 33.510 63.820 ;
        RECT 5.130 63.620 5.450 63.680 ;
        RECT 13.410 63.620 13.730 63.680 ;
        RECT 33.190 63.620 33.510 63.680 ;
        RECT 18.930 63.480 19.250 63.540 ;
        RECT 19.850 63.480 20.170 63.540 ;
        RECT 18.930 63.340 20.170 63.480 ;
        RECT 18.930 63.280 19.250 63.340 ;
        RECT 19.850 63.280 20.170 63.340 ;
        RECT 23.085 63.480 23.375 63.525 ;
        RECT 23.530 63.480 23.850 63.540 ;
        RECT 23.085 63.340 23.850 63.480 ;
        RECT 23.085 63.295 23.375 63.340 ;
        RECT 23.530 63.280 23.850 63.340 ;
        RECT 25.385 63.480 25.675 63.525 ;
        RECT 29.510 63.480 29.830 63.540 ;
        RECT 25.385 63.340 29.830 63.480 ;
        RECT 25.385 63.295 25.675 63.340 ;
        RECT 29.510 63.280 29.830 63.340 ;
        RECT 29.970 63.280 30.290 63.540 ;
        RECT 30.905 63.480 31.195 63.525 ;
        RECT 37.420 63.480 37.560 64.020 ;
        RECT 38.265 63.975 38.555 64.205 ;
        RECT 41.930 64.160 42.250 64.220 ;
        RECT 43.770 64.160 44.090 64.220 ;
        RECT 41.930 64.020 44.090 64.160 ;
        RECT 38.365 63.540 38.505 63.975 ;
        RECT 41.930 63.960 42.250 64.020 ;
        RECT 43.770 63.960 44.090 64.020 ;
        RECT 47.450 63.960 47.770 64.220 ;
        RECT 48.370 64.160 48.690 64.220 ;
        RECT 52.510 64.160 52.830 64.220 ;
        RECT 55.730 64.160 56.050 64.220 ;
        RECT 48.370 64.020 56.050 64.160 ;
        RECT 48.370 63.960 48.690 64.020 ;
        RECT 52.510 63.960 52.830 64.020 ;
        RECT 55.730 63.960 56.050 64.020 ;
        RECT 56.650 63.960 56.970 64.220 ;
        RECT 58.950 63.960 59.270 64.220 ;
        RECT 59.500 64.205 59.640 64.700 ;
        RECT 62.170 64.640 62.490 64.700 ;
        RECT 63.090 64.840 63.410 64.900 ;
        RECT 69.530 64.840 69.850 64.900 ;
        RECT 63.090 64.700 69.850 64.840 ;
        RECT 63.090 64.640 63.410 64.700 ;
        RECT 69.530 64.640 69.850 64.700 ;
        RECT 70.910 64.500 71.230 64.560 ;
        RECT 60.420 64.360 71.230 64.500 ;
        RECT 60.420 64.205 60.560 64.360 ;
        RECT 70.910 64.300 71.230 64.360 ;
        RECT 59.425 63.975 59.715 64.205 ;
        RECT 60.345 63.975 60.635 64.205 ;
        RECT 60.805 63.975 61.095 64.205 ;
        RECT 47.910 63.820 48.230 63.880 ;
        RECT 60.880 63.820 61.020 63.975 ;
        RECT 63.090 63.960 63.410 64.220 ;
        RECT 64.010 63.960 64.330 64.220 ;
        RECT 64.930 63.960 65.250 64.220 ;
        RECT 66.325 64.160 66.615 64.205 ;
        RECT 66.770 64.160 67.090 64.220 ;
        RECT 66.325 64.020 67.090 64.160 ;
        RECT 66.325 63.975 66.615 64.020 ;
        RECT 66.770 63.960 67.090 64.020 ;
        RECT 47.910 63.680 61.020 63.820 ;
        RECT 47.910 63.620 48.230 63.680 ;
        RECT 62.630 63.620 62.950 63.880 ;
        RECT 63.565 63.820 63.855 63.865 ;
        RECT 74.590 63.820 74.910 63.880 ;
        RECT 63.565 63.680 74.910 63.820 ;
        RECT 63.565 63.635 63.855 63.680 ;
        RECT 74.590 63.620 74.910 63.680 ;
        RECT 30.905 63.340 37.560 63.480 ;
        RECT 30.905 63.295 31.195 63.340 ;
        RECT 3.750 63.140 4.070 63.200 ;
        RECT 7.445 63.140 7.735 63.185 ;
        RECT 3.750 63.000 7.735 63.140 ;
        RECT 3.750 62.940 4.070 63.000 ;
        RECT 7.445 62.955 7.735 63.000 ;
        RECT 10.190 62.940 10.510 63.200 ;
        RECT 20.310 62.940 20.630 63.200 ;
        RECT 22.625 63.140 22.915 63.185 ;
        RECT 29.050 63.140 29.370 63.200 ;
        RECT 22.625 63.000 29.370 63.140 ;
        RECT 22.625 62.955 22.915 63.000 ;
        RECT 29.050 62.940 29.370 63.000 ;
        RECT 32.730 63.140 33.050 63.200 ;
        RECT 33.650 63.140 33.970 63.200 ;
        RECT 32.730 63.000 33.970 63.140 ;
        RECT 32.730 62.940 33.050 63.000 ;
        RECT 33.650 62.940 33.970 63.000 ;
        RECT 35.045 63.140 35.335 63.185 ;
        RECT 36.410 63.140 36.730 63.200 ;
        RECT 35.045 63.000 36.730 63.140 ;
        RECT 37.420 63.140 37.560 63.340 ;
        RECT 38.250 63.480 38.570 63.540 ;
        RECT 56.190 63.480 56.510 63.540 ;
        RECT 38.250 63.340 56.510 63.480 ;
        RECT 38.250 63.280 38.570 63.340 ;
        RECT 56.190 63.280 56.510 63.340 ;
        RECT 64.930 63.480 65.250 63.540 ;
        RECT 70.450 63.480 70.770 63.540 ;
        RECT 64.930 63.340 70.770 63.480 ;
        RECT 64.930 63.280 65.250 63.340 ;
        RECT 70.450 63.280 70.770 63.340 ;
        RECT 49.750 63.140 50.070 63.200 ;
        RECT 37.420 63.000 50.070 63.140 ;
        RECT 35.045 62.955 35.335 63.000 ;
        RECT 36.410 62.940 36.730 63.000 ;
        RECT 49.750 62.940 50.070 63.000 ;
        RECT 50.225 63.140 50.515 63.185 ;
        RECT 54.810 63.140 55.130 63.200 ;
        RECT 50.225 63.000 55.130 63.140 ;
        RECT 50.225 62.955 50.515 63.000 ;
        RECT 54.810 62.940 55.130 63.000 ;
        RECT 58.030 62.940 58.350 63.200 ;
        RECT 61.725 63.140 62.015 63.185 ;
        RECT 63.090 63.140 63.410 63.200 ;
        RECT 61.725 63.000 63.410 63.140 ;
        RECT 61.725 62.955 62.015 63.000 ;
        RECT 63.090 62.940 63.410 63.000 ;
        RECT 66.770 63.140 67.090 63.200 ;
        RECT 71.830 63.140 72.150 63.200 ;
        RECT 66.770 63.000 72.150 63.140 ;
        RECT 66.770 62.940 67.090 63.000 ;
        RECT 71.830 62.940 72.150 63.000 ;
        RECT 73.670 62.940 73.990 63.200 ;
        RECT 5.520 62.320 76.820 62.800 ;
        RECT 8.350 62.120 8.670 62.180 ;
        RECT 9.285 62.120 9.575 62.165 ;
        RECT 8.350 61.980 9.575 62.120 ;
        RECT 8.350 61.920 8.670 61.980 ;
        RECT 9.285 61.935 9.575 61.980 ;
        RECT 10.665 62.120 10.955 62.165 ;
        RECT 11.110 62.120 11.430 62.180 ;
        RECT 10.665 61.980 11.430 62.120 ;
        RECT 10.665 61.935 10.955 61.980 ;
        RECT 11.110 61.920 11.430 61.980 ;
        RECT 18.470 62.120 18.790 62.180 ;
        RECT 25.830 62.120 26.150 62.180 ;
        RECT 26.305 62.120 26.595 62.165 ;
        RECT 29.065 62.120 29.355 62.165 ;
        RECT 31.810 62.120 32.130 62.180 ;
        RECT 18.470 61.980 26.595 62.120 ;
        RECT 18.470 61.920 18.790 61.980 ;
        RECT 25.830 61.920 26.150 61.980 ;
        RECT 26.305 61.935 26.595 61.980 ;
        RECT 26.840 61.980 28.820 62.120 ;
        RECT 8.810 61.780 9.130 61.840 ;
        RECT 12.045 61.780 12.335 61.825 ;
        RECT 8.810 61.640 12.335 61.780 ;
        RECT 8.810 61.580 9.130 61.640 ;
        RECT 12.045 61.595 12.335 61.640 ;
        RECT 15.265 61.780 15.555 61.825 ;
        RECT 15.710 61.780 16.030 61.840 ;
        RECT 15.265 61.640 16.030 61.780 ;
        RECT 15.265 61.595 15.555 61.640 ;
        RECT 15.710 61.580 16.030 61.640 ;
        RECT 18.930 61.780 19.250 61.840 ;
        RECT 19.865 61.780 20.155 61.825 ;
        RECT 26.840 61.780 26.980 61.980 ;
        RECT 28.130 61.780 28.450 61.840 ;
        RECT 18.930 61.640 20.155 61.780 ;
        RECT 18.930 61.580 19.250 61.640 ;
        RECT 19.865 61.595 20.155 61.640 ;
        RECT 26.380 61.640 26.980 61.780 ;
        RECT 27.300 61.640 28.450 61.780 ;
        RECT 28.680 61.780 28.820 61.980 ;
        RECT 29.065 61.980 32.130 62.120 ;
        RECT 29.065 61.935 29.355 61.980 ;
        RECT 31.810 61.920 32.130 61.980 ;
        RECT 32.285 62.120 32.575 62.165 ;
        RECT 35.950 62.120 36.270 62.180 ;
        RECT 32.285 61.980 36.270 62.120 ;
        RECT 32.285 61.935 32.575 61.980 ;
        RECT 35.950 61.920 36.270 61.980 ;
        RECT 47.465 62.120 47.755 62.165 ;
        RECT 47.910 62.120 48.230 62.180 ;
        RECT 72.765 62.120 73.055 62.165 ;
        RECT 47.465 61.980 48.230 62.120 ;
        RECT 47.465 61.935 47.755 61.980 ;
        RECT 47.910 61.920 48.230 61.980 ;
        RECT 48.460 61.980 73.055 62.120 ;
        RECT 33.650 61.780 33.970 61.840 ;
        RECT 45.150 61.780 45.470 61.840 ;
        RECT 28.680 61.640 35.260 61.780 ;
        RECT 14.790 61.440 15.110 61.500 ;
        RECT 20.770 61.440 21.090 61.500 ;
        RECT 22.625 61.440 22.915 61.485 ;
        RECT 13.040 61.300 20.540 61.440 ;
        RECT 8.825 60.915 9.115 61.145 ;
        RECT 9.730 61.100 10.050 61.160 ;
        RECT 10.205 61.100 10.495 61.145 ;
        RECT 11.110 61.100 11.430 61.160 ;
        RECT 13.040 61.145 13.180 61.300 ;
        RECT 14.790 61.240 15.110 61.300 ;
        RECT 9.730 60.960 11.430 61.100 ;
        RECT 8.900 60.760 9.040 60.915 ;
        RECT 9.730 60.900 10.050 60.960 ;
        RECT 10.205 60.915 10.495 60.960 ;
        RECT 11.110 60.900 11.430 60.960 ;
        RECT 11.585 61.100 11.875 61.145 ;
        RECT 11.585 60.960 12.720 61.100 ;
        RECT 11.585 60.915 11.875 60.960 ;
        RECT 12.030 60.760 12.350 60.820 ;
        RECT 8.900 60.620 12.350 60.760 ;
        RECT 12.030 60.560 12.350 60.620 ;
        RECT 7.905 60.420 8.195 60.465 ;
        RECT 8.350 60.420 8.670 60.480 ;
        RECT 7.905 60.280 8.670 60.420 ;
        RECT 7.905 60.235 8.195 60.280 ;
        RECT 8.350 60.220 8.670 60.280 ;
        RECT 8.810 60.420 9.130 60.480 ;
        RECT 12.580 60.420 12.720 60.960 ;
        RECT 12.965 60.915 13.255 61.145 ;
        RECT 14.345 61.100 14.635 61.145 ;
        RECT 15.250 61.100 15.570 61.160 ;
        RECT 14.345 60.960 15.570 61.100 ;
        RECT 14.345 60.915 14.635 60.960 ;
        RECT 15.250 60.900 15.570 60.960 ;
        RECT 17.105 61.100 17.395 61.145 ;
        RECT 17.640 61.100 18.680 61.110 ;
        RECT 19.850 61.100 20.170 61.160 ;
        RECT 17.105 60.970 20.170 61.100 ;
        RECT 17.105 60.960 17.780 60.970 ;
        RECT 18.540 60.960 20.170 60.970 ;
        RECT 20.400 61.100 20.540 61.300 ;
        RECT 20.770 61.300 22.915 61.440 ;
        RECT 20.770 61.240 21.090 61.300 ;
        RECT 22.625 61.255 22.915 61.300 ;
        RECT 23.990 61.440 24.310 61.500 ;
        RECT 26.380 61.440 26.520 61.640 ;
        RECT 23.990 61.300 26.520 61.440 ;
        RECT 23.990 61.240 24.310 61.300 ;
        RECT 26.750 61.240 27.070 61.500 ;
        RECT 23.070 61.100 23.390 61.160 ;
        RECT 20.400 60.960 23.390 61.100 ;
        RECT 17.105 60.915 17.395 60.960 ;
        RECT 19.850 60.900 20.170 60.960 ;
        RECT 23.070 60.900 23.390 60.960 ;
        RECT 24.925 61.100 25.215 61.145 ;
        RECT 26.840 61.100 26.980 61.240 ;
        RECT 27.300 61.145 27.440 61.640 ;
        RECT 28.130 61.580 28.450 61.640 ;
        RECT 33.650 61.580 33.970 61.640 ;
        RECT 29.050 61.440 29.370 61.500 ;
        RECT 35.120 61.485 35.260 61.640 ;
        RECT 43.860 61.640 45.470 61.780 ;
        RECT 30.445 61.440 30.735 61.485 ;
        RECT 27.755 61.300 28.820 61.440 ;
        RECT 24.925 60.960 26.980 61.100 ;
        RECT 24.925 60.915 25.215 60.960 ;
        RECT 27.225 60.915 27.515 61.145 ;
        RECT 13.410 60.560 13.730 60.820 ;
        RECT 20.770 60.760 21.090 60.820 ;
        RECT 14.420 60.620 21.090 60.760 ;
        RECT 23.160 60.760 23.300 60.900 ;
        RECT 27.755 60.760 27.895 61.300 ;
        RECT 28.680 61.145 28.820 61.300 ;
        RECT 29.050 61.300 30.735 61.440 ;
        RECT 29.050 61.240 29.370 61.300 ;
        RECT 30.445 61.255 30.735 61.300 ;
        RECT 35.045 61.255 35.335 61.485 ;
        RECT 28.145 60.915 28.435 61.145 ;
        RECT 28.605 60.915 28.895 61.145 ;
        RECT 29.525 60.915 29.815 61.145 ;
        RECT 23.160 60.620 27.895 60.760 ;
        RECT 14.420 60.420 14.560 60.620 ;
        RECT 20.770 60.560 21.090 60.620 ;
        RECT 8.810 60.280 14.560 60.420 ;
        RECT 14.790 60.420 15.110 60.480 ;
        RECT 16.185 60.420 16.475 60.465 ;
        RECT 14.790 60.280 16.475 60.420 ;
        RECT 8.810 60.220 9.130 60.280 ;
        RECT 14.790 60.220 15.110 60.280 ;
        RECT 16.185 60.235 16.475 60.280 ;
        RECT 18.470 60.420 18.790 60.480 ;
        RECT 19.390 60.420 19.710 60.480 ;
        RECT 18.470 60.280 19.710 60.420 ;
        RECT 18.470 60.220 18.790 60.280 ;
        RECT 19.390 60.220 19.710 60.280 ;
        RECT 21.690 60.220 22.010 60.480 ;
        RECT 22.165 60.420 22.455 60.465 ;
        RECT 23.990 60.420 24.310 60.480 ;
        RECT 22.165 60.280 24.310 60.420 ;
        RECT 22.165 60.235 22.455 60.280 ;
        RECT 23.990 60.220 24.310 60.280 ;
        RECT 24.910 60.420 25.230 60.480 ;
        RECT 25.845 60.420 26.135 60.465 ;
        RECT 24.910 60.280 26.135 60.420 ;
        RECT 28.200 60.420 28.340 60.915 ;
        RECT 29.600 60.760 29.740 60.915 ;
        RECT 29.970 60.900 30.290 61.160 ;
        RECT 31.350 60.900 31.670 61.160 ;
        RECT 32.730 61.100 33.050 61.160 ;
        RECT 33.205 61.100 33.495 61.145 ;
        RECT 32.730 60.960 33.495 61.100 ;
        RECT 32.730 60.900 33.050 60.960 ;
        RECT 33.205 60.915 33.495 60.960 ;
        RECT 34.110 60.900 34.430 61.160 ;
        RECT 43.860 61.145 44.000 61.640 ;
        RECT 45.150 61.580 45.470 61.640 ;
        RECT 46.530 61.780 46.850 61.840 ;
        RECT 48.460 61.780 48.600 61.980 ;
        RECT 72.765 61.935 73.055 61.980 ;
        RECT 51.590 61.780 51.910 61.840 ;
        RECT 46.530 61.640 48.600 61.780 ;
        RECT 48.960 61.640 51.910 61.780 ;
        RECT 46.530 61.580 46.850 61.640 ;
        RECT 48.370 61.440 48.690 61.500 ;
        RECT 48.960 61.485 49.100 61.640 ;
        RECT 51.590 61.580 51.910 61.640 ;
        RECT 53.430 61.580 53.750 61.840 ;
        RECT 46.620 61.300 48.690 61.440 ;
        RECT 43.785 60.915 44.075 61.145 ;
        RECT 44.230 61.100 44.550 61.160 ;
        RECT 46.620 61.145 46.760 61.300 ;
        RECT 48.370 61.240 48.690 61.300 ;
        RECT 48.845 61.255 49.135 61.485 ;
        RECT 57.110 61.440 57.430 61.500 ;
        RECT 49.380 61.300 57.430 61.440 ;
        RECT 49.380 61.145 49.520 61.300 ;
        RECT 57.110 61.240 57.430 61.300 ;
        RECT 45.165 61.100 45.455 61.145 ;
        RECT 44.230 60.960 45.455 61.100 ;
        RECT 44.230 60.900 44.550 60.960 ;
        RECT 45.165 60.915 45.455 60.960 ;
        RECT 46.545 60.915 46.835 61.145 ;
        RECT 47.925 61.100 48.215 61.145 ;
        RECT 47.925 60.960 49.060 61.100 ;
        RECT 47.925 60.915 48.215 60.960 ;
        RECT 34.200 60.760 34.340 60.900 ;
        RECT 29.600 60.620 34.340 60.760 ;
        RECT 35.030 60.760 35.350 60.820 ;
        RECT 40.550 60.760 40.870 60.820 ;
        RECT 35.030 60.620 40.870 60.760 ;
        RECT 35.030 60.560 35.350 60.620 ;
        RECT 40.550 60.560 40.870 60.620 ;
        RECT 43.310 60.760 43.630 60.820 ;
        RECT 44.705 60.760 44.995 60.805 ;
        RECT 43.310 60.620 44.995 60.760 ;
        RECT 43.310 60.560 43.630 60.620 ;
        RECT 44.705 60.575 44.995 60.620 ;
        RECT 29.510 60.420 29.830 60.480 ;
        RECT 28.200 60.280 29.830 60.420 ;
        RECT 24.910 60.220 25.230 60.280 ;
        RECT 25.845 60.235 26.135 60.280 ;
        RECT 29.510 60.220 29.830 60.280 ;
        RECT 31.810 60.420 32.130 60.480 ;
        RECT 33.205 60.420 33.495 60.465 ;
        RECT 31.810 60.280 33.495 60.420 ;
        RECT 31.810 60.220 32.130 60.280 ;
        RECT 33.205 60.235 33.495 60.280 ;
        RECT 35.950 60.420 36.270 60.480 ;
        RECT 42.850 60.420 43.170 60.480 ;
        RECT 35.950 60.280 43.170 60.420 ;
        RECT 45.240 60.420 45.380 60.915 ;
        RECT 48.920 60.480 49.060 60.960 ;
        RECT 49.305 60.915 49.595 61.145 ;
        RECT 49.945 60.970 50.235 61.115 ;
        RECT 49.945 60.885 50.440 60.970 ;
        RECT 50.685 60.915 50.975 61.145 ;
        RECT 61.710 61.100 62.030 61.160 ;
        RECT 71.845 61.100 72.135 61.145 ;
        RECT 61.710 60.960 72.135 61.100 ;
        RECT 50.020 60.830 50.440 60.885 ;
        RECT 48.370 60.420 48.690 60.480 ;
        RECT 45.240 60.280 48.690 60.420 ;
        RECT 35.950 60.220 36.270 60.280 ;
        RECT 42.850 60.220 43.170 60.280 ;
        RECT 48.370 60.220 48.690 60.280 ;
        RECT 48.830 60.220 49.150 60.480 ;
        RECT 50.300 60.420 50.440 60.830 ;
        RECT 50.760 60.760 50.900 60.915 ;
        RECT 61.710 60.900 62.030 60.960 ;
        RECT 71.845 60.915 72.135 60.960 ;
        RECT 74.130 60.900 74.450 61.160 ;
        RECT 52.510 60.760 52.830 60.820 ;
        RECT 50.760 60.620 52.830 60.760 ;
        RECT 52.510 60.560 52.830 60.620 ;
        RECT 59.885 60.760 60.175 60.805 ;
        RECT 61.250 60.760 61.570 60.820 ;
        RECT 59.885 60.620 61.570 60.760 ;
        RECT 59.885 60.575 60.175 60.620 ;
        RECT 61.250 60.560 61.570 60.620 ;
        RECT 62.170 60.760 62.490 60.820 ;
        RECT 62.170 60.620 66.080 60.760 ;
        RECT 62.170 60.560 62.490 60.620 ;
        RECT 65.940 60.480 66.080 60.620 ;
        RECT 69.070 60.560 69.390 60.820 ;
        RECT 70.465 60.760 70.755 60.805 ;
        RECT 74.220 60.760 74.360 60.900 ;
        RECT 70.465 60.620 74.360 60.760 ;
        RECT 74.605 60.760 74.895 60.805 ;
        RECT 75.970 60.760 76.290 60.820 ;
        RECT 74.605 60.620 76.290 60.760 ;
        RECT 70.465 60.575 70.755 60.620 ;
        RECT 74.605 60.575 74.895 60.620 ;
        RECT 75.970 60.560 76.290 60.620 ;
        RECT 63.550 60.420 63.870 60.480 ;
        RECT 50.300 60.280 63.870 60.420 ;
        RECT 63.550 60.220 63.870 60.280 ;
        RECT 65.850 60.420 66.170 60.480 ;
        RECT 70.925 60.420 71.215 60.465 ;
        RECT 65.850 60.280 71.215 60.420 ;
        RECT 65.850 60.220 66.170 60.280 ;
        RECT 70.925 60.235 71.215 60.280 ;
        RECT 73.210 60.420 73.530 60.480 ;
        RECT 74.145 60.420 74.435 60.465 ;
        RECT 76.430 60.420 76.750 60.480 ;
        RECT 73.210 60.280 76.750 60.420 ;
        RECT 73.210 60.220 73.530 60.280 ;
        RECT 74.145 60.235 74.435 60.280 ;
        RECT 76.430 60.220 76.750 60.280 ;
        RECT 5.520 59.600 76.820 60.080 ;
        RECT 9.730 59.200 10.050 59.460 ;
        RECT 10.650 59.400 10.970 59.460 ;
        RECT 15.250 59.400 15.570 59.460 ;
        RECT 10.650 59.260 15.570 59.400 ;
        RECT 10.650 59.200 10.970 59.260 ;
        RECT 15.250 59.200 15.570 59.260 ;
        RECT 16.630 59.400 16.950 59.460 ;
        RECT 19.865 59.400 20.155 59.445 ;
        RECT 16.630 59.260 20.155 59.400 ;
        RECT 16.630 59.200 16.950 59.260 ;
        RECT 19.865 59.215 20.155 59.260 ;
        RECT 20.785 59.400 21.075 59.445 ;
        RECT 21.690 59.400 22.010 59.460 ;
        RECT 20.785 59.260 22.010 59.400 ;
        RECT 20.785 59.215 21.075 59.260 ;
        RECT 21.690 59.200 22.010 59.260 ;
        RECT 22.625 59.400 22.915 59.445 ;
        RECT 24.450 59.400 24.770 59.460 ;
        RECT 26.765 59.400 27.055 59.445 ;
        RECT 22.625 59.260 27.055 59.400 ;
        RECT 22.625 59.215 22.915 59.260 ;
        RECT 24.450 59.200 24.770 59.260 ;
        RECT 26.765 59.215 27.055 59.260 ;
        RECT 32.270 59.200 32.590 59.460 ;
        RECT 33.650 59.200 33.970 59.460 ;
        RECT 47.910 59.400 48.230 59.460 ;
        RECT 49.750 59.400 50.070 59.460 ;
        RECT 35.120 59.260 38.935 59.400 ;
        RECT 9.820 59.060 9.960 59.200 ;
        RECT 13.410 59.060 13.730 59.120 ;
        RECT 23.085 59.060 23.375 59.105 ;
        RECT 25.830 59.060 26.150 59.120 ;
        RECT 35.120 59.060 35.260 59.260 ;
        RECT 9.820 58.920 11.340 59.060 ;
        RECT 8.350 58.520 8.670 58.780 ;
        RECT 8.825 58.535 9.115 58.765 ;
        RECT 3.750 58.040 4.070 58.100 ;
        RECT 7.445 58.040 7.735 58.085 ;
        RECT 3.750 57.900 7.735 58.040 ;
        RECT 8.900 58.040 9.040 58.535 ;
        RECT 9.730 58.520 10.050 58.780 ;
        RECT 11.200 58.765 11.340 58.920 ;
        RECT 12.120 58.920 13.730 59.060 ;
        RECT 12.120 58.765 12.260 58.920 ;
        RECT 13.410 58.860 13.730 58.920 ;
        RECT 14.090 58.920 22.840 59.060 ;
        RECT 10.665 58.535 10.955 58.765 ;
        RECT 11.125 58.535 11.415 58.765 ;
        RECT 12.045 58.535 12.335 58.765 ;
        RECT 12.965 58.710 13.255 58.765 ;
        RECT 14.090 58.710 14.230 58.920 ;
        RECT 12.965 58.570 14.230 58.710 ;
        RECT 12.965 58.535 13.255 58.570 ;
        RECT 14.970 58.535 15.260 58.765 ;
        RECT 19.405 58.720 19.695 58.765 ;
        RECT 19.850 58.720 20.170 58.780 ;
        RECT 19.405 58.580 20.170 58.720 ;
        RECT 19.405 58.535 19.695 58.580 ;
        RECT 9.285 58.380 9.575 58.425 ;
        RECT 10.740 58.380 10.880 58.535 ;
        RECT 15.045 58.380 15.185 58.535 ;
        RECT 19.850 58.520 20.170 58.580 ;
        RECT 20.325 58.710 20.615 58.765 ;
        RECT 20.770 58.710 21.090 58.780 ;
        RECT 20.325 58.570 21.090 58.710 ;
        RECT 22.700 58.720 22.840 58.920 ;
        RECT 23.085 58.920 25.600 59.060 ;
        RECT 23.085 58.875 23.375 58.920 ;
        RECT 24.910 58.720 25.230 58.780 ;
        RECT 22.700 58.580 25.230 58.720 ;
        RECT 25.460 58.720 25.600 58.920 ;
        RECT 25.830 58.920 35.260 59.060 ;
        RECT 35.490 59.060 35.810 59.120 ;
        RECT 35.490 58.920 37.560 59.060 ;
        RECT 25.830 58.860 26.150 58.920 ;
        RECT 35.490 58.860 35.810 58.920 ;
        RECT 27.225 58.720 27.515 58.765 ;
        RECT 25.460 58.580 28.360 58.720 ;
        RECT 20.325 58.535 20.615 58.570 ;
        RECT 20.770 58.520 21.090 58.570 ;
        RECT 24.910 58.520 25.230 58.580 ;
        RECT 27.225 58.535 27.515 58.580 ;
        RECT 9.285 58.240 10.880 58.380 ;
        RECT 13.500 58.240 15.185 58.380 ;
        RECT 9.285 58.195 9.575 58.240 ;
        RECT 11.570 58.040 11.890 58.100 ;
        RECT 8.900 57.900 11.890 58.040 ;
        RECT 3.750 57.840 4.070 57.900 ;
        RECT 7.445 57.855 7.735 57.900 ;
        RECT 11.570 57.840 11.890 57.900 ;
        RECT 9.730 57.700 10.050 57.760 ;
        RECT 13.500 57.700 13.640 58.240 ;
        RECT 17.565 58.195 17.855 58.425 ;
        RECT 21.230 58.380 21.550 58.440 ;
        RECT 23.545 58.380 23.835 58.425 ;
        RECT 21.230 58.240 23.835 58.380 ;
        RECT 15.710 58.040 16.030 58.100 ;
        RECT 17.105 58.040 17.395 58.085 ;
        RECT 15.710 57.900 17.395 58.040 ;
        RECT 17.640 58.040 17.780 58.195 ;
        RECT 21.230 58.180 21.550 58.240 ;
        RECT 23.545 58.195 23.835 58.240 ;
        RECT 25.830 58.380 26.150 58.440 ;
        RECT 27.685 58.380 27.975 58.425 ;
        RECT 25.830 58.240 27.975 58.380 ;
        RECT 28.220 58.380 28.360 58.580 ;
        RECT 30.890 58.520 31.210 58.780 ;
        RECT 37.420 58.765 37.560 58.920 ;
        RECT 38.795 58.795 38.935 59.260 ;
        RECT 47.910 59.260 50.070 59.400 ;
        RECT 47.910 59.200 48.230 59.260 ;
        RECT 49.750 59.200 50.070 59.260 ;
        RECT 50.210 59.400 50.530 59.460 ;
        RECT 57.570 59.400 57.890 59.460 ;
        RECT 50.210 59.260 57.890 59.400 ;
        RECT 50.210 59.200 50.530 59.260 ;
        RECT 57.570 59.200 57.890 59.260 ;
        RECT 58.490 59.400 58.810 59.460 ;
        RECT 58.490 59.260 63.780 59.400 ;
        RECT 58.490 59.200 58.810 59.260 ;
        RECT 42.405 59.060 42.695 59.105 ;
        RECT 47.005 59.060 47.295 59.105 ;
        RECT 53.890 59.060 54.210 59.120 ;
        RECT 42.405 58.920 46.760 59.060 ;
        RECT 42.405 58.875 42.695 58.920 ;
        RECT 37.345 58.535 37.635 58.765 ;
        RECT 37.805 58.535 38.095 58.765 ;
        RECT 38.720 58.565 39.010 58.795 ;
        RECT 32.270 58.380 32.590 58.440 ;
        RECT 28.220 58.240 32.590 58.380 ;
        RECT 25.830 58.180 26.150 58.240 ;
        RECT 27.685 58.195 27.975 58.240 ;
        RECT 32.270 58.180 32.590 58.240 ;
        RECT 33.205 58.195 33.495 58.425 ;
        RECT 18.470 58.040 18.790 58.100 ;
        RECT 17.640 57.900 18.790 58.040 ;
        RECT 15.710 57.840 16.030 57.900 ;
        RECT 17.105 57.855 17.395 57.900 ;
        RECT 18.470 57.840 18.790 57.900 ;
        RECT 18.930 57.840 19.250 58.100 ;
        RECT 24.910 57.840 25.230 58.100 ;
        RECT 30.890 58.040 31.210 58.100 ;
        RECT 33.280 58.040 33.420 58.195 ;
        RECT 34.570 58.180 34.890 58.440 ;
        RECT 30.890 57.900 33.420 58.040 ;
        RECT 35.045 58.040 35.335 58.085 ;
        RECT 35.490 58.040 35.810 58.100 ;
        RECT 35.045 57.900 35.810 58.040 ;
        RECT 30.890 57.840 31.210 57.900 ;
        RECT 35.045 57.855 35.335 57.900 ;
        RECT 35.490 57.840 35.810 57.900 ;
        RECT 36.410 57.840 36.730 58.100 ;
        RECT 37.880 58.040 38.020 58.535 ;
        RECT 40.550 58.520 40.870 58.780 ;
        RECT 41.485 58.720 41.775 58.765 ;
        RECT 41.945 58.720 42.235 58.765 ;
        RECT 41.485 58.580 42.235 58.720 ;
        RECT 41.485 58.535 41.775 58.580 ;
        RECT 41.945 58.535 42.235 58.580 ;
        RECT 43.310 58.720 43.630 58.780 ;
        RECT 43.785 58.720 44.075 58.765 ;
        RECT 43.310 58.580 44.075 58.720 ;
        RECT 46.620 58.720 46.760 58.920 ;
        RECT 47.005 58.920 54.210 59.060 ;
        RECT 47.005 58.875 47.295 58.920 ;
        RECT 53.890 58.860 54.210 58.920 ;
        RECT 56.665 59.060 56.955 59.105 ;
        RECT 62.170 59.060 62.490 59.120 ;
        RECT 56.665 58.920 62.490 59.060 ;
        RECT 56.665 58.875 56.955 58.920 ;
        RECT 62.170 58.860 62.490 58.920 ;
        RECT 52.970 58.720 53.290 58.780 ;
        RECT 46.620 58.580 53.290 58.720 ;
        RECT 43.310 58.520 43.630 58.580 ;
        RECT 43.785 58.535 44.075 58.580 ;
        RECT 52.970 58.520 53.290 58.580 ;
        RECT 55.730 58.720 56.050 58.780 ;
        RECT 59.885 58.720 60.175 58.765 ;
        RECT 55.730 58.580 60.175 58.720 ;
        RECT 55.730 58.520 56.050 58.580 ;
        RECT 59.885 58.535 60.175 58.580 ;
        RECT 60.790 58.520 61.110 58.780 ;
        RECT 63.090 58.520 63.410 58.780 ;
        RECT 63.640 58.765 63.780 59.260 ;
        RECT 74.590 59.200 74.910 59.460 ;
        RECT 63.565 58.535 63.855 58.765 ;
        RECT 71.830 58.720 72.150 58.780 ;
        RECT 73.685 58.720 73.975 58.765 ;
        RECT 71.830 58.580 73.975 58.720 ;
        RECT 71.830 58.520 72.150 58.580 ;
        RECT 73.685 58.535 73.975 58.580 ;
        RECT 74.145 58.535 74.435 58.765 ;
        RECT 38.250 58.380 38.570 58.440 ;
        RECT 39.185 58.380 39.475 58.425 ;
        RECT 38.250 58.240 39.475 58.380 ;
        RECT 38.250 58.180 38.570 58.240 ;
        RECT 39.185 58.195 39.475 58.240 ;
        RECT 39.630 58.180 39.950 58.440 ;
        RECT 42.850 58.180 43.170 58.440 ;
        RECT 49.290 58.380 49.610 58.440 ;
        RECT 58.490 58.380 58.810 58.440 ;
        RECT 49.290 58.240 58.810 58.380 ;
        RECT 49.290 58.180 49.610 58.240 ;
        RECT 58.490 58.180 58.810 58.240 ;
        RECT 59.405 58.380 59.695 58.425 ;
        RECT 62.185 58.380 62.475 58.425 ;
        RECT 59.405 58.240 62.475 58.380 ;
        RECT 59.405 58.195 59.695 58.240 ;
        RECT 62.185 58.195 62.475 58.240 ;
        RECT 73.210 58.380 73.530 58.440 ;
        RECT 74.220 58.380 74.360 58.535 ;
        RECT 73.210 58.240 74.360 58.380 ;
        RECT 73.210 58.180 73.530 58.240 ;
        RECT 65.850 58.040 66.170 58.100 ;
        RECT 37.880 57.900 66.170 58.040 ;
        RECT 65.850 57.840 66.170 57.900 ;
        RECT 9.730 57.560 13.640 57.700 ;
        RECT 14.345 57.700 14.635 57.745 ;
        RECT 28.590 57.700 28.910 57.760 ;
        RECT 14.345 57.560 28.910 57.700 ;
        RECT 9.730 57.500 10.050 57.560 ;
        RECT 14.345 57.515 14.635 57.560 ;
        RECT 28.590 57.500 28.910 57.560 ;
        RECT 29.985 57.700 30.275 57.745 ;
        RECT 31.810 57.700 32.130 57.760 ;
        RECT 29.985 57.560 32.130 57.700 ;
        RECT 29.985 57.515 30.275 57.560 ;
        RECT 31.810 57.500 32.130 57.560 ;
        RECT 32.730 57.700 33.050 57.760 ;
        RECT 36.005 57.700 36.295 57.745 ;
        RECT 38.250 57.700 38.570 57.760 ;
        RECT 32.730 57.560 38.570 57.700 ;
        RECT 32.730 57.500 33.050 57.560 ;
        RECT 36.005 57.515 36.295 57.560 ;
        RECT 38.250 57.500 38.570 57.560 ;
        RECT 38.710 57.700 39.030 57.760 ;
        RECT 42.850 57.700 43.170 57.760 ;
        RECT 38.710 57.560 43.170 57.700 ;
        RECT 38.710 57.500 39.030 57.560 ;
        RECT 42.850 57.500 43.170 57.560 ;
        RECT 50.225 57.700 50.515 57.745 ;
        RECT 53.430 57.700 53.750 57.760 ;
        RECT 50.225 57.560 53.750 57.700 ;
        RECT 50.225 57.515 50.515 57.560 ;
        RECT 53.430 57.500 53.750 57.560 ;
        RECT 57.570 57.700 57.890 57.760 ;
        RECT 58.505 57.700 58.795 57.745 ;
        RECT 57.570 57.560 58.795 57.700 ;
        RECT 57.570 57.500 57.890 57.560 ;
        RECT 58.505 57.515 58.795 57.560 ;
        RECT 66.310 57.500 66.630 57.760 ;
        RECT 5.520 56.880 76.820 57.360 ;
        RECT 7.430 56.680 7.750 56.740 ;
        RECT 7.905 56.680 8.195 56.725 ;
        RECT 7.430 56.540 8.195 56.680 ;
        RECT 7.430 56.480 7.750 56.540 ;
        RECT 7.905 56.495 8.195 56.540 ;
        RECT 12.950 56.680 13.270 56.740 ;
        RECT 14.345 56.680 14.635 56.725 ;
        RECT 12.950 56.540 14.635 56.680 ;
        RECT 12.950 56.480 13.270 56.540 ;
        RECT 14.345 56.495 14.635 56.540 ;
        RECT 16.170 56.680 16.490 56.740 ;
        RECT 18.945 56.680 19.235 56.725 ;
        RECT 16.170 56.540 19.235 56.680 ;
        RECT 16.170 56.480 16.490 56.540 ;
        RECT 18.945 56.495 19.235 56.540 ;
        RECT 22.610 56.680 22.930 56.740 ;
        RECT 24.450 56.680 24.770 56.740 ;
        RECT 22.610 56.540 24.770 56.680 ;
        RECT 22.610 56.480 22.930 56.540 ;
        RECT 24.450 56.480 24.770 56.540 ;
        RECT 26.305 56.680 26.595 56.725 ;
        RECT 27.670 56.680 27.990 56.740 ;
        RECT 26.305 56.540 27.990 56.680 ;
        RECT 26.305 56.495 26.595 56.540 ;
        RECT 27.670 56.480 27.990 56.540 ;
        RECT 30.890 56.480 31.210 56.740 ;
        RECT 31.350 56.680 31.670 56.740 ;
        RECT 32.285 56.680 32.575 56.725 ;
        RECT 31.350 56.540 32.575 56.680 ;
        RECT 31.350 56.480 31.670 56.540 ;
        RECT 32.285 56.495 32.575 56.540 ;
        RECT 38.250 56.680 38.570 56.740 ;
        RECT 43.325 56.680 43.615 56.725 ;
        RECT 38.250 56.540 43.615 56.680 ;
        RECT 38.250 56.480 38.570 56.540 ;
        RECT 6.970 56.340 7.290 56.400 ;
        RECT 11.125 56.340 11.415 56.385 ;
        RECT 6.970 56.200 11.415 56.340 ;
        RECT 6.970 56.140 7.290 56.200 ;
        RECT 11.125 56.155 11.415 56.200 ;
        RECT 11.570 56.140 11.890 56.400 ;
        RECT 17.105 56.340 17.395 56.385 ;
        RECT 24.910 56.340 25.230 56.400 ;
        RECT 17.105 56.200 25.230 56.340 ;
        RECT 17.105 56.155 17.395 56.200 ;
        RECT 24.910 56.140 25.230 56.200 ;
        RECT 25.385 56.340 25.675 56.385 ;
        RECT 26.750 56.340 27.070 56.400 ;
        RECT 25.385 56.200 27.070 56.340 ;
        RECT 25.385 56.155 25.675 56.200 ;
        RECT 26.750 56.140 27.070 56.200 ;
        RECT 28.590 56.140 28.910 56.400 ;
        RECT 29.970 56.340 30.290 56.400 ;
        RECT 38.710 56.340 39.030 56.400 ;
        RECT 29.970 56.200 39.030 56.340 ;
        RECT 29.970 56.140 30.290 56.200 ;
        RECT 38.710 56.140 39.030 56.200 ;
        RECT 39.185 56.340 39.475 56.385 ;
        RECT 40.090 56.340 40.410 56.400 ;
        RECT 39.185 56.200 40.410 56.340 ;
        RECT 39.185 56.155 39.475 56.200 ;
        RECT 40.090 56.140 40.410 56.200 ;
        RECT 40.550 56.340 40.870 56.400 ;
        RECT 41.945 56.340 42.235 56.385 ;
        RECT 40.550 56.200 42.235 56.340 ;
        RECT 40.550 56.140 40.870 56.200 ;
        RECT 41.945 56.155 42.235 56.200 ;
        RECT 11.660 56.000 11.800 56.140 ;
        RECT 8.900 55.860 11.800 56.000 ;
        RECT 15.710 56.000 16.030 56.060 ;
        RECT 17.565 56.000 17.855 56.045 ;
        RECT 15.710 55.860 17.855 56.000 ;
        RECT 3.750 55.660 4.070 55.720 ;
        RECT 8.900 55.705 9.040 55.860 ;
        RECT 15.710 55.800 16.030 55.860 ;
        RECT 17.565 55.815 17.855 55.860 ;
        RECT 20.770 56.000 21.090 56.060 ;
        RECT 23.085 56.000 23.375 56.045 ;
        RECT 25.830 56.000 26.150 56.060 ;
        RECT 20.770 55.860 26.150 56.000 ;
        RECT 28.680 56.000 28.820 56.140 ;
        RECT 33.665 56.000 33.955 56.045 ;
        RECT 28.680 55.860 33.955 56.000 ;
        RECT 20.770 55.800 21.090 55.860 ;
        RECT 23.085 55.815 23.375 55.860 ;
        RECT 25.830 55.800 26.150 55.860 ;
        RECT 33.665 55.815 33.955 55.860 ;
        RECT 34.110 55.800 34.430 56.060 ;
        RECT 35.030 56.000 35.350 56.060 ;
        RECT 39.645 56.000 39.935 56.045 ;
        RECT 42.480 56.000 42.620 56.540 ;
        RECT 43.325 56.495 43.615 56.540 ;
        RECT 52.510 56.680 52.830 56.740 ;
        RECT 54.365 56.680 54.655 56.725 ;
        RECT 52.510 56.540 54.655 56.680 ;
        RECT 52.510 56.480 52.830 56.540 ;
        RECT 54.365 56.495 54.655 56.540 ;
        RECT 56.650 56.680 56.970 56.740 ;
        RECT 60.790 56.680 61.110 56.740 ;
        RECT 62.185 56.680 62.475 56.725 ;
        RECT 70.450 56.680 70.770 56.740 ;
        RECT 74.145 56.680 74.435 56.725 ;
        RECT 56.650 56.540 62.475 56.680 ;
        RECT 56.650 56.480 56.970 56.540 ;
        RECT 60.790 56.480 61.110 56.540 ;
        RECT 62.185 56.495 62.475 56.540 ;
        RECT 63.180 56.540 74.435 56.680 ;
        RECT 47.450 56.340 47.770 56.400 ;
        RECT 57.570 56.340 57.890 56.400 ;
        RECT 47.450 56.200 57.890 56.340 ;
        RECT 47.450 56.140 47.770 56.200 ;
        RECT 57.570 56.140 57.890 56.200 ;
        RECT 34.665 55.860 35.350 56.000 ;
        RECT 6.985 55.660 7.275 55.705 ;
        RECT 3.750 55.520 7.275 55.660 ;
        RECT 3.750 55.460 4.070 55.520 ;
        RECT 6.985 55.475 7.275 55.520 ;
        RECT 8.825 55.475 9.115 55.705 ;
        RECT 9.730 55.460 10.050 55.720 ;
        RECT 10.665 55.475 10.955 55.705 ;
        RECT 12.045 55.660 12.335 55.705 ;
        RECT 13.410 55.660 13.730 55.720 ;
        RECT 15.250 55.660 15.570 55.720 ;
        RECT 12.045 55.520 13.730 55.660 ;
        RECT 15.055 55.520 15.570 55.660 ;
        RECT 12.045 55.475 12.335 55.520 ;
        RECT 9.285 55.320 9.575 55.365 ;
        RECT 10.740 55.320 10.880 55.475 ;
        RECT 13.410 55.460 13.730 55.520 ;
        RECT 15.250 55.460 15.570 55.520 ;
        RECT 19.390 55.660 19.710 55.720 ;
        RECT 19.865 55.660 20.155 55.705 ;
        RECT 19.390 55.520 20.155 55.660 ;
        RECT 19.390 55.460 19.710 55.520 ;
        RECT 19.865 55.475 20.155 55.520 ;
        RECT 22.625 55.660 22.915 55.705 ;
        RECT 23.530 55.660 23.850 55.720 ;
        RECT 22.625 55.520 23.850 55.660 ;
        RECT 22.625 55.475 22.915 55.520 ;
        RECT 23.530 55.460 23.850 55.520 ;
        RECT 23.990 55.660 24.310 55.720 ;
        RECT 24.465 55.660 24.755 55.705 ;
        RECT 23.990 55.520 24.755 55.660 ;
        RECT 23.990 55.460 24.310 55.520 ;
        RECT 24.465 55.475 24.755 55.520 ;
        RECT 27.210 55.460 27.530 55.720 ;
        RECT 28.590 55.460 28.910 55.720 ;
        RECT 29.050 55.460 29.370 55.720 ;
        RECT 29.970 55.460 30.290 55.720 ;
        RECT 32.730 55.460 33.050 55.720 ;
        RECT 34.665 55.705 34.805 55.860 ;
        RECT 35.030 55.800 35.350 55.860 ;
        RECT 36.960 55.860 39.935 56.000 ;
        RECT 36.960 55.705 37.100 55.860 ;
        RECT 39.645 55.815 39.935 55.860 ;
        RECT 41.100 55.860 42.620 56.000 ;
        RECT 42.850 56.000 43.170 56.060 ;
        RECT 55.730 56.000 56.050 56.060 ;
        RECT 42.850 55.860 56.050 56.000 ;
        RECT 34.590 55.475 34.880 55.705 ;
        RECT 35.505 55.660 35.795 55.705 ;
        RECT 35.965 55.660 36.255 55.705 ;
        RECT 35.505 55.520 36.255 55.660 ;
        RECT 35.505 55.475 35.795 55.520 ;
        RECT 35.965 55.475 36.255 55.520 ;
        RECT 36.885 55.475 37.175 55.705 ;
        RECT 9.285 55.180 10.880 55.320 ;
        RECT 11.570 55.320 11.890 55.380 ;
        RECT 12.490 55.320 12.810 55.380 ;
        RECT 11.570 55.180 12.810 55.320 ;
        RECT 9.285 55.135 9.575 55.180 ;
        RECT 11.570 55.120 11.890 55.180 ;
        RECT 12.490 55.120 12.810 55.180 ;
        RECT 12.965 55.320 13.255 55.365 ;
        RECT 21.230 55.320 21.550 55.380 ;
        RECT 12.965 55.180 21.550 55.320 ;
        RECT 12.965 55.135 13.255 55.180 ;
        RECT 21.230 55.120 21.550 55.180 ;
        RECT 22.165 55.320 22.455 55.365 ;
        RECT 23.070 55.320 23.390 55.380 ;
        RECT 22.165 55.180 23.390 55.320 ;
        RECT 22.165 55.135 22.455 55.180 ;
        RECT 23.070 55.120 23.390 55.180 ;
        RECT 33.650 55.320 33.970 55.380 ;
        RECT 35.580 55.320 35.720 55.475 ;
        RECT 37.330 55.460 37.650 55.720 ;
        RECT 37.975 55.660 38.265 55.705 ;
        RECT 38.710 55.660 39.030 55.720 ;
        RECT 41.100 55.705 41.240 55.860 ;
        RECT 42.850 55.800 43.170 55.860 ;
        RECT 55.730 55.800 56.050 55.860 ;
        RECT 57.110 56.000 57.430 56.060 ;
        RECT 63.180 56.000 63.320 56.540 ;
        RECT 70.450 56.480 70.770 56.540 ;
        RECT 74.145 56.495 74.435 56.540 ;
        RECT 69.530 56.340 69.850 56.400 ;
        RECT 72.750 56.340 73.070 56.400 ;
        RECT 73.685 56.340 73.975 56.385 ;
        RECT 69.530 56.200 72.060 56.340 ;
        RECT 69.530 56.140 69.850 56.200 ;
        RECT 57.110 55.860 63.320 56.000 ;
        RECT 63.550 56.000 63.870 56.060 ;
        RECT 68.150 56.000 68.470 56.060 ;
        RECT 71.920 56.000 72.060 56.200 ;
        RECT 72.750 56.200 73.975 56.340 ;
        RECT 72.750 56.140 73.070 56.200 ;
        RECT 73.685 56.155 73.975 56.200 ;
        RECT 63.550 55.860 71.600 56.000 ;
        RECT 57.110 55.800 57.430 55.860 ;
        RECT 37.975 55.520 39.030 55.660 ;
        RECT 37.975 55.475 38.265 55.520 ;
        RECT 38.710 55.460 39.030 55.520 ;
        RECT 40.565 55.475 40.855 55.705 ;
        RECT 41.025 55.475 41.315 55.705 ;
        RECT 41.470 55.660 41.790 55.720 ;
        RECT 42.405 55.660 42.695 55.705 ;
        RECT 43.785 55.660 44.075 55.705 ;
        RECT 48.830 55.660 49.150 55.720 ;
        RECT 52.510 55.660 52.830 55.720 ;
        RECT 57.660 55.705 57.800 55.860 ;
        RECT 63.550 55.800 63.870 55.860 ;
        RECT 68.150 55.800 68.470 55.860 ;
        RECT 41.470 55.520 42.695 55.660 ;
        RECT 33.650 55.180 35.720 55.320 ;
        RECT 36.410 55.320 36.730 55.380 ;
        RECT 40.640 55.320 40.780 55.475 ;
        RECT 41.470 55.460 41.790 55.520 ;
        RECT 42.405 55.475 42.695 55.520 ;
        RECT 42.940 55.520 52.830 55.660 ;
        RECT 41.560 55.320 41.700 55.460 ;
        RECT 42.940 55.320 43.080 55.520 ;
        RECT 43.785 55.475 44.075 55.520 ;
        RECT 48.830 55.460 49.150 55.520 ;
        RECT 52.510 55.460 52.830 55.520 ;
        RECT 55.285 55.475 55.575 55.705 ;
        RECT 57.585 55.475 57.875 55.705 ;
        RECT 59.885 55.660 60.175 55.705 ;
        RECT 65.850 55.660 66.170 55.720 ;
        RECT 59.885 55.520 66.170 55.660 ;
        RECT 59.885 55.475 60.175 55.520 ;
        RECT 36.410 55.180 40.780 55.320 ;
        RECT 41.100 55.180 41.700 55.320 ;
        RECT 42.020 55.180 43.080 55.320 ;
        RECT 43.310 55.320 43.630 55.380 ;
        RECT 44.230 55.320 44.550 55.380 ;
        RECT 43.310 55.180 44.550 55.320 ;
        RECT 33.650 55.120 33.970 55.180 ;
        RECT 36.410 55.120 36.730 55.180 ;
        RECT 10.650 54.980 10.970 55.040 ;
        RECT 15.265 54.980 15.555 55.025 ;
        RECT 10.650 54.840 15.555 54.980 ;
        RECT 10.650 54.780 10.970 54.840 ;
        RECT 15.265 54.795 15.555 54.840 ;
        RECT 18.470 54.980 18.790 55.040 ;
        RECT 20.325 54.980 20.615 55.025 ;
        RECT 18.470 54.840 20.615 54.980 ;
        RECT 18.470 54.780 18.790 54.840 ;
        RECT 20.325 54.795 20.615 54.840 ;
        RECT 20.770 54.980 21.090 55.040 ;
        RECT 35.490 54.980 35.810 55.040 ;
        RECT 20.770 54.840 35.810 54.980 ;
        RECT 20.770 54.780 21.090 54.840 ;
        RECT 35.490 54.780 35.810 54.840 ;
        RECT 40.090 54.980 40.410 55.040 ;
        RECT 41.100 54.980 41.240 55.180 ;
        RECT 40.090 54.840 41.240 54.980 ;
        RECT 41.470 54.980 41.790 55.040 ;
        RECT 42.020 54.980 42.160 55.180 ;
        RECT 43.310 55.120 43.630 55.180 ;
        RECT 44.230 55.120 44.550 55.180 ;
        RECT 53.890 55.120 54.210 55.380 ;
        RECT 55.360 55.320 55.500 55.475 ;
        RECT 65.850 55.460 66.170 55.520 ;
        RECT 70.450 55.460 70.770 55.720 ;
        RECT 71.460 55.705 71.600 55.860 ;
        RECT 71.920 55.860 72.980 56.000 ;
        RECT 71.920 55.705 72.060 55.860 ;
        RECT 72.840 55.720 72.980 55.860 ;
        RECT 71.385 55.475 71.675 55.705 ;
        RECT 71.845 55.475 72.135 55.705 ;
        RECT 56.650 55.320 56.970 55.380 ;
        RECT 66.770 55.320 67.090 55.380 ;
        RECT 55.360 55.180 67.090 55.320 ;
        RECT 56.650 55.120 56.970 55.180 ;
        RECT 66.770 55.120 67.090 55.180 ;
        RECT 69.530 55.120 69.850 55.380 ;
        RECT 72.310 55.365 72.600 55.595 ;
        RECT 72.750 55.460 73.070 55.720 ;
        RECT 74.145 55.660 74.435 55.705 ;
        RECT 74.590 55.660 74.910 55.720 ;
        RECT 74.145 55.520 74.910 55.660 ;
        RECT 74.145 55.475 74.435 55.520 ;
        RECT 74.590 55.460 74.910 55.520 ;
        RECT 75.050 55.460 75.370 55.720 ;
        RECT 41.470 54.840 42.160 54.980 ;
        RECT 42.850 54.980 43.170 55.040 ;
        RECT 55.270 54.980 55.590 55.040 ;
        RECT 42.850 54.840 55.590 54.980 ;
        RECT 40.090 54.780 40.410 54.840 ;
        RECT 41.470 54.780 41.790 54.840 ;
        RECT 42.850 54.780 43.170 54.840 ;
        RECT 55.270 54.780 55.590 54.840 ;
        RECT 62.630 54.980 62.950 55.040 ;
        RECT 72.385 54.980 72.525 55.365 ;
        RECT 62.630 54.840 72.525 54.980 ;
        RECT 62.630 54.780 62.950 54.840 ;
        RECT 5.520 54.160 76.820 54.640 ;
        RECT 6.050 53.960 6.370 54.020 ;
        RECT 9.285 53.960 9.575 54.005 ;
        RECT 6.050 53.820 9.575 53.960 ;
        RECT 6.050 53.760 6.370 53.820 ;
        RECT 9.285 53.775 9.575 53.820 ;
        RECT 12.965 53.960 13.255 54.005 ;
        RECT 13.410 53.960 13.730 54.020 ;
        RECT 12.965 53.820 13.730 53.960 ;
        RECT 12.965 53.775 13.255 53.820 ;
        RECT 13.410 53.760 13.730 53.820 ;
        RECT 15.250 53.960 15.570 54.020 ;
        RECT 16.185 53.960 16.475 54.005 ;
        RECT 15.250 53.820 16.475 53.960 ;
        RECT 15.250 53.760 15.570 53.820 ;
        RECT 16.185 53.775 16.475 53.820 ;
        RECT 17.550 53.760 17.870 54.020 ;
        RECT 19.405 53.775 19.695 54.005 ;
        RECT 6.510 53.620 6.830 53.680 ;
        RECT 19.480 53.620 19.620 53.775 ;
        RECT 22.610 53.760 22.930 54.020 ;
        RECT 28.590 53.960 28.910 54.020 ;
        RECT 31.825 53.960 32.115 54.005 ;
        RECT 28.590 53.820 32.115 53.960 ;
        RECT 28.590 53.760 28.910 53.820 ;
        RECT 31.825 53.775 32.115 53.820 ;
        RECT 35.505 53.960 35.795 54.005 ;
        RECT 39.170 53.960 39.490 54.020 ;
        RECT 35.505 53.820 39.490 53.960 ;
        RECT 35.505 53.775 35.795 53.820 ;
        RECT 39.170 53.760 39.490 53.820 ;
        RECT 40.105 53.960 40.395 54.005 ;
        RECT 41.470 53.960 41.790 54.020 ;
        RECT 45.610 53.960 45.930 54.020 ;
        RECT 40.105 53.820 41.790 53.960 ;
        RECT 40.105 53.775 40.395 53.820 ;
        RECT 41.470 53.760 41.790 53.820 ;
        RECT 42.940 53.820 45.930 53.960 ;
        RECT 6.510 53.480 19.620 53.620 ;
        RECT 22.150 53.620 22.470 53.680 ;
        RECT 31.350 53.620 31.670 53.680 ;
        RECT 33.190 53.620 33.510 53.680 ;
        RECT 38.710 53.620 39.030 53.680 ;
        RECT 42.940 53.665 43.080 53.820 ;
        RECT 45.610 53.760 45.930 53.820 ;
        RECT 48.370 53.960 48.690 54.020 ;
        RECT 55.730 53.960 56.050 54.020 ;
        RECT 75.050 53.960 75.370 54.020 ;
        RECT 48.370 53.820 53.200 53.960 ;
        RECT 48.370 53.760 48.690 53.820 ;
        RECT 41.025 53.620 41.315 53.665 ;
        RECT 22.150 53.480 32.960 53.620 ;
        RECT 6.510 53.420 6.830 53.480 ;
        RECT 22.150 53.420 22.470 53.480 ;
        RECT 31.350 53.420 31.670 53.480 ;
        RECT 7.890 53.080 8.210 53.340 ;
        RECT 10.190 53.080 10.510 53.340 ;
        RECT 10.650 53.280 10.970 53.340 ;
        RECT 11.125 53.280 11.415 53.325 ;
        RECT 10.650 53.140 11.415 53.280 ;
        RECT 10.650 53.080 10.970 53.140 ;
        RECT 11.125 53.095 11.415 53.140 ;
        RECT 12.490 53.080 12.810 53.340 ;
        RECT 12.950 53.280 13.270 53.340 ;
        RECT 13.425 53.280 13.715 53.325 ;
        RECT 12.950 53.140 13.715 53.280 ;
        RECT 12.950 53.080 13.270 53.140 ;
        RECT 13.425 53.095 13.715 53.140 ;
        RECT 13.870 53.280 14.190 53.340 ;
        RECT 14.805 53.280 15.095 53.325 ;
        RECT 13.870 53.140 15.095 53.280 ;
        RECT 13.870 53.080 14.190 53.140 ;
        RECT 14.805 53.095 15.095 53.140 ;
        RECT 15.265 53.095 15.555 53.325 ;
        RECT 3.290 52.940 3.610 53.000 ;
        RECT 15.340 52.940 15.480 53.095 ;
        RECT 16.630 53.080 16.950 53.340 ;
        RECT 18.010 53.080 18.330 53.340 ;
        RECT 20.310 53.080 20.630 53.340 ;
        RECT 21.705 53.095 21.995 53.325 ;
        RECT 22.625 53.280 22.915 53.325 ;
        RECT 27.670 53.280 27.990 53.340 ;
        RECT 32.820 53.325 32.960 53.480 ;
        RECT 33.190 53.480 37.100 53.620 ;
        RECT 33.190 53.420 33.510 53.480 ;
        RECT 22.625 53.140 27.990 53.280 ;
        RECT 22.625 53.095 22.915 53.140 ;
        RECT 3.290 52.800 15.480 52.940 ;
        RECT 17.090 52.940 17.410 53.000 ;
        RECT 18.485 52.940 18.775 52.985 ;
        RECT 17.090 52.800 18.775 52.940 ;
        RECT 21.780 52.940 21.920 53.095 ;
        RECT 27.670 53.080 27.990 53.140 ;
        RECT 32.745 53.095 33.035 53.325 ;
        RECT 34.110 53.080 34.430 53.340 ;
        RECT 36.410 53.080 36.730 53.340 ;
        RECT 36.960 53.325 37.100 53.480 ;
        RECT 38.710 53.480 41.315 53.620 ;
        RECT 38.710 53.420 39.030 53.480 ;
        RECT 41.025 53.435 41.315 53.480 ;
        RECT 42.865 53.435 43.155 53.665 ;
        RECT 45.150 53.620 45.470 53.680 ;
        RECT 43.400 53.480 45.470 53.620 ;
        RECT 45.700 53.620 45.840 53.760 ;
        RECT 47.910 53.620 48.230 53.680 ;
        RECT 48.830 53.620 49.150 53.680 ;
        RECT 45.700 53.480 47.220 53.620 ;
        RECT 43.400 53.340 43.540 53.480 ;
        RECT 45.150 53.420 45.470 53.480 ;
        RECT 36.885 53.095 37.175 53.325 ;
        RECT 38.250 53.080 38.570 53.340 ;
        RECT 39.645 53.095 39.935 53.325 ;
        RECT 23.530 52.940 23.850 53.000 ;
        RECT 32.285 52.940 32.575 52.985 ;
        RECT 21.780 52.800 32.575 52.940 ;
        RECT 39.720 52.940 39.860 53.095 ;
        RECT 41.470 53.080 41.790 53.340 ;
        RECT 42.405 53.095 42.695 53.325 ;
        RECT 42.480 52.940 42.620 53.095 ;
        RECT 43.310 53.080 43.630 53.340 ;
        RECT 45.625 53.280 45.915 53.325 ;
        RECT 45.240 53.140 45.915 53.280 ;
        RECT 45.240 53.000 45.380 53.140 ;
        RECT 45.625 53.095 45.915 53.140 ;
        RECT 46.530 53.080 46.850 53.340 ;
        RECT 47.080 53.325 47.220 53.480 ;
        RECT 47.910 53.480 49.150 53.620 ;
        RECT 47.910 53.420 48.230 53.480 ;
        RECT 48.830 53.420 49.150 53.480 ;
        RECT 50.210 53.420 50.530 53.680 ;
        RECT 50.670 53.420 50.990 53.680 ;
        RECT 52.510 53.420 52.830 53.680 ;
        RECT 47.005 53.095 47.295 53.325 ;
        RECT 47.465 53.095 47.755 53.325 ;
        RECT 45.150 52.940 45.470 53.000 ;
        RECT 39.720 52.800 42.160 52.940 ;
        RECT 42.480 52.800 45.470 52.940 ;
        RECT 3.290 52.740 3.610 52.800 ;
        RECT 17.090 52.740 17.410 52.800 ;
        RECT 18.485 52.755 18.775 52.800 ;
        RECT 23.530 52.740 23.850 52.800 ;
        RECT 32.285 52.755 32.575 52.800 ;
        RECT 0.070 52.600 0.390 52.660 ;
        RECT 13.885 52.600 14.175 52.645 ;
        RECT 0.070 52.460 14.175 52.600 ;
        RECT 0.070 52.400 0.390 52.460 ;
        RECT 13.885 52.415 14.175 52.460 ;
        RECT 18.010 52.600 18.330 52.660 ;
        RECT 26.290 52.600 26.610 52.660 ;
        RECT 18.010 52.460 26.610 52.600 ;
        RECT 18.010 52.400 18.330 52.460 ;
        RECT 26.290 52.400 26.610 52.460 ;
        RECT 27.670 52.600 27.990 52.660 ;
        RECT 35.950 52.600 36.270 52.660 ;
        RECT 27.670 52.460 36.270 52.600 ;
        RECT 27.670 52.400 27.990 52.460 ;
        RECT 35.950 52.400 36.270 52.460 ;
        RECT 39.185 52.600 39.475 52.645 ;
        RECT 41.470 52.600 41.790 52.660 ;
        RECT 39.185 52.460 41.790 52.600 ;
        RECT 42.020 52.600 42.160 52.800 ;
        RECT 45.150 52.740 45.470 52.800 ;
        RECT 44.705 52.600 44.995 52.645 ;
        RECT 42.020 52.460 44.995 52.600 ;
        RECT 47.540 52.600 47.680 53.095 ;
        RECT 48.370 53.080 48.690 53.340 ;
        RECT 49.750 53.080 50.070 53.340 ;
        RECT 51.605 53.280 51.895 53.325 ;
        RECT 50.760 53.140 51.895 53.280 ;
        RECT 50.760 53.000 50.900 53.140 ;
        RECT 51.605 53.095 51.895 53.140 ;
        RECT 52.050 53.080 52.370 53.340 ;
        RECT 53.060 53.325 53.200 53.820 ;
        RECT 54.900 53.820 56.050 53.960 ;
        RECT 54.900 53.325 55.040 53.820 ;
        RECT 55.730 53.760 56.050 53.820 ;
        RECT 57.200 53.820 75.370 53.960 ;
        RECT 57.200 53.620 57.340 53.820 ;
        RECT 75.050 53.760 75.370 53.820 ;
        RECT 55.360 53.480 57.340 53.620 ;
        RECT 55.360 53.340 55.500 53.480 ;
        RECT 57.570 53.420 57.890 53.680 ;
        RECT 70.910 53.620 71.230 53.680 ;
        RECT 73.225 53.620 73.515 53.665 ;
        RECT 73.670 53.620 73.990 53.680 ;
        RECT 70.910 53.480 73.990 53.620 ;
        RECT 70.910 53.420 71.230 53.480 ;
        RECT 73.225 53.435 73.515 53.480 ;
        RECT 73.670 53.420 73.990 53.480 ;
        RECT 52.985 53.095 53.275 53.325 ;
        RECT 54.825 53.095 55.115 53.325 ;
        RECT 55.270 53.080 55.590 53.340 ;
        RECT 56.650 53.325 56.970 53.340 ;
        RECT 55.745 53.095 56.035 53.325 ;
        RECT 56.635 53.280 56.970 53.325 ;
        RECT 66.770 53.280 67.090 53.340 ;
        RECT 68.165 53.280 68.455 53.325 ;
        RECT 56.635 53.140 57.135 53.280 ;
        RECT 66.770 53.140 68.455 53.280 ;
        RECT 56.635 53.095 56.970 53.140 ;
        RECT 50.670 52.740 50.990 53.000 ;
        RECT 51.590 52.600 51.910 52.660 ;
        RECT 52.970 52.600 53.290 52.660 ;
        RECT 53.445 52.600 53.735 52.645 ;
        RECT 47.540 52.460 52.740 52.600 ;
        RECT 39.185 52.415 39.475 52.460 ;
        RECT 41.470 52.400 41.790 52.460 ;
        RECT 44.705 52.415 44.995 52.460 ;
        RECT 51.590 52.400 51.910 52.460 ;
        RECT 5.590 52.260 5.910 52.320 ;
        RECT 8.825 52.260 9.115 52.305 ;
        RECT 5.590 52.120 9.115 52.260 ;
        RECT 5.590 52.060 5.910 52.120 ;
        RECT 8.825 52.075 9.115 52.120 ;
        RECT 11.585 52.260 11.875 52.305 ;
        RECT 12.950 52.260 13.270 52.320 ;
        RECT 15.250 52.260 15.570 52.320 ;
        RECT 11.585 52.120 15.570 52.260 ;
        RECT 11.585 52.075 11.875 52.120 ;
        RECT 12.950 52.060 13.270 52.120 ;
        RECT 15.250 52.060 15.570 52.120 ;
        RECT 16.170 52.260 16.490 52.320 ;
        RECT 22.150 52.260 22.470 52.320 ;
        RECT 16.170 52.120 22.470 52.260 ;
        RECT 16.170 52.060 16.490 52.120 ;
        RECT 22.150 52.060 22.470 52.120 ;
        RECT 33.650 52.060 33.970 52.320 ;
        RECT 37.345 52.260 37.635 52.305 ;
        RECT 38.710 52.260 39.030 52.320 ;
        RECT 37.345 52.120 39.030 52.260 ;
        RECT 37.345 52.075 37.635 52.120 ;
        RECT 38.710 52.060 39.030 52.120 ;
        RECT 41.025 52.260 41.315 52.305 ;
        RECT 42.850 52.260 43.170 52.320 ;
        RECT 41.025 52.120 43.170 52.260 ;
        RECT 41.025 52.075 41.315 52.120 ;
        RECT 42.850 52.060 43.170 52.120 ;
        RECT 44.245 52.260 44.535 52.305 ;
        RECT 47.910 52.260 48.230 52.320 ;
        RECT 44.245 52.120 48.230 52.260 ;
        RECT 44.245 52.075 44.535 52.120 ;
        RECT 47.910 52.060 48.230 52.120 ;
        RECT 48.830 52.060 49.150 52.320 ;
        RECT 52.600 52.260 52.740 52.460 ;
        RECT 52.970 52.460 53.735 52.600 ;
        RECT 55.820 52.600 55.960 53.095 ;
        RECT 56.650 53.080 56.970 53.095 ;
        RECT 66.770 53.080 67.090 53.140 ;
        RECT 68.165 53.095 68.455 53.140 ;
        RECT 68.610 53.280 68.930 53.340 ;
        RECT 71.385 53.280 71.675 53.325 ;
        RECT 68.610 53.140 71.675 53.280 ;
        RECT 68.610 53.080 68.930 53.140 ;
        RECT 71.385 53.095 71.675 53.140 ;
        RECT 74.145 53.280 74.435 53.325 ;
        RECT 76.890 53.280 77.210 53.340 ;
        RECT 74.145 53.140 77.210 53.280 ;
        RECT 74.145 53.095 74.435 53.140 ;
        RECT 76.890 53.080 77.210 53.140 ;
        RECT 66.325 52.755 66.615 52.985 ;
        RECT 57.110 52.600 57.430 52.660 ;
        RECT 55.820 52.460 57.430 52.600 ;
        RECT 52.970 52.400 53.290 52.460 ;
        RECT 53.445 52.415 53.735 52.460 ;
        RECT 57.110 52.400 57.430 52.460 ;
        RECT 60.330 52.600 60.650 52.660 ;
        RECT 66.400 52.600 66.540 52.755 ;
        RECT 69.990 52.740 70.310 53.000 ;
        RECT 71.830 52.740 72.150 53.000 ;
        RECT 70.080 52.600 70.220 52.740 ;
        RECT 73.670 52.600 73.990 52.660 ;
        RECT 60.330 52.460 73.990 52.600 ;
        RECT 60.330 52.400 60.650 52.460 ;
        RECT 73.670 52.400 73.990 52.460 ;
        RECT 57.570 52.260 57.890 52.320 ;
        RECT 52.600 52.120 57.890 52.260 ;
        RECT 57.570 52.060 57.890 52.120 ;
        RECT 69.990 52.260 70.310 52.320 ;
        RECT 74.605 52.260 74.895 52.305 ;
        RECT 69.990 52.120 74.895 52.260 ;
        RECT 69.990 52.060 70.310 52.120 ;
        RECT 74.605 52.075 74.895 52.120 ;
        RECT 5.520 51.440 76.820 51.920 ;
        RECT 9.730 51.240 10.050 51.300 ;
        RECT 10.665 51.240 10.955 51.285 ;
        RECT 13.870 51.240 14.190 51.300 ;
        RECT 9.730 51.100 14.190 51.240 ;
        RECT 9.730 51.040 10.050 51.100 ;
        RECT 10.665 51.055 10.955 51.100 ;
        RECT 13.870 51.040 14.190 51.100 ;
        RECT 18.010 51.040 18.330 51.300 ;
        RECT 23.990 51.040 24.310 51.300 ;
        RECT 24.540 51.100 25.600 51.240 ;
        RECT 11.585 50.900 11.875 50.945 ;
        RECT 12.490 50.900 12.810 50.960 ;
        RECT 14.790 50.900 15.110 50.960 ;
        RECT 11.585 50.760 15.110 50.900 ;
        RECT 11.585 50.715 11.875 50.760 ;
        RECT 12.490 50.700 12.810 50.760 ;
        RECT 13.410 50.360 13.730 50.620 ;
        RECT 7.905 50.220 8.195 50.265 ;
        RECT 9.270 50.220 9.590 50.280 ;
        RECT 13.500 50.220 13.640 50.360 ;
        RECT 7.905 50.080 13.640 50.220 ;
        RECT 7.905 50.035 8.195 50.080 ;
        RECT 9.270 50.020 9.590 50.080 ;
        RECT 8.825 49.880 9.115 49.925 ;
        RECT 11.110 49.880 11.430 49.940 ;
        RECT 8.825 49.740 11.430 49.880 ;
        RECT 8.825 49.695 9.115 49.740 ;
        RECT 11.110 49.680 11.430 49.740 ;
        RECT 12.965 49.695 13.255 49.925 ;
        RECT 13.425 49.880 13.715 49.925 ;
        RECT 13.960 49.880 14.100 50.760 ;
        RECT 14.790 50.700 15.110 50.760 ;
        RECT 15.250 50.700 15.570 50.960 ;
        RECT 15.710 50.900 16.030 50.960 ;
        RECT 19.390 50.900 19.710 50.960 ;
        RECT 15.710 50.760 19.710 50.900 ;
        RECT 15.710 50.700 16.030 50.760 ;
        RECT 19.390 50.700 19.710 50.760 ;
        RECT 19.865 50.375 20.155 50.605 ;
        RECT 20.310 50.560 20.630 50.620 ;
        RECT 24.540 50.605 24.680 51.100 ;
        RECT 24.925 50.715 25.215 50.945 ;
        RECT 25.460 50.900 25.600 51.100 ;
        RECT 28.590 51.040 28.910 51.300 ;
        RECT 31.810 51.240 32.130 51.300 ;
        RECT 29.140 51.100 32.130 51.240 ;
        RECT 29.140 50.900 29.280 51.100 ;
        RECT 31.810 51.040 32.130 51.100 ;
        RECT 32.285 51.240 32.575 51.285 ;
        RECT 33.650 51.240 33.970 51.300 ;
        RECT 32.285 51.100 33.970 51.240 ;
        RECT 32.285 51.055 32.575 51.100 ;
        RECT 33.650 51.040 33.970 51.100 ;
        RECT 36.410 51.240 36.730 51.300 ;
        RECT 36.885 51.240 37.175 51.285 ;
        RECT 43.325 51.240 43.615 51.285 ;
        RECT 45.610 51.240 45.930 51.300 ;
        RECT 36.410 51.100 37.175 51.240 ;
        RECT 36.410 51.040 36.730 51.100 ;
        RECT 36.885 51.055 37.175 51.100 ;
        RECT 37.420 51.100 45.930 51.240 ;
        RECT 37.420 50.900 37.560 51.100 ;
        RECT 43.325 51.055 43.615 51.100 ;
        RECT 45.610 51.040 45.930 51.100 ;
        RECT 46.530 51.240 46.850 51.300 ;
        RECT 48.370 51.240 48.690 51.300 ;
        RECT 50.670 51.240 50.990 51.300 ;
        RECT 51.590 51.240 51.910 51.300 ;
        RECT 46.530 51.100 48.140 51.240 ;
        RECT 46.530 51.040 46.850 51.100 ;
        RECT 25.460 50.760 29.280 50.900 ;
        RECT 33.740 50.760 37.560 50.900 ;
        RECT 39.170 50.900 39.490 50.960 ;
        RECT 41.470 50.900 41.790 50.960 ;
        RECT 42.405 50.900 42.695 50.945 ;
        RECT 39.170 50.760 41.240 50.900 ;
        RECT 22.165 50.560 22.455 50.605 ;
        RECT 20.310 50.420 22.455 50.560 ;
        RECT 16.645 50.220 16.935 50.265 ;
        RECT 19.940 50.220 20.080 50.375 ;
        RECT 20.310 50.360 20.630 50.420 ;
        RECT 22.165 50.375 22.455 50.420 ;
        RECT 24.465 50.375 24.755 50.605 ;
        RECT 25.000 50.560 25.140 50.715 ;
        RECT 31.810 50.560 32.130 50.620 ;
        RECT 33.740 50.560 33.880 50.760 ;
        RECT 39.170 50.700 39.490 50.760 ;
        RECT 25.000 50.420 30.750 50.560 ;
        RECT 16.645 50.080 20.080 50.220 ;
        RECT 16.645 50.035 16.935 50.080 ;
        RECT 20.770 50.020 21.090 50.280 ;
        RECT 21.230 50.020 21.550 50.280 ;
        RECT 21.690 50.020 22.010 50.280 ;
        RECT 25.830 50.265 26.150 50.280 ;
        RECT 23.085 50.035 23.375 50.265 ;
        RECT 23.545 50.035 23.835 50.265 ;
        RECT 25.820 50.035 26.150 50.265 ;
        RECT 13.425 49.740 14.100 49.880 ;
        RECT 16.170 49.880 16.490 49.940 ;
        RECT 17.105 49.880 17.395 49.925 ;
        RECT 16.170 49.740 17.395 49.880 ;
        RECT 13.425 49.695 13.715 49.740 ;
        RECT 9.730 49.340 10.050 49.600 ;
        RECT 13.040 49.540 13.180 49.695 ;
        RECT 16.170 49.680 16.490 49.740 ;
        RECT 17.105 49.695 17.395 49.740 ;
        RECT 18.025 49.880 18.315 49.925 ;
        RECT 22.610 49.880 22.930 49.940 ;
        RECT 18.025 49.740 22.930 49.880 ;
        RECT 18.025 49.695 18.315 49.740 ;
        RECT 22.610 49.680 22.930 49.740 ;
        RECT 15.250 49.540 15.570 49.600 ;
        RECT 13.040 49.400 15.570 49.540 ;
        RECT 15.250 49.340 15.570 49.400 ;
        RECT 20.310 49.540 20.630 49.600 ;
        RECT 23.160 49.540 23.300 50.035 ;
        RECT 23.620 49.880 23.760 50.035 ;
        RECT 25.830 50.020 26.150 50.035 ;
        RECT 26.290 50.020 26.610 50.280 ;
        RECT 27.670 50.220 27.990 50.280 ;
        RECT 27.475 50.080 27.990 50.220 ;
        RECT 27.670 50.020 27.990 50.080 ;
        RECT 28.130 50.020 28.450 50.280 ;
        RECT 30.610 50.270 30.750 50.420 ;
        RECT 31.810 50.420 33.880 50.560 ;
        RECT 35.045 50.560 35.335 50.605 ;
        RECT 35.950 50.560 36.270 50.620 ;
        RECT 41.100 50.605 41.240 50.760 ;
        RECT 41.470 50.760 42.695 50.900 ;
        RECT 41.470 50.700 41.790 50.760 ;
        RECT 42.405 50.715 42.695 50.760 ;
        RECT 35.045 50.420 36.270 50.560 ;
        RECT 31.810 50.360 32.130 50.420 ;
        RECT 35.045 50.375 35.335 50.420 ;
        RECT 35.950 50.360 36.270 50.420 ;
        RECT 37.805 50.560 38.095 50.605 ;
        RECT 38.265 50.560 38.555 50.605 ;
        RECT 37.805 50.420 38.555 50.560 ;
        RECT 37.805 50.375 38.095 50.420 ;
        RECT 38.265 50.375 38.555 50.420 ;
        RECT 41.025 50.375 41.315 50.605 ;
        RECT 30.610 50.265 31.250 50.270 ;
        RECT 29.525 50.035 29.815 50.265 ;
        RECT 30.610 50.130 31.325 50.265 ;
        RECT 31.035 50.035 31.325 50.130 ;
        RECT 32.730 50.220 33.050 50.280 ;
        RECT 33.205 50.220 33.495 50.265 ;
        RECT 32.730 50.080 33.495 50.220 ;
        RECT 26.380 49.880 26.520 50.020 ;
        RECT 23.620 49.740 26.520 49.880 ;
        RECT 26.765 49.695 27.055 49.925 ;
        RECT 27.210 49.880 27.530 49.940 ;
        RECT 29.600 49.880 29.740 50.035 ;
        RECT 32.730 50.020 33.050 50.080 ;
        RECT 33.205 50.035 33.495 50.080 ;
        RECT 33.650 50.020 33.970 50.280 ;
        RECT 35.490 50.020 35.810 50.280 ;
        RECT 36.425 50.220 36.715 50.265 ;
        RECT 36.870 50.220 37.190 50.280 ;
        RECT 36.425 50.080 37.190 50.220 ;
        RECT 38.340 50.220 38.480 50.375 ;
        RECT 44.705 50.220 44.995 50.265 ;
        RECT 45.150 50.220 45.470 50.280 ;
        RECT 38.340 50.080 45.470 50.220 ;
        RECT 45.700 50.220 45.840 51.040 ;
        RECT 48.000 50.900 48.140 51.100 ;
        RECT 48.370 51.100 51.910 51.240 ;
        RECT 48.370 51.040 48.690 51.100 ;
        RECT 50.670 51.040 50.990 51.100 ;
        RECT 51.590 51.040 51.910 51.100 ;
        RECT 71.830 51.240 72.150 51.300 ;
        RECT 75.050 51.240 75.370 51.300 ;
        RECT 71.830 51.100 75.370 51.240 ;
        RECT 71.830 51.040 72.150 51.100 ;
        RECT 75.050 51.040 75.370 51.100 ;
        RECT 49.305 50.900 49.595 50.945 ;
        RECT 48.000 50.760 49.595 50.900 ;
        RECT 49.305 50.715 49.595 50.760 ;
        RECT 69.530 50.900 69.850 50.960 ;
        RECT 69.530 50.760 72.060 50.900 ;
        RECT 69.530 50.700 69.850 50.760 ;
        RECT 50.210 50.560 50.530 50.620 ;
        RECT 47.540 50.420 50.530 50.560 ;
        RECT 46.545 50.220 46.835 50.265 ;
        RECT 45.700 50.080 46.835 50.220 ;
        RECT 36.425 50.035 36.715 50.080 ;
        RECT 36.870 50.020 37.190 50.080 ;
        RECT 44.705 50.035 44.995 50.080 ;
        RECT 45.150 50.020 45.470 50.080 ;
        RECT 46.545 50.035 46.835 50.080 ;
        RECT 27.210 49.740 29.740 49.880 ;
        RECT 20.310 49.400 23.300 49.540 ;
        RECT 25.370 49.540 25.690 49.600 ;
        RECT 26.840 49.540 26.980 49.695 ;
        RECT 27.210 49.680 27.530 49.740 ;
        RECT 29.970 49.680 30.290 49.940 ;
        RECT 30.430 49.880 30.750 49.940 ;
        RECT 40.565 49.880 40.855 49.925 ;
        RECT 41.470 49.880 41.790 49.940 ;
        RECT 30.430 49.740 41.790 49.880 ;
        RECT 30.430 49.680 30.750 49.740 ;
        RECT 40.565 49.695 40.855 49.740 ;
        RECT 41.470 49.680 41.790 49.740 ;
        RECT 43.310 49.880 43.630 49.940 ;
        RECT 45.625 49.880 45.915 49.925 ;
        RECT 43.310 49.740 45.915 49.880 ;
        RECT 43.310 49.680 43.630 49.740 ;
        RECT 45.625 49.695 45.915 49.740 ;
        RECT 46.085 49.880 46.375 49.925 ;
        RECT 47.540 49.880 47.680 50.420 ;
        RECT 50.210 50.360 50.530 50.420 ;
        RECT 52.050 50.560 52.370 50.620 ;
        RECT 71.920 50.560 72.060 50.760 ;
        RECT 72.750 50.560 73.070 50.620 ;
        RECT 75.050 50.560 75.370 50.620 ;
        RECT 52.050 50.420 71.140 50.560 ;
        RECT 52.050 50.360 52.370 50.420 ;
        RECT 47.910 50.220 48.230 50.280 ;
        RECT 48.830 50.220 49.150 50.280 ;
        RECT 50.685 50.220 50.975 50.265 ;
        RECT 47.910 50.080 48.600 50.220 ;
        RECT 47.910 50.020 48.230 50.080 ;
        RECT 46.085 49.740 47.680 49.880 ;
        RECT 48.460 49.880 48.600 50.080 ;
        RECT 48.830 50.080 50.975 50.220 ;
        RECT 48.830 50.020 49.150 50.080 ;
        RECT 50.685 50.035 50.975 50.080 ;
        RECT 51.325 50.220 51.615 50.265 ;
        RECT 52.510 50.220 52.830 50.280 ;
        RECT 51.325 50.080 52.830 50.220 ;
        RECT 51.325 50.035 51.615 50.080 ;
        RECT 52.510 50.020 52.830 50.080 ;
        RECT 52.970 50.265 53.290 50.280 ;
        RECT 52.970 50.035 53.425 50.265 ;
        RECT 53.905 50.220 54.195 50.265 ;
        RECT 58.490 50.220 58.810 50.280 ;
        RECT 53.905 50.080 58.810 50.220 ;
        RECT 53.905 50.035 54.195 50.080 ;
        RECT 52.970 50.020 53.290 50.035 ;
        RECT 58.490 50.020 58.810 50.080 ;
        RECT 60.330 50.020 60.650 50.280 ;
        RECT 60.790 50.020 61.110 50.280 ;
        RECT 49.305 49.880 49.595 49.925 ;
        RECT 48.460 49.740 49.595 49.880 ;
        RECT 46.085 49.695 46.375 49.740 ;
        RECT 49.305 49.695 49.595 49.740 ;
        RECT 50.210 49.880 50.530 49.940 ;
        RECT 50.210 49.740 70.680 49.880 ;
        RECT 31.810 49.540 32.130 49.600 ;
        RECT 25.370 49.400 32.130 49.540 ;
        RECT 20.310 49.340 20.630 49.400 ;
        RECT 25.370 49.340 25.690 49.400 ;
        RECT 31.810 49.340 32.130 49.400 ;
        RECT 32.270 49.540 32.590 49.600 ;
        RECT 37.805 49.540 38.095 49.585 ;
        RECT 32.270 49.400 38.095 49.540 ;
        RECT 32.270 49.340 32.590 49.400 ;
        RECT 37.805 49.355 38.095 49.400 ;
        RECT 41.010 49.540 41.330 49.600 ;
        RECT 46.160 49.540 46.300 49.695 ;
        RECT 50.210 49.680 50.530 49.740 ;
        RECT 41.010 49.400 46.300 49.540 ;
        RECT 47.465 49.540 47.755 49.585 ;
        RECT 47.910 49.540 48.230 49.600 ;
        RECT 47.465 49.400 48.230 49.540 ;
        RECT 41.010 49.340 41.330 49.400 ;
        RECT 47.465 49.355 47.755 49.400 ;
        RECT 47.910 49.340 48.230 49.400 ;
        RECT 48.385 49.540 48.675 49.585 ;
        RECT 48.830 49.540 49.150 49.600 ;
        RECT 48.385 49.400 49.150 49.540 ;
        RECT 48.385 49.355 48.675 49.400 ;
        RECT 48.830 49.340 49.150 49.400 ;
        RECT 52.065 49.540 52.355 49.585 ;
        RECT 55.730 49.540 56.050 49.600 ;
        RECT 52.065 49.400 56.050 49.540 ;
        RECT 52.065 49.355 52.355 49.400 ;
        RECT 55.730 49.340 56.050 49.400 ;
        RECT 66.770 49.540 67.090 49.600 ;
        RECT 70.540 49.585 70.680 49.740 ;
        RECT 67.245 49.540 67.535 49.585 ;
        RECT 66.770 49.400 67.535 49.540 ;
        RECT 66.770 49.340 67.090 49.400 ;
        RECT 67.245 49.355 67.535 49.400 ;
        RECT 70.465 49.355 70.755 49.585 ;
        RECT 71.000 49.540 71.140 50.420 ;
        RECT 71.920 50.420 73.070 50.560 ;
        RECT 71.385 50.220 71.675 50.265 ;
        RECT 71.920 50.220 72.060 50.420 ;
        RECT 72.750 50.360 73.070 50.420 ;
        RECT 73.300 50.420 75.370 50.560 ;
        RECT 73.300 50.265 73.440 50.420 ;
        RECT 75.050 50.360 75.370 50.420 ;
        RECT 71.385 50.080 72.060 50.220 ;
        RECT 71.385 50.035 71.675 50.080 ;
        RECT 73.225 50.035 73.515 50.265 ;
        RECT 73.685 50.035 73.975 50.265 ;
        RECT 71.830 49.680 72.150 49.940 ;
        RECT 72.305 49.695 72.595 49.925 ;
        RECT 72.750 49.880 73.070 49.940 ;
        RECT 73.760 49.880 73.900 50.035 ;
        RECT 72.750 49.740 73.900 49.880 ;
        RECT 72.380 49.540 72.520 49.695 ;
        RECT 72.750 49.680 73.070 49.740 ;
        RECT 71.000 49.400 72.520 49.540 ;
        RECT 74.590 49.340 74.910 49.600 ;
        RECT 5.520 48.720 76.820 49.200 ;
        RECT 22.165 48.520 22.455 48.565 ;
        RECT 23.070 48.520 23.390 48.580 ;
        RECT 22.165 48.380 23.390 48.520 ;
        RECT 22.165 48.335 22.455 48.380 ;
        RECT 23.070 48.320 23.390 48.380 ;
        RECT 28.130 48.520 28.450 48.580 ;
        RECT 35.965 48.520 36.255 48.565 ;
        RECT 36.870 48.520 37.190 48.580 ;
        RECT 37.790 48.520 38.110 48.580 ;
        RECT 45.610 48.520 45.930 48.580 ;
        RECT 47.465 48.520 47.755 48.565 ;
        RECT 28.130 48.380 35.260 48.520 ;
        RECT 28.130 48.320 28.450 48.380 ;
        RECT 17.090 48.180 17.410 48.240 ;
        RECT 14.420 48.040 17.410 48.180 ;
        RECT 0.990 47.840 1.310 47.900 ;
        RECT 6.985 47.840 7.275 47.885 ;
        RECT 0.990 47.700 7.275 47.840 ;
        RECT 0.990 47.640 1.310 47.700 ;
        RECT 6.985 47.655 7.275 47.700 ;
        RECT 9.270 47.640 9.590 47.900 ;
        RECT 10.055 47.840 10.345 47.885 ;
        RECT 12.030 47.840 12.350 47.900 ;
        RECT 10.055 47.700 12.350 47.840 ;
        RECT 10.055 47.655 10.345 47.700 ;
        RECT 12.030 47.640 12.350 47.700 ;
        RECT 12.950 47.640 13.270 47.900 ;
        RECT 14.420 47.885 14.560 48.040 ;
        RECT 17.090 47.980 17.410 48.040 ;
        RECT 31.810 48.180 32.130 48.240 ;
        RECT 33.665 48.180 33.955 48.225 ;
        RECT 31.810 48.040 33.955 48.180 ;
        RECT 31.810 47.980 32.130 48.040 ;
        RECT 33.665 47.995 33.955 48.040 ;
        RECT 34.110 48.180 34.430 48.240 ;
        RECT 34.585 48.180 34.875 48.225 ;
        RECT 34.110 48.040 34.875 48.180 ;
        RECT 34.110 47.980 34.430 48.040 ;
        RECT 34.585 47.995 34.875 48.040 ;
        RECT 14.345 47.655 14.635 47.885 ;
        RECT 14.805 47.655 15.095 47.885 ;
        RECT 4.210 47.500 4.530 47.560 ;
        RECT 14.880 47.500 15.020 47.655 ;
        RECT 21.230 47.640 21.550 47.900 ;
        RECT 22.150 47.840 22.470 47.900 ;
        RECT 24.450 47.840 24.770 47.900 ;
        RECT 22.150 47.700 24.770 47.840 ;
        RECT 22.150 47.640 22.470 47.700 ;
        RECT 24.450 47.640 24.770 47.700 ;
        RECT 32.730 47.640 33.050 47.900 ;
        RECT 33.190 47.640 33.510 47.900 ;
        RECT 35.120 47.885 35.260 48.380 ;
        RECT 35.965 48.380 41.240 48.520 ;
        RECT 35.965 48.335 36.255 48.380 ;
        RECT 36.870 48.320 37.190 48.380 ;
        RECT 37.790 48.320 38.110 48.380 ;
        RECT 35.490 48.180 35.810 48.240 ;
        RECT 39.185 48.180 39.475 48.225 ;
        RECT 35.490 48.040 39.475 48.180 ;
        RECT 41.100 48.180 41.240 48.380 ;
        RECT 45.610 48.380 47.755 48.520 ;
        RECT 45.610 48.320 45.930 48.380 ;
        RECT 46.160 48.180 46.300 48.380 ;
        RECT 47.465 48.335 47.755 48.380 ;
        RECT 47.910 48.520 48.230 48.580 ;
        RECT 47.910 48.380 49.520 48.520 ;
        RECT 47.910 48.320 48.230 48.380 ;
        RECT 49.380 48.225 49.520 48.380 ;
        RECT 41.100 48.040 46.300 48.180 ;
        RECT 35.490 47.980 35.810 48.040 ;
        RECT 39.185 47.995 39.475 48.040 ;
        RECT 49.305 47.995 49.595 48.225 ;
        RECT 50.210 48.170 50.530 48.430 ;
        RECT 52.510 48.320 52.830 48.580 ;
        RECT 57.570 48.520 57.890 48.580 ;
        RECT 75.050 48.520 75.370 48.580 ;
        RECT 57.570 48.380 75.370 48.520 ;
        RECT 57.570 48.320 57.890 48.380 ;
        RECT 75.050 48.320 75.370 48.380 ;
        RECT 50.225 47.995 50.515 48.170 ;
        RECT 35.045 47.840 35.335 47.885 ;
        RECT 35.045 47.700 35.720 47.840 ;
        RECT 35.045 47.655 35.335 47.700 ;
        RECT 4.210 47.360 15.020 47.500 ;
        RECT 21.320 47.500 21.460 47.640 ;
        RECT 23.530 47.500 23.850 47.560 ;
        RECT 21.320 47.360 23.850 47.500 ;
        RECT 4.210 47.300 4.530 47.360 ;
        RECT 23.530 47.300 23.850 47.360 ;
        RECT 27.670 47.500 27.990 47.560 ;
        RECT 29.050 47.500 29.370 47.560 ;
        RECT 27.670 47.360 29.370 47.500 ;
        RECT 27.670 47.300 27.990 47.360 ;
        RECT 29.050 47.300 29.370 47.360 ;
        RECT 29.970 47.500 30.290 47.560 ;
        RECT 33.280 47.500 33.420 47.640 ;
        RECT 29.970 47.360 33.420 47.500 ;
        RECT 29.970 47.300 30.290 47.360 ;
        RECT 11.110 46.960 11.430 47.220 ;
        RECT 13.410 46.960 13.730 47.220 ;
        RECT 15.710 46.960 16.030 47.220 ;
        RECT 31.825 46.975 32.115 47.205 ;
        RECT 33.650 47.160 33.970 47.220 ;
        RECT 35.045 47.160 35.335 47.205 ;
        RECT 33.650 47.020 35.335 47.160 ;
        RECT 35.580 47.160 35.720 47.700 ;
        RECT 36.410 47.640 36.730 47.900 ;
        RECT 38.710 47.640 39.030 47.900 ;
        RECT 39.645 47.655 39.935 47.885 ;
        RECT 36.870 47.500 37.190 47.560 ;
        RECT 39.720 47.500 39.860 47.655 ;
        RECT 41.010 47.640 41.330 47.900 ;
        RECT 41.470 47.640 41.790 47.900 ;
        RECT 42.390 47.640 42.710 47.900 ;
        RECT 43.310 47.640 43.630 47.900 ;
        RECT 43.770 47.640 44.090 47.900 ;
        RECT 45.165 47.840 45.455 47.885 ;
        RECT 45.700 47.840 46.760 47.845 ;
        RECT 45.165 47.705 46.760 47.840 ;
        RECT 45.165 47.700 45.840 47.705 ;
        RECT 45.165 47.655 45.455 47.700 ;
        RECT 36.870 47.360 39.860 47.500 ;
        RECT 41.560 47.500 41.700 47.640 ;
        RECT 43.400 47.500 43.540 47.640 ;
        RECT 41.560 47.360 43.540 47.500 ;
        RECT 36.870 47.300 37.190 47.360 ;
        RECT 45.625 47.315 45.915 47.545 ;
        RECT 46.620 47.500 46.760 47.705 ;
        RECT 47.910 47.640 48.230 47.900 ;
        RECT 50.685 47.840 50.975 47.885 ;
        RECT 48.845 47.740 49.135 47.835 ;
        RECT 48.845 47.605 49.520 47.740 ;
        RECT 48.920 47.600 49.520 47.605 ;
        RECT 49.380 47.500 49.520 47.600 ;
        RECT 50.300 47.700 50.975 47.840 ;
        RECT 50.300 47.560 50.440 47.700 ;
        RECT 50.685 47.655 50.975 47.700 ;
        RECT 51.325 47.840 51.615 47.885 ;
        RECT 52.600 47.840 52.740 48.320 ;
        RECT 60.345 48.180 60.635 48.225 ;
        RECT 61.250 48.180 61.570 48.240 ;
        RECT 60.345 48.040 61.570 48.180 ;
        RECT 60.345 47.995 60.635 48.040 ;
        RECT 61.250 47.980 61.570 48.040 ;
        RECT 68.150 47.980 68.470 48.240 ;
        RECT 51.325 47.700 52.740 47.840 ;
        RECT 52.970 47.840 53.290 47.900 ;
        RECT 53.905 47.840 54.195 47.885 ;
        RECT 52.970 47.700 54.195 47.840 ;
        RECT 51.325 47.655 51.615 47.700 ;
        RECT 52.970 47.640 53.290 47.700 ;
        RECT 53.905 47.655 54.195 47.700 ;
        RECT 55.745 47.840 56.035 47.885 ;
        RECT 57.110 47.840 57.430 47.900 ;
        RECT 55.745 47.700 57.430 47.840 ;
        RECT 55.745 47.655 56.035 47.700 ;
        RECT 57.110 47.640 57.430 47.700 ;
        RECT 59.425 47.655 59.715 47.885 ;
        RECT 66.770 47.840 67.090 47.900 ;
        RECT 70.465 47.840 70.755 47.885 ;
        RECT 72.765 47.840 73.055 47.885 ;
        RECT 66.770 47.700 70.755 47.840 ;
        RECT 50.210 47.500 50.530 47.560 ;
        RECT 46.620 47.360 47.220 47.500 ;
        RECT 49.380 47.360 50.530 47.500 ;
        RECT 38.710 47.160 39.030 47.220 ;
        RECT 35.580 47.020 39.030 47.160 ;
        RECT 7.905 46.820 8.195 46.865 ;
        RECT 8.350 46.820 8.670 46.880 ;
        RECT 10.650 46.820 10.970 46.880 ;
        RECT 7.905 46.680 10.970 46.820 ;
        RECT 7.905 46.635 8.195 46.680 ;
        RECT 8.350 46.620 8.670 46.680 ;
        RECT 10.650 46.620 10.970 46.680 ;
        RECT 12.030 46.820 12.350 46.880 ;
        RECT 27.210 46.820 27.530 46.880 ;
        RECT 12.030 46.680 27.530 46.820 ;
        RECT 31.900 46.820 32.040 46.975 ;
        RECT 33.650 46.960 33.970 47.020 ;
        RECT 35.045 46.975 35.335 47.020 ;
        RECT 38.710 46.960 39.030 47.020 ;
        RECT 40.105 47.160 40.395 47.205 ;
        RECT 41.010 47.160 41.330 47.220 ;
        RECT 40.105 47.020 41.330 47.160 ;
        RECT 40.105 46.975 40.395 47.020 ;
        RECT 41.010 46.960 41.330 47.020 ;
        RECT 41.485 47.160 41.775 47.205 ;
        RECT 41.930 47.160 42.250 47.220 ;
        RECT 41.485 47.020 42.250 47.160 ;
        RECT 41.485 46.975 41.775 47.020 ;
        RECT 41.930 46.960 42.250 47.020 ;
        RECT 42.865 47.160 43.155 47.205 ;
        RECT 44.690 47.160 45.010 47.220 ;
        RECT 42.865 47.020 45.010 47.160 ;
        RECT 42.865 46.975 43.155 47.020 ;
        RECT 44.690 46.960 45.010 47.020 ;
        RECT 34.110 46.820 34.430 46.880 ;
        RECT 39.170 46.820 39.490 46.880 ;
        RECT 31.900 46.680 39.490 46.820 ;
        RECT 12.030 46.620 12.350 46.680 ;
        RECT 27.210 46.620 27.530 46.680 ;
        RECT 34.110 46.620 34.430 46.680 ;
        RECT 39.170 46.620 39.490 46.680 ;
        RECT 43.310 46.820 43.630 46.880 ;
        RECT 44.245 46.820 44.535 46.865 ;
        RECT 43.310 46.680 44.535 46.820 ;
        RECT 45.700 46.820 45.840 47.315 ;
        RECT 47.080 47.160 47.220 47.360 ;
        RECT 50.210 47.300 50.530 47.360 ;
        RECT 52.510 47.500 52.830 47.560 ;
        RECT 53.445 47.500 53.735 47.545 ;
        RECT 52.510 47.360 53.735 47.500 ;
        RECT 52.510 47.300 52.830 47.360 ;
        RECT 53.445 47.315 53.735 47.360 ;
        RECT 54.810 47.500 55.130 47.560 ;
        RECT 55.285 47.500 55.575 47.545 ;
        RECT 54.810 47.360 55.575 47.500 ;
        RECT 54.810 47.300 55.130 47.360 ;
        RECT 55.285 47.315 55.575 47.360 ;
        RECT 49.305 47.160 49.595 47.205 ;
        RECT 47.080 47.020 49.595 47.160 ;
        RECT 49.305 46.975 49.595 47.020 ;
        RECT 50.670 47.160 50.990 47.220 ;
        RECT 52.600 47.160 52.740 47.300 ;
        RECT 50.670 47.020 52.740 47.160 ;
        RECT 50.670 46.960 50.990 47.020 ;
        RECT 47.910 46.820 48.230 46.880 ;
        RECT 45.700 46.680 48.230 46.820 ;
        RECT 43.310 46.620 43.630 46.680 ;
        RECT 44.245 46.635 44.535 46.680 ;
        RECT 47.910 46.620 48.230 46.680 ;
        RECT 48.370 46.620 48.690 46.880 ;
        RECT 48.830 46.820 49.150 46.880 ;
        RECT 49.750 46.820 50.070 46.880 ;
        RECT 48.830 46.680 50.070 46.820 ;
        RECT 55.360 46.820 55.500 47.315 ;
        RECT 59.500 47.160 59.640 47.655 ;
        RECT 66.770 47.640 67.090 47.700 ;
        RECT 70.465 47.655 70.755 47.700 ;
        RECT 71.460 47.700 73.055 47.840 ;
        RECT 69.070 47.500 69.390 47.560 ;
        RECT 70.925 47.500 71.215 47.545 ;
        RECT 69.070 47.360 71.215 47.500 ;
        RECT 69.070 47.300 69.390 47.360 ;
        RECT 70.925 47.315 71.215 47.360 ;
        RECT 70.450 47.160 70.770 47.220 ;
        RECT 59.500 47.020 70.770 47.160 ;
        RECT 70.450 46.960 70.770 47.020 ;
        RECT 62.630 46.820 62.950 46.880 ;
        RECT 55.360 46.680 62.950 46.820 ;
        RECT 48.830 46.620 49.150 46.680 ;
        RECT 49.750 46.620 50.070 46.680 ;
        RECT 62.630 46.620 62.950 46.680 ;
        RECT 68.150 46.820 68.470 46.880 ;
        RECT 71.460 46.820 71.600 47.700 ;
        RECT 72.765 47.655 73.055 47.700 ;
        RECT 68.150 46.680 71.600 46.820 ;
        RECT 68.150 46.620 68.470 46.680 ;
        RECT 5.520 46.000 76.820 46.480 ;
        RECT 21.245 45.800 21.535 45.845 ;
        RECT 27.670 45.800 27.990 45.860 ;
        RECT 21.245 45.660 27.990 45.800 ;
        RECT 21.245 45.615 21.535 45.660 ;
        RECT 27.670 45.600 27.990 45.660 ;
        RECT 30.890 45.800 31.210 45.860 ;
        RECT 36.410 45.800 36.730 45.860 ;
        RECT 30.890 45.660 36.730 45.800 ;
        RECT 30.890 45.600 31.210 45.660 ;
        RECT 36.410 45.600 36.730 45.660 ;
        RECT 40.550 45.800 40.870 45.860 ;
        RECT 41.025 45.800 41.315 45.845 ;
        RECT 40.550 45.660 41.315 45.800 ;
        RECT 40.550 45.600 40.870 45.660 ;
        RECT 41.025 45.615 41.315 45.660 ;
        RECT 41.560 45.660 42.620 45.800 ;
        RECT 21.690 45.460 22.010 45.520 ;
        RECT 32.270 45.460 32.590 45.520 ;
        RECT 9.360 45.320 32.590 45.460 ;
        RECT 7.890 45.120 8.210 45.180 ;
        RECT 9.360 45.120 9.500 45.320 ;
        RECT 21.690 45.260 22.010 45.320 ;
        RECT 32.270 45.260 32.590 45.320 ;
        RECT 35.490 45.460 35.810 45.520 ;
        RECT 40.090 45.460 40.410 45.520 ;
        RECT 41.560 45.460 41.700 45.660 ;
        RECT 35.490 45.320 41.700 45.460 ;
        RECT 35.490 45.260 35.810 45.320 ;
        RECT 40.090 45.260 40.410 45.320 ;
        RECT 41.945 45.275 42.235 45.505 ;
        RECT 7.890 44.980 9.500 45.120 ;
        RECT 7.890 44.920 8.210 44.980 ;
        RECT 8.810 44.580 9.130 44.840 ;
        RECT 9.360 44.825 9.500 44.980 ;
        RECT 10.190 44.920 10.510 45.180 ;
        RECT 14.330 45.120 14.650 45.180 ;
        RECT 17.550 45.120 17.870 45.180 ;
        RECT 14.330 44.980 20.540 45.120 ;
        RECT 14.330 44.920 14.650 44.980 ;
        RECT 17.550 44.920 17.870 44.980 ;
        RECT 9.285 44.595 9.575 44.825 ;
        RECT 10.650 44.580 10.970 44.840 ;
        RECT 18.930 44.580 19.250 44.840 ;
        RECT 20.400 44.825 20.540 44.980 ;
        RECT 26.290 44.920 26.610 45.180 ;
        RECT 27.210 45.120 27.530 45.180 ;
        RECT 41.470 45.120 41.790 45.180 ;
        RECT 27.210 44.980 41.790 45.120 ;
        RECT 27.210 44.920 27.530 44.980 ;
        RECT 41.470 44.920 41.790 44.980 ;
        RECT 20.325 44.595 20.615 44.825 ;
        RECT 23.530 44.780 23.850 44.840 ;
        RECT 25.845 44.780 26.135 44.825 ;
        RECT 23.530 44.640 26.135 44.780 ;
        RECT 23.530 44.580 23.850 44.640 ;
        RECT 25.845 44.595 26.135 44.640 ;
        RECT 26.750 44.580 27.070 44.840 ;
        RECT 39.645 44.730 39.935 44.825 ;
        RECT 41.025 44.780 41.315 44.825 ;
        RECT 42.020 44.780 42.160 45.275 ;
        RECT 42.480 45.120 42.620 45.660 ;
        RECT 47.450 45.600 47.770 45.860 ;
        RECT 49.305 45.800 49.595 45.845 ;
        RECT 50.210 45.800 50.530 45.860 ;
        RECT 49.305 45.660 50.530 45.800 ;
        RECT 49.305 45.615 49.595 45.660 ;
        RECT 50.210 45.600 50.530 45.660 ;
        RECT 50.670 45.800 50.990 45.860 ;
        RECT 51.590 45.800 51.910 45.860 ;
        RECT 50.670 45.660 51.910 45.800 ;
        RECT 50.670 45.600 50.990 45.660 ;
        RECT 51.590 45.600 51.910 45.660 ;
        RECT 54.365 45.800 54.655 45.845 ;
        RECT 54.365 45.660 58.260 45.800 ;
        RECT 54.365 45.615 54.655 45.660 ;
        RECT 46.070 45.460 46.390 45.520 ;
        RECT 47.925 45.460 48.215 45.505 ;
        RECT 46.070 45.320 48.215 45.460 ;
        RECT 46.070 45.260 46.390 45.320 ;
        RECT 47.925 45.275 48.215 45.320 ;
        RECT 54.350 45.120 54.670 45.180 ;
        RECT 58.120 45.165 58.260 45.660 ;
        RECT 62.170 45.600 62.490 45.860 ;
        RECT 69.530 45.800 69.850 45.860 ;
        RECT 71.385 45.800 71.675 45.845 ;
        RECT 69.530 45.660 71.675 45.800 ;
        RECT 69.530 45.600 69.850 45.660 ;
        RECT 71.385 45.615 71.675 45.660 ;
        RECT 74.145 45.800 74.435 45.845 ;
        RECT 75.510 45.800 75.830 45.860 ;
        RECT 74.145 45.660 75.830 45.800 ;
        RECT 74.145 45.615 74.435 45.660 ;
        RECT 75.510 45.600 75.830 45.660 ;
        RECT 58.950 45.260 59.270 45.520 ;
        RECT 64.010 45.460 64.330 45.520 ;
        RECT 72.750 45.460 73.070 45.520 ;
        RECT 59.500 45.320 64.330 45.460 ;
        RECT 55.285 45.120 55.575 45.165 ;
        RECT 58.045 45.120 58.335 45.165 ;
        RECT 59.500 45.120 59.640 45.320 ;
        RECT 64.010 45.260 64.330 45.320 ;
        RECT 64.560 45.320 73.070 45.460 ;
        RECT 42.480 44.980 54.120 45.120 ;
        RECT 39.645 44.595 40.320 44.730 ;
        RECT 41.025 44.640 42.160 44.780 ;
        RECT 41.025 44.595 41.315 44.640 ;
        RECT 39.720 44.590 40.320 44.595 ;
        RECT 8.350 44.440 8.670 44.500 ;
        RECT 27.210 44.440 27.530 44.500 ;
        RECT 36.870 44.440 37.190 44.500 ;
        RECT 39.170 44.440 39.490 44.500 ;
        RECT 8.350 44.300 27.530 44.440 ;
        RECT 8.350 44.240 8.670 44.300 ;
        RECT 27.210 44.240 27.530 44.300 ;
        RECT 30.980 44.300 39.490 44.440 ;
        RECT 40.180 44.440 40.320 44.590 ;
        RECT 43.310 44.580 43.630 44.840 ;
        RECT 45.150 44.580 45.470 44.840 ;
        RECT 46.545 44.780 46.835 44.825 ;
        RECT 46.990 44.780 47.310 44.840 ;
        RECT 46.545 44.640 47.310 44.780 ;
        RECT 46.545 44.595 46.835 44.640 ;
        RECT 46.990 44.580 47.310 44.640 ;
        RECT 48.830 44.580 49.150 44.840 ;
        RECT 49.290 44.780 49.610 44.840 ;
        RECT 50.225 44.780 50.515 44.825 ;
        RECT 49.290 44.640 50.515 44.780 ;
        RECT 49.290 44.580 49.610 44.640 ;
        RECT 50.225 44.595 50.515 44.640 ;
        RECT 51.130 44.580 51.450 44.840 ;
        RECT 52.065 44.595 52.355 44.825 ;
        RECT 41.470 44.440 41.790 44.500 ;
        RECT 40.180 44.300 41.790 44.440 ;
        RECT 7.905 44.100 8.195 44.145 ;
        RECT 16.170 44.100 16.490 44.160 ;
        RECT 7.905 43.960 16.490 44.100 ;
        RECT 7.905 43.915 8.195 43.960 ;
        RECT 16.170 43.900 16.490 43.960 ;
        RECT 18.010 44.100 18.330 44.160 ;
        RECT 19.405 44.100 19.695 44.145 ;
        RECT 18.010 43.960 19.695 44.100 ;
        RECT 18.010 43.900 18.330 43.960 ;
        RECT 19.405 43.915 19.695 43.960 ;
        RECT 19.850 44.100 20.170 44.160 ;
        RECT 30.980 44.100 31.120 44.300 ;
        RECT 36.870 44.240 37.190 44.300 ;
        RECT 39.170 44.240 39.490 44.300 ;
        RECT 41.470 44.240 41.790 44.300 ;
        RECT 41.930 44.240 42.250 44.500 ;
        RECT 47.910 44.440 48.230 44.500 ;
        RECT 49.380 44.440 49.520 44.580 ;
        RECT 42.480 44.300 49.520 44.440 ;
        RECT 19.850 43.960 31.120 44.100 ;
        RECT 31.350 44.100 31.670 44.160 ;
        RECT 40.105 44.100 40.395 44.145 ;
        RECT 40.550 44.100 40.870 44.160 ;
        RECT 31.350 43.960 40.870 44.100 ;
        RECT 19.850 43.900 20.170 43.960 ;
        RECT 31.350 43.900 31.670 43.960 ;
        RECT 40.105 43.915 40.395 43.960 ;
        RECT 40.550 43.900 40.870 43.960 ;
        RECT 41.010 44.100 41.330 44.160 ;
        RECT 42.480 44.100 42.620 44.300 ;
        RECT 47.910 44.240 48.230 44.300 ;
        RECT 50.670 44.240 50.990 44.500 ;
        RECT 52.140 44.440 52.280 44.595 ;
        RECT 53.430 44.580 53.750 44.840 ;
        RECT 53.980 44.825 54.120 44.980 ;
        RECT 54.350 44.980 55.575 45.120 ;
        RECT 54.350 44.920 54.670 44.980 ;
        RECT 55.285 44.935 55.575 44.980 ;
        RECT 56.280 44.980 57.340 45.120 ;
        RECT 56.280 44.825 56.420 44.980 ;
        RECT 53.905 44.595 54.195 44.825 ;
        RECT 56.205 44.595 56.495 44.825 ;
        RECT 56.665 44.595 56.955 44.825 ;
        RECT 57.200 44.780 57.340 44.980 ;
        RECT 58.045 44.980 59.640 45.120 ;
        RECT 59.885 45.120 60.175 45.165 ;
        RECT 60.790 45.120 61.110 45.180 ;
        RECT 59.885 44.980 61.110 45.120 ;
        RECT 58.045 44.935 58.335 44.980 ;
        RECT 59.885 44.935 60.175 44.980 ;
        RECT 60.790 44.920 61.110 44.980 ;
        RECT 61.250 45.120 61.570 45.180 ;
        RECT 64.560 45.120 64.700 45.320 ;
        RECT 72.750 45.260 73.070 45.320 ;
        RECT 74.590 45.260 74.910 45.520 ;
        RECT 61.250 44.980 64.700 45.120 ;
        RECT 69.070 45.120 69.390 45.180 ;
        RECT 73.685 45.120 73.975 45.165 ;
        RECT 76.890 45.120 77.210 45.180 ;
        RECT 69.070 44.980 73.975 45.120 ;
        RECT 61.250 44.920 61.570 44.980 ;
        RECT 69.070 44.920 69.390 44.980 ;
        RECT 73.685 44.935 73.975 44.980 ;
        RECT 74.220 44.980 77.210 45.120 ;
        RECT 58.490 44.780 58.810 44.840 ;
        RECT 58.965 44.780 59.255 44.825 ;
        RECT 57.200 44.640 58.260 44.780 ;
        RECT 54.350 44.440 54.670 44.500 ;
        RECT 51.245 44.300 54.670 44.440 ;
        RECT 41.010 43.960 42.620 44.100 ;
        RECT 41.010 43.900 41.330 43.960 ;
        RECT 42.850 43.900 43.170 44.160 ;
        RECT 46.070 43.900 46.390 44.160 ;
        RECT 47.450 44.100 47.770 44.160 ;
        RECT 51.245 44.100 51.385 44.300 ;
        RECT 54.350 44.240 54.670 44.300 ;
        RECT 55.270 44.440 55.590 44.500 ;
        RECT 56.740 44.440 56.880 44.595 ;
        RECT 55.270 44.300 56.880 44.440 ;
        RECT 58.120 44.440 58.260 44.640 ;
        RECT 58.490 44.640 59.255 44.780 ;
        RECT 58.490 44.580 58.810 44.640 ;
        RECT 58.965 44.595 59.255 44.640 ;
        RECT 60.330 44.580 60.650 44.840 ;
        RECT 63.550 44.780 63.870 44.840 ;
        RECT 69.545 44.780 69.835 44.825 ;
        RECT 69.990 44.780 70.310 44.840 ;
        RECT 63.550 44.640 69.300 44.780 ;
        RECT 63.550 44.580 63.870 44.640 ;
        RECT 59.870 44.440 60.190 44.500 ;
        RECT 62.630 44.440 62.950 44.500 ;
        RECT 58.120 44.300 60.190 44.440 ;
        RECT 55.270 44.240 55.590 44.300 ;
        RECT 59.870 44.240 60.190 44.300 ;
        RECT 60.420 44.300 62.950 44.440 ;
        RECT 69.160 44.440 69.300 44.640 ;
        RECT 69.545 44.640 70.310 44.780 ;
        RECT 69.545 44.595 69.835 44.640 ;
        RECT 69.990 44.580 70.310 44.640 ;
        RECT 70.925 44.595 71.215 44.825 ;
        RECT 71.830 44.780 72.150 44.840 ;
        RECT 73.225 44.780 73.515 44.825 ;
        RECT 74.220 44.780 74.360 44.980 ;
        RECT 76.890 44.920 77.210 44.980 ;
        RECT 71.830 44.640 74.360 44.780 ;
        RECT 71.000 44.440 71.140 44.595 ;
        RECT 71.830 44.580 72.150 44.640 ;
        RECT 73.225 44.595 73.515 44.640 ;
        RECT 75.050 44.580 75.370 44.840 ;
        RECT 69.160 44.300 71.140 44.440 ;
        RECT 47.450 43.960 51.385 44.100 ;
        RECT 51.590 44.100 51.910 44.160 ;
        RECT 58.505 44.100 58.795 44.145 ;
        RECT 60.420 44.100 60.560 44.300 ;
        RECT 62.630 44.240 62.950 44.300 ;
        RECT 51.590 43.960 60.560 44.100 ;
        RECT 47.450 43.900 47.770 43.960 ;
        RECT 51.590 43.900 51.910 43.960 ;
        RECT 58.505 43.915 58.795 43.960 ;
        RECT 5.520 43.280 76.820 43.760 ;
        RECT 9.285 43.080 9.575 43.125 ;
        RECT 10.190 43.080 10.510 43.140 ;
        RECT 9.285 42.940 10.510 43.080 ;
        RECT 9.285 42.895 9.575 42.940 ;
        RECT 10.190 42.880 10.510 42.940 ;
        RECT 11.110 42.880 11.430 43.140 ;
        RECT 16.645 43.080 16.935 43.125 ;
        RECT 18.010 43.080 18.330 43.140 ;
        RECT 16.645 42.940 18.330 43.080 ;
        RECT 16.645 42.895 16.935 42.940 ;
        RECT 18.010 42.880 18.330 42.940 ;
        RECT 18.930 43.080 19.250 43.140 ;
        RECT 23.085 43.080 23.375 43.125 ;
        RECT 18.930 42.940 23.375 43.080 ;
        RECT 18.930 42.880 19.250 42.940 ;
        RECT 23.085 42.895 23.375 42.940 ;
        RECT 23.990 43.080 24.310 43.140 ;
        RECT 25.830 43.080 26.150 43.140 ;
        RECT 23.990 42.940 26.150 43.080 ;
        RECT 23.990 42.880 24.310 42.940 ;
        RECT 25.830 42.880 26.150 42.940 ;
        RECT 26.290 42.880 26.610 43.140 ;
        RECT 31.350 43.080 31.670 43.140 ;
        RECT 32.285 43.080 32.575 43.125 ;
        RECT 31.350 42.940 32.575 43.080 ;
        RECT 31.350 42.880 31.670 42.940 ;
        RECT 32.285 42.895 32.575 42.940 ;
        RECT 34.125 43.080 34.415 43.125 ;
        RECT 34.570 43.080 34.890 43.140 ;
        RECT 44.230 43.080 44.550 43.140 ;
        RECT 34.125 42.940 34.890 43.080 ;
        RECT 34.125 42.895 34.415 42.940 ;
        RECT 34.570 42.880 34.890 42.940 ;
        RECT 35.580 42.940 44.550 43.080 ;
        RECT 10.650 42.740 10.970 42.800 ;
        RECT 20.770 42.740 21.090 42.800 ;
        RECT 24.450 42.740 24.770 42.800 ;
        RECT 33.205 42.740 33.495 42.785 ;
        RECT 35.580 42.740 35.720 42.940 ;
        RECT 44.230 42.880 44.550 42.940 ;
        RECT 45.610 43.080 45.930 43.140 ;
        RECT 49.765 43.080 50.055 43.125 ;
        RECT 50.210 43.080 50.530 43.140 ;
        RECT 45.610 42.940 50.530 43.080 ;
        RECT 45.610 42.880 45.930 42.940 ;
        RECT 49.765 42.895 50.055 42.940 ;
        RECT 50.210 42.880 50.530 42.940 ;
        RECT 51.605 43.080 51.895 43.125 ;
        RECT 52.970 43.080 53.290 43.140 ;
        RECT 51.605 42.940 53.290 43.080 ;
        RECT 51.605 42.895 51.895 42.940 ;
        RECT 52.970 42.880 53.290 42.940 ;
        RECT 54.350 42.880 54.670 43.140 ;
        RECT 58.950 43.080 59.270 43.140 ;
        RECT 55.820 42.940 59.270 43.080 ;
        RECT 10.650 42.600 20.540 42.740 ;
        RECT 10.650 42.540 10.970 42.600 ;
        RECT 16.170 42.200 16.490 42.460 ;
        RECT 17.550 42.200 17.870 42.460 ;
        RECT 18.930 42.200 19.250 42.460 ;
        RECT 19.850 42.200 20.170 42.460 ;
        RECT 20.400 42.445 20.540 42.600 ;
        RECT 20.770 42.600 24.770 42.740 ;
        RECT 20.770 42.540 21.090 42.600 ;
        RECT 24.450 42.540 24.770 42.600 ;
        RECT 25.460 42.600 33.495 42.740 ;
        RECT 20.325 42.215 20.615 42.445 ;
        RECT 21.690 42.200 22.010 42.460 ;
        RECT 22.165 42.400 22.455 42.445 ;
        RECT 23.990 42.400 24.310 42.460 ;
        RECT 22.165 42.260 24.310 42.400 ;
        RECT 22.165 42.215 22.455 42.260 ;
        RECT 23.990 42.200 24.310 42.260 ;
        RECT 11.570 41.860 11.890 42.120 ;
        RECT 12.030 41.860 12.350 42.120 ;
        RECT 25.460 42.060 25.600 42.600 ;
        RECT 33.205 42.555 33.495 42.600 ;
        RECT 34.665 42.600 35.720 42.740 ;
        RECT 35.965 42.740 36.255 42.785 ;
        RECT 40.090 42.740 40.410 42.800 ;
        RECT 35.965 42.600 40.410 42.740 ;
        RECT 25.845 42.400 26.135 42.445 ;
        RECT 30.890 42.400 31.210 42.460 ;
        RECT 25.845 42.260 31.210 42.400 ;
        RECT 25.845 42.215 26.135 42.260 ;
        RECT 30.890 42.200 31.210 42.260 ;
        RECT 31.810 42.200 32.130 42.460 ;
        RECT 34.665 42.400 34.805 42.600 ;
        RECT 35.965 42.555 36.255 42.600 ;
        RECT 40.090 42.540 40.410 42.600 ;
        RECT 40.550 42.540 40.870 42.800 ;
        RECT 41.470 42.740 41.790 42.800 ;
        RECT 54.440 42.740 54.580 42.880 ;
        RECT 54.825 42.740 55.115 42.785 ;
        RECT 41.470 42.600 49.060 42.740 ;
        RECT 54.440 42.600 55.115 42.740 ;
        RECT 41.470 42.540 41.790 42.600 ;
        RECT 33.280 42.260 34.805 42.400 ;
        RECT 35.045 42.400 35.335 42.445 ;
        RECT 35.490 42.400 35.810 42.460 ;
        RECT 35.045 42.260 35.810 42.400 ;
        RECT 17.640 41.920 25.600 42.060 ;
        RECT 17.640 41.765 17.780 41.920 ;
        RECT 26.750 41.860 27.070 42.120 ;
        RECT 17.565 41.535 17.855 41.765 ;
        RECT 20.785 41.720 21.075 41.765 ;
        RECT 24.005 41.720 24.295 41.765 ;
        RECT 20.785 41.580 24.295 41.720 ;
        RECT 20.785 41.535 21.075 41.580 ;
        RECT 24.005 41.535 24.295 41.580 ;
        RECT 24.450 41.720 24.770 41.780 ;
        RECT 26.840 41.720 26.980 41.860 ;
        RECT 33.280 41.765 33.420 42.260 ;
        RECT 35.045 42.215 35.335 42.260 ;
        RECT 35.490 42.200 35.810 42.260 ;
        RECT 36.410 42.200 36.730 42.460 ;
        RECT 39.645 42.215 39.935 42.445 ;
        RECT 39.720 42.060 39.860 42.215 ;
        RECT 41.010 42.200 41.330 42.460 ;
        RECT 41.930 42.400 42.250 42.460 ;
        RECT 42.405 42.400 42.695 42.445 ;
        RECT 41.930 42.260 42.695 42.400 ;
        RECT 41.930 42.200 42.250 42.260 ;
        RECT 42.405 42.215 42.695 42.260 ;
        RECT 43.310 42.200 43.630 42.460 ;
        RECT 43.785 42.400 44.075 42.445 ;
        RECT 46.545 42.400 46.835 42.445 ;
        RECT 43.785 42.260 46.835 42.400 ;
        RECT 43.785 42.215 44.075 42.260 ;
        RECT 46.545 42.215 46.835 42.260 ;
        RECT 46.990 42.400 47.310 42.460 ;
        RECT 47.465 42.400 47.755 42.445 ;
        RECT 46.990 42.260 47.755 42.400 ;
        RECT 46.990 42.200 47.310 42.260 ;
        RECT 47.465 42.215 47.755 42.260 ;
        RECT 47.925 42.400 48.215 42.445 ;
        RECT 48.370 42.400 48.690 42.460 ;
        RECT 47.925 42.260 48.690 42.400 ;
        RECT 47.925 42.215 48.215 42.260 ;
        RECT 48.370 42.200 48.690 42.260 ;
        RECT 39.720 41.920 42.620 42.060 ;
        RECT 24.450 41.580 26.980 41.720 ;
        RECT 24.450 41.520 24.770 41.580 ;
        RECT 33.205 41.535 33.495 41.765 ;
        RECT 39.170 41.520 39.490 41.780 ;
        RECT 39.630 41.520 39.950 41.780 ;
        RECT 42.480 41.765 42.620 41.920 ;
        RECT 42.405 41.535 42.695 41.765 ;
        RECT 48.920 41.720 49.060 42.600 ;
        RECT 54.825 42.555 55.115 42.600 ;
        RECT 55.285 42.740 55.575 42.785 ;
        RECT 55.820 42.740 55.960 42.940 ;
        RECT 58.950 42.880 59.270 42.940 ;
        RECT 59.410 43.080 59.730 43.140 ;
        RECT 59.410 42.940 62.170 43.080 ;
        RECT 59.410 42.880 59.730 42.940 ;
        RECT 59.870 42.740 60.190 42.800 ;
        RECT 55.285 42.600 55.960 42.740 ;
        RECT 56.280 42.600 60.190 42.740 ;
        RECT 62.030 42.740 62.170 42.940 ;
        RECT 65.390 42.880 65.710 43.140 ;
        RECT 70.450 43.080 70.770 43.140 ;
        RECT 72.765 43.080 73.055 43.125 ;
        RECT 70.450 42.940 73.055 43.080 ;
        RECT 70.450 42.880 70.770 42.940 ;
        RECT 72.765 42.895 73.055 42.940 ;
        RECT 62.030 42.600 65.160 42.740 ;
        RECT 55.285 42.555 55.575 42.600 ;
        RECT 50.685 42.400 50.975 42.445 ;
        RECT 51.590 42.400 51.910 42.460 ;
        RECT 50.685 42.260 51.910 42.400 ;
        RECT 50.685 42.215 50.975 42.260 ;
        RECT 51.590 42.200 51.910 42.260 ;
        RECT 52.065 42.215 52.355 42.445 ;
        RECT 52.970 42.400 53.290 42.460 ;
        RECT 56.280 42.445 56.420 42.600 ;
        RECT 59.870 42.540 60.190 42.600 ;
        RECT 54.135 42.400 54.425 42.445 ;
        RECT 52.970 42.260 54.425 42.400 ;
        RECT 52.140 42.060 52.280 42.215 ;
        RECT 52.970 42.200 53.290 42.260 ;
        RECT 54.135 42.215 54.425 42.260 ;
        RECT 56.200 42.215 56.490 42.445 ;
        RECT 56.650 42.200 56.970 42.460 ;
        RECT 57.570 42.400 57.890 42.460 ;
        RECT 58.490 42.400 58.810 42.460 ;
        RECT 57.570 42.260 58.810 42.400 ;
        RECT 57.570 42.200 57.890 42.260 ;
        RECT 58.490 42.200 58.810 42.260 ;
        RECT 59.410 42.200 59.730 42.460 ;
        RECT 60.805 42.400 61.095 42.445 ;
        RECT 61.250 42.400 61.570 42.460 ;
        RECT 60.805 42.260 61.570 42.400 ;
        RECT 60.805 42.215 61.095 42.260 ;
        RECT 61.250 42.200 61.570 42.260 ;
        RECT 61.710 42.200 62.030 42.460 ;
        RECT 63.180 42.445 63.320 42.600 ;
        RECT 63.105 42.215 63.395 42.445 ;
        RECT 64.470 42.200 64.790 42.460 ;
        RECT 65.020 42.400 65.160 42.600 ;
        RECT 66.310 42.540 66.630 42.800 ;
        RECT 69.070 42.400 69.390 42.460 ;
        RECT 71.830 42.400 72.150 42.460 ;
        RECT 65.020 42.260 72.150 42.400 ;
        RECT 69.070 42.200 69.390 42.260 ;
        RECT 71.830 42.200 72.150 42.260 ;
        RECT 58.030 42.060 58.350 42.120 ;
        RECT 52.140 41.920 58.350 42.060 ;
        RECT 58.030 41.860 58.350 41.920 ;
        RECT 60.345 42.060 60.635 42.105 ;
        RECT 70.450 42.060 70.770 42.120 ;
        RECT 60.345 41.920 70.770 42.060 ;
        RECT 60.345 41.875 60.635 41.920 ;
        RECT 70.450 41.860 70.770 41.920 ;
        RECT 52.985 41.720 53.275 41.765 ;
        RECT 71.370 41.720 71.690 41.780 ;
        RECT 42.940 41.580 48.370 41.720 ;
        RECT 48.920 41.580 52.740 41.720 ;
        RECT 21.230 41.380 21.550 41.440 ;
        RECT 28.590 41.380 28.910 41.440 ;
        RECT 37.790 41.380 38.110 41.440 ;
        RECT 21.230 41.240 38.110 41.380 ;
        RECT 39.260 41.380 39.400 41.520 ;
        RECT 42.940 41.380 43.080 41.580 ;
        RECT 39.260 41.240 43.080 41.380 ;
        RECT 48.230 41.380 48.370 41.580 ;
        RECT 48.830 41.380 49.150 41.440 ;
        RECT 51.590 41.380 51.910 41.440 ;
        RECT 48.230 41.240 51.910 41.380 ;
        RECT 52.600 41.380 52.740 41.580 ;
        RECT 52.985 41.580 71.690 41.720 ;
        RECT 52.985 41.535 53.275 41.580 ;
        RECT 71.370 41.520 71.690 41.580 ;
        RECT 53.445 41.380 53.735 41.425 ;
        RECT 52.600 41.240 53.735 41.380 ;
        RECT 21.230 41.180 21.550 41.240 ;
        RECT 28.590 41.180 28.910 41.240 ;
        RECT 37.790 41.180 38.110 41.240 ;
        RECT 48.830 41.180 49.150 41.240 ;
        RECT 51.590 41.180 51.910 41.240 ;
        RECT 53.445 41.195 53.735 41.240 ;
        RECT 64.010 41.180 64.330 41.440 ;
        RECT 64.470 41.380 64.790 41.440 ;
        RECT 66.310 41.380 66.630 41.440 ;
        RECT 64.470 41.240 66.630 41.380 ;
        RECT 64.470 41.180 64.790 41.240 ;
        RECT 66.310 41.180 66.630 41.240 ;
        RECT 5.520 40.560 76.820 41.040 ;
        RECT 8.810 40.160 9.130 40.420 ;
        RECT 22.625 40.360 22.915 40.405 ;
        RECT 23.070 40.360 23.390 40.420 ;
        RECT 22.625 40.220 23.390 40.360 ;
        RECT 22.625 40.175 22.915 40.220 ;
        RECT 23.070 40.160 23.390 40.220 ;
        RECT 23.990 40.160 24.310 40.420 ;
        RECT 36.410 40.360 36.730 40.420 ;
        RECT 36.885 40.360 37.175 40.405 ;
        RECT 36.410 40.220 37.175 40.360 ;
        RECT 36.410 40.160 36.730 40.220 ;
        RECT 36.885 40.175 37.175 40.220 ;
        RECT 45.610 40.160 45.930 40.420 ;
        RECT 47.910 40.360 48.230 40.420 ;
        RECT 53.430 40.360 53.750 40.420 ;
        RECT 47.910 40.220 53.750 40.360 ;
        RECT 47.910 40.160 48.230 40.220 ;
        RECT 53.430 40.160 53.750 40.220 ;
        RECT 53.890 40.360 54.210 40.420 ;
        RECT 57.125 40.360 57.415 40.405 ;
        RECT 53.890 40.220 57.415 40.360 ;
        RECT 53.890 40.160 54.210 40.220 ;
        RECT 57.125 40.175 57.415 40.220 ;
        RECT 58.030 40.360 58.350 40.420 ;
        RECT 59.410 40.360 59.730 40.420 ;
        RECT 58.030 40.220 59.730 40.360 ;
        RECT 58.030 40.160 58.350 40.220 ;
        RECT 59.410 40.160 59.730 40.220 ;
        RECT 59.870 40.360 60.190 40.420 ;
        RECT 59.870 40.220 60.560 40.360 ;
        RECT 59.870 40.160 60.190 40.220 ;
        RECT 16.645 39.835 16.935 40.065 ;
        RECT 18.930 40.020 19.250 40.080 ;
        RECT 27.670 40.020 27.990 40.080 ;
        RECT 30.430 40.020 30.750 40.080 ;
        RECT 18.930 39.880 25.140 40.020 ;
        RECT 11.110 39.480 11.430 39.740 ;
        RECT 12.030 39.480 12.350 39.740 ;
        RECT 16.720 39.680 16.860 39.835 ;
        RECT 18.930 39.820 19.250 39.880 ;
        RECT 16.720 39.540 24.680 39.680 ;
        RECT 15.250 39.140 15.570 39.400 ;
        RECT 16.630 39.140 16.950 39.400 ;
        RECT 18.930 39.340 19.250 39.400 ;
        RECT 19.865 39.340 20.155 39.385 ;
        RECT 18.930 39.200 20.155 39.340 ;
        RECT 18.930 39.140 19.250 39.200 ;
        RECT 19.865 39.155 20.155 39.200 ;
        RECT 20.770 39.140 21.090 39.400 ;
        RECT 21.245 39.340 21.535 39.385 ;
        RECT 23.070 39.340 23.390 39.400 ;
        RECT 21.245 39.200 23.390 39.340 ;
        RECT 21.245 39.155 21.535 39.200 ;
        RECT 23.070 39.140 23.390 39.200 ;
        RECT 16.720 39.000 16.860 39.140 ;
        RECT 20.310 39.000 20.630 39.060 ;
        RECT 22.625 39.000 22.915 39.045 ;
        RECT 16.720 38.860 22.915 39.000 ;
        RECT 24.540 39.000 24.680 39.540 ;
        RECT 25.000 39.340 25.140 39.880 ;
        RECT 27.670 39.880 30.750 40.020 ;
        RECT 27.670 39.820 27.990 39.880 ;
        RECT 30.430 39.820 30.750 39.880 ;
        RECT 32.285 40.020 32.575 40.065 ;
        RECT 37.330 40.020 37.650 40.080 ;
        RECT 32.285 39.880 37.650 40.020 ;
        RECT 32.285 39.835 32.575 39.880 ;
        RECT 37.330 39.820 37.650 39.880 ;
        RECT 41.010 40.020 41.330 40.080 ;
        RECT 52.065 40.020 52.355 40.065 ;
        RECT 41.010 39.880 52.355 40.020 ;
        RECT 41.010 39.820 41.330 39.880 ;
        RECT 52.065 39.835 52.355 39.880 ;
        RECT 26.290 39.480 26.610 39.740 ;
        RECT 27.210 39.480 27.530 39.740 ;
        RECT 29.985 39.680 30.275 39.725 ;
        RECT 28.220 39.540 30.275 39.680 ;
        RECT 28.220 39.385 28.360 39.540 ;
        RECT 29.985 39.495 30.275 39.540 ;
        RECT 34.110 39.680 34.430 39.740 ;
        RECT 46.070 39.680 46.390 39.740 ;
        RECT 53.890 39.680 54.210 39.740 ;
        RECT 34.110 39.540 46.390 39.680 ;
        RECT 34.110 39.480 34.430 39.540 ;
        RECT 46.070 39.480 46.390 39.540 ;
        RECT 53.060 39.540 54.210 39.680 ;
        RECT 28.145 39.340 28.435 39.385 ;
        RECT 25.000 39.200 28.435 39.340 ;
        RECT 28.145 39.155 28.435 39.200 ;
        RECT 28.590 39.340 28.910 39.400 ;
        RECT 29.525 39.340 29.815 39.385 ;
        RECT 28.590 39.200 29.815 39.340 ;
        RECT 28.590 39.140 28.910 39.200 ;
        RECT 29.525 39.155 29.815 39.200 ;
        RECT 30.445 39.340 30.735 39.385 ;
        RECT 30.890 39.340 31.210 39.400 ;
        RECT 30.445 39.200 31.210 39.340 ;
        RECT 30.445 39.155 30.735 39.200 ;
        RECT 30.890 39.140 31.210 39.200 ;
        RECT 31.350 39.340 31.670 39.400 ;
        RECT 33.205 39.340 33.495 39.385 ;
        RECT 31.350 39.200 33.495 39.340 ;
        RECT 31.350 39.140 31.670 39.200 ;
        RECT 32.285 39.000 32.575 39.045 ;
        RECT 24.540 38.860 32.575 39.000 ;
        RECT 32.820 39.000 32.960 39.200 ;
        RECT 33.205 39.155 33.495 39.200 ;
        RECT 33.665 39.340 33.955 39.385 ;
        RECT 34.570 39.340 34.890 39.400 ;
        RECT 33.665 39.200 34.890 39.340 ;
        RECT 33.665 39.155 33.955 39.200 ;
        RECT 34.570 39.140 34.890 39.200 ;
        RECT 36.425 39.155 36.715 39.385 ;
        RECT 37.345 39.340 37.635 39.385 ;
        RECT 37.790 39.340 38.110 39.400 ;
        RECT 37.345 39.200 38.110 39.340 ;
        RECT 37.345 39.155 37.635 39.200 ;
        RECT 36.500 39.000 36.640 39.155 ;
        RECT 37.790 39.140 38.110 39.200 ;
        RECT 47.450 39.140 47.770 39.400 ;
        RECT 53.060 39.385 53.200 39.540 ;
        RECT 53.890 39.480 54.210 39.540 ;
        RECT 55.270 39.680 55.590 39.740 ;
        RECT 58.965 39.680 59.255 39.725 ;
        RECT 59.870 39.680 60.190 39.740 ;
        RECT 55.270 39.540 60.190 39.680 ;
        RECT 60.420 39.680 60.560 40.220 ;
        RECT 61.710 40.160 62.030 40.420 ;
        RECT 63.105 40.360 63.395 40.405 ;
        RECT 64.010 40.360 64.330 40.420 ;
        RECT 63.105 40.220 64.330 40.360 ;
        RECT 63.105 40.175 63.395 40.220 ;
        RECT 64.010 40.160 64.330 40.220 ;
        RECT 68.610 40.360 68.930 40.420 ;
        RECT 70.925 40.360 71.215 40.405 ;
        RECT 68.610 40.220 71.215 40.360 ;
        RECT 68.610 40.160 68.930 40.220 ;
        RECT 70.925 40.175 71.215 40.220 ;
        RECT 61.265 40.020 61.555 40.065 ;
        RECT 61.800 40.020 61.940 40.160 ;
        RECT 62.630 40.020 62.950 40.080 ;
        RECT 61.265 39.880 62.400 40.020 ;
        RECT 61.265 39.835 61.555 39.880 ;
        RECT 60.420 39.540 61.480 39.680 ;
        RECT 55.270 39.480 55.590 39.540 ;
        RECT 58.965 39.495 59.255 39.540 ;
        RECT 59.870 39.480 60.190 39.540 ;
        RECT 61.340 39.400 61.480 39.540 ;
        RECT 52.985 39.155 53.275 39.385 ;
        RECT 53.445 39.155 53.735 39.385 ;
        RECT 54.365 39.155 54.655 39.385 ;
        RECT 54.825 39.340 55.115 39.385 ;
        RECT 57.110 39.340 57.430 39.400 ;
        RECT 54.825 39.200 57.430 39.340 ;
        RECT 54.825 39.155 55.115 39.200 ;
        RECT 32.820 38.860 36.640 39.000 ;
        RECT 20.310 38.800 20.630 38.860 ;
        RECT 22.625 38.815 22.915 38.860 ;
        RECT 32.285 38.815 32.575 38.860 ;
        RECT 8.810 38.660 9.130 38.720 ;
        RECT 10.665 38.660 10.955 38.705 ;
        RECT 11.570 38.660 11.890 38.720 ;
        RECT 8.810 38.520 11.890 38.660 ;
        RECT 8.810 38.460 9.130 38.520 ;
        RECT 10.665 38.475 10.955 38.520 ;
        RECT 11.570 38.460 11.890 38.520 ;
        RECT 15.725 38.660 16.015 38.705 ;
        RECT 18.945 38.660 19.235 38.705 ;
        RECT 21.705 38.660 21.995 38.705 ;
        RECT 15.725 38.520 21.995 38.660 ;
        RECT 15.725 38.475 16.015 38.520 ;
        RECT 18.945 38.475 19.235 38.520 ;
        RECT 21.705 38.475 21.995 38.520 ;
        RECT 25.845 38.660 26.135 38.705 ;
        RECT 27.670 38.660 27.990 38.720 ;
        RECT 25.845 38.520 27.990 38.660 ;
        RECT 25.845 38.475 26.135 38.520 ;
        RECT 27.670 38.460 27.990 38.520 ;
        RECT 28.605 38.660 28.895 38.705 ;
        RECT 33.190 38.660 33.510 38.720 ;
        RECT 28.605 38.520 33.510 38.660 ;
        RECT 36.500 38.660 36.640 38.860 ;
        RECT 49.290 39.000 49.610 39.060 ;
        RECT 50.670 39.000 50.990 39.060 ;
        RECT 53.520 39.000 53.660 39.155 ;
        RECT 49.290 38.860 53.660 39.000 ;
        RECT 54.440 39.000 54.580 39.155 ;
        RECT 57.110 39.140 57.430 39.200 ;
        RECT 58.030 39.140 58.350 39.400 ;
        RECT 59.425 39.340 59.715 39.385 ;
        RECT 58.580 39.200 59.715 39.340 ;
        RECT 58.580 39.000 58.720 39.200 ;
        RECT 59.425 39.155 59.715 39.200 ;
        RECT 60.330 39.140 60.650 39.400 ;
        RECT 60.805 39.155 61.095 39.385 ;
        RECT 61.250 39.340 61.570 39.400 ;
        RECT 61.725 39.340 62.015 39.385 ;
        RECT 61.250 39.200 62.015 39.340 ;
        RECT 54.440 38.860 58.720 39.000 ;
        RECT 60.880 39.000 61.020 39.155 ;
        RECT 61.250 39.140 61.570 39.200 ;
        RECT 61.725 39.155 62.015 39.200 ;
        RECT 62.260 39.000 62.400 39.880 ;
        RECT 62.630 39.880 64.700 40.020 ;
        RECT 62.630 39.820 62.950 39.880 ;
        RECT 64.010 39.480 64.330 39.740 ;
        RECT 64.560 39.725 64.700 39.880 ;
        RECT 64.485 39.495 64.775 39.725 ;
        RECT 65.405 39.680 65.695 39.725 ;
        RECT 74.130 39.680 74.450 39.740 ;
        RECT 65.405 39.540 74.450 39.680 ;
        RECT 65.405 39.495 65.695 39.540 ;
        RECT 74.130 39.480 74.450 39.540 ;
        RECT 62.645 39.340 62.935 39.385 ;
        RECT 63.090 39.340 63.410 39.400 ;
        RECT 62.645 39.200 63.410 39.340 ;
        RECT 62.645 39.155 62.935 39.200 ;
        RECT 63.090 39.140 63.410 39.200 ;
        RECT 64.945 39.340 65.235 39.385 ;
        RECT 66.310 39.340 66.630 39.400 ;
        RECT 64.945 39.200 66.630 39.340 ;
        RECT 64.945 39.155 65.235 39.200 ;
        RECT 66.310 39.140 66.630 39.200 ;
        RECT 66.770 39.140 67.090 39.400 ;
        RECT 69.085 39.340 69.375 39.385 ;
        RECT 70.910 39.340 71.230 39.400 ;
        RECT 69.085 39.200 71.230 39.340 ;
        RECT 69.085 39.155 69.375 39.200 ;
        RECT 70.910 39.140 71.230 39.200 ;
        RECT 71.385 39.340 71.675 39.385 ;
        RECT 71.830 39.340 72.150 39.400 ;
        RECT 71.385 39.200 72.150 39.340 ;
        RECT 71.385 39.155 71.675 39.200 ;
        RECT 71.830 39.140 72.150 39.200 ;
        RECT 72.750 39.140 73.070 39.400 ;
        RECT 65.390 39.000 65.710 39.060 ;
        RECT 60.880 38.860 61.940 39.000 ;
        RECT 62.260 38.860 65.710 39.000 ;
        RECT 49.290 38.800 49.610 38.860 ;
        RECT 50.670 38.800 50.990 38.860 ;
        RECT 61.800 38.720 61.940 38.860 ;
        RECT 65.390 38.800 65.710 38.860 ;
        RECT 36.870 38.660 37.190 38.720 ;
        RECT 36.500 38.520 37.190 38.660 ;
        RECT 28.605 38.475 28.895 38.520 ;
        RECT 33.190 38.460 33.510 38.520 ;
        RECT 36.870 38.460 37.190 38.520 ;
        RECT 42.390 38.660 42.710 38.720 ;
        RECT 44.705 38.660 44.995 38.705 ;
        RECT 42.390 38.520 44.995 38.660 ;
        RECT 42.390 38.460 42.710 38.520 ;
        RECT 44.705 38.475 44.995 38.520 ;
        RECT 61.710 38.460 62.030 38.720 ;
        RECT 5.520 37.840 76.820 38.320 ;
        RECT 9.730 37.640 10.050 37.700 ;
        RECT 12.045 37.640 12.335 37.685 ;
        RECT 15.725 37.640 16.015 37.685 ;
        RECT 9.730 37.500 16.015 37.640 ;
        RECT 9.730 37.440 10.050 37.500 ;
        RECT 12.045 37.455 12.335 37.500 ;
        RECT 15.725 37.455 16.015 37.500 ;
        RECT 20.770 37.640 21.090 37.700 ;
        RECT 27.210 37.640 27.530 37.700 ;
        RECT 20.770 37.500 27.530 37.640 ;
        RECT 20.770 37.440 21.090 37.500 ;
        RECT 27.210 37.440 27.530 37.500 ;
        RECT 32.270 37.640 32.590 37.700 ;
        RECT 34.110 37.640 34.430 37.700 ;
        RECT 32.270 37.500 34.430 37.640 ;
        RECT 32.270 37.440 32.590 37.500 ;
        RECT 34.110 37.440 34.430 37.500 ;
        RECT 35.030 37.440 35.350 37.700 ;
        RECT 35.950 37.440 36.270 37.700 ;
        RECT 40.090 37.640 40.410 37.700 ;
        RECT 40.565 37.640 40.855 37.685 ;
        RECT 40.090 37.500 40.855 37.640 ;
        RECT 40.090 37.440 40.410 37.500 ;
        RECT 40.565 37.455 40.855 37.500 ;
        RECT 41.470 37.640 41.790 37.700 ;
        RECT 42.850 37.640 43.170 37.700 ;
        RECT 49.305 37.640 49.595 37.685 ;
        RECT 41.470 37.500 49.595 37.640 ;
        RECT 41.470 37.440 41.790 37.500 ;
        RECT 42.850 37.440 43.170 37.500 ;
        RECT 49.305 37.455 49.595 37.500 ;
        RECT 53.445 37.640 53.735 37.685 ;
        RECT 68.610 37.640 68.930 37.700 ;
        RECT 53.445 37.500 68.930 37.640 ;
        RECT 53.445 37.455 53.735 37.500 ;
        RECT 68.610 37.440 68.930 37.500 ;
        RECT 11.585 37.300 11.875 37.345 ;
        RECT 13.410 37.300 13.730 37.360 ;
        RECT 16.185 37.300 16.475 37.345 ;
        RECT 11.585 37.160 16.475 37.300 ;
        RECT 11.585 37.115 11.875 37.160 ;
        RECT 13.410 37.100 13.730 37.160 ;
        RECT 16.185 37.115 16.475 37.160 ;
        RECT 20.310 37.300 20.630 37.360 ;
        RECT 41.930 37.300 42.250 37.360 ;
        RECT 47.465 37.300 47.755 37.345 ;
        RECT 20.310 37.160 43.080 37.300 ;
        RECT 20.310 37.100 20.630 37.160 ;
        RECT 26.290 36.960 26.610 37.020 ;
        RECT 31.825 36.960 32.115 37.005 ;
        RECT 26.290 36.820 32.115 36.960 ;
        RECT 26.290 36.760 26.610 36.820 ;
        RECT 12.030 36.620 12.350 36.680 ;
        RECT 12.965 36.620 13.255 36.665 ;
        RECT 17.105 36.620 17.395 36.665 ;
        RECT 20.770 36.620 21.090 36.680 ;
        RECT 12.030 36.480 21.090 36.620 ;
        RECT 12.030 36.420 12.350 36.480 ;
        RECT 12.965 36.435 13.255 36.480 ;
        RECT 17.105 36.435 17.395 36.480 ;
        RECT 20.770 36.420 21.090 36.480 ;
        RECT 30.980 36.280 31.120 36.820 ;
        RECT 31.825 36.775 32.115 36.820 ;
        RECT 35.950 36.960 36.240 37.005 ;
        RECT 36.870 36.960 37.190 37.020 ;
        RECT 38.340 37.005 38.480 37.160 ;
        RECT 41.930 37.100 42.250 37.160 ;
        RECT 35.950 36.820 37.190 36.960 ;
        RECT 35.950 36.775 36.240 36.820 ;
        RECT 36.870 36.760 37.190 36.820 ;
        RECT 38.265 36.775 38.555 37.005 ;
        RECT 41.470 36.760 41.790 37.020 ;
        RECT 42.390 36.760 42.710 37.020 ;
        RECT 42.940 37.005 43.080 37.160 ;
        RECT 45.240 37.160 47.755 37.300 ;
        RECT 45.240 37.020 45.380 37.160 ;
        RECT 47.465 37.115 47.755 37.160 ;
        RECT 48.370 37.300 48.690 37.360 ;
        RECT 51.590 37.300 51.910 37.360 ;
        RECT 55.285 37.300 55.575 37.345 ;
        RECT 58.045 37.300 58.335 37.345 ;
        RECT 48.370 37.160 50.900 37.300 ;
        RECT 48.370 37.100 48.690 37.160 ;
        RECT 42.865 36.775 43.155 37.005 ;
        RECT 43.310 36.960 43.630 37.020 ;
        RECT 43.785 36.960 44.075 37.005 ;
        RECT 43.310 36.820 44.075 36.960 ;
        RECT 43.310 36.760 43.630 36.820 ;
        RECT 43.785 36.775 44.075 36.820 ;
        RECT 44.690 36.760 45.010 37.020 ;
        RECT 45.150 36.760 45.470 37.020 ;
        RECT 45.610 36.760 45.930 37.020 ;
        RECT 49.750 36.760 50.070 37.020 ;
        RECT 50.760 37.005 50.900 37.160 ;
        RECT 51.590 37.160 55.575 37.300 ;
        RECT 51.590 37.100 51.910 37.160 ;
        RECT 55.285 37.115 55.575 37.160 ;
        RECT 56.280 37.160 58.335 37.300 ;
        RECT 50.685 36.775 50.975 37.005 ;
        RECT 52.525 36.775 52.815 37.005 ;
        RECT 40.090 36.620 40.410 36.680 ;
        RECT 37.420 36.480 40.410 36.620 ;
        RECT 37.420 36.280 37.560 36.480 ;
        RECT 40.090 36.420 40.410 36.480 ;
        RECT 41.930 36.420 42.250 36.680 ;
        RECT 45.700 36.620 45.840 36.760 ;
        RECT 50.225 36.620 50.515 36.665 ;
        RECT 45.700 36.480 50.515 36.620 ;
        RECT 52.600 36.620 52.740 36.775 ;
        RECT 53.890 36.760 54.210 37.020 ;
        RECT 55.730 36.960 56.050 37.020 ;
        RECT 56.280 37.005 56.420 37.160 ;
        RECT 58.045 37.115 58.335 37.160 ;
        RECT 58.950 37.100 59.270 37.360 ;
        RECT 60.790 37.300 61.110 37.360 ;
        RECT 61.725 37.300 62.015 37.345 ;
        RECT 60.790 37.160 62.015 37.300 ;
        RECT 60.790 37.100 61.110 37.160 ;
        RECT 61.725 37.115 62.015 37.160 ;
        RECT 62.170 37.300 62.490 37.360 ;
        RECT 66.325 37.300 66.615 37.345 ;
        RECT 62.170 37.160 66.615 37.300 ;
        RECT 62.170 37.100 62.490 37.160 ;
        RECT 66.325 37.115 66.615 37.160 ;
        RECT 56.205 36.960 56.495 37.005 ;
        RECT 55.730 36.820 56.495 36.960 ;
        RECT 55.730 36.760 56.050 36.820 ;
        RECT 56.205 36.775 56.495 36.820 ;
        RECT 56.665 36.960 56.955 37.005 ;
        RECT 57.570 36.960 57.890 37.020 ;
        RECT 56.665 36.820 57.890 36.960 ;
        RECT 56.665 36.775 56.955 36.820 ;
        RECT 57.570 36.760 57.890 36.820 ;
        RECT 59.410 36.760 59.730 37.020 ;
        RECT 59.870 36.960 60.190 37.020 ;
        RECT 60.345 36.960 60.635 37.005 ;
        RECT 59.870 36.820 60.635 36.960 ;
        RECT 59.870 36.760 60.190 36.820 ;
        RECT 60.345 36.775 60.635 36.820 ;
        RECT 62.645 36.960 62.935 37.005 ;
        RECT 63.550 36.960 63.870 37.020 ;
        RECT 62.645 36.820 63.870 36.960 ;
        RECT 62.645 36.775 62.935 36.820 ;
        RECT 63.550 36.760 63.870 36.820 ;
        RECT 64.025 36.960 64.315 37.005 ;
        RECT 64.470 36.960 64.790 37.020 ;
        RECT 64.025 36.820 64.790 36.960 ;
        RECT 64.025 36.775 64.315 36.820 ;
        RECT 64.470 36.760 64.790 36.820 ;
        RECT 64.945 36.960 65.235 37.005 ;
        RECT 65.850 36.960 66.170 37.020 ;
        RECT 64.945 36.820 66.170 36.960 ;
        RECT 64.945 36.775 65.235 36.820 ;
        RECT 65.850 36.760 66.170 36.820 ;
        RECT 67.690 36.620 68.010 36.680 ;
        RECT 52.600 36.480 68.010 36.620 ;
        RECT 50.225 36.435 50.515 36.480 ;
        RECT 67.690 36.420 68.010 36.480 ;
        RECT 30.980 36.140 37.560 36.280 ;
        RECT 37.805 36.280 38.095 36.325 ;
        RECT 47.005 36.280 47.295 36.325 ;
        RECT 37.805 36.140 47.295 36.280 ;
        RECT 37.805 36.095 38.095 36.140 ;
        RECT 47.005 36.095 47.295 36.140 ;
        RECT 54.825 36.280 55.115 36.325 ;
        RECT 64.010 36.280 64.330 36.340 ;
        RECT 54.825 36.140 64.330 36.280 ;
        RECT 54.825 36.095 55.115 36.140 ;
        RECT 64.010 36.080 64.330 36.140 ;
        RECT 9.730 35.740 10.050 36.000 ;
        RECT 13.870 35.740 14.190 36.000 ;
        RECT 20.310 35.940 20.630 36.000 ;
        RECT 30.890 35.940 31.210 36.000 ;
        RECT 38.250 35.940 38.570 36.000 ;
        RECT 40.550 35.940 40.870 36.000 ;
        RECT 20.310 35.800 40.870 35.940 ;
        RECT 20.310 35.740 20.630 35.800 ;
        RECT 30.890 35.740 31.210 35.800 ;
        RECT 38.250 35.740 38.570 35.800 ;
        RECT 40.550 35.740 40.870 35.800 ;
        RECT 55.285 35.940 55.575 35.985 ;
        RECT 56.650 35.940 56.970 36.000 ;
        RECT 55.285 35.800 56.970 35.940 ;
        RECT 55.285 35.755 55.575 35.800 ;
        RECT 56.650 35.740 56.970 35.800 ;
        RECT 57.110 35.940 57.430 36.000 ;
        RECT 58.965 35.940 59.255 35.985 ;
        RECT 57.110 35.800 59.255 35.940 ;
        RECT 57.110 35.740 57.430 35.800 ;
        RECT 58.965 35.755 59.255 35.800 ;
        RECT 59.870 35.740 60.190 36.000 ;
        RECT 72.750 35.740 73.070 36.000 ;
        RECT 5.520 35.120 76.820 35.600 ;
        RECT 9.285 34.920 9.575 34.965 ;
        RECT 9.730 34.920 10.050 34.980 ;
        RECT 26.305 34.920 26.595 34.965 ;
        RECT 9.285 34.780 10.050 34.920 ;
        RECT 9.285 34.735 9.575 34.780 ;
        RECT 9.730 34.720 10.050 34.780 ;
        RECT 24.540 34.780 26.595 34.920 ;
        RECT 7.890 34.580 8.210 34.640 ;
        RECT 19.390 34.580 19.710 34.640 ;
        RECT 7.890 34.440 19.710 34.580 ;
        RECT 7.890 34.380 8.210 34.440 ;
        RECT 8.900 33.945 9.040 34.440 ;
        RECT 19.390 34.380 19.710 34.440 ;
        RECT 11.585 34.240 11.875 34.285 ;
        RECT 15.250 34.240 15.570 34.300 ;
        RECT 11.585 34.100 15.570 34.240 ;
        RECT 11.585 34.055 11.875 34.100 ;
        RECT 15.250 34.040 15.570 34.100 ;
        RECT 23.990 34.240 24.310 34.300 ;
        RECT 24.540 34.240 24.680 34.780 ;
        RECT 26.305 34.735 26.595 34.780 ;
        RECT 30.905 34.920 31.195 34.965 ;
        RECT 31.810 34.920 32.130 34.980 ;
        RECT 30.905 34.780 32.130 34.920 ;
        RECT 30.905 34.735 31.195 34.780 ;
        RECT 31.810 34.720 32.130 34.780 ;
        RECT 43.310 34.920 43.630 34.980 ;
        RECT 44.705 34.920 44.995 34.965 ;
        RECT 43.310 34.780 44.995 34.920 ;
        RECT 43.310 34.720 43.630 34.780 ;
        RECT 44.705 34.735 44.995 34.780 ;
        RECT 47.005 34.920 47.295 34.965 ;
        RECT 49.750 34.920 50.070 34.980 ;
        RECT 47.005 34.780 50.070 34.920 ;
        RECT 47.005 34.735 47.295 34.780 ;
        RECT 49.750 34.720 50.070 34.780 ;
        RECT 53.890 34.720 54.210 34.980 ;
        RECT 56.665 34.920 56.955 34.965 ;
        RECT 58.490 34.920 58.810 34.980 ;
        RECT 61.265 34.920 61.555 34.965 ;
        RECT 56.665 34.780 58.810 34.920 ;
        RECT 56.665 34.735 56.955 34.780 ;
        RECT 58.490 34.720 58.810 34.780 ;
        RECT 60.880 34.780 61.555 34.920 ;
        RECT 33.190 34.580 33.510 34.640 ;
        RECT 36.870 34.580 37.190 34.640 ;
        RECT 58.950 34.580 59.270 34.640 ;
        RECT 60.880 34.580 61.020 34.780 ;
        RECT 61.265 34.735 61.555 34.780 ;
        RECT 61.710 34.920 62.030 34.980 ;
        RECT 63.565 34.920 63.855 34.965 ;
        RECT 61.710 34.780 63.855 34.920 ;
        RECT 61.710 34.720 62.030 34.780 ;
        RECT 63.565 34.735 63.855 34.780 ;
        RECT 73.210 34.580 73.530 34.640 ;
        RECT 33.190 34.440 37.190 34.580 ;
        RECT 33.190 34.380 33.510 34.440 ;
        RECT 36.870 34.380 37.190 34.440 ;
        RECT 55.820 34.440 61.020 34.580 ;
        RECT 72.380 34.440 73.530 34.580 ;
        RECT 23.990 34.100 24.680 34.240 ;
        RECT 24.925 34.240 25.215 34.285 ;
        RECT 26.290 34.240 26.610 34.300 ;
        RECT 24.925 34.100 26.610 34.240 ;
        RECT 23.990 34.040 24.310 34.100 ;
        RECT 24.925 34.055 25.215 34.100 ;
        RECT 26.290 34.040 26.610 34.100 ;
        RECT 35.030 34.240 35.350 34.300 ;
        RECT 36.410 34.240 36.730 34.300 ;
        RECT 35.030 34.100 36.730 34.240 ;
        RECT 35.030 34.040 35.350 34.100 ;
        RECT 36.410 34.040 36.730 34.100 ;
        RECT 46.070 34.040 46.390 34.300 ;
        RECT 50.685 34.240 50.975 34.285 ;
        RECT 47.080 34.100 49.980 34.240 ;
        RECT 8.825 33.715 9.115 33.945 ;
        RECT 10.190 33.700 10.510 33.960 ;
        RECT 10.665 33.900 10.955 33.945 ;
        RECT 13.870 33.900 14.190 33.960 ;
        RECT 10.665 33.760 14.190 33.900 ;
        RECT 10.665 33.715 10.955 33.760 ;
        RECT 13.870 33.700 14.190 33.760 ;
        RECT 18.930 33.900 19.250 33.960 ;
        RECT 19.865 33.900 20.155 33.945 ;
        RECT 20.310 33.900 20.630 33.960 ;
        RECT 18.930 33.760 20.630 33.900 ;
        RECT 18.930 33.700 19.250 33.760 ;
        RECT 19.865 33.715 20.155 33.760 ;
        RECT 20.310 33.700 20.630 33.760 ;
        RECT 23.530 33.900 23.850 33.960 ;
        RECT 25.845 33.900 26.135 33.945 ;
        RECT 23.530 33.760 26.135 33.900 ;
        RECT 23.530 33.700 23.850 33.760 ;
        RECT 25.845 33.715 26.135 33.760 ;
        RECT 26.765 33.900 27.055 33.945 ;
        RECT 28.130 33.900 28.450 33.960 ;
        RECT 26.765 33.760 28.450 33.900 ;
        RECT 26.765 33.715 27.055 33.760 ;
        RECT 28.130 33.700 28.450 33.760 ;
        RECT 31.810 33.700 32.130 33.960 ;
        RECT 32.270 33.700 32.590 33.960 ;
        RECT 33.190 33.700 33.510 33.960 ;
        RECT 33.665 33.900 33.955 33.945 ;
        RECT 39.170 33.900 39.490 33.960 ;
        RECT 33.665 33.760 39.490 33.900 ;
        RECT 33.665 33.715 33.955 33.760 ;
        RECT 39.170 33.700 39.490 33.760 ;
        RECT 40.090 33.900 40.410 33.960 ;
        RECT 47.080 33.900 47.220 34.100 ;
        RECT 40.090 33.760 47.220 33.900 ;
        RECT 40.090 33.700 40.410 33.760 ;
        RECT 47.450 33.700 47.770 33.960 ;
        RECT 49.840 33.945 49.980 34.100 ;
        RECT 50.685 34.100 55.040 34.240 ;
        RECT 50.685 34.055 50.975 34.100 ;
        RECT 54.900 33.960 55.040 34.100 ;
        RECT 48.845 33.715 49.135 33.945 ;
        RECT 49.765 33.715 50.055 33.945 ;
        RECT 51.145 33.715 51.435 33.945 ;
        RECT 51.590 33.900 51.910 33.960 ;
        RECT 52.065 33.900 52.355 33.945 ;
        RECT 52.510 33.900 52.830 33.960 ;
        RECT 51.590 33.760 52.830 33.900 ;
        RECT 41.010 33.560 41.330 33.620 ;
        RECT 48.920 33.560 49.060 33.715 ;
        RECT 50.210 33.560 50.530 33.620 ;
        RECT 41.010 33.420 50.530 33.560 ;
        RECT 41.010 33.360 41.330 33.420 ;
        RECT 50.210 33.360 50.530 33.420 ;
        RECT 19.405 33.220 19.695 33.265 ;
        RECT 19.850 33.220 20.170 33.280 ;
        RECT 19.405 33.080 20.170 33.220 ;
        RECT 19.405 33.035 19.695 33.080 ;
        RECT 19.850 33.020 20.170 33.080 ;
        RECT 20.310 33.220 20.630 33.280 ;
        RECT 21.705 33.220 21.995 33.265 ;
        RECT 20.310 33.080 21.995 33.220 ;
        RECT 20.310 33.020 20.630 33.080 ;
        RECT 21.705 33.035 21.995 33.080 ;
        RECT 22.610 33.220 22.930 33.280 ;
        RECT 23.545 33.220 23.835 33.265 ;
        RECT 30.890 33.220 31.210 33.280 ;
        RECT 22.610 33.080 31.210 33.220 ;
        RECT 22.610 33.020 22.930 33.080 ;
        RECT 23.545 33.035 23.835 33.080 ;
        RECT 30.890 33.020 31.210 33.080 ;
        RECT 44.230 33.220 44.550 33.280 ;
        RECT 47.450 33.220 47.770 33.280 ;
        RECT 44.230 33.080 47.770 33.220 ;
        RECT 44.230 33.020 44.550 33.080 ;
        RECT 47.450 33.020 47.770 33.080 ;
        RECT 49.750 33.220 50.070 33.280 ;
        RECT 51.220 33.220 51.360 33.715 ;
        RECT 51.590 33.700 51.910 33.760 ;
        RECT 52.065 33.715 52.355 33.760 ;
        RECT 52.510 33.700 52.830 33.760 ;
        RECT 54.810 33.700 55.130 33.960 ;
        RECT 55.820 33.945 55.960 34.440 ;
        RECT 58.950 34.380 59.270 34.440 ;
        RECT 60.790 34.240 61.110 34.300 ;
        RECT 64.025 34.240 64.315 34.285 ;
        RECT 72.380 34.240 72.520 34.440 ;
        RECT 73.210 34.380 73.530 34.440 ;
        RECT 57.200 34.100 64.315 34.240 ;
        RECT 55.745 33.715 56.035 33.945 ;
        RECT 55.285 33.560 55.575 33.605 ;
        RECT 57.200 33.560 57.340 34.100 ;
        RECT 60.790 34.040 61.110 34.100 ;
        RECT 64.025 34.055 64.315 34.100 ;
        RECT 69.160 34.100 72.520 34.240 ;
        RECT 57.585 33.715 57.875 33.945 ;
        RECT 55.285 33.420 57.340 33.560 ;
        RECT 57.660 33.560 57.800 33.715 ;
        RECT 58.030 33.700 58.350 33.960 ;
        RECT 63.565 33.900 63.855 33.945 ;
        RECT 65.390 33.900 65.710 33.960 ;
        RECT 63.565 33.760 65.710 33.900 ;
        RECT 63.565 33.715 63.855 33.760 ;
        RECT 65.390 33.700 65.710 33.760 ;
        RECT 65.865 33.900 66.155 33.945 ;
        RECT 67.230 33.900 67.550 33.960 ;
        RECT 69.160 33.945 69.300 34.100 ;
        RECT 72.750 34.040 73.070 34.300 ;
        RECT 65.865 33.760 67.550 33.900 ;
        RECT 65.865 33.715 66.155 33.760 ;
        RECT 67.230 33.700 67.550 33.760 ;
        RECT 69.085 33.715 69.375 33.945 ;
        RECT 70.450 33.700 70.770 33.960 ;
        RECT 70.910 33.900 71.230 33.960 ;
        RECT 73.225 33.900 73.515 33.945 ;
        RECT 70.910 33.760 73.515 33.900 ;
        RECT 70.910 33.700 71.230 33.760 ;
        RECT 73.225 33.715 73.515 33.760 ;
        RECT 75.050 33.700 75.370 33.960 ;
        RECT 59.870 33.560 60.190 33.620 ;
        RECT 60.345 33.560 60.635 33.605 ;
        RECT 69.990 33.560 70.310 33.620 ;
        RECT 71.845 33.560 72.135 33.605 ;
        RECT 57.660 33.420 59.640 33.560 ;
        RECT 55.285 33.375 55.575 33.420 ;
        RECT 49.750 33.080 51.360 33.220 ;
        RECT 53.430 33.220 53.750 33.280 ;
        RECT 58.030 33.220 58.350 33.280 ;
        RECT 58.965 33.220 59.255 33.265 ;
        RECT 53.430 33.080 59.255 33.220 ;
        RECT 59.500 33.220 59.640 33.420 ;
        RECT 59.870 33.420 60.635 33.560 ;
        RECT 59.870 33.360 60.190 33.420 ;
        RECT 60.345 33.375 60.635 33.420 ;
        RECT 62.260 33.420 66.080 33.560 ;
        RECT 60.790 33.220 61.110 33.280 ;
        RECT 59.500 33.080 61.110 33.220 ;
        RECT 49.750 33.020 50.070 33.080 ;
        RECT 53.430 33.020 53.750 33.080 ;
        RECT 58.030 33.020 58.350 33.080 ;
        RECT 58.965 33.035 59.255 33.080 ;
        RECT 60.790 33.020 61.110 33.080 ;
        RECT 61.250 33.265 61.570 33.280 ;
        RECT 62.260 33.265 62.400 33.420 ;
        RECT 65.940 33.280 66.080 33.420 ;
        RECT 69.990 33.420 72.135 33.560 ;
        RECT 69.990 33.360 70.310 33.420 ;
        RECT 71.845 33.375 72.135 33.420 ;
        RECT 61.250 33.035 61.635 33.265 ;
        RECT 62.185 33.035 62.475 33.265 ;
        RECT 62.630 33.220 62.950 33.280 ;
        RECT 65.405 33.220 65.695 33.265 ;
        RECT 62.630 33.080 65.695 33.220 ;
        RECT 61.250 33.020 61.570 33.035 ;
        RECT 62.630 33.020 62.950 33.080 ;
        RECT 65.405 33.035 65.695 33.080 ;
        RECT 65.850 33.020 66.170 33.280 ;
        RECT 66.785 33.220 67.075 33.265 ;
        RECT 68.150 33.220 68.470 33.280 ;
        RECT 66.785 33.080 68.470 33.220 ;
        RECT 66.785 33.035 67.075 33.080 ;
        RECT 68.150 33.020 68.470 33.080 ;
        RECT 71.385 33.220 71.675 33.265 ;
        RECT 72.290 33.220 72.610 33.280 ;
        RECT 71.385 33.080 72.610 33.220 ;
        RECT 71.385 33.035 71.675 33.080 ;
        RECT 72.290 33.020 72.610 33.080 ;
        RECT 5.520 32.400 76.820 32.880 ;
        RECT 10.665 32.015 10.955 32.245 ;
        RECT 12.030 32.200 12.350 32.260 ;
        RECT 18.470 32.200 18.790 32.260 ;
        RECT 20.785 32.200 21.075 32.245 ;
        RECT 23.070 32.200 23.390 32.260 ;
        RECT 12.030 32.060 20.540 32.200 ;
        RECT 10.740 31.860 10.880 32.015 ;
        RECT 12.030 32.000 12.350 32.060 ;
        RECT 18.470 32.000 18.790 32.060 ;
        RECT 17.105 31.860 17.395 31.905 ;
        RECT 20.400 31.860 20.540 32.060 ;
        RECT 20.785 32.060 23.390 32.200 ;
        RECT 20.785 32.015 21.075 32.060 ;
        RECT 23.070 32.000 23.390 32.060 ;
        RECT 23.545 32.200 23.835 32.245 ;
        RECT 23.990 32.200 24.310 32.260 ;
        RECT 23.545 32.060 24.310 32.200 ;
        RECT 23.545 32.015 23.835 32.060 ;
        RECT 23.990 32.000 24.310 32.060 ;
        RECT 25.830 32.200 26.150 32.260 ;
        RECT 28.590 32.200 28.910 32.260 ;
        RECT 25.830 32.060 28.910 32.200 ;
        RECT 25.830 32.000 26.150 32.060 ;
        RECT 28.590 32.000 28.910 32.060 ;
        RECT 31.825 32.200 32.115 32.245 ;
        RECT 33.190 32.200 33.510 32.260 ;
        RECT 34.110 32.200 34.430 32.260 ;
        RECT 31.825 32.060 33.510 32.200 ;
        RECT 31.825 32.015 32.115 32.060 ;
        RECT 33.190 32.000 33.510 32.060 ;
        RECT 33.740 32.060 34.430 32.200 ;
        RECT 25.370 31.860 25.690 31.920 ;
        RECT 27.225 31.860 27.515 31.905 ;
        RECT 28.145 31.860 28.435 31.905 ;
        RECT 33.740 31.860 33.880 32.060 ;
        RECT 34.110 32.000 34.430 32.060 ;
        RECT 35.120 32.060 38.480 32.200 ;
        RECT 8.440 31.720 10.880 31.860 ;
        RECT 11.200 31.720 18.700 31.860 ;
        RECT 20.400 31.720 26.520 31.860 ;
        RECT 8.440 31.565 8.580 31.720 ;
        RECT 8.365 31.335 8.655 31.565 ;
        RECT 9.285 31.335 9.575 31.565 ;
        RECT 10.650 31.520 10.970 31.580 ;
        RECT 11.200 31.520 11.340 31.720 ;
        RECT 17.105 31.675 17.395 31.720 ;
        RECT 10.650 31.380 11.340 31.520 ;
        RECT 11.585 31.520 11.875 31.565 ;
        RECT 16.645 31.520 16.935 31.565 ;
        RECT 11.585 31.380 16.935 31.520 ;
        RECT 4.670 31.180 4.990 31.240 ;
        RECT 9.360 31.180 9.500 31.335 ;
        RECT 10.650 31.320 10.970 31.380 ;
        RECT 11.585 31.335 11.875 31.380 ;
        RECT 16.645 31.335 16.935 31.380 ;
        RECT 4.670 31.040 9.500 31.180 ;
        RECT 4.670 30.980 4.990 31.040 ;
        RECT 3.750 30.840 4.070 30.900 ;
        RECT 7.445 30.840 7.735 30.885 ;
        RECT 3.750 30.700 7.735 30.840 ;
        RECT 3.750 30.640 4.070 30.700 ;
        RECT 7.445 30.655 7.735 30.700 ;
        RECT 10.190 30.640 10.510 30.900 ;
        RECT 16.720 30.840 16.860 31.335 ;
        RECT 17.550 31.320 17.870 31.580 ;
        RECT 18.025 31.510 18.315 31.565 ;
        RECT 18.560 31.510 18.700 31.720 ;
        RECT 25.370 31.660 25.690 31.720 ;
        RECT 18.025 31.370 18.700 31.510 ;
        RECT 18.025 31.335 18.315 31.370 ;
        RECT 19.390 31.320 19.710 31.580 ;
        RECT 19.865 31.520 20.155 31.565 ;
        RECT 22.610 31.520 22.930 31.580 ;
        RECT 23.085 31.520 23.375 31.565 ;
        RECT 19.865 31.380 21.460 31.520 ;
        RECT 19.865 31.335 20.155 31.380 ;
        RECT 18.485 31.180 18.775 31.225 ;
        RECT 20.310 31.180 20.630 31.240 ;
        RECT 18.485 31.040 20.630 31.180 ;
        RECT 18.485 30.995 18.775 31.040 ;
        RECT 20.310 30.980 20.630 31.040 ;
        RECT 19.850 30.840 20.170 30.900 ;
        RECT 21.320 30.885 21.460 31.380 ;
        RECT 22.610 31.380 23.375 31.520 ;
        RECT 22.610 31.320 22.930 31.380 ;
        RECT 23.085 31.335 23.375 31.380 ;
        RECT 24.910 31.520 25.230 31.580 ;
        RECT 26.380 31.565 26.520 31.720 ;
        RECT 27.225 31.720 33.880 31.860 ;
        RECT 27.225 31.675 27.515 31.720 ;
        RECT 28.145 31.675 28.435 31.720 ;
        RECT 24.910 31.380 26.035 31.520 ;
        RECT 24.910 31.320 25.230 31.380 ;
        RECT 24.005 30.995 24.295 31.225 ;
        RECT 24.450 31.180 24.770 31.240 ;
        RECT 25.385 31.180 25.675 31.225 ;
        RECT 24.450 31.040 25.675 31.180 ;
        RECT 25.895 31.180 26.035 31.380 ;
        RECT 26.305 31.335 26.595 31.565 ;
        RECT 26.750 31.520 27.070 31.580 ;
        RECT 29.065 31.520 29.355 31.565 ;
        RECT 26.750 31.380 29.355 31.520 ;
        RECT 26.750 31.320 27.070 31.380 ;
        RECT 29.065 31.335 29.355 31.380 ;
        RECT 32.270 31.520 32.590 31.580 ;
        RECT 32.745 31.520 33.035 31.565 ;
        RECT 32.270 31.380 33.035 31.520 ;
        RECT 32.270 31.320 32.590 31.380 ;
        RECT 32.745 31.335 33.035 31.380 ;
        RECT 34.645 31.550 34.935 31.595 ;
        RECT 35.120 31.550 35.260 32.060 ;
        RECT 36.755 31.860 37.045 31.905 ;
        RECT 36.755 31.675 37.100 31.860 ;
        RECT 34.645 31.410 35.260 31.550 ;
        RECT 34.645 31.365 34.935 31.410 ;
        RECT 35.490 31.310 35.810 31.570 ;
        RECT 35.965 31.520 36.255 31.565 ;
        RECT 36.410 31.520 36.730 31.530 ;
        RECT 35.965 31.380 36.730 31.520 ;
        RECT 35.965 31.335 36.255 31.380 ;
        RECT 36.410 31.270 36.730 31.380 ;
        RECT 33.190 31.180 33.510 31.240 ;
        RECT 33.665 31.180 33.955 31.225 ;
        RECT 25.895 31.040 33.955 31.180 ;
        RECT 16.720 30.700 20.170 30.840 ;
        RECT 19.850 30.640 20.170 30.700 ;
        RECT 21.245 30.655 21.535 30.885 ;
        RECT 24.080 30.840 24.220 30.995 ;
        RECT 24.450 30.980 24.770 31.040 ;
        RECT 25.385 30.995 25.675 31.040 ;
        RECT 33.190 30.980 33.510 31.040 ;
        RECT 33.665 30.995 33.955 31.040 ;
        RECT 34.110 30.980 34.430 31.240 ;
        RECT 27.210 30.840 27.530 30.900 ;
        RECT 24.080 30.700 27.530 30.840 ;
        RECT 27.210 30.640 27.530 30.700 ;
        RECT 29.985 30.840 30.275 30.885 ;
        RECT 36.960 30.840 37.100 31.675 ;
        RECT 38.340 31.580 38.480 32.060 ;
        RECT 39.170 32.000 39.490 32.260 ;
        RECT 40.090 32.200 40.410 32.260 ;
        RECT 43.785 32.200 44.075 32.245 ;
        RECT 40.090 32.060 44.075 32.200 ;
        RECT 40.090 32.000 40.410 32.060 ;
        RECT 43.785 32.015 44.075 32.060 ;
        RECT 44.245 32.200 44.535 32.245 ;
        RECT 45.150 32.200 45.470 32.260 ;
        RECT 44.245 32.060 45.470 32.200 ;
        RECT 44.245 32.015 44.535 32.060 ;
        RECT 45.150 32.000 45.470 32.060 ;
        RECT 50.670 32.000 50.990 32.260 ;
        RECT 55.285 32.200 55.575 32.245 ;
        RECT 56.190 32.200 56.510 32.260 ;
        RECT 55.285 32.060 56.510 32.200 ;
        RECT 55.285 32.015 55.575 32.060 ;
        RECT 56.190 32.000 56.510 32.060 ;
        RECT 57.570 32.000 57.890 32.260 ;
        RECT 60.330 32.200 60.650 32.260 ;
        RECT 60.805 32.200 61.095 32.245 ;
        RECT 60.330 32.060 61.095 32.200 ;
        RECT 60.330 32.000 60.650 32.060 ;
        RECT 60.805 32.015 61.095 32.060 ;
        RECT 64.945 32.200 65.235 32.245 ;
        RECT 65.390 32.200 65.710 32.260 ;
        RECT 64.945 32.060 65.710 32.200 ;
        RECT 64.945 32.015 65.235 32.060 ;
        RECT 65.390 32.000 65.710 32.060 ;
        RECT 67.230 32.000 67.550 32.260 ;
        RECT 69.070 32.200 69.390 32.260 ;
        RECT 71.845 32.200 72.135 32.245 ;
        RECT 73.670 32.200 73.990 32.260 ;
        RECT 69.070 32.060 73.990 32.200 ;
        RECT 69.070 32.000 69.390 32.060 ;
        RECT 71.845 32.015 72.135 32.060 ;
        RECT 73.670 32.000 73.990 32.060 ;
        RECT 39.630 31.860 39.950 31.920 ;
        RECT 64.470 31.905 64.790 31.920 ;
        RECT 43.325 31.860 43.615 31.905 ;
        RECT 52.525 31.860 52.815 31.905 ;
        RECT 52.985 31.860 53.275 31.905 ;
        RECT 61.565 31.860 61.855 31.905 ;
        RECT 62.645 31.860 62.935 31.905 ;
        RECT 39.630 31.720 43.615 31.860 ;
        RECT 39.630 31.660 39.950 31.720 ;
        RECT 43.325 31.675 43.615 31.720 ;
        RECT 44.320 31.720 51.820 31.860 ;
        RECT 37.345 31.335 37.635 31.565 ;
        RECT 37.805 31.335 38.095 31.565 ;
        RECT 38.250 31.520 38.570 31.580 ;
        RECT 41.010 31.520 41.330 31.580 ;
        RECT 42.865 31.520 43.155 31.565 ;
        RECT 38.250 31.380 43.155 31.520 ;
        RECT 29.985 30.700 37.100 30.840 ;
        RECT 29.985 30.655 30.275 30.700 ;
        RECT 31.350 30.500 31.670 30.560 ;
        RECT 35.490 30.500 35.810 30.560 ;
        RECT 37.420 30.500 37.560 31.335 ;
        RECT 37.880 31.180 38.020 31.335 ;
        RECT 38.250 31.320 38.570 31.380 ;
        RECT 41.010 31.320 41.330 31.380 ;
        RECT 42.865 31.335 43.155 31.380 ;
        RECT 38.710 31.180 39.030 31.240 ;
        RECT 37.880 31.040 39.030 31.180 ;
        RECT 38.710 30.980 39.030 31.040 ;
        RECT 39.630 31.180 39.950 31.240 ;
        RECT 44.320 31.225 44.460 31.720 ;
        RECT 45.165 31.520 45.455 31.565 ;
        RECT 49.290 31.520 49.610 31.580 ;
        RECT 44.780 31.380 49.610 31.520 ;
        RECT 44.245 31.180 44.535 31.225 ;
        RECT 39.630 31.040 44.535 31.180 ;
        RECT 39.630 30.980 39.950 31.040 ;
        RECT 44.245 30.995 44.535 31.040 ;
        RECT 41.010 30.840 41.330 30.900 ;
        RECT 44.780 30.840 44.920 31.380 ;
        RECT 45.165 31.335 45.455 31.380 ;
        RECT 49.290 31.320 49.610 31.380 ;
        RECT 50.210 31.320 50.530 31.580 ;
        RECT 51.130 31.520 51.450 31.580 ;
        RECT 51.680 31.565 51.820 31.720 ;
        RECT 52.525 31.720 61.855 31.860 ;
        RECT 52.525 31.675 52.815 31.720 ;
        RECT 52.985 31.675 53.275 31.720 ;
        RECT 61.565 31.675 61.855 31.720 ;
        RECT 62.030 31.720 62.935 31.860 ;
        RECT 51.605 31.520 51.895 31.565 ;
        RECT 51.130 31.380 51.895 31.520 ;
        RECT 51.130 31.320 51.450 31.380 ;
        RECT 51.605 31.335 51.895 31.380 ;
        RECT 54.350 31.320 54.670 31.580 ;
        RECT 54.900 31.380 58.260 31.520 ;
        RECT 45.610 31.180 45.930 31.240 ;
        RECT 53.905 31.180 54.195 31.225 ;
        RECT 54.900 31.180 55.040 31.380 ;
        RECT 45.610 31.040 55.040 31.180 ;
        RECT 58.120 31.180 58.260 31.380 ;
        RECT 58.490 31.320 58.810 31.580 ;
        RECT 58.950 31.320 59.270 31.580 ;
        RECT 59.870 31.520 60.190 31.580 ;
        RECT 60.345 31.520 60.635 31.565 ;
        RECT 62.030 31.520 62.170 31.720 ;
        RECT 62.645 31.675 62.935 31.720 ;
        RECT 63.105 31.675 63.395 31.905 ;
        RECT 64.185 31.675 64.790 31.905 ;
        RECT 69.545 31.860 69.835 31.905 ;
        RECT 69.545 31.720 75.280 31.860 ;
        RECT 69.545 31.675 69.835 31.720 ;
        RECT 59.870 31.380 62.170 31.520 ;
        RECT 59.870 31.320 60.190 31.380 ;
        RECT 60.345 31.335 60.635 31.380 ;
        RECT 61.250 31.180 61.570 31.240 ;
        RECT 58.120 31.040 61.570 31.180 ;
        RECT 45.610 30.980 45.930 31.040 ;
        RECT 53.905 30.995 54.195 31.040 ;
        RECT 61.250 30.980 61.570 31.040 ;
        RECT 62.170 31.180 62.490 31.240 ;
        RECT 63.180 31.180 63.320 31.675 ;
        RECT 64.470 31.660 64.790 31.675 ;
        RECT 70.910 31.520 71.230 31.580 ;
        RECT 71.385 31.520 71.675 31.565 ;
        RECT 62.170 31.040 63.320 31.180 ;
        RECT 68.240 31.380 71.675 31.520 ;
        RECT 62.170 30.980 62.490 31.040 ;
        RECT 68.240 30.900 68.380 31.380 ;
        RECT 70.910 31.320 71.230 31.380 ;
        RECT 71.385 31.335 71.675 31.380 ;
        RECT 57.110 30.840 57.430 30.900 ;
        RECT 41.010 30.700 44.920 30.840 ;
        RECT 54.440 30.700 57.430 30.840 ;
        RECT 41.010 30.640 41.330 30.700 ;
        RECT 54.440 30.545 54.580 30.700 ;
        RECT 57.110 30.640 57.430 30.700 ;
        RECT 58.950 30.840 59.270 30.900 ;
        RECT 58.950 30.700 61.560 30.840 ;
        RECT 58.950 30.640 59.270 30.700 ;
        RECT 31.350 30.360 37.560 30.500 ;
        RECT 31.350 30.300 31.670 30.360 ;
        RECT 35.490 30.300 35.810 30.360 ;
        RECT 54.365 30.315 54.655 30.545 ;
        RECT 54.810 30.500 55.130 30.560 ;
        RECT 59.885 30.500 60.175 30.545 ;
        RECT 60.330 30.500 60.650 30.560 ;
        RECT 54.810 30.360 60.650 30.500 ;
        RECT 61.420 30.500 61.560 30.700 ;
        RECT 68.150 30.640 68.470 30.900 ;
        RECT 71.920 30.840 72.060 31.720 ;
        RECT 75.140 31.580 75.280 31.720 ;
        RECT 72.305 31.520 72.595 31.565 ;
        RECT 73.210 31.520 73.530 31.580 ;
        RECT 72.305 31.380 73.530 31.520 ;
        RECT 72.305 31.335 72.595 31.380 ;
        RECT 73.210 31.320 73.530 31.380 ;
        RECT 75.050 31.320 75.370 31.580 ;
        RECT 74.130 30.980 74.450 31.240 ;
        RECT 72.290 30.840 72.610 30.900 ;
        RECT 71.920 30.700 72.610 30.840 ;
        RECT 72.290 30.640 72.610 30.700 ;
        RECT 61.725 30.500 62.015 30.545 ;
        RECT 61.420 30.360 62.015 30.500 ;
        RECT 54.810 30.300 55.130 30.360 ;
        RECT 59.885 30.315 60.175 30.360 ;
        RECT 60.330 30.300 60.650 30.360 ;
        RECT 61.725 30.315 62.015 30.360 ;
        RECT 64.010 30.300 64.330 30.560 ;
        RECT 5.520 29.680 76.820 30.160 ;
        RECT 8.810 29.280 9.130 29.540 ;
        RECT 13.410 29.280 13.730 29.540 ;
        RECT 21.245 29.480 21.535 29.525 ;
        RECT 31.350 29.480 31.670 29.540 ;
        RECT 21.245 29.340 31.670 29.480 ;
        RECT 21.245 29.295 21.535 29.340 ;
        RECT 31.350 29.280 31.670 29.340 ;
        RECT 31.810 29.480 32.130 29.540 ;
        RECT 35.965 29.480 36.255 29.525 ;
        RECT 45.610 29.480 45.930 29.540 ;
        RECT 31.810 29.340 45.930 29.480 ;
        RECT 31.810 29.280 32.130 29.340 ;
        RECT 35.965 29.295 36.255 29.340 ;
        RECT 45.610 29.280 45.930 29.340 ;
        RECT 51.145 29.480 51.435 29.525 ;
        RECT 58.490 29.480 58.810 29.540 ;
        RECT 51.145 29.340 58.810 29.480 ;
        RECT 51.145 29.295 51.435 29.340 ;
        RECT 58.490 29.280 58.810 29.340 ;
        RECT 60.330 29.480 60.650 29.540 ;
        RECT 61.265 29.480 61.555 29.525 ;
        RECT 64.010 29.480 64.330 29.540 ;
        RECT 60.330 29.340 64.330 29.480 ;
        RECT 60.330 29.280 60.650 29.340 ;
        RECT 61.265 29.295 61.555 29.340 ;
        RECT 64.010 29.280 64.330 29.340 ;
        RECT 64.930 29.480 65.250 29.540 ;
        RECT 65.405 29.480 65.695 29.525 ;
        RECT 64.930 29.340 65.695 29.480 ;
        RECT 64.930 29.280 65.250 29.340 ;
        RECT 65.405 29.295 65.695 29.340 ;
        RECT 66.770 29.480 67.090 29.540 ;
        RECT 67.245 29.480 67.535 29.525 ;
        RECT 66.770 29.340 67.535 29.480 ;
        RECT 66.770 29.280 67.090 29.340 ;
        RECT 67.245 29.295 67.535 29.340 ;
        RECT 71.370 29.280 71.690 29.540 ;
        RECT 73.225 29.295 73.515 29.525 ;
        RECT 10.190 29.140 10.510 29.200 ;
        RECT 11.585 29.140 11.875 29.185 ;
        RECT 14.330 29.140 14.650 29.200 ;
        RECT 24.910 29.140 25.230 29.200 ;
        RECT 7.980 29.000 14.650 29.140 ;
        RECT 7.980 28.505 8.120 29.000 ;
        RECT 10.190 28.940 10.510 29.000 ;
        RECT 11.585 28.955 11.875 29.000 ;
        RECT 14.330 28.940 14.650 29.000 ;
        RECT 15.325 29.000 25.230 29.140 ;
        RECT 9.285 28.800 9.575 28.845 ;
        RECT 12.030 28.800 12.350 28.860 ;
        RECT 9.285 28.660 12.350 28.800 ;
        RECT 9.285 28.615 9.575 28.660 ;
        RECT 12.030 28.600 12.350 28.660 ;
        RECT 12.965 28.800 13.255 28.845 ;
        RECT 13.410 28.800 13.730 28.860 ;
        RECT 15.325 28.800 15.465 29.000 ;
        RECT 24.910 28.940 25.230 29.000 ;
        RECT 33.190 29.140 33.510 29.200 ;
        RECT 35.045 29.140 35.335 29.185 ;
        RECT 40.090 29.140 40.410 29.200 ;
        RECT 33.190 29.000 35.335 29.140 ;
        RECT 33.190 28.940 33.510 29.000 ;
        RECT 35.045 28.955 35.335 29.000 ;
        RECT 37.880 29.000 40.410 29.140 ;
        RECT 12.965 28.660 15.465 28.800 ;
        RECT 17.550 28.800 17.870 28.860 ;
        RECT 19.405 28.800 19.695 28.845 ;
        RECT 21.230 28.800 21.550 28.860 ;
        RECT 17.550 28.660 37.560 28.800 ;
        RECT 12.965 28.615 13.255 28.660 ;
        RECT 13.410 28.600 13.730 28.660 ;
        RECT 17.550 28.600 17.870 28.660 ;
        RECT 19.405 28.615 19.695 28.660 ;
        RECT 21.230 28.600 21.550 28.660 ;
        RECT 7.905 28.275 8.195 28.505 ;
        RECT 8.365 28.460 8.655 28.505 ;
        RECT 9.745 28.460 10.035 28.505 ;
        RECT 13.870 28.460 14.190 28.520 ;
        RECT 8.365 28.320 14.190 28.460 ;
        RECT 8.365 28.275 8.655 28.320 ;
        RECT 9.745 28.275 10.035 28.320 ;
        RECT 13.870 28.260 14.190 28.320 ;
        RECT 14.330 28.260 14.650 28.520 ;
        RECT 19.850 28.460 20.170 28.520 ;
        RECT 20.325 28.460 20.615 28.505 ;
        RECT 19.850 28.320 20.615 28.460 ;
        RECT 19.850 28.260 20.170 28.320 ;
        RECT 20.325 28.275 20.615 28.320 ;
        RECT 23.530 28.260 23.850 28.520 ;
        RECT 34.125 28.460 34.415 28.505 ;
        RECT 35.030 28.460 35.350 28.520 ;
        RECT 34.125 28.320 35.350 28.460 ;
        RECT 34.125 28.275 34.415 28.320 ;
        RECT 35.030 28.260 35.350 28.320 ;
        RECT 35.490 28.260 35.810 28.520 ;
        RECT 36.885 28.275 37.175 28.505 ;
        RECT 36.960 28.120 37.100 28.275 ;
        RECT 37.420 28.165 37.560 28.660 ;
        RECT 37.880 28.505 38.020 29.000 ;
        RECT 40.090 28.940 40.410 29.000 ;
        RECT 40.550 28.940 40.870 29.200 ;
        RECT 41.485 28.955 41.775 29.185 ;
        RECT 58.030 29.140 58.350 29.200 ;
        RECT 73.300 29.140 73.440 29.295 ;
        RECT 58.030 29.000 73.440 29.140 ;
        RECT 40.180 28.800 40.320 28.940 ;
        RECT 41.560 28.800 41.700 28.955 ;
        RECT 58.030 28.940 58.350 29.000 ;
        RECT 40.180 28.660 41.700 28.800 ;
        RECT 50.210 28.800 50.530 28.860 ;
        RECT 64.470 28.800 64.790 28.860 ;
        RECT 50.210 28.660 52.740 28.800 ;
        RECT 50.210 28.600 50.530 28.660 ;
        RECT 37.805 28.275 38.095 28.505 ;
        RECT 38.250 28.460 38.570 28.520 ;
        RECT 38.725 28.460 39.015 28.505 ;
        RECT 38.250 28.320 39.015 28.460 ;
        RECT 38.250 28.260 38.570 28.320 ;
        RECT 38.725 28.275 39.015 28.320 ;
        RECT 51.130 28.260 51.450 28.520 ;
        RECT 52.600 28.505 52.740 28.660 ;
        RECT 61.420 28.660 65.160 28.800 ;
        RECT 52.525 28.275 52.815 28.505 ;
        RECT 58.490 28.460 58.810 28.520 ;
        RECT 61.420 28.460 61.560 28.660 ;
        RECT 64.470 28.600 64.790 28.660 ;
        RECT 65.020 28.505 65.160 28.660 ;
        RECT 65.850 28.600 66.170 28.860 ;
        RECT 67.690 28.600 68.010 28.860 ;
        RECT 72.750 28.800 73.070 28.860 ;
        RECT 68.700 28.660 73.070 28.800 ;
        RECT 68.700 28.505 68.840 28.660 ;
        RECT 72.750 28.600 73.070 28.660 ;
        RECT 64.025 28.460 64.315 28.505 ;
        RECT 58.490 28.320 61.560 28.460 ;
        RECT 58.490 28.260 58.810 28.320 ;
        RECT 21.780 27.980 37.100 28.120 ;
        RECT 37.345 28.120 37.635 28.165 ;
        RECT 39.185 28.120 39.475 28.165 ;
        RECT 41.010 28.120 41.330 28.180 ;
        RECT 50.670 28.120 50.990 28.180 ;
        RECT 52.065 28.120 52.355 28.165 ;
        RECT 37.345 27.980 39.860 28.120 ;
        RECT 5.130 27.780 5.450 27.840 ;
        RECT 12.045 27.780 12.335 27.825 ;
        RECT 21.780 27.780 21.920 27.980 ;
        RECT 35.580 27.840 35.720 27.980 ;
        RECT 37.345 27.935 37.635 27.980 ;
        RECT 39.185 27.935 39.475 27.980 ;
        RECT 5.130 27.640 21.920 27.780 ;
        RECT 22.150 27.780 22.470 27.840 ;
        RECT 22.625 27.780 22.915 27.825 ;
        RECT 25.830 27.780 26.150 27.840 ;
        RECT 22.150 27.640 26.150 27.780 ;
        RECT 5.130 27.580 5.450 27.640 ;
        RECT 12.045 27.595 12.335 27.640 ;
        RECT 22.150 27.580 22.470 27.640 ;
        RECT 22.625 27.595 22.915 27.640 ;
        RECT 25.830 27.580 26.150 27.640 ;
        RECT 32.270 27.780 32.590 27.840 ;
        RECT 33.205 27.780 33.495 27.825 ;
        RECT 32.270 27.640 33.495 27.780 ;
        RECT 32.270 27.580 32.590 27.640 ;
        RECT 33.205 27.595 33.495 27.640 ;
        RECT 35.490 27.580 35.810 27.840 ;
        RECT 39.720 27.780 39.860 27.980 ;
        RECT 41.010 27.980 50.440 28.120 ;
        RECT 41.010 27.920 41.330 27.980 ;
        RECT 49.750 27.780 50.070 27.840 ;
        RECT 39.720 27.640 50.070 27.780 ;
        RECT 50.300 27.780 50.440 27.980 ;
        RECT 50.670 27.980 52.355 28.120 ;
        RECT 50.670 27.920 50.990 27.980 ;
        RECT 52.065 27.935 52.355 27.980 ;
        RECT 57.110 28.120 57.430 28.180 ;
        RECT 61.420 28.165 61.560 28.320 ;
        RECT 61.800 28.320 64.315 28.460 ;
        RECT 60.345 28.120 60.635 28.165 ;
        RECT 57.110 27.980 60.635 28.120 ;
        RECT 57.110 27.920 57.430 27.980 ;
        RECT 60.345 27.935 60.635 27.980 ;
        RECT 61.345 27.935 61.635 28.165 ;
        RECT 51.590 27.780 51.910 27.840 ;
        RECT 50.300 27.640 51.910 27.780 ;
        RECT 49.750 27.580 50.070 27.640 ;
        RECT 51.590 27.580 51.910 27.640 ;
        RECT 55.270 27.780 55.590 27.840 ;
        RECT 58.490 27.780 58.810 27.840 ;
        RECT 55.270 27.640 58.810 27.780 ;
        RECT 55.270 27.580 55.590 27.640 ;
        RECT 58.490 27.580 58.810 27.640 ;
        RECT 59.870 27.780 60.190 27.840 ;
        RECT 61.800 27.780 61.940 28.320 ;
        RECT 64.025 28.275 64.315 28.320 ;
        RECT 64.945 28.275 65.235 28.505 ;
        RECT 65.405 28.275 65.695 28.505 ;
        RECT 68.625 28.275 68.915 28.505 ;
        RECT 63.090 28.120 63.410 28.180 ;
        RECT 64.485 28.120 64.775 28.165 ;
        RECT 65.480 28.120 65.620 28.275 ;
        RECT 69.070 28.260 69.390 28.520 ;
        RECT 70.465 28.460 70.755 28.505 ;
        RECT 71.845 28.460 72.135 28.505 ;
        RECT 70.465 28.320 72.135 28.460 ;
        RECT 70.465 28.275 70.755 28.320 ;
        RECT 71.845 28.275 72.135 28.320 ;
        RECT 63.090 27.980 65.620 28.120 ;
        RECT 63.090 27.920 63.410 27.980 ;
        RECT 64.485 27.935 64.775 27.980 ;
        RECT 73.210 27.920 73.530 28.180 ;
        RECT 73.670 28.120 73.990 28.180 ;
        RECT 74.145 28.120 74.435 28.165 ;
        RECT 73.670 27.980 74.435 28.120 ;
        RECT 73.670 27.920 73.990 27.980 ;
        RECT 74.145 27.935 74.435 27.980 ;
        RECT 59.870 27.640 61.940 27.780 ;
        RECT 62.185 27.780 62.475 27.825 ;
        RECT 64.010 27.780 64.330 27.840 ;
        RECT 62.185 27.640 64.330 27.780 ;
        RECT 59.870 27.580 60.190 27.640 ;
        RECT 62.185 27.595 62.475 27.640 ;
        RECT 64.010 27.580 64.330 27.640 ;
        RECT 5.520 26.960 76.820 27.440 ;
        RECT 11.110 26.760 11.430 26.820 ;
        RECT 12.045 26.760 12.335 26.805 ;
        RECT 23.990 26.760 24.310 26.820 ;
        RECT 38.250 26.760 38.570 26.820 ;
        RECT 11.110 26.620 25.140 26.760 ;
        RECT 11.110 26.560 11.430 26.620 ;
        RECT 12.045 26.575 12.335 26.620 ;
        RECT 23.990 26.560 24.310 26.620 ;
        RECT 13.870 26.220 14.190 26.480 ;
        RECT 19.865 26.420 20.155 26.465 ;
        RECT 21.230 26.420 21.550 26.480 ;
        RECT 19.865 26.280 21.550 26.420 ;
        RECT 19.865 26.235 20.155 26.280 ;
        RECT 21.230 26.220 21.550 26.280 ;
        RECT 8.365 26.080 8.655 26.125 ;
        RECT 12.965 26.080 13.255 26.125 ;
        RECT 13.960 26.080 14.100 26.220 ;
        RECT 8.365 25.940 16.400 26.080 ;
        RECT 8.365 25.895 8.655 25.940 ;
        RECT 12.965 25.895 13.255 25.940 ;
        RECT 3.750 25.740 4.070 25.800 ;
        RECT 16.260 25.785 16.400 25.940 ;
        RECT 18.930 25.880 19.250 26.140 ;
        RECT 19.390 25.880 19.710 26.140 ;
        RECT 22.150 25.880 22.470 26.140 ;
        RECT 23.545 26.080 23.835 26.125 ;
        RECT 23.990 26.080 24.310 26.140 ;
        RECT 23.545 25.940 24.310 26.080 ;
        RECT 23.545 25.895 23.835 25.940 ;
        RECT 23.990 25.880 24.310 25.940 ;
        RECT 24.450 25.880 24.770 26.140 ;
        RECT 25.000 26.080 25.140 26.620 ;
        RECT 33.280 26.620 38.570 26.760 ;
        RECT 26.765 26.420 27.055 26.465 ;
        RECT 31.350 26.420 31.670 26.480 ;
        RECT 26.765 26.280 31.670 26.420 ;
        RECT 26.765 26.235 27.055 26.280 ;
        RECT 31.350 26.220 31.670 26.280 ;
        RECT 25.845 26.080 26.135 26.125 ;
        RECT 25.000 25.940 26.135 26.080 ;
        RECT 25.845 25.895 26.135 25.940 ;
        RECT 30.890 26.080 31.210 26.140 ;
        RECT 31.825 26.080 32.115 26.125 ;
        RECT 30.890 25.940 32.115 26.080 ;
        RECT 30.890 25.880 31.210 25.940 ;
        RECT 31.825 25.895 32.115 25.940 ;
        RECT 32.270 25.880 32.590 26.140 ;
        RECT 33.280 26.125 33.420 26.620 ;
        RECT 38.250 26.560 38.570 26.620 ;
        RECT 39.630 26.760 39.950 26.820 ;
        RECT 41.470 26.760 41.790 26.820 ;
        RECT 39.630 26.620 41.790 26.760 ;
        RECT 39.630 26.560 39.950 26.620 ;
        RECT 41.470 26.560 41.790 26.620 ;
        RECT 41.930 26.760 42.250 26.820 ;
        RECT 44.705 26.760 44.995 26.805 ;
        RECT 58.950 26.760 59.270 26.820 ;
        RECT 59.885 26.760 60.175 26.805 ;
        RECT 63.550 26.760 63.870 26.820 ;
        RECT 41.930 26.620 44.995 26.760 ;
        RECT 41.930 26.560 42.250 26.620 ;
        RECT 44.705 26.575 44.995 26.620 ;
        RECT 45.240 26.620 58.720 26.760 ;
        RECT 35.490 26.420 35.810 26.480 ;
        RECT 44.230 26.420 44.550 26.480 ;
        RECT 35.490 26.280 44.550 26.420 ;
        RECT 35.490 26.220 35.810 26.280 ;
        RECT 44.230 26.220 44.550 26.280 ;
        RECT 33.205 25.895 33.495 26.125 ;
        RECT 33.665 26.080 33.955 26.125 ;
        RECT 35.045 26.080 35.335 26.125 ;
        RECT 33.665 25.940 35.335 26.080 ;
        RECT 33.665 25.895 33.955 25.940 ;
        RECT 35.045 25.895 35.335 25.940 ;
        RECT 35.965 25.895 36.255 26.125 ;
        RECT 6.985 25.740 7.275 25.785 ;
        RECT 3.750 25.600 7.275 25.740 ;
        RECT 3.750 25.540 4.070 25.600 ;
        RECT 6.985 25.555 7.275 25.600 ;
        RECT 13.885 25.555 14.175 25.785 ;
        RECT 16.185 25.740 16.475 25.785 ;
        RECT 16.630 25.740 16.950 25.800 ;
        RECT 16.185 25.600 16.950 25.740 ;
        RECT 16.185 25.555 16.475 25.600 ;
        RECT 13.960 25.400 14.100 25.555 ;
        RECT 16.630 25.540 16.950 25.600 ;
        RECT 17.105 25.740 17.395 25.785 ;
        RECT 35.490 25.740 35.810 25.800 ;
        RECT 36.040 25.740 36.180 25.895 ;
        RECT 36.870 25.880 37.190 26.140 ;
        RECT 37.330 25.880 37.650 26.140 ;
        RECT 39.630 25.880 39.950 26.140 ;
        RECT 40.565 26.080 40.855 26.125 ;
        RECT 41.010 26.080 41.330 26.140 ;
        RECT 40.565 25.940 41.330 26.080 ;
        RECT 40.565 25.895 40.855 25.940 ;
        RECT 41.010 25.880 41.330 25.940 ;
        RECT 17.105 25.600 36.180 25.740 ;
        RECT 38.250 25.740 38.570 25.800 ;
        RECT 45.240 25.740 45.380 26.620 ;
        RECT 58.580 26.420 58.720 26.620 ;
        RECT 58.950 26.620 60.175 26.760 ;
        RECT 58.950 26.560 59.270 26.620 ;
        RECT 59.885 26.575 60.175 26.620 ;
        RECT 62.260 26.620 63.870 26.760 ;
        RECT 59.410 26.420 59.730 26.480 ;
        RECT 61.265 26.420 61.555 26.465 ;
        RECT 51.220 26.280 58.260 26.420 ;
        RECT 58.580 26.280 61.555 26.420 ;
        RECT 45.610 25.880 45.930 26.140 ;
        RECT 46.070 25.880 46.390 26.140 ;
        RECT 47.465 25.895 47.755 26.125 ;
        RECT 50.670 26.080 50.990 26.140 ;
        RECT 51.220 26.125 51.360 26.280 ;
        RECT 58.120 26.140 58.260 26.280 ;
        RECT 59.410 26.220 59.730 26.280 ;
        RECT 61.265 26.235 61.555 26.280 ;
        RECT 51.145 26.080 51.435 26.125 ;
        RECT 50.670 25.940 51.435 26.080 ;
        RECT 38.250 25.600 45.380 25.740 ;
        RECT 46.530 25.740 46.850 25.800 ;
        RECT 47.540 25.740 47.680 25.895 ;
        RECT 50.670 25.880 50.990 25.940 ;
        RECT 51.145 25.895 51.435 25.940 ;
        RECT 57.585 25.895 57.875 26.125 ;
        RECT 48.830 25.740 49.150 25.800 ;
        RECT 54.810 25.740 55.130 25.800 ;
        RECT 46.530 25.600 55.130 25.740 ;
        RECT 57.660 25.740 57.800 25.895 ;
        RECT 58.030 25.880 58.350 26.140 ;
        RECT 58.950 25.880 59.270 26.140 ;
        RECT 62.260 26.125 62.400 26.620 ;
        RECT 63.550 26.560 63.870 26.620 ;
        RECT 66.785 26.575 67.075 26.805 ;
        RECT 66.860 26.420 67.000 26.575 ;
        RECT 70.910 26.560 71.230 26.820 ;
        RECT 72.290 26.560 72.610 26.820 ;
        RECT 73.670 26.760 73.990 26.820 ;
        RECT 74.145 26.760 74.435 26.805 ;
        RECT 73.670 26.620 74.435 26.760 ;
        RECT 73.670 26.560 73.990 26.620 ;
        RECT 74.145 26.575 74.435 26.620 ;
        RECT 74.605 26.420 74.895 26.465 ;
        RECT 62.720 26.280 74.895 26.420 ;
        RECT 62.185 25.895 62.475 26.125 ;
        RECT 58.490 25.740 58.810 25.800 ;
        RECT 57.660 25.600 58.810 25.740 ;
        RECT 17.105 25.555 17.395 25.600 ;
        RECT 35.490 25.540 35.810 25.600 ;
        RECT 38.250 25.540 38.570 25.600 ;
        RECT 46.530 25.540 46.850 25.600 ;
        RECT 48.830 25.540 49.150 25.600 ;
        RECT 54.810 25.540 55.130 25.600 ;
        RECT 58.490 25.540 58.810 25.600 ;
        RECT 14.330 25.400 14.650 25.460 ;
        RECT 19.390 25.400 19.710 25.460 ;
        RECT 13.960 25.260 19.710 25.400 ;
        RECT 14.330 25.200 14.650 25.260 ;
        RECT 19.390 25.200 19.710 25.260 ;
        RECT 21.230 25.200 21.550 25.460 ;
        RECT 28.130 25.400 28.450 25.460 ;
        RECT 62.720 25.400 62.860 26.280 ;
        RECT 74.605 26.235 74.895 26.280 ;
        RECT 67.690 25.880 68.010 26.140 ;
        RECT 69.530 25.880 69.850 26.140 ;
        RECT 69.990 25.880 70.310 26.140 ;
        RECT 71.830 26.080 72.150 26.140 ;
        RECT 73.210 26.080 73.530 26.140 ;
        RECT 71.830 25.940 73.530 26.080 ;
        RECT 71.830 25.880 72.150 25.940 ;
        RECT 73.210 25.880 73.530 25.940 ;
        RECT 63.105 25.740 63.395 25.785 ;
        RECT 73.670 25.740 73.990 25.800 ;
        RECT 63.105 25.600 73.990 25.740 ;
        RECT 63.105 25.555 63.395 25.600 ;
        RECT 73.670 25.540 73.990 25.600 ;
        RECT 28.130 25.260 62.860 25.400 ;
        RECT 28.130 25.200 28.450 25.260 ;
        RECT 12.030 25.060 12.350 25.120 ;
        RECT 20.310 25.060 20.630 25.120 ;
        RECT 12.030 24.920 20.630 25.060 ;
        RECT 12.030 24.860 12.350 24.920 ;
        RECT 20.310 24.860 20.630 24.920 ;
        RECT 34.570 24.860 34.890 25.120 ;
        RECT 40.550 24.860 40.870 25.120 ;
        RECT 47.005 25.060 47.295 25.105 ;
        RECT 49.290 25.060 49.610 25.120 ;
        RECT 50.210 25.060 50.530 25.120 ;
        RECT 47.005 24.920 50.530 25.060 ;
        RECT 47.005 24.875 47.295 24.920 ;
        RECT 49.290 24.860 49.610 24.920 ;
        RECT 50.210 24.860 50.530 24.920 ;
        RECT 50.685 25.060 50.975 25.105 ;
        RECT 51.130 25.060 51.450 25.120 ;
        RECT 50.685 24.920 51.450 25.060 ;
        RECT 50.685 24.875 50.975 24.920 ;
        RECT 51.130 24.860 51.450 24.920 ;
        RECT 53.430 25.060 53.750 25.120 ;
        RECT 68.150 25.060 68.470 25.120 ;
        RECT 68.625 25.060 68.915 25.105 ;
        RECT 53.430 24.920 68.915 25.060 ;
        RECT 53.430 24.860 53.750 24.920 ;
        RECT 68.150 24.860 68.470 24.920 ;
        RECT 68.625 24.875 68.915 24.920 ;
        RECT 5.520 24.240 76.820 24.720 ;
        RECT 12.030 23.840 12.350 24.100 ;
        RECT 15.710 24.040 16.030 24.100 ;
        RECT 17.105 24.040 17.395 24.085 ;
        RECT 20.770 24.040 21.090 24.100 ;
        RECT 15.710 23.900 21.090 24.040 ;
        RECT 15.710 23.840 16.030 23.900 ;
        RECT 17.105 23.855 17.395 23.900 ;
        RECT 20.770 23.840 21.090 23.900 ;
        RECT 22.165 24.040 22.455 24.085 ;
        RECT 24.925 24.040 25.215 24.085 ;
        RECT 26.750 24.040 27.070 24.100 ;
        RECT 22.165 23.900 27.070 24.040 ;
        RECT 22.165 23.855 22.455 23.900 ;
        RECT 24.925 23.855 25.215 23.900 ;
        RECT 26.750 23.840 27.070 23.900 ;
        RECT 30.890 23.840 31.210 24.100 ;
        RECT 35.950 24.040 36.270 24.100 ;
        RECT 37.805 24.040 38.095 24.085 ;
        RECT 43.770 24.040 44.090 24.100 ;
        RECT 35.950 23.900 38.095 24.040 ;
        RECT 35.950 23.840 36.270 23.900 ;
        RECT 37.805 23.855 38.095 23.900 ;
        RECT 38.800 23.900 44.090 24.040 ;
        RECT 11.585 23.700 11.875 23.745 ;
        RECT 16.630 23.700 16.950 23.760 ;
        RECT 11.585 23.560 16.950 23.700 ;
        RECT 11.585 23.515 11.875 23.560 ;
        RECT 16.630 23.500 16.950 23.560 ;
        RECT 18.025 23.700 18.315 23.745 ;
        RECT 23.990 23.700 24.310 23.760 ;
        RECT 24.465 23.700 24.755 23.745 ;
        RECT 18.025 23.560 24.755 23.700 ;
        RECT 18.025 23.515 18.315 23.560 ;
        RECT 23.990 23.500 24.310 23.560 ;
        RECT 24.465 23.515 24.755 23.560 ;
        RECT 27.670 23.700 27.990 23.760 ;
        RECT 29.985 23.700 30.275 23.745 ;
        RECT 37.330 23.700 37.650 23.760 ;
        RECT 27.670 23.560 37.650 23.700 ;
        RECT 27.670 23.500 27.990 23.560 ;
        RECT 29.985 23.515 30.275 23.560 ;
        RECT 37.330 23.500 37.650 23.560 ;
        RECT 14.790 23.360 15.110 23.420 ;
        RECT 15.265 23.360 15.555 23.405 ;
        RECT 14.790 23.220 15.555 23.360 ;
        RECT 14.790 23.160 15.110 23.220 ;
        RECT 15.265 23.175 15.555 23.220 ;
        RECT 20.310 23.360 20.630 23.420 ;
        RECT 30.430 23.360 30.750 23.420 ;
        RECT 35.045 23.360 35.335 23.405 ;
        RECT 38.800 23.360 38.940 23.900 ;
        RECT 43.770 23.840 44.090 23.900 ;
        RECT 49.765 24.040 50.055 24.085 ;
        RECT 53.430 24.040 53.750 24.100 ;
        RECT 49.765 23.900 53.750 24.040 ;
        RECT 49.765 23.855 50.055 23.900 ;
        RECT 53.430 23.840 53.750 23.900 ;
        RECT 62.170 24.040 62.490 24.100 ;
        RECT 70.465 24.040 70.755 24.085 ;
        RECT 62.170 23.900 70.755 24.040 ;
        RECT 62.170 23.840 62.490 23.900 ;
        RECT 70.465 23.855 70.755 23.900 ;
        RECT 75.050 23.840 75.370 24.100 ;
        RECT 39.170 23.700 39.490 23.760 ;
        RECT 48.830 23.700 49.150 23.760 ;
        RECT 39.170 23.560 49.150 23.700 ;
        RECT 39.170 23.500 39.490 23.560 ;
        RECT 48.830 23.500 49.150 23.560 ;
        RECT 50.670 23.500 50.990 23.760 ;
        RECT 57.110 23.500 57.430 23.760 ;
        RECT 69.530 23.700 69.850 23.760 ;
        RECT 72.765 23.700 73.055 23.745 ;
        RECT 75.970 23.700 76.290 23.760 ;
        RECT 69.530 23.560 76.290 23.700 ;
        RECT 69.530 23.500 69.850 23.560 ;
        RECT 72.765 23.515 73.055 23.560 ;
        RECT 75.970 23.500 76.290 23.560 ;
        RECT 47.465 23.360 47.755 23.405 ;
        RECT 48.370 23.360 48.690 23.420 ;
        RECT 55.285 23.360 55.575 23.405 ;
        RECT 20.310 23.220 29.280 23.360 ;
        RECT 20.310 23.160 20.630 23.220 ;
        RECT 8.350 22.820 8.670 23.080 ;
        RECT 16.630 23.020 16.950 23.080 ;
        RECT 18.945 23.020 19.235 23.065 ;
        RECT 16.630 22.880 19.235 23.020 ;
        RECT 16.630 22.820 16.950 22.880 ;
        RECT 18.945 22.835 19.235 22.880 ;
        RECT 19.850 23.020 20.170 23.080 ;
        RECT 22.610 23.020 22.930 23.080 ;
        RECT 24.450 23.020 24.770 23.080 ;
        RECT 25.385 23.020 25.675 23.065 ;
        RECT 19.850 22.880 22.380 23.020 ;
        RECT 19.850 22.820 20.170 22.880 ;
        RECT 7.890 22.680 8.210 22.740 ;
        RECT 9.745 22.680 10.035 22.725 ;
        RECT 17.105 22.680 17.395 22.725 ;
        RECT 19.390 22.680 19.710 22.740 ;
        RECT 21.370 22.680 21.660 22.725 ;
        RECT 7.890 22.540 21.660 22.680 ;
        RECT 22.240 22.680 22.380 22.880 ;
        RECT 22.610 22.880 25.675 23.020 ;
        RECT 22.610 22.820 22.930 22.880 ;
        RECT 24.450 22.820 24.770 22.880 ;
        RECT 25.385 22.835 25.675 22.880 ;
        RECT 26.765 23.020 27.055 23.065 ;
        RECT 27.670 23.020 27.990 23.080 ;
        RECT 26.765 22.880 27.990 23.020 ;
        RECT 26.765 22.835 27.055 22.880 ;
        RECT 25.460 22.680 25.600 22.835 ;
        RECT 27.670 22.820 27.990 22.880 ;
        RECT 28.130 22.820 28.450 23.080 ;
        RECT 29.140 23.065 29.280 23.220 ;
        RECT 30.430 23.220 33.885 23.360 ;
        RECT 30.430 23.160 30.750 23.220 ;
        RECT 29.065 22.835 29.355 23.065 ;
        RECT 31.825 22.835 32.115 23.065 ;
        RECT 32.745 22.835 33.035 23.065 ;
        RECT 31.900 22.680 32.040 22.835 ;
        RECT 22.240 22.540 23.760 22.680 ;
        RECT 25.460 22.540 32.040 22.680 ;
        RECT 7.890 22.480 8.210 22.540 ;
        RECT 9.745 22.495 10.035 22.540 ;
        RECT 17.105 22.495 17.395 22.540 ;
        RECT 19.390 22.480 19.710 22.540 ;
        RECT 21.370 22.495 21.660 22.540 ;
        RECT 1.910 22.340 2.230 22.400 ;
        RECT 7.445 22.340 7.735 22.385 ;
        RECT 1.910 22.200 7.735 22.340 ;
        RECT 1.910 22.140 2.230 22.200 ;
        RECT 7.445 22.155 7.735 22.200 ;
        RECT 14.790 22.340 15.110 22.400 ;
        RECT 19.850 22.340 20.170 22.400 ;
        RECT 20.325 22.340 20.615 22.385 ;
        RECT 14.790 22.200 20.615 22.340 ;
        RECT 14.790 22.140 15.110 22.200 ;
        RECT 19.850 22.140 20.170 22.200 ;
        RECT 20.325 22.155 20.615 22.200 ;
        RECT 20.770 22.140 21.090 22.400 ;
        RECT 23.070 22.140 23.390 22.400 ;
        RECT 23.620 22.340 23.760 22.540 ;
        RECT 26.305 22.340 26.595 22.385 ;
        RECT 27.685 22.340 27.975 22.385 ;
        RECT 23.620 22.200 27.975 22.340 ;
        RECT 32.820 22.340 32.960 22.835 ;
        RECT 33.190 22.820 33.510 23.080 ;
        RECT 33.745 23.065 33.885 23.220 ;
        RECT 35.045 23.220 38.940 23.360 ;
        RECT 41.100 23.220 47.220 23.360 ;
        RECT 35.045 23.175 35.335 23.220 ;
        RECT 33.670 22.835 33.960 23.065 ;
        RECT 38.730 23.020 39.020 23.065 ;
        RECT 38.730 22.880 40.320 23.020 ;
        RECT 38.730 22.835 39.020 22.880 ;
        RECT 33.745 22.680 33.885 22.835 ;
        RECT 39.170 22.680 39.490 22.740 ;
        RECT 33.745 22.540 39.490 22.680 ;
        RECT 39.170 22.480 39.490 22.540 ;
        RECT 39.630 22.480 39.950 22.740 ;
        RECT 40.180 22.680 40.320 22.880 ;
        RECT 40.550 22.820 40.870 23.080 ;
        RECT 41.100 23.065 41.240 23.220 ;
        RECT 41.025 22.835 41.315 23.065 ;
        RECT 42.865 23.020 43.155 23.065 ;
        RECT 43.770 23.020 44.090 23.080 ;
        RECT 42.865 22.880 44.090 23.020 ;
        RECT 42.865 22.835 43.155 22.880 ;
        RECT 43.770 22.820 44.090 22.880 ;
        RECT 43.310 22.680 43.630 22.740 ;
        RECT 40.180 22.540 43.630 22.680 ;
        RECT 47.080 22.680 47.220 23.220 ;
        RECT 47.465 23.220 48.690 23.360 ;
        RECT 47.465 23.175 47.755 23.220 ;
        RECT 48.370 23.160 48.690 23.220 ;
        RECT 49.840 23.220 52.740 23.360 ;
        RECT 49.840 23.080 49.980 23.220 ;
        RECT 47.910 22.820 48.230 23.080 ;
        RECT 49.750 22.820 50.070 23.080 ;
        RECT 52.050 22.820 52.370 23.080 ;
        RECT 52.600 23.065 52.740 23.220 ;
        RECT 55.285 23.220 58.720 23.360 ;
        RECT 55.285 23.175 55.575 23.220 ;
        RECT 58.580 23.080 58.720 23.220 ;
        RECT 52.525 22.835 52.815 23.065 ;
        RECT 53.430 22.820 53.750 23.080 ;
        RECT 58.030 22.820 58.350 23.080 ;
        RECT 58.490 22.820 58.810 23.080 ;
        RECT 66.310 23.020 66.630 23.080 ;
        RECT 71.385 23.020 71.675 23.065 ;
        RECT 66.310 22.880 71.675 23.020 ;
        RECT 66.310 22.820 66.630 22.880 ;
        RECT 71.385 22.835 71.675 22.880 ;
        RECT 73.670 22.820 73.990 23.080 ;
        RECT 74.130 22.820 74.450 23.080 ;
        RECT 56.650 22.680 56.970 22.740 ;
        RECT 47.080 22.540 56.970 22.680 ;
        RECT 43.310 22.480 43.630 22.540 ;
        RECT 56.650 22.480 56.970 22.540 ;
        RECT 57.125 22.680 57.415 22.725 ;
        RECT 58.950 22.680 59.270 22.740 ;
        RECT 57.125 22.540 59.270 22.680 ;
        RECT 57.125 22.495 57.415 22.540 ;
        RECT 34.570 22.340 34.890 22.400 ;
        RECT 32.820 22.200 34.890 22.340 ;
        RECT 26.305 22.155 26.595 22.200 ;
        RECT 27.685 22.155 27.975 22.200 ;
        RECT 34.570 22.140 34.890 22.200 ;
        RECT 41.470 22.340 41.790 22.400 ;
        RECT 41.945 22.340 42.235 22.385 ;
        RECT 46.070 22.340 46.390 22.400 ;
        RECT 46.990 22.340 47.310 22.400 ;
        RECT 57.200 22.340 57.340 22.495 ;
        RECT 58.950 22.480 59.270 22.540 ;
        RECT 41.470 22.200 57.340 22.340 ;
        RECT 41.470 22.140 41.790 22.200 ;
        RECT 41.945 22.155 42.235 22.200 ;
        RECT 46.070 22.140 46.390 22.200 ;
        RECT 46.990 22.140 47.310 22.200 ;
        RECT 5.520 21.520 76.820 22.000 ;
        RECT 8.350 21.320 8.670 21.380 ;
        RECT 9.285 21.320 9.575 21.365 ;
        RECT 8.350 21.180 9.575 21.320 ;
        RECT 8.350 21.120 8.670 21.180 ;
        RECT 9.285 21.135 9.575 21.180 ;
        RECT 16.630 21.120 16.950 21.380 ;
        RECT 23.990 21.120 24.310 21.380 ;
        RECT 34.570 21.320 34.890 21.380 ;
        RECT 40.090 21.320 40.410 21.380 ;
        RECT 34.570 21.180 40.410 21.320 ;
        RECT 34.570 21.120 34.890 21.180 ;
        RECT 40.090 21.120 40.410 21.180 ;
        RECT 43.310 21.320 43.630 21.380 ;
        RECT 49.765 21.320 50.055 21.365 ;
        RECT 43.310 21.180 50.055 21.320 ;
        RECT 43.310 21.120 43.630 21.180 ;
        RECT 49.765 21.135 50.055 21.180 ;
        RECT 50.670 21.320 50.990 21.380 ;
        RECT 55.745 21.320 56.035 21.365 ;
        RECT 58.045 21.320 58.335 21.365 ;
        RECT 50.670 21.180 58.335 21.320 ;
        RECT 50.670 21.120 50.990 21.180 ;
        RECT 55.745 21.135 56.035 21.180 ;
        RECT 58.045 21.135 58.335 21.180 ;
        RECT 23.085 20.795 23.375 21.025 ;
        RECT 24.080 20.980 24.220 21.120 ;
        RECT 42.405 20.980 42.695 21.025 ;
        RECT 45.150 20.980 45.470 21.040 ;
        RECT 47.450 20.980 47.770 21.040 ;
        RECT 48.830 20.980 49.150 21.040 ;
        RECT 24.080 20.840 26.060 20.980 ;
        RECT 7.890 20.440 8.210 20.700 ;
        RECT 8.365 20.640 8.655 20.685 ;
        RECT 10.205 20.640 10.495 20.685 ;
        RECT 8.365 20.500 10.495 20.640 ;
        RECT 8.365 20.455 8.655 20.500 ;
        RECT 10.205 20.455 10.495 20.500 ;
        RECT 14.805 20.640 15.095 20.685 ;
        RECT 15.710 20.640 16.030 20.700 ;
        RECT 22.610 20.640 22.930 20.700 ;
        RECT 23.160 20.640 23.300 20.795 ;
        RECT 25.920 20.685 26.060 20.840 ;
        RECT 38.800 20.840 45.470 20.980 ;
        RECT 14.805 20.500 16.030 20.640 ;
        RECT 14.805 20.455 15.095 20.500 ;
        RECT 15.710 20.440 16.030 20.500 ;
        RECT 17.640 20.500 23.300 20.640 ;
        RECT 17.640 20.005 17.780 20.500 ;
        RECT 22.610 20.440 22.930 20.500 ;
        RECT 24.005 20.455 24.295 20.685 ;
        RECT 24.465 20.455 24.755 20.685 ;
        RECT 25.845 20.455 26.135 20.685 ;
        RECT 24.080 20.300 24.220 20.455 ;
        RECT 21.780 20.160 24.220 20.300 ;
        RECT 24.540 20.300 24.680 20.455 ;
        RECT 26.750 20.440 27.070 20.700 ;
        RECT 38.800 20.685 38.940 20.840 ;
        RECT 42.405 20.795 42.695 20.840 ;
        RECT 45.150 20.780 45.470 20.840 ;
        RECT 46.160 20.840 49.150 20.980 ;
        RECT 38.725 20.455 39.015 20.685 ;
        RECT 39.170 20.440 39.490 20.700 ;
        RECT 39.630 20.440 39.950 20.700 ;
        RECT 40.565 20.455 40.855 20.685 ;
        RECT 41.025 20.640 41.315 20.685 ;
        RECT 42.850 20.640 43.170 20.700 ;
        RECT 41.025 20.500 43.170 20.640 ;
        RECT 41.025 20.455 41.315 20.500 ;
        RECT 27.670 20.300 27.990 20.360 ;
        RECT 24.540 20.160 27.990 20.300 ;
        RECT 17.565 19.775 17.855 20.005 ;
        RECT 14.790 19.620 15.110 19.680 ;
        RECT 16.645 19.620 16.935 19.665 ;
        RECT 21.780 19.620 21.920 20.160 ;
        RECT 27.670 20.100 27.990 20.160 ;
        RECT 33.650 20.300 33.970 20.360 ;
        RECT 39.720 20.300 39.860 20.440 ;
        RECT 33.650 20.160 39.860 20.300 ;
        RECT 40.640 20.300 40.780 20.455 ;
        RECT 42.850 20.440 43.170 20.500 ;
        RECT 43.310 20.440 43.630 20.700 ;
        RECT 43.770 20.440 44.090 20.700 ;
        RECT 44.705 20.455 44.995 20.685 ;
        RECT 45.610 20.640 45.930 20.700 ;
        RECT 46.160 20.685 46.300 20.840 ;
        RECT 47.450 20.780 47.770 20.840 ;
        RECT 48.830 20.780 49.150 20.840 ;
        RECT 54.810 20.980 55.130 21.040 ;
        RECT 56.665 20.980 56.955 21.025 ;
        RECT 54.810 20.840 59.180 20.980 ;
        RECT 54.810 20.780 55.130 20.840 ;
        RECT 56.665 20.795 56.955 20.840 ;
        RECT 46.085 20.640 46.375 20.685 ;
        RECT 45.610 20.500 46.375 20.640 ;
        RECT 44.245 20.300 44.535 20.345 ;
        RECT 40.640 20.160 44.535 20.300 ;
        RECT 44.780 20.300 44.920 20.455 ;
        RECT 45.610 20.440 45.930 20.500 ;
        RECT 46.085 20.455 46.375 20.500 ;
        RECT 46.530 20.440 46.850 20.700 ;
        RECT 46.990 20.640 47.310 20.700 ;
        RECT 47.925 20.640 48.215 20.685 ;
        RECT 49.290 20.640 49.610 20.730 ;
        RECT 46.990 20.500 48.215 20.640 ;
        RECT 46.990 20.440 47.310 20.500 ;
        RECT 47.925 20.455 48.215 20.500 ;
        RECT 48.920 20.500 49.775 20.640 ;
        RECT 46.620 20.300 46.760 20.440 ;
        RECT 44.780 20.160 46.760 20.300 ;
        RECT 47.465 20.300 47.755 20.345 ;
        RECT 48.920 20.300 49.060 20.500 ;
        RECT 49.290 20.470 49.610 20.500 ;
        RECT 49.305 20.455 49.595 20.470 ;
        RECT 50.210 20.440 50.530 20.700 ;
        RECT 50.670 20.440 50.990 20.700 ;
        RECT 51.590 20.640 51.910 20.700 ;
        RECT 59.040 20.685 59.180 20.840 ;
        RECT 55.285 20.670 55.575 20.685 ;
        RECT 55.285 20.640 56.275 20.670 ;
        RECT 57.585 20.640 57.875 20.685 ;
        RECT 51.590 20.530 57.875 20.640 ;
        RECT 51.590 20.500 55.575 20.530 ;
        RECT 56.135 20.500 57.875 20.530 ;
        RECT 51.590 20.440 51.910 20.500 ;
        RECT 55.285 20.455 55.575 20.500 ;
        RECT 57.585 20.455 57.875 20.500 ;
        RECT 58.965 20.455 59.255 20.685 ;
        RECT 59.870 20.440 60.190 20.700 ;
        RECT 47.465 20.160 49.060 20.300 ;
        RECT 33.650 20.100 33.970 20.160 ;
        RECT 44.245 20.115 44.535 20.160 ;
        RECT 47.465 20.115 47.755 20.160 ;
        RECT 22.150 19.960 22.470 20.020 ;
        RECT 24.450 19.960 24.770 20.020 ;
        RECT 22.150 19.820 24.770 19.960 ;
        RECT 22.150 19.760 22.470 19.820 ;
        RECT 24.450 19.760 24.770 19.820 ;
        RECT 37.790 19.760 38.110 20.020 ;
        RECT 41.010 19.960 41.330 20.020 ;
        RECT 41.485 19.960 41.775 20.005 ;
        RECT 43.770 19.960 44.090 20.020 ;
        RECT 41.010 19.820 44.090 19.960 ;
        RECT 41.010 19.760 41.330 19.820 ;
        RECT 41.485 19.775 41.775 19.820 ;
        RECT 43.770 19.760 44.090 19.820 ;
        RECT 44.690 19.960 45.010 20.020 ;
        RECT 45.165 19.960 45.455 20.005 ;
        RECT 44.690 19.820 45.455 19.960 ;
        RECT 44.690 19.760 45.010 19.820 ;
        RECT 45.165 19.775 45.455 19.820 ;
        RECT 45.610 19.960 45.930 20.020 ;
        RECT 51.145 19.960 51.435 20.005 ;
        RECT 45.610 19.820 51.435 19.960 ;
        RECT 45.610 19.760 45.930 19.820 ;
        RECT 51.145 19.775 51.435 19.820 ;
        RECT 56.650 19.760 56.970 20.020 ;
        RECT 14.790 19.480 21.920 19.620 ;
        RECT 23.085 19.620 23.375 19.665 ;
        RECT 23.990 19.620 24.310 19.680 ;
        RECT 23.085 19.480 24.310 19.620 ;
        RECT 14.790 19.420 15.110 19.480 ;
        RECT 16.645 19.435 16.935 19.480 ;
        RECT 23.085 19.435 23.375 19.480 ;
        RECT 23.990 19.420 24.310 19.480 ;
        RECT 26.750 19.420 27.070 19.680 ;
        RECT 42.850 19.620 43.170 19.680 ;
        RECT 57.110 19.620 57.430 19.680 ;
        RECT 42.850 19.480 57.430 19.620 ;
        RECT 42.850 19.420 43.170 19.480 ;
        RECT 57.110 19.420 57.430 19.480 ;
        RECT 5.520 18.800 76.820 19.280 ;
        RECT 23.545 18.600 23.835 18.645 ;
        RECT 26.290 18.600 26.610 18.660 ;
        RECT 23.545 18.460 26.610 18.600 ;
        RECT 23.545 18.415 23.835 18.460 ;
        RECT 26.290 18.400 26.610 18.460 ;
        RECT 28.145 18.600 28.435 18.645 ;
        RECT 29.050 18.600 29.370 18.660 ;
        RECT 28.145 18.460 29.370 18.600 ;
        RECT 28.145 18.415 28.435 18.460 ;
        RECT 29.050 18.400 29.370 18.460 ;
        RECT 35.045 18.600 35.335 18.645 ;
        RECT 46.530 18.600 46.850 18.660 ;
        RECT 48.370 18.600 48.690 18.660 ;
        RECT 35.045 18.460 46.850 18.600 ;
        RECT 35.045 18.415 35.335 18.460 ;
        RECT 46.530 18.400 46.850 18.460 ;
        RECT 47.080 18.460 48.690 18.600 ;
        RECT 24.450 18.060 24.770 18.320 ;
        RECT 24.925 18.260 25.215 18.305 ;
        RECT 27.670 18.260 27.990 18.320 ;
        RECT 24.925 18.120 27.990 18.260 ;
        RECT 24.925 18.075 25.215 18.120 ;
        RECT 27.670 18.060 27.990 18.120 ;
        RECT 30.430 18.260 30.750 18.320 ;
        RECT 47.080 18.260 47.220 18.460 ;
        RECT 48.370 18.400 48.690 18.460 ;
        RECT 49.305 18.600 49.595 18.645 ;
        RECT 50.670 18.600 50.990 18.660 ;
        RECT 49.305 18.460 50.990 18.600 ;
        RECT 49.305 18.415 49.595 18.460 ;
        RECT 50.670 18.400 50.990 18.460 ;
        RECT 30.430 18.120 47.220 18.260 ;
        RECT 47.450 18.260 47.770 18.320 ;
        RECT 50.225 18.260 50.515 18.305 ;
        RECT 47.450 18.120 50.515 18.260 ;
        RECT 30.430 18.060 30.750 18.120 ;
        RECT 47.450 18.060 47.770 18.120 ;
        RECT 50.225 18.075 50.515 18.120 ;
        RECT 73.210 18.260 73.530 18.320 ;
        RECT 73.685 18.260 73.975 18.305 ;
        RECT 73.210 18.120 73.975 18.260 ;
        RECT 73.210 18.060 73.530 18.120 ;
        RECT 73.685 18.075 73.975 18.120 ;
        RECT 24.540 17.920 24.680 18.060 ;
        RECT 27.225 17.920 27.515 17.965 ;
        RECT 28.130 17.920 28.450 17.980 ;
        RECT 24.540 17.780 28.450 17.920 ;
        RECT 27.225 17.735 27.515 17.780 ;
        RECT 28.130 17.720 28.450 17.780 ;
        RECT 40.090 17.920 40.410 17.980 ;
        RECT 40.090 17.780 46.760 17.920 ;
        RECT 40.090 17.720 40.410 17.780 ;
        RECT 23.070 17.580 23.390 17.640 ;
        RECT 24.465 17.580 24.755 17.625 ;
        RECT 23.070 17.440 24.755 17.580 ;
        RECT 23.070 17.380 23.390 17.440 ;
        RECT 24.465 17.395 24.755 17.440 ;
        RECT 25.385 17.395 25.675 17.625 ;
        RECT 25.845 17.395 26.135 17.625 ;
        RECT 25.460 16.900 25.600 17.395 ;
        RECT 25.920 17.240 26.060 17.395 ;
        RECT 26.750 17.380 27.070 17.640 ;
        RECT 28.605 17.580 28.895 17.625 ;
        RECT 29.510 17.580 29.830 17.640 ;
        RECT 28.605 17.440 29.830 17.580 ;
        RECT 28.605 17.395 28.895 17.440 ;
        RECT 29.510 17.380 29.830 17.440 ;
        RECT 33.650 17.380 33.970 17.640 ;
        RECT 35.490 17.580 35.810 17.640 ;
        RECT 39.170 17.580 39.490 17.640 ;
        RECT 46.620 17.625 46.760 17.780 ;
        RECT 49.840 17.780 52.740 17.920 ;
        RECT 49.840 17.640 49.980 17.780 ;
        RECT 35.490 17.440 39.490 17.580 ;
        RECT 35.490 17.380 35.810 17.440 ;
        RECT 39.170 17.380 39.490 17.440 ;
        RECT 46.085 17.395 46.375 17.625 ;
        RECT 46.545 17.580 46.835 17.625 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 46.545 17.440 48.230 17.580 ;
        RECT 46.545 17.395 46.835 17.440 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 27.225 17.240 27.515 17.285 ;
        RECT 25.920 17.100 27.515 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 27.225 17.055 27.515 17.100 ;
        RECT 29.050 17.240 29.370 17.300 ;
        RECT 46.160 17.240 46.300 17.395 ;
        RECT 47.910 17.380 48.230 17.440 ;
        RECT 48.385 17.580 48.675 17.625 ;
        RECT 49.750 17.580 50.070 17.640 ;
        RECT 48.385 17.440 50.070 17.580 ;
        RECT 48.385 17.395 48.675 17.440 ;
        RECT 49.750 17.380 50.070 17.440 ;
        RECT 52.050 17.380 52.370 17.640 ;
        RECT 52.600 17.625 52.740 17.780 ;
        RECT 52.525 17.395 52.815 17.625 ;
        RECT 53.430 17.380 53.750 17.640 ;
        RECT 53.520 17.240 53.660 17.380 ;
        RECT 29.050 17.100 53.660 17.240 ;
        RECT 29.050 17.040 29.370 17.100 ;
        RECT 74.590 17.040 74.910 17.300 ;
        RECT 26.750 16.900 27.070 16.960 ;
        RECT 25.460 16.760 27.070 16.900 ;
        RECT 26.750 16.700 27.070 16.760 ;
        RECT 5.520 16.080 76.820 16.560 ;
        RECT 23.085 15.880 23.375 15.925 ;
        RECT 27.210 15.880 27.530 15.940 ;
        RECT 23.085 15.740 27.530 15.880 ;
        RECT 23.085 15.695 23.375 15.740 ;
        RECT 27.210 15.680 27.530 15.740 ;
        RECT 29.510 15.880 29.830 15.940 ;
        RECT 32.745 15.880 33.035 15.925 ;
        RECT 35.490 15.880 35.810 15.940 ;
        RECT 29.510 15.740 35.810 15.880 ;
        RECT 29.510 15.680 29.830 15.740 ;
        RECT 32.745 15.695 33.035 15.740 ;
        RECT 35.490 15.680 35.810 15.740 ;
        RECT 26.765 15.540 27.055 15.585 ;
        RECT 30.445 15.540 30.735 15.585 ;
        RECT 33.190 15.540 33.510 15.600 ;
        RECT 24.540 15.400 27.055 15.540 ;
        RECT 23.070 15.200 23.390 15.260 ;
        RECT 24.540 15.245 24.680 15.400 ;
        RECT 26.765 15.355 27.055 15.400 ;
        RECT 27.760 15.400 30.735 15.540 ;
        RECT 27.760 15.260 27.900 15.400 ;
        RECT 30.445 15.355 30.735 15.400 ;
        RECT 30.980 15.400 33.510 15.540 ;
        RECT 24.005 15.200 24.295 15.245 ;
        RECT 23.070 15.060 24.295 15.200 ;
        RECT 23.070 15.000 23.390 15.060 ;
        RECT 24.005 15.015 24.295 15.060 ;
        RECT 24.465 15.015 24.755 15.245 ;
        RECT 25.830 15.000 26.150 15.260 ;
        RECT 26.305 15.015 26.595 15.245 ;
        RECT 27.225 15.200 27.515 15.245 ;
        RECT 27.670 15.200 27.990 15.260 ;
        RECT 27.225 15.060 27.990 15.200 ;
        RECT 27.225 15.015 27.515 15.060 ;
        RECT 26.380 14.860 26.520 15.015 ;
        RECT 27.670 15.000 27.990 15.060 ;
        RECT 28.605 15.015 28.895 15.245 ;
        RECT 26.750 14.860 27.070 14.920 ;
        RECT 26.380 14.720 27.070 14.860 ;
        RECT 28.680 14.860 28.820 15.015 ;
        RECT 29.510 15.000 29.830 15.260 ;
        RECT 29.970 15.000 30.290 15.260 ;
        RECT 30.980 15.245 31.120 15.400 ;
        RECT 33.190 15.340 33.510 15.400 ;
        RECT 30.905 15.015 31.195 15.245 ;
        RECT 32.285 15.200 32.575 15.245 ;
        RECT 32.730 15.200 33.050 15.260 ;
        RECT 32.285 15.060 33.050 15.200 ;
        RECT 32.285 15.015 32.575 15.060 ;
        RECT 30.980 14.860 31.120 15.015 ;
        RECT 32.730 15.000 33.050 15.060 ;
        RECT 33.665 15.200 33.955 15.245 ;
        RECT 36.870 15.200 37.190 15.260 ;
        RECT 33.665 15.060 37.190 15.200 ;
        RECT 33.665 15.015 33.955 15.060 ;
        RECT 36.870 15.000 37.190 15.060 ;
        RECT 28.680 14.720 31.120 14.860 ;
        RECT 26.750 14.660 27.070 14.720 ;
        RECT 75.050 14.660 75.370 14.920 ;
        RECT 23.990 14.520 24.310 14.580 ;
        RECT 25.385 14.520 25.675 14.565 ;
        RECT 23.990 14.380 25.675 14.520 ;
        RECT 23.990 14.320 24.310 14.380 ;
        RECT 25.385 14.335 25.675 14.380 ;
        RECT 27.685 14.520 27.975 14.565 ;
        RECT 28.130 14.520 28.450 14.580 ;
        RECT 27.685 14.380 28.450 14.520 ;
        RECT 27.685 14.335 27.975 14.380 ;
        RECT 28.130 14.320 28.450 14.380 ;
        RECT 34.585 14.180 34.875 14.225 ;
        RECT 35.950 14.180 36.270 14.240 ;
        RECT 34.585 14.040 36.270 14.180 ;
        RECT 34.585 13.995 34.875 14.040 ;
        RECT 35.950 13.980 36.270 14.040 ;
        RECT 5.520 13.360 76.820 13.840 ;
        RECT 23.530 13.160 23.850 13.220 ;
        RECT 24.005 13.160 24.295 13.205 ;
        RECT 23.530 13.020 24.295 13.160 ;
        RECT 23.530 12.960 23.850 13.020 ;
        RECT 24.005 12.975 24.295 13.020 ;
        RECT 25.845 13.160 26.135 13.205 ;
        RECT 26.750 13.160 27.070 13.220 ;
        RECT 29.510 13.160 29.830 13.220 ;
        RECT 25.845 13.020 27.070 13.160 ;
        RECT 25.845 12.975 26.135 13.020 ;
        RECT 26.750 12.960 27.070 13.020 ;
        RECT 27.300 13.020 29.830 13.160 ;
        RECT 12.950 12.140 13.270 12.200 ;
        RECT 13.425 12.140 13.715 12.185 ;
        RECT 12.950 12.000 13.715 12.140 ;
        RECT 12.950 11.940 13.270 12.000 ;
        RECT 13.425 11.955 13.715 12.000 ;
        RECT 22.610 12.140 22.930 12.200 ;
        RECT 23.085 12.140 23.375 12.185 ;
        RECT 22.610 12.000 23.375 12.140 ;
        RECT 22.610 11.940 22.930 12.000 ;
        RECT 23.085 11.955 23.375 12.000 ;
        RECT 26.765 12.140 27.055 12.185 ;
        RECT 27.300 12.140 27.440 13.020 ;
        RECT 29.510 12.960 29.830 13.020 ;
        RECT 30.905 13.160 31.195 13.205 ;
        RECT 32.730 13.160 33.050 13.220 ;
        RECT 30.905 13.020 33.050 13.160 ;
        RECT 30.905 12.975 31.195 13.020 ;
        RECT 32.730 12.960 33.050 13.020 ;
        RECT 33.650 12.960 33.970 13.220 ;
        RECT 29.065 12.820 29.355 12.865 ;
        RECT 34.570 12.820 34.890 12.880 ;
        RECT 29.065 12.680 34.890 12.820 ;
        RECT 29.065 12.635 29.355 12.680 ;
        RECT 34.570 12.620 34.890 12.680 ;
        RECT 27.685 12.480 27.975 12.525 ;
        RECT 30.430 12.480 30.750 12.540 ;
        RECT 27.685 12.340 30.750 12.480 ;
        RECT 27.685 12.295 27.975 12.340 ;
        RECT 30.430 12.280 30.750 12.340 ;
        RECT 26.765 12.000 27.440 12.140 ;
        RECT 26.765 11.955 27.055 12.000 ;
        RECT 28.145 11.955 28.435 12.185 ;
        RECT 29.050 12.140 29.370 12.200 ;
        RECT 29.985 12.140 30.275 12.185 ;
        RECT 29.050 12.000 30.275 12.140 ;
        RECT 26.290 11.800 26.610 11.860 ;
        RECT 28.220 11.800 28.360 11.955 ;
        RECT 29.050 11.940 29.370 12.000 ;
        RECT 29.985 11.955 30.275 12.000 ;
        RECT 35.950 11.940 36.270 12.200 ;
        RECT 26.290 11.660 28.360 11.800 ;
        RECT 32.270 11.800 32.590 11.860 ;
        RECT 33.205 11.800 33.495 11.845 ;
        RECT 32.270 11.660 33.495 11.800 ;
        RECT 26.290 11.600 26.610 11.660 ;
        RECT 32.270 11.600 32.590 11.660 ;
        RECT 33.205 11.615 33.495 11.660 ;
        RECT 35.490 11.460 35.810 11.520 ;
        RECT 36.885 11.460 37.175 11.505 ;
        RECT 35.490 11.320 37.175 11.460 ;
        RECT 35.490 11.260 35.810 11.320 ;
        RECT 36.885 11.275 37.175 11.320 ;
        RECT 5.520 10.640 76.820 11.120 ;
      LAYER met2 ;
        RECT 0.160 52.690 0.300 92.570 ;
        RECT 2.860 68.350 3.120 68.670 ;
        RECT 0.100 52.370 0.360 52.690 ;
        RECT 1.010 47.755 1.290 48.125 ;
        RECT 1.020 47.610 1.280 47.755 ;
        RECT 2.920 42.685 3.060 68.350 ;
        RECT 3.380 53.030 3.520 92.570 ;
        RECT 4.240 87.390 4.500 87.710 ;
        RECT 3.770 71.555 4.050 71.925 ;
        RECT 3.840 71.390 3.980 71.555 ;
        RECT 3.780 71.070 4.040 71.390 ;
        RECT 3.780 62.910 4.040 63.230 ;
        RECT 3.840 61.725 3.980 62.910 ;
        RECT 3.770 61.355 4.050 61.725 ;
        RECT 3.770 57.955 4.050 58.325 ;
        RECT 3.780 57.810 4.040 57.955 ;
        RECT 3.780 55.430 4.040 55.750 ;
        RECT 3.840 54.925 3.980 55.430 ;
        RECT 3.770 54.555 4.050 54.925 ;
        RECT 3.320 52.710 3.580 53.030 ;
        RECT 4.300 47.590 4.440 87.390 ;
        RECT 6.070 81.755 6.350 82.125 ;
        RECT 5.160 80.250 5.420 80.570 ;
        RECT 5.220 67.050 5.360 80.250 ;
        RECT 6.140 79.890 6.280 81.755 ;
        RECT 6.600 81.250 6.740 92.570 ;
        RECT 9.820 87.710 9.960 92.570 ;
        RECT 11.140 92.490 11.400 92.810 ;
        RECT 10.220 90.790 10.480 91.110 ;
        RECT 9.760 87.390 10.020 87.710 ;
        RECT 6.540 80.930 6.800 81.250 ;
        RECT 9.760 79.910 10.020 80.230 ;
        RECT 6.080 79.570 6.340 79.890 ;
        RECT 6.530 78.355 6.810 78.725 ;
        RECT 6.070 74.955 6.350 75.325 ;
        RECT 5.610 68.155 5.890 68.525 ;
        RECT 5.680 67.650 5.820 68.155 ;
        RECT 5.620 67.330 5.880 67.650 ;
        RECT 5.220 66.910 5.820 67.050 ;
        RECT 4.690 64.755 4.970 65.125 ;
        RECT 4.760 64.590 4.900 64.755 ;
        RECT 4.700 64.270 4.960 64.590 ;
        RECT 5.160 63.590 5.420 63.910 ;
        RECT 4.240 47.270 4.500 47.590 ;
        RECT 2.850 42.315 3.130 42.685 ;
        RECT 3.770 30.755 4.050 31.125 ;
        RECT 4.700 30.950 4.960 31.270 ;
        RECT 3.780 30.610 4.040 30.755 ;
        RECT 4.760 27.725 4.900 30.950 ;
        RECT 5.220 27.870 5.360 63.590 ;
        RECT 5.680 52.350 5.820 66.910 ;
        RECT 6.140 54.050 6.280 74.955 ;
        RECT 6.080 53.730 6.340 54.050 ;
        RECT 6.600 53.710 6.740 78.355 ;
        RECT 9.300 77.530 9.560 77.850 ;
        RECT 7.920 76.510 8.180 76.830 ;
        RECT 7.460 72.090 7.720 72.410 ;
        RECT 7.520 70.030 7.660 72.090 ;
        RECT 7.460 69.710 7.720 70.030 ;
        RECT 7.520 66.630 7.660 69.710 ;
        RECT 7.460 66.310 7.720 66.630 ;
        RECT 6.990 62.715 7.270 63.085 ;
        RECT 7.060 56.430 7.200 62.715 ;
        RECT 7.520 56.770 7.660 66.310 ;
        RECT 7.460 56.450 7.720 56.770 ;
        RECT 7.000 56.110 7.260 56.430 ;
        RECT 6.540 53.390 6.800 53.710 ;
        RECT 7.980 53.370 8.120 76.510 ;
        RECT 8.840 71.750 9.100 72.070 ;
        RECT 8.380 63.930 8.640 64.250 ;
        RECT 8.440 62.210 8.580 63.930 ;
        RECT 8.380 61.890 8.640 62.210 ;
        RECT 8.900 61.870 9.040 71.750 ;
        RECT 9.360 70.565 9.500 77.530 ;
        RECT 9.820 77.170 9.960 79.910 ;
        RECT 9.760 76.850 10.020 77.170 ;
        RECT 9.290 70.195 9.570 70.565 ;
        RECT 9.300 69.030 9.560 69.350 ;
        RECT 9.360 67.310 9.500 69.030 ;
        RECT 9.300 66.990 9.560 67.310 ;
        RECT 9.820 64.330 9.960 76.850 ;
        RECT 10.280 74.790 10.420 90.790 ;
        RECT 11.200 80.910 11.340 92.490 ;
        RECT 12.060 83.990 12.320 84.310 ;
        RECT 12.120 80.910 12.260 83.990 ;
        RECT 13.040 83.485 13.180 92.570 ;
        RECT 14.810 83.795 15.090 84.165 ;
        RECT 12.970 83.115 13.250 83.485 ;
        RECT 12.510 82.435 12.790 82.805 ;
        RECT 11.140 80.590 11.400 80.910 ;
        RECT 12.060 80.590 12.320 80.910 ;
        RECT 11.600 80.250 11.860 80.570 ;
        RECT 11.130 79.715 11.410 80.085 ;
        RECT 11.200 77.510 11.340 79.715 ;
        RECT 11.140 77.190 11.400 77.510 ;
        RECT 10.220 74.470 10.480 74.790 ;
        RECT 10.680 71.750 10.940 72.070 ;
        RECT 10.220 69.370 10.480 69.690 ;
        RECT 9.360 64.190 9.960 64.330 ;
        RECT 8.840 61.550 9.100 61.870 ;
        RECT 8.380 60.190 8.640 60.510 ;
        RECT 8.840 60.190 9.100 60.510 ;
        RECT 8.440 58.810 8.580 60.190 ;
        RECT 8.380 58.490 8.640 58.810 ;
        RECT 8.900 58.210 9.040 60.190 ;
        RECT 8.440 58.070 9.040 58.210 ;
        RECT 7.920 53.050 8.180 53.370 ;
        RECT 5.620 52.030 5.880 52.350 ;
        RECT 8.440 48.370 8.580 58.070 ;
        RECT 9.360 56.285 9.500 64.190 ;
        RECT 9.750 63.395 10.030 63.765 ;
        RECT 9.820 61.190 9.960 63.395 ;
        RECT 10.280 63.230 10.420 69.370 ;
        RECT 10.740 67.650 10.880 71.750 ;
        RECT 11.660 71.245 11.800 80.250 ;
        RECT 12.060 77.420 12.320 77.510 ;
        RECT 12.580 77.420 12.720 82.435 ;
        RECT 14.880 79.890 15.020 83.795 ;
        RECT 15.740 80.250 16.000 80.570 ;
        RECT 14.820 79.570 15.080 79.890 ;
        RECT 12.060 77.280 12.720 77.420 ;
        RECT 12.060 77.190 12.320 77.280 ;
        RECT 12.980 77.190 13.240 77.510 ;
        RECT 13.440 77.190 13.700 77.510 ;
        RECT 12.520 76.510 12.780 76.830 ;
        RECT 11.590 70.875 11.870 71.245 ;
        RECT 12.060 69.030 12.320 69.350 ;
        RECT 12.580 69.090 12.720 76.510 ;
        RECT 13.040 75.325 13.180 77.190 ;
        RECT 12.970 74.955 13.250 75.325 ;
        RECT 13.500 74.645 13.640 77.190 ;
        RECT 14.360 76.850 14.620 77.170 ;
        RECT 14.820 76.850 15.080 77.170 ;
        RECT 15.270 76.995 15.550 77.365 ;
        RECT 14.420 75.470 14.560 76.850 ;
        RECT 14.880 75.810 15.020 76.850 ;
        RECT 14.820 75.490 15.080 75.810 ;
        RECT 14.360 75.150 14.620 75.470 ;
        RECT 13.430 74.275 13.710 74.645 ;
        RECT 13.900 73.790 14.160 74.110 ;
        RECT 12.980 71.750 13.240 72.070 ;
        RECT 13.040 71.245 13.180 71.750 ;
        RECT 12.970 70.875 13.250 71.245 ;
        RECT 12.980 69.600 13.240 69.690 ;
        RECT 12.980 69.460 13.640 69.600 ;
        RECT 12.980 69.370 13.240 69.460 ;
        RECT 11.600 68.690 11.860 69.010 ;
        RECT 10.680 67.330 10.940 67.650 ;
        RECT 11.660 67.310 11.800 68.690 ;
        RECT 11.600 66.990 11.860 67.310 ;
        RECT 10.680 66.650 10.940 66.970 ;
        RECT 10.220 62.910 10.480 63.230 ;
        RECT 9.760 60.870 10.020 61.190 ;
        RECT 9.750 59.995 10.030 60.365 ;
        RECT 9.820 59.490 9.960 59.995 ;
        RECT 9.760 59.170 10.020 59.490 ;
        RECT 9.750 58.635 10.030 59.005 ;
        RECT 9.760 58.490 10.020 58.635 ;
        RECT 9.760 57.470 10.020 57.790 ;
        RECT 9.290 55.915 9.570 56.285 ;
        RECT 9.820 55.750 9.960 57.470 ;
        RECT 10.280 56.965 10.420 62.910 ;
        RECT 10.740 60.365 10.880 66.650 ;
        RECT 11.140 66.310 11.400 66.630 ;
        RECT 11.200 62.210 11.340 66.310 ;
        RECT 12.120 66.290 12.260 69.030 ;
        RECT 12.580 68.950 13.180 69.090 ;
        RECT 13.500 69.010 13.640 69.460 ;
        RECT 12.520 68.350 12.780 68.670 ;
        RECT 12.580 66.630 12.720 68.350 ;
        RECT 12.520 66.310 12.780 66.630 ;
        RECT 12.060 65.970 12.320 66.290 ;
        RECT 11.600 65.630 11.860 65.950 ;
        RECT 11.140 61.890 11.400 62.210 ;
        RECT 11.140 60.870 11.400 61.190 ;
        RECT 10.670 59.995 10.950 60.365 ;
        RECT 10.680 59.170 10.940 59.490 ;
        RECT 10.210 56.595 10.490 56.965 ;
        RECT 9.760 55.430 10.020 55.750 ;
        RECT 9.820 51.330 9.960 55.430 ;
        RECT 10.740 55.070 10.880 59.170 ;
        RECT 10.680 54.750 10.940 55.070 ;
        RECT 10.210 53.195 10.490 53.565 ;
        RECT 10.220 53.050 10.480 53.195 ;
        RECT 10.680 53.050 10.940 53.370 ;
        RECT 9.760 51.010 10.020 51.330 ;
        RECT 9.300 49.990 9.560 50.310 ;
        RECT 7.980 48.230 8.580 48.370 ;
        RECT 7.980 45.210 8.120 48.230 ;
        RECT 9.360 47.930 9.500 49.990 ;
        RECT 9.760 49.310 10.020 49.630 ;
        RECT 9.300 47.610 9.560 47.930 ;
        RECT 8.380 46.590 8.640 46.910 ;
        RECT 7.920 44.890 8.180 45.210 ;
        RECT 7.980 34.670 8.120 44.890 ;
        RECT 8.440 44.530 8.580 46.590 ;
        RECT 8.840 44.550 9.100 44.870 ;
        RECT 8.380 44.210 8.640 44.530 ;
        RECT 8.900 40.450 9.040 44.550 ;
        RECT 8.840 40.130 9.100 40.450 ;
        RECT 8.840 38.430 9.100 38.750 ;
        RECT 7.920 34.350 8.180 34.670 ;
        RECT 8.900 29.570 9.040 38.430 ;
        RECT 9.820 37.730 9.960 49.310 ;
        RECT 10.740 46.910 10.880 53.050 ;
        RECT 11.200 49.970 11.340 60.870 ;
        RECT 11.660 58.130 11.800 65.630 ;
        RECT 12.120 60.850 12.260 65.970 ;
        RECT 12.510 65.435 12.790 65.805 ;
        RECT 12.580 64.250 12.720 65.435 ;
        RECT 12.520 63.930 12.780 64.250 ;
        RECT 12.060 60.530 12.320 60.850 ;
        RECT 11.600 57.810 11.860 58.130 ;
        RECT 11.660 56.430 11.800 57.810 ;
        RECT 11.600 56.110 11.860 56.430 ;
        RECT 11.600 55.090 11.860 55.410 ;
        RECT 11.140 49.650 11.400 49.970 ;
        RECT 11.660 47.840 11.800 55.090 ;
        RECT 12.120 48.370 12.260 60.530 ;
        RECT 12.580 55.410 12.720 63.930 ;
        RECT 13.040 63.820 13.180 68.950 ;
        RECT 13.440 68.690 13.700 69.010 ;
        RECT 13.500 66.970 13.640 68.690 ;
        RECT 13.440 66.650 13.700 66.970 ;
        RECT 13.440 64.445 13.700 64.590 ;
        RECT 13.430 64.075 13.710 64.445 ;
        RECT 13.440 63.820 13.700 63.910 ;
        RECT 13.040 63.680 13.700 63.820 ;
        RECT 13.440 63.590 13.700 63.680 ;
        RECT 13.440 60.530 13.700 60.850 ;
        RECT 13.500 59.150 13.640 60.530 ;
        RECT 13.440 58.830 13.700 59.150 ;
        RECT 12.970 57.275 13.250 57.645 ;
        RECT 13.040 56.770 13.180 57.275 ;
        RECT 12.980 56.450 13.240 56.770 ;
        RECT 13.500 55.750 13.640 58.830 ;
        RECT 13.440 55.430 13.700 55.750 ;
        RECT 12.520 55.090 12.780 55.410 ;
        RECT 13.500 54.050 13.640 55.430 ;
        RECT 13.440 53.730 13.700 54.050 ;
        RECT 12.520 53.050 12.780 53.370 ;
        RECT 12.980 53.050 13.240 53.370 ;
        RECT 12.580 50.990 12.720 53.050 ;
        RECT 13.040 52.350 13.180 53.050 ;
        RECT 12.980 52.030 13.240 52.350 ;
        RECT 12.520 50.670 12.780 50.990 ;
        RECT 13.500 50.650 13.640 53.730 ;
        RECT 13.960 53.370 14.100 73.790 ;
        RECT 14.420 61.725 14.560 75.150 ;
        RECT 15.340 75.130 15.480 76.995 ;
        RECT 15.800 76.685 15.940 80.250 ;
        RECT 15.730 76.315 16.010 76.685 ;
        RECT 15.730 75.635 16.010 76.005 ;
        RECT 15.280 74.810 15.540 75.130 ;
        RECT 15.800 73.000 15.940 75.635 ;
        RECT 15.340 72.860 15.940 73.000 ;
        RECT 15.340 72.410 15.480 72.860 ;
        RECT 15.280 72.090 15.540 72.410 ;
        RECT 15.740 72.090 16.000 72.410 ;
        RECT 15.800 71.925 15.940 72.090 ;
        RECT 15.280 71.410 15.540 71.730 ;
        RECT 15.730 71.555 16.010 71.925 ;
        RECT 15.340 69.885 15.480 71.410 ;
        RECT 14.820 69.370 15.080 69.690 ;
        RECT 15.270 69.515 15.550 69.885 ;
        RECT 14.880 66.630 15.020 69.370 ;
        RECT 15.740 68.350 16.000 68.670 ;
        RECT 15.800 66.630 15.940 68.350 ;
        RECT 14.820 66.485 15.080 66.630 ;
        RECT 14.810 66.115 15.090 66.485 ;
        RECT 15.740 66.310 16.000 66.630 ;
        RECT 14.880 64.930 15.020 66.115 ;
        RECT 15.280 65.630 15.540 65.950 ;
        RECT 14.820 64.610 15.080 64.930 ;
        RECT 14.350 61.355 14.630 61.725 ;
        RECT 14.820 61.210 15.080 61.530 ;
        RECT 14.880 60.930 15.020 61.210 ;
        RECT 15.340 61.190 15.480 65.630 ;
        RECT 15.740 61.550 16.000 61.870 ;
        RECT 14.420 60.790 15.020 60.930 ;
        RECT 15.280 60.870 15.540 61.190 ;
        RECT 13.900 53.050 14.160 53.370 ;
        RECT 13.900 51.010 14.160 51.330 ;
        RECT 13.440 50.330 13.700 50.650 ;
        RECT 12.120 48.230 12.720 48.370 ;
        RECT 12.060 47.840 12.320 47.930 ;
        RECT 11.660 47.700 12.320 47.840 ;
        RECT 12.060 47.610 12.320 47.700 ;
        RECT 11.140 46.930 11.400 47.250 ;
        RECT 10.680 46.590 10.940 46.910 ;
        RECT 10.220 44.890 10.480 45.210 ;
        RECT 10.280 43.170 10.420 44.890 ;
        RECT 10.680 44.550 10.940 44.870 ;
        RECT 10.220 42.850 10.480 43.170 ;
        RECT 10.740 42.830 10.880 44.550 ;
        RECT 11.200 43.170 11.340 46.930 ;
        RECT 12.120 46.910 12.260 47.610 ;
        RECT 12.060 46.590 12.320 46.910 ;
        RECT 11.140 42.850 11.400 43.170 ;
        RECT 10.680 42.510 10.940 42.830 ;
        RECT 9.760 37.410 10.020 37.730 ;
        RECT 9.760 35.710 10.020 36.030 ;
        RECT 9.820 35.010 9.960 35.710 ;
        RECT 9.760 34.690 10.020 35.010 ;
        RECT 10.220 33.900 10.480 33.990 ;
        RECT 10.740 33.900 10.880 42.510 ;
        RECT 11.200 39.770 11.340 42.850 ;
        RECT 11.600 41.830 11.860 42.150 ;
        RECT 12.060 41.830 12.320 42.150 ;
        RECT 11.140 39.450 11.400 39.770 ;
        RECT 11.660 38.750 11.800 41.830 ;
        RECT 12.120 39.770 12.260 41.830 ;
        RECT 12.060 39.450 12.320 39.770 ;
        RECT 11.600 38.430 11.860 38.750 ;
        RECT 12.120 36.710 12.260 39.450 ;
        RECT 12.060 36.390 12.320 36.710 ;
        RECT 12.580 34.410 12.720 48.230 ;
        RECT 12.980 47.610 13.240 47.930 ;
        RECT 10.220 33.760 10.880 33.900 ;
        RECT 10.220 33.670 10.480 33.760 ;
        RECT 10.740 31.610 10.880 33.760 ;
        RECT 11.200 34.270 12.720 34.410 ;
        RECT 10.680 31.290 10.940 31.610 ;
        RECT 10.220 30.610 10.480 30.930 ;
        RECT 8.840 29.250 9.100 29.570 ;
        RECT 10.280 29.230 10.420 30.610 ;
        RECT 10.220 28.910 10.480 29.230 ;
        RECT 4.690 27.355 4.970 27.725 ;
        RECT 5.160 27.550 5.420 27.870 ;
        RECT 11.200 26.850 11.340 34.270 ;
        RECT 12.060 31.970 12.320 32.290 ;
        RECT 12.120 28.890 12.260 31.970 ;
        RECT 13.040 31.010 13.180 47.610 ;
        RECT 13.430 47.075 13.710 47.445 ;
        RECT 13.440 46.930 13.700 47.075 ;
        RECT 13.960 44.610 14.100 51.010 ;
        RECT 14.420 45.210 14.560 60.790 ;
        RECT 14.820 60.190 15.080 60.510 ;
        RECT 14.880 59.005 15.020 60.190 ;
        RECT 15.340 59.490 15.480 60.870 ;
        RECT 15.280 59.170 15.540 59.490 ;
        RECT 14.810 58.890 15.090 59.005 ;
        RECT 14.810 58.750 15.480 58.890 ;
        RECT 14.810 58.635 15.090 58.750 ;
        RECT 14.810 57.955 15.090 58.325 ;
        RECT 14.880 50.990 15.020 57.955 ;
        RECT 15.340 55.750 15.480 58.750 ;
        RECT 15.800 58.130 15.940 61.550 ;
        RECT 15.740 57.810 16.000 58.130 ;
        RECT 15.800 56.090 15.940 57.810 ;
        RECT 16.260 56.770 16.400 92.570 ;
        RECT 18.950 91.955 19.230 92.325 ;
        RECT 18.040 82.290 18.300 82.610 ;
        RECT 16.660 81.950 16.920 82.270 ;
        RECT 16.720 80.570 16.860 81.950 ;
        RECT 18.100 80.570 18.240 82.290 ;
        RECT 16.660 80.250 16.920 80.570 ;
        RECT 17.120 80.250 17.380 80.570 ;
        RECT 18.040 80.250 18.300 80.570 ;
        RECT 17.180 79.550 17.320 80.250 ;
        RECT 17.120 79.230 17.380 79.550 ;
        RECT 17.180 77.850 17.320 79.230 ;
        RECT 17.580 78.210 17.840 78.530 ;
        RECT 17.120 77.530 17.380 77.850 ;
        RECT 17.110 72.235 17.390 72.605 ;
        RECT 17.180 72.070 17.320 72.235 ;
        RECT 17.120 71.750 17.380 72.070 ;
        RECT 16.660 71.070 16.920 71.390 ;
        RECT 16.720 70.370 16.860 71.070 ;
        RECT 17.110 70.875 17.390 71.245 ;
        RECT 16.660 70.050 16.920 70.370 ;
        RECT 16.660 69.030 16.920 69.350 ;
        RECT 16.720 67.165 16.860 69.030 ;
        RECT 17.180 68.670 17.320 70.875 ;
        RECT 17.120 68.350 17.380 68.670 ;
        RECT 17.120 67.330 17.380 67.650 ;
        RECT 16.650 66.795 16.930 67.165 ;
        RECT 16.720 65.805 16.860 66.795 ;
        RECT 16.650 65.435 16.930 65.805 ;
        RECT 16.650 64.755 16.930 65.125 ;
        RECT 16.720 64.250 16.860 64.755 ;
        RECT 16.660 63.930 16.920 64.250 ;
        RECT 16.720 59.490 16.860 63.930 ;
        RECT 17.180 60.930 17.320 67.330 ;
        RECT 17.640 67.220 17.780 78.210 ;
        RECT 18.040 73.790 18.300 74.110 ;
        RECT 18.100 69.010 18.240 73.790 ;
        RECT 18.500 69.205 18.760 69.350 ;
        RECT 18.040 68.690 18.300 69.010 ;
        RECT 18.490 68.835 18.770 69.205 ;
        RECT 19.020 68.580 19.160 91.955 ;
        RECT 19.480 78.045 19.620 92.570 ;
        RECT 20.330 86.515 20.610 86.885 ;
        RECT 19.880 83.310 20.140 83.630 ;
        RECT 19.940 79.890 20.080 83.310 ;
        RECT 20.400 81.250 20.540 86.515 ;
        RECT 22.700 84.845 22.840 92.570 ;
        RECT 22.630 84.475 22.910 84.845 ;
        RECT 24.020 84.670 24.280 84.990 ;
        RECT 23.100 83.650 23.360 83.970 ;
        RECT 22.640 82.630 22.900 82.950 ;
        RECT 21.720 82.290 21.980 82.610 ;
        RECT 20.340 80.930 20.600 81.250 ;
        RECT 21.780 80.570 21.920 82.290 ;
        RECT 22.180 80.930 22.440 81.250 ;
        RECT 21.720 80.250 21.980 80.570 ;
        RECT 22.240 80.230 22.380 80.930 ;
        RECT 22.700 80.570 22.840 82.630 ;
        RECT 22.640 80.250 22.900 80.570 ;
        RECT 21.260 79.910 21.520 80.230 ;
        RECT 22.180 79.910 22.440 80.230 ;
        RECT 19.880 79.570 20.140 79.890 ;
        RECT 21.320 79.550 21.460 79.910 ;
        RECT 21.260 79.230 21.520 79.550 ;
        RECT 21.070 78.695 22.610 79.065 ;
        RECT 19.410 77.675 19.690 78.045 ;
        RECT 21.720 77.530 21.980 77.850 ;
        RECT 22.170 77.675 22.450 78.045 ;
        RECT 19.420 77.190 19.680 77.510 ;
        RECT 21.260 77.190 21.520 77.510 ;
        RECT 18.560 68.440 19.160 68.580 ;
        RECT 18.040 67.220 18.300 67.310 ;
        RECT 17.640 67.080 18.300 67.220 ;
        RECT 18.040 66.990 18.300 67.080 ;
        RECT 17.570 65.435 17.850 65.805 ;
        RECT 17.640 64.930 17.780 65.435 ;
        RECT 17.580 64.610 17.840 64.930 ;
        RECT 18.100 63.650 18.240 66.990 ;
        RECT 18.560 64.250 18.700 68.440 ;
        RECT 18.960 66.990 19.220 67.310 ;
        RECT 18.500 63.930 18.760 64.250 ;
        RECT 18.100 63.510 18.700 63.650 ;
        RECT 19.020 63.570 19.160 66.990 ;
        RECT 18.560 62.210 18.700 63.510 ;
        RECT 18.960 63.250 19.220 63.570 ;
        RECT 18.950 62.715 19.230 63.085 ;
        RECT 18.500 61.890 18.760 62.210 ;
        RECT 19.020 61.870 19.160 62.715 ;
        RECT 18.960 61.550 19.220 61.870 ;
        RECT 17.180 60.790 19.160 60.930 ;
        RECT 16.660 59.170 16.920 59.490 ;
        RECT 16.650 58.635 16.930 59.005 ;
        RECT 16.200 56.450 16.460 56.770 ;
        RECT 15.740 55.770 16.000 56.090 ;
        RECT 15.280 55.605 15.540 55.750 ;
        RECT 15.270 55.235 15.550 55.605 ;
        RECT 16.720 55.320 16.860 58.635 ;
        RECT 16.260 55.180 16.860 55.320 ;
        RECT 15.270 53.875 15.550 54.245 ;
        RECT 15.280 53.730 15.540 53.875 ;
        RECT 16.260 52.350 16.400 55.180 ;
        RECT 16.650 54.555 16.930 54.925 ;
        RECT 16.720 53.370 16.860 54.555 ;
        RECT 16.660 53.050 16.920 53.370 ;
        RECT 17.180 53.030 17.320 60.790 ;
        RECT 18.500 60.190 18.760 60.510 ;
        RECT 18.560 59.060 18.700 60.190 ;
        RECT 19.020 59.400 19.160 60.790 ;
        RECT 19.480 60.510 19.620 77.190 ;
        RECT 20.340 76.850 20.600 77.170 ;
        RECT 19.880 76.510 20.140 76.830 ;
        RECT 19.940 67.845 20.080 76.510 ;
        RECT 20.400 75.130 20.540 76.850 ;
        RECT 20.800 76.510 21.060 76.830 ;
        RECT 21.320 76.685 21.460 77.190 ;
        RECT 20.340 74.810 20.600 75.130 ;
        RECT 20.860 74.020 21.000 76.510 ;
        RECT 21.250 76.315 21.530 76.685 ;
        RECT 21.780 76.005 21.920 77.530 ;
        RECT 22.240 77.510 22.380 77.675 ;
        RECT 22.180 77.190 22.440 77.510 ;
        RECT 21.260 75.490 21.520 75.810 ;
        RECT 21.710 75.635 21.990 76.005 ;
        RECT 23.160 75.810 23.300 83.650 ;
        RECT 23.550 80.395 23.830 80.765 ;
        RECT 21.320 75.130 21.460 75.490 ;
        RECT 21.780 75.130 21.920 75.635 ;
        RECT 22.640 75.490 22.900 75.810 ;
        RECT 23.100 75.490 23.360 75.810 ;
        RECT 22.700 75.210 22.840 75.490 ;
        RECT 23.620 75.210 23.760 80.395 ;
        RECT 24.080 77.850 24.220 84.670 ;
        RECT 25.920 83.485 26.060 92.570 ;
        RECT 29.140 86.885 29.280 92.570 ;
        RECT 32.360 91.110 32.500 92.570 ;
        RECT 32.300 90.790 32.560 91.110 ;
        RECT 29.070 86.515 29.350 86.885 ;
        RECT 25.850 83.115 26.130 83.485 ;
        RECT 26.320 82.970 26.580 83.290 ;
        RECT 24.370 81.415 25.910 81.785 ;
        RECT 26.380 80.570 26.520 82.970 ;
        RECT 34.600 82.290 34.860 82.610 ;
        RECT 31.380 80.590 31.640 80.910 ;
        RECT 24.940 80.250 25.200 80.570 ;
        RECT 26.320 80.250 26.580 80.570 ;
        RECT 28.160 80.250 28.420 80.570 ;
        RECT 24.480 79.910 24.740 80.230 ;
        RECT 24.020 77.530 24.280 77.850 ;
        RECT 24.540 77.080 24.680 79.910 ;
        RECT 25.000 78.725 25.140 80.250 ;
        RECT 26.780 79.570 27.040 79.890 ;
        RECT 24.930 78.355 25.210 78.725 ;
        RECT 25.860 77.080 26.120 77.170 ;
        RECT 24.540 76.940 26.120 77.080 ;
        RECT 25.860 76.850 26.120 76.940 ;
        RECT 24.370 75.975 25.910 76.345 ;
        RECT 24.940 75.720 25.200 75.810 ;
        RECT 21.260 74.810 21.520 75.130 ;
        RECT 21.720 74.810 21.980 75.130 ;
        RECT 22.700 75.070 23.760 75.210 ;
        RECT 24.080 75.580 25.600 75.720 ;
        RECT 23.560 74.360 23.820 74.450 ;
        RECT 24.080 74.360 24.220 75.580 ;
        RECT 24.940 75.490 25.200 75.580 ;
        RECT 25.460 75.325 25.600 75.580 ;
        RECT 25.860 75.490 26.120 75.810 ;
        RECT 24.470 74.955 24.750 75.325 ;
        RECT 25.390 74.955 25.670 75.325 ;
        RECT 24.540 74.700 24.680 74.955 ;
        RECT 25.920 74.700 26.060 75.490 ;
        RECT 24.540 74.560 26.060 74.700 ;
        RECT 23.560 74.220 24.220 74.360 ;
        RECT 26.310 74.275 26.590 74.645 ;
        RECT 23.560 74.130 23.820 74.220 ;
        RECT 26.320 74.130 26.580 74.275 ;
        RECT 20.400 73.880 21.000 74.020 ;
        RECT 20.400 71.245 20.540 73.880 ;
        RECT 21.070 73.255 22.610 73.625 ;
        RECT 23.550 73.595 23.830 73.965 ;
        RECT 24.940 73.790 25.200 74.110 ;
        RECT 23.620 72.070 23.760 73.595 ;
        RECT 25.000 72.070 25.140 73.790 ;
        RECT 26.840 72.750 26.980 79.570 ;
        RECT 27.230 79.035 27.510 79.405 ;
        RECT 27.700 79.230 27.960 79.550 ;
        RECT 27.300 78.530 27.440 79.035 ;
        RECT 27.760 78.530 27.900 79.230 ;
        RECT 27.240 78.210 27.500 78.530 ;
        RECT 27.700 78.210 27.960 78.530 ;
        RECT 27.700 76.850 27.960 77.170 ;
        RECT 27.760 75.130 27.900 76.850 ;
        RECT 27.700 75.040 27.960 75.130 ;
        RECT 27.300 74.900 27.960 75.040 ;
        RECT 25.860 72.430 26.120 72.750 ;
        RECT 26.780 72.430 27.040 72.750 ;
        RECT 21.720 71.750 21.980 72.070 ;
        RECT 23.100 71.750 23.360 72.070 ;
        RECT 23.560 71.750 23.820 72.070 ;
        RECT 24.940 71.750 25.200 72.070 ;
        RECT 20.330 70.875 20.610 71.245 ;
        RECT 21.780 70.565 21.920 71.750 ;
        RECT 21.710 70.195 21.990 70.565 ;
        RECT 20.340 69.600 20.600 69.690 ;
        RECT 20.340 69.460 21.000 69.600 ;
        RECT 20.340 69.370 20.600 69.460 ;
        RECT 20.860 69.205 21.000 69.460 ;
        RECT 21.260 69.370 21.520 69.690 ;
        RECT 22.170 69.515 22.450 69.885 ;
        RECT 22.640 69.710 22.900 70.030 ;
        RECT 22.180 69.370 22.440 69.515 ;
        RECT 20.340 68.690 20.600 69.010 ;
        RECT 20.790 68.835 21.070 69.205 ;
        RECT 21.320 69.010 21.460 69.370 ;
        RECT 22.700 69.260 22.840 69.710 ;
        RECT 23.160 69.590 23.300 71.750 ;
        RECT 25.920 71.730 26.060 72.430 ;
        RECT 27.300 71.810 27.440 74.900 ;
        RECT 27.700 74.810 27.960 74.900 ;
        RECT 27.700 74.130 27.960 74.450 ;
        RECT 27.760 73.090 27.900 74.130 ;
        RECT 28.220 74.110 28.360 80.250 ;
        RECT 29.080 79.910 29.340 80.230 ;
        RECT 29.540 79.910 29.800 80.230 ;
        RECT 30.460 79.910 30.720 80.230 ;
        RECT 30.920 79.910 31.180 80.230 ;
        RECT 28.620 74.470 28.880 74.790 ;
        RECT 28.160 73.790 28.420 74.110 ;
        RECT 27.700 72.770 27.960 73.090 ;
        RECT 28.680 72.410 28.820 74.470 ;
        RECT 28.620 72.090 28.880 72.410 ;
        RECT 28.680 71.810 28.820 72.090 ;
        RECT 25.860 71.410 26.120 71.730 ;
        RECT 26.780 71.410 27.040 71.730 ;
        RECT 27.300 71.670 27.900 71.810 ;
        RECT 28.220 71.730 28.820 71.810 ;
        RECT 23.560 71.070 23.820 71.390 ;
        RECT 23.620 69.940 23.760 71.070 ;
        RECT 24.370 70.535 25.910 70.905 ;
        RECT 26.840 70.565 26.980 71.410 ;
        RECT 27.240 71.070 27.500 71.390 ;
        RECT 26.770 70.195 27.050 70.565 ;
        RECT 23.620 69.800 24.680 69.940 ;
        RECT 23.160 69.450 24.220 69.590 ;
        RECT 22.700 69.120 23.300 69.260 ;
        RECT 21.260 68.690 21.520 69.010 ;
        RECT 19.870 67.475 20.150 67.845 ;
        RECT 20.400 66.630 20.540 68.690 ;
        RECT 21.070 67.815 22.610 68.185 ;
        RECT 22.180 67.330 22.440 67.650 ;
        RECT 20.800 66.650 21.060 66.970 ;
        RECT 20.340 66.310 20.600 66.630 ;
        RECT 19.880 65.630 20.140 65.950 ;
        RECT 20.340 65.630 20.600 65.950 ;
        RECT 19.940 64.590 20.080 65.630 ;
        RECT 20.400 64.590 20.540 65.630 ;
        RECT 19.880 64.270 20.140 64.590 ;
        RECT 20.340 64.270 20.600 64.590 ;
        RECT 20.860 64.250 21.000 66.650 ;
        RECT 22.240 66.630 22.380 67.330 ;
        RECT 22.180 66.310 22.440 66.630 ;
        RECT 22.640 66.485 22.900 66.630 ;
        RECT 21.260 65.630 21.520 65.950 ;
        RECT 22.240 65.805 22.380 66.310 ;
        RECT 22.630 66.115 22.910 66.485 ;
        RECT 23.160 66.290 23.300 69.120 ;
        RECT 23.560 68.350 23.820 68.670 ;
        RECT 23.620 67.310 23.760 68.350 ;
        RECT 23.560 66.990 23.820 67.310 ;
        RECT 23.100 65.970 23.360 66.290 ;
        RECT 23.550 66.115 23.830 66.485 ;
        RECT 20.800 63.930 21.060 64.250 ;
        RECT 19.880 63.250 20.140 63.570 ;
        RECT 19.940 61.610 20.080 63.250 ;
        RECT 20.340 62.910 20.600 63.230 ;
        RECT 21.320 63.140 21.460 65.630 ;
        RECT 22.170 65.435 22.450 65.805 ;
        RECT 23.160 65.125 23.300 65.970 ;
        RECT 22.180 64.610 22.440 64.930 ;
        RECT 23.090 64.755 23.370 65.125 ;
        RECT 22.240 64.250 22.380 64.610 ;
        RECT 23.620 64.250 23.760 66.115 ;
        RECT 22.180 63.930 22.440 64.250 ;
        RECT 23.560 63.930 23.820 64.250 ;
        RECT 23.550 63.395 23.830 63.765 ;
        RECT 23.560 63.250 23.820 63.395 ;
        RECT 21.320 63.000 23.300 63.140 ;
        RECT 20.400 62.120 20.540 62.910 ;
        RECT 21.070 62.375 22.610 62.745 ;
        RECT 20.400 61.980 21.000 62.120 ;
        RECT 19.940 61.470 20.540 61.610 ;
        RECT 20.860 61.530 21.000 61.980 ;
        RECT 19.880 60.870 20.140 61.190 ;
        RECT 19.420 60.190 19.680 60.510 ;
        RECT 19.940 60.365 20.080 60.870 ;
        RECT 19.870 59.995 20.150 60.365 ;
        RECT 19.020 59.260 20.080 59.400 ;
        RECT 18.560 58.920 19.620 59.060 ;
        RECT 18.500 57.810 18.760 58.130 ;
        RECT 18.960 57.810 19.220 58.130 ;
        RECT 18.030 56.595 18.310 56.965 ;
        RECT 17.570 55.915 17.850 56.285 ;
        RECT 17.640 54.050 17.780 55.915 ;
        RECT 17.580 53.730 17.840 54.050 ;
        RECT 18.100 53.370 18.240 56.595 ;
        RECT 18.560 55.070 18.700 57.810 ;
        RECT 19.020 56.965 19.160 57.810 ;
        RECT 18.950 56.595 19.230 56.965 ;
        RECT 19.480 55.750 19.620 58.920 ;
        RECT 19.940 58.810 20.080 59.260 ;
        RECT 19.880 58.490 20.140 58.810 ;
        RECT 20.400 58.380 20.540 61.470 ;
        RECT 20.800 61.440 21.060 61.530 ;
        RECT 20.800 61.300 21.460 61.440 ;
        RECT 22.170 61.355 22.450 61.725 ;
        RECT 20.800 61.210 21.060 61.300 ;
        RECT 20.790 60.675 21.070 61.045 ;
        RECT 20.800 60.530 21.060 60.675 ;
        RECT 20.790 59.315 21.070 59.685 ;
        RECT 20.860 58.810 21.000 59.315 ;
        RECT 20.800 58.490 21.060 58.810 ;
        RECT 21.320 58.470 21.460 61.300 ;
        RECT 21.720 60.365 21.980 60.510 ;
        RECT 21.710 59.995 21.990 60.365 ;
        RECT 22.240 59.570 22.380 61.355 ;
        RECT 23.160 61.190 23.300 63.000 ;
        RECT 24.080 61.530 24.220 69.450 ;
        RECT 24.540 68.670 24.680 69.800 ;
        RECT 25.400 69.600 25.660 69.690 ;
        RECT 26.310 69.600 26.590 69.885 ;
        RECT 25.400 69.460 26.060 69.600 ;
        RECT 26.310 69.515 26.980 69.600 ;
        RECT 25.400 69.370 25.660 69.460 ;
        RECT 25.920 69.220 26.060 69.460 ;
        RECT 26.320 69.460 26.980 69.515 ;
        RECT 26.320 69.370 26.580 69.460 ;
        RECT 25.920 69.080 26.520 69.220 ;
        RECT 26.380 68.670 26.520 69.080 ;
        RECT 24.480 68.350 24.740 68.670 ;
        RECT 26.320 68.350 26.580 68.670 ;
        RECT 26.840 67.310 26.980 69.460 ;
        RECT 26.310 66.795 26.590 67.165 ;
        RECT 26.780 66.990 27.040 67.310 ;
        RECT 25.860 66.540 26.120 66.630 ;
        RECT 25.000 66.400 26.120 66.540 ;
        RECT 25.000 65.950 25.140 66.400 ;
        RECT 25.860 66.310 26.120 66.400 ;
        RECT 26.380 66.200 26.520 66.795 ;
        RECT 26.380 66.060 26.980 66.200 ;
        RECT 24.940 65.630 25.200 65.950 ;
        RECT 25.860 65.860 26.120 65.950 ;
        RECT 25.860 65.720 26.520 65.860 ;
        RECT 25.860 65.630 26.120 65.720 ;
        RECT 24.370 65.095 25.910 65.465 ;
        RECT 26.380 65.125 26.520 65.720 ;
        RECT 25.400 64.840 25.660 64.930 ;
        RECT 25.400 64.700 26.060 64.840 ;
        RECT 26.310 64.755 26.590 65.125 ;
        RECT 25.400 64.610 25.660 64.700 ;
        RECT 25.920 64.500 26.060 64.700 ;
        RECT 26.840 64.500 26.980 66.060 ;
        RECT 25.920 64.360 26.980 64.500 ;
        RECT 24.480 63.930 24.740 64.250 ;
        RECT 24.540 63.085 24.680 63.930 ;
        RECT 27.300 63.480 27.440 71.070 ;
        RECT 27.760 69.885 27.900 71.670 ;
        RECT 28.160 71.670 28.820 71.730 ;
        RECT 28.160 71.410 28.420 71.670 ;
        RECT 28.620 71.070 28.880 71.390 ;
        RECT 29.140 71.245 29.280 79.910 ;
        RECT 29.600 75.325 29.740 79.910 ;
        RECT 30.000 76.510 30.260 76.830 ;
        RECT 30.520 76.685 30.660 79.910 ;
        RECT 30.980 77.510 31.120 79.910 ;
        RECT 30.920 77.190 31.180 77.510 ;
        RECT 29.530 74.955 29.810 75.325 ;
        RECT 30.060 75.130 30.200 76.510 ;
        RECT 30.450 76.315 30.730 76.685 ;
        RECT 30.920 76.510 31.180 76.830 ;
        RECT 30.980 75.470 31.120 76.510 ;
        RECT 30.920 75.150 31.180 75.470 ;
        RECT 30.000 74.810 30.260 75.130 ;
        RECT 29.540 73.790 29.800 74.110 ;
        RECT 28.680 70.370 28.820 71.070 ;
        RECT 29.070 70.875 29.350 71.245 ;
        RECT 28.620 70.050 28.880 70.370 ;
        RECT 27.690 69.515 27.970 69.885 ;
        RECT 29.080 69.370 29.340 69.690 ;
        RECT 27.700 69.030 27.960 69.350 ;
        RECT 28.160 69.030 28.420 69.350 ;
        RECT 27.760 67.845 27.900 69.030 ;
        RECT 27.690 67.475 27.970 67.845 ;
        RECT 28.220 66.290 28.360 69.030 ;
        RECT 29.140 67.310 29.280 69.370 ;
        RECT 29.080 66.990 29.340 67.310 ;
        RECT 28.620 66.650 28.880 66.970 ;
        RECT 28.160 65.970 28.420 66.290 ;
        RECT 28.680 64.250 28.820 66.650 ;
        RECT 29.600 65.690 29.740 73.790 ;
        RECT 30.060 66.970 30.200 74.810 ;
        RECT 30.460 74.130 30.720 74.450 ;
        RECT 30.520 72.070 30.660 74.130 ;
        RECT 30.920 73.790 31.180 74.110 ;
        RECT 30.460 71.750 30.720 72.070 ;
        RECT 30.450 70.875 30.730 71.245 ;
        RECT 30.000 66.650 30.260 66.970 ;
        RECT 29.140 65.550 29.740 65.690 ;
        RECT 28.160 63.930 28.420 64.250 ;
        RECT 28.620 63.930 28.880 64.250 ;
        RECT 28.220 63.765 28.360 63.930 ;
        RECT 25.460 63.340 27.440 63.480 ;
        RECT 28.150 63.395 28.430 63.765 ;
        RECT 24.470 62.715 24.750 63.085 ;
        RECT 24.930 62.035 25.210 62.405 ;
        RECT 24.020 61.210 24.280 61.530 ;
        RECT 23.100 60.870 23.360 61.190 ;
        RECT 25.000 60.510 25.140 62.035 ;
        RECT 25.460 60.930 25.600 63.340 ;
        RECT 29.140 63.230 29.280 65.550 ;
        RECT 29.990 64.755 30.270 65.125 ;
        RECT 30.520 64.930 30.660 70.875 ;
        RECT 30.980 68.670 31.120 73.790 ;
        RECT 31.440 71.245 31.580 80.590 ;
        RECT 33.220 80.250 33.480 80.570 ;
        RECT 32.750 77.675 33.030 78.045 ;
        RECT 32.820 72.605 32.960 77.675 ;
        RECT 33.280 75.130 33.420 80.250 ;
        RECT 34.140 78.210 34.400 78.530 ;
        RECT 33.680 77.530 33.940 77.850 ;
        RECT 33.220 74.810 33.480 75.130 ;
        RECT 32.300 72.090 32.560 72.410 ;
        RECT 32.750 72.235 33.030 72.605 ;
        RECT 33.740 72.410 33.880 77.530 ;
        RECT 34.200 75.810 34.340 78.210 ;
        RECT 34.140 75.490 34.400 75.810 ;
        RECT 34.140 74.470 34.400 74.790 ;
        RECT 34.200 72.750 34.340 74.470 ;
        RECT 34.140 72.430 34.400 72.750 ;
        RECT 31.370 70.875 31.650 71.245 ;
        RECT 32.360 69.350 32.500 72.090 ;
        RECT 32.300 69.260 32.560 69.350 ;
        RECT 31.900 69.120 32.560 69.260 ;
        RECT 32.820 69.205 32.960 72.235 ;
        RECT 33.680 72.090 33.940 72.410 ;
        RECT 33.680 71.410 33.940 71.730 ;
        RECT 30.920 68.350 31.180 68.670 ;
        RECT 31.380 68.350 31.640 68.670 ;
        RECT 31.440 66.630 31.580 68.350 ;
        RECT 31.380 66.310 31.640 66.630 ;
        RECT 30.920 65.970 31.180 66.290 ;
        RECT 30.980 65.805 31.120 65.970 ;
        RECT 30.910 65.435 31.190 65.805 ;
        RECT 30.060 63.570 30.200 64.755 ;
        RECT 30.460 64.610 30.720 64.930 ;
        RECT 30.460 63.930 30.720 64.250 ;
        RECT 29.540 63.250 29.800 63.570 ;
        RECT 30.000 63.250 30.260 63.570 ;
        RECT 29.080 62.910 29.340 63.230 ;
        RECT 25.860 61.890 26.120 62.210 ;
        RECT 26.310 62.170 26.590 62.405 ;
        RECT 26.310 62.035 28.820 62.170 ;
        RECT 26.380 62.030 28.820 62.035 ;
        RECT 25.920 61.725 26.060 61.890 ;
        RECT 25.850 61.355 26.130 61.725 ;
        RECT 28.160 61.550 28.420 61.870 ;
        RECT 26.780 61.440 27.040 61.530 ;
        RECT 26.780 61.300 27.900 61.440 ;
        RECT 26.780 61.210 27.040 61.300 ;
        RECT 27.760 61.100 27.900 61.300 ;
        RECT 28.220 61.100 28.360 61.550 ;
        RECT 27.755 60.960 27.900 61.100 ;
        RECT 28.200 60.960 28.360 61.100 ;
        RECT 25.460 60.790 27.440 60.930 ;
        RECT 23.090 59.995 23.370 60.365 ;
        RECT 24.020 60.190 24.280 60.510 ;
        RECT 24.940 60.190 25.200 60.510 ;
        RECT 21.780 59.490 22.380 59.570 ;
        RECT 21.720 59.430 22.380 59.490 ;
        RECT 21.720 59.170 21.980 59.430 ;
        RECT 20.400 58.240 20.600 58.380 ;
        RECT 20.460 58.040 20.600 58.240 ;
        RECT 21.260 58.150 21.520 58.470 ;
        RECT 20.400 57.900 20.600 58.040 ;
        RECT 19.870 57.275 20.150 57.645 ;
        RECT 18.950 55.235 19.230 55.605 ;
        RECT 19.420 55.430 19.680 55.750 ;
        RECT 19.940 55.490 20.080 57.275 ;
        RECT 20.400 56.000 20.540 57.900 ;
        RECT 21.070 56.935 22.610 57.305 ;
        RECT 22.640 56.450 22.900 56.770 ;
        RECT 20.800 56.000 21.060 56.090 ;
        RECT 20.400 55.860 21.060 56.000 ;
        RECT 21.250 55.915 21.530 56.285 ;
        RECT 20.800 55.770 21.060 55.860 ;
        RECT 19.940 55.350 21.000 55.490 ;
        RECT 21.320 55.410 21.460 55.915 ;
        RECT 18.500 54.750 18.760 55.070 ;
        RECT 18.040 53.050 18.300 53.370 ;
        RECT 17.120 52.710 17.380 53.030 ;
        RECT 15.280 52.030 15.540 52.350 ;
        RECT 16.200 52.030 16.460 52.350 ;
        RECT 15.340 50.990 15.480 52.030 ;
        RECT 15.730 51.155 16.010 51.525 ;
        RECT 15.800 50.990 15.940 51.155 ;
        RECT 14.820 50.670 15.080 50.990 ;
        RECT 15.280 50.845 15.540 50.990 ;
        RECT 14.360 44.890 14.620 45.210 ;
        RECT 13.960 44.470 14.560 44.610 ;
        RECT 13.440 37.070 13.700 37.390 ;
        RECT 12.580 30.870 13.180 31.010 ;
        RECT 12.060 28.570 12.320 28.890 ;
        RECT 11.140 26.530 11.400 26.850 ;
        RECT 3.780 25.510 4.040 25.830 ;
        RECT 3.840 24.325 3.980 25.510 ;
        RECT 12.060 25.060 12.320 25.150 ;
        RECT 12.580 25.060 12.720 30.870 ;
        RECT 13.500 29.570 13.640 37.070 ;
        RECT 13.900 35.710 14.160 36.030 ;
        RECT 13.960 33.990 14.100 35.710 ;
        RECT 13.900 33.670 14.160 33.990 ;
        RECT 14.420 33.220 14.560 44.470 ;
        RECT 13.960 33.080 14.560 33.220 ;
        RECT 13.440 29.250 13.700 29.570 ;
        RECT 13.960 28.970 14.100 33.080 ;
        RECT 13.500 28.890 14.100 28.970 ;
        RECT 14.360 28.910 14.620 29.230 ;
        RECT 13.440 28.830 14.100 28.890 ;
        RECT 13.440 28.570 13.700 28.830 ;
        RECT 14.420 28.550 14.560 28.910 ;
        RECT 13.900 28.230 14.160 28.550 ;
        RECT 14.360 28.230 14.620 28.550 ;
        RECT 13.960 26.510 14.100 28.230 ;
        RECT 13.900 26.190 14.160 26.510 ;
        RECT 14.420 25.490 14.560 28.230 ;
        RECT 14.360 25.170 14.620 25.490 ;
        RECT 12.060 24.920 12.720 25.060 ;
        RECT 12.060 24.830 12.320 24.920 ;
        RECT 3.770 23.955 4.050 24.325 ;
        RECT 12.120 24.130 12.260 24.830 ;
        RECT 12.060 23.810 12.320 24.130 ;
        RECT 14.880 23.450 15.020 50.670 ;
        RECT 15.270 50.475 15.550 50.845 ;
        RECT 15.740 50.670 16.000 50.990 ;
        RECT 15.340 49.630 15.480 50.475 ;
        RECT 16.260 49.970 16.400 52.030 ;
        RECT 16.200 49.650 16.460 49.970 ;
        RECT 15.280 49.310 15.540 49.630 ;
        RECT 15.340 39.850 15.480 49.310 ;
        RECT 15.730 48.435 16.010 48.805 ;
        RECT 15.800 47.250 15.940 48.435 ;
        RECT 17.180 48.270 17.320 52.710 ;
        RECT 18.040 52.370 18.300 52.690 ;
        RECT 18.100 51.330 18.240 52.370 ;
        RECT 18.040 51.010 18.300 51.330 ;
        RECT 17.120 47.950 17.380 48.270 ;
        RECT 15.740 46.930 16.000 47.250 ;
        RECT 19.020 45.290 19.160 55.235 ;
        RECT 20.860 55.070 21.000 55.350 ;
        RECT 21.260 55.090 21.520 55.410 ;
        RECT 20.800 54.750 21.060 55.070 ;
        RECT 20.330 53.875 20.610 54.245 ;
        RECT 22.700 54.050 22.840 56.450 ;
        RECT 23.160 55.410 23.300 59.995 ;
        RECT 24.080 58.040 24.220 60.190 ;
        RECT 24.370 59.655 25.910 60.025 ;
        RECT 24.480 59.170 24.740 59.490 ;
        RECT 26.310 59.315 26.590 59.685 ;
        RECT 23.620 57.900 24.220 58.040 ;
        RECT 23.620 55.750 23.760 57.900 ;
        RECT 24.010 57.275 24.290 57.645 ;
        RECT 24.080 55.750 24.220 57.275 ;
        RECT 24.540 56.770 24.680 59.170 ;
        RECT 25.860 58.890 26.120 59.150 ;
        RECT 25.460 58.830 26.120 58.890 ;
        RECT 24.940 58.720 25.200 58.810 ;
        RECT 25.460 58.750 26.060 58.830 ;
        RECT 25.460 58.720 25.600 58.750 ;
        RECT 24.940 58.580 25.600 58.720 ;
        RECT 24.940 58.490 25.200 58.580 ;
        RECT 25.860 58.150 26.120 58.470 ;
        RECT 24.940 57.810 25.200 58.130 ;
        RECT 24.480 56.450 24.740 56.770 ;
        RECT 25.000 56.430 25.140 57.810 ;
        RECT 24.940 56.110 25.200 56.430 ;
        RECT 25.920 56.090 26.060 58.150 ;
        RECT 25.860 55.770 26.120 56.090 ;
        RECT 23.560 55.430 23.820 55.750 ;
        RECT 24.020 55.430 24.280 55.750 ;
        RECT 23.100 55.090 23.360 55.410 ;
        RECT 20.400 53.370 20.540 53.875 ;
        RECT 22.640 53.730 22.900 54.050 ;
        RECT 22.180 53.390 22.440 53.710 ;
        RECT 20.340 53.050 20.600 53.370 ;
        RECT 20.330 52.515 20.610 52.885 ;
        RECT 19.420 50.670 19.680 50.990 ;
        RECT 19.480 48.370 19.620 50.670 ;
        RECT 20.400 50.650 20.540 52.515 ;
        RECT 22.240 52.350 22.380 53.390 ;
        RECT 22.180 52.030 22.440 52.350 ;
        RECT 21.070 51.495 22.610 51.865 ;
        RECT 20.340 50.330 20.600 50.650 ;
        RECT 20.800 50.165 21.060 50.310 ;
        RECT 20.790 49.795 21.070 50.165 ;
        RECT 21.260 49.990 21.520 50.310 ;
        RECT 21.720 49.990 21.980 50.310 ;
        RECT 20.340 49.310 20.600 49.630 ;
        RECT 19.480 48.230 20.080 48.370 ;
        RECT 17.580 44.890 17.840 45.210 ;
        RECT 18.560 45.150 19.160 45.290 ;
        RECT 16.200 43.870 16.460 44.190 ;
        RECT 16.260 42.490 16.400 43.870 ;
        RECT 17.640 42.490 17.780 44.890 ;
        RECT 18.040 43.870 18.300 44.190 ;
        RECT 18.100 43.170 18.240 43.870 ;
        RECT 18.040 42.850 18.300 43.170 ;
        RECT 16.200 42.170 16.460 42.490 ;
        RECT 17.580 42.400 17.840 42.490 ;
        RECT 16.720 42.260 17.840 42.400 ;
        RECT 15.340 39.710 15.940 39.850 ;
        RECT 15.280 39.110 15.540 39.430 ;
        RECT 15.340 34.330 15.480 39.110 ;
        RECT 15.280 34.010 15.540 34.330 ;
        RECT 15.800 24.130 15.940 39.710 ;
        RECT 16.720 39.430 16.860 42.260 ;
        RECT 17.580 42.170 17.840 42.260 ;
        RECT 16.660 39.110 16.920 39.430 ;
        RECT 18.560 32.290 18.700 45.150 ;
        RECT 18.960 44.550 19.220 44.870 ;
        RECT 19.020 43.170 19.160 44.550 ;
        RECT 19.940 44.190 20.080 48.230 ;
        RECT 20.400 45.800 20.540 49.310 ;
        RECT 21.320 47.930 21.460 49.990 ;
        RECT 21.260 47.610 21.520 47.930 ;
        RECT 21.780 47.840 21.920 49.990 ;
        RECT 22.640 49.650 22.900 49.970 ;
        RECT 22.180 47.840 22.440 47.930 ;
        RECT 21.780 47.700 22.440 47.840 ;
        RECT 22.180 47.610 22.440 47.700 ;
        RECT 22.700 47.330 22.840 49.650 ;
        RECT 23.160 48.610 23.300 55.090 ;
        RECT 23.620 54.980 23.760 55.430 ;
        RECT 23.620 54.840 24.220 54.980 ;
        RECT 23.560 52.710 23.820 53.030 ;
        RECT 23.100 48.290 23.360 48.610 ;
        RECT 23.620 47.590 23.760 52.710 ;
        RECT 24.080 51.330 24.220 54.840 ;
        RECT 24.370 54.215 25.910 54.585 ;
        RECT 26.380 52.690 26.520 59.315 ;
        RECT 26.780 56.110 27.040 56.430 ;
        RECT 26.840 54.925 26.980 56.110 ;
        RECT 27.300 55.750 27.440 60.790 ;
        RECT 27.755 60.420 27.895 60.960 ;
        RECT 28.200 60.760 28.340 60.960 ;
        RECT 28.200 60.620 28.360 60.760 ;
        RECT 27.755 60.280 27.900 60.420 ;
        RECT 27.760 59.005 27.900 60.280 ;
        RECT 27.690 58.635 27.970 59.005 ;
        RECT 27.690 56.595 27.970 56.965 ;
        RECT 27.700 56.450 27.960 56.595 ;
        RECT 27.240 55.430 27.500 55.750 ;
        RECT 26.770 54.555 27.050 54.925 ;
        RECT 27.700 53.050 27.960 53.370 ;
        RECT 27.760 52.690 27.900 53.050 ;
        RECT 26.320 52.370 26.580 52.690 ;
        RECT 27.700 52.370 27.960 52.690 ;
        RECT 25.850 51.835 26.130 52.205 ;
        RECT 24.020 51.010 24.280 51.330 ;
        RECT 25.920 50.310 26.060 51.835 ;
        RECT 27.230 50.475 27.510 50.845 ;
        RECT 25.390 49.795 25.670 50.165 ;
        RECT 25.860 49.990 26.120 50.310 ;
        RECT 26.320 50.165 26.580 50.310 ;
        RECT 26.310 49.795 26.590 50.165 ;
        RECT 27.300 49.970 27.440 50.475 ;
        RECT 27.760 50.310 27.900 52.370 ;
        RECT 28.220 50.730 28.360 60.620 ;
        RECT 28.680 58.210 28.820 62.030 ;
        RECT 29.600 61.725 29.740 63.250 ;
        RECT 29.080 61.210 29.340 61.530 ;
        RECT 29.530 61.355 29.810 61.725 ;
        RECT 29.140 59.685 29.280 61.210 ;
        RECT 30.000 60.870 30.260 61.190 ;
        RECT 29.540 60.190 29.800 60.510 ;
        RECT 29.070 59.315 29.350 59.685 ;
        RECT 28.680 58.070 29.280 58.210 ;
        RECT 28.620 57.470 28.880 57.790 ;
        RECT 28.680 56.430 28.820 57.470 ;
        RECT 29.140 56.965 29.280 58.070 ;
        RECT 29.070 56.595 29.350 56.965 ;
        RECT 28.620 56.110 28.880 56.430 ;
        RECT 28.620 55.430 28.880 55.750 ;
        RECT 29.080 55.430 29.340 55.750 ;
        RECT 28.680 54.050 28.820 55.430 ;
        RECT 28.620 53.730 28.880 54.050 ;
        RECT 28.610 52.515 28.890 52.885 ;
        RECT 28.680 51.330 28.820 52.515 ;
        RECT 28.620 51.010 28.880 51.330 ;
        RECT 28.220 50.590 28.820 50.730 ;
        RECT 27.700 49.990 27.960 50.310 ;
        RECT 28.160 49.990 28.420 50.310 ;
        RECT 27.240 49.880 27.500 49.970 ;
        RECT 25.460 49.630 25.600 49.795 ;
        RECT 26.840 49.740 27.500 49.880 ;
        RECT 25.400 49.310 25.660 49.630 ;
        RECT 24.370 48.775 25.910 49.145 ;
        RECT 24.480 47.610 24.740 47.930 ;
        RECT 22.700 47.190 23.300 47.330 ;
        RECT 23.560 47.270 23.820 47.590 ;
        RECT 21.070 46.055 22.610 46.425 ;
        RECT 20.400 45.660 21.460 45.800 ;
        RECT 19.880 43.870 20.140 44.190 ;
        RECT 18.960 42.850 19.220 43.170 ;
        RECT 20.800 42.570 21.060 42.830 ;
        RECT 19.940 42.510 21.060 42.570 ;
        RECT 19.940 42.490 21.000 42.510 ;
        RECT 18.960 42.170 19.220 42.490 ;
        RECT 19.880 42.430 21.000 42.490 ;
        RECT 19.880 42.170 20.140 42.430 ;
        RECT 19.020 40.110 19.160 42.170 ;
        RECT 21.320 41.470 21.460 45.660 ;
        RECT 21.720 45.230 21.980 45.550 ;
        RECT 21.780 42.490 21.920 45.230 ;
        RECT 21.720 42.170 21.980 42.490 ;
        RECT 21.260 41.150 21.520 41.470 ;
        RECT 21.070 40.615 22.610 40.985 ;
        RECT 23.160 40.450 23.300 47.190 ;
        RECT 23.620 44.870 23.760 47.270 ;
        RECT 23.560 44.550 23.820 44.870 ;
        RECT 24.540 44.610 24.680 47.610 ;
        RECT 26.320 44.890 26.580 45.210 ;
        RECT 23.100 40.130 23.360 40.450 ;
        RECT 18.960 39.790 19.220 40.110 ;
        RECT 19.020 39.430 19.160 39.790 ;
        RECT 18.960 39.110 19.220 39.430 ;
        RECT 20.800 39.110 21.060 39.430 ;
        RECT 23.100 39.110 23.360 39.430 ;
        RECT 20.340 38.770 20.600 39.090 ;
        RECT 20.400 37.390 20.540 38.770 ;
        RECT 20.860 37.730 21.000 39.110 ;
        RECT 20.800 37.410 21.060 37.730 ;
        RECT 20.340 37.070 20.600 37.390 ;
        RECT 20.860 36.710 21.000 37.410 ;
        RECT 20.800 36.390 21.060 36.710 ;
        RECT 20.340 35.710 20.600 36.030 ;
        RECT 19.420 34.350 19.680 34.670 ;
        RECT 18.960 33.670 19.220 33.990 ;
        RECT 18.500 31.970 18.760 32.290 ;
        RECT 17.580 31.290 17.840 31.610 ;
        RECT 17.640 28.890 17.780 31.290 ;
        RECT 17.580 28.570 17.840 28.890 ;
        RECT 19.020 26.170 19.160 33.670 ;
        RECT 19.480 31.610 19.620 34.350 ;
        RECT 20.400 33.990 20.540 35.710 ;
        RECT 21.070 35.175 22.610 35.545 ;
        RECT 20.340 33.670 20.600 33.990 ;
        RECT 19.880 32.990 20.140 33.310 ;
        RECT 20.340 32.990 20.600 33.310 ;
        RECT 22.640 32.990 22.900 33.310 ;
        RECT 19.420 31.290 19.680 31.610 ;
        RECT 19.940 30.930 20.080 32.990 ;
        RECT 20.400 31.270 20.540 32.990 ;
        RECT 22.700 31.610 22.840 32.990 ;
        RECT 23.160 32.290 23.300 39.110 ;
        RECT 23.620 33.990 23.760 44.550 ;
        RECT 24.080 44.470 24.680 44.610 ;
        RECT 24.080 43.170 24.220 44.470 ;
        RECT 24.370 43.335 25.910 43.705 ;
        RECT 26.380 43.170 26.520 44.890 ;
        RECT 26.840 44.870 26.980 49.740 ;
        RECT 27.240 49.650 27.500 49.740 ;
        RECT 28.220 48.610 28.360 49.990 ;
        RECT 28.160 48.290 28.420 48.610 ;
        RECT 27.700 47.270 27.960 47.590 ;
        RECT 27.240 46.590 27.500 46.910 ;
        RECT 27.300 45.210 27.440 46.590 ;
        RECT 27.760 45.890 27.900 47.270 ;
        RECT 28.680 46.820 28.820 50.590 ;
        RECT 29.140 47.590 29.280 55.430 ;
        RECT 29.080 47.270 29.340 47.590 ;
        RECT 28.680 46.680 29.280 46.820 ;
        RECT 27.700 45.570 27.960 45.890 ;
        RECT 27.240 44.890 27.500 45.210 ;
        RECT 28.150 45.035 28.430 45.405 ;
        RECT 26.780 44.550 27.040 44.870 ;
        RECT 27.240 44.210 27.500 44.530 ;
        RECT 24.020 42.850 24.280 43.170 ;
        RECT 25.860 42.850 26.120 43.170 ;
        RECT 26.320 42.850 26.580 43.170 ;
        RECT 24.480 42.510 24.740 42.830 ;
        RECT 24.020 42.170 24.280 42.490 ;
        RECT 24.080 40.450 24.220 42.170 ;
        RECT 24.540 41.810 24.680 42.510 ;
        RECT 24.480 41.490 24.740 41.810 ;
        RECT 24.020 40.130 24.280 40.450 ;
        RECT 25.920 38.660 26.060 42.850 ;
        RECT 26.380 39.770 26.520 42.850 ;
        RECT 26.780 41.830 27.040 42.150 ;
        RECT 26.320 39.450 26.580 39.770 ;
        RECT 25.920 38.520 26.520 38.660 ;
        RECT 24.370 37.895 25.910 38.265 ;
        RECT 26.380 37.050 26.520 38.520 ;
        RECT 26.320 36.730 26.580 37.050 ;
        RECT 26.840 34.410 26.980 41.830 ;
        RECT 27.300 40.645 27.440 44.210 ;
        RECT 27.230 40.275 27.510 40.645 ;
        RECT 27.700 39.790 27.960 40.110 ;
        RECT 27.240 39.450 27.500 39.770 ;
        RECT 27.300 37.730 27.440 39.450 ;
        RECT 27.760 38.750 27.900 39.790 ;
        RECT 27.700 38.430 27.960 38.750 ;
        RECT 27.240 37.410 27.500 37.730 ;
        RECT 26.380 34.330 26.980 34.410 ;
        RECT 24.020 34.010 24.280 34.330 ;
        RECT 26.320 34.270 26.980 34.330 ;
        RECT 26.320 34.010 26.580 34.270 ;
        RECT 23.560 33.670 23.820 33.990 ;
        RECT 23.100 31.970 23.360 32.290 ;
        RECT 23.620 31.690 23.760 33.670 ;
        RECT 24.080 32.290 24.220 34.010 ;
        RECT 24.370 32.455 25.910 32.825 ;
        RECT 24.020 31.970 24.280 32.290 ;
        RECT 25.860 31.970 26.120 32.290 ;
        RECT 25.400 31.805 25.660 31.950 ;
        RECT 22.640 31.290 22.900 31.610 ;
        RECT 23.160 31.550 23.760 31.690 ;
        RECT 20.340 30.950 20.600 31.270 ;
        RECT 19.880 30.610 20.140 30.930 ;
        RECT 19.940 28.550 20.080 30.610 ;
        RECT 21.070 29.735 22.610 30.105 ;
        RECT 21.260 28.570 21.520 28.890 ;
        RECT 19.880 28.230 20.140 28.550 ;
        RECT 21.320 26.510 21.460 28.570 ;
        RECT 22.180 27.550 22.440 27.870 ;
        RECT 21.260 26.190 21.520 26.510 ;
        RECT 18.960 25.850 19.220 26.170 ;
        RECT 19.420 25.850 19.680 26.170 ;
        RECT 16.660 25.510 16.920 25.830 ;
        RECT 15.740 23.810 16.000 24.130 ;
        RECT 14.820 23.130 15.080 23.450 ;
        RECT 8.380 22.790 8.640 23.110 ;
        RECT 7.920 22.450 8.180 22.770 ;
        RECT 1.940 22.110 2.200 22.430 ;
        RECT 2.000 20.925 2.140 22.110 ;
        RECT 1.930 20.555 2.210 20.925 ;
        RECT 7.980 20.730 8.120 22.450 ;
        RECT 8.440 21.410 8.580 22.790 ;
        RECT 14.880 22.430 15.020 23.130 ;
        RECT 14.820 22.110 15.080 22.430 ;
        RECT 8.380 21.090 8.640 21.410 ;
        RECT 7.920 20.410 8.180 20.730 ;
        RECT 14.880 19.710 15.020 22.110 ;
        RECT 15.800 20.730 15.940 23.810 ;
        RECT 16.720 23.790 16.860 25.510 ;
        RECT 19.480 25.490 19.620 25.850 ;
        RECT 21.320 25.490 21.460 26.190 ;
        RECT 22.240 26.170 22.380 27.550 ;
        RECT 22.180 25.850 22.440 26.170 ;
        RECT 19.420 25.170 19.680 25.490 ;
        RECT 21.260 25.170 21.520 25.490 ;
        RECT 16.660 23.470 16.920 23.790 ;
        RECT 16.720 23.110 16.860 23.470 ;
        RECT 16.660 22.790 16.920 23.110 ;
        RECT 16.720 21.410 16.860 22.790 ;
        RECT 19.480 22.770 19.620 25.170 ;
        RECT 20.340 24.830 20.600 25.150 ;
        RECT 20.400 23.450 20.540 24.830 ;
        RECT 21.070 24.295 22.610 24.665 ;
        RECT 20.800 23.810 21.060 24.130 ;
        RECT 23.160 24.040 23.300 31.550 ;
        RECT 24.940 31.290 25.200 31.610 ;
        RECT 25.390 31.435 25.670 31.805 ;
        RECT 24.480 31.180 24.740 31.270 ;
        RECT 24.080 31.040 24.740 31.180 ;
        RECT 23.560 28.230 23.820 28.550 ;
        RECT 22.240 23.900 23.300 24.040 ;
        RECT 20.340 23.130 20.600 23.450 ;
        RECT 19.880 22.790 20.140 23.110 ;
        RECT 19.420 22.450 19.680 22.770 ;
        RECT 19.940 22.430 20.080 22.790 ;
        RECT 20.860 22.430 21.000 23.810 ;
        RECT 19.880 22.110 20.140 22.430 ;
        RECT 20.800 22.110 21.060 22.430 ;
        RECT 16.660 21.090 16.920 21.410 ;
        RECT 15.740 20.410 16.000 20.730 ;
        RECT 22.240 20.050 22.380 23.900 ;
        RECT 22.640 22.790 22.900 23.110 ;
        RECT 22.700 20.730 22.840 22.790 ;
        RECT 23.100 22.110 23.360 22.430 ;
        RECT 22.640 20.410 22.900 20.730 ;
        RECT 22.180 19.730 22.440 20.050 ;
        RECT 14.820 19.390 15.080 19.710 ;
        RECT 21.070 18.855 22.610 19.225 ;
        RECT 23.160 17.670 23.300 22.110 ;
        RECT 23.100 17.350 23.360 17.670 ;
        RECT 23.160 15.290 23.300 17.350 ;
        RECT 23.100 14.970 23.360 15.290 ;
        RECT 21.070 13.415 22.610 13.785 ;
        RECT 23.620 13.250 23.760 28.230 ;
        RECT 24.080 26.850 24.220 31.040 ;
        RECT 24.480 30.950 24.740 31.040 ;
        RECT 25.000 29.230 25.140 31.290 ;
        RECT 24.940 28.910 25.200 29.230 ;
        RECT 25.920 27.870 26.060 31.970 ;
        RECT 25.860 27.550 26.120 27.870 ;
        RECT 24.370 27.015 25.910 27.385 ;
        RECT 24.020 26.530 24.280 26.850 ;
        RECT 24.020 25.850 24.280 26.170 ;
        RECT 24.480 25.850 24.740 26.170 ;
        RECT 24.080 23.790 24.220 25.850 ;
        RECT 24.020 23.470 24.280 23.790 ;
        RECT 24.080 21.410 24.220 23.470 ;
        RECT 24.540 23.110 24.680 25.850 ;
        RECT 24.480 22.790 24.740 23.110 ;
        RECT 24.370 21.575 25.910 21.945 ;
        RECT 24.020 21.090 24.280 21.410 ;
        RECT 24.480 19.730 24.740 20.050 ;
        RECT 24.020 19.390 24.280 19.710 ;
        RECT 24.080 14.610 24.220 19.390 ;
        RECT 24.540 18.350 24.680 19.730 ;
        RECT 26.380 18.690 26.520 34.010 ;
        RECT 26.780 31.290 27.040 31.610 ;
        RECT 26.840 24.130 26.980 31.290 ;
        RECT 27.300 30.930 27.440 37.410 ;
        RECT 28.220 33.990 28.360 45.035 ;
        RECT 28.620 41.150 28.880 41.470 ;
        RECT 28.680 39.430 28.820 41.150 ;
        RECT 28.620 39.110 28.880 39.430 ;
        RECT 28.160 33.670 28.420 33.990 ;
        RECT 28.680 32.290 28.820 39.110 ;
        RECT 28.620 31.970 28.880 32.290 ;
        RECT 27.240 30.610 27.500 30.930 ;
        RECT 26.780 23.810 27.040 24.130 ;
        RECT 26.840 20.730 26.980 23.810 ;
        RECT 26.780 20.410 27.040 20.730 ;
        RECT 26.780 19.390 27.040 19.710 ;
        RECT 26.320 18.370 26.580 18.690 ;
        RECT 24.480 18.030 24.740 18.350 ;
        RECT 26.840 17.670 26.980 19.390 ;
        RECT 26.780 17.350 27.040 17.670 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 24.370 16.135 25.910 16.505 ;
        RECT 26.380 15.370 26.520 17.010 ;
        RECT 26.780 16.670 27.040 16.990 ;
        RECT 25.920 15.290 26.520 15.370 ;
        RECT 25.860 15.230 26.520 15.290 ;
        RECT 25.860 14.970 26.120 15.230 ;
        RECT 26.840 14.950 26.980 16.670 ;
        RECT 27.300 15.970 27.440 30.610 ;
        RECT 28.160 25.170 28.420 25.490 ;
        RECT 27.700 23.470 27.960 23.790 ;
        RECT 27.760 23.110 27.900 23.470 ;
        RECT 28.220 23.110 28.360 25.170 ;
        RECT 27.700 22.790 27.960 23.110 ;
        RECT 28.160 22.790 28.420 23.110 ;
        RECT 27.760 20.390 27.900 22.790 ;
        RECT 27.700 20.070 27.960 20.390 ;
        RECT 29.140 18.690 29.280 46.680 ;
        RECT 29.080 18.370 29.340 18.690 ;
        RECT 27.700 18.030 27.960 18.350 ;
        RECT 27.240 15.650 27.500 15.970 ;
        RECT 27.760 15.290 27.900 18.030 ;
        RECT 28.160 17.690 28.420 18.010 ;
        RECT 27.700 14.970 27.960 15.290 ;
        RECT 26.780 14.630 27.040 14.950 ;
        RECT 24.020 14.290 24.280 14.610 ;
        RECT 26.840 13.250 26.980 14.630 ;
        RECT 28.220 14.610 28.360 17.690 ;
        RECT 29.140 17.330 29.280 18.370 ;
        RECT 29.600 17.670 29.740 60.190 ;
        RECT 30.060 56.430 30.200 60.870 ;
        RECT 30.000 56.110 30.260 56.430 ;
        RECT 30.520 56.170 30.660 63.930 ;
        RECT 30.980 61.610 31.120 65.435 ;
        RECT 31.900 62.210 32.040 69.120 ;
        RECT 32.300 69.030 32.560 69.120 ;
        RECT 32.750 68.835 33.030 69.205 ;
        RECT 32.290 68.155 32.570 68.525 ;
        RECT 32.760 68.410 33.020 68.670 ;
        RECT 32.760 68.350 33.420 68.410 ;
        RECT 32.820 68.270 33.420 68.350 ;
        RECT 32.360 64.840 32.500 68.155 ;
        RECT 33.280 67.310 33.420 68.270 ;
        RECT 33.740 67.310 33.880 71.410 ;
        RECT 34.660 71.390 34.800 82.290 ;
        RECT 35.060 76.850 35.320 77.170 ;
        RECT 35.120 72.070 35.260 76.850 ;
        RECT 35.580 73.090 35.720 92.570 ;
        RECT 38.800 84.165 38.940 92.570 ;
        RECT 38.730 83.795 39.010 84.165 ;
        RECT 41.040 83.990 41.300 84.310 ;
        RECT 41.100 82.610 41.240 83.990 ;
        RECT 42.020 83.630 42.160 92.570 ;
        RECT 45.240 85.410 45.380 92.570 ;
        RECT 45.240 85.270 45.840 85.410 ;
        RECT 41.960 83.310 42.220 83.630 ;
        RECT 41.040 82.290 41.300 82.610 ;
        RECT 37.360 81.950 37.620 82.270 ;
        RECT 36.440 80.930 36.700 81.250 ;
        RECT 35.980 77.190 36.240 77.510 ;
        RECT 35.520 72.770 35.780 73.090 ;
        RECT 35.060 71.750 35.320 72.070 ;
        RECT 34.600 71.070 34.860 71.390 ;
        RECT 35.050 70.875 35.330 71.245 ;
        RECT 35.520 71.070 35.780 71.390 ;
        RECT 34.590 69.515 34.870 69.885 ;
        RECT 34.600 69.370 34.860 69.515 ;
        RECT 34.140 69.030 34.400 69.350 ;
        RECT 33.220 66.990 33.480 67.310 ;
        RECT 33.680 66.990 33.940 67.310 ;
        RECT 34.200 65.690 34.340 69.030 ;
        RECT 34.600 68.690 34.860 69.010 ;
        RECT 34.660 67.650 34.800 68.690 ;
        RECT 34.600 67.330 34.860 67.650 ;
        RECT 33.740 65.550 34.340 65.690 ;
        RECT 34.600 65.630 34.860 65.950 ;
        RECT 32.360 64.700 32.960 64.840 ;
        RECT 32.290 64.075 32.570 64.445 ;
        RECT 32.820 64.250 32.960 64.700 ;
        RECT 32.300 63.930 32.560 64.075 ;
        RECT 32.760 63.930 33.020 64.250 ;
        RECT 31.840 61.890 32.100 62.210 ;
        RECT 30.980 61.470 32.040 61.610 ;
        RECT 31.380 60.870 31.640 61.190 ;
        RECT 30.910 59.995 31.190 60.365 ;
        RECT 30.980 58.810 31.120 59.995 ;
        RECT 30.920 58.490 31.180 58.810 ;
        RECT 30.920 57.810 31.180 58.130 ;
        RECT 30.980 56.770 31.120 57.810 ;
        RECT 31.440 56.770 31.580 60.870 ;
        RECT 31.900 60.510 32.040 61.470 ;
        RECT 32.360 61.045 32.500 63.930 ;
        RECT 32.750 63.395 33.030 63.765 ;
        RECT 33.220 63.590 33.480 63.910 ;
        RECT 32.820 63.230 32.960 63.395 ;
        RECT 32.760 62.910 33.020 63.230 ;
        RECT 32.820 61.190 32.960 62.910 ;
        RECT 32.290 60.675 32.570 61.045 ;
        RECT 32.760 60.870 33.020 61.190 ;
        RECT 31.840 60.190 32.100 60.510 ;
        RECT 32.290 59.315 32.570 59.685 ;
        RECT 32.300 59.170 32.560 59.315 ;
        RECT 32.300 58.150 32.560 58.470 ;
        RECT 31.840 57.645 32.100 57.790 ;
        RECT 31.830 57.275 32.110 57.645 ;
        RECT 30.920 56.450 31.180 56.770 ;
        RECT 31.380 56.450 31.640 56.770 ;
        RECT 30.060 55.750 30.200 56.110 ;
        RECT 30.520 56.030 31.120 56.170 ;
        RECT 30.000 55.430 30.260 55.750 ;
        RECT 30.000 49.650 30.260 49.970 ;
        RECT 30.460 49.650 30.720 49.970 ;
        RECT 30.060 47.590 30.200 49.650 ;
        RECT 30.000 47.270 30.260 47.590 ;
        RECT 30.520 40.110 30.660 49.650 ;
        RECT 30.980 45.890 31.120 56.030 ;
        RECT 31.380 53.390 31.640 53.710 ;
        RECT 30.920 45.570 31.180 45.890 ;
        RECT 31.440 44.190 31.580 53.390 ;
        RECT 31.840 51.010 32.100 51.330 ;
        RECT 31.900 50.650 32.040 51.010 ;
        RECT 31.840 50.330 32.100 50.650 ;
        RECT 32.360 49.630 32.500 58.150 ;
        RECT 32.760 57.470 33.020 57.790 ;
        RECT 32.820 55.750 32.960 57.470 ;
        RECT 32.760 55.430 33.020 55.750 ;
        RECT 33.280 53.710 33.420 63.590 ;
        RECT 33.740 63.230 33.880 65.550 ;
        RECT 34.140 64.610 34.400 64.930 ;
        RECT 33.680 62.910 33.940 63.230 ;
        RECT 33.680 61.550 33.940 61.870 ;
        RECT 33.740 59.490 33.880 61.550 ;
        RECT 34.200 61.190 34.340 64.610 ;
        RECT 34.660 64.590 34.800 65.630 ;
        RECT 34.600 64.270 34.860 64.590 ;
        RECT 34.140 60.870 34.400 61.190 ;
        RECT 35.120 60.850 35.260 70.875 ;
        RECT 35.060 60.530 35.320 60.850 ;
        RECT 35.120 59.570 35.260 60.530 ;
        RECT 33.680 59.170 33.940 59.490 ;
        RECT 34.200 59.430 35.260 59.570 ;
        RECT 33.740 55.410 33.880 59.170 ;
        RECT 34.200 56.090 34.340 59.430 ;
        RECT 35.580 59.150 35.720 71.070 ;
        RECT 36.040 62.210 36.180 77.190 ;
        RECT 36.500 71.390 36.640 80.930 ;
        RECT 36.900 76.850 37.160 77.170 ;
        RECT 36.440 71.070 36.700 71.390 ;
        RECT 36.960 69.770 37.100 76.850 ;
        RECT 37.420 72.070 37.560 81.950 ;
        RECT 38.730 81.755 39.010 82.125 ;
        RECT 43.340 81.950 43.600 82.270 ;
        RECT 38.800 80.765 38.940 81.755 ;
        RECT 38.730 80.395 39.010 80.765 ;
        RECT 41.500 80.250 41.760 80.570 ;
        RECT 38.740 79.570 39.000 79.890 ;
        RECT 37.820 76.850 38.080 77.170 ;
        RECT 37.880 76.685 38.020 76.850 ;
        RECT 37.810 76.315 38.090 76.685 ;
        RECT 37.820 75.490 38.080 75.810 ;
        RECT 38.270 75.635 38.550 76.005 ;
        RECT 37.360 71.750 37.620 72.070 ;
        RECT 36.500 69.630 37.100 69.770 ;
        RECT 36.500 69.350 36.640 69.630 ;
        RECT 36.440 69.030 36.700 69.350 ;
        RECT 37.420 68.525 37.560 71.750 ;
        RECT 37.350 68.155 37.630 68.525 ;
        RECT 37.420 67.560 37.560 68.155 ;
        RECT 36.960 67.420 37.560 67.560 ;
        RECT 36.430 66.795 36.710 67.165 ;
        RECT 36.500 66.290 36.640 66.795 ;
        RECT 36.440 65.970 36.700 66.290 ;
        RECT 36.440 64.610 36.700 64.930 ;
        RECT 36.500 63.230 36.640 64.610 ;
        RECT 36.960 64.590 37.100 67.420 ;
        RECT 37.880 67.220 38.020 75.490 ;
        RECT 38.340 71.390 38.480 75.635 ;
        RECT 38.800 72.070 38.940 79.570 ;
        RECT 41.040 77.530 41.300 77.850 ;
        RECT 39.190 76.995 39.470 77.365 ;
        RECT 40.120 77.190 40.380 77.510 ;
        RECT 40.580 77.190 40.840 77.510 ;
        RECT 39.260 76.830 39.400 76.995 ;
        RECT 39.200 76.510 39.460 76.830 ;
        RECT 39.650 75.635 39.930 76.005 ;
        RECT 39.190 74.275 39.470 74.645 ;
        RECT 38.740 71.750 39.000 72.070 ;
        RECT 38.280 71.245 38.540 71.390 ;
        RECT 39.260 71.245 39.400 74.275 ;
        RECT 39.720 72.070 39.860 75.635 ;
        RECT 39.660 71.750 39.920 72.070 ;
        RECT 38.270 70.875 38.550 71.245 ;
        RECT 39.190 71.130 39.470 71.245 ;
        RECT 39.190 70.990 39.860 71.130 ;
        RECT 39.190 70.875 39.470 70.990 ;
        RECT 38.280 69.370 38.540 69.690 ;
        RECT 38.740 69.370 39.000 69.690 ;
        RECT 39.200 69.370 39.460 69.690 ;
        RECT 38.340 67.650 38.480 69.370 ;
        RECT 38.800 69.010 38.940 69.370 ;
        RECT 38.740 68.690 39.000 69.010 ;
        RECT 38.280 67.330 38.540 67.650 ;
        RECT 37.420 67.080 38.020 67.220 ;
        RECT 37.420 64.590 37.560 67.080 ;
        RECT 38.280 66.310 38.540 66.630 ;
        RECT 38.340 65.950 38.480 66.310 ;
        RECT 38.280 65.860 38.540 65.950 ;
        RECT 37.880 65.720 38.540 65.860 ;
        RECT 36.900 64.270 37.160 64.590 ;
        RECT 37.360 64.270 37.620 64.590 ;
        RECT 36.440 62.910 36.700 63.230 ;
        RECT 35.980 61.890 36.240 62.210 ;
        RECT 35.980 60.190 36.240 60.510 ;
        RECT 35.520 58.830 35.780 59.150 ;
        RECT 34.600 58.150 34.860 58.470 ;
        RECT 34.140 55.770 34.400 56.090 ;
        RECT 33.680 55.090 33.940 55.410 ;
        RECT 33.220 53.390 33.480 53.710 ;
        RECT 34.140 53.050 34.400 53.370 ;
        RECT 33.680 52.030 33.940 52.350 ;
        RECT 33.740 51.330 33.880 52.030 ;
        RECT 33.680 51.010 33.940 51.330 ;
        RECT 32.760 49.990 33.020 50.310 ;
        RECT 33.680 49.990 33.940 50.310 ;
        RECT 31.840 49.310 32.100 49.630 ;
        RECT 32.300 49.310 32.560 49.630 ;
        RECT 31.900 48.270 32.040 49.310 ;
        RECT 31.840 47.950 32.100 48.270 ;
        RECT 31.900 45.405 32.040 47.950 ;
        RECT 32.820 47.930 32.960 49.990 ;
        RECT 32.760 47.610 33.020 47.930 ;
        RECT 33.220 47.610 33.480 47.930 ;
        RECT 31.830 45.035 32.110 45.405 ;
        RECT 32.300 45.230 32.560 45.550 ;
        RECT 31.380 43.870 31.640 44.190 ;
        RECT 31.440 43.170 31.580 43.870 ;
        RECT 31.380 42.850 31.640 43.170 ;
        RECT 30.920 42.170 31.180 42.490 ;
        RECT 30.980 42.005 31.120 42.170 ;
        RECT 30.910 41.635 31.190 42.005 ;
        RECT 30.460 39.790 30.720 40.110 ;
        RECT 30.520 23.450 30.660 39.790 ;
        RECT 31.440 39.430 31.580 42.850 ;
        RECT 31.840 42.170 32.100 42.490 ;
        RECT 30.920 39.110 31.180 39.430 ;
        RECT 31.380 39.110 31.640 39.430 ;
        RECT 30.980 36.030 31.120 39.110 ;
        RECT 30.920 35.710 31.180 36.030 ;
        RECT 31.900 35.010 32.040 42.170 ;
        RECT 32.360 37.730 32.500 45.230 ;
        RECT 32.300 37.410 32.560 37.730 ;
        RECT 31.840 34.690 32.100 35.010 ;
        RECT 31.840 33.670 32.100 33.990 ;
        RECT 32.300 33.670 32.560 33.990 ;
        RECT 30.920 32.990 31.180 33.310 ;
        RECT 30.980 27.045 31.120 32.990 ;
        RECT 31.380 30.270 31.640 30.590 ;
        RECT 31.440 29.570 31.580 30.270 ;
        RECT 31.900 29.570 32.040 33.670 ;
        RECT 32.360 31.805 32.500 33.670 ;
        RECT 32.290 31.435 32.570 31.805 ;
        RECT 32.300 31.290 32.560 31.435 ;
        RECT 31.380 29.250 31.640 29.570 ;
        RECT 31.840 29.250 32.100 29.570 ;
        RECT 32.300 27.550 32.560 27.870 ;
        RECT 30.910 26.675 31.190 27.045 ;
        RECT 31.380 26.365 31.640 26.510 ;
        RECT 30.920 25.850 31.180 26.170 ;
        RECT 31.370 25.995 31.650 26.365 ;
        RECT 32.360 26.170 32.500 27.550 ;
        RECT 32.300 25.850 32.560 26.170 ;
        RECT 30.980 24.130 31.120 25.850 ;
        RECT 30.920 23.810 31.180 24.130 ;
        RECT 30.460 23.130 30.720 23.450 ;
        RECT 30.460 18.030 30.720 18.350 ;
        RECT 29.540 17.410 29.800 17.670 ;
        RECT 30.520 17.410 30.660 18.030 ;
        RECT 29.540 17.350 30.660 17.410 ;
        RECT 29.080 17.010 29.340 17.330 ;
        RECT 29.600 17.270 30.660 17.350 ;
        RECT 29.140 16.730 29.280 17.010 ;
        RECT 29.140 16.590 30.200 16.730 ;
        RECT 29.540 15.650 29.800 15.970 ;
        RECT 29.600 15.290 29.740 15.650 ;
        RECT 30.060 15.290 30.200 16.590 ;
        RECT 29.540 14.970 29.800 15.290 ;
        RECT 30.000 14.970 30.260 15.290 ;
        RECT 28.160 14.290 28.420 14.610 ;
        RECT 29.600 13.250 29.740 14.970 ;
        RECT 23.560 12.930 23.820 13.250 ;
        RECT 26.780 12.930 27.040 13.250 ;
        RECT 29.540 12.930 29.800 13.250 ;
        RECT 30.520 12.570 30.660 17.270 ;
        RECT 32.820 15.290 32.960 47.610 ;
        RECT 33.280 38.750 33.420 47.610 ;
        RECT 33.740 47.250 33.880 49.990 ;
        RECT 34.200 48.270 34.340 53.050 ;
        RECT 34.140 47.950 34.400 48.270 ;
        RECT 33.680 46.930 33.940 47.250 ;
        RECT 34.140 46.590 34.400 46.910 ;
        RECT 34.200 41.470 34.340 46.590 ;
        RECT 34.660 43.170 34.800 58.150 ;
        RECT 35.520 57.810 35.780 58.130 ;
        RECT 35.060 55.770 35.320 56.090 ;
        RECT 34.600 42.850 34.860 43.170 ;
        RECT 33.740 41.330 34.340 41.470 ;
        RECT 33.220 38.430 33.480 38.750 ;
        RECT 33.280 34.670 33.420 38.430 ;
        RECT 33.220 34.350 33.480 34.670 ;
        RECT 33.220 33.670 33.480 33.990 ;
        RECT 33.280 32.290 33.420 33.670 ;
        RECT 33.220 31.970 33.480 32.290 ;
        RECT 33.220 31.125 33.480 31.270 ;
        RECT 33.210 30.755 33.490 31.125 ;
        RECT 33.280 29.230 33.420 30.755 ;
        RECT 33.220 28.910 33.480 29.230 ;
        RECT 33.220 23.020 33.480 23.110 ;
        RECT 33.740 23.020 33.880 41.330 ;
        RECT 34.140 39.450 34.400 39.770 ;
        RECT 34.200 37.730 34.340 39.450 ;
        RECT 34.600 39.110 34.860 39.430 ;
        RECT 34.140 37.410 34.400 37.730 ;
        RECT 34.140 31.970 34.400 32.290 ;
        RECT 34.200 31.270 34.340 31.970 ;
        RECT 34.140 30.950 34.400 31.270 ;
        RECT 34.660 25.150 34.800 39.110 ;
        RECT 35.120 37.730 35.260 55.770 ;
        RECT 35.580 55.070 35.720 57.810 ;
        RECT 35.520 54.750 35.780 55.070 ;
        RECT 36.040 53.565 36.180 60.190 ;
        RECT 37.880 59.400 38.020 65.720 ;
        RECT 38.280 65.630 38.540 65.720 ;
        RECT 39.260 64.445 39.400 69.370 ;
        RECT 39.190 64.075 39.470 64.445 ;
        RECT 38.280 63.250 38.540 63.570 ;
        RECT 36.960 59.260 38.020 59.400 ;
        RECT 36.430 57.955 36.710 58.325 ;
        RECT 36.440 57.810 36.700 57.955 ;
        RECT 36.430 55.915 36.710 56.285 ;
        RECT 36.500 55.410 36.640 55.915 ;
        RECT 36.440 55.090 36.700 55.410 ;
        RECT 36.430 54.555 36.710 54.925 ;
        RECT 35.970 53.195 36.250 53.565 ;
        RECT 36.500 53.370 36.640 54.555 ;
        RECT 36.440 53.050 36.700 53.370 ;
        RECT 35.980 52.370 36.240 52.690 ;
        RECT 36.040 52.090 36.180 52.370 ;
        RECT 36.960 52.090 37.100 59.260 ;
        RECT 38.340 58.890 38.480 63.250 ;
        RECT 39.720 58.890 39.860 70.990 ;
        RECT 40.180 67.650 40.320 77.190 ;
        RECT 40.640 70.030 40.780 77.190 ;
        RECT 41.100 74.790 41.240 77.530 ;
        RECT 41.560 75.810 41.700 80.250 ;
        RECT 41.950 79.715 42.230 80.085 ;
        RECT 42.020 79.550 42.160 79.715 ;
        RECT 41.960 79.230 42.220 79.550 ;
        RECT 42.020 78.530 42.160 79.230 ;
        RECT 41.960 78.210 42.220 78.530 ;
        RECT 41.960 76.510 42.220 76.830 ;
        RECT 42.880 76.510 43.140 76.830 ;
        RECT 41.500 75.490 41.760 75.810 ;
        RECT 41.040 74.470 41.300 74.790 ;
        RECT 41.100 71.730 41.240 74.470 ;
        RECT 41.040 71.410 41.300 71.730 ;
        RECT 40.580 69.710 40.840 70.030 ;
        RECT 41.030 68.155 41.310 68.525 ;
        RECT 41.500 68.350 41.760 68.670 ;
        RECT 40.120 67.330 40.380 67.650 ;
        RECT 41.100 66.630 41.240 68.155 ;
        RECT 41.560 67.650 41.700 68.350 ;
        RECT 41.500 67.330 41.760 67.650 ;
        RECT 40.120 66.310 40.380 66.630 ;
        RECT 40.580 66.310 40.840 66.630 ;
        RECT 41.040 66.310 41.300 66.630 ;
        RECT 41.500 66.310 41.760 66.630 ;
        RECT 37.880 58.750 38.480 58.890 ;
        RECT 39.260 58.750 39.860 58.890 ;
        RECT 37.360 55.430 37.620 55.750 ;
        RECT 37.880 55.605 38.020 58.750 ;
        RECT 38.280 58.150 38.540 58.470 ;
        RECT 38.340 57.790 38.480 58.150 ;
        RECT 38.280 57.470 38.540 57.790 ;
        RECT 38.740 57.470 39.000 57.790 ;
        RECT 38.340 56.770 38.480 57.470 ;
        RECT 38.280 56.450 38.540 56.770 ;
        RECT 36.040 51.950 37.100 52.090 ;
        RECT 35.510 50.475 35.790 50.845 ;
        RECT 36.040 50.650 36.180 51.950 ;
        RECT 36.440 51.010 36.700 51.330 ;
        RECT 35.580 50.310 35.720 50.475 ;
        RECT 35.980 50.330 36.240 50.650 ;
        RECT 35.520 49.990 35.780 50.310 ;
        RECT 35.520 48.125 35.780 48.270 ;
        RECT 35.510 47.755 35.790 48.125 ;
        RECT 35.520 45.230 35.780 45.550 ;
        RECT 35.580 42.490 35.720 45.230 ;
        RECT 35.520 42.170 35.780 42.490 ;
        RECT 36.040 41.470 36.180 50.330 ;
        RECT 36.500 50.165 36.640 51.010 ;
        RECT 36.430 49.795 36.710 50.165 ;
        RECT 36.900 49.990 37.160 50.310 ;
        RECT 36.960 48.610 37.100 49.990 ;
        RECT 36.900 48.290 37.160 48.610 ;
        RECT 36.440 47.610 36.700 47.930 ;
        RECT 36.500 45.890 36.640 47.610 ;
        RECT 36.900 47.270 37.160 47.590 ;
        RECT 36.960 46.765 37.100 47.270 ;
        RECT 36.890 46.395 37.170 46.765 ;
        RECT 36.440 45.570 36.700 45.890 ;
        RECT 36.500 43.365 36.640 45.570 ;
        RECT 36.900 44.210 37.160 44.530 ;
        RECT 36.430 42.995 36.710 43.365 ;
        RECT 36.440 42.170 36.700 42.490 ;
        RECT 35.580 41.330 36.180 41.470 ;
        RECT 35.060 37.410 35.320 37.730 ;
        RECT 35.060 34.010 35.320 34.330 ;
        RECT 35.120 29.140 35.260 34.010 ;
        RECT 35.580 31.600 35.720 41.330 ;
        RECT 36.500 40.450 36.640 42.170 ;
        RECT 36.440 40.130 36.700 40.450 ;
        RECT 36.960 39.170 37.100 44.210 ;
        RECT 37.420 40.110 37.560 55.430 ;
        RECT 37.810 55.235 38.090 55.605 ;
        RECT 38.340 53.370 38.480 56.450 ;
        RECT 38.800 56.430 38.940 57.470 ;
        RECT 38.740 56.110 39.000 56.430 ;
        RECT 38.800 55.750 38.940 56.110 ;
        RECT 38.740 55.430 39.000 55.750 ;
        RECT 39.260 54.050 39.400 58.750 ;
        RECT 39.660 58.150 39.920 58.470 ;
        RECT 39.200 53.730 39.460 54.050 ;
        RECT 38.740 53.565 39.000 53.710 ;
        RECT 38.280 53.050 38.540 53.370 ;
        RECT 38.730 53.195 39.010 53.565 ;
        RECT 38.740 52.030 39.000 52.350 ;
        RECT 38.270 49.795 38.550 50.165 ;
        RECT 37.820 48.290 38.080 48.610 ;
        RECT 37.880 41.470 38.020 48.290 ;
        RECT 37.820 41.150 38.080 41.470 ;
        RECT 37.360 39.790 37.620 40.110 ;
        RECT 36.500 39.030 37.100 39.170 ;
        RECT 37.820 39.110 38.080 39.430 ;
        RECT 35.980 37.410 36.240 37.730 ;
        RECT 35.520 31.280 35.780 31.600 ;
        RECT 35.580 30.590 35.720 31.280 ;
        RECT 35.520 30.270 35.780 30.590 ;
        RECT 35.120 29.000 35.720 29.140 ;
        RECT 35.580 28.550 35.720 29.000 ;
        RECT 35.060 28.405 35.320 28.550 ;
        RECT 35.050 28.035 35.330 28.405 ;
        RECT 35.520 28.230 35.780 28.550 ;
        RECT 35.120 25.740 35.260 28.035 ;
        RECT 35.520 27.725 35.780 27.870 ;
        RECT 35.510 27.355 35.790 27.725 ;
        RECT 35.520 26.365 35.780 26.510 ;
        RECT 35.510 25.995 35.790 26.365 ;
        RECT 35.520 25.740 35.780 25.830 ;
        RECT 35.120 25.600 35.780 25.740 ;
        RECT 35.520 25.510 35.780 25.600 ;
        RECT 34.600 24.830 34.860 25.150 ;
        RECT 36.040 24.130 36.180 37.410 ;
        RECT 36.500 34.330 36.640 39.030 ;
        RECT 36.900 38.430 37.160 38.750 ;
        RECT 36.960 37.050 37.100 38.430 ;
        RECT 36.900 36.730 37.160 37.050 ;
        RECT 36.900 34.350 37.160 34.670 ;
        RECT 36.440 34.010 36.700 34.330 ;
        RECT 36.440 31.520 36.700 31.560 ;
        RECT 36.960 31.520 37.100 34.350 ;
        RECT 36.440 31.380 37.100 31.520 ;
        RECT 36.440 31.240 36.700 31.380 ;
        RECT 36.960 26.170 37.100 31.380 ;
        RECT 37.350 28.715 37.630 29.085 ;
        RECT 37.420 26.170 37.560 28.715 ;
        RECT 36.900 25.850 37.160 26.170 ;
        RECT 37.360 25.850 37.620 26.170 ;
        RECT 35.980 23.810 36.240 24.130 ;
        RECT 33.220 22.880 33.880 23.020 ;
        RECT 33.220 22.790 33.480 22.880 ;
        RECT 33.740 20.390 33.880 22.880 ;
        RECT 34.600 22.110 34.860 22.430 ;
        RECT 34.660 21.410 34.800 22.110 ;
        RECT 34.600 21.090 34.860 21.410 ;
        RECT 33.680 20.070 33.940 20.390 ;
        RECT 33.740 17.670 33.880 20.070 ;
        RECT 33.680 17.350 33.940 17.670 ;
        RECT 33.220 15.540 33.480 15.630 ;
        RECT 33.740 15.540 33.880 17.350 ;
        RECT 33.220 15.400 33.880 15.540 ;
        RECT 33.220 15.310 33.480 15.400 ;
        RECT 32.760 14.970 33.020 15.290 ;
        RECT 32.820 13.250 32.960 14.970 ;
        RECT 33.740 13.250 33.880 15.400 ;
        RECT 32.760 12.930 33.020 13.250 ;
        RECT 33.680 12.930 33.940 13.250 ;
        RECT 34.660 12.910 34.800 21.090 ;
        RECT 35.520 17.350 35.780 17.670 ;
        RECT 35.580 15.970 35.720 17.350 ;
        RECT 35.520 15.650 35.780 15.970 ;
        RECT 36.960 15.290 37.100 25.850 ;
        RECT 37.420 23.790 37.560 25.850 ;
        RECT 37.360 23.470 37.620 23.790 ;
        RECT 37.880 20.050 38.020 39.110 ;
        RECT 38.340 36.030 38.480 49.795 ;
        RECT 38.800 48.805 38.940 52.030 ;
        RECT 39.200 50.670 39.460 50.990 ;
        RECT 38.730 48.435 39.010 48.805 ;
        RECT 38.730 47.755 39.010 48.125 ;
        RECT 38.740 47.610 39.000 47.755 ;
        RECT 38.740 46.930 39.000 47.250 ;
        RECT 38.280 35.710 38.540 36.030 ;
        RECT 38.800 31.690 38.940 46.930 ;
        RECT 39.260 46.910 39.400 50.670 ;
        RECT 39.200 46.590 39.460 46.910 ;
        RECT 39.190 44.355 39.470 44.725 ;
        RECT 39.200 44.210 39.460 44.355 ;
        RECT 39.190 41.635 39.470 42.005 ;
        RECT 39.720 41.810 39.860 58.150 ;
        RECT 40.180 56.430 40.320 66.310 ;
        RECT 40.640 64.930 40.780 66.310 ;
        RECT 40.580 64.610 40.840 64.930 ;
        RECT 41.560 64.590 41.700 66.310 ;
        RECT 42.020 64.930 42.160 76.510 ;
        RECT 41.960 64.610 42.220 64.930 ;
        RECT 42.410 64.755 42.690 65.125 ;
        RECT 41.500 64.270 41.760 64.590 ;
        RECT 41.960 63.930 42.220 64.250 ;
        RECT 40.580 60.530 40.840 60.850 ;
        RECT 40.640 58.810 40.780 60.530 ;
        RECT 40.580 58.720 40.840 58.810 ;
        RECT 40.580 58.580 41.700 58.720 ;
        RECT 40.580 58.490 40.840 58.580 ;
        RECT 40.120 56.110 40.380 56.430 ;
        RECT 40.580 56.110 40.840 56.430 ;
        RECT 40.120 54.750 40.380 55.070 ;
        RECT 40.180 45.550 40.320 54.750 ;
        RECT 40.640 45.890 40.780 56.110 ;
        RECT 41.560 55.750 41.700 58.580 ;
        RECT 41.500 55.430 41.760 55.750 ;
        RECT 41.500 54.750 41.760 55.070 ;
        RECT 41.560 54.050 41.700 54.750 ;
        RECT 41.500 53.730 41.760 54.050 ;
        RECT 41.500 53.280 41.760 53.370 ;
        RECT 41.100 53.140 41.760 53.280 ;
        RECT 41.100 49.630 41.240 53.140 ;
        RECT 41.500 53.050 41.760 53.140 ;
        RECT 41.490 52.515 41.770 52.885 ;
        RECT 41.500 52.370 41.760 52.515 ;
        RECT 41.500 50.670 41.760 50.990 ;
        RECT 41.560 49.970 41.700 50.670 ;
        RECT 41.500 49.650 41.760 49.970 ;
        RECT 41.040 49.310 41.300 49.630 ;
        RECT 41.030 47.755 41.310 48.125 ;
        RECT 41.040 47.610 41.300 47.755 ;
        RECT 41.500 47.610 41.760 47.930 ;
        RECT 41.030 47.075 41.310 47.445 ;
        RECT 41.040 46.930 41.300 47.075 ;
        RECT 40.580 45.570 40.840 45.890 ;
        RECT 40.120 45.230 40.380 45.550 ;
        RECT 41.030 45.035 41.310 45.405 ;
        RECT 41.560 45.210 41.700 47.610 ;
        RECT 42.020 47.250 42.160 63.930 ;
        RECT 42.480 51.410 42.620 64.755 ;
        RECT 42.940 60.510 43.080 76.510 ;
        RECT 43.400 66.630 43.540 81.950 ;
        RECT 44.720 80.250 44.980 80.570 ;
        RECT 43.800 75.150 44.060 75.470 ;
        RECT 43.860 69.885 44.000 75.150 ;
        RECT 44.780 73.090 44.920 80.250 ;
        RECT 45.180 79.910 45.440 80.230 ;
        RECT 45.240 79.405 45.380 79.910 ;
        RECT 45.170 79.035 45.450 79.405 ;
        RECT 45.700 78.190 45.840 85.270 ;
        RECT 48.460 83.370 48.600 92.570 ;
        RECT 48.000 83.230 48.600 83.370 ;
        RECT 46.100 79.910 46.360 80.230 ;
        RECT 45.640 77.870 45.900 78.190 ;
        RECT 45.180 75.490 45.440 75.810 ;
        RECT 44.720 72.770 44.980 73.090 ;
        RECT 44.260 71.750 44.520 72.070 ;
        RECT 43.790 69.515 44.070 69.885 ;
        RECT 43.340 66.310 43.600 66.630 ;
        RECT 43.400 62.170 43.540 66.310 ;
        RECT 43.860 64.250 44.000 69.515 ;
        RECT 44.320 69.350 44.460 71.750 ;
        RECT 44.780 70.565 44.920 72.770 ;
        RECT 45.240 72.070 45.380 75.490 ;
        RECT 46.160 74.645 46.300 79.910 ;
        RECT 48.000 77.850 48.140 83.230 ;
        RECT 48.860 82.630 49.120 82.950 ;
        RECT 47.940 77.530 48.200 77.850 ;
        RECT 48.920 77.510 49.060 82.630 ;
        RECT 51.680 80.910 51.820 92.570 ;
        RECT 54.900 86.770 55.040 92.570 ;
        RECT 54.440 86.630 55.040 86.770 ;
        RECT 54.440 81.250 54.580 86.630 ;
        RECT 56.680 83.650 56.940 83.970 ;
        RECT 54.380 80.930 54.640 81.250 ;
        RECT 54.840 80.930 55.100 81.250 ;
        RECT 51.620 80.590 51.880 80.910 ;
        RECT 53.450 80.395 53.730 80.765 ;
        RECT 53.520 79.890 53.660 80.395 ;
        RECT 53.460 79.570 53.720 79.890 ;
        RECT 53.920 79.570 54.180 79.890 ;
        RECT 48.860 77.190 49.120 77.510 ;
        RECT 51.620 77.190 51.880 77.510 ;
        RECT 51.160 76.850 51.420 77.170 ;
        RECT 48.860 74.810 49.120 75.130 ;
        RECT 49.380 75.070 50.440 75.210 ;
        RECT 46.090 74.275 46.370 74.645 ;
        RECT 47.020 74.130 47.280 74.450 ;
        RECT 45.180 71.750 45.440 72.070 ;
        RECT 45.640 71.750 45.900 72.070 ;
        RECT 46.560 71.750 46.820 72.070 ;
        RECT 44.710 70.195 44.990 70.565 ;
        RECT 44.260 69.030 44.520 69.350 ;
        RECT 44.250 66.795 44.530 67.165 ;
        RECT 44.320 66.290 44.460 66.795 ;
        RECT 44.260 65.970 44.520 66.290 ;
        RECT 44.260 64.270 44.520 64.590 ;
        RECT 43.800 63.930 44.060 64.250 ;
        RECT 43.400 62.030 44.000 62.170 ;
        RECT 43.340 60.530 43.600 60.850 ;
        RECT 42.880 60.190 43.140 60.510 ;
        RECT 43.400 59.570 43.540 60.530 ;
        RECT 42.940 59.430 43.540 59.570 ;
        RECT 42.940 58.470 43.080 59.430 ;
        RECT 43.340 58.490 43.600 58.810 ;
        RECT 42.880 58.150 43.140 58.470 ;
        RECT 42.940 57.790 43.080 58.150 ;
        RECT 42.880 57.470 43.140 57.790 ;
        RECT 42.940 56.090 43.080 57.470 ;
        RECT 42.880 55.770 43.140 56.090 ;
        RECT 43.400 55.410 43.540 58.490 ;
        RECT 43.340 55.090 43.600 55.410 ;
        RECT 42.880 54.750 43.140 55.070 ;
        RECT 42.940 52.350 43.080 54.750 ;
        RECT 43.340 53.050 43.600 53.370 ;
        RECT 42.880 52.030 43.140 52.350 ;
        RECT 42.480 51.270 43.080 51.410 ;
        RECT 42.410 49.795 42.690 50.165 ;
        RECT 42.480 47.930 42.620 49.795 ;
        RECT 42.420 47.610 42.680 47.930 ;
        RECT 42.940 47.330 43.080 51.270 ;
        RECT 43.400 49.970 43.540 53.050 ;
        RECT 43.860 52.205 44.000 62.030 ;
        RECT 44.320 61.190 44.460 64.270 ;
        RECT 44.260 60.870 44.520 61.190 ;
        RECT 44.260 55.090 44.520 55.410 ;
        RECT 43.790 51.835 44.070 52.205 ;
        RECT 43.340 49.650 43.600 49.970 ;
        RECT 43.400 49.485 43.540 49.650 ;
        RECT 43.330 49.115 43.610 49.485 ;
        RECT 43.400 47.930 43.540 49.115 ;
        RECT 43.340 47.610 43.600 47.930 ;
        RECT 43.790 47.755 44.070 48.125 ;
        RECT 43.800 47.610 44.060 47.755 ;
        RECT 41.960 46.930 42.220 47.250 ;
        RECT 42.940 47.190 44.000 47.330 ;
        RECT 43.340 46.590 43.600 46.910 ;
        RECT 41.100 44.190 41.240 45.035 ;
        RECT 41.500 44.890 41.760 45.210 ;
        RECT 43.400 44.870 43.540 46.590 ;
        RECT 43.340 44.550 43.600 44.870 ;
        RECT 41.500 44.210 41.760 44.530 ;
        RECT 41.960 44.210 42.220 44.530 ;
        RECT 40.580 43.870 40.840 44.190 ;
        RECT 41.040 43.870 41.300 44.190 ;
        RECT 40.640 42.830 40.780 43.870 ;
        RECT 41.560 42.830 41.700 44.210 ;
        RECT 40.120 42.510 40.380 42.830 ;
        RECT 40.580 42.510 40.840 42.830 ;
        RECT 41.500 42.510 41.760 42.830 ;
        RECT 39.200 41.490 39.460 41.635 ;
        RECT 39.660 41.490 39.920 41.810 ;
        RECT 40.180 37.730 40.320 42.510 ;
        RECT 42.020 42.490 42.160 44.210 ;
        RECT 42.880 43.870 43.140 44.190 ;
        RECT 41.040 42.170 41.300 42.490 ;
        RECT 41.960 42.170 42.220 42.490 ;
        RECT 41.100 40.110 41.240 42.170 ;
        RECT 41.040 39.790 41.300 40.110 ;
        RECT 40.120 37.410 40.380 37.730 ;
        RECT 41.500 37.410 41.760 37.730 ;
        RECT 41.560 37.050 41.700 37.410 ;
        RECT 42.020 37.390 42.160 42.170 ;
        RECT 42.420 38.430 42.680 38.750 ;
        RECT 41.960 37.070 42.220 37.390 ;
        RECT 42.480 37.050 42.620 38.430 ;
        RECT 42.940 37.730 43.080 43.870 ;
        RECT 43.860 42.570 44.000 47.190 ;
        RECT 44.320 43.170 44.460 55.090 ;
        RECT 44.780 47.250 44.920 70.195 ;
        RECT 45.700 69.770 45.840 71.750 ;
        RECT 46.620 70.370 46.760 71.750 ;
        RECT 46.560 70.050 46.820 70.370 ;
        RECT 45.700 69.690 46.760 69.770 ;
        RECT 45.700 69.630 46.820 69.690 ;
        RECT 46.560 69.370 46.820 69.630 ;
        RECT 45.640 69.030 45.900 69.350 ;
        RECT 45.180 67.330 45.440 67.650 ;
        RECT 45.240 61.870 45.380 67.330 ;
        RECT 45.180 61.550 45.440 61.870 ;
        RECT 45.700 54.810 45.840 69.030 ;
        RECT 46.090 68.835 46.370 69.205 ;
        RECT 45.240 54.670 45.840 54.810 ;
        RECT 45.240 53.710 45.380 54.670 ;
        RECT 45.640 53.730 45.900 54.050 ;
        RECT 45.180 53.390 45.440 53.710 ;
        RECT 45.180 52.710 45.440 53.030 ;
        RECT 45.240 50.310 45.380 52.710 ;
        RECT 45.700 51.330 45.840 53.730 ;
        RECT 45.640 51.010 45.900 51.330 ;
        RECT 45.180 49.990 45.440 50.310 ;
        RECT 45.640 48.290 45.900 48.610 ;
        RECT 45.170 47.755 45.450 48.125 ;
        RECT 44.720 46.930 44.980 47.250 ;
        RECT 45.240 44.870 45.380 47.755 ;
        RECT 45.180 44.550 45.440 44.870 ;
        RECT 45.700 43.170 45.840 48.290 ;
        RECT 46.160 45.550 46.300 68.835 ;
        RECT 46.550 62.715 46.830 63.085 ;
        RECT 46.620 61.870 46.760 62.715 ;
        RECT 46.560 61.550 46.820 61.870 ;
        RECT 46.560 53.050 46.820 53.370 ;
        RECT 46.620 52.205 46.760 53.050 ;
        RECT 46.550 51.835 46.830 52.205 ;
        RECT 46.560 51.010 46.820 51.330 ;
        RECT 46.100 45.230 46.360 45.550 ;
        RECT 46.100 44.045 46.360 44.190 ;
        RECT 46.090 43.675 46.370 44.045 ;
        RECT 44.260 42.850 44.520 43.170 ;
        RECT 45.640 42.850 45.900 43.170 ;
        RECT 43.340 42.170 43.600 42.490 ;
        RECT 43.860 42.430 44.460 42.570 ;
        RECT 42.880 37.410 43.140 37.730 ;
        RECT 43.400 37.050 43.540 42.170 ;
        RECT 43.790 41.635 44.070 42.005 ;
        RECT 41.500 36.730 41.760 37.050 ;
        RECT 42.420 36.730 42.680 37.050 ;
        RECT 43.340 36.730 43.600 37.050 ;
        RECT 40.120 36.390 40.380 36.710 ;
        RECT 41.960 36.390 42.220 36.710 ;
        RECT 40.180 33.990 40.320 36.390 ;
        RECT 40.580 35.710 40.840 36.030 ;
        RECT 39.200 33.670 39.460 33.990 ;
        RECT 40.120 33.670 40.380 33.990 ;
        RECT 39.260 32.290 39.400 33.670 ;
        RECT 40.180 32.290 40.320 33.670 ;
        RECT 39.200 31.970 39.460 32.290 ;
        RECT 40.120 31.970 40.380 32.290 ;
        RECT 39.660 31.805 39.920 31.950 ;
        RECT 38.280 31.290 38.540 31.610 ;
        RECT 38.800 31.550 39.400 31.690 ;
        RECT 38.340 29.085 38.480 31.290 ;
        RECT 38.740 30.950 39.000 31.270 ;
        RECT 38.270 28.715 38.550 29.085 ;
        RECT 38.340 28.550 38.480 28.715 ;
        RECT 38.280 28.230 38.540 28.550 ;
        RECT 38.280 26.760 38.540 26.850 ;
        RECT 38.800 26.760 38.940 30.950 ;
        RECT 38.280 26.620 38.940 26.760 ;
        RECT 38.280 26.530 38.540 26.620 ;
        RECT 38.340 25.830 38.480 26.530 ;
        RECT 38.280 25.510 38.540 25.830 ;
        RECT 39.260 23.790 39.400 31.550 ;
        RECT 39.650 31.435 39.930 31.805 ;
        RECT 39.660 30.950 39.920 31.270 ;
        RECT 39.720 28.405 39.860 30.950 ;
        RECT 40.180 29.230 40.320 31.970 ;
        RECT 40.640 29.230 40.780 35.710 ;
        RECT 41.040 33.330 41.300 33.650 ;
        RECT 41.100 31.610 41.240 33.330 ;
        RECT 41.040 31.290 41.300 31.610 ;
        RECT 41.030 30.755 41.310 31.125 ;
        RECT 41.040 30.610 41.300 30.755 ;
        RECT 40.120 28.910 40.380 29.230 ;
        RECT 40.580 28.910 40.840 29.230 ;
        RECT 39.650 28.035 39.930 28.405 ;
        RECT 40.640 28.290 40.780 28.910 ;
        RECT 40.180 28.150 40.780 28.290 ;
        RECT 39.650 26.675 39.930 27.045 ;
        RECT 39.660 26.530 39.920 26.675 ;
        RECT 39.720 26.170 39.860 26.530 ;
        RECT 39.660 25.850 39.920 26.170 ;
        RECT 39.200 23.470 39.460 23.790 ;
        RECT 39.200 22.450 39.460 22.770 ;
        RECT 39.660 22.450 39.920 22.770 ;
        RECT 39.260 20.730 39.400 22.450 ;
        RECT 39.720 20.730 39.860 22.450 ;
        RECT 40.180 21.410 40.320 28.150 ;
        RECT 41.040 27.890 41.300 28.210 ;
        RECT 41.100 27.725 41.240 27.890 ;
        RECT 41.030 27.355 41.310 27.725 ;
        RECT 42.020 26.850 42.160 36.390 ;
        RECT 43.400 35.010 43.540 36.730 ;
        RECT 43.340 34.690 43.600 35.010 ;
        RECT 41.500 26.530 41.760 26.850 ;
        RECT 41.960 26.530 42.220 26.850 ;
        RECT 41.040 25.850 41.300 26.170 ;
        RECT 40.580 24.830 40.840 25.150 ;
        RECT 40.640 23.110 40.780 24.830 ;
        RECT 40.580 22.790 40.840 23.110 ;
        RECT 40.120 21.090 40.380 21.410 ;
        RECT 39.200 20.410 39.460 20.730 ;
        RECT 39.660 20.410 39.920 20.730 ;
        RECT 37.820 19.730 38.080 20.050 ;
        RECT 39.260 17.670 39.400 20.410 ;
        RECT 40.180 18.010 40.320 21.090 ;
        RECT 41.100 20.050 41.240 25.850 ;
        RECT 41.560 22.430 41.700 26.530 ;
        RECT 43.860 24.130 44.000 41.635 ;
        RECT 44.320 33.845 44.460 42.430 ;
        RECT 46.620 42.400 46.760 51.010 ;
        RECT 47.080 44.870 47.220 74.130 ;
        RECT 48.920 73.285 49.060 74.810 ;
        RECT 49.380 74.790 49.520 75.070 ;
        RECT 49.320 74.470 49.580 74.790 ;
        RECT 49.780 74.470 50.040 74.790 ;
        RECT 48.850 72.915 49.130 73.285 ;
        RECT 48.400 72.090 48.660 72.410 ;
        RECT 47.480 71.750 47.740 72.070 ;
        RECT 47.540 69.010 47.680 71.750 ;
        RECT 47.940 71.070 48.200 71.390 ;
        RECT 47.480 68.690 47.740 69.010 ;
        RECT 47.480 63.930 47.740 64.250 ;
        RECT 47.540 56.430 47.680 63.930 ;
        RECT 48.000 63.910 48.140 71.070 ;
        RECT 48.460 69.690 48.600 72.090 ;
        RECT 48.860 71.750 49.120 72.070 ;
        RECT 48.400 69.370 48.660 69.690 ;
        RECT 48.400 68.690 48.660 69.010 ;
        RECT 48.460 65.950 48.600 68.690 ;
        RECT 48.400 65.630 48.660 65.950 ;
        RECT 48.400 63.930 48.660 64.250 ;
        RECT 47.940 63.590 48.200 63.910 ;
        RECT 47.940 61.890 48.200 62.210 ;
        RECT 48.000 59.490 48.140 61.890 ;
        RECT 48.460 61.530 48.600 63.930 ;
        RECT 48.400 61.210 48.660 61.530 ;
        RECT 48.920 60.510 49.060 71.750 ;
        RECT 49.320 71.070 49.580 71.390 ;
        RECT 48.400 60.190 48.660 60.510 ;
        RECT 48.860 60.190 49.120 60.510 ;
        RECT 47.940 59.170 48.200 59.490 ;
        RECT 47.480 56.110 47.740 56.430 ;
        RECT 48.460 54.050 48.600 60.190 ;
        RECT 48.920 55.750 49.060 60.190 ;
        RECT 49.380 58.470 49.520 71.070 ;
        RECT 49.840 63.230 49.980 74.470 ;
        RECT 50.300 69.350 50.440 75.070 ;
        RECT 50.700 74.810 50.960 75.130 ;
        RECT 50.240 69.030 50.500 69.350 ;
        RECT 49.780 62.910 50.040 63.230 ;
        RECT 50.300 59.490 50.440 69.030 ;
        RECT 49.780 59.170 50.040 59.490 ;
        RECT 50.240 59.170 50.500 59.490 ;
        RECT 49.840 58.890 49.980 59.170 ;
        RECT 50.760 58.890 50.900 74.810 ;
        RECT 51.220 71.390 51.360 76.850 ;
        RECT 51.160 71.070 51.420 71.390 ;
        RECT 51.220 69.350 51.360 71.070 ;
        RECT 51.160 69.030 51.420 69.350 ;
        RECT 51.160 66.990 51.420 67.310 ;
        RECT 49.840 58.750 50.900 58.890 ;
        RECT 49.320 58.150 49.580 58.470 ;
        RECT 48.860 55.430 49.120 55.750 ;
        RECT 48.400 53.730 48.660 54.050 ;
        RECT 50.230 53.875 50.510 54.245 ;
        RECT 50.300 53.710 50.440 53.875 ;
        RECT 47.940 53.565 48.200 53.710 ;
        RECT 48.860 53.565 49.120 53.710 ;
        RECT 47.930 53.195 48.210 53.565 ;
        RECT 48.400 53.050 48.660 53.370 ;
        RECT 48.850 53.195 49.130 53.565 ;
        RECT 50.240 53.390 50.500 53.710 ;
        RECT 50.700 53.620 50.960 53.710 ;
        RECT 51.220 53.620 51.360 66.990 ;
        RECT 51.680 65.950 51.820 77.190 ;
        RECT 52.540 76.510 52.800 76.830 ;
        RECT 52.080 71.750 52.340 72.070 ;
        RECT 51.620 65.630 51.880 65.950 ;
        RECT 51.680 64.590 51.820 65.630 ;
        RECT 51.620 64.270 51.880 64.590 ;
        RECT 51.620 61.780 51.880 61.870 ;
        RECT 52.140 61.780 52.280 71.750 ;
        RECT 52.600 71.730 52.740 76.510 ;
        RECT 53.000 74.810 53.260 75.130 ;
        RECT 52.540 71.410 52.800 71.730 ;
        RECT 52.600 66.290 52.740 71.410 ;
        RECT 52.540 65.970 52.800 66.290 ;
        RECT 52.540 63.930 52.800 64.250 ;
        RECT 51.620 61.640 52.280 61.780 ;
        RECT 51.620 61.550 51.880 61.640 ;
        RECT 50.700 53.480 51.360 53.620 ;
        RECT 50.700 53.390 50.960 53.480 ;
        RECT 49.780 53.280 50.040 53.370 ;
        RECT 49.380 53.140 50.040 53.280 ;
        RECT 47.940 52.030 48.200 52.350 ;
        RECT 48.000 50.310 48.140 52.030 ;
        RECT 48.460 51.330 48.600 53.050 ;
        RECT 48.860 52.030 49.120 52.350 ;
        RECT 48.400 51.010 48.660 51.330 ;
        RECT 48.920 50.310 49.060 52.030 ;
        RECT 47.940 49.990 48.200 50.310 ;
        RECT 48.860 49.990 49.120 50.310 ;
        RECT 47.940 49.310 48.200 49.630 ;
        RECT 48.860 49.310 49.120 49.630 ;
        RECT 48.000 48.610 48.140 49.310 ;
        RECT 47.940 48.290 48.200 48.610 ;
        RECT 47.470 47.755 47.750 48.125 ;
        RECT 48.000 47.930 48.140 48.290 ;
        RECT 47.540 45.890 47.680 47.755 ;
        RECT 47.940 47.610 48.200 47.930 ;
        RECT 48.920 47.330 49.060 49.310 ;
        RECT 48.000 47.190 49.060 47.330 ;
        RECT 48.000 46.910 48.140 47.190 ;
        RECT 48.920 46.910 49.060 47.190 ;
        RECT 47.940 46.590 48.200 46.910 ;
        RECT 48.400 46.590 48.660 46.910 ;
        RECT 48.860 46.590 49.120 46.910 ;
        RECT 47.480 45.570 47.740 45.890 ;
        RECT 47.020 44.550 47.280 44.870 ;
        RECT 47.470 44.355 47.750 44.725 ;
        RECT 47.540 44.190 47.680 44.355 ;
        RECT 47.940 44.210 48.200 44.530 ;
        RECT 47.480 43.870 47.740 44.190 ;
        RECT 47.020 42.400 47.280 42.490 ;
        RECT 46.620 42.260 47.280 42.400 ;
        RECT 47.020 42.170 47.280 42.260 ;
        RECT 48.000 40.450 48.140 44.210 ;
        RECT 48.460 42.490 48.600 46.590 ;
        RECT 48.850 45.035 49.130 45.405 ;
        RECT 48.920 44.870 49.060 45.035 ;
        RECT 49.380 44.870 49.520 53.140 ;
        RECT 49.780 53.050 50.040 53.140 ;
        RECT 50.700 52.710 50.960 53.030 ;
        RECT 50.760 51.330 50.900 52.710 ;
        RECT 50.700 51.010 50.960 51.330 ;
        RECT 51.220 50.845 51.360 53.480 ;
        RECT 51.680 52.690 51.820 61.550 ;
        RECT 52.600 61.440 52.740 63.930 ;
        RECT 52.140 61.300 52.740 61.440 ;
        RECT 52.140 53.370 52.280 61.300 ;
        RECT 52.540 60.530 52.800 60.850 ;
        RECT 52.600 56.770 52.740 60.530 ;
        RECT 53.060 58.810 53.200 74.810 ;
        RECT 53.980 74.530 54.120 79.570 ;
        RECT 54.380 77.190 54.640 77.510 ;
        RECT 53.520 74.390 54.120 74.530 ;
        RECT 53.520 66.970 53.660 74.390 ;
        RECT 53.920 73.790 54.180 74.110 ;
        RECT 53.980 67.310 54.120 73.790 ;
        RECT 54.440 69.770 54.580 77.190 ;
        RECT 54.900 75.130 55.040 80.930 ;
        RECT 55.290 78.355 55.570 78.725 ;
        RECT 55.360 77.510 55.500 78.355 ;
        RECT 55.300 77.190 55.560 77.510 ;
        RECT 55.360 76.005 55.500 77.190 ;
        RECT 56.220 76.850 56.480 77.170 ;
        RECT 55.760 76.510 56.020 76.830 ;
        RECT 55.290 75.635 55.570 76.005 ;
        RECT 54.840 74.810 55.100 75.130 ;
        RECT 55.300 74.130 55.560 74.450 ;
        RECT 55.360 73.090 55.500 74.130 ;
        RECT 55.300 72.770 55.560 73.090 ;
        RECT 54.440 69.630 55.500 69.770 ;
        RECT 53.920 67.050 54.180 67.310 ;
        RECT 53.920 66.990 54.580 67.050 ;
        RECT 53.460 66.650 53.720 66.970 ;
        RECT 53.980 66.910 54.580 66.990 ;
        RECT 54.440 66.630 54.580 66.910 ;
        RECT 53.920 66.485 54.180 66.630 ;
        RECT 53.460 65.970 53.720 66.290 ;
        RECT 53.910 66.115 54.190 66.485 ;
        RECT 54.380 66.310 54.640 66.630 ;
        RECT 53.520 65.010 53.660 65.970 ;
        RECT 53.520 64.870 54.580 65.010 ;
        RECT 53.920 64.270 54.180 64.590 ;
        RECT 53.460 61.550 53.720 61.870 ;
        RECT 53.520 59.005 53.660 61.550 ;
        RECT 53.980 59.150 54.120 64.270 ;
        RECT 53.000 58.490 53.260 58.810 ;
        RECT 53.450 58.635 53.730 59.005 ;
        RECT 53.920 58.830 54.180 59.150 ;
        RECT 53.460 57.470 53.720 57.790 ;
        RECT 52.540 56.450 52.800 56.770 ;
        RECT 52.540 55.430 52.800 55.750 ;
        RECT 52.600 53.710 52.740 55.430 ;
        RECT 52.540 53.390 52.800 53.710 ;
        RECT 52.080 53.050 52.340 53.370 ;
        RECT 52.990 53.195 53.270 53.565 ;
        RECT 53.060 52.690 53.200 53.195 ;
        RECT 51.620 52.370 51.880 52.690 ;
        RECT 53.000 52.370 53.260 52.690 ;
        RECT 52.070 51.835 52.350 52.205 ;
        RECT 51.620 51.010 51.880 51.330 ;
        RECT 50.240 50.560 50.500 50.650 ;
        RECT 50.240 50.420 50.900 50.560 ;
        RECT 51.150 50.475 51.430 50.845 ;
        RECT 50.240 50.330 50.500 50.420 ;
        RECT 50.240 49.650 50.500 49.970 ;
        RECT 50.300 48.460 50.440 49.650 ;
        RECT 50.240 48.140 50.500 48.460 ;
        RECT 50.240 47.270 50.500 47.590 ;
        RECT 49.780 46.590 50.040 46.910 ;
        RECT 48.860 44.550 49.120 44.870 ;
        RECT 49.320 44.550 49.580 44.870 ;
        RECT 48.400 42.170 48.660 42.490 ;
        RECT 45.640 40.130 45.900 40.450 ;
        RECT 47.940 40.130 48.200 40.450 ;
        RECT 45.700 37.050 45.840 40.130 ;
        RECT 46.100 39.450 46.360 39.770 ;
        RECT 44.720 36.730 44.980 37.050 ;
        RECT 45.180 36.730 45.440 37.050 ;
        RECT 45.640 36.730 45.900 37.050 ;
        RECT 44.250 33.475 44.530 33.845 ;
        RECT 44.260 32.990 44.520 33.310 ;
        RECT 44.320 26.510 44.460 32.990 ;
        RECT 44.260 26.190 44.520 26.510 ;
        RECT 43.800 23.810 44.060 24.130 ;
        RECT 43.860 23.110 44.000 23.810 ;
        RECT 43.800 22.790 44.060 23.110 ;
        RECT 43.340 22.450 43.600 22.770 ;
        RECT 41.500 22.110 41.760 22.430 ;
        RECT 43.400 21.410 43.540 22.450 ;
        RECT 43.340 21.090 43.600 21.410 ;
        RECT 43.400 20.730 43.540 21.090 ;
        RECT 42.880 20.410 43.140 20.730 ;
        RECT 43.340 20.410 43.600 20.730 ;
        RECT 43.800 20.410 44.060 20.730 ;
        RECT 41.040 19.730 41.300 20.050 ;
        RECT 42.940 19.710 43.080 20.410 ;
        RECT 43.860 20.050 44.000 20.410 ;
        RECT 44.780 20.050 44.920 36.730 ;
        RECT 45.240 32.290 45.380 36.730 ;
        RECT 46.160 34.330 46.300 39.450 ;
        RECT 47.480 39.110 47.740 39.430 ;
        RECT 46.100 34.010 46.360 34.330 ;
        RECT 47.540 33.990 47.680 39.110 ;
        RECT 48.460 37.390 48.600 42.170 ;
        RECT 48.860 41.150 49.120 41.470 ;
        RECT 48.400 37.070 48.660 37.390 ;
        RECT 47.480 33.670 47.740 33.990 ;
        RECT 47.540 33.310 47.680 33.670 ;
        RECT 47.480 32.990 47.740 33.310 ;
        RECT 45.180 31.970 45.440 32.290 ;
        RECT 45.640 30.950 45.900 31.270 ;
        RECT 45.700 29.570 45.840 30.950 ;
        RECT 45.640 29.250 45.900 29.570 ;
        RECT 45.640 25.850 45.900 26.170 ;
        RECT 46.100 25.850 46.360 26.170 ;
        RECT 45.180 20.750 45.440 21.070 ;
        RECT 45.240 20.130 45.380 20.750 ;
        RECT 45.700 20.730 45.840 25.850 ;
        RECT 46.160 22.430 46.300 25.850 ;
        RECT 48.920 25.830 49.060 41.150 ;
        RECT 49.320 38.770 49.580 39.090 ;
        RECT 49.380 31.610 49.520 38.770 ;
        RECT 49.840 37.050 49.980 46.590 ;
        RECT 50.300 45.890 50.440 47.270 ;
        RECT 50.760 47.250 50.900 50.420 ;
        RECT 50.700 46.930 50.960 47.250 ;
        RECT 50.240 45.570 50.500 45.890 ;
        RECT 50.700 45.570 50.960 45.890 ;
        RECT 50.760 44.530 50.900 45.570 ;
        RECT 51.220 44.870 51.360 50.475 ;
        RECT 51.680 45.890 51.820 51.010 ;
        RECT 52.140 50.650 52.280 51.835 ;
        RECT 52.990 51.155 53.270 51.525 ;
        RECT 52.080 50.330 52.340 50.650 ;
        RECT 51.620 45.570 51.880 45.890 ;
        RECT 51.160 44.550 51.420 44.870 ;
        RECT 50.700 44.210 50.960 44.530 ;
        RECT 50.240 42.850 50.500 43.170 ;
        RECT 49.780 36.730 50.040 37.050 ;
        RECT 49.840 35.010 49.980 36.730 ;
        RECT 50.300 36.280 50.440 42.850 ;
        RECT 50.760 39.090 50.900 44.210 ;
        RECT 51.620 43.870 51.880 44.190 ;
        RECT 51.680 42.685 51.820 43.870 ;
        RECT 51.610 42.315 51.890 42.685 ;
        RECT 51.620 42.170 51.880 42.315 ;
        RECT 51.610 41.635 51.890 42.005 ;
        RECT 51.680 41.470 51.820 41.635 ;
        RECT 51.620 41.150 51.880 41.470 ;
        RECT 50.700 38.770 50.960 39.090 ;
        RECT 51.620 37.070 51.880 37.390 ;
        RECT 50.300 36.140 50.900 36.280 ;
        RECT 49.780 34.690 50.040 35.010 ;
        RECT 50.240 33.330 50.500 33.650 ;
        RECT 49.780 32.990 50.040 33.310 ;
        RECT 49.320 31.290 49.580 31.610 ;
        RECT 49.840 27.870 49.980 32.990 ;
        RECT 50.300 31.610 50.440 33.330 ;
        RECT 50.760 32.290 50.900 36.140 ;
        RECT 51.680 35.885 51.820 37.070 ;
        RECT 51.610 35.515 51.890 35.885 ;
        RECT 51.620 33.670 51.880 33.990 ;
        RECT 50.700 31.970 50.960 32.290 ;
        RECT 50.240 31.290 50.500 31.610 ;
        RECT 50.300 28.890 50.440 31.290 ;
        RECT 50.240 28.570 50.500 28.890 ;
        RECT 50.760 28.210 50.900 31.970 ;
        RECT 51.160 31.290 51.420 31.610 ;
        RECT 51.220 28.550 51.360 31.290 ;
        RECT 51.160 28.230 51.420 28.550 ;
        RECT 50.700 27.890 50.960 28.210 ;
        RECT 51.680 27.870 51.820 33.670 ;
        RECT 52.140 31.805 52.280 50.330 ;
        RECT 53.060 50.310 53.200 51.155 ;
        RECT 52.540 49.990 52.800 50.310 ;
        RECT 53.000 49.990 53.260 50.310 ;
        RECT 52.600 48.610 52.740 49.990 ;
        RECT 52.990 49.115 53.270 49.485 ;
        RECT 52.540 48.290 52.800 48.610 ;
        RECT 53.060 47.930 53.200 49.115 ;
        RECT 53.000 47.610 53.260 47.930 ;
        RECT 52.540 47.270 52.800 47.590 ;
        RECT 52.600 33.990 52.740 47.270 ;
        RECT 53.520 44.870 53.660 57.470 ;
        RECT 53.920 55.090 54.180 55.410 ;
        RECT 52.990 44.355 53.270 44.725 ;
        RECT 53.460 44.550 53.720 44.870 ;
        RECT 53.060 43.170 53.200 44.355 ;
        RECT 53.000 42.850 53.260 43.170 ;
        RECT 53.520 42.685 53.660 44.550 ;
        RECT 53.000 42.170 53.260 42.490 ;
        RECT 53.450 42.315 53.730 42.685 ;
        RECT 53.060 34.525 53.200 42.170 ;
        RECT 53.980 40.450 54.120 55.090 ;
        RECT 54.440 45.210 54.580 64.870 ;
        RECT 54.840 62.910 55.100 63.230 ;
        RECT 54.900 48.690 55.040 62.910 ;
        RECT 55.360 55.070 55.500 69.630 ;
        RECT 55.820 66.630 55.960 76.510 ;
        RECT 56.280 75.130 56.420 76.850 ;
        RECT 56.220 74.810 56.480 75.130 ;
        RECT 56.220 69.370 56.480 69.690 ;
        RECT 56.280 67.845 56.420 69.370 ;
        RECT 56.740 69.350 56.880 83.650 ;
        RECT 58.120 80.650 58.260 92.570 ;
        RECT 61.340 83.485 61.480 92.570 ;
        RECT 64.560 87.565 64.700 92.570 ;
        RECT 67.780 88.245 67.920 92.570 ;
        RECT 67.710 87.875 67.990 88.245 ;
        RECT 64.490 87.195 64.770 87.565 ;
        RECT 71.000 86.885 71.140 92.570 ;
        RECT 73.700 92.490 73.960 92.810 ;
        RECT 73.760 92.210 73.900 92.490 ;
        RECT 74.220 92.210 74.360 92.570 ;
        RECT 73.760 92.070 74.360 92.210 ;
        RECT 77.440 89.605 77.580 92.570 ;
        RECT 80.660 90.965 80.800 92.570 ;
        RECT 80.590 90.595 80.870 90.965 ;
        RECT 77.370 89.235 77.650 89.605 ;
        RECT 70.930 86.515 71.210 86.885 ;
        RECT 69.560 84.670 69.820 84.990 ;
        RECT 61.270 83.115 61.550 83.485 ;
        RECT 62.200 82.630 62.460 82.950 ;
        RECT 69.620 82.870 69.760 84.670 ;
        RECT 69.160 82.730 69.760 82.870 ;
        RECT 59.900 82.290 60.160 82.610 ;
        RECT 57.200 80.510 58.260 80.650 ;
        RECT 56.680 69.030 56.940 69.350 ;
        RECT 56.210 67.475 56.490 67.845 ;
        RECT 56.280 67.310 56.420 67.475 ;
        RECT 56.220 66.990 56.480 67.310 ;
        RECT 57.200 67.165 57.340 80.510 ;
        RECT 58.510 80.395 58.790 80.765 ;
        RECT 58.060 79.910 58.320 80.230 ;
        RECT 58.120 74.020 58.260 79.910 ;
        RECT 58.580 77.420 58.720 80.395 ;
        RECT 59.960 79.890 60.100 82.290 ;
        RECT 60.820 80.250 61.080 80.570 ;
        RECT 59.900 79.570 60.160 79.890 ;
        RECT 58.980 79.460 59.240 79.550 ;
        RECT 58.980 79.320 59.640 79.460 ;
        RECT 58.980 79.230 59.240 79.320 ;
        RECT 59.500 77.510 59.640 79.320 ;
        RECT 59.960 78.725 60.100 79.570 ;
        RECT 59.890 78.355 60.170 78.725 ;
        RECT 58.980 77.420 59.240 77.510 ;
        RECT 58.580 77.280 59.240 77.420 ;
        RECT 58.980 77.190 59.240 77.280 ;
        RECT 59.440 77.190 59.700 77.510 ;
        RECT 58.520 76.510 58.780 76.830 ;
        RECT 58.980 76.510 59.240 76.830 ;
        RECT 60.880 76.685 61.020 80.250 ;
        RECT 58.580 75.130 58.720 76.510 ;
        RECT 58.520 74.810 58.780 75.130 ;
        RECT 59.040 74.790 59.180 76.510 ;
        RECT 60.810 76.315 61.090 76.685 ;
        RECT 61.740 76.510 62.000 76.830 ;
        RECT 60.820 75.150 61.080 75.470 ;
        RECT 58.980 74.470 59.240 74.790 ;
        RECT 58.520 74.020 58.780 74.110 ;
        RECT 58.120 73.880 58.780 74.020 ;
        RECT 60.880 73.965 61.020 75.150 ;
        RECT 61.800 75.130 61.940 76.510 ;
        RECT 61.740 74.810 62.000 75.130 ;
        RECT 58.520 73.790 58.780 73.880 ;
        RECT 60.810 73.850 61.090 73.965 ;
        RECT 58.060 71.750 58.320 72.070 ;
        RECT 57.600 69.370 57.860 69.690 ;
        RECT 57.660 67.650 57.800 69.370 ;
        RECT 57.600 67.330 57.860 67.650 ;
        RECT 57.130 66.795 57.410 67.165 ;
        RECT 55.760 66.310 56.020 66.630 ;
        RECT 56.220 66.310 56.480 66.630 ;
        RECT 55.820 64.250 55.960 66.310 ;
        RECT 55.760 63.930 56.020 64.250 ;
        RECT 56.280 63.570 56.420 66.310 ;
        RECT 57.140 65.970 57.400 66.290 ;
        RECT 57.200 64.590 57.340 65.970 ;
        RECT 58.120 65.805 58.260 71.750 ;
        RECT 58.580 66.290 58.720 73.790 ;
        RECT 60.420 73.710 61.090 73.850 ;
        RECT 58.980 71.070 59.240 71.390 ;
        RECT 59.040 69.885 59.180 71.070 ;
        RECT 58.970 69.515 59.250 69.885 ;
        RECT 59.900 68.690 60.160 69.010 ;
        RECT 59.960 67.730 60.100 68.690 ;
        RECT 59.040 67.590 60.100 67.730 ;
        RECT 59.040 66.630 59.180 67.590 ;
        RECT 59.440 66.990 59.700 67.310 ;
        RECT 58.980 66.310 59.240 66.630 ;
        RECT 58.520 65.970 58.780 66.290 ;
        RECT 58.050 65.690 58.330 65.805 ;
        RECT 58.980 65.690 59.240 65.950 ;
        RECT 59.500 65.860 59.640 66.990 ;
        RECT 59.900 65.860 60.160 65.950 ;
        RECT 59.500 65.720 60.160 65.860 ;
        RECT 58.050 65.630 59.240 65.690 ;
        RECT 59.900 65.630 60.160 65.720 ;
        RECT 58.050 65.550 59.180 65.630 ;
        RECT 58.050 65.435 58.330 65.550 ;
        RECT 57.140 64.270 57.400 64.590 ;
        RECT 56.680 63.930 56.940 64.250 ;
        RECT 58.980 63.930 59.240 64.250 ;
        RECT 56.220 63.250 56.480 63.570 ;
        RECT 55.760 58.490 56.020 58.810 ;
        RECT 55.820 56.090 55.960 58.490 ;
        RECT 55.760 55.770 56.020 56.090 ;
        RECT 55.300 54.750 55.560 55.070 ;
        RECT 55.820 54.050 55.960 55.770 ;
        RECT 56.280 54.245 56.420 63.250 ;
        RECT 56.740 56.770 56.880 63.930 ;
        RECT 58.060 62.910 58.320 63.230 ;
        RECT 57.140 61.210 57.400 61.530 ;
        RECT 56.680 56.450 56.940 56.770 ;
        RECT 57.200 56.090 57.340 61.210 ;
        RECT 57.600 59.170 57.860 59.490 ;
        RECT 57.660 57.790 57.800 59.170 ;
        RECT 57.600 57.470 57.860 57.790 ;
        RECT 57.600 56.110 57.860 56.430 ;
        RECT 57.140 55.770 57.400 56.090 ;
        RECT 56.680 55.090 56.940 55.410 ;
        RECT 55.760 53.730 56.020 54.050 ;
        RECT 56.210 53.875 56.490 54.245 ;
        RECT 56.740 53.370 56.880 55.090 ;
        RECT 57.660 53.710 57.800 56.110 ;
        RECT 57.600 53.390 57.860 53.710 ;
        RECT 55.300 53.280 55.560 53.370 ;
        RECT 55.300 53.140 55.960 53.280 ;
        RECT 55.300 53.050 55.560 53.140 ;
        RECT 55.820 49.630 55.960 53.140 ;
        RECT 56.680 53.050 56.940 53.370 ;
        RECT 55.760 49.310 56.020 49.630 ;
        RECT 54.900 48.550 55.500 48.690 ;
        RECT 54.840 47.270 55.100 47.590 ;
        RECT 54.380 44.890 54.640 45.210 ;
        RECT 54.380 44.210 54.640 44.530 ;
        RECT 54.440 43.170 54.580 44.210 ;
        RECT 54.380 42.850 54.640 43.170 ;
        RECT 53.460 40.130 53.720 40.450 ;
        RECT 53.920 40.130 54.180 40.450 ;
        RECT 52.990 34.155 53.270 34.525 ;
        RECT 52.540 33.670 52.800 33.990 ;
        RECT 53.520 33.310 53.660 40.130 ;
        RECT 53.920 39.450 54.180 39.770 ;
        RECT 53.980 38.605 54.120 39.450 ;
        RECT 53.910 38.235 54.190 38.605 ;
        RECT 53.910 36.875 54.190 37.245 ;
        RECT 53.920 36.730 54.180 36.875 ;
        RECT 53.980 35.010 54.120 36.730 ;
        RECT 53.920 34.690 54.180 35.010 ;
        RECT 54.900 34.410 55.040 47.270 ;
        RECT 55.360 44.530 55.500 48.550 ;
        RECT 55.300 44.210 55.560 44.530 ;
        RECT 55.360 39.770 55.500 44.210 ;
        RECT 55.300 39.450 55.560 39.770 ;
        RECT 55.820 37.925 55.960 49.310 ;
        RECT 56.740 48.370 56.880 53.050 ;
        RECT 57.130 52.515 57.410 52.885 ;
        RECT 57.140 52.370 57.400 52.515 ;
        RECT 56.280 48.230 56.880 48.370 ;
        RECT 55.750 37.555 56.030 37.925 ;
        RECT 55.760 36.730 56.020 37.050 ;
        RECT 55.820 35.940 55.960 36.730 ;
        RECT 56.280 36.565 56.420 48.230 ;
        RECT 57.200 47.930 57.340 52.370 ;
        RECT 57.600 52.030 57.860 52.350 ;
        RECT 57.660 48.610 57.800 52.030 ;
        RECT 57.600 48.290 57.860 48.610 ;
        RECT 57.140 47.610 57.400 47.930 ;
        RECT 56.680 42.170 56.940 42.490 ;
        RECT 56.210 36.195 56.490 36.565 ;
        RECT 56.740 36.030 56.880 42.170 ;
        RECT 57.200 42.005 57.340 47.610 ;
        RECT 57.660 42.490 57.800 48.290 ;
        RECT 57.600 42.170 57.860 42.490 ;
        RECT 58.120 42.150 58.260 62.910 ;
        RECT 58.520 59.170 58.780 59.490 ;
        RECT 58.580 58.470 58.720 59.170 ;
        RECT 58.520 58.150 58.780 58.470 ;
        RECT 58.520 49.990 58.780 50.310 ;
        RECT 58.580 44.870 58.720 49.990 ;
        RECT 59.040 45.550 59.180 63.930 ;
        RECT 60.420 62.170 60.560 73.710 ;
        RECT 60.810 73.595 61.090 73.710 ;
        RECT 62.260 70.370 62.400 82.630 ;
        RECT 66.330 81.075 66.610 81.445 ;
        RECT 64.960 78.210 65.220 78.530 ;
        RECT 64.040 77.420 64.300 77.510 ;
        RECT 64.040 77.280 64.700 77.420 ;
        RECT 64.040 77.190 64.300 77.280 ;
        RECT 62.660 75.325 62.920 75.470 ;
        RECT 62.650 74.955 62.930 75.325 ;
        RECT 64.560 74.790 64.700 77.280 ;
        RECT 65.020 77.170 65.160 78.210 ;
        RECT 66.400 77.510 66.540 81.075 ;
        RECT 66.800 79.910 67.060 80.230 ;
        RECT 66.860 79.550 67.000 79.910 ;
        RECT 66.800 79.230 67.060 79.550 ;
        RECT 66.340 77.190 66.600 77.510 ;
        RECT 64.960 76.850 65.220 77.170 ;
        RECT 65.410 74.955 65.690 75.325 ;
        RECT 64.500 74.470 64.760 74.790 ;
        RECT 62.200 70.050 62.460 70.370 ;
        RECT 60.820 66.650 61.080 66.970 ;
        RECT 59.960 62.030 60.560 62.170 ;
        RECT 58.980 45.230 59.240 45.550 ;
        RECT 58.520 44.610 58.780 44.870 ;
        RECT 58.520 44.550 59.640 44.610 ;
        RECT 58.580 44.470 59.640 44.550 ;
        RECT 59.960 44.530 60.100 62.030 ;
        RECT 60.880 58.810 61.020 66.650 ;
        RECT 61.740 65.970 62.000 66.290 ;
        RECT 61.800 61.190 61.940 65.970 ;
        RECT 62.260 64.930 62.400 70.050 ;
        RECT 64.560 69.885 64.700 74.470 ;
        RECT 64.490 69.515 64.770 69.885 ;
        RECT 63.120 68.350 63.380 68.670 ;
        RECT 63.180 64.930 63.320 68.350 ;
        RECT 63.570 68.155 63.850 68.525 ;
        RECT 62.200 64.610 62.460 64.930 ;
        RECT 63.120 64.610 63.380 64.930 ;
        RECT 61.740 60.870 62.000 61.190 ;
        RECT 62.260 60.850 62.400 64.610 ;
        RECT 63.180 64.250 63.320 64.610 ;
        RECT 63.120 63.930 63.380 64.250 ;
        RECT 62.660 63.590 62.920 63.910 ;
        RECT 61.280 60.530 61.540 60.850 ;
        RECT 62.200 60.530 62.460 60.850 ;
        RECT 60.820 58.490 61.080 58.810 ;
        RECT 60.820 56.450 61.080 56.770 ;
        RECT 60.360 52.370 60.620 52.690 ;
        RECT 60.420 50.310 60.560 52.370 ;
        RECT 60.880 50.310 61.020 56.450 ;
        RECT 60.360 49.990 60.620 50.310 ;
        RECT 60.820 49.990 61.080 50.310 ;
        RECT 61.340 48.270 61.480 60.530 ;
        RECT 62.200 58.830 62.460 59.150 ;
        RECT 61.280 47.950 61.540 48.270 ;
        RECT 62.260 45.890 62.400 58.830 ;
        RECT 62.720 55.070 62.860 63.590 ;
        RECT 63.120 62.910 63.380 63.230 ;
        RECT 63.180 58.810 63.320 62.910 ;
        RECT 63.640 60.930 63.780 68.155 ;
        RECT 64.040 65.630 64.300 65.950 ;
        RECT 64.100 64.250 64.240 65.630 ;
        RECT 64.040 63.930 64.300 64.250 ;
        RECT 64.560 62.970 64.700 69.515 ;
        RECT 64.960 63.930 65.220 64.250 ;
        RECT 65.020 63.570 65.160 63.930 ;
        RECT 64.960 63.250 65.220 63.570 ;
        RECT 64.560 62.830 65.160 62.970 ;
        RECT 63.640 60.790 64.240 60.930 ;
        RECT 64.100 60.760 64.240 60.790 ;
        RECT 64.100 60.620 64.700 60.760 ;
        RECT 63.580 60.190 63.840 60.510 ;
        RECT 63.120 58.490 63.380 58.810 ;
        RECT 63.640 56.090 63.780 60.190 ;
        RECT 64.560 56.965 64.700 60.620 ;
        RECT 64.490 56.595 64.770 56.965 ;
        RECT 63.580 55.770 63.840 56.090 ;
        RECT 62.660 54.750 62.920 55.070 ;
        RECT 62.720 46.910 62.860 54.750 ;
        RECT 64.490 51.835 64.770 52.205 ;
        RECT 63.570 51.155 63.850 51.525 ;
        RECT 62.660 46.590 62.920 46.910 ;
        RECT 62.200 45.570 62.460 45.890 ;
        RECT 60.820 44.890 61.080 45.210 ;
        RECT 61.280 44.890 61.540 45.210 ;
        RECT 60.360 44.550 60.620 44.870 ;
        RECT 59.500 43.170 59.640 44.470 ;
        RECT 59.900 44.210 60.160 44.530 ;
        RECT 58.980 42.850 59.240 43.170 ;
        RECT 59.440 42.850 59.700 43.170 ;
        RECT 58.520 42.170 58.780 42.490 ;
        RECT 57.130 41.635 57.410 42.005 ;
        RECT 58.060 41.830 58.320 42.150 ;
        RECT 58.580 42.005 58.720 42.170 ;
        RECT 58.510 41.635 58.790 42.005 ;
        RECT 57.590 40.955 57.870 41.325 ;
        RECT 57.140 39.110 57.400 39.430 ;
        RECT 57.200 36.030 57.340 39.110 ;
        RECT 57.660 37.810 57.800 40.955 ;
        RECT 58.060 40.130 58.320 40.450 ;
        RECT 58.120 39.965 58.260 40.130 ;
        RECT 58.050 39.595 58.330 39.965 ;
        RECT 58.120 39.430 58.260 39.595 ;
        RECT 58.060 39.110 58.320 39.430 ;
        RECT 59.040 38.605 59.180 42.850 ;
        RECT 59.430 42.315 59.710 42.685 ;
        RECT 59.900 42.510 60.160 42.830 ;
        RECT 59.440 42.170 59.700 42.315 ;
        RECT 59.960 40.450 60.100 42.510 ;
        RECT 59.440 40.130 59.700 40.450 ;
        RECT 59.900 40.130 60.160 40.450 ;
        RECT 58.970 38.235 59.250 38.605 ;
        RECT 57.660 37.670 58.720 37.810 ;
        RECT 57.600 36.730 57.860 37.050 ;
        RECT 55.820 35.800 56.420 35.940 ;
        RECT 54.900 34.270 55.500 34.410 ;
        RECT 54.840 33.670 55.100 33.990 ;
        RECT 53.460 32.990 53.720 33.310 ;
        RECT 52.070 31.435 52.350 31.805 ;
        RECT 54.380 31.290 54.640 31.610 ;
        RECT 54.440 31.125 54.580 31.290 ;
        RECT 54.370 30.755 54.650 31.125 ;
        RECT 54.900 30.590 55.040 33.670 ;
        RECT 54.840 30.270 55.100 30.590 ;
        RECT 55.360 27.870 55.500 34.270 ;
        RECT 56.280 32.290 56.420 35.800 ;
        RECT 56.680 35.710 56.940 36.030 ;
        RECT 57.140 35.710 57.400 36.030 ;
        RECT 57.660 32.290 57.800 36.730 ;
        RECT 58.050 36.195 58.330 36.565 ;
        RECT 58.120 33.990 58.260 36.195 ;
        RECT 58.580 35.010 58.720 37.670 ;
        RECT 58.970 37.555 59.250 37.925 ;
        RECT 59.040 37.390 59.180 37.555 ;
        RECT 58.980 37.070 59.240 37.390 ;
        RECT 59.500 37.050 59.640 40.130 ;
        RECT 59.900 39.450 60.160 39.770 ;
        RECT 59.960 37.050 60.100 39.450 ;
        RECT 60.420 39.430 60.560 44.550 ;
        RECT 60.360 39.110 60.620 39.430 ;
        RECT 59.440 36.730 59.700 37.050 ;
        RECT 59.900 36.730 60.160 37.050 ;
        RECT 60.420 36.620 60.560 39.110 ;
        RECT 60.880 37.390 61.020 44.890 ;
        RECT 61.340 44.725 61.480 44.890 ;
        RECT 61.270 44.355 61.550 44.725 ;
        RECT 61.280 42.170 61.540 42.490 ;
        RECT 61.740 42.170 62.000 42.490 ;
        RECT 61.340 39.850 61.480 42.170 ;
        RECT 61.800 40.450 61.940 42.170 ;
        RECT 61.740 40.130 62.000 40.450 ;
        RECT 61.340 39.710 61.940 39.850 ;
        RECT 61.280 39.110 61.540 39.430 ;
        RECT 60.820 37.070 61.080 37.390 ;
        RECT 59.890 36.195 60.170 36.565 ;
        RECT 60.420 36.480 61.020 36.620 ;
        RECT 59.960 36.030 60.100 36.195 ;
        RECT 59.900 35.710 60.160 36.030 ;
        RECT 58.520 34.690 58.780 35.010 ;
        RECT 59.430 34.835 59.710 35.205 ;
        RECT 58.980 34.350 59.240 34.670 ;
        RECT 58.060 33.900 58.320 33.990 ;
        RECT 58.060 33.760 58.720 33.900 ;
        RECT 58.060 33.670 58.320 33.760 ;
        RECT 58.060 32.990 58.320 33.310 ;
        RECT 56.220 31.970 56.480 32.290 ;
        RECT 57.600 31.970 57.860 32.290 ;
        RECT 56.670 30.755 56.950 31.125 ;
        RECT 49.780 27.550 50.040 27.870 ;
        RECT 51.620 27.550 51.880 27.870 ;
        RECT 55.300 27.550 55.560 27.870 ;
        RECT 46.560 25.510 46.820 25.830 ;
        RECT 48.860 25.510 49.120 25.830 ;
        RECT 46.100 22.110 46.360 22.430 ;
        RECT 46.620 20.730 46.760 25.510 ;
        RECT 49.320 24.830 49.580 25.150 ;
        RECT 48.850 23.955 49.130 24.325 ;
        RECT 48.920 23.790 49.060 23.955 ;
        RECT 48.390 23.275 48.670 23.645 ;
        RECT 48.860 23.470 49.120 23.790 ;
        RECT 48.400 23.130 48.660 23.275 ;
        RECT 47.940 22.790 48.200 23.110 ;
        RECT 47.020 22.110 47.280 22.430 ;
        RECT 47.080 20.730 47.220 22.110 ;
        RECT 47.480 20.750 47.740 21.070 ;
        RECT 45.640 20.410 45.900 20.730 ;
        RECT 46.560 20.410 46.820 20.730 ;
        RECT 47.020 20.410 47.280 20.730 ;
        RECT 45.240 20.050 45.840 20.130 ;
        RECT 43.800 19.730 44.060 20.050 ;
        RECT 44.720 19.730 44.980 20.050 ;
        RECT 45.240 19.990 45.900 20.050 ;
        RECT 45.640 19.730 45.900 19.990 ;
        RECT 42.880 19.390 43.140 19.710 ;
        RECT 46.620 18.690 46.760 20.410 ;
        RECT 46.560 18.370 46.820 18.690 ;
        RECT 47.540 18.350 47.680 20.750 ;
        RECT 47.480 18.030 47.740 18.350 ;
        RECT 40.120 17.690 40.380 18.010 ;
        RECT 48.000 17.670 48.140 22.790 ;
        RECT 48.860 20.925 49.120 21.070 ;
        RECT 48.850 20.555 49.130 20.925 ;
        RECT 49.380 20.760 49.520 24.830 ;
        RECT 49.840 23.110 49.980 27.550 ;
        RECT 50.700 25.850 50.960 26.170 ;
        RECT 50.240 25.005 50.500 25.150 ;
        RECT 50.230 24.635 50.510 25.005 ;
        RECT 50.760 23.790 50.900 25.850 ;
        RECT 54.840 25.510 55.100 25.830 ;
        RECT 51.160 24.830 51.420 25.150 ;
        RECT 53.460 24.830 53.720 25.150 ;
        RECT 51.220 24.325 51.360 24.830 ;
        RECT 51.150 23.955 51.430 24.325 ;
        RECT 53.520 24.130 53.660 24.830 ;
        RECT 53.460 23.810 53.720 24.130 ;
        RECT 50.700 23.700 50.960 23.790 ;
        RECT 50.300 23.560 50.960 23.700 ;
        RECT 49.780 22.790 50.040 23.110 ;
        RECT 49.320 20.440 49.580 20.760 ;
        RECT 48.390 18.515 48.670 18.885 ;
        RECT 48.400 18.370 48.660 18.515 ;
        RECT 49.840 17.670 49.980 22.790 ;
        RECT 50.300 20.730 50.440 23.560 ;
        RECT 50.700 23.470 50.960 23.560 ;
        RECT 52.070 23.275 52.350 23.645 ;
        RECT 52.140 23.110 52.280 23.275 ;
        RECT 53.520 23.110 53.660 23.810 ;
        RECT 52.080 22.790 52.340 23.110 ;
        RECT 53.460 22.790 53.720 23.110 ;
        RECT 50.700 21.090 50.960 21.410 ;
        RECT 50.760 20.730 50.900 21.090 ;
        RECT 50.240 20.410 50.500 20.730 ;
        RECT 50.700 20.410 50.960 20.730 ;
        RECT 51.610 20.555 51.890 20.925 ;
        RECT 51.620 20.410 51.880 20.555 ;
        RECT 50.760 18.690 50.900 20.410 ;
        RECT 52.140 18.885 52.280 22.790 ;
        RECT 50.700 18.370 50.960 18.690 ;
        RECT 52.070 18.515 52.350 18.885 ;
        RECT 52.140 17.670 52.280 18.515 ;
        RECT 53.520 17.670 53.660 22.790 ;
        RECT 54.900 21.070 55.040 25.510 ;
        RECT 56.740 22.770 56.880 30.755 ;
        RECT 57.140 30.610 57.400 30.930 ;
        RECT 57.200 28.210 57.340 30.610 ;
        RECT 58.120 29.230 58.260 32.990 ;
        RECT 58.580 32.485 58.720 33.760 ;
        RECT 58.510 32.115 58.790 32.485 ;
        RECT 59.040 31.610 59.180 34.350 ;
        RECT 58.520 31.290 58.780 31.610 ;
        RECT 58.980 31.290 59.240 31.610 ;
        RECT 58.580 29.570 58.720 31.290 ;
        RECT 59.040 30.930 59.180 31.290 ;
        RECT 58.980 30.610 59.240 30.930 ;
        RECT 58.520 29.250 58.780 29.570 ;
        RECT 58.060 28.910 58.320 29.230 ;
        RECT 58.580 28.550 58.720 29.250 ;
        RECT 58.520 28.230 58.780 28.550 ;
        RECT 57.140 27.890 57.400 28.210 ;
        RECT 57.200 23.790 57.340 27.890 ;
        RECT 58.520 27.550 58.780 27.870 ;
        RECT 58.580 26.250 58.720 27.550 ;
        RECT 59.040 26.850 59.180 30.610 ;
        RECT 58.980 26.530 59.240 26.850 ;
        RECT 59.500 26.510 59.640 34.835 ;
        RECT 60.880 34.330 61.020 36.480 ;
        RECT 61.340 35.205 61.480 39.110 ;
        RECT 61.800 38.750 61.940 39.710 ;
        RECT 61.740 38.430 62.000 38.750 ;
        RECT 61.270 34.835 61.550 35.205 ;
        RECT 61.800 35.010 61.940 38.430 ;
        RECT 62.260 37.390 62.400 45.570 ;
        RECT 63.640 44.870 63.780 51.155 ;
        RECT 64.040 45.230 64.300 45.550 ;
        RECT 63.580 44.550 63.840 44.870 ;
        RECT 62.660 44.210 62.920 44.530 ;
        RECT 62.720 40.110 62.860 44.210 ;
        RECT 62.660 39.790 62.920 40.110 ;
        RECT 63.120 39.110 63.380 39.430 ;
        RECT 62.200 37.070 62.460 37.390 ;
        RECT 61.740 34.690 62.000 35.010 ;
        RECT 61.800 34.410 61.940 34.690 ;
        RECT 60.820 34.010 61.080 34.330 ;
        RECT 61.340 34.270 61.940 34.410 ;
        RECT 61.340 33.730 61.480 34.270 ;
        RECT 62.650 34.155 62.930 34.525 ;
        RECT 59.900 33.330 60.160 33.650 ;
        RECT 60.420 33.590 61.480 33.730 ;
        RECT 59.960 31.610 60.100 33.330 ;
        RECT 60.420 32.290 60.560 33.590 ;
        RECT 62.720 33.310 62.860 34.155 ;
        RECT 60.820 32.990 61.080 33.310 ;
        RECT 61.280 32.990 61.540 33.310 ;
        RECT 62.660 32.990 62.920 33.310 ;
        RECT 60.360 31.970 60.620 32.290 ;
        RECT 59.900 31.290 60.160 31.610 ;
        RECT 59.960 27.870 60.100 31.290 ;
        RECT 60.360 30.270 60.620 30.590 ;
        RECT 60.420 29.570 60.560 30.270 ;
        RECT 60.360 29.250 60.620 29.570 ;
        RECT 59.900 27.550 60.160 27.870 ;
        RECT 60.880 27.610 61.020 32.990 ;
        RECT 61.340 31.270 61.480 32.990 ;
        RECT 61.280 30.950 61.540 31.270 ;
        RECT 62.200 31.125 62.460 31.270 ;
        RECT 62.190 30.755 62.470 31.125 ;
        RECT 63.180 28.210 63.320 39.110 ;
        RECT 63.640 37.050 63.780 44.550 ;
        RECT 64.100 41.890 64.240 45.230 ;
        RECT 64.560 42.490 64.700 51.835 ;
        RECT 64.500 42.170 64.760 42.490 ;
        RECT 64.100 41.750 64.700 41.890 ;
        RECT 64.560 41.470 64.700 41.750 ;
        RECT 64.040 41.150 64.300 41.470 ;
        RECT 64.500 41.150 64.760 41.470 ;
        RECT 64.100 40.450 64.240 41.150 ;
        RECT 64.040 40.130 64.300 40.450 ;
        RECT 64.030 39.595 64.310 39.965 ;
        RECT 64.040 39.450 64.300 39.595 ;
        RECT 65.020 37.810 65.160 62.830 ;
        RECT 65.480 50.165 65.620 74.955 ;
        RECT 66.340 65.970 66.600 66.290 ;
        RECT 65.880 60.190 66.140 60.510 ;
        RECT 65.940 58.130 66.080 60.190 ;
        RECT 65.880 57.810 66.140 58.130 ;
        RECT 65.940 55.750 66.080 57.810 ;
        RECT 66.400 57.790 66.540 65.970 ;
        RECT 66.860 64.250 67.000 79.230 ;
        RECT 68.170 79.035 68.450 79.405 ;
        RECT 67.260 77.190 67.520 77.510 ;
        RECT 67.320 75.810 67.460 77.190 ;
        RECT 67.720 76.850 67.980 77.170 ;
        RECT 67.260 75.490 67.520 75.810 ;
        RECT 67.260 74.645 67.520 74.790 ;
        RECT 67.250 74.275 67.530 74.645 ;
        RECT 67.780 67.650 67.920 76.850 ;
        RECT 68.240 71.730 68.380 79.035 ;
        RECT 68.180 71.410 68.440 71.730 ;
        RECT 68.240 69.690 68.380 71.410 ;
        RECT 69.160 69.690 69.300 82.730 ;
        RECT 70.940 81.950 71.200 82.270 ;
        RECT 71.000 80.230 71.140 81.950 ;
        RECT 71.860 80.480 72.120 80.570 ;
        RECT 71.460 80.340 72.120 80.480 ;
        RECT 70.940 79.910 71.200 80.230 ;
        RECT 70.470 77.675 70.750 78.045 ;
        RECT 70.480 77.530 70.740 77.675 ;
        RECT 70.940 76.510 71.200 76.830 ;
        RECT 71.000 75.130 71.140 76.510 ;
        RECT 70.940 74.810 71.200 75.130 ;
        RECT 69.560 73.965 69.820 74.110 ;
        RECT 69.550 73.595 69.830 73.965 ;
        RECT 68.180 69.370 68.440 69.690 ;
        RECT 69.100 69.370 69.360 69.690 ;
        RECT 70.020 69.370 70.280 69.690 ;
        RECT 67.720 67.330 67.980 67.650 ;
        RECT 66.800 63.930 67.060 64.250 ;
        RECT 66.800 62.910 67.060 63.230 ;
        RECT 66.340 57.470 66.600 57.790 ;
        RECT 65.880 55.430 66.140 55.750 ;
        RECT 65.410 49.795 65.690 50.165 ;
        RECT 65.870 45.715 66.150 46.085 ;
        RECT 65.410 44.355 65.690 44.725 ;
        RECT 65.480 43.170 65.620 44.355 ;
        RECT 65.940 44.045 66.080 45.715 ;
        RECT 65.870 43.675 66.150 44.045 ;
        RECT 65.420 42.850 65.680 43.170 ;
        RECT 66.400 42.830 66.540 57.470 ;
        RECT 66.860 55.410 67.000 62.910 ;
        RECT 66.800 55.090 67.060 55.410 ;
        RECT 67.250 54.555 67.530 54.925 ;
        RECT 66.800 53.050 67.060 53.370 ;
        RECT 66.860 49.630 67.000 53.050 ;
        RECT 66.800 49.310 67.060 49.630 ;
        RECT 66.860 47.930 67.000 49.310 ;
        RECT 66.800 47.610 67.060 47.930 ;
        RECT 66.340 42.510 66.600 42.830 ;
        RECT 66.340 41.150 66.600 41.470 ;
        RECT 66.400 39.430 66.540 41.150 ;
        RECT 66.860 39.430 67.000 47.610 ;
        RECT 66.340 39.110 66.600 39.430 ;
        RECT 66.800 39.110 67.060 39.430 ;
        RECT 65.420 38.770 65.680 39.090 ;
        RECT 64.100 37.670 65.160 37.810 ;
        RECT 63.580 36.730 63.840 37.050 ;
        RECT 63.120 27.890 63.380 28.210 ;
        RECT 58.580 26.170 59.180 26.250 ;
        RECT 59.440 26.190 59.700 26.510 ;
        RECT 58.060 25.850 58.320 26.170 ;
        RECT 58.580 26.110 59.240 26.170 ;
        RECT 58.980 25.850 59.240 26.110 ;
        RECT 57.140 23.470 57.400 23.790 ;
        RECT 56.680 22.450 56.940 22.770 ;
        RECT 54.840 20.750 55.100 21.070 ;
        RECT 56.740 20.050 56.880 22.450 ;
        RECT 56.680 19.730 56.940 20.050 ;
        RECT 57.200 19.710 57.340 23.470 ;
        RECT 58.120 23.110 58.260 25.850 ;
        RECT 58.520 25.510 58.780 25.830 ;
        RECT 58.580 25.005 58.720 25.510 ;
        RECT 58.510 24.635 58.790 25.005 ;
        RECT 58.580 23.110 58.720 24.635 ;
        RECT 58.060 22.790 58.320 23.110 ;
        RECT 58.520 22.790 58.780 23.110 ;
        RECT 59.040 22.770 59.180 25.850 ;
        RECT 58.980 22.450 59.240 22.770 ;
        RECT 59.960 20.730 60.100 27.550 ;
        RECT 60.880 27.470 62.400 27.610 ;
        RECT 62.260 24.130 62.400 27.470 ;
        RECT 63.640 26.850 63.780 36.730 ;
        RECT 64.100 36.370 64.240 37.670 ;
        RECT 64.500 36.960 64.760 37.050 ;
        RECT 64.500 36.820 65.160 36.960 ;
        RECT 64.500 36.730 64.760 36.820 ;
        RECT 64.040 36.050 64.300 36.370 ;
        RECT 64.500 31.630 64.760 31.950 ;
        RECT 64.040 30.270 64.300 30.590 ;
        RECT 64.100 29.570 64.240 30.270 ;
        RECT 64.040 29.250 64.300 29.570 ;
        RECT 64.560 28.890 64.700 31.630 ;
        RECT 65.020 29.570 65.160 36.820 ;
        RECT 65.480 33.990 65.620 38.770 ;
        RECT 65.880 36.730 66.140 37.050 ;
        RECT 65.420 33.670 65.680 33.990 ;
        RECT 65.480 32.290 65.620 33.670 ;
        RECT 65.940 33.310 66.080 36.730 ;
        RECT 65.880 32.990 66.140 33.310 ;
        RECT 65.420 31.970 65.680 32.290 ;
        RECT 64.960 29.250 65.220 29.570 ;
        RECT 64.500 28.570 64.760 28.890 ;
        RECT 65.020 28.290 65.160 29.250 ;
        RECT 65.940 28.890 66.080 32.990 ;
        RECT 65.880 28.570 66.140 28.890 ;
        RECT 64.100 28.150 65.160 28.290 ;
        RECT 64.100 27.870 64.240 28.150 ;
        RECT 64.040 27.550 64.300 27.870 ;
        RECT 63.580 26.530 63.840 26.850 ;
        RECT 62.200 23.810 62.460 24.130 ;
        RECT 66.400 23.110 66.540 39.110 ;
        RECT 66.790 38.235 67.070 38.605 ;
        RECT 66.860 29.570 67.000 38.235 ;
        RECT 67.320 33.990 67.460 54.555 ;
        RECT 67.780 46.085 67.920 67.330 ;
        RECT 69.560 64.610 69.820 64.930 ;
        RECT 69.100 60.530 69.360 60.850 ;
        RECT 68.180 55.770 68.440 56.090 ;
        RECT 68.240 48.270 68.380 55.770 ;
        RECT 68.640 53.050 68.900 53.370 ;
        RECT 68.180 47.950 68.440 48.270 ;
        RECT 68.700 47.330 68.840 53.050 ;
        RECT 69.160 47.590 69.300 60.530 ;
        RECT 69.620 56.430 69.760 64.610 ;
        RECT 69.560 56.110 69.820 56.430 ;
        RECT 69.560 55.090 69.820 55.410 ;
        RECT 69.620 51.525 69.760 55.090 ;
        RECT 70.080 53.030 70.220 69.370 ;
        RECT 70.940 68.350 71.200 68.670 ;
        RECT 70.480 65.970 70.740 66.290 ;
        RECT 70.540 63.570 70.680 65.970 ;
        RECT 71.000 64.590 71.140 68.350 ;
        RECT 70.940 64.270 71.200 64.590 ;
        RECT 70.480 63.250 70.740 63.570 ;
        RECT 70.540 56.770 70.680 63.250 ;
        RECT 71.460 63.085 71.600 80.340 ;
        RECT 71.860 80.250 72.120 80.340 ;
        RECT 73.700 80.250 73.960 80.570 ;
        RECT 73.240 79.910 73.500 80.230 ;
        RECT 71.860 79.570 72.120 79.890 ;
        RECT 71.920 75.130 72.060 79.570 ;
        RECT 72.320 77.365 72.580 77.510 ;
        RECT 72.310 76.995 72.590 77.365 ;
        RECT 72.780 77.190 73.040 77.510 ;
        RECT 72.840 75.810 72.980 77.190 ;
        RECT 72.780 75.490 73.040 75.810 ;
        RECT 71.860 74.810 72.120 75.130 ;
        RECT 72.320 74.470 72.580 74.790 ;
        RECT 72.380 73.285 72.520 74.470 ;
        RECT 72.310 72.915 72.590 73.285 ;
        RECT 72.320 71.750 72.580 72.070 ;
        RECT 71.860 71.410 72.120 71.730 ;
        RECT 71.920 69.690 72.060 71.410 ;
        RECT 72.380 71.245 72.520 71.750 ;
        RECT 72.310 70.875 72.590 71.245 ;
        RECT 71.860 69.370 72.120 69.690 ;
        RECT 71.860 66.310 72.120 66.630 ;
        RECT 72.780 66.310 73.040 66.630 ;
        RECT 71.920 63.230 72.060 66.310 ;
        RECT 72.310 64.755 72.590 65.125 ;
        RECT 71.390 62.715 71.670 63.085 ;
        RECT 71.860 62.910 72.120 63.230 ;
        RECT 72.380 62.170 72.520 64.755 ;
        RECT 71.460 62.030 72.520 62.170 ;
        RECT 70.480 56.450 70.740 56.770 ;
        RECT 70.480 55.430 70.740 55.750 ;
        RECT 70.020 52.710 70.280 53.030 ;
        RECT 70.020 52.030 70.280 52.350 ;
        RECT 69.550 51.155 69.830 51.525 ;
        RECT 69.560 50.670 69.820 50.990 ;
        RECT 68.240 47.190 68.840 47.330 ;
        RECT 69.100 47.270 69.360 47.590 ;
        RECT 68.240 46.910 68.380 47.190 ;
        RECT 68.180 46.590 68.440 46.910 ;
        RECT 67.710 45.715 67.990 46.085 ;
        RECT 67.720 36.390 67.980 36.710 ;
        RECT 67.260 33.670 67.520 33.990 ;
        RECT 67.250 32.115 67.530 32.485 ;
        RECT 67.260 31.970 67.520 32.115 ;
        RECT 66.800 29.250 67.060 29.570 ;
        RECT 67.780 28.890 67.920 36.390 ;
        RECT 68.240 33.310 68.380 46.590 ;
        RECT 69.090 46.395 69.370 46.765 ;
        RECT 69.160 45.210 69.300 46.395 ;
        RECT 69.620 45.890 69.760 50.670 ;
        RECT 69.560 45.570 69.820 45.890 ;
        RECT 69.100 44.890 69.360 45.210 ;
        RECT 69.100 42.170 69.360 42.490 ;
        RECT 68.630 41.635 68.910 42.005 ;
        RECT 68.700 40.450 68.840 41.635 ;
        RECT 68.640 40.130 68.900 40.450 ;
        RECT 68.630 37.555 68.910 37.925 ;
        RECT 68.640 37.410 68.900 37.555 ;
        RECT 68.180 32.990 68.440 33.310 ;
        RECT 69.160 32.290 69.300 42.170 ;
        RECT 69.620 36.565 69.760 45.570 ;
        RECT 70.080 44.870 70.220 52.030 ;
        RECT 70.540 47.250 70.680 55.430 ;
        RECT 70.940 53.390 71.200 53.710 ;
        RECT 70.480 46.930 70.740 47.250 ;
        RECT 70.020 44.550 70.280 44.870 ;
        RECT 70.540 43.170 70.680 46.930 ;
        RECT 70.480 42.850 70.740 43.170 ;
        RECT 70.480 41.830 70.740 42.150 ;
        RECT 69.550 36.195 69.830 36.565 ;
        RECT 70.540 33.990 70.680 41.830 ;
        RECT 71.000 39.430 71.140 53.390 ;
        RECT 71.460 41.810 71.600 62.030 ;
        RECT 71.860 58.490 72.120 58.810 ;
        RECT 71.920 53.030 72.060 58.490 ;
        RECT 72.310 57.955 72.590 58.325 ;
        RECT 71.860 52.710 72.120 53.030 ;
        RECT 71.860 51.010 72.120 51.330 ;
        RECT 71.920 49.970 72.060 51.010 ;
        RECT 71.860 49.650 72.120 49.970 ;
        RECT 71.860 44.550 72.120 44.870 ;
        RECT 71.920 42.490 72.060 44.550 ;
        RECT 71.860 42.170 72.120 42.490 ;
        RECT 71.400 41.490 71.660 41.810 ;
        RECT 70.940 39.110 71.200 39.430 ;
        RECT 71.860 39.110 72.120 39.430 ;
        RECT 71.390 34.155 71.670 34.525 ;
        RECT 70.480 33.670 70.740 33.990 ;
        RECT 70.940 33.670 71.200 33.990 ;
        RECT 70.020 33.330 70.280 33.650 ;
        RECT 69.100 31.970 69.360 32.290 ;
        RECT 69.090 31.435 69.370 31.805 ;
        RECT 68.180 30.610 68.440 30.930 ;
        RECT 67.720 28.570 67.980 28.890 ;
        RECT 67.720 25.850 67.980 26.170 ;
        RECT 67.780 24.325 67.920 25.850 ;
        RECT 68.240 25.150 68.380 30.610 ;
        RECT 69.160 28.550 69.300 31.435 ;
        RECT 69.100 28.230 69.360 28.550 ;
        RECT 70.080 26.170 70.220 33.330 ;
        RECT 71.000 31.610 71.140 33.670 ;
        RECT 70.940 31.290 71.200 31.610 ;
        RECT 70.930 30.755 71.210 31.125 ;
        RECT 71.000 26.850 71.140 30.755 ;
        RECT 71.460 29.570 71.600 34.155 ;
        RECT 71.920 33.845 72.060 39.110 ;
        RECT 71.850 33.475 72.130 33.845 ;
        RECT 71.400 29.250 71.660 29.570 ;
        RECT 70.940 26.530 71.200 26.850 ;
        RECT 71.920 26.170 72.060 33.475 ;
        RECT 72.380 33.310 72.520 57.955 ;
        RECT 72.840 56.430 72.980 66.310 ;
        RECT 73.300 60.510 73.440 79.910 ;
        RECT 73.760 78.530 73.900 80.250 ;
        RECT 73.700 78.210 73.960 78.530 ;
        RECT 74.160 76.510 74.420 76.830 ;
        RECT 74.220 76.005 74.360 76.510 ;
        RECT 74.150 75.635 74.430 76.005 ;
        RECT 74.620 74.810 74.880 75.130 ;
        RECT 73.700 74.470 73.960 74.790 ;
        RECT 73.760 73.090 73.900 74.470 ;
        RECT 73.700 72.770 73.960 73.090 ;
        RECT 74.160 70.050 74.420 70.370 ;
        RECT 73.700 69.370 73.960 69.690 ;
        RECT 73.760 67.650 73.900 69.370 ;
        RECT 73.700 67.330 73.960 67.650 ;
        RECT 74.220 66.630 74.360 70.050 ;
        RECT 74.680 66.630 74.820 74.810 ;
        RECT 75.080 71.750 75.340 72.070 ;
        RECT 74.160 66.310 74.420 66.630 ;
        RECT 74.620 66.310 74.880 66.630 ;
        RECT 74.620 63.590 74.880 63.910 ;
        RECT 73.700 62.910 73.960 63.230 ;
        RECT 73.240 60.190 73.500 60.510 ;
        RECT 73.230 58.635 73.510 59.005 ;
        RECT 73.300 58.470 73.440 58.635 ;
        RECT 73.240 58.150 73.500 58.470 ;
        RECT 72.780 56.110 73.040 56.430 ;
        RECT 72.780 55.430 73.040 55.750 ;
        RECT 72.840 50.650 72.980 55.430 ;
        RECT 72.780 50.330 73.040 50.650 ;
        RECT 72.780 49.650 73.040 49.970 ;
        RECT 72.840 45.550 72.980 49.650 ;
        RECT 72.780 45.230 73.040 45.550 ;
        RECT 72.770 42.995 73.050 43.365 ;
        RECT 72.840 39.430 72.980 42.995 ;
        RECT 72.780 39.110 73.040 39.430 ;
        RECT 72.780 35.710 73.040 36.030 ;
        RECT 72.840 34.330 72.980 35.710 ;
        RECT 73.300 34.670 73.440 58.150 ;
        RECT 73.760 53.710 73.900 62.910 ;
        RECT 74.160 60.870 74.420 61.190 ;
        RECT 73.700 53.390 73.960 53.710 ;
        RECT 73.700 52.370 73.960 52.690 ;
        RECT 73.240 34.350 73.500 34.670 ;
        RECT 72.780 34.010 73.040 34.330 ;
        RECT 72.320 32.990 72.580 33.310 ;
        RECT 72.320 30.610 72.580 30.930 ;
        RECT 72.380 26.850 72.520 30.610 ;
        RECT 72.840 28.890 72.980 34.010 ;
        RECT 73.760 33.900 73.900 52.370 ;
        RECT 74.220 39.770 74.360 60.870 ;
        RECT 74.680 59.490 74.820 63.590 ;
        RECT 75.140 62.170 75.280 71.750 ;
        RECT 75.530 69.515 75.810 69.885 ;
        RECT 75.540 69.370 75.800 69.515 ;
        RECT 75.140 62.030 75.740 62.170 ;
        RECT 74.620 59.170 74.880 59.490 ;
        RECT 74.620 55.430 74.880 55.750 ;
        RECT 75.080 55.430 75.340 55.750 ;
        RECT 74.680 52.885 74.820 55.430 ;
        RECT 75.140 54.050 75.280 55.430 ;
        RECT 75.080 53.730 75.340 54.050 ;
        RECT 74.610 52.515 74.890 52.885 ;
        RECT 75.140 51.330 75.280 53.730 ;
        RECT 75.080 51.010 75.340 51.330 ;
        RECT 75.080 50.330 75.340 50.650 ;
        RECT 74.620 49.310 74.880 49.630 ;
        RECT 74.680 48.125 74.820 49.310 ;
        RECT 75.140 48.610 75.280 50.330 ;
        RECT 75.080 48.290 75.340 48.610 ;
        RECT 74.610 47.755 74.890 48.125 ;
        RECT 75.070 47.075 75.350 47.445 ;
        RECT 74.620 45.405 74.880 45.550 ;
        RECT 74.610 45.035 74.890 45.405 ;
        RECT 75.140 44.870 75.280 47.075 ;
        RECT 75.600 45.890 75.740 62.030 ;
        RECT 76.000 60.530 76.260 60.850 ;
        RECT 75.540 45.570 75.800 45.890 ;
        RECT 75.080 44.550 75.340 44.870 ;
        RECT 74.160 39.450 74.420 39.770 ;
        RECT 73.300 33.760 73.900 33.900 ;
        RECT 73.300 31.610 73.440 33.760 ;
        RECT 75.080 33.670 75.340 33.990 ;
        RECT 73.700 31.970 73.960 32.290 ;
        RECT 73.240 31.290 73.500 31.610 ;
        RECT 72.780 28.570 73.040 28.890 ;
        RECT 73.300 28.210 73.440 31.290 ;
        RECT 73.760 28.210 73.900 31.970 ;
        RECT 75.140 31.610 75.280 33.670 ;
        RECT 75.080 31.290 75.340 31.610 ;
        RECT 74.160 30.950 74.420 31.270 ;
        RECT 73.240 27.890 73.500 28.210 ;
        RECT 73.700 27.890 73.960 28.210 ;
        RECT 73.760 26.850 73.900 27.890 ;
        RECT 72.320 26.530 72.580 26.850 ;
        RECT 73.700 26.530 73.960 26.850 ;
        RECT 69.560 25.850 69.820 26.170 ;
        RECT 70.020 25.850 70.280 26.170 ;
        RECT 71.860 25.850 72.120 26.170 ;
        RECT 68.180 24.830 68.440 25.150 ;
        RECT 67.710 23.955 67.990 24.325 ;
        RECT 69.620 23.790 69.760 25.850 ;
        RECT 69.560 23.470 69.820 23.790 ;
        RECT 72.380 23.645 72.520 26.530 ;
        RECT 73.240 25.850 73.500 26.170 ;
        RECT 72.310 23.275 72.590 23.645 ;
        RECT 66.340 22.790 66.600 23.110 ;
        RECT 59.900 20.410 60.160 20.730 ;
        RECT 57.140 19.390 57.400 19.710 ;
        RECT 73.300 18.350 73.440 25.850 ;
        RECT 73.760 25.830 73.900 26.530 ;
        RECT 73.700 25.510 73.960 25.830 ;
        RECT 74.220 23.110 74.360 30.950 ;
        RECT 75.070 27.355 75.350 27.725 ;
        RECT 75.140 24.130 75.280 27.355 ;
        RECT 75.080 23.810 75.340 24.130 ;
        RECT 76.060 23.790 76.200 60.530 ;
        RECT 76.460 60.190 76.720 60.510 ;
        RECT 76.520 43.365 76.660 60.190 ;
        RECT 76.920 53.050 77.180 53.370 ;
        RECT 76.980 45.210 77.120 53.050 ;
        RECT 76.920 44.890 77.180 45.210 ;
        RECT 76.450 42.995 76.730 43.365 ;
        RECT 76.000 23.470 76.260 23.790 ;
        RECT 73.700 22.790 73.960 23.110 ;
        RECT 74.160 22.790 74.420 23.110 ;
        RECT 73.760 20.925 73.900 22.790 ;
        RECT 73.690 20.555 73.970 20.925 ;
        RECT 73.240 18.030 73.500 18.350 ;
        RECT 39.200 17.350 39.460 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 49.780 17.350 50.040 17.670 ;
        RECT 52.080 17.350 52.340 17.670 ;
        RECT 53.460 17.350 53.720 17.670 ;
        RECT 74.610 17.155 74.890 17.525 ;
        RECT 74.620 17.010 74.880 17.155 ;
        RECT 36.900 14.970 37.160 15.290 ;
        RECT 75.080 14.630 75.340 14.950 ;
        RECT 35.980 13.950 36.240 14.270 ;
        RECT 75.140 14.125 75.280 14.630 ;
        RECT 34.600 12.590 34.860 12.910 ;
        RECT 30.460 12.250 30.720 12.570 ;
        RECT 36.040 12.230 36.180 13.950 ;
        RECT 75.070 13.755 75.350 14.125 ;
        RECT 12.980 11.910 13.240 12.230 ;
        RECT 22.640 11.910 22.900 12.230 ;
        RECT 29.080 11.910 29.340 12.230 ;
        RECT 35.980 11.910 36.240 12.230 ;
        RECT 13.040 0.500 13.180 11.910 ;
        RECT 22.700 0.500 22.840 11.910 ;
        RECT 26.320 11.570 26.580 11.890 ;
        RECT 24.370 10.695 25.910 11.065 ;
        RECT 26.380 6.530 26.520 11.570 ;
        RECT 25.920 6.390 26.520 6.530 ;
        RECT 25.920 0.500 26.060 6.390 ;
        RECT 29.140 0.500 29.280 11.910 ;
        RECT 32.300 11.570 32.560 11.890 ;
        RECT 32.360 0.500 32.500 11.570 ;
        RECT 35.520 11.230 35.780 11.550 ;
        RECT 35.580 0.500 35.720 11.230 ;
      LAYER met3 ;
        RECT 18.925 92.290 19.255 92.305 ;
        RECT 18.925 91.990 81.850 92.290 ;
        RECT 18.925 91.975 19.255 91.990 ;
        RECT 33.390 90.930 33.770 90.940 ;
        RECT 80.565 90.930 80.895 90.945 ;
        RECT 33.390 90.630 80.895 90.930 ;
        RECT 33.390 90.620 33.770 90.630 ;
        RECT 80.565 90.615 80.895 90.630 ;
        RECT 40.750 89.570 41.130 89.580 ;
        RECT 77.345 89.570 77.675 89.585 ;
        RECT 40.750 89.270 77.675 89.570 ;
        RECT 40.750 89.260 41.130 89.270 ;
        RECT 77.345 89.255 77.675 89.270 ;
        RECT 39.830 88.890 40.210 88.900 ;
        RECT 39.830 88.590 81.850 88.890 ;
        RECT 39.830 88.580 40.210 88.590 ;
        RECT 67.685 88.210 68.015 88.225 ;
        RECT 68.350 88.210 68.730 88.220 ;
        RECT 67.685 87.910 68.730 88.210 ;
        RECT 67.685 87.895 68.015 87.910 ;
        RECT 68.350 87.900 68.730 87.910 ;
        RECT 44.430 87.530 44.810 87.540 ;
        RECT 64.465 87.530 64.795 87.545 ;
        RECT 44.430 87.230 64.795 87.530 ;
        RECT 44.430 87.220 44.810 87.230 ;
        RECT 64.465 87.215 64.795 87.230 ;
        RECT 20.305 86.850 20.635 86.865 ;
        RECT 29.045 86.850 29.375 86.865 ;
        RECT 20.305 86.550 29.375 86.850 ;
        RECT 20.305 86.535 20.635 86.550 ;
        RECT 29.045 86.535 29.375 86.550 ;
        RECT 45.350 86.850 45.730 86.860 ;
        RECT 70.905 86.850 71.235 86.865 ;
        RECT 45.350 86.550 71.235 86.850 ;
        RECT 45.350 86.540 45.730 86.550 ;
        RECT 70.905 86.535 71.235 86.550 ;
        RECT 30.630 85.490 31.010 85.500 ;
        RECT 30.630 85.190 81.850 85.490 ;
        RECT 30.630 85.180 31.010 85.190 ;
        RECT 22.605 84.810 22.935 84.825 ;
        RECT 28.790 84.810 29.170 84.820 ;
        RECT 22.605 84.510 29.170 84.810 ;
        RECT 22.605 84.495 22.935 84.510 ;
        RECT 28.790 84.500 29.170 84.510 ;
        RECT 14.785 84.130 15.115 84.145 ;
        RECT 38.705 84.130 39.035 84.145 ;
        RECT 14.785 83.830 39.035 84.130 ;
        RECT 14.785 83.815 15.115 83.830 ;
        RECT 38.705 83.815 39.035 83.830 ;
        RECT 12.945 83.460 13.275 83.465 ;
        RECT 12.945 83.450 13.530 83.460 ;
        RECT 12.720 83.150 13.530 83.450 ;
        RECT 12.945 83.140 13.530 83.150 ;
        RECT 25.825 83.450 26.155 83.465 ;
        RECT 27.870 83.450 28.250 83.460 ;
        RECT 25.825 83.150 28.250 83.450 ;
        RECT 12.945 83.135 13.275 83.140 ;
        RECT 25.825 83.135 26.155 83.150 ;
        RECT 27.870 83.140 28.250 83.150 ;
        RECT 60.070 83.450 60.450 83.460 ;
        RECT 61.245 83.450 61.575 83.465 ;
        RECT 60.070 83.150 61.575 83.450 ;
        RECT 60.070 83.140 60.450 83.150 ;
        RECT 61.245 83.135 61.575 83.150 ;
        RECT 12.485 82.770 12.815 82.785 ;
        RECT 12.485 82.470 26.600 82.770 ;
        RECT 12.485 82.455 12.815 82.470 ;
        RECT 6.045 82.090 6.375 82.105 ;
        RECT 0.500 81.790 6.375 82.090 ;
        RECT 6.045 81.775 6.375 81.790 ;
        RECT 24.350 81.435 25.930 81.765 ;
        RECT 26.300 81.410 26.600 82.470 ;
        RECT 38.705 82.090 39.035 82.105 ;
        RECT 38.705 81.790 81.850 82.090 ;
        RECT 38.705 81.775 39.035 81.790 ;
        RECT 26.950 81.410 27.330 81.420 ;
        RECT 66.305 81.410 66.635 81.425 ;
        RECT 26.300 81.110 66.635 81.410 ;
        RECT 26.950 81.100 27.330 81.110 ;
        RECT 66.305 81.095 66.635 81.110 ;
        RECT 23.525 80.730 23.855 80.745 ;
        RECT 38.705 80.730 39.035 80.745 ;
        RECT 23.525 80.430 39.035 80.730 ;
        RECT 23.525 80.415 23.855 80.430 ;
        RECT 38.705 80.415 39.035 80.430 ;
        RECT 53.425 80.730 53.755 80.745 ;
        RECT 58.485 80.730 58.815 80.745 ;
        RECT 53.425 80.430 58.815 80.730 ;
        RECT 53.425 80.415 53.755 80.430 ;
        RECT 58.485 80.415 58.815 80.430 ;
        RECT 11.105 80.050 11.435 80.065 ;
        RECT 41.925 80.050 42.255 80.065 ;
        RECT 11.105 79.750 42.255 80.050 ;
        RECT 11.105 79.735 11.435 79.750 ;
        RECT 41.925 79.735 42.255 79.750 ;
        RECT 27.205 79.370 27.535 79.385 ;
        RECT 45.145 79.370 45.475 79.385 ;
        RECT 68.145 79.370 68.475 79.385 ;
        RECT 27.205 79.070 68.475 79.370 ;
        RECT 27.205 79.055 27.535 79.070 ;
        RECT 45.145 79.055 45.475 79.070 ;
        RECT 68.145 79.055 68.475 79.070 ;
        RECT 21.050 78.715 22.630 79.045 ;
        RECT 6.505 78.690 6.835 78.705 ;
        RECT 0.500 78.390 6.835 78.690 ;
        RECT 6.505 78.375 6.835 78.390 ;
        RECT 24.905 78.690 25.235 78.705 ;
        RECT 55.265 78.690 55.595 78.705 ;
        RECT 24.905 78.390 55.595 78.690 ;
        RECT 24.905 78.375 25.235 78.390 ;
        RECT 55.265 78.375 55.595 78.390 ;
        RECT 58.230 78.690 58.610 78.700 ;
        RECT 59.865 78.690 60.195 78.705 ;
        RECT 58.230 78.390 60.195 78.690 ;
        RECT 58.230 78.380 58.610 78.390 ;
        RECT 59.865 78.375 60.195 78.390 ;
        RECT 63.750 78.690 64.130 78.700 ;
        RECT 63.750 78.390 81.850 78.690 ;
        RECT 63.750 78.380 64.130 78.390 ;
        RECT 18.670 78.010 19.050 78.020 ;
        RECT 19.385 78.010 19.715 78.025 ;
        RECT 18.670 77.710 19.715 78.010 ;
        RECT 18.670 77.700 19.050 77.710 ;
        RECT 19.385 77.695 19.715 77.710 ;
        RECT 22.145 78.010 22.475 78.025 ;
        RECT 31.550 78.010 31.930 78.020 ;
        RECT 22.145 77.710 31.930 78.010 ;
        RECT 22.145 77.695 22.475 77.710 ;
        RECT 31.550 77.700 31.930 77.710 ;
        RECT 32.725 78.010 33.055 78.025 ;
        RECT 70.445 78.010 70.775 78.025 ;
        RECT 32.725 77.710 70.775 78.010 ;
        RECT 32.725 77.695 33.055 77.710 ;
        RECT 70.445 77.695 70.775 77.710 ;
        RECT 15.245 77.330 15.575 77.345 ;
        RECT 39.165 77.330 39.495 77.345 ;
        RECT 72.285 77.330 72.615 77.345 ;
        RECT 15.245 77.030 39.495 77.330 ;
        RECT 15.245 77.015 15.575 77.030 ;
        RECT 39.165 77.015 39.495 77.030 ;
        RECT 39.870 77.030 72.615 77.330 ;
        RECT 15.705 76.650 16.035 76.665 ;
        RECT 17.750 76.650 18.130 76.660 ;
        RECT 15.705 76.350 18.130 76.650 ;
        RECT 15.705 76.335 16.035 76.350 ;
        RECT 17.750 76.340 18.130 76.350 ;
        RECT 21.225 76.650 21.555 76.665 ;
        RECT 23.270 76.650 23.650 76.660 ;
        RECT 21.225 76.350 23.650 76.650 ;
        RECT 21.225 76.335 21.555 76.350 ;
        RECT 23.270 76.340 23.650 76.350 ;
        RECT 30.425 76.650 30.755 76.665 ;
        RECT 32.470 76.650 32.850 76.660 ;
        RECT 30.425 76.350 32.850 76.650 ;
        RECT 30.425 76.335 30.755 76.350 ;
        RECT 32.470 76.340 32.850 76.350 ;
        RECT 35.230 76.650 35.610 76.660 ;
        RECT 37.785 76.650 38.115 76.665 ;
        RECT 39.870 76.650 40.170 77.030 ;
        RECT 72.285 77.015 72.615 77.030 ;
        RECT 35.230 76.350 38.115 76.650 ;
        RECT 35.230 76.340 35.610 76.350 ;
        RECT 37.785 76.335 38.115 76.350 ;
        RECT 38.950 76.350 40.170 76.650 ;
        RECT 60.785 76.660 61.115 76.665 ;
        RECT 60.785 76.650 61.370 76.660 ;
        RECT 60.785 76.350 61.570 76.650 ;
        RECT 24.350 75.995 25.930 76.325 ;
        RECT 15.705 75.970 16.035 75.985 ;
        RECT 21.685 75.970 22.015 75.985 ;
        RECT 15.705 75.670 22.015 75.970 ;
        RECT 15.705 75.655 16.035 75.670 ;
        RECT 21.685 75.655 22.015 75.670 ;
        RECT 38.245 75.970 38.575 75.985 ;
        RECT 38.950 75.970 39.250 76.350 ;
        RECT 60.785 76.340 61.370 76.350 ;
        RECT 60.785 76.335 61.115 76.340 ;
        RECT 38.245 75.670 39.250 75.970 ;
        RECT 39.625 75.970 39.955 75.985 ;
        RECT 40.750 75.970 41.130 75.980 ;
        RECT 39.625 75.670 41.130 75.970 ;
        RECT 38.245 75.655 38.575 75.670 ;
        RECT 39.625 75.655 39.955 75.670 ;
        RECT 40.750 75.660 41.130 75.670 ;
        RECT 55.265 75.970 55.595 75.985 ;
        RECT 74.125 75.970 74.455 75.985 ;
        RECT 55.265 75.670 74.455 75.970 ;
        RECT 55.265 75.655 55.595 75.670 ;
        RECT 74.125 75.655 74.455 75.670 ;
        RECT 6.045 75.290 6.375 75.305 ;
        RECT 0.500 74.990 6.375 75.290 ;
        RECT 6.045 74.975 6.375 74.990 ;
        RECT 12.945 75.290 13.275 75.305 ;
        RECT 24.445 75.290 24.775 75.305 ;
        RECT 12.945 74.990 24.775 75.290 ;
        RECT 12.945 74.975 13.275 74.990 ;
        RECT 24.445 74.975 24.775 74.990 ;
        RECT 25.365 75.290 25.695 75.305 ;
        RECT 29.505 75.290 29.835 75.305 ;
        RECT 62.625 75.290 62.955 75.305 ;
        RECT 25.365 74.990 62.955 75.290 ;
        RECT 25.365 74.975 25.695 74.990 ;
        RECT 29.505 74.975 29.835 74.990 ;
        RECT 62.625 74.975 62.955 74.990 ;
        RECT 65.385 75.290 65.715 75.305 ;
        RECT 65.385 74.990 81.850 75.290 ;
        RECT 65.385 74.975 65.715 74.990 ;
        RECT 13.405 74.610 13.735 74.625 ;
        RECT 26.285 74.610 26.615 74.625 ;
        RECT 39.165 74.610 39.495 74.625 ;
        RECT 46.065 74.620 46.395 74.625 ;
        RECT 46.065 74.610 46.650 74.620 ;
        RECT 67.225 74.610 67.555 74.625 ;
        RECT 13.405 74.310 39.495 74.610 ;
        RECT 45.660 74.310 67.555 74.610 ;
        RECT 13.405 74.295 13.735 74.310 ;
        RECT 26.285 74.295 26.615 74.310 ;
        RECT 39.165 74.295 39.495 74.310 ;
        RECT 46.065 74.300 46.650 74.310 ;
        RECT 46.065 74.295 46.395 74.300 ;
        RECT 67.225 74.295 67.555 74.310 ;
        RECT 23.525 73.930 23.855 73.945 ;
        RECT 46.080 73.930 46.380 74.295 ;
        RECT 23.525 73.630 46.380 73.930 ;
        RECT 60.785 73.930 61.115 73.945 ;
        RECT 69.525 73.930 69.855 73.945 ;
        RECT 60.785 73.630 69.855 73.930 ;
        RECT 23.525 73.615 23.855 73.630 ;
        RECT 60.785 73.615 61.115 73.630 ;
        RECT 69.525 73.615 69.855 73.630 ;
        RECT 21.050 73.275 22.630 73.605 ;
        RECT 48.825 73.250 49.155 73.265 ;
        RECT 72.285 73.250 72.615 73.265 ;
        RECT 48.825 72.950 72.615 73.250 ;
        RECT 48.825 72.935 49.155 72.950 ;
        RECT 72.285 72.935 72.615 72.950 ;
        RECT 17.085 72.570 17.415 72.585 ;
        RECT 32.725 72.570 33.055 72.585 ;
        RECT 17.085 72.270 33.055 72.570 ;
        RECT 17.085 72.255 17.415 72.270 ;
        RECT 32.725 72.255 33.055 72.270 ;
        RECT 3.745 71.890 4.075 71.905 ;
        RECT 0.500 71.590 4.075 71.890 ;
        RECT 3.745 71.575 4.075 71.590 ;
        RECT 15.705 71.890 16.035 71.905 ;
        RECT 40.750 71.890 41.130 71.900 ;
        RECT 15.705 71.590 36.490 71.890 ;
        RECT 15.705 71.575 16.035 71.590 ;
        RECT 11.565 71.210 11.895 71.225 ;
        RECT 12.230 71.210 12.610 71.220 ;
        RECT 11.565 70.910 12.610 71.210 ;
        RECT 11.565 70.895 11.895 70.910 ;
        RECT 12.230 70.900 12.610 70.910 ;
        RECT 12.945 71.210 13.275 71.225 ;
        RECT 17.085 71.210 17.415 71.225 ;
        RECT 20.305 71.210 20.635 71.225 ;
        RECT 12.945 70.910 20.635 71.210 ;
        RECT 12.945 70.895 13.275 70.910 ;
        RECT 17.085 70.895 17.415 70.910 ;
        RECT 20.305 70.895 20.635 70.910 ;
        RECT 29.045 71.210 29.375 71.225 ;
        RECT 30.425 71.210 30.755 71.225 ;
        RECT 29.045 70.910 30.755 71.210 ;
        RECT 29.045 70.895 29.375 70.910 ;
        RECT 30.425 70.895 30.755 70.910 ;
        RECT 31.345 71.210 31.675 71.225 ;
        RECT 35.025 71.210 35.355 71.225 ;
        RECT 36.190 71.220 36.490 71.590 ;
        RECT 40.750 71.590 81.850 71.890 ;
        RECT 40.750 71.580 41.130 71.590 ;
        RECT 31.345 70.910 35.355 71.210 ;
        RECT 31.345 70.895 31.675 70.910 ;
        RECT 35.025 70.895 35.355 70.910 ;
        RECT 36.150 71.210 36.530 71.220 ;
        RECT 38.245 71.210 38.575 71.225 ;
        RECT 36.150 70.910 38.575 71.210 ;
        RECT 36.150 70.900 36.530 70.910 ;
        RECT 38.245 70.895 38.575 70.910 ;
        RECT 39.165 71.210 39.495 71.225 ;
        RECT 72.285 71.210 72.615 71.225 ;
        RECT 39.165 70.910 72.615 71.210 ;
        RECT 39.165 70.895 39.495 70.910 ;
        RECT 72.285 70.895 72.615 70.910 ;
        RECT 24.350 70.555 25.930 70.885 ;
        RECT 9.265 70.530 9.595 70.545 ;
        RECT 11.310 70.530 11.690 70.540 ;
        RECT 21.685 70.530 22.015 70.545 ;
        RECT 9.265 70.230 22.015 70.530 ;
        RECT 9.265 70.215 9.595 70.230 ;
        RECT 11.310 70.220 11.690 70.230 ;
        RECT 21.685 70.215 22.015 70.230 ;
        RECT 26.745 70.530 27.075 70.545 ;
        RECT 44.685 70.530 45.015 70.545 ;
        RECT 26.745 70.230 45.015 70.530 ;
        RECT 26.745 70.215 27.075 70.230 ;
        RECT 44.685 70.215 45.015 70.230 ;
        RECT 15.245 69.850 15.575 69.865 ;
        RECT 22.145 69.850 22.475 69.865 ;
        RECT 26.285 69.850 26.615 69.865 ;
        RECT 15.245 69.550 26.615 69.850 ;
        RECT 15.245 69.535 15.575 69.550 ;
        RECT 22.145 69.535 22.475 69.550 ;
        RECT 26.285 69.535 26.615 69.550 ;
        RECT 27.665 69.850 27.995 69.865 ;
        RECT 34.565 69.850 34.895 69.865 ;
        RECT 27.665 69.550 34.895 69.850 ;
        RECT 27.665 69.535 27.995 69.550 ;
        RECT 34.565 69.535 34.895 69.550 ;
        RECT 43.765 69.850 44.095 69.865 ;
        RECT 58.945 69.850 59.275 69.865 ;
        RECT 43.765 69.550 59.275 69.850 ;
        RECT 43.765 69.535 44.095 69.550 ;
        RECT 58.945 69.535 59.275 69.550 ;
        RECT 64.465 69.850 64.795 69.865 ;
        RECT 75.505 69.850 75.835 69.865 ;
        RECT 64.465 69.550 75.835 69.850 ;
        RECT 64.465 69.535 64.795 69.550 ;
        RECT 75.505 69.535 75.835 69.550 ;
        RECT 16.830 69.170 17.210 69.180 ;
        RECT 18.465 69.170 18.795 69.185 ;
        RECT 16.830 68.870 18.795 69.170 ;
        RECT 16.830 68.860 17.210 68.870 ;
        RECT 18.465 68.855 18.795 68.870 ;
        RECT 20.765 69.170 21.095 69.185 ;
        RECT 29.710 69.170 30.090 69.180 ;
        RECT 32.725 69.170 33.055 69.185 ;
        RECT 20.765 68.870 29.360 69.170 ;
        RECT 20.765 68.855 21.095 68.870 ;
        RECT 5.585 68.490 5.915 68.505 ;
        RECT 0.500 68.190 5.915 68.490 ;
        RECT 29.060 68.490 29.360 68.870 ;
        RECT 29.710 68.870 33.055 69.170 ;
        RECT 29.710 68.860 30.090 68.870 ;
        RECT 32.725 68.855 33.055 68.870 ;
        RECT 46.065 69.180 46.395 69.185 ;
        RECT 46.065 69.170 46.650 69.180 ;
        RECT 46.065 68.870 46.850 69.170 ;
        RECT 46.065 68.860 46.650 68.870 ;
        RECT 46.065 68.855 46.395 68.860 ;
        RECT 32.265 68.490 32.595 68.505 ;
        RECT 37.325 68.490 37.655 68.505 ;
        RECT 41.005 68.490 41.335 68.505 ;
        RECT 29.060 68.190 34.650 68.490 ;
        RECT 5.585 68.175 5.915 68.190 ;
        RECT 32.265 68.175 32.595 68.190 ;
        RECT 21.050 67.835 22.630 68.165 ;
        RECT 19.845 67.820 20.175 67.825 ;
        RECT 19.590 67.810 20.175 67.820 ;
        RECT 27.665 67.810 27.995 67.825 ;
        RECT 19.390 67.510 20.175 67.810 ;
        RECT 19.590 67.500 20.175 67.510 ;
        RECT 19.845 67.495 20.175 67.500 ;
        RECT 25.380 67.510 27.995 67.810 ;
        RECT 34.350 67.810 34.650 68.190 ;
        RECT 37.325 68.190 41.335 68.490 ;
        RECT 37.325 68.175 37.655 68.190 ;
        RECT 41.005 68.175 41.335 68.190 ;
        RECT 63.545 68.490 63.875 68.505 ;
        RECT 63.545 68.190 81.850 68.490 ;
        RECT 63.545 68.175 63.875 68.190 ;
        RECT 56.185 67.810 56.515 67.825 ;
        RECT 34.350 67.510 56.515 67.810 ;
        RECT 16.625 67.130 16.955 67.145 ;
        RECT 25.380 67.130 25.680 67.510 ;
        RECT 27.665 67.495 27.995 67.510 ;
        RECT 56.185 67.495 56.515 67.510 ;
        RECT 16.625 66.830 25.680 67.130 ;
        RECT 26.285 67.130 26.615 67.145 ;
        RECT 30.630 67.130 31.010 67.140 ;
        RECT 26.285 66.830 31.010 67.130 ;
        RECT 16.625 66.815 16.955 66.830 ;
        RECT 26.285 66.815 26.615 66.830 ;
        RECT 30.630 66.820 31.010 66.830 ;
        RECT 36.405 67.130 36.735 67.145 ;
        RECT 44.225 67.130 44.555 67.145 ;
        RECT 57.105 67.130 57.435 67.145 ;
        RECT 36.405 66.830 44.555 67.130 ;
        RECT 36.405 66.815 36.735 66.830 ;
        RECT 44.225 66.815 44.555 66.830 ;
        RECT 45.160 66.830 57.435 67.130 ;
        RECT 14.785 66.450 15.115 66.465 ;
        RECT 22.605 66.450 22.935 66.465 ;
        RECT 14.785 66.150 22.935 66.450 ;
        RECT 14.785 66.135 15.115 66.150 ;
        RECT 22.605 66.135 22.935 66.150 ;
        RECT 23.525 66.450 23.855 66.465 ;
        RECT 45.160 66.450 45.460 66.830 ;
        RECT 57.105 66.815 57.435 66.830 ;
        RECT 23.525 66.150 45.460 66.450 ;
        RECT 48.110 66.450 48.490 66.460 ;
        RECT 53.885 66.450 54.215 66.465 ;
        RECT 48.110 66.150 54.215 66.450 ;
        RECT 23.525 66.135 23.855 66.150 ;
        RECT 48.110 66.140 48.490 66.150 ;
        RECT 53.885 66.135 54.215 66.150 ;
        RECT 12.485 65.770 12.815 65.785 ;
        RECT 16.625 65.770 16.955 65.785 ;
        RECT 12.485 65.470 16.955 65.770 ;
        RECT 12.485 65.455 12.815 65.470 ;
        RECT 16.625 65.455 16.955 65.470 ;
        RECT 17.545 65.770 17.875 65.785 ;
        RECT 22.145 65.770 22.475 65.785 ;
        RECT 17.545 65.470 22.475 65.770 ;
        RECT 17.545 65.455 17.875 65.470 ;
        RECT 22.145 65.455 22.475 65.470 ;
        RECT 30.885 65.770 31.215 65.785 ;
        RECT 58.025 65.770 58.355 65.785 ;
        RECT 30.885 65.470 58.355 65.770 ;
        RECT 30.885 65.455 31.215 65.470 ;
        RECT 58.025 65.455 58.355 65.470 ;
        RECT 24.350 65.115 25.930 65.445 ;
        RECT 4.665 65.090 4.995 65.105 ;
        RECT 0.500 64.790 4.995 65.090 ;
        RECT 4.665 64.775 4.995 64.790 ;
        RECT 16.625 65.090 16.955 65.105 ;
        RECT 23.065 65.090 23.395 65.105 ;
        RECT 16.625 64.790 23.395 65.090 ;
        RECT 16.625 64.775 16.955 64.790 ;
        RECT 23.065 64.775 23.395 64.790 ;
        RECT 26.285 65.090 26.615 65.105 ;
        RECT 29.965 65.090 30.295 65.105 ;
        RECT 42.385 65.090 42.715 65.105 ;
        RECT 72.285 65.090 72.615 65.105 ;
        RECT 26.285 64.790 48.450 65.090 ;
        RECT 26.285 64.775 26.615 64.790 ;
        RECT 29.965 64.775 30.295 64.790 ;
        RECT 42.385 64.775 42.715 64.790 ;
        RECT 13.405 64.410 13.735 64.425 ;
        RECT 32.265 64.410 32.595 64.425 ;
        RECT 39.165 64.410 39.495 64.425 ;
        RECT 13.405 64.110 31.890 64.410 ;
        RECT 13.405 64.095 13.735 64.110 ;
        RECT 9.725 63.730 10.055 63.745 ;
        RECT 13.420 63.730 13.720 64.095 ;
        RECT 9.725 63.430 13.720 63.730 ;
        RECT 23.525 63.730 23.855 63.745 ;
        RECT 26.950 63.730 27.330 63.740 ;
        RECT 23.525 63.430 27.330 63.730 ;
        RECT 9.725 63.415 10.055 63.430 ;
        RECT 23.525 63.415 23.855 63.430 ;
        RECT 26.950 63.420 27.330 63.430 ;
        RECT 28.125 63.730 28.455 63.745 ;
        RECT 30.630 63.730 31.010 63.740 ;
        RECT 28.125 63.430 31.010 63.730 ;
        RECT 31.590 63.730 31.890 64.110 ;
        RECT 32.265 64.110 39.495 64.410 ;
        RECT 32.265 64.095 32.595 64.110 ;
        RECT 39.165 64.095 39.495 64.110 ;
        RECT 32.725 63.730 33.055 63.745 ;
        RECT 31.590 63.430 33.055 63.730 ;
        RECT 28.125 63.415 28.455 63.430 ;
        RECT 30.630 63.420 31.010 63.430 ;
        RECT 32.725 63.415 33.055 63.430 ;
        RECT 6.965 63.050 7.295 63.065 ;
        RECT 18.925 63.050 19.255 63.065 ;
        RECT 6.965 62.750 19.255 63.050 ;
        RECT 6.965 62.735 7.295 62.750 ;
        RECT 18.925 62.735 19.255 62.750 ;
        RECT 24.445 63.050 24.775 63.065 ;
        RECT 46.525 63.050 46.855 63.065 ;
        RECT 24.445 62.750 46.855 63.050 ;
        RECT 48.150 63.050 48.450 64.790 ;
        RECT 72.285 64.790 81.850 65.090 ;
        RECT 72.285 64.775 72.615 64.790 ;
        RECT 71.365 63.050 71.695 63.065 ;
        RECT 48.150 62.750 71.695 63.050 ;
        RECT 24.445 62.735 24.775 62.750 ;
        RECT 46.525 62.735 46.855 62.750 ;
        RECT 71.365 62.735 71.695 62.750 ;
        RECT 21.050 62.395 22.630 62.725 ;
        RECT 24.905 62.370 25.235 62.385 ;
        RECT 26.285 62.370 26.615 62.385 ;
        RECT 24.905 62.070 26.615 62.370 ;
        RECT 24.905 62.055 25.235 62.070 ;
        RECT 26.285 62.055 26.615 62.070 ;
        RECT 3.745 61.690 4.075 61.705 ;
        RECT 0.500 61.390 4.075 61.690 ;
        RECT 3.745 61.375 4.075 61.390 ;
        RECT 14.325 61.690 14.655 61.705 ;
        RECT 14.990 61.690 15.370 61.700 ;
        RECT 22.145 61.690 22.475 61.705 ;
        RECT 14.325 61.390 15.370 61.690 ;
        RECT 14.325 61.375 14.655 61.390 ;
        RECT 14.990 61.380 15.370 61.390 ;
        RECT 15.720 61.390 22.475 61.690 ;
        RECT 15.720 61.010 16.020 61.390 ;
        RECT 22.145 61.375 22.475 61.390 ;
        RECT 25.825 61.690 26.155 61.705 ;
        RECT 27.870 61.690 28.250 61.700 ;
        RECT 25.825 61.390 28.250 61.690 ;
        RECT 25.825 61.375 26.155 61.390 ;
        RECT 27.870 61.380 28.250 61.390 ;
        RECT 29.505 61.690 29.835 61.705 ;
        RECT 29.505 61.390 81.850 61.690 ;
        RECT 29.505 61.375 29.835 61.390 ;
        RECT 9.740 60.710 16.020 61.010 ;
        RECT 20.765 61.010 21.095 61.025 ;
        RECT 32.265 61.010 32.595 61.025 ;
        RECT 20.765 60.710 32.595 61.010 ;
        RECT 9.740 60.345 10.040 60.710 ;
        RECT 20.765 60.695 21.095 60.710 ;
        RECT 32.265 60.695 32.595 60.710 ;
        RECT 9.725 60.015 10.055 60.345 ;
        RECT 10.645 60.015 10.975 60.345 ;
        RECT 15.910 60.330 16.290 60.340 ;
        RECT 19.845 60.330 20.175 60.345 ;
        RECT 15.910 60.030 20.175 60.330 ;
        RECT 15.910 60.020 16.290 60.030 ;
        RECT 19.845 60.015 20.175 60.030 ;
        RECT 21.685 60.330 22.015 60.345 ;
        RECT 23.065 60.330 23.395 60.345 ;
        RECT 21.685 60.030 23.395 60.330 ;
        RECT 21.685 60.015 22.015 60.030 ;
        RECT 23.065 60.015 23.395 60.030 ;
        RECT 30.885 60.330 31.215 60.345 ;
        RECT 33.390 60.330 33.770 60.340 ;
        RECT 30.885 60.030 33.770 60.330 ;
        RECT 30.885 60.015 31.215 60.030 ;
        RECT 33.390 60.020 33.770 60.030 ;
        RECT 10.660 59.650 10.960 60.015 ;
        RECT 24.350 59.675 25.930 60.005 ;
        RECT 20.765 59.650 21.095 59.665 ;
        RECT 10.660 59.350 21.095 59.650 ;
        RECT 16.640 58.985 16.940 59.350 ;
        RECT 20.765 59.335 21.095 59.350 ;
        RECT 26.285 59.650 26.615 59.665 ;
        RECT 29.045 59.650 29.375 59.665 ;
        RECT 26.285 59.350 29.375 59.650 ;
        RECT 26.285 59.335 26.615 59.350 ;
        RECT 29.045 59.335 29.375 59.350 ;
        RECT 31.550 59.650 31.930 59.660 ;
        RECT 32.265 59.650 32.595 59.665 ;
        RECT 31.550 59.350 32.595 59.650 ;
        RECT 31.550 59.340 31.930 59.350 ;
        RECT 32.265 59.335 32.595 59.350 ;
        RECT 9.725 58.970 10.055 58.985 ;
        RECT 14.785 58.970 15.115 58.985 ;
        RECT 9.725 58.670 15.115 58.970 ;
        RECT 9.725 58.655 10.055 58.670 ;
        RECT 14.785 58.655 15.115 58.670 ;
        RECT 16.625 58.655 16.955 58.985 ;
        RECT 27.665 58.970 27.995 58.985 ;
        RECT 53.425 58.970 53.755 58.985 ;
        RECT 73.205 58.970 73.535 58.985 ;
        RECT 27.665 58.670 48.450 58.970 ;
        RECT 27.665 58.655 27.995 58.670 ;
        RECT 3.745 58.290 4.075 58.305 ;
        RECT 14.785 58.300 15.115 58.305 ;
        RECT 14.785 58.290 15.370 58.300 ;
        RECT 0.500 57.990 4.075 58.290 ;
        RECT 14.560 57.990 15.370 58.290 ;
        RECT 3.745 57.975 4.075 57.990 ;
        RECT 14.785 57.980 15.370 57.990 ;
        RECT 17.750 58.290 18.130 58.300 ;
        RECT 36.405 58.290 36.735 58.305 ;
        RECT 17.750 57.990 36.735 58.290 ;
        RECT 17.750 57.980 18.130 57.990 ;
        RECT 14.785 57.975 15.115 57.980 ;
        RECT 36.405 57.975 36.735 57.990 ;
        RECT 12.945 57.610 13.275 57.625 ;
        RECT 19.845 57.610 20.175 57.625 ;
        RECT 12.945 57.310 20.175 57.610 ;
        RECT 12.945 57.295 13.275 57.310 ;
        RECT 19.845 57.295 20.175 57.310 ;
        RECT 23.985 57.610 24.315 57.625 ;
        RECT 28.790 57.610 29.170 57.620 ;
        RECT 23.985 57.310 29.170 57.610 ;
        RECT 23.985 57.295 24.315 57.310 ;
        RECT 28.790 57.300 29.170 57.310 ;
        RECT 29.710 57.610 30.090 57.620 ;
        RECT 31.805 57.610 32.135 57.625 ;
        RECT 33.390 57.610 33.770 57.620 ;
        RECT 29.710 57.310 33.770 57.610 ;
        RECT 29.710 57.300 30.090 57.310 ;
        RECT 31.805 57.295 32.135 57.310 ;
        RECT 33.390 57.300 33.770 57.310 ;
        RECT 21.050 56.955 22.630 57.285 ;
        RECT 10.185 56.930 10.515 56.945 ;
        RECT 18.005 56.930 18.335 56.945 ;
        RECT 18.925 56.940 19.255 56.945 ;
        RECT 10.185 56.630 18.335 56.930 ;
        RECT 10.185 56.615 10.515 56.630 ;
        RECT 18.005 56.615 18.335 56.630 ;
        RECT 18.670 56.930 19.255 56.940 ;
        RECT 26.950 56.930 27.330 56.940 ;
        RECT 27.665 56.930 27.995 56.945 ;
        RECT 18.670 56.630 19.480 56.930 ;
        RECT 26.950 56.630 27.995 56.930 ;
        RECT 18.670 56.620 19.255 56.630 ;
        RECT 26.950 56.620 27.330 56.630 ;
        RECT 18.925 56.615 19.255 56.620 ;
        RECT 27.665 56.615 27.995 56.630 ;
        RECT 29.045 56.930 29.375 56.945 ;
        RECT 34.310 56.930 34.690 56.940 ;
        RECT 29.045 56.630 34.690 56.930 ;
        RECT 48.150 56.930 48.450 58.670 ;
        RECT 53.425 58.670 73.535 58.970 ;
        RECT 53.425 58.655 53.755 58.670 ;
        RECT 73.205 58.655 73.535 58.670 ;
        RECT 72.285 58.290 72.615 58.305 ;
        RECT 72.285 57.990 81.850 58.290 ;
        RECT 72.285 57.975 72.615 57.990 ;
        RECT 64.465 56.930 64.795 56.945 ;
        RECT 48.150 56.630 64.795 56.930 ;
        RECT 29.045 56.615 29.375 56.630 ;
        RECT 34.310 56.620 34.690 56.630 ;
        RECT 64.465 56.615 64.795 56.630 ;
        RECT 9.265 56.250 9.595 56.265 ;
        RECT 17.545 56.250 17.875 56.265 ;
        RECT 9.265 55.950 17.875 56.250 ;
        RECT 9.265 55.935 9.595 55.950 ;
        RECT 17.545 55.935 17.875 55.950 ;
        RECT 21.225 56.250 21.555 56.265 ;
        RECT 36.405 56.250 36.735 56.265 ;
        RECT 21.225 55.950 36.735 56.250 ;
        RECT 21.225 55.935 21.555 55.950 ;
        RECT 36.405 55.935 36.735 55.950 ;
        RECT 15.245 55.570 15.575 55.585 ;
        RECT 18.925 55.570 19.255 55.585 ;
        RECT 37.785 55.570 38.115 55.585 ;
        RECT 15.245 55.270 38.115 55.570 ;
        RECT 15.245 55.255 15.575 55.270 ;
        RECT 18.925 55.255 19.255 55.270 ;
        RECT 37.785 55.255 38.115 55.270 ;
        RECT 3.745 54.890 4.075 54.905 ;
        RECT 0.500 54.590 4.075 54.890 ;
        RECT 3.745 54.575 4.075 54.590 ;
        RECT 14.070 54.890 14.450 54.900 ;
        RECT 16.625 54.890 16.955 54.905 ;
        RECT 14.070 54.590 16.955 54.890 ;
        RECT 14.070 54.580 14.450 54.590 ;
        RECT 16.625 54.575 16.955 54.590 ;
        RECT 26.745 54.890 27.075 54.905 ;
        RECT 35.230 54.890 35.610 54.900 ;
        RECT 26.745 54.590 35.610 54.890 ;
        RECT 26.745 54.575 27.075 54.590 ;
        RECT 35.230 54.580 35.610 54.590 ;
        RECT 36.405 54.890 36.735 54.905 ;
        RECT 39.830 54.890 40.210 54.900 ;
        RECT 36.405 54.590 40.210 54.890 ;
        RECT 36.405 54.575 36.735 54.590 ;
        RECT 39.830 54.580 40.210 54.590 ;
        RECT 67.225 54.890 67.555 54.905 ;
        RECT 67.225 54.590 81.850 54.890 ;
        RECT 67.225 54.575 67.555 54.590 ;
        RECT 24.350 54.235 25.930 54.565 ;
        RECT 11.310 54.210 11.690 54.220 ;
        RECT 15.245 54.210 15.575 54.225 ;
        RECT 11.310 53.910 15.575 54.210 ;
        RECT 11.310 53.900 11.690 53.910 ;
        RECT 15.245 53.895 15.575 53.910 ;
        RECT 19.590 54.210 19.970 54.220 ;
        RECT 20.305 54.210 20.635 54.225 ;
        RECT 19.590 53.910 20.635 54.210 ;
        RECT 19.590 53.900 19.970 53.910 ;
        RECT 20.305 53.895 20.635 53.910 ;
        RECT 50.205 54.210 50.535 54.225 ;
        RECT 56.185 54.210 56.515 54.225 ;
        RECT 50.205 53.910 56.515 54.210 ;
        RECT 50.205 53.895 50.535 53.910 ;
        RECT 56.185 53.895 56.515 53.910 ;
        RECT 10.185 53.530 10.515 53.545 ;
        RECT 35.945 53.530 36.275 53.545 ;
        RECT 10.185 53.230 36.275 53.530 ;
        RECT 10.185 53.215 10.515 53.230 ;
        RECT 35.945 53.215 36.275 53.230 ;
        RECT 38.705 53.530 39.035 53.545 ;
        RECT 47.905 53.530 48.235 53.545 ;
        RECT 38.705 53.230 48.235 53.530 ;
        RECT 38.705 53.215 39.035 53.230 ;
        RECT 47.905 53.215 48.235 53.230 ;
        RECT 48.825 53.530 49.155 53.545 ;
        RECT 52.965 53.530 53.295 53.545 ;
        RECT 48.825 53.230 53.295 53.530 ;
        RECT 48.825 53.215 49.155 53.230 ;
        RECT 52.965 53.215 53.295 53.230 ;
        RECT 20.305 52.850 20.635 52.865 ;
        RECT 28.585 52.850 28.915 52.865 ;
        RECT 20.305 52.550 28.915 52.850 ;
        RECT 20.305 52.535 20.635 52.550 ;
        RECT 28.585 52.535 28.915 52.550 ;
        RECT 41.465 52.850 41.795 52.865 ;
        RECT 57.105 52.850 57.435 52.865 ;
        RECT 74.585 52.850 74.915 52.865 ;
        RECT 41.465 52.550 53.050 52.850 ;
        RECT 41.465 52.535 41.795 52.550 ;
        RECT 25.825 52.170 26.155 52.185 ;
        RECT 27.870 52.170 28.250 52.180 ;
        RECT 25.825 51.870 28.250 52.170 ;
        RECT 25.825 51.855 26.155 51.870 ;
        RECT 27.870 51.860 28.250 51.870 ;
        RECT 43.765 52.170 44.095 52.185 ;
        RECT 46.525 52.170 46.855 52.185 ;
        RECT 52.045 52.170 52.375 52.185 ;
        RECT 43.765 51.870 52.375 52.170 ;
        RECT 52.750 52.170 53.050 52.550 ;
        RECT 57.105 52.550 74.915 52.850 ;
        RECT 57.105 52.535 57.435 52.550 ;
        RECT 74.585 52.535 74.915 52.550 ;
        RECT 64.465 52.170 64.795 52.185 ;
        RECT 52.750 51.870 64.795 52.170 ;
        RECT 43.765 51.855 44.095 51.870 ;
        RECT 46.525 51.855 46.855 51.870 ;
        RECT 52.045 51.855 52.375 51.870 ;
        RECT 64.465 51.855 64.795 51.870 ;
        RECT 21.050 51.515 22.630 51.845 ;
        RECT 15.705 51.500 16.035 51.505 ;
        RECT 15.705 51.490 16.290 51.500 ;
        RECT 52.965 51.490 53.295 51.505 ;
        RECT 63.545 51.490 63.875 51.505 ;
        RECT 15.480 51.190 16.290 51.490 ;
        RECT 15.705 51.180 16.290 51.190 ;
        RECT 23.310 51.190 63.875 51.490 ;
        RECT 15.705 51.175 16.035 51.180 ;
        RECT 15.245 50.810 15.575 50.825 ;
        RECT 23.310 50.810 23.610 51.190 ;
        RECT 52.965 51.175 53.295 51.190 ;
        RECT 63.545 51.175 63.875 51.190 ;
        RECT 69.525 51.490 69.855 51.505 ;
        RECT 69.525 51.190 81.850 51.490 ;
        RECT 69.525 51.175 69.855 51.190 ;
        RECT 15.245 50.510 23.610 50.810 ;
        RECT 27.205 50.810 27.535 50.825 ;
        RECT 35.485 50.810 35.815 50.825 ;
        RECT 51.125 50.810 51.455 50.825 ;
        RECT 27.205 50.510 51.455 50.810 ;
        RECT 15.245 50.495 15.575 50.510 ;
        RECT 27.205 50.495 27.535 50.510 ;
        RECT 35.485 50.495 35.815 50.510 ;
        RECT 51.125 50.495 51.455 50.510 ;
        RECT 16.830 50.130 17.210 50.140 ;
        RECT 20.765 50.130 21.095 50.145 ;
        RECT 25.365 50.130 25.695 50.145 ;
        RECT 16.830 49.830 25.695 50.130 ;
        RECT 16.830 49.820 17.210 49.830 ;
        RECT 20.765 49.815 21.095 49.830 ;
        RECT 25.365 49.815 25.695 49.830 ;
        RECT 26.285 50.130 26.615 50.145 ;
        RECT 36.405 50.130 36.735 50.145 ;
        RECT 38.245 50.130 38.575 50.145 ;
        RECT 26.285 49.830 38.575 50.130 ;
        RECT 26.285 49.815 26.615 49.830 ;
        RECT 36.405 49.815 36.735 49.830 ;
        RECT 38.245 49.815 38.575 49.830 ;
        RECT 42.385 50.130 42.715 50.145 ;
        RECT 65.385 50.130 65.715 50.145 ;
        RECT 42.385 49.830 65.715 50.130 ;
        RECT 42.385 49.815 42.715 49.830 ;
        RECT 65.385 49.815 65.715 49.830 ;
        RECT 43.305 49.450 43.635 49.465 ;
        RECT 52.965 49.450 53.295 49.465 ;
        RECT 43.305 49.150 53.295 49.450 ;
        RECT 43.305 49.135 43.635 49.150 ;
        RECT 52.965 49.135 53.295 49.150 ;
        RECT 24.350 48.795 25.930 49.125 ;
        RECT 15.705 48.770 16.035 48.785 ;
        RECT 23.270 48.770 23.650 48.780 ;
        RECT 15.705 48.470 23.650 48.770 ;
        RECT 15.705 48.455 16.035 48.470 ;
        RECT 23.270 48.460 23.650 48.470 ;
        RECT 38.705 48.770 39.035 48.785 ;
        RECT 63.750 48.770 64.130 48.780 ;
        RECT 38.705 48.470 46.610 48.770 ;
        RECT 38.705 48.455 39.035 48.470 ;
        RECT 0.985 48.090 1.315 48.105 ;
        RECT 0.500 47.790 1.315 48.090 ;
        RECT 0.985 47.775 1.315 47.790 ;
        RECT 32.470 48.090 32.850 48.100 ;
        RECT 35.485 48.090 35.815 48.105 ;
        RECT 32.470 47.790 35.815 48.090 ;
        RECT 32.470 47.780 32.850 47.790 ;
        RECT 35.485 47.775 35.815 47.790 ;
        RECT 36.150 48.090 36.530 48.100 ;
        RECT 38.705 48.090 39.035 48.105 ;
        RECT 41.005 48.100 41.335 48.105 ;
        RECT 40.750 48.090 41.335 48.100 ;
        RECT 36.150 47.790 39.035 48.090 ;
        RECT 40.550 47.790 41.335 48.090 ;
        RECT 36.150 47.780 36.530 47.790 ;
        RECT 38.705 47.775 39.035 47.790 ;
        RECT 40.750 47.780 41.335 47.790 ;
        RECT 41.005 47.775 41.335 47.780 ;
        RECT 43.765 48.090 44.095 48.105 ;
        RECT 45.145 48.100 45.475 48.105 ;
        RECT 44.430 48.090 44.810 48.100 ;
        RECT 43.765 47.790 44.810 48.090 ;
        RECT 43.765 47.775 44.095 47.790 ;
        RECT 44.430 47.780 44.810 47.790 ;
        RECT 45.145 48.090 45.730 48.100 ;
        RECT 45.145 47.790 45.930 48.090 ;
        RECT 45.145 47.780 45.730 47.790 ;
        RECT 45.145 47.775 45.475 47.780 ;
        RECT 12.230 47.410 12.610 47.420 ;
        RECT 13.405 47.410 13.735 47.425 ;
        RECT 12.230 47.110 13.735 47.410 ;
        RECT 12.230 47.100 12.610 47.110 ;
        RECT 13.405 47.095 13.735 47.110 ;
        RECT 30.630 47.410 31.010 47.420 ;
        RECT 41.005 47.410 41.335 47.425 ;
        RECT 30.630 47.110 41.335 47.410 ;
        RECT 46.310 47.410 46.610 48.470 ;
        RECT 48.150 48.470 64.130 48.770 ;
        RECT 47.445 48.090 47.775 48.105 ;
        RECT 48.150 48.090 48.450 48.470 ;
        RECT 63.750 48.460 64.130 48.470 ;
        RECT 47.445 47.790 48.450 48.090 ;
        RECT 74.585 48.090 74.915 48.105 ;
        RECT 74.585 47.790 81.850 48.090 ;
        RECT 47.445 47.775 47.775 47.790 ;
        RECT 74.585 47.775 74.915 47.790 ;
        RECT 75.045 47.410 75.375 47.425 ;
        RECT 46.310 47.110 75.375 47.410 ;
        RECT 30.630 47.100 31.010 47.110 ;
        RECT 41.005 47.095 41.335 47.110 ;
        RECT 75.045 47.095 75.375 47.110 ;
        RECT 33.390 46.730 33.770 46.740 ;
        RECT 36.865 46.730 37.195 46.745 ;
        RECT 33.390 46.430 37.195 46.730 ;
        RECT 41.020 46.730 41.320 47.095 ;
        RECT 69.065 46.730 69.395 46.745 ;
        RECT 41.020 46.430 69.395 46.730 ;
        RECT 33.390 46.420 33.770 46.430 ;
        RECT 36.865 46.415 37.195 46.430 ;
        RECT 69.065 46.415 69.395 46.430 ;
        RECT 21.050 46.075 22.630 46.405 ;
        RECT 34.310 46.050 34.690 46.060 ;
        RECT 65.845 46.050 66.175 46.065 ;
        RECT 67.685 46.050 68.015 46.065 ;
        RECT 34.310 45.750 62.250 46.050 ;
        RECT 34.310 45.740 34.690 45.750 ;
        RECT 28.125 45.370 28.455 45.385 ;
        RECT 31.805 45.370 32.135 45.385 ;
        RECT 41.005 45.370 41.335 45.385 ;
        RECT 28.125 45.070 41.335 45.370 ;
        RECT 28.125 45.055 28.455 45.070 ;
        RECT 31.805 45.055 32.135 45.070 ;
        RECT 41.005 45.055 41.335 45.070 ;
        RECT 48.825 45.370 49.155 45.385 ;
        RECT 60.070 45.370 60.450 45.380 ;
        RECT 48.825 45.070 60.450 45.370 ;
        RECT 61.950 45.370 62.250 45.750 ;
        RECT 65.845 45.750 68.015 46.050 ;
        RECT 65.845 45.735 66.175 45.750 ;
        RECT 67.685 45.735 68.015 45.750 ;
        RECT 74.585 45.370 74.915 45.385 ;
        RECT 61.950 45.070 74.915 45.370 ;
        RECT 48.825 45.055 49.155 45.070 ;
        RECT 60.070 45.060 60.450 45.070 ;
        RECT 74.585 45.055 74.915 45.070 ;
        RECT 39.165 44.690 39.495 44.705 ;
        RECT 47.445 44.690 47.775 44.705 ;
        RECT 39.165 44.390 47.775 44.690 ;
        RECT 39.165 44.375 39.495 44.390 ;
        RECT 47.445 44.375 47.775 44.390 ;
        RECT 52.965 44.690 53.295 44.705 ;
        RECT 61.245 44.690 61.575 44.705 ;
        RECT 52.965 44.390 61.575 44.690 ;
        RECT 52.965 44.375 53.295 44.390 ;
        RECT 61.245 44.375 61.575 44.390 ;
        RECT 65.385 44.690 65.715 44.705 ;
        RECT 65.385 44.390 81.850 44.690 ;
        RECT 65.385 44.375 65.715 44.390 ;
        RECT 46.065 44.010 46.395 44.025 ;
        RECT 65.845 44.010 66.175 44.025 ;
        RECT 46.065 43.710 66.175 44.010 ;
        RECT 46.065 43.695 46.395 43.710 ;
        RECT 65.845 43.695 66.175 43.710 ;
        RECT 24.350 43.355 25.930 43.685 ;
        RECT 36.405 43.330 36.735 43.345 ;
        RECT 72.745 43.330 73.075 43.345 ;
        RECT 76.425 43.330 76.755 43.345 ;
        RECT 36.405 43.030 76.755 43.330 ;
        RECT 36.405 43.015 36.735 43.030 ;
        RECT 72.745 43.015 73.075 43.030 ;
        RECT 76.425 43.015 76.755 43.030 ;
        RECT 2.825 42.650 3.155 42.665 ;
        RECT 51.585 42.650 51.915 42.665 ;
        RECT 2.825 42.350 51.915 42.650 ;
        RECT 2.825 42.335 3.155 42.350 ;
        RECT 51.585 42.335 51.915 42.350 ;
        RECT 53.425 42.650 53.755 42.665 ;
        RECT 59.405 42.650 59.735 42.665 ;
        RECT 53.425 42.350 59.735 42.650 ;
        RECT 53.425 42.335 53.755 42.350 ;
        RECT 59.405 42.335 59.735 42.350 ;
        RECT 30.885 41.970 31.215 41.985 ;
        RECT 39.165 41.970 39.495 41.985 ;
        RECT 30.885 41.670 39.495 41.970 ;
        RECT 30.885 41.655 31.215 41.670 ;
        RECT 39.165 41.655 39.495 41.670 ;
        RECT 43.765 41.970 44.095 41.985 ;
        RECT 48.110 41.970 48.490 41.980 ;
        RECT 43.765 41.670 48.490 41.970 ;
        RECT 43.765 41.655 44.095 41.670 ;
        RECT 48.110 41.660 48.490 41.670 ;
        RECT 51.585 41.970 51.915 41.985 ;
        RECT 57.105 41.970 57.435 41.985 ;
        RECT 51.585 41.670 57.435 41.970 ;
        RECT 51.585 41.655 51.915 41.670 ;
        RECT 57.105 41.655 57.435 41.670 ;
        RECT 58.485 41.970 58.815 41.985 ;
        RECT 68.605 41.970 68.935 41.985 ;
        RECT 58.485 41.670 68.935 41.970 ;
        RECT 58.485 41.655 58.815 41.670 ;
        RECT 68.605 41.655 68.935 41.670 ;
        RECT 57.565 41.290 57.895 41.305 ;
        RECT 57.565 40.990 81.850 41.290 ;
        RECT 57.565 40.975 57.895 40.990 ;
        RECT 21.050 40.635 22.630 40.965 ;
        RECT 27.205 40.610 27.535 40.625 ;
        RECT 27.205 40.310 59.490 40.610 ;
        RECT 27.205 40.295 27.535 40.310 ;
        RECT 58.025 39.940 58.355 39.945 ;
        RECT 58.025 39.930 58.610 39.940 ;
        RECT 57.800 39.630 58.610 39.930 ;
        RECT 59.190 39.930 59.490 40.310 ;
        RECT 64.005 39.930 64.335 39.945 ;
        RECT 59.190 39.630 64.335 39.930 ;
        RECT 58.025 39.620 58.610 39.630 ;
        RECT 58.025 39.615 58.355 39.620 ;
        RECT 64.005 39.615 64.335 39.630 ;
        RECT 53.885 38.570 54.215 38.585 ;
        RECT 58.945 38.570 59.275 38.585 ;
        RECT 66.765 38.570 67.095 38.585 ;
        RECT 53.885 38.270 67.095 38.570 ;
        RECT 53.885 38.255 54.215 38.270 ;
        RECT 58.945 38.255 59.275 38.270 ;
        RECT 66.765 38.255 67.095 38.270 ;
        RECT 24.350 37.915 25.930 38.245 ;
        RECT 55.725 37.890 56.055 37.905 ;
        RECT 58.945 37.890 59.275 37.905 ;
        RECT 55.725 37.590 59.275 37.890 ;
        RECT 55.725 37.575 56.055 37.590 ;
        RECT 58.945 37.575 59.275 37.590 ;
        RECT 68.605 37.890 68.935 37.905 ;
        RECT 68.605 37.590 81.850 37.890 ;
        RECT 68.605 37.575 68.935 37.590 ;
        RECT 53.885 37.210 54.215 37.225 ;
        RECT 68.350 37.210 68.730 37.220 ;
        RECT 53.885 36.910 68.730 37.210 ;
        RECT 53.885 36.895 54.215 36.910 ;
        RECT 68.350 36.900 68.730 36.910 ;
        RECT 56.185 36.530 56.515 36.545 ;
        RECT 58.025 36.530 58.355 36.545 ;
        RECT 56.185 36.230 58.355 36.530 ;
        RECT 56.185 36.215 56.515 36.230 ;
        RECT 58.025 36.215 58.355 36.230 ;
        RECT 59.865 36.530 60.195 36.545 ;
        RECT 60.990 36.530 61.370 36.540 ;
        RECT 69.525 36.530 69.855 36.545 ;
        RECT 59.865 36.230 61.370 36.530 ;
        RECT 59.865 36.215 60.195 36.230 ;
        RECT 60.990 36.220 61.370 36.230 ;
        RECT 61.950 36.230 69.855 36.530 ;
        RECT 51.585 35.850 51.915 35.865 ;
        RECT 61.950 35.850 62.250 36.230 ;
        RECT 69.525 36.215 69.855 36.230 ;
        RECT 51.585 35.550 62.250 35.850 ;
        RECT 51.585 35.535 51.915 35.550 ;
        RECT 21.050 35.195 22.630 35.525 ;
        RECT 59.405 35.170 59.735 35.185 ;
        RECT 61.245 35.170 61.575 35.185 ;
        RECT 59.405 34.870 61.575 35.170 ;
        RECT 59.405 34.855 59.735 34.870 ;
        RECT 61.245 34.855 61.575 34.870 ;
        RECT 52.965 34.490 53.295 34.505 ;
        RECT 62.625 34.490 62.955 34.505 ;
        RECT 52.965 34.190 62.955 34.490 ;
        RECT 52.965 34.175 53.295 34.190 ;
        RECT 62.625 34.175 62.955 34.190 ;
        RECT 71.365 34.490 71.695 34.505 ;
        RECT 71.365 34.190 81.850 34.490 ;
        RECT 71.365 34.175 71.695 34.190 ;
        RECT 44.225 33.810 44.555 33.825 ;
        RECT 71.825 33.810 72.155 33.825 ;
        RECT 44.225 33.510 72.155 33.810 ;
        RECT 44.225 33.495 44.555 33.510 ;
        RECT 71.825 33.495 72.155 33.510 ;
        RECT 24.350 32.475 25.930 32.805 ;
        RECT 58.485 32.450 58.815 32.465 ;
        RECT 67.225 32.450 67.555 32.465 ;
        RECT 58.485 32.150 67.555 32.450 ;
        RECT 58.485 32.135 58.815 32.150 ;
        RECT 67.225 32.135 67.555 32.150 ;
        RECT 25.365 31.770 25.695 31.785 ;
        RECT 32.265 31.770 32.595 31.785 ;
        RECT 39.625 31.770 39.955 31.785 ;
        RECT 25.365 31.470 39.955 31.770 ;
        RECT 25.365 31.455 25.695 31.470 ;
        RECT 32.265 31.455 32.595 31.470 ;
        RECT 39.625 31.455 39.955 31.470 ;
        RECT 52.045 31.770 52.375 31.785 ;
        RECT 69.065 31.770 69.395 31.785 ;
        RECT 52.045 31.470 69.395 31.770 ;
        RECT 52.045 31.455 52.375 31.470 ;
        RECT 69.065 31.455 69.395 31.470 ;
        RECT 3.745 31.090 4.075 31.105 ;
        RECT 0.500 30.790 4.075 31.090 ;
        RECT 3.745 30.775 4.075 30.790 ;
        RECT 33.185 31.090 33.515 31.105 ;
        RECT 41.005 31.090 41.335 31.105 ;
        RECT 33.185 30.790 41.335 31.090 ;
        RECT 33.185 30.775 33.515 30.790 ;
        RECT 41.005 30.775 41.335 30.790 ;
        RECT 54.345 31.090 54.675 31.105 ;
        RECT 56.645 31.090 56.975 31.105 ;
        RECT 62.165 31.090 62.495 31.105 ;
        RECT 54.345 30.790 62.495 31.090 ;
        RECT 54.345 30.775 54.675 30.790 ;
        RECT 56.645 30.775 56.975 30.790 ;
        RECT 62.165 30.775 62.495 30.790 ;
        RECT 70.905 31.090 71.235 31.105 ;
        RECT 70.905 30.790 81.850 31.090 ;
        RECT 70.905 30.775 71.235 30.790 ;
        RECT 21.050 29.755 22.630 30.085 ;
        RECT 37.325 29.050 37.655 29.065 ;
        RECT 38.245 29.050 38.575 29.065 ;
        RECT 37.325 28.750 38.575 29.050 ;
        RECT 37.325 28.735 37.655 28.750 ;
        RECT 38.245 28.735 38.575 28.750 ;
        RECT 35.025 28.370 35.355 28.385 ;
        RECT 39.625 28.370 39.955 28.385 ;
        RECT 35.025 28.070 39.955 28.370 ;
        RECT 35.025 28.055 35.355 28.070 ;
        RECT 39.625 28.055 39.955 28.070 ;
        RECT 4.665 27.690 4.995 27.705 ;
        RECT 0.500 27.390 4.995 27.690 ;
        RECT 4.665 27.375 4.995 27.390 ;
        RECT 35.485 27.690 35.815 27.705 ;
        RECT 41.005 27.690 41.335 27.705 ;
        RECT 35.485 27.390 41.335 27.690 ;
        RECT 35.485 27.375 35.815 27.390 ;
        RECT 41.005 27.375 41.335 27.390 ;
        RECT 75.045 27.690 75.375 27.705 ;
        RECT 75.045 27.390 81.850 27.690 ;
        RECT 75.045 27.375 75.375 27.390 ;
        RECT 24.350 27.035 25.930 27.365 ;
        RECT 30.885 27.010 31.215 27.025 ;
        RECT 39.625 27.010 39.955 27.025 ;
        RECT 30.885 26.710 39.955 27.010 ;
        RECT 30.885 26.695 31.215 26.710 ;
        RECT 39.625 26.695 39.955 26.710 ;
        RECT 31.345 26.330 31.675 26.345 ;
        RECT 35.485 26.330 35.815 26.345 ;
        RECT 31.345 26.030 35.815 26.330 ;
        RECT 31.345 26.015 31.675 26.030 ;
        RECT 35.485 26.015 35.815 26.030 ;
        RECT 50.205 24.970 50.535 24.985 ;
        RECT 58.485 24.970 58.815 24.985 ;
        RECT 50.205 24.670 58.815 24.970 ;
        RECT 50.205 24.655 50.535 24.670 ;
        RECT 58.485 24.655 58.815 24.670 ;
        RECT 21.050 24.315 22.630 24.645 ;
        RECT 3.745 24.290 4.075 24.305 ;
        RECT 0.500 23.990 4.075 24.290 ;
        RECT 3.745 23.975 4.075 23.990 ;
        RECT 48.825 24.290 49.155 24.305 ;
        RECT 51.125 24.290 51.455 24.305 ;
        RECT 48.825 23.990 51.455 24.290 ;
        RECT 48.825 23.975 49.155 23.990 ;
        RECT 51.125 23.975 51.455 23.990 ;
        RECT 67.685 24.290 68.015 24.305 ;
        RECT 67.685 23.990 81.850 24.290 ;
        RECT 67.685 23.975 68.015 23.990 ;
        RECT 48.365 23.610 48.695 23.625 ;
        RECT 52.045 23.610 52.375 23.625 ;
        RECT 72.285 23.610 72.615 23.625 ;
        RECT 48.365 23.310 72.615 23.610 ;
        RECT 48.365 23.295 48.695 23.310 ;
        RECT 52.045 23.295 52.375 23.310 ;
        RECT 72.285 23.295 72.615 23.310 ;
        RECT 24.350 21.595 25.930 21.925 ;
        RECT 1.905 20.890 2.235 20.905 ;
        RECT 0.500 20.590 2.235 20.890 ;
        RECT 1.905 20.575 2.235 20.590 ;
        RECT 48.825 20.890 49.155 20.905 ;
        RECT 51.585 20.890 51.915 20.905 ;
        RECT 48.825 20.590 51.915 20.890 ;
        RECT 48.825 20.575 49.155 20.590 ;
        RECT 51.585 20.575 51.915 20.590 ;
        RECT 73.665 20.890 73.995 20.905 ;
        RECT 73.665 20.590 81.850 20.890 ;
        RECT 73.665 20.575 73.995 20.590 ;
        RECT 21.050 18.875 22.630 19.205 ;
        RECT 48.365 18.850 48.695 18.865 ;
        RECT 52.045 18.850 52.375 18.865 ;
        RECT 48.365 18.550 52.375 18.850 ;
        RECT 48.365 18.535 48.695 18.550 ;
        RECT 52.045 18.535 52.375 18.550 ;
        RECT 74.585 17.490 74.915 17.505 ;
        RECT 74.585 17.190 81.850 17.490 ;
        RECT 74.585 17.175 74.915 17.190 ;
        RECT 24.350 16.155 25.930 16.485 ;
        RECT 75.045 14.090 75.375 14.105 ;
        RECT 75.045 13.790 81.850 14.090 ;
        RECT 75.045 13.775 75.375 13.790 ;
        RECT 21.050 13.435 22.630 13.765 ;
        RECT 24.350 10.715 25.930 11.045 ;
      LAYER met4 ;
        RECT 33.415 90.615 33.745 90.945 ;
        RECT 30.655 85.175 30.985 85.505 ;
        RECT 28.815 84.495 29.145 84.825 ;
        RECT 13.175 83.135 13.505 83.465 ;
        RECT 27.895 83.135 28.225 83.465 ;
        RECT 12.255 70.895 12.585 71.225 ;
        RECT 11.335 70.215 11.665 70.545 ;
        RECT 11.350 54.225 11.650 70.215 ;
        RECT 11.335 53.895 11.665 54.225 ;
        RECT 12.270 47.425 12.570 70.895 ;
        RECT 13.190 66.450 13.490 83.135 ;
        RECT 26.975 81.095 27.305 81.425 ;
        RECT 18.695 77.695 19.025 78.025 ;
        RECT 17.775 76.335 18.105 76.665 ;
        RECT 16.855 68.855 17.185 69.185 ;
        RECT 13.190 66.150 14.410 66.450 ;
        RECT 14.110 54.905 14.410 66.150 ;
        RECT 15.015 61.375 15.345 61.705 ;
        RECT 15.030 58.305 15.330 61.375 ;
        RECT 15.935 60.015 16.265 60.345 ;
        RECT 15.015 57.975 15.345 58.305 ;
        RECT 14.095 54.575 14.425 54.905 ;
        RECT 15.950 51.505 16.250 60.015 ;
        RECT 15.935 51.175 16.265 51.505 ;
        RECT 16.870 50.145 17.170 68.855 ;
        RECT 17.790 58.305 18.090 76.335 ;
        RECT 17.775 57.975 18.105 58.305 ;
        RECT 18.710 56.945 19.010 77.695 ;
        RECT 23.295 76.335 23.625 76.665 ;
        RECT 19.615 67.495 19.945 67.825 ;
        RECT 18.695 56.615 19.025 56.945 ;
        RECT 19.630 54.225 19.930 67.495 ;
        RECT 19.615 53.895 19.945 54.225 ;
        RECT 16.855 49.815 17.185 50.145 ;
        RECT 23.310 48.785 23.610 76.335 ;
        RECT 26.990 63.745 27.290 81.095 ;
        RECT 26.975 63.415 27.305 63.745 ;
        RECT 27.910 63.050 28.210 83.135 ;
        RECT 26.300 62.750 28.210 63.050 ;
        RECT 26.300 59.650 26.600 62.750 ;
        RECT 27.895 61.375 28.225 61.705 ;
        RECT 26.300 59.350 27.290 59.650 ;
        RECT 26.990 56.945 27.290 59.350 ;
        RECT 26.975 56.615 27.305 56.945 ;
        RECT 27.910 52.185 28.210 61.375 ;
        RECT 28.830 57.625 29.130 84.495 ;
        RECT 29.735 68.855 30.065 69.185 ;
        RECT 29.750 57.625 30.050 68.855 ;
        RECT 30.670 67.145 30.970 85.175 ;
        RECT 31.575 77.695 31.905 78.025 ;
        RECT 30.655 66.815 30.985 67.145 ;
        RECT 30.655 63.415 30.985 63.745 ;
        RECT 28.815 57.295 29.145 57.625 ;
        RECT 29.735 57.295 30.065 57.625 ;
        RECT 27.895 51.855 28.225 52.185 ;
        RECT 23.295 48.455 23.625 48.785 ;
        RECT 30.670 47.425 30.970 63.415 ;
        RECT 31.590 59.665 31.890 77.695 ;
        RECT 32.495 76.335 32.825 76.665 ;
        RECT 31.575 59.335 31.905 59.665 ;
        RECT 32.510 48.105 32.810 76.335 ;
        RECT 33.430 60.345 33.730 90.615 ;
        RECT 40.775 89.255 41.105 89.585 ;
        RECT 39.855 88.575 40.185 88.905 ;
        RECT 35.255 76.335 35.585 76.665 ;
        RECT 33.415 60.015 33.745 60.345 ;
        RECT 33.415 57.295 33.745 57.625 ;
        RECT 32.495 47.775 32.825 48.105 ;
        RECT 12.255 47.095 12.585 47.425 ;
        RECT 30.655 47.095 30.985 47.425 ;
        RECT 33.430 46.745 33.730 57.295 ;
        RECT 34.335 56.615 34.665 56.945 ;
        RECT 33.415 46.415 33.745 46.745 ;
        RECT 34.350 46.065 34.650 56.615 ;
        RECT 35.270 54.905 35.570 76.335 ;
        RECT 36.175 70.895 36.505 71.225 ;
        RECT 35.255 54.575 35.585 54.905 ;
        RECT 36.190 48.105 36.490 70.895 ;
        RECT 39.870 54.905 40.170 88.575 ;
        RECT 40.790 75.985 41.090 89.255 ;
        RECT 68.375 87.895 68.705 88.225 ;
        RECT 44.455 87.215 44.785 87.545 ;
        RECT 40.775 75.655 41.105 75.985 ;
        RECT 40.775 71.575 41.105 71.905 ;
        RECT 39.855 54.575 40.185 54.905 ;
        RECT 40.790 48.105 41.090 71.575 ;
        RECT 44.470 48.105 44.770 87.215 ;
        RECT 45.375 86.535 45.705 86.865 ;
        RECT 45.390 48.105 45.690 86.535 ;
        RECT 60.095 83.135 60.425 83.465 ;
        RECT 58.255 78.375 58.585 78.705 ;
        RECT 46.295 74.295 46.625 74.625 ;
        RECT 46.310 69.185 46.610 74.295 ;
        RECT 46.295 68.855 46.625 69.185 ;
        RECT 48.135 66.135 48.465 66.465 ;
        RECT 36.175 47.775 36.505 48.105 ;
        RECT 40.775 47.775 41.105 48.105 ;
        RECT 44.455 47.775 44.785 48.105 ;
        RECT 45.375 47.775 45.705 48.105 ;
        RECT 34.335 45.735 34.665 46.065 ;
        RECT 48.150 41.985 48.450 66.135 ;
        RECT 48.135 41.655 48.465 41.985 ;
        RECT 58.270 39.945 58.570 78.375 ;
        RECT 60.110 45.385 60.410 83.135 ;
        RECT 63.775 78.375 64.105 78.705 ;
        RECT 61.015 76.335 61.345 76.665 ;
        RECT 60.095 45.055 60.425 45.385 ;
        RECT 58.255 39.615 58.585 39.945 ;
        RECT 61.030 36.545 61.330 76.335 ;
        RECT 63.790 48.785 64.090 78.375 ;
        RECT 63.775 48.455 64.105 48.785 ;
        RECT 68.390 37.225 68.690 87.895 ;
        RECT 68.375 36.895 68.705 37.225 ;
        RECT 61.015 36.215 61.345 36.545 ;
  END
END digital
END LIBRARY

