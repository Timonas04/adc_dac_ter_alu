VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 18.245 209.755 18.415 209.945 ;
        RECT 20.545 209.755 20.715 209.945 ;
        RECT 21.005 209.755 21.175 209.945 ;
        RECT 24.225 209.755 24.395 209.945 ;
        RECT 26.065 209.755 26.235 209.945 ;
        RECT 26.525 209.775 26.695 209.945 ;
        RECT 26.530 209.755 26.695 209.775 ;
        RECT 30.660 209.755 30.830 209.945 ;
        RECT 33.420 209.755 33.590 209.945 ;
        RECT 33.885 209.775 34.055 209.945 ;
        RECT 33.915 209.755 34.055 209.775 ;
        RECT 36.645 209.755 36.815 209.945 ;
        RECT 39.840 209.755 40.010 209.945 ;
        RECT 44.475 209.800 44.635 209.910 ;
        RECT 54.125 209.755 54.295 209.945 ;
        RECT 54.590 209.755 54.760 209.945 ;
        RECT 60.100 209.755 60.270 209.945 ;
        RECT 69.305 209.755 69.475 209.945 ;
        RECT 71.605 209.755 71.775 209.945 ;
        RECT 72.065 209.755 72.235 209.945 ;
        RECT 81.265 209.755 81.435 209.945 ;
        RECT 83.105 209.775 83.275 209.945 ;
        RECT 83.105 209.755 83.305 209.775 ;
        RECT 87.695 209.755 87.865 209.945 ;
        RECT 89.085 209.755 89.255 209.945 ;
        RECT 18.105 208.945 19.475 209.755 ;
        RECT 19.495 208.845 20.845 209.755 ;
        RECT 20.865 209.075 22.695 209.755 ;
        RECT 21.350 208.845 22.695 209.075 ;
        RECT 22.705 209.075 24.535 209.755 ;
        RECT 24.545 209.075 26.375 209.755 ;
        RECT 26.530 209.075 28.365 209.755 ;
        RECT 22.705 208.845 24.050 209.075 ;
        RECT 24.545 208.845 25.890 209.075 ;
        RECT 27.435 208.845 28.365 209.075 ;
        RECT 28.785 208.845 30.975 209.755 ;
        RECT 30.995 208.885 31.425 209.670 ;
        RECT 31.545 208.845 33.735 209.755 ;
        RECT 33.915 208.935 36.485 209.755 ;
        RECT 36.505 209.075 39.715 209.755 ;
        RECT 34.895 208.845 36.485 208.935 ;
        RECT 38.580 208.845 39.715 209.075 ;
        RECT 39.780 208.845 43.855 209.755 ;
        RECT 43.875 208.885 44.305 209.670 ;
        RECT 45.330 209.075 54.435 209.755 ;
        RECT 54.445 209.075 56.720 209.755 ;
        RECT 55.350 208.845 56.720 209.075 ;
        RECT 56.755 208.885 57.185 209.670 ;
        RECT 57.495 208.845 60.415 209.755 ;
        RECT 60.510 209.075 69.615 209.755 ;
        RECT 69.635 208.885 70.065 209.670 ;
        RECT 70.085 208.845 71.900 209.755 ;
        RECT 71.925 209.075 81.030 209.755 ;
        RECT 81.135 208.845 82.485 209.755 ;
        RECT 82.515 208.885 82.945 209.670 ;
        RECT 83.105 209.075 86.635 209.755 ;
        RECT 83.810 208.845 86.635 209.075 ;
        RECT 86.645 208.975 88.015 209.755 ;
        RECT 88.025 208.945 89.395 209.755 ;
      LAYER nwell ;
        RECT 17.910 205.725 89.590 208.555 ;
      LAYER pwell ;
        RECT 20.605 205.345 21.555 205.435 ;
        RECT 18.105 204.525 19.475 205.335 ;
        RECT 20.605 204.525 22.535 205.345 ;
        RECT 22.705 205.205 24.050 205.435 ;
        RECT 25.685 205.345 26.635 205.435 ;
        RECT 22.705 204.525 24.535 205.205 ;
        RECT 24.705 204.525 26.635 205.345 ;
        RECT 29.130 205.235 30.515 205.435 ;
        RECT 26.845 204.555 30.515 205.235 ;
        RECT 30.995 204.610 31.425 205.395 ;
        RECT 18.245 204.315 18.415 204.525 ;
        RECT 22.385 204.505 22.535 204.525 ;
        RECT 19.635 204.370 19.795 204.480 ;
        RECT 21.005 204.315 21.175 204.505 ;
        RECT 21.460 204.315 21.630 204.505 ;
        RECT 22.385 204.335 22.555 204.505 ;
        RECT 22.840 204.315 23.010 204.505 ;
        RECT 24.225 204.335 24.395 204.525 ;
        RECT 24.705 204.505 24.855 204.525 ;
        RECT 24.685 204.335 24.855 204.505 ;
        RECT 26.060 204.315 26.230 204.505 ;
        RECT 26.985 204.335 27.155 204.555 ;
        RECT 29.145 204.525 30.515 204.555 ;
        RECT 31.905 204.525 35.575 205.435 ;
        RECT 35.585 205.205 37.175 205.435 ;
        RECT 35.585 204.525 39.255 205.205 ;
        RECT 39.350 204.525 48.455 205.205 ;
        RECT 48.465 204.525 52.565 205.435 ;
        RECT 52.605 204.525 56.275 205.435 ;
        RECT 56.755 204.610 57.185 205.395 ;
        RECT 60.625 205.205 64.555 205.435 ;
        RECT 74.610 205.205 77.435 205.435 ;
        RECT 78.290 205.205 81.115 205.435 ;
        RECT 57.205 204.525 59.945 205.205 ;
        RECT 60.140 204.525 64.555 205.205 ;
        RECT 64.565 204.525 73.670 205.205 ;
        RECT 73.905 204.525 77.435 205.205 ;
        RECT 77.585 204.525 81.115 205.205 ;
        RECT 81.135 204.525 82.485 205.435 ;
        RECT 82.515 204.610 82.945 205.395 ;
        RECT 83.810 205.205 86.635 205.435 ;
        RECT 83.105 204.525 86.635 205.205 ;
        RECT 86.645 204.525 88.015 205.305 ;
        RECT 88.025 204.525 89.395 205.335 ;
        RECT 18.105 203.505 19.475 204.315 ;
        RECT 19.485 203.635 21.315 204.315 ;
        RECT 19.485 203.405 20.830 203.635 ;
        RECT 21.345 203.405 22.695 204.315 ;
        RECT 22.725 203.405 24.075 204.315 ;
        RECT 24.540 204.085 26.230 204.315 ;
        RECT 26.385 204.285 27.780 204.315 ;
        RECT 28.825 204.285 28.995 204.505 ;
        RECT 29.285 204.335 29.455 204.505 ;
        RECT 30.660 204.365 30.780 204.475 ;
        RECT 31.580 204.365 31.700 204.475 ;
        RECT 32.050 204.335 32.220 204.525 ;
        RECT 29.315 204.315 29.455 204.335 ;
        RECT 34.345 204.315 34.515 204.505 ;
        RECT 38.940 204.335 39.110 204.525 ;
        RECT 43.545 204.315 43.715 204.505 ;
        RECT 44.475 204.360 44.635 204.470 ;
        RECT 45.385 204.315 45.555 204.505 ;
        RECT 48.145 204.335 48.315 204.525 ;
        RECT 48.610 204.335 48.780 204.525 ;
        RECT 55.960 204.335 56.130 204.525 ;
        RECT 56.420 204.365 56.540 204.475 ;
        RECT 57.345 204.335 57.515 204.525 ;
        RECT 60.140 204.505 60.250 204.525 ;
        RECT 64.705 204.505 64.875 204.525 ;
        RECT 73.905 204.505 74.105 204.525 ;
        RECT 77.585 204.505 77.785 204.525 ;
        RECT 60.080 204.335 60.250 204.505 ;
        RECT 63.325 204.315 63.495 204.505 ;
        RECT 64.700 204.335 64.875 204.505 ;
        RECT 64.700 204.315 64.870 204.335 ;
        RECT 65.170 204.315 65.340 204.505 ;
        RECT 68.855 204.360 69.015 204.470 ;
        RECT 73.445 204.335 73.615 204.505 ;
        RECT 73.415 204.315 73.615 204.335 ;
        RECT 73.905 204.315 74.075 204.505 ;
        RECT 77.585 204.335 77.755 204.505 ;
        RECT 82.185 204.335 82.355 204.525 ;
        RECT 83.105 204.505 83.305 204.525 ;
        RECT 83.105 204.335 83.275 204.505 ;
        RECT 84.025 204.315 84.195 204.505 ;
        RECT 87.240 204.315 87.410 204.505 ;
        RECT 87.705 204.475 87.875 204.525 ;
        RECT 87.700 204.365 87.875 204.475 ;
        RECT 87.705 204.335 87.875 204.365 ;
        RECT 89.085 204.315 89.255 204.525 ;
        RECT 24.540 203.405 26.375 204.085 ;
        RECT 26.385 203.605 29.120 204.285 ;
        RECT 26.385 203.405 27.795 203.605 ;
        RECT 29.315 203.495 31.885 204.315 ;
        RECT 31.915 203.635 34.655 204.315 ;
        RECT 34.750 203.635 43.855 204.315 ;
        RECT 30.295 203.405 31.885 203.495 ;
        RECT 43.875 203.445 44.305 204.230 ;
        RECT 45.245 203.635 54.350 204.315 ;
        RECT 54.530 203.635 63.635 204.315 ;
        RECT 63.665 203.405 65.015 204.315 ;
        RECT 65.025 203.405 68.625 204.315 ;
        RECT 69.635 203.445 70.065 204.230 ;
        RECT 70.085 203.635 73.615 204.315 ;
        RECT 70.085 203.405 72.910 203.635 ;
        RECT 73.775 203.405 75.125 204.315 ;
        RECT 75.230 203.635 84.335 204.315 ;
        RECT 84.345 203.405 87.555 204.315 ;
        RECT 88.025 203.505 89.395 204.315 ;
      LAYER nwell ;
        RECT 17.910 200.285 89.590 203.115 ;
      LAYER pwell ;
        RECT 18.105 199.085 19.475 199.895 ;
        RECT 20.890 199.765 22.235 199.995 ;
        RECT 20.405 199.085 22.235 199.765 ;
        RECT 22.245 199.765 23.590 199.995 ;
        RECT 22.245 199.085 24.075 199.765 ;
        RECT 25.025 199.085 26.375 199.995 ;
        RECT 27.525 199.905 28.475 199.995 ;
        RECT 26.545 199.085 28.475 199.905 ;
        RECT 28.685 199.085 30.975 199.995 ;
        RECT 30.995 199.170 31.425 199.955 ;
        RECT 31.445 199.085 32.815 199.865 ;
        RECT 32.835 199.085 35.565 199.995 ;
        RECT 35.585 199.085 38.325 199.765 ;
        RECT 38.430 199.085 47.535 199.765 ;
        RECT 47.630 199.085 56.735 199.765 ;
        RECT 56.755 199.170 57.185 199.955 ;
        RECT 57.205 199.085 61.335 199.995 ;
        RECT 61.365 199.085 62.715 199.995 ;
        RECT 62.725 199.085 71.830 199.765 ;
        RECT 71.925 199.085 81.030 199.765 ;
        RECT 81.125 199.085 82.495 199.865 ;
        RECT 82.515 199.170 82.945 199.955 ;
        RECT 82.975 199.315 86.175 199.995 ;
        RECT 86.670 199.765 88.015 199.995 ;
        RECT 82.975 199.085 86.030 199.315 ;
        RECT 86.185 199.085 88.015 199.765 ;
        RECT 88.025 199.085 89.395 199.895 ;
        RECT 18.245 198.875 18.415 199.085 ;
        RECT 19.635 198.930 19.795 199.040 ;
        RECT 20.545 198.895 20.715 199.085 ;
        RECT 21.005 198.875 21.175 199.065 ;
        RECT 21.460 198.925 21.580 199.035 ;
        RECT 22.385 198.915 22.555 199.065 ;
        RECT 18.105 198.065 19.475 198.875 ;
        RECT 19.485 198.195 21.315 198.875 ;
        RECT 19.485 197.965 20.830 198.195 ;
        RECT 21.785 197.965 22.675 198.915 ;
        RECT 22.855 198.875 23.025 199.065 ;
        RECT 23.765 198.895 23.935 199.085 ;
        RECT 24.230 198.875 24.400 199.065 ;
        RECT 25.140 198.895 25.310 199.085 ;
        RECT 26.545 199.065 26.695 199.085 ;
        RECT 26.525 198.895 26.695 199.065 ;
        RECT 27.905 198.875 28.075 199.065 ;
        RECT 30.660 198.895 30.830 199.085 ;
        RECT 32.505 198.895 32.675 199.085 ;
        RECT 32.505 198.875 32.670 198.895 ;
        RECT 32.965 198.875 33.135 199.065 ;
        RECT 35.265 198.895 35.435 199.085 ;
        RECT 35.725 198.895 35.895 199.085 ;
        RECT 38.945 198.875 39.115 199.065 ;
        RECT 40.330 198.875 40.500 199.065 ;
        RECT 40.790 198.875 40.960 199.065 ;
        RECT 22.705 198.095 24.075 198.875 ;
        RECT 24.085 197.965 27.755 198.875 ;
        RECT 27.765 197.965 30.515 198.875 ;
        RECT 30.835 198.195 32.670 198.875 ;
        RECT 30.835 197.965 31.765 198.195 ;
        RECT 32.825 197.965 36.035 198.875 ;
        RECT 36.045 197.965 39.255 198.875 ;
        RECT 39.265 197.965 40.615 198.875 ;
        RECT 40.645 197.965 43.565 198.875 ;
        RECT 43.875 198.005 44.305 198.790 ;
        RECT 44.470 198.645 44.640 199.065 ;
        RECT 47.225 198.895 47.395 199.085 ;
        RECT 49.070 198.875 49.240 199.065 ;
        RECT 52.745 198.875 52.915 199.065 ;
        RECT 56.425 198.895 56.595 199.085 ;
        RECT 61.020 198.895 61.190 199.085 ;
        RECT 62.400 198.895 62.570 199.085 ;
        RECT 62.865 198.895 63.035 199.085 ;
        RECT 65.620 198.875 65.790 199.065 ;
        RECT 66.090 198.895 66.260 199.065 ;
        RECT 69.300 198.925 69.420 199.035 ;
        RECT 66.115 198.875 66.260 198.895 ;
        RECT 70.225 198.875 70.395 199.065 ;
        RECT 72.065 198.895 72.235 199.085 ;
        RECT 79.430 198.875 79.600 199.065 ;
        RECT 81.265 198.895 81.435 199.085 ;
        RECT 83.110 198.875 83.280 199.065 ;
        RECT 85.860 198.895 86.030 199.085 ;
        RECT 86.325 198.895 86.495 199.085 ;
        RECT 87.695 198.875 87.865 199.065 ;
        RECT 89.085 198.875 89.255 199.085 ;
        RECT 45.750 198.645 48.910 198.875 ;
        RECT 44.365 198.195 48.910 198.645 ;
        RECT 44.365 197.965 45.740 198.195 ;
        RECT 47.530 197.965 48.910 198.195 ;
        RECT 48.925 197.965 52.580 198.875 ;
        RECT 52.605 198.195 61.710 198.875 ;
        RECT 61.805 197.965 65.935 198.875 ;
        RECT 66.115 197.965 69.155 198.875 ;
        RECT 69.635 198.005 70.065 198.790 ;
        RECT 70.085 198.195 79.190 198.875 ;
        RECT 79.285 197.965 82.830 198.875 ;
        RECT 82.965 197.965 86.510 198.875 ;
        RECT 86.645 198.095 88.015 198.875 ;
        RECT 88.025 198.065 89.395 198.875 ;
      LAYER nwell ;
        RECT 17.910 194.845 89.590 197.675 ;
      LAYER pwell ;
        RECT 19.955 194.465 21.545 194.555 ;
        RECT 18.105 193.645 19.475 194.455 ;
        RECT 19.955 193.645 22.525 194.465 ;
        RECT 23.755 194.325 24.685 194.555 ;
        RECT 18.245 193.435 18.415 193.645 ;
        RECT 22.385 193.625 22.525 193.645 ;
        RECT 22.850 193.645 24.685 194.325 ;
        RECT 25.005 193.645 28.675 194.555 ;
        RECT 29.605 193.645 30.975 194.425 ;
        RECT 30.995 193.730 31.425 194.515 ;
        RECT 31.445 193.645 32.795 194.555 ;
        RECT 32.825 193.645 34.655 194.555 ;
        RECT 34.815 193.645 38.470 194.555 ;
        RECT 39.265 193.645 42.475 194.555 ;
        RECT 42.570 193.645 51.675 194.325 ;
        RECT 51.685 193.645 55.815 194.555 ;
        RECT 56.755 193.730 57.185 194.515 ;
        RECT 57.290 193.645 66.395 194.325 ;
        RECT 66.405 193.645 69.615 194.555 ;
        RECT 69.625 193.645 73.295 194.555 ;
        RECT 73.390 193.645 82.495 194.325 ;
        RECT 82.515 193.730 82.945 194.515 ;
        RECT 83.810 194.325 86.635 194.555 ;
        RECT 83.105 193.645 86.635 194.325 ;
        RECT 86.655 193.645 88.005 194.555 ;
        RECT 88.025 193.645 89.395 194.455 ;
        RECT 22.850 193.625 23.015 193.645 ;
        RECT 19.620 193.485 19.740 193.595 ;
        RECT 21.005 193.435 21.175 193.625 ;
        RECT 21.475 193.435 21.645 193.625 ;
        RECT 22.385 193.455 22.555 193.625 ;
        RECT 22.845 193.455 23.015 193.625 ;
        RECT 23.765 193.435 23.935 193.625 ;
        RECT 25.145 193.435 25.315 193.625 ;
        RECT 25.600 193.485 25.720 193.595 ;
        RECT 26.065 193.435 26.235 193.625 ;
        RECT 28.360 193.455 28.530 193.645 ;
        RECT 28.835 193.490 28.995 193.600 ;
        RECT 30.665 193.455 30.835 193.645 ;
        RECT 31.120 193.485 31.240 193.595 ;
        RECT 30.665 193.435 30.830 193.455 ;
        RECT 31.595 193.435 31.765 193.625 ;
        RECT 32.510 193.455 32.680 193.645 ;
        RECT 32.970 193.455 33.140 193.645 ;
        RECT 34.815 193.625 34.975 193.645 ;
        RECT 34.345 193.435 34.515 193.625 ;
        RECT 34.805 193.455 34.975 193.625 ;
        RECT 37.565 193.455 37.735 193.625 ;
        RECT 37.565 193.435 37.715 193.455 ;
        RECT 38.025 193.435 38.195 193.625 ;
        RECT 38.940 193.485 39.060 193.595 ;
        RECT 39.405 193.455 39.575 193.645 ;
        RECT 43.540 193.435 43.710 193.625 ;
        RECT 47.225 193.435 47.395 193.625 ;
        RECT 47.685 193.435 47.855 193.625 ;
        RECT 51.365 193.455 51.535 193.645 ;
        RECT 51.830 193.455 52.000 193.645 ;
        RECT 55.975 193.490 56.135 193.600 ;
        RECT 59.645 193.435 59.815 193.625 ;
        RECT 60.100 193.485 60.220 193.595 ;
        RECT 66.085 193.455 66.255 193.645 ;
        RECT 69.300 193.625 69.470 193.645 ;
        RECT 69.300 193.455 69.475 193.625 ;
        RECT 69.770 193.455 69.940 193.645 ;
        RECT 69.305 193.435 69.475 193.455 ;
        RECT 70.225 193.435 70.395 193.625 ;
        RECT 73.440 193.485 73.560 193.595 ;
        RECT 73.910 193.435 74.080 193.625 ;
        RECT 78.055 193.480 78.215 193.590 ;
        RECT 82.185 193.455 82.355 193.645 ;
        RECT 83.105 193.625 83.305 193.645 ;
        RECT 83.105 193.455 83.275 193.625 ;
        RECT 86.785 193.455 86.955 193.645 ;
        RECT 87.705 193.435 87.875 193.625 ;
        RECT 89.085 193.435 89.255 193.645 ;
        RECT 18.105 192.625 19.475 193.435 ;
        RECT 19.485 192.755 21.315 193.435 ;
        RECT 19.485 192.525 20.830 192.755 ;
        RECT 21.325 192.655 22.695 193.435 ;
        RECT 22.705 192.655 24.075 193.435 ;
        RECT 24.095 192.525 25.445 193.435 ;
        RECT 25.935 192.525 28.665 193.435 ;
        RECT 28.995 192.755 30.830 193.435 ;
        RECT 28.995 192.525 29.925 192.755 ;
        RECT 31.445 192.655 32.815 193.435 ;
        RECT 32.825 192.525 34.640 193.435 ;
        RECT 35.785 192.615 37.715 193.435 ;
        RECT 37.885 192.755 40.635 193.435 ;
        RECT 35.785 192.525 36.735 192.615 ;
        RECT 39.705 192.525 40.635 192.755 ;
        RECT 40.645 192.525 43.855 193.435 ;
        RECT 43.875 192.565 44.305 193.350 ;
        RECT 44.325 192.525 47.535 193.435 ;
        RECT 47.545 192.525 50.755 193.435 ;
        RECT 50.850 192.755 59.955 193.435 ;
        RECT 60.510 192.755 69.615 193.435 ;
        RECT 70.085 193.405 71.925 193.435 ;
        RECT 69.635 192.565 70.065 193.350 ;
        RECT 70.085 192.755 73.250 193.405 ;
        RECT 70.570 192.725 73.250 192.755 ;
        RECT 70.570 192.525 71.925 192.725 ;
        RECT 73.765 192.525 77.895 193.435 ;
        RECT 78.910 192.755 88.015 193.435 ;
        RECT 88.025 192.625 89.395 193.435 ;
      LAYER nwell ;
        RECT 17.910 189.405 89.590 192.235 ;
      LAYER pwell ;
        RECT 18.105 188.205 19.475 189.015 ;
        RECT 20.405 188.205 21.775 188.985 ;
        RECT 21.785 188.205 23.155 188.985 ;
        RECT 23.165 188.205 24.535 188.985 ;
        RECT 26.975 188.885 27.905 189.115 ;
        RECT 26.070 188.205 27.905 188.885 ;
        RECT 28.225 188.885 29.570 189.115 ;
        RECT 28.225 188.205 30.055 188.885 ;
        RECT 30.995 188.290 31.425 189.075 ;
        RECT 32.365 188.885 33.295 189.115 ;
        RECT 32.365 188.205 36.265 188.885 ;
        RECT 36.965 188.205 38.335 188.985 ;
        RECT 38.345 188.205 40.160 189.115 ;
        RECT 40.270 188.205 49.375 188.885 ;
        RECT 49.385 188.205 53.040 189.115 ;
        RECT 53.065 188.205 56.735 189.115 ;
        RECT 56.755 188.290 57.185 189.075 ;
        RECT 57.215 188.205 59.955 188.885 ;
        RECT 59.965 188.205 64.040 189.115 ;
        RECT 64.105 188.205 73.210 188.885 ;
        RECT 73.390 188.205 82.495 188.885 ;
        RECT 82.515 188.290 82.945 189.075 ;
        RECT 82.965 188.205 86.005 189.115 ;
        RECT 86.185 188.205 88.015 189.115 ;
        RECT 88.025 188.205 89.395 189.015 ;
        RECT 18.245 187.995 18.415 188.205 ;
        RECT 21.465 188.185 21.635 188.205 ;
        RECT 19.635 188.050 19.795 188.160 ;
        RECT 21.005 187.995 21.175 188.185 ;
        RECT 21.460 188.015 21.635 188.185 ;
        RECT 22.845 188.015 23.015 188.205 ;
        RECT 24.225 188.015 24.395 188.205 ;
        RECT 26.070 188.185 26.235 188.205 ;
        RECT 24.685 188.015 24.855 188.185 ;
        RECT 21.460 187.995 21.630 188.015 ;
        RECT 25.605 187.995 25.775 188.185 ;
        RECT 26.065 188.015 26.235 188.185 ;
        RECT 26.990 187.995 27.160 188.185 ;
        RECT 29.745 188.015 29.915 188.205 ;
        RECT 30.215 188.050 30.375 188.160 ;
        RECT 30.670 187.995 30.840 188.185 ;
        RECT 31.595 188.050 31.755 188.160 ;
        RECT 32.045 187.995 32.215 188.185 ;
        RECT 32.780 188.015 32.950 188.205 ;
        RECT 33.700 187.995 33.870 188.185 ;
        RECT 36.640 188.045 36.760 188.155 ;
        RECT 37.105 188.015 37.275 188.205 ;
        RECT 37.840 187.995 38.010 188.185 ;
        RECT 39.865 188.015 40.035 188.205 ;
        RECT 41.700 188.045 41.820 188.155 ;
        RECT 42.165 187.995 42.335 188.185 ;
        RECT 44.470 187.995 44.640 188.185 ;
        RECT 49.065 188.015 49.235 188.205 ;
        RECT 49.530 188.015 49.700 188.205 ;
        RECT 49.990 187.995 50.160 188.185 ;
        RECT 50.420 187.995 50.590 188.185 ;
        RECT 56.420 188.015 56.590 188.205 ;
        RECT 57.350 187.995 57.520 188.185 ;
        RECT 59.645 188.015 59.815 188.205 ;
        RECT 60.105 187.995 60.275 188.185 ;
        RECT 63.810 188.015 63.980 188.205 ;
        RECT 64.245 188.015 64.415 188.205 ;
        RECT 69.305 187.995 69.475 188.185 ;
        RECT 70.215 187.995 70.385 188.185 ;
        RECT 76.665 188.015 76.835 188.185 ;
        RECT 82.185 188.015 82.355 188.205 ;
        RECT 85.860 188.185 86.005 188.205 ;
        RECT 87.700 188.185 87.870 188.205 ;
        RECT 85.860 188.015 86.035 188.185 ;
        RECT 87.700 188.015 87.875 188.185 ;
        RECT 76.665 187.995 76.805 188.015 ;
        RECT 85.865 187.995 86.035 188.015 ;
        RECT 87.705 187.995 87.875 188.015 ;
        RECT 89.085 187.995 89.255 188.205 ;
        RECT 18.105 187.185 19.475 187.995 ;
        RECT 19.485 187.315 21.315 187.995 ;
        RECT 19.485 187.085 20.830 187.315 ;
        RECT 21.345 187.085 22.695 187.995 ;
        RECT 22.835 187.085 25.835 187.995 ;
        RECT 26.845 187.315 30.515 187.995 ;
        RECT 26.845 187.085 27.770 187.315 ;
        RECT 30.525 187.085 31.875 187.995 ;
        RECT 31.915 187.085 33.265 187.995 ;
        RECT 33.285 187.315 37.185 187.995 ;
        RECT 37.425 187.315 41.325 187.995 ;
        RECT 42.025 187.315 43.855 187.995 ;
        RECT 33.285 187.085 34.215 187.315 ;
        RECT 37.425 187.085 38.355 187.315 ;
        RECT 42.510 187.085 43.855 187.315 ;
        RECT 43.875 187.125 44.305 187.910 ;
        RECT 44.325 187.085 48.625 187.995 ;
        RECT 48.925 187.085 50.275 187.995 ;
        RECT 50.360 187.085 54.435 187.995 ;
        RECT 54.445 187.085 57.645 187.995 ;
        RECT 57.675 187.315 60.415 187.995 ;
        RECT 60.510 187.315 69.615 187.995 ;
        RECT 69.635 187.125 70.065 187.910 ;
        RECT 70.085 187.315 74.215 187.995 ;
        RECT 70.085 187.085 71.455 187.315 ;
        RECT 74.235 187.175 76.805 187.995 ;
        RECT 77.070 187.315 86.175 187.995 ;
        RECT 86.185 187.315 88.015 187.995 ;
        RECT 88.025 187.185 89.395 187.995 ;
        RECT 74.235 187.085 75.825 187.175 ;
      LAYER nwell ;
        RECT 17.910 183.965 89.590 186.795 ;
      LAYER pwell ;
        RECT 18.105 182.765 19.475 183.575 ;
        RECT 19.485 182.765 20.855 183.545 ;
        RECT 21.345 182.765 22.695 183.675 ;
        RECT 22.835 182.765 25.835 183.675 ;
        RECT 26.385 183.445 27.310 183.675 ;
        RECT 26.385 182.765 30.055 183.445 ;
        RECT 30.995 182.850 31.425 183.635 ;
        RECT 31.445 182.765 32.815 183.545 ;
        RECT 32.825 183.445 33.755 183.675 ;
        RECT 32.825 182.765 36.725 183.445 ;
        RECT 36.965 182.765 38.335 183.545 ;
        RECT 38.805 182.765 40.175 183.545 ;
        RECT 41.115 182.765 43.845 183.675 ;
        RECT 44.325 182.765 48.400 183.675 ;
        RECT 49.385 182.765 52.595 183.675 ;
        RECT 52.605 182.765 54.420 183.675 ;
        RECT 54.545 182.765 56.735 183.675 ;
        RECT 56.755 182.850 57.185 183.635 ;
        RECT 57.290 182.765 66.395 183.445 ;
        RECT 66.415 182.765 69.155 183.445 ;
        RECT 69.165 182.765 78.270 183.445 ;
        RECT 78.365 182.765 82.020 183.675 ;
        RECT 82.515 182.850 82.945 183.635 ;
        RECT 82.965 182.995 86.165 183.675 ;
        RECT 83.110 182.765 86.165 182.995 ;
        RECT 86.185 182.765 87.535 183.675 ;
        RECT 88.025 182.765 89.395 183.575 ;
        RECT 18.245 182.555 18.415 182.765 ;
        RECT 19.635 182.575 19.805 182.765 ;
        RECT 21.460 182.745 21.630 182.765 ;
        RECT 21.000 182.605 21.120 182.715 ;
        RECT 21.460 182.575 21.635 182.745 ;
        RECT 21.465 182.555 21.635 182.575 ;
        RECT 22.835 182.555 23.005 182.745 ;
        RECT 23.305 182.555 23.475 182.745 ;
        RECT 25.150 182.555 25.320 182.745 ;
        RECT 25.605 182.575 25.775 182.765 ;
        RECT 26.060 182.605 26.180 182.715 ;
        RECT 26.530 182.575 26.700 182.765 ;
        RECT 27.435 182.555 27.605 182.745 ;
        RECT 27.915 182.555 28.085 182.745 ;
        RECT 29.295 182.555 29.465 182.745 ;
        RECT 30.215 182.610 30.375 182.720 ;
        RECT 30.665 182.555 30.835 182.745 ;
        RECT 32.495 182.575 32.665 182.765 ;
        RECT 32.955 182.555 33.125 182.745 ;
        RECT 33.240 182.575 33.410 182.765 ;
        RECT 33.435 182.600 33.595 182.710 ;
        RECT 34.340 182.555 34.510 182.745 ;
        RECT 35.725 182.555 35.895 182.745 ;
        RECT 37.105 182.575 37.275 182.765 ;
        RECT 38.480 182.605 38.600 182.715 ;
        RECT 39.855 182.575 40.025 182.765 ;
        RECT 40.335 182.610 40.495 182.720 ;
        RECT 41.245 182.555 41.415 182.745 ;
        RECT 43.545 182.575 43.715 182.765 ;
        RECT 48.170 182.745 48.340 182.765 ;
        RECT 49.525 182.745 49.695 182.765 ;
        RECT 44.000 182.605 44.120 182.715 ;
        RECT 46.765 182.555 46.935 182.745 ;
        RECT 48.135 182.575 48.340 182.745 ;
        RECT 48.615 182.610 48.775 182.720 ;
        RECT 49.515 182.575 49.695 182.745 ;
        RECT 48.135 182.555 48.305 182.575 ;
        RECT 49.515 182.555 49.685 182.575 ;
        RECT 49.995 182.555 50.165 182.745 ;
        RECT 52.275 182.555 52.445 182.745 ;
        RECT 53.655 182.555 53.825 182.745 ;
        RECT 54.125 182.555 54.295 182.765 ;
        RECT 56.420 182.575 56.590 182.765 ;
        RECT 61.025 182.575 61.195 182.745 ;
        RECT 61.025 182.555 61.185 182.575 ;
        RECT 64.245 182.555 64.415 182.745 ;
        RECT 64.715 182.600 64.875 182.710 ;
        RECT 66.085 182.575 66.255 182.765 ;
        RECT 68.845 182.575 69.015 182.765 ;
        RECT 69.305 182.715 69.475 182.765 ;
        RECT 69.300 182.605 69.475 182.715 ;
        RECT 69.305 182.575 69.475 182.605 ;
        RECT 68.815 182.555 69.015 182.575 ;
        RECT 76.200 182.555 76.370 182.745 ;
        RECT 76.670 182.555 76.840 182.745 ;
        RECT 78.510 182.575 78.680 182.765 ;
        RECT 82.180 182.605 82.300 182.715 ;
        RECT 83.110 182.575 83.280 182.765 ;
        RECT 86.330 182.575 86.500 182.765 ;
        RECT 87.705 182.715 87.875 182.745 ;
        RECT 87.700 182.605 87.875 182.715 ;
        RECT 87.705 182.555 87.875 182.605 ;
        RECT 89.085 182.555 89.255 182.765 ;
        RECT 18.105 181.745 19.475 182.555 ;
        RECT 20.405 181.775 21.775 182.555 ;
        RECT 21.785 181.775 23.155 182.555 ;
        RECT 23.165 181.875 24.995 182.555 ;
        RECT 25.005 181.645 26.355 182.555 ;
        RECT 26.385 181.775 27.755 182.555 ;
        RECT 27.765 181.775 29.135 182.555 ;
        RECT 29.145 181.775 30.515 182.555 ;
        RECT 30.535 181.645 31.885 182.555 ;
        RECT 31.905 181.775 33.275 182.555 ;
        RECT 34.225 181.645 35.575 182.555 ;
        RECT 35.585 181.745 41.095 182.555 ;
        RECT 41.105 181.745 43.855 182.555 ;
        RECT 43.875 181.685 44.305 182.470 ;
        RECT 44.355 181.645 47.075 182.555 ;
        RECT 47.085 181.775 48.455 182.555 ;
        RECT 48.465 181.775 49.835 182.555 ;
        RECT 49.845 181.775 51.215 182.555 ;
        RECT 51.225 181.775 52.595 182.555 ;
        RECT 52.605 181.775 53.975 182.555 ;
        RECT 53.985 181.645 57.195 182.555 ;
        RECT 57.530 181.645 61.185 182.555 ;
        RECT 61.345 181.645 64.555 182.555 ;
        RECT 65.485 181.875 69.015 182.555 ;
        RECT 65.485 181.645 68.310 181.875 ;
        RECT 69.635 181.685 70.065 182.470 ;
        RECT 70.445 181.645 76.515 182.555 ;
        RECT 76.670 182.325 78.360 182.555 ;
        RECT 76.525 181.645 78.360 182.325 ;
        RECT 78.910 181.875 88.015 182.555 ;
        RECT 88.025 181.745 89.395 182.555 ;
      LAYER nwell ;
        RECT 17.910 178.525 89.590 181.355 ;
      LAYER pwell ;
        RECT 18.105 177.325 19.475 178.135 ;
        RECT 21.455 178.005 22.385 178.235 ;
        RECT 20.550 177.325 22.385 178.005 ;
        RECT 22.705 178.005 24.070 178.235 ;
        RECT 27.745 178.005 28.675 178.235 ;
        RECT 22.705 177.325 25.915 178.005 ;
        RECT 25.925 177.325 28.675 178.005 ;
        RECT 29.145 177.325 30.960 178.235 ;
        RECT 30.995 177.410 31.425 178.195 ;
        RECT 32.365 177.325 35.285 178.235 ;
        RECT 35.585 177.325 37.415 178.235 ;
        RECT 37.440 177.325 41.095 178.235 ;
        RECT 41.105 177.325 44.775 178.235 ;
        RECT 44.785 178.005 45.705 178.235 ;
        RECT 44.785 177.325 48.370 178.005 ;
        RECT 48.925 177.325 50.755 178.235 ;
        RECT 50.765 178.005 51.695 178.235 ;
        RECT 55.345 178.005 56.275 178.235 ;
        RECT 50.765 177.325 53.515 178.005 ;
        RECT 53.525 177.325 56.275 178.005 ;
        RECT 56.755 177.410 57.185 178.195 ;
        RECT 57.205 177.325 60.415 178.235 ;
        RECT 61.345 177.325 64.095 178.235 ;
        RECT 64.590 178.005 65.935 178.235 ;
        RECT 64.105 177.325 65.935 178.005 ;
        RECT 65.945 177.325 69.420 178.235 ;
        RECT 69.635 177.325 70.985 178.235 ;
        RECT 71.005 177.325 80.110 178.005 ;
        RECT 80.205 177.325 82.415 178.235 ;
        RECT 82.515 177.410 82.945 178.195 ;
        RECT 82.965 177.325 86.175 178.235 ;
        RECT 86.670 178.005 88.015 178.235 ;
        RECT 86.185 177.325 88.015 178.005 ;
        RECT 88.025 177.325 89.395 178.135 ;
        RECT 18.245 177.115 18.415 177.325 ;
        RECT 20.550 177.305 20.715 177.325 ;
        RECT 25.600 177.305 25.770 177.325 ;
        RECT 19.635 177.115 19.805 177.305 ;
        RECT 20.545 177.135 20.715 177.305 ;
        RECT 21.015 177.160 21.175 177.270 ;
        RECT 21.930 177.115 22.100 177.305 ;
        RECT 25.600 177.135 25.775 177.305 ;
        RECT 26.065 177.135 26.235 177.325 ;
        RECT 25.605 177.115 25.775 177.135 ;
        RECT 26.985 177.115 27.155 177.305 ;
        RECT 27.445 177.115 27.615 177.305 ;
        RECT 28.825 177.275 28.995 177.305 ;
        RECT 28.820 177.165 28.995 177.275 ;
        RECT 28.825 177.115 28.995 177.165 ;
        RECT 30.665 177.135 30.835 177.325 ;
        RECT 31.595 177.170 31.755 177.280 ;
        RECT 32.510 177.135 32.680 177.325 ;
        RECT 33.420 177.115 33.590 177.305 ;
        RECT 34.805 177.115 34.975 177.305 ;
        RECT 35.730 177.135 35.900 177.325 ;
        RECT 40.325 177.115 40.495 177.305 ;
        RECT 40.780 177.135 40.950 177.325 ;
        RECT 41.250 177.135 41.420 177.325 ;
        RECT 44.465 177.115 44.635 177.305 ;
        RECT 44.930 177.135 45.100 177.325 ;
        RECT 47.685 177.115 47.855 177.305 ;
        RECT 48.600 177.165 48.720 177.275 ;
        RECT 49.520 177.165 49.640 177.275 ;
        RECT 50.440 177.135 50.610 177.325 ;
        RECT 50.910 177.115 51.080 177.305 ;
        RECT 52.285 177.115 52.455 177.305 ;
        RECT 53.205 177.135 53.375 177.325 ;
        RECT 53.665 177.305 53.835 177.325 ;
        RECT 53.655 177.135 53.835 177.305 ;
        RECT 53.655 177.115 53.825 177.135 ;
        RECT 55.050 177.115 55.220 177.305 ;
        RECT 56.415 177.115 56.585 177.305 ;
        RECT 57.345 177.135 57.515 177.325 ;
        RECT 60.105 177.135 60.275 177.305 ;
        RECT 60.575 177.170 60.735 177.280 ;
        RECT 60.075 177.115 60.275 177.135 ;
        RECT 61.490 177.115 61.660 177.325 ;
        RECT 61.950 177.115 62.120 177.305 ;
        RECT 64.245 177.135 64.415 177.325 ;
        RECT 64.700 177.165 64.820 177.275 ;
        RECT 65.170 177.115 65.340 177.305 ;
        RECT 66.090 177.135 66.260 177.325 ;
        RECT 68.855 177.160 69.015 177.270 ;
        RECT 69.765 177.135 69.935 177.325 ;
        RECT 71.145 177.135 71.315 177.325 ;
        RECT 72.985 177.115 73.155 177.305 ;
        RECT 73.440 177.165 73.560 177.275 ;
        RECT 73.910 177.115 74.080 177.305 ;
        RECT 77.135 177.160 77.295 177.270 ;
        RECT 78.045 177.115 78.215 177.305 ;
        RECT 80.350 177.135 80.520 177.325 ;
        RECT 83.110 177.135 83.280 177.325 ;
        RECT 86.325 177.135 86.495 177.325 ;
        RECT 87.255 177.160 87.415 177.270 ;
        RECT 89.085 177.115 89.255 177.325 ;
        RECT 18.105 176.305 19.475 177.115 ;
        RECT 19.485 176.335 20.855 177.115 ;
        RECT 21.930 176.885 23.620 177.115 ;
        RECT 21.785 176.205 23.620 176.885 ;
        RECT 24.085 176.435 25.915 177.115 ;
        RECT 24.085 176.205 25.430 176.435 ;
        RECT 25.925 176.335 27.295 177.115 ;
        RECT 27.305 176.335 28.675 177.115 ;
        RECT 28.685 176.305 32.355 177.115 ;
        RECT 33.305 176.205 34.655 177.115 ;
        RECT 34.665 176.305 40.175 177.115 ;
        RECT 40.185 176.305 43.855 177.115 ;
        RECT 43.875 176.245 44.305 177.030 ;
        RECT 44.325 176.435 47.535 177.115 ;
        RECT 46.400 176.205 47.535 176.435 ;
        RECT 47.560 176.205 49.375 177.115 ;
        RECT 49.845 176.205 51.195 177.115 ;
        RECT 51.225 176.335 52.595 177.115 ;
        RECT 52.605 176.335 53.975 177.115 ;
        RECT 53.985 176.205 55.335 177.115 ;
        RECT 55.365 176.335 56.735 177.115 ;
        RECT 56.745 176.435 60.275 177.115 ;
        RECT 56.745 176.205 59.570 176.435 ;
        RECT 60.425 176.205 61.775 177.115 ;
        RECT 61.805 176.205 64.555 177.115 ;
        RECT 65.025 176.435 68.610 177.115 ;
        RECT 65.025 176.205 65.945 176.435 ;
        RECT 69.635 176.245 70.065 177.030 ;
        RECT 70.085 176.205 73.295 177.115 ;
        RECT 73.910 176.885 76.965 177.115 ;
        RECT 73.765 176.205 76.965 176.885 ;
        RECT 77.905 176.435 87.010 177.115 ;
        RECT 88.025 176.305 89.395 177.115 ;
      LAYER nwell ;
        RECT 17.910 173.085 89.590 175.915 ;
      LAYER pwell ;
        RECT 18.105 171.885 19.475 172.695 ;
        RECT 20.405 171.885 23.615 172.795 ;
        RECT 23.625 171.885 29.135 172.695 ;
        RECT 29.145 171.885 30.975 172.695 ;
        RECT 30.995 171.970 31.425 172.755 ;
        RECT 31.455 171.885 34.185 172.795 ;
        RECT 34.205 171.885 37.875 172.695 ;
        RECT 38.345 171.885 39.695 172.795 ;
        RECT 39.725 171.885 45.235 172.695 ;
        RECT 45.245 171.885 50.755 172.695 ;
        RECT 51.700 171.885 53.515 172.795 ;
        RECT 54.460 171.885 56.275 172.795 ;
        RECT 56.755 171.970 57.185 172.755 ;
        RECT 57.665 171.885 59.035 172.665 ;
        RECT 59.055 171.885 60.405 172.795 ;
        RECT 60.445 171.885 61.795 172.795 ;
        RECT 61.805 171.885 65.015 172.795 ;
        RECT 65.485 171.885 66.855 172.665 ;
        RECT 66.885 171.885 68.235 172.795 ;
        RECT 68.255 171.885 69.605 172.795 ;
        RECT 69.725 171.885 71.915 172.795 ;
        RECT 72.190 171.885 75.125 172.795 ;
        RECT 75.155 171.885 78.090 172.795 ;
        RECT 78.835 172.115 82.035 172.795 ;
        RECT 78.835 171.885 81.890 172.115 ;
        RECT 82.515 171.970 82.945 172.755 ;
        RECT 82.975 172.115 86.175 172.795 ;
        RECT 86.670 172.565 88.015 172.795 ;
        RECT 82.975 171.885 86.030 172.115 ;
        RECT 86.185 171.885 88.015 172.565 ;
        RECT 88.025 171.885 89.395 172.695 ;
        RECT 18.245 171.675 18.415 171.885 ;
        RECT 19.625 171.675 19.795 171.865 ;
        RECT 20.545 171.695 20.715 171.885 ;
        RECT 21.460 171.725 21.580 171.835 ;
        RECT 22.200 171.675 22.370 171.865 ;
        RECT 23.765 171.695 23.935 171.885 ;
        RECT 26.065 171.675 26.235 171.865 ;
        RECT 29.285 171.695 29.455 171.885 ;
        RECT 30.205 171.675 30.375 171.865 ;
        RECT 32.505 171.695 32.675 171.865 ;
        RECT 33.885 171.695 34.055 171.885 ;
        RECT 34.345 171.695 34.515 171.885 ;
        RECT 32.505 171.675 32.670 171.695 ;
        RECT 35.725 171.675 35.895 171.865 ;
        RECT 36.195 171.720 36.355 171.830 ;
        RECT 37.380 171.675 37.550 171.865 ;
        RECT 38.020 171.725 38.140 171.835 ;
        RECT 39.410 171.695 39.580 171.885 ;
        RECT 39.865 171.695 40.035 171.885 ;
        RECT 41.245 171.675 41.415 171.865 ;
        RECT 45.385 171.695 45.555 171.885 ;
        RECT 45.845 171.675 46.015 171.865 ;
        RECT 46.300 171.725 46.420 171.835 ;
        RECT 46.765 171.675 46.935 171.865 ;
        RECT 49.525 171.675 49.695 171.865 ;
        RECT 50.915 171.730 51.075 171.840 ;
        RECT 51.825 171.695 51.995 171.885 ;
        RECT 52.285 171.675 52.455 171.865 ;
        RECT 53.675 171.730 53.835 171.840 ;
        RECT 54.135 171.720 54.295 171.830 ;
        RECT 54.585 171.695 54.755 171.885 ;
        RECT 55.045 171.675 55.215 171.865 ;
        RECT 56.420 171.725 56.540 171.835 ;
        RECT 56.895 171.720 57.055 171.830 ;
        RECT 57.340 171.725 57.460 171.835 ;
        RECT 58.715 171.675 58.885 171.885 ;
        RECT 59.185 171.695 59.355 171.885 ;
        RECT 60.560 171.695 60.730 171.885 ;
        RECT 62.405 171.695 62.575 171.865 ;
        RECT 62.375 171.675 62.575 171.695 ;
        RECT 62.865 171.675 63.035 171.865 ;
        RECT 64.705 171.695 64.875 171.885 ;
        RECT 65.165 171.835 65.335 171.865 ;
        RECT 65.160 171.725 65.335 171.835 ;
        RECT 65.165 171.675 65.335 171.725 ;
        RECT 65.635 171.675 65.805 171.865 ;
        RECT 66.535 171.695 66.705 171.885 ;
        RECT 67.920 171.865 68.090 171.885 ;
        RECT 67.915 171.695 68.090 171.865 ;
        RECT 67.915 171.675 68.085 171.695 ;
        RECT 68.385 171.675 68.555 171.885 ;
        RECT 70.220 171.725 70.340 171.835 ;
        RECT 70.695 171.675 70.865 171.865 ;
        RECT 71.600 171.695 71.770 171.885 ;
        RECT 72.190 171.865 72.235 171.885 ;
        RECT 78.045 171.865 78.090 171.885 ;
        RECT 72.065 171.695 72.235 171.865 ;
        RECT 72.985 171.675 73.155 171.865 ;
        RECT 76.665 171.675 76.835 171.865 ;
        RECT 77.125 171.675 77.295 171.865 ;
        RECT 78.045 171.695 78.215 171.865 ;
        RECT 78.500 171.725 78.620 171.835 ;
        RECT 78.965 171.675 79.135 171.865 ;
        RECT 81.720 171.695 81.890 171.885 ;
        RECT 82.180 171.725 82.300 171.835 ;
        RECT 85.860 171.695 86.030 171.885 ;
        RECT 86.325 171.695 86.495 171.885 ;
        RECT 89.085 171.675 89.255 171.885 ;
        RECT 18.105 170.865 19.475 171.675 ;
        RECT 19.485 170.865 21.315 171.675 ;
        RECT 21.785 170.995 25.685 171.675 ;
        RECT 21.785 170.765 22.715 170.995 ;
        RECT 25.925 170.865 28.675 171.675 ;
        RECT 28.685 170.765 30.500 171.675 ;
        RECT 30.835 170.995 32.670 171.675 ;
        RECT 30.835 170.765 31.765 170.995 ;
        RECT 32.825 170.765 36.035 171.675 ;
        RECT 36.965 170.995 40.865 171.675 ;
        RECT 36.965 170.765 37.895 170.995 ;
        RECT 41.105 170.865 43.855 171.675 ;
        RECT 43.875 170.805 44.305 171.590 ;
        RECT 44.325 170.765 46.140 171.675 ;
        RECT 46.635 170.765 49.365 171.675 ;
        RECT 49.385 170.865 52.135 171.675 ;
        RECT 52.160 170.765 53.975 171.675 ;
        RECT 54.920 170.765 56.735 171.675 ;
        RECT 57.665 170.895 59.035 171.675 ;
        RECT 59.045 170.995 62.575 171.675 ;
        RECT 59.045 170.765 61.870 170.995 ;
        RECT 62.725 170.895 64.095 171.675 ;
        RECT 64.105 170.895 65.475 171.675 ;
        RECT 65.485 170.895 66.855 171.675 ;
        RECT 66.865 170.895 68.235 171.675 ;
        RECT 68.245 170.895 69.615 171.675 ;
        RECT 69.635 170.805 70.065 171.590 ;
        RECT 70.545 170.895 71.915 171.675 ;
        RECT 71.935 170.765 73.285 171.675 ;
        RECT 73.445 170.765 76.895 171.675 ;
        RECT 76.985 170.995 78.815 171.675 ;
        RECT 78.825 170.995 87.930 171.675 ;
        RECT 77.470 170.765 78.815 170.995 ;
        RECT 88.025 170.865 89.395 171.675 ;
      LAYER nwell ;
        RECT 17.910 167.645 89.590 170.475 ;
      LAYER pwell ;
        RECT 18.105 166.445 19.475 167.255 ;
        RECT 19.485 166.445 21.315 167.255 ;
        RECT 21.325 167.125 22.255 167.355 ;
        RECT 21.325 166.445 25.225 167.125 ;
        RECT 25.465 166.445 28.215 167.255 ;
        RECT 28.225 166.445 30.040 167.355 ;
        RECT 30.995 166.530 31.425 167.315 ;
        RECT 31.755 167.125 32.685 167.355 ;
        RECT 31.755 166.445 33.590 167.125 ;
        RECT 33.745 166.445 35.560 167.355 ;
        RECT 36.505 167.125 37.435 167.355 ;
        RECT 36.505 166.445 40.405 167.125 ;
        RECT 40.655 166.445 42.005 167.355 ;
        RECT 42.025 166.445 43.375 167.355 ;
        RECT 44.325 166.445 46.140 167.355 ;
        RECT 46.175 166.445 47.525 167.355 ;
        RECT 47.545 166.445 48.915 167.255 ;
        RECT 48.925 166.445 50.275 167.355 ;
        RECT 50.305 166.445 55.815 167.255 ;
        RECT 56.755 166.530 57.185 167.315 ;
        RECT 57.205 167.155 58.150 167.355 ;
        RECT 59.485 167.155 60.415 167.355 ;
        RECT 57.205 166.675 60.415 167.155 ;
        RECT 57.205 166.475 60.275 166.675 ;
        RECT 57.205 166.445 58.150 166.475 ;
        RECT 18.245 166.235 18.415 166.445 ;
        RECT 19.625 166.235 19.795 166.445 ;
        RECT 21.740 166.255 21.910 166.445 ;
        RECT 25.605 166.255 25.775 166.445 ;
        RECT 25.790 166.235 25.960 166.425 ;
        RECT 29.285 166.235 29.455 166.425 ;
        RECT 29.745 166.235 29.915 166.445 ;
        RECT 33.425 166.425 33.590 166.445 ;
        RECT 30.215 166.290 30.375 166.400 ;
        RECT 33.425 166.255 33.595 166.425 ;
        RECT 35.265 166.235 35.435 166.445 ;
        RECT 35.735 166.290 35.895 166.400 ;
        RECT 36.920 166.255 37.090 166.445 ;
        RECT 40.785 166.235 40.955 166.445 ;
        RECT 43.090 166.255 43.260 166.445 ;
        RECT 43.555 166.395 43.715 166.400 ;
        RECT 43.540 166.290 43.715 166.395 ;
        RECT 43.540 166.285 43.660 166.290 ;
        RECT 44.465 166.235 44.635 166.425 ;
        RECT 45.845 166.255 46.015 166.445 ;
        RECT 46.305 166.255 46.475 166.445 ;
        RECT 47.685 166.425 47.855 166.445 ;
        RECT 47.220 166.285 47.340 166.395 ;
        RECT 47.685 166.255 47.860 166.425 ;
        RECT 49.990 166.255 50.160 166.445 ;
        RECT 50.445 166.255 50.615 166.445 ;
        RECT 47.690 166.235 47.860 166.255 ;
        RECT 51.365 166.235 51.535 166.425 ;
        RECT 53.210 166.235 53.380 166.425 ;
        RECT 55.975 166.290 56.135 166.400 ;
        RECT 59.640 166.235 59.810 166.425 ;
        RECT 60.105 166.255 60.275 166.475 ;
        RECT 60.425 166.445 62.255 167.255 ;
        RECT 62.725 166.445 65.935 167.355 ;
        RECT 65.960 166.445 69.615 167.355 ;
        RECT 69.625 166.445 71.440 167.355 ;
        RECT 72.515 166.445 75.515 167.355 ;
        RECT 77.430 167.125 78.800 167.355 ;
        RECT 76.525 166.445 78.800 167.125 ;
        RECT 78.835 166.445 81.575 167.125 ;
        RECT 82.515 166.530 82.945 167.315 ;
        RECT 83.045 166.445 85.255 167.355 ;
        RECT 85.265 166.445 88.005 167.125 ;
        RECT 88.025 166.445 89.395 167.255 ;
        RECT 60.565 166.255 60.735 166.445 ;
        RECT 62.400 166.285 62.520 166.395 ;
        RECT 62.855 166.255 63.025 166.445 ;
        RECT 60.110 166.235 60.275 166.255 ;
        RECT 63.330 166.235 63.500 166.425 ;
        RECT 63.785 166.235 63.955 166.425 ;
        RECT 66.545 166.235 66.715 166.425 ;
        RECT 68.395 166.235 68.565 166.425 ;
        RECT 69.300 166.255 69.470 166.445 ;
        RECT 70.235 166.280 70.395 166.390 ;
        RECT 71.145 166.235 71.315 166.445 ;
        RECT 71.615 166.290 71.775 166.400 ;
        RECT 72.525 166.235 72.695 166.425 ;
        RECT 73.905 166.235 74.075 166.425 ;
        RECT 75.285 166.255 75.455 166.445 ;
        RECT 75.755 166.290 75.915 166.400 ;
        RECT 76.670 166.255 76.840 166.445 ;
        RECT 18.105 165.425 19.475 166.235 ;
        RECT 19.485 165.425 22.235 166.235 ;
        RECT 22.475 165.555 26.375 166.235 ;
        RECT 25.445 165.325 26.375 165.555 ;
        RECT 26.385 165.325 29.595 166.235 ;
        RECT 29.605 165.425 35.115 166.235 ;
        RECT 35.125 165.425 40.635 166.235 ;
        RECT 40.645 165.425 43.395 166.235 ;
        RECT 43.875 165.365 44.305 166.150 ;
        RECT 44.325 165.425 47.075 166.235 ;
        RECT 47.545 165.555 51.215 166.235 ;
        RECT 47.545 165.325 48.470 165.555 ;
        RECT 51.225 165.425 53.055 166.235 ;
        RECT 53.065 165.325 55.985 166.235 ;
        RECT 56.480 165.325 59.955 166.235 ;
        RECT 60.110 165.555 61.945 166.235 ;
        RECT 61.015 165.325 61.945 165.555 ;
        RECT 62.265 165.325 63.615 166.235 ;
        RECT 63.645 165.425 66.395 166.235 ;
        RECT 66.420 165.325 68.235 166.235 ;
        RECT 68.245 165.455 69.615 166.235 ;
        RECT 69.635 165.365 70.065 166.150 ;
        RECT 71.005 165.455 72.375 166.235 ;
        RECT 72.385 165.455 73.755 166.235 ;
        RECT 73.845 165.325 77.295 166.235 ;
        RECT 77.580 166.205 77.750 166.425 ;
        RECT 79.895 166.280 80.055 166.390 ;
        RECT 80.805 166.235 80.975 166.425 ;
        RECT 81.265 166.255 81.435 166.445 ;
        RECT 81.735 166.290 81.895 166.400 ;
        RECT 84.940 166.255 85.110 166.445 ;
        RECT 85.405 166.255 85.575 166.445 ;
        RECT 78.780 166.205 79.735 166.235 ;
        RECT 77.455 165.525 79.735 166.205 ;
        RECT 80.665 165.555 83.415 166.235 ;
        RECT 78.780 165.325 79.735 165.525 ;
        RECT 82.485 165.325 83.415 165.555 ;
        RECT 83.425 166.205 84.820 166.235 ;
        RECT 85.865 166.205 86.035 166.425 ;
        RECT 86.325 166.235 86.495 166.425 ;
        RECT 89.085 166.235 89.255 166.445 ;
        RECT 83.425 165.525 86.160 166.205 ;
        RECT 86.185 165.555 88.015 166.235 ;
        RECT 83.425 165.325 84.835 165.525 ;
        RECT 86.670 165.325 88.015 165.555 ;
        RECT 88.025 165.425 89.395 166.235 ;
      LAYER nwell ;
        RECT 17.910 162.205 89.590 165.035 ;
      LAYER pwell ;
        RECT 18.105 161.005 19.475 161.815 ;
        RECT 19.485 161.005 22.235 161.815 ;
        RECT 25.445 161.685 26.375 161.915 ;
        RECT 22.475 161.005 26.375 161.685 ;
        RECT 26.385 161.005 29.135 161.815 ;
        RECT 29.605 161.005 30.955 161.915 ;
        RECT 30.995 161.090 31.425 161.875 ;
        RECT 31.445 161.005 34.655 161.915 ;
        RECT 35.125 161.685 36.055 161.915 ;
        RECT 35.125 161.005 39.025 161.685 ;
        RECT 39.265 161.005 40.615 161.915 ;
        RECT 40.645 161.005 43.395 161.815 ;
        RECT 43.405 161.005 46.615 161.915 ;
        RECT 46.625 161.005 52.135 161.815 ;
        RECT 52.145 161.005 55.815 161.815 ;
        RECT 56.755 161.090 57.185 161.875 ;
        RECT 57.205 161.715 58.150 161.915 ;
        RECT 59.485 161.715 60.415 161.915 ;
        RECT 57.205 161.235 60.415 161.715 ;
        RECT 57.205 161.035 60.275 161.235 ;
        RECT 57.205 161.005 58.150 161.035 ;
        RECT 18.245 160.795 18.415 161.005 ;
        RECT 19.625 160.815 19.795 161.005 ;
        RECT 21.005 160.795 21.175 160.985 ;
        RECT 21.465 160.795 21.635 160.985 ;
        RECT 24.225 160.795 24.395 160.985 ;
        RECT 24.685 160.795 24.855 160.985 ;
        RECT 25.790 160.815 25.960 161.005 ;
        RECT 26.525 160.815 26.695 161.005 ;
        RECT 29.280 160.845 29.400 160.955 ;
        RECT 30.200 160.845 30.320 160.955 ;
        RECT 30.670 160.815 30.840 161.005 ;
        RECT 31.585 160.795 31.755 160.985 ;
        RECT 32.045 160.815 32.215 160.985 ;
        RECT 34.345 160.815 34.515 161.005 ;
        RECT 34.800 160.845 34.920 160.955 ;
        RECT 32.075 160.795 32.215 160.815 ;
        RECT 35.080 160.795 35.250 160.985 ;
        RECT 35.540 160.815 35.710 161.005 ;
        RECT 38.945 160.795 39.115 160.985 ;
        RECT 40.330 160.815 40.500 161.005 ;
        RECT 40.785 160.815 40.955 161.005 ;
        RECT 43.095 160.840 43.255 160.950 ;
        RECT 43.535 160.815 43.705 161.005 ;
        RECT 46.765 160.815 46.935 161.005 ;
        RECT 48.145 160.815 48.315 160.985 ;
        RECT 40.790 160.795 40.955 160.815 ;
        RECT 48.145 160.795 48.305 160.815 ;
        RECT 51.820 160.795 51.990 160.985 ;
        RECT 52.285 160.795 52.455 161.005 ;
        RECT 55.505 160.795 55.675 160.985 ;
        RECT 55.975 160.850 56.135 160.960 ;
        RECT 60.105 160.815 60.275 161.035 ;
        RECT 60.425 161.005 65.935 161.815 ;
        RECT 65.945 161.005 69.615 161.815 ;
        RECT 69.625 161.005 70.995 161.815 ;
        RECT 60.565 160.815 60.735 161.005 ;
        RECT 61.030 160.795 61.200 160.985 ;
        RECT 66.085 160.815 66.255 161.005 ;
        RECT 67.925 160.795 68.095 160.985 ;
        RECT 68.385 160.795 68.555 160.985 ;
        RECT 69.765 160.815 69.935 161.005 ;
        RECT 70.225 160.795 70.395 160.985 ;
        RECT 71.005 160.965 71.895 161.915 ;
        RECT 73.295 161.685 74.215 161.915 ;
        RECT 71.925 161.005 74.215 161.685 ;
        RECT 74.245 161.005 75.595 161.915 ;
        RECT 76.065 161.005 77.435 161.785 ;
        RECT 78.780 161.715 79.735 161.915 ;
        RECT 77.455 161.035 79.735 161.715 ;
        RECT 71.605 160.815 71.775 160.965 ;
        RECT 72.065 160.815 72.235 161.005 ;
        RECT 73.445 160.795 73.615 160.985 ;
        RECT 75.280 160.815 75.450 161.005 ;
        RECT 75.745 160.955 75.915 160.985 ;
        RECT 75.740 160.845 75.915 160.955 ;
        RECT 75.745 160.795 75.915 160.845 ;
        RECT 76.215 160.815 76.385 161.005 ;
        RECT 77.580 160.815 77.750 161.035 ;
        RECT 78.780 161.005 79.735 161.035 ;
        RECT 80.285 161.005 82.495 161.915 ;
        RECT 82.515 161.090 82.945 161.875 ;
        RECT 82.975 161.005 84.325 161.915 ;
        RECT 84.425 161.005 88.010 161.915 ;
        RECT 88.025 161.005 89.395 161.815 ;
        RECT 78.055 160.840 78.215 160.950 ;
        RECT 78.965 160.795 79.135 160.985 ;
        RECT 79.880 160.845 80.000 160.955 ;
        RECT 82.180 160.815 82.350 161.005 ;
        RECT 83.105 160.815 83.275 161.005 ;
        RECT 87.700 160.815 87.870 161.005 ;
        RECT 89.085 160.795 89.255 161.005 ;
        RECT 18.105 159.985 19.475 160.795 ;
        RECT 19.485 160.115 21.315 160.795 ;
        RECT 21.325 160.115 23.155 160.795 ;
        RECT 19.485 159.885 20.830 160.115 ;
        RECT 23.165 160.015 24.535 160.795 ;
        RECT 24.545 159.985 30.055 160.795 ;
        RECT 30.535 159.885 31.885 160.795 ;
        RECT 32.075 159.975 34.645 160.795 ;
        RECT 33.055 159.885 34.645 159.975 ;
        RECT 34.665 160.115 38.565 160.795 ;
        RECT 34.665 159.885 35.595 160.115 ;
        RECT 38.805 159.985 40.635 160.795 ;
        RECT 40.790 160.115 42.625 160.795 ;
        RECT 41.695 159.885 42.625 160.115 ;
        RECT 43.875 159.925 44.305 160.710 ;
        RECT 44.650 159.885 48.305 160.795 ;
        RECT 48.465 159.885 52.135 160.795 ;
        RECT 52.145 159.885 55.355 160.795 ;
        RECT 55.365 159.985 60.875 160.795 ;
        RECT 60.885 159.885 65.275 160.795 ;
        RECT 65.495 159.885 68.225 160.795 ;
        RECT 68.245 159.985 69.615 160.795 ;
        RECT 69.635 159.925 70.065 160.710 ;
        RECT 70.085 159.885 73.295 160.795 ;
        RECT 73.305 160.115 75.595 160.795 ;
        RECT 75.605 160.115 77.895 160.795 ;
        RECT 78.825 160.115 87.930 160.795 ;
        RECT 74.675 159.885 75.595 160.115 ;
        RECT 76.975 159.885 77.895 160.115 ;
        RECT 88.025 159.985 89.395 160.795 ;
      LAYER nwell ;
        RECT 17.910 156.765 89.590 159.595 ;
      LAYER pwell ;
        RECT 18.105 155.565 19.475 156.375 ;
        RECT 20.405 155.565 22.235 156.475 ;
        RECT 24.090 156.245 25.455 156.475 ;
        RECT 22.245 155.565 25.455 156.245 ;
        RECT 25.465 155.565 27.295 156.475 ;
        RECT 27.305 155.565 30.975 156.375 ;
        RECT 30.995 155.650 31.425 156.435 ;
        RECT 31.445 156.245 32.790 156.475 ;
        RECT 39.025 156.385 39.975 156.475 ;
        RECT 31.445 155.565 33.275 156.245 ;
        RECT 33.285 155.565 36.955 156.375 ;
        RECT 38.045 155.565 39.975 156.385 ;
        RECT 40.185 155.565 45.695 156.375 ;
        RECT 45.705 155.565 47.535 156.375 ;
        RECT 47.545 155.565 50.295 156.475 ;
        RECT 50.305 155.565 52.135 156.375 ;
        RECT 53.990 156.245 55.355 156.475 ;
        RECT 52.145 155.565 55.355 156.245 ;
        RECT 55.365 155.565 56.735 156.375 ;
        RECT 56.755 155.650 57.185 156.435 ;
        RECT 57.635 155.565 60.415 156.475 ;
        RECT 60.425 155.565 62.255 156.375 ;
        RECT 62.725 155.565 64.540 156.475 ;
        RECT 66.830 156.275 67.775 156.475 ;
        RECT 65.025 155.595 67.775 156.275 ;
        RECT 18.245 155.355 18.415 155.565 ;
        RECT 19.600 155.520 19.770 155.545 ;
        RECT 19.600 155.410 19.795 155.520 ;
        RECT 19.600 155.375 19.770 155.410 ;
        RECT 20.550 155.375 20.720 155.565 ;
        RECT 22.390 155.375 22.560 155.565 ;
        RECT 24.235 155.400 24.395 155.510 ;
        RECT 19.660 155.355 19.770 155.375 ;
        RECT 25.145 155.355 25.315 155.545 ;
        RECT 26.980 155.375 27.150 155.565 ;
        RECT 27.445 155.375 27.615 155.565 ;
        RECT 28.825 155.355 28.995 155.545 ;
        RECT 32.965 155.375 33.135 155.565 ;
        RECT 33.425 155.355 33.595 155.565 ;
        RECT 38.045 155.545 38.195 155.565 ;
        RECT 37.115 155.410 37.275 155.520 ;
        RECT 38.025 155.375 38.195 155.545 ;
        RECT 39.405 155.355 39.575 155.545 ;
        RECT 39.865 155.355 40.035 155.545 ;
        RECT 40.325 155.375 40.495 155.565 ;
        RECT 43.540 155.405 43.660 155.515 ;
        RECT 44.455 155.355 44.625 155.545 ;
        RECT 45.845 155.375 46.015 155.565 ;
        RECT 47.685 155.355 47.855 155.565 ;
        RECT 50.445 155.355 50.615 155.565 ;
        RECT 52.290 155.375 52.460 155.565 ;
        RECT 53.200 155.355 53.370 155.545 ;
        RECT 53.665 155.355 53.835 155.545 ;
        RECT 55.505 155.375 55.675 155.565 ;
        RECT 59.185 155.355 59.355 155.545 ;
        RECT 60.105 155.375 60.275 155.565 ;
        RECT 60.565 155.375 60.735 155.565 ;
        RECT 62.400 155.405 62.520 155.515 ;
        RECT 62.865 155.355 63.035 155.545 ;
        RECT 64.245 155.375 64.415 155.565 ;
        RECT 65.170 155.545 65.340 155.595 ;
        RECT 66.830 155.565 67.775 155.595 ;
        RECT 67.785 155.565 70.535 156.375 ;
        RECT 72.375 156.245 73.295 156.475 ;
        RECT 71.005 155.565 73.295 156.245 ;
        RECT 73.325 155.565 74.675 156.475 ;
        RECT 74.685 155.565 78.355 156.375 ;
        RECT 79.285 155.565 80.655 156.345 ;
        RECT 80.665 155.565 82.495 156.245 ;
        RECT 82.515 155.650 82.945 156.435 ;
        RECT 83.910 156.245 85.250 156.475 ;
        RECT 83.425 155.565 88.015 156.245 ;
        RECT 88.025 155.565 89.395 156.375 ;
        RECT 64.700 155.405 64.820 155.515 ;
        RECT 65.165 155.375 65.340 155.545 ;
        RECT 65.165 155.355 65.335 155.375 ;
        RECT 65.625 155.355 65.795 155.545 ;
        RECT 67.925 155.375 68.095 155.565 ;
        RECT 69.300 155.405 69.420 155.515 ;
        RECT 70.680 155.405 70.800 155.515 ;
        RECT 71.145 155.375 71.315 155.565 ;
        RECT 72.525 155.355 72.695 155.545 ;
        RECT 74.360 155.375 74.530 155.565 ;
        RECT 74.825 155.375 74.995 155.565 ;
        RECT 74.825 155.355 74.975 155.375 ;
        RECT 75.285 155.355 75.455 155.545 ;
        RECT 78.515 155.410 78.675 155.520 ;
        RECT 79.435 155.375 79.605 155.565 ;
        RECT 80.815 155.400 80.975 155.510 ;
        RECT 82.185 155.375 82.355 155.565 ;
        RECT 82.635 155.355 82.805 155.545 ;
        RECT 83.115 155.515 83.285 155.545 ;
        RECT 83.100 155.405 83.285 155.515 ;
        RECT 83.115 155.355 83.285 155.405 ;
        RECT 83.570 155.375 83.740 155.565 ;
        RECT 85.865 155.355 86.035 155.545 ;
        RECT 86.325 155.355 86.495 155.545 ;
        RECT 89.085 155.355 89.255 155.565 ;
        RECT 18.105 154.545 19.475 155.355 ;
        RECT 19.660 154.675 24.075 155.355 ;
        RECT 25.005 154.675 28.675 155.355 ;
        RECT 28.685 155.125 30.255 155.355 ;
        RECT 32.345 155.315 33.265 155.355 ;
        RECT 32.345 155.125 33.275 155.315 ;
        RECT 28.685 154.765 33.275 155.125 ;
        RECT 28.685 154.675 33.265 154.765 ;
        RECT 20.145 154.445 24.075 154.675 ;
        RECT 27.745 154.445 28.675 154.675 ;
        RECT 30.265 154.445 33.265 154.675 ;
        RECT 33.285 154.545 36.035 155.355 ;
        RECT 36.185 154.445 39.635 155.355 ;
        RECT 39.725 154.545 43.395 155.355 ;
        RECT 43.875 154.485 44.305 155.270 ;
        RECT 44.325 154.445 47.535 155.355 ;
        RECT 47.555 154.445 50.285 155.355 ;
        RECT 50.305 154.545 52.135 155.355 ;
        RECT 52.165 154.445 53.515 155.355 ;
        RECT 53.525 154.545 59.035 155.355 ;
        RECT 59.045 154.545 62.715 155.355 ;
        RECT 62.725 154.545 64.095 155.355 ;
        RECT 64.115 154.445 65.465 155.355 ;
        RECT 65.485 154.545 69.155 155.355 ;
        RECT 69.635 154.485 70.065 155.270 ;
        RECT 70.095 154.445 72.825 155.355 ;
        RECT 73.045 154.535 74.975 155.355 ;
        RECT 75.145 154.545 80.655 155.355 ;
        RECT 81.585 154.575 82.955 155.355 ;
        RECT 82.965 154.575 84.335 155.355 ;
        RECT 84.345 154.675 86.175 155.355 ;
        RECT 86.185 154.675 88.015 155.355 ;
        RECT 73.045 154.445 73.995 154.535 ;
        RECT 84.345 154.445 85.690 154.675 ;
        RECT 86.670 154.445 88.015 154.675 ;
        RECT 88.025 154.545 89.395 155.355 ;
      LAYER nwell ;
        RECT 17.910 151.325 89.590 154.155 ;
      LAYER pwell ;
        RECT 19.495 150.945 21.085 151.035 ;
        RECT 18.105 150.125 19.475 150.935 ;
        RECT 19.495 150.125 22.065 150.945 ;
        RECT 24.065 150.805 24.995 151.035 ;
        RECT 22.245 150.125 24.995 150.805 ;
        RECT 25.005 150.125 26.835 150.935 ;
        RECT 27.305 150.835 28.235 151.035 ;
        RECT 29.565 150.835 30.515 151.035 ;
        RECT 27.305 150.355 30.515 150.835 ;
        RECT 27.450 150.155 30.515 150.355 ;
        RECT 30.995 150.210 31.425 150.995 ;
        RECT 31.445 150.835 32.375 151.035 ;
        RECT 33.705 150.835 34.655 151.035 ;
        RECT 31.445 150.355 34.655 150.835 ;
        RECT 18.245 149.915 18.415 150.125 ;
        RECT 21.925 150.105 22.065 150.125 ;
        RECT 21.005 149.915 21.175 150.105 ;
        RECT 21.465 149.915 21.635 150.105 ;
        RECT 21.925 149.935 22.095 150.105 ;
        RECT 22.385 149.935 22.555 150.125 ;
        RECT 23.765 149.915 23.935 150.105 ;
        RECT 24.225 149.915 24.395 150.105 ;
        RECT 25.145 149.935 25.315 150.125 ;
        RECT 26.980 149.965 27.100 150.075 ;
        RECT 27.450 149.935 27.620 150.155 ;
        RECT 29.580 150.125 30.515 150.155 ;
        RECT 31.590 150.155 34.655 150.355 ;
        RECT 29.745 149.915 29.915 150.105 ;
        RECT 30.660 149.965 30.780 150.075 ;
        RECT 31.590 149.935 31.760 150.155 ;
        RECT 33.720 150.125 34.655 150.155 ;
        RECT 35.595 150.125 39.715 151.035 ;
        RECT 39.725 150.125 41.555 150.805 ;
        RECT 41.585 150.125 42.935 151.035 ;
        RECT 44.545 150.945 45.495 151.035 ;
        RECT 43.565 150.125 45.495 150.945 ;
        RECT 45.705 150.355 47.540 151.035 ;
        RECT 45.850 150.125 47.540 150.355 ;
        RECT 48.005 150.125 49.835 150.935 ;
        RECT 50.305 150.125 53.975 151.035 ;
        RECT 54.470 150.805 55.815 151.035 ;
        RECT 53.985 150.125 55.815 150.805 ;
        RECT 56.755 150.210 57.185 150.995 ;
        RECT 57.205 150.125 60.415 151.035 ;
        RECT 60.465 150.805 61.840 151.035 ;
        RECT 63.630 150.805 65.010 151.035 ;
        RECT 60.465 150.355 65.010 150.805 ;
        RECT 34.815 149.970 34.975 150.080 ;
        RECT 35.265 149.915 35.435 150.105 ;
        RECT 37.105 149.915 37.275 150.105 ;
        RECT 37.565 149.935 37.735 150.125 ;
        RECT 38.945 149.915 39.115 150.105 ;
        RECT 39.405 149.935 39.575 150.125 ;
        RECT 41.245 149.935 41.415 150.125 ;
        RECT 42.620 150.105 42.790 150.125 ;
        RECT 43.565 150.105 43.715 150.125 ;
        RECT 42.620 149.935 42.795 150.105 ;
        RECT 43.080 149.965 43.200 150.075 ;
        RECT 43.545 149.935 43.715 150.105 ;
        RECT 42.625 149.915 42.795 149.935 ;
        RECT 44.465 149.915 44.635 150.105 ;
        RECT 45.850 149.935 46.020 150.125 ;
        RECT 48.145 149.935 48.315 150.125 ;
        RECT 49.980 149.965 50.100 150.075 ;
        RECT 50.445 149.915 50.615 150.125 ;
        RECT 54.125 149.935 54.295 150.125 ;
        RECT 55.965 149.935 56.135 150.105 ;
        RECT 55.965 149.915 56.130 149.935 ;
        RECT 56.430 149.915 56.600 150.105 ;
        RECT 57.345 149.935 57.515 150.125 ;
        RECT 57.805 149.915 57.975 150.105 ;
        RECT 60.570 149.935 60.740 150.355 ;
        RECT 61.850 150.125 65.010 150.355 ;
        RECT 65.025 150.125 66.375 151.035 ;
        RECT 66.405 150.125 67.775 150.935 ;
        RECT 67.795 150.125 70.525 151.035 ;
        RECT 70.545 150.125 72.360 151.035 ;
        RECT 72.385 150.125 77.895 150.935 ;
        RECT 77.905 150.125 81.575 150.935 ;
        RECT 82.515 150.210 82.945 150.995 ;
        RECT 82.965 150.125 84.795 150.935 ;
        RECT 84.805 150.125 86.175 150.905 ;
        RECT 86.185 150.125 88.015 150.805 ;
        RECT 88.025 150.125 89.395 150.935 ;
        RECT 61.020 149.915 61.190 150.105 ;
        RECT 62.405 149.915 62.575 150.105 ;
        RECT 66.090 149.935 66.260 150.125 ;
        RECT 66.545 149.935 66.715 150.125 ;
        RECT 69.305 149.915 69.475 150.105 ;
        RECT 70.225 149.915 70.395 150.125 ;
        RECT 72.065 149.935 72.235 150.125 ;
        RECT 72.525 149.935 72.695 150.125 ;
        RECT 75.745 149.915 75.915 150.105 ;
        RECT 78.045 149.935 78.215 150.125 ;
        RECT 81.265 149.915 81.435 150.105 ;
        RECT 81.735 149.970 81.895 150.080 ;
        RECT 83.105 149.935 83.275 150.125 ;
        RECT 84.955 149.935 85.125 150.125 ;
        RECT 86.325 149.935 86.495 150.125 ;
        RECT 87.705 149.915 87.875 150.105 ;
        RECT 89.085 149.915 89.255 150.125 ;
        RECT 18.105 149.105 19.475 149.915 ;
        RECT 19.485 149.235 21.315 149.915 ;
        RECT 19.485 149.005 20.830 149.235 ;
        RECT 21.335 149.005 22.685 149.915 ;
        RECT 22.705 149.135 24.075 149.915 ;
        RECT 24.085 149.105 29.595 149.915 ;
        RECT 29.605 149.105 35.115 149.915 ;
        RECT 35.140 149.005 36.955 149.915 ;
        RECT 36.965 149.235 38.795 149.915 ;
        RECT 37.450 149.005 38.795 149.235 ;
        RECT 38.805 149.105 42.475 149.915 ;
        RECT 42.485 149.105 43.855 149.915 ;
        RECT 43.875 149.045 44.305 149.830 ;
        RECT 44.325 149.105 49.835 149.915 ;
        RECT 50.305 149.005 53.975 149.915 ;
        RECT 54.295 149.235 56.130 149.915 ;
        RECT 54.295 149.005 55.225 149.235 ;
        RECT 56.285 149.005 57.635 149.915 ;
        RECT 57.665 149.005 60.875 149.915 ;
        RECT 60.905 149.005 62.255 149.915 ;
        RECT 62.265 149.105 67.775 149.915 ;
        RECT 67.785 149.005 69.600 149.915 ;
        RECT 69.635 149.045 70.065 149.830 ;
        RECT 70.085 149.105 75.595 149.915 ;
        RECT 75.605 149.105 81.115 149.915 ;
        RECT 81.125 149.105 86.635 149.915 ;
        RECT 86.645 149.135 88.015 149.915 ;
        RECT 88.025 149.105 89.395 149.915 ;
      LAYER nwell ;
        RECT 17.910 145.885 89.590 148.715 ;
      LAYER pwell ;
        RECT 18.105 144.685 19.475 145.495 ;
        RECT 19.485 144.685 24.995 145.495 ;
        RECT 25.005 144.685 30.515 145.495 ;
        RECT 30.995 144.770 31.425 145.555 ;
        RECT 31.445 144.685 33.275 145.495 ;
        RECT 33.765 144.685 35.115 145.595 ;
        RECT 35.125 144.685 38.785 145.595 ;
        RECT 38.975 144.685 42.475 145.595 ;
        RECT 42.485 144.685 45.235 145.495 ;
        RECT 45.255 144.915 48.455 145.595 ;
        RECT 45.255 144.685 48.310 144.915 ;
        RECT 48.465 144.685 53.975 145.495 ;
        RECT 53.985 144.685 56.735 145.495 ;
        RECT 56.755 144.770 57.185 145.555 ;
        RECT 57.700 145.365 59.075 145.595 ;
        RECT 60.845 145.365 61.795 145.595 ;
        RECT 62.290 145.365 63.635 145.595 ;
        RECT 64.130 145.365 67.740 145.595 ;
        RECT 57.700 144.915 61.795 145.365 ;
        RECT 18.245 144.475 18.415 144.685 ;
        RECT 19.625 144.475 19.795 144.685 ;
        RECT 25.145 144.475 25.315 144.685 ;
        RECT 30.665 144.635 30.835 144.665 ;
        RECT 30.660 144.525 30.835 144.635 ;
        RECT 30.665 144.475 30.835 144.525 ;
        RECT 31.585 144.495 31.755 144.685 ;
        RECT 33.420 144.525 33.540 144.635 ;
        RECT 33.880 144.495 34.050 144.685 ;
        RECT 37.560 144.475 37.730 144.665 ;
        RECT 38.500 144.495 38.670 144.685 ;
        RECT 38.975 144.665 39.110 144.685 ;
        RECT 38.940 144.495 39.110 144.665 ;
        RECT 39.865 144.495 40.035 144.665 ;
        RECT 40.335 144.520 40.495 144.630 ;
        RECT 39.865 144.475 40.015 144.495 ;
        RECT 41.250 144.475 41.420 144.665 ;
        RECT 42.625 144.495 42.795 144.685 ;
        RECT 43.540 144.525 43.660 144.635 ;
        RECT 45.845 144.475 46.015 144.665 ;
        RECT 46.305 144.475 46.475 144.665 ;
        RECT 47.685 144.475 47.855 144.665 ;
        RECT 48.140 144.495 48.310 144.685 ;
        RECT 48.605 144.495 48.775 144.685 ;
        RECT 53.205 144.475 53.375 144.665 ;
        RECT 54.125 144.495 54.295 144.685 ;
        RECT 57.340 144.525 57.460 144.635 ;
        RECT 57.805 144.495 57.975 144.915 ;
        RECT 59.085 144.685 61.795 144.915 ;
        RECT 61.805 144.685 63.635 145.365 ;
        RECT 63.645 144.685 67.740 145.365 ;
        RECT 67.785 144.685 73.295 145.495 ;
        RECT 73.305 144.685 78.815 145.495 ;
        RECT 78.825 144.685 82.495 145.495 ;
        RECT 82.515 144.770 82.945 145.555 ;
        RECT 82.965 144.685 85.715 145.495 ;
        RECT 86.185 144.685 88.015 145.365 ;
        RECT 88.025 144.685 89.395 145.495 ;
        RECT 58.725 144.475 58.895 144.665 ;
        RECT 61.945 144.495 62.115 144.685 ;
        RECT 62.400 144.525 62.520 144.635 ;
        RECT 63.790 144.495 63.960 144.685 ;
        RECT 66.540 144.475 66.710 144.665 ;
        RECT 67.005 144.475 67.175 144.665 ;
        RECT 67.925 144.495 68.095 144.685 ;
        RECT 70.225 144.475 70.395 144.665 ;
        RECT 73.445 144.495 73.615 144.685 ;
        RECT 75.745 144.475 75.915 144.665 ;
        RECT 78.965 144.495 79.135 144.685 ;
        RECT 81.265 144.475 81.435 144.665 ;
        RECT 83.105 144.495 83.275 144.685 ;
        RECT 85.860 144.525 85.980 144.635 ;
        RECT 87.705 144.495 87.875 144.685 ;
        RECT 89.085 144.475 89.255 144.685 ;
        RECT 18.105 143.665 19.475 144.475 ;
        RECT 19.485 143.665 24.995 144.475 ;
        RECT 25.005 143.665 30.515 144.475 ;
        RECT 30.525 143.665 36.035 144.475 ;
        RECT 36.045 143.565 37.875 144.475 ;
        RECT 38.085 143.655 40.015 144.475 ;
        RECT 41.105 143.795 43.380 144.475 ;
        RECT 38.085 143.565 39.035 143.655 ;
        RECT 42.010 143.565 43.380 143.795 ;
        RECT 43.875 143.605 44.305 144.390 ;
        RECT 44.325 143.795 46.155 144.475 ;
        RECT 46.165 143.695 47.535 144.475 ;
        RECT 47.545 143.665 53.055 144.475 ;
        RECT 53.065 143.665 58.575 144.475 ;
        RECT 58.585 143.665 62.255 144.475 ;
        RECT 62.760 143.795 66.855 144.475 ;
        RECT 62.760 143.565 66.370 143.795 ;
        RECT 66.865 143.665 69.615 144.475 ;
        RECT 69.635 143.605 70.065 144.390 ;
        RECT 70.085 143.665 75.595 144.475 ;
        RECT 75.605 143.665 81.115 144.475 ;
        RECT 81.125 143.665 86.635 144.475 ;
        RECT 88.025 143.665 89.395 144.475 ;
      LAYER nwell ;
        RECT 17.910 140.445 89.590 143.275 ;
      LAYER pwell ;
        RECT 18.105 139.245 19.475 140.055 ;
        RECT 19.485 139.245 24.995 140.055 ;
        RECT 27.305 139.245 30.975 140.055 ;
        RECT 30.995 139.330 31.425 140.115 ;
        RECT 31.445 139.245 35.115 140.055 ;
        RECT 35.585 139.245 36.955 140.025 ;
        RECT 36.965 139.245 38.795 140.055 ;
        RECT 39.290 139.925 40.635 140.155 ;
        RECT 38.805 139.245 40.635 139.925 ;
        RECT 40.645 139.245 41.995 140.155 ;
        RECT 42.025 139.245 43.395 140.025 ;
        RECT 43.875 139.330 44.305 140.115 ;
        RECT 45.245 139.245 47.075 139.925 ;
        RECT 47.085 139.245 48.455 140.055 ;
        RECT 48.950 139.925 50.295 140.155 ;
        RECT 48.465 139.245 50.295 139.925 ;
        RECT 50.305 139.245 55.815 140.055 ;
        RECT 56.755 139.330 57.185 140.115 ;
        RECT 57.205 139.245 62.715 140.055 ;
        RECT 62.725 139.245 68.235 140.055 ;
        RECT 68.245 139.245 69.615 140.055 ;
        RECT 69.635 139.330 70.065 140.115 ;
        RECT 70.085 139.245 75.595 140.055 ;
        RECT 75.605 139.245 81.115 140.055 ;
        RECT 81.125 139.245 82.495 140.055 ;
        RECT 82.515 139.330 82.945 140.115 ;
        RECT 82.965 139.245 86.635 140.055 ;
        RECT 86.645 139.245 88.015 140.055 ;
        RECT 88.025 139.245 89.395 140.055 ;
        RECT 18.245 139.055 18.415 139.245 ;
        RECT 19.625 139.055 19.795 139.245 ;
        RECT 25.155 139.090 25.315 139.200 ;
        RECT 26.985 139.055 27.155 139.225 ;
        RECT 27.445 139.055 27.615 139.245 ;
        RECT 31.585 139.055 31.755 139.245 ;
        RECT 35.260 139.085 35.380 139.195 ;
        RECT 36.645 139.055 36.815 139.245 ;
        RECT 37.105 139.055 37.275 139.245 ;
        RECT 38.945 139.055 39.115 139.245 ;
        RECT 41.710 139.055 41.880 139.245 ;
        RECT 42.175 139.055 42.345 139.245 ;
        RECT 43.540 139.085 43.660 139.195 ;
        RECT 44.475 139.090 44.635 139.200 ;
        RECT 45.385 139.055 45.555 139.245 ;
        RECT 47.225 139.055 47.395 139.245 ;
        RECT 48.605 139.055 48.775 139.245 ;
        RECT 50.445 139.055 50.615 139.245 ;
        RECT 55.975 139.090 56.135 139.200 ;
        RECT 57.345 139.055 57.515 139.245 ;
        RECT 62.865 139.055 63.035 139.245 ;
        RECT 68.385 139.055 68.555 139.245 ;
        RECT 70.225 139.055 70.395 139.245 ;
        RECT 75.745 139.055 75.915 139.245 ;
        RECT 81.265 139.055 81.435 139.245 ;
        RECT 83.105 139.055 83.275 139.245 ;
        RECT 86.785 139.055 86.955 139.245 ;
        RECT 89.085 139.055 89.255 139.245 ;
      LAYER li1 ;
        RECT 18.100 209.775 89.400 209.945 ;
        RECT 18.185 209.025 19.395 209.775 ;
        RECT 18.185 208.485 18.705 209.025 ;
        RECT 19.625 208.955 19.835 209.775 ;
        RECT 20.005 208.975 20.335 209.605 ;
        RECT 18.875 208.315 19.395 208.855 ;
        RECT 20.005 208.375 20.255 208.975 ;
        RECT 20.505 208.955 20.735 209.775 ;
        RECT 21.035 209.225 21.205 209.605 ;
        RECT 21.420 209.395 21.750 209.775 ;
        RECT 21.035 209.055 21.750 209.225 ;
        RECT 20.425 208.535 20.755 208.785 ;
        RECT 20.945 208.505 21.300 208.875 ;
        RECT 21.580 208.865 21.750 209.055 ;
        RECT 21.920 209.030 22.175 209.605 ;
        RECT 21.580 208.535 21.835 208.865 ;
        RECT 18.185 207.225 19.395 208.315 ;
        RECT 19.625 207.225 19.835 208.365 ;
        RECT 20.005 207.395 20.335 208.375 ;
        RECT 20.505 207.225 20.735 208.365 ;
        RECT 21.580 208.325 21.750 208.535 ;
        RECT 21.035 208.155 21.750 208.325 ;
        RECT 22.005 208.300 22.175 209.030 ;
        RECT 22.350 208.935 22.610 209.775 ;
        RECT 22.790 208.935 23.050 209.775 ;
        RECT 23.225 209.030 23.480 209.605 ;
        RECT 23.650 209.395 23.980 209.775 ;
        RECT 24.195 209.225 24.365 209.605 ;
        RECT 23.650 209.055 24.365 209.225 ;
        RECT 21.035 207.395 21.205 208.155 ;
        RECT 21.420 207.225 21.750 207.985 ;
        RECT 21.920 207.395 22.175 208.300 ;
        RECT 22.350 207.225 22.610 208.375 ;
        RECT 22.790 207.225 23.050 208.375 ;
        RECT 23.225 208.300 23.395 209.030 ;
        RECT 23.650 208.865 23.820 209.055 ;
        RECT 24.630 208.935 24.890 209.775 ;
        RECT 25.065 209.030 25.320 209.605 ;
        RECT 25.490 209.395 25.820 209.775 ;
        RECT 26.035 209.225 26.205 209.605 ;
        RECT 26.630 209.265 26.870 209.775 ;
        RECT 27.050 209.265 27.330 209.595 ;
        RECT 27.560 209.265 27.775 209.775 ;
        RECT 25.490 209.055 26.205 209.225 ;
        RECT 23.565 208.535 23.820 208.865 ;
        RECT 23.650 208.325 23.820 208.535 ;
        RECT 24.100 208.505 24.455 208.875 ;
        RECT 23.225 207.395 23.480 208.300 ;
        RECT 23.650 208.155 24.365 208.325 ;
        RECT 23.650 207.225 23.980 207.985 ;
        RECT 24.195 207.395 24.365 208.155 ;
        RECT 24.630 207.225 24.890 208.375 ;
        RECT 25.065 208.300 25.235 209.030 ;
        RECT 25.490 208.865 25.660 209.055 ;
        RECT 25.405 208.535 25.660 208.865 ;
        RECT 25.490 208.325 25.660 208.535 ;
        RECT 25.940 208.505 26.295 208.875 ;
        RECT 26.525 208.535 26.880 209.095 ;
        RECT 27.050 208.365 27.220 209.265 ;
        RECT 27.390 208.535 27.655 209.095 ;
        RECT 27.945 209.035 28.560 209.605 ;
        RECT 28.875 209.395 30.045 209.605 ;
        RECT 28.875 209.375 29.205 209.395 ;
        RECT 27.905 208.365 28.075 208.865 ;
        RECT 25.065 207.395 25.320 208.300 ;
        RECT 25.490 208.155 26.205 208.325 ;
        RECT 25.490 207.225 25.820 207.985 ;
        RECT 26.035 207.395 26.205 208.155 ;
        RECT 26.650 208.195 28.075 208.365 ;
        RECT 26.650 208.020 27.040 208.195 ;
        RECT 27.525 207.225 27.855 208.025 ;
        RECT 28.245 208.015 28.560 209.035 ;
        RECT 28.765 208.955 29.625 209.205 ;
        RECT 29.795 209.145 30.045 209.395 ;
        RECT 30.215 209.315 30.385 209.775 ;
        RECT 30.555 209.145 30.895 209.605 ;
        RECT 29.795 208.975 30.895 209.145 ;
        RECT 31.065 209.050 31.355 209.775 ;
        RECT 31.635 209.395 32.805 209.605 ;
        RECT 31.635 209.375 31.965 209.395 ;
        RECT 31.525 208.955 32.385 209.205 ;
        RECT 32.555 209.145 32.805 209.395 ;
        RECT 32.975 209.315 33.145 209.775 ;
        RECT 33.315 209.145 33.655 209.605 ;
        RECT 32.555 208.975 33.655 209.145 ;
        RECT 34.025 209.145 34.355 209.505 ;
        RECT 34.985 209.315 35.235 209.775 ;
        RECT 35.405 209.315 35.955 209.605 ;
        RECT 34.025 208.955 35.415 209.145 ;
        RECT 28.765 208.365 29.045 208.955 ;
        RECT 29.215 208.535 29.965 208.785 ;
        RECT 30.135 208.535 30.895 208.785 ;
        RECT 28.765 208.195 30.465 208.365 ;
        RECT 28.025 207.395 28.560 208.015 ;
        RECT 28.870 207.225 29.125 208.025 ;
        RECT 29.295 207.395 29.625 208.195 ;
        RECT 29.795 207.225 29.965 208.025 ;
        RECT 30.135 207.395 30.465 208.195 ;
        RECT 30.635 207.225 30.895 208.365 ;
        RECT 31.065 207.225 31.355 208.390 ;
        RECT 31.525 208.365 31.805 208.955 ;
        RECT 35.245 208.865 35.415 208.955 ;
        RECT 31.975 208.535 32.725 208.785 ;
        RECT 32.895 208.535 33.655 208.785 ;
        RECT 33.825 208.535 34.515 208.785 ;
        RECT 34.745 208.535 35.075 208.785 ;
        RECT 35.245 208.535 35.535 208.865 ;
        RECT 31.525 208.195 33.225 208.365 ;
        RECT 31.630 207.225 31.885 208.025 ;
        RECT 32.055 207.395 32.385 208.195 ;
        RECT 32.555 207.225 32.725 208.025 ;
        RECT 32.895 207.395 33.225 208.195 ;
        RECT 33.395 207.225 33.655 208.365 ;
        RECT 33.825 208.095 34.140 208.535 ;
        RECT 35.245 208.285 35.415 208.535 ;
        RECT 34.475 208.115 35.415 208.285 ;
        RECT 34.025 207.225 34.305 207.895 ;
        RECT 34.475 207.565 34.775 208.115 ;
        RECT 35.705 207.945 35.955 209.315 ;
        RECT 36.125 208.975 36.415 209.775 ;
        RECT 36.670 209.275 37.165 209.605 ;
        RECT 34.985 207.225 35.315 207.945 ;
        RECT 35.505 207.395 35.955 207.945 ;
        RECT 36.125 207.225 36.415 208.365 ;
        RECT 36.585 207.785 36.825 209.095 ;
        RECT 36.995 208.365 37.165 209.275 ;
        RECT 37.385 208.535 37.735 209.500 ;
        RECT 37.915 208.535 38.215 209.505 ;
        RECT 38.395 208.535 38.675 209.505 ;
        RECT 38.855 208.975 39.125 209.775 ;
        RECT 39.295 209.055 39.635 209.565 ;
        RECT 39.890 209.225 40.220 209.605 ;
        RECT 40.390 209.395 41.575 209.565 ;
        RECT 41.835 209.305 42.005 209.775 ;
        RECT 39.890 209.055 40.435 209.225 ;
        RECT 38.870 208.535 39.200 208.785 ;
        RECT 38.870 208.365 39.185 208.535 ;
        RECT 36.995 208.195 39.185 208.365 ;
        RECT 36.590 207.225 36.925 207.605 ;
        RECT 37.095 207.395 37.345 208.195 ;
        RECT 37.565 207.225 37.895 207.945 ;
        RECT 38.080 207.395 38.330 208.195 ;
        RECT 38.795 207.225 39.125 208.025 ;
        RECT 39.375 207.655 39.635 209.055 ;
        RECT 39.805 208.535 40.065 208.885 ;
        RECT 40.265 208.415 40.435 209.055 ;
        RECT 40.805 209.125 41.190 209.215 ;
        RECT 42.175 209.125 42.505 209.590 ;
        RECT 40.805 208.955 42.505 209.125 ;
        RECT 42.675 208.955 42.845 209.775 ;
        RECT 43.015 209.125 43.345 209.595 ;
        RECT 43.515 209.295 43.685 209.775 ;
        RECT 43.015 208.955 43.775 209.125 ;
        RECT 43.945 209.050 44.235 209.775 ;
        RECT 45.415 209.295 45.715 209.775 ;
        RECT 45.885 209.125 46.145 209.580 ;
        RECT 46.315 209.295 46.575 209.775 ;
        RECT 46.755 209.125 47.015 209.580 ;
        RECT 47.185 209.295 47.435 209.775 ;
        RECT 47.615 209.125 47.875 209.580 ;
        RECT 48.045 209.295 48.295 209.775 ;
        RECT 48.475 209.125 48.735 209.580 ;
        RECT 48.905 209.295 49.150 209.775 ;
        RECT 49.320 209.125 49.595 209.580 ;
        RECT 49.765 209.295 50.010 209.775 ;
        RECT 50.180 209.125 50.440 209.580 ;
        RECT 50.610 209.295 50.870 209.775 ;
        RECT 51.040 209.125 51.300 209.580 ;
        RECT 51.470 209.295 51.730 209.775 ;
        RECT 51.900 209.125 52.160 209.580 ;
        RECT 52.330 209.215 52.590 209.775 ;
        RECT 45.415 209.095 52.160 209.125 ;
        RECT 40.605 208.585 40.950 208.785 ;
        RECT 41.120 208.585 41.510 208.785 ;
        RECT 40.265 208.365 41.050 208.415 ;
        RECT 39.295 207.395 39.635 207.655 ;
        RECT 39.970 208.190 41.050 208.365 ;
        RECT 39.970 207.395 40.300 208.190 ;
        RECT 40.470 207.225 40.710 208.010 ;
        RECT 40.880 207.985 41.050 208.190 ;
        RECT 41.220 208.155 41.510 208.585 ;
        RECT 41.700 208.575 42.185 208.785 ;
        RECT 42.355 208.575 42.795 208.785 ;
        RECT 42.965 208.575 43.295 208.785 ;
        RECT 41.700 208.155 42.005 208.575 ;
        RECT 42.965 208.405 43.135 208.575 ;
        RECT 42.175 208.235 43.135 208.405 ;
        RECT 42.175 207.985 42.345 208.235 ;
        RECT 40.880 207.815 42.345 207.985 ;
        RECT 41.270 207.395 42.025 207.815 ;
        RECT 42.515 207.225 42.845 208.065 ;
        RECT 43.465 207.985 43.775 208.955 ;
        RECT 45.385 208.955 52.160 209.095 ;
        RECT 45.385 208.925 46.580 208.955 ;
        RECT 43.015 207.815 43.775 207.985 ;
        RECT 43.015 207.395 43.265 207.815 ;
        RECT 43.435 207.225 43.775 207.645 ;
        RECT 43.945 207.225 44.235 208.390 ;
        RECT 45.415 208.365 46.580 208.925 ;
        RECT 52.760 208.785 53.010 209.595 ;
        RECT 53.190 209.250 53.450 209.775 ;
        RECT 53.620 208.785 53.870 209.595 ;
        RECT 54.050 209.265 54.355 209.775 ;
        RECT 54.545 209.265 54.785 209.775 ;
        RECT 54.955 209.265 55.245 209.605 ;
        RECT 55.475 209.265 55.790 209.775 ;
        RECT 46.750 208.535 53.870 208.785 ;
        RECT 54.040 208.535 54.355 209.095 ;
        RECT 54.590 208.755 54.785 209.095 ;
        RECT 54.585 208.585 54.785 208.755 ;
        RECT 54.590 208.535 54.785 208.585 ;
        RECT 45.415 208.140 52.160 208.365 ;
        RECT 45.415 207.225 45.685 207.970 ;
        RECT 45.855 207.400 46.145 208.140 ;
        RECT 46.755 208.125 52.160 208.140 ;
        RECT 46.315 207.230 46.570 207.955 ;
        RECT 46.755 207.400 47.015 208.125 ;
        RECT 47.185 207.230 47.430 207.955 ;
        RECT 47.615 207.400 47.875 208.125 ;
        RECT 48.045 207.230 48.290 207.955 ;
        RECT 48.475 207.400 48.735 208.125 ;
        RECT 48.905 207.230 49.150 207.955 ;
        RECT 49.320 207.400 49.580 208.125 ;
        RECT 49.750 207.230 50.010 207.955 ;
        RECT 50.180 207.400 50.440 208.125 ;
        RECT 50.610 207.230 50.870 207.955 ;
        RECT 51.040 207.400 51.300 208.125 ;
        RECT 51.470 207.230 51.730 207.955 ;
        RECT 51.900 207.400 52.160 208.125 ;
        RECT 52.330 207.230 52.590 208.025 ;
        RECT 52.760 207.400 53.010 208.535 ;
        RECT 46.315 207.225 52.590 207.230 ;
        RECT 53.190 207.225 53.450 208.035 ;
        RECT 53.625 207.395 53.870 208.535 ;
        RECT 54.955 208.365 55.135 209.265 ;
        RECT 55.960 209.205 56.130 209.475 ;
        RECT 56.300 209.375 56.630 209.775 ;
        RECT 55.305 208.535 55.715 209.095 ;
        RECT 55.960 209.035 56.655 209.205 ;
        RECT 56.825 209.050 57.115 209.775 ;
        RECT 57.615 209.375 57.945 209.775 ;
        RECT 58.115 209.205 58.445 209.545 ;
        RECT 59.495 209.375 59.825 209.775 ;
        RECT 55.885 208.365 56.055 208.865 ;
        RECT 54.595 208.195 56.055 208.365 ;
        RECT 54.050 207.225 54.345 208.035 ;
        RECT 54.595 208.020 54.955 208.195 ;
        RECT 56.225 208.025 56.655 209.035 ;
        RECT 57.460 209.035 59.825 209.205 ;
        RECT 59.995 209.050 60.325 209.560 ;
        RECT 60.595 209.295 60.895 209.775 ;
        RECT 61.065 209.125 61.325 209.580 ;
        RECT 61.495 209.295 61.755 209.775 ;
        RECT 61.935 209.125 62.195 209.580 ;
        RECT 62.365 209.295 62.615 209.775 ;
        RECT 62.795 209.125 63.055 209.580 ;
        RECT 63.225 209.295 63.475 209.775 ;
        RECT 63.655 209.125 63.915 209.580 ;
        RECT 64.085 209.295 64.330 209.775 ;
        RECT 64.500 209.125 64.775 209.580 ;
        RECT 64.945 209.295 65.190 209.775 ;
        RECT 65.360 209.125 65.620 209.580 ;
        RECT 65.790 209.295 66.050 209.775 ;
        RECT 66.220 209.125 66.480 209.580 ;
        RECT 66.650 209.295 66.910 209.775 ;
        RECT 67.080 209.125 67.340 209.580 ;
        RECT 67.510 209.215 67.770 209.775 ;
        RECT 55.540 207.225 55.710 208.025 ;
        RECT 55.880 207.855 56.655 208.025 ;
        RECT 55.880 207.395 56.210 207.855 ;
        RECT 56.380 207.225 56.550 207.685 ;
        RECT 56.825 207.225 57.115 208.390 ;
        RECT 57.460 208.035 57.630 209.035 ;
        RECT 59.655 208.865 59.825 209.035 ;
        RECT 57.800 208.205 58.045 208.865 ;
        RECT 58.260 208.205 58.525 208.865 ;
        RECT 58.720 208.205 59.005 208.865 ;
        RECT 59.180 208.535 59.485 208.865 ;
        RECT 59.655 208.535 59.965 208.865 ;
        RECT 59.180 208.205 59.395 208.535 ;
        RECT 60.135 208.415 60.325 209.050 ;
        RECT 57.460 207.865 57.915 208.035 ;
        RECT 57.585 207.435 57.915 207.865 ;
        RECT 58.095 207.865 59.385 208.035 ;
        RECT 58.095 207.445 58.345 207.865 ;
        RECT 58.575 207.225 58.905 207.695 ;
        RECT 59.135 207.445 59.385 207.865 ;
        RECT 59.575 207.225 59.825 208.365 ;
        RECT 60.105 208.285 60.325 208.415 ;
        RECT 59.995 207.435 60.325 208.285 ;
        RECT 60.595 208.955 67.340 209.125 ;
        RECT 60.595 208.365 61.760 208.955 ;
        RECT 67.940 208.785 68.190 209.595 ;
        RECT 68.370 209.250 68.630 209.775 ;
        RECT 68.800 208.785 69.050 209.595 ;
        RECT 69.230 209.265 69.535 209.775 ;
        RECT 61.930 208.535 69.050 208.785 ;
        RECT 69.220 208.535 69.535 209.095 ;
        RECT 69.705 209.050 69.995 209.775 ;
        RECT 70.175 209.045 70.475 209.775 ;
        RECT 70.655 208.865 70.885 209.485 ;
        RECT 71.085 209.215 71.310 209.595 ;
        RECT 71.480 209.385 71.810 209.775 ;
        RECT 72.005 209.265 72.310 209.775 ;
        RECT 71.085 209.035 71.415 209.215 ;
        RECT 70.180 208.535 70.475 208.865 ;
        RECT 70.655 208.535 71.070 208.865 ;
        RECT 60.595 208.140 67.340 208.365 ;
        RECT 60.595 207.225 60.865 207.970 ;
        RECT 61.035 207.400 61.325 208.140 ;
        RECT 61.935 208.125 67.340 208.140 ;
        RECT 61.495 207.230 61.750 207.955 ;
        RECT 61.935 207.400 62.195 208.125 ;
        RECT 62.365 207.230 62.610 207.955 ;
        RECT 62.795 207.400 63.055 208.125 ;
        RECT 63.225 207.230 63.470 207.955 ;
        RECT 63.655 207.400 63.915 208.125 ;
        RECT 64.085 207.230 64.330 207.955 ;
        RECT 64.500 207.400 64.760 208.125 ;
        RECT 64.930 207.230 65.190 207.955 ;
        RECT 65.360 207.400 65.620 208.125 ;
        RECT 65.790 207.230 66.050 207.955 ;
        RECT 66.220 207.400 66.480 208.125 ;
        RECT 66.650 207.230 66.910 207.955 ;
        RECT 67.080 207.400 67.340 208.125 ;
        RECT 67.510 207.230 67.770 208.025 ;
        RECT 67.940 207.400 68.190 208.535 ;
        RECT 61.495 207.225 67.770 207.230 ;
        RECT 68.370 207.225 68.630 208.035 ;
        RECT 68.805 207.395 69.050 208.535 ;
        RECT 69.230 207.225 69.525 208.035 ;
        RECT 69.705 207.225 69.995 208.390 ;
        RECT 71.240 208.365 71.415 209.035 ;
        RECT 71.585 208.535 71.825 209.185 ;
        RECT 72.005 208.535 72.320 209.095 ;
        RECT 72.490 208.785 72.740 209.595 ;
        RECT 72.910 209.250 73.170 209.775 ;
        RECT 73.350 208.785 73.600 209.595 ;
        RECT 73.770 209.215 74.030 209.775 ;
        RECT 74.200 209.125 74.460 209.580 ;
        RECT 74.630 209.295 74.890 209.775 ;
        RECT 75.060 209.125 75.320 209.580 ;
        RECT 75.490 209.295 75.750 209.775 ;
        RECT 75.920 209.125 76.180 209.580 ;
        RECT 76.350 209.295 76.595 209.775 ;
        RECT 76.765 209.125 77.040 209.580 ;
        RECT 77.210 209.295 77.455 209.775 ;
        RECT 77.625 209.125 77.885 209.580 ;
        RECT 78.065 209.295 78.315 209.775 ;
        RECT 78.485 209.125 78.745 209.580 ;
        RECT 78.925 209.295 79.175 209.775 ;
        RECT 79.345 209.125 79.605 209.580 ;
        RECT 79.785 209.295 80.045 209.775 ;
        RECT 80.215 209.125 80.475 209.580 ;
        RECT 80.645 209.295 80.945 209.775 ;
        RECT 74.200 208.955 80.945 209.125 ;
        RECT 81.245 208.955 81.475 209.775 ;
        RECT 81.645 208.975 81.975 209.605 ;
        RECT 72.490 208.535 79.610 208.785 ;
        RECT 70.175 208.005 71.070 208.335 ;
        RECT 71.240 208.175 71.825 208.365 ;
        RECT 70.175 207.835 71.380 208.005 ;
        RECT 70.175 207.405 70.505 207.835 ;
        RECT 70.685 207.225 70.880 207.665 ;
        RECT 71.050 207.405 71.380 207.835 ;
        RECT 71.550 207.405 71.825 208.175 ;
        RECT 72.015 207.225 72.310 208.035 ;
        RECT 72.490 207.395 72.735 208.535 ;
        RECT 72.910 207.225 73.170 208.035 ;
        RECT 73.350 207.400 73.600 208.535 ;
        RECT 79.780 208.415 80.945 208.955 ;
        RECT 81.225 208.535 81.555 208.785 ;
        RECT 79.780 208.365 80.975 208.415 ;
        RECT 81.725 208.375 81.975 208.975 ;
        RECT 82.145 208.955 82.355 209.775 ;
        RECT 82.585 209.050 82.875 209.775 ;
        RECT 74.200 208.245 80.975 208.365 ;
        RECT 74.200 208.140 80.945 208.245 ;
        RECT 74.200 208.125 79.605 208.140 ;
        RECT 73.770 207.230 74.030 208.025 ;
        RECT 74.200 207.400 74.460 208.125 ;
        RECT 74.630 207.230 74.890 207.955 ;
        RECT 75.060 207.400 75.320 208.125 ;
        RECT 75.490 207.230 75.750 207.955 ;
        RECT 75.920 207.400 76.180 208.125 ;
        RECT 76.350 207.230 76.610 207.955 ;
        RECT 76.780 207.400 77.040 208.125 ;
        RECT 77.210 207.230 77.455 207.955 ;
        RECT 77.625 207.400 77.885 208.125 ;
        RECT 78.070 207.230 78.315 207.955 ;
        RECT 78.485 207.400 78.745 208.125 ;
        RECT 78.930 207.230 79.175 207.955 ;
        RECT 79.345 207.400 79.605 208.125 ;
        RECT 79.790 207.230 80.045 207.955 ;
        RECT 80.215 207.400 80.505 208.140 ;
        RECT 73.770 207.225 80.045 207.230 ;
        RECT 80.675 207.225 80.945 207.970 ;
        RECT 81.245 207.225 81.475 208.365 ;
        RECT 81.645 207.395 81.975 208.375 ;
        RECT 82.145 207.225 82.355 208.365 ;
        RECT 82.585 207.225 82.875 208.390 ;
        RECT 83.065 208.195 83.295 209.535 ;
        RECT 83.475 208.695 83.705 209.595 ;
        RECT 83.905 208.995 84.150 209.775 ;
        RECT 84.320 209.235 84.750 209.595 ;
        RECT 85.330 209.405 86.060 209.775 ;
        RECT 84.320 209.045 86.060 209.235 ;
        RECT 84.320 208.815 84.540 209.045 ;
        RECT 83.475 208.015 83.815 208.695 ;
        RECT 83.065 207.815 83.815 208.015 ;
        RECT 83.995 208.515 84.540 208.815 ;
        RECT 83.065 207.425 83.305 207.815 ;
        RECT 83.475 207.225 83.825 207.635 ;
        RECT 83.995 207.405 84.325 208.515 ;
        RECT 84.710 208.245 85.135 208.865 ;
        RECT 85.330 208.245 85.590 208.865 ;
        RECT 85.800 208.535 86.060 209.045 ;
        RECT 84.495 207.875 85.520 208.075 ;
        RECT 84.495 207.405 84.675 207.875 ;
        RECT 84.845 207.225 85.175 207.705 ;
        RECT 85.350 207.405 85.520 207.875 ;
        RECT 85.785 207.225 86.070 208.365 ;
        RECT 86.260 207.405 86.540 209.595 ;
        RECT 86.725 209.100 86.985 209.605 ;
        RECT 87.165 209.395 87.495 209.775 ;
        RECT 87.675 209.225 87.845 209.605 ;
        RECT 86.725 208.300 86.905 209.100 ;
        RECT 87.180 209.055 87.845 209.225 ;
        RECT 87.180 208.800 87.350 209.055 ;
        RECT 88.105 209.025 89.315 209.775 ;
        RECT 87.075 208.470 87.350 208.800 ;
        RECT 87.575 208.505 87.915 208.875 ;
        RECT 87.180 208.325 87.350 208.470 ;
        RECT 86.725 207.395 86.995 208.300 ;
        RECT 87.180 208.155 87.855 208.325 ;
        RECT 87.165 207.225 87.495 207.985 ;
        RECT 87.675 207.395 87.855 208.155 ;
        RECT 88.105 208.315 88.625 208.855 ;
        RECT 88.795 208.485 89.315 209.025 ;
        RECT 88.105 207.225 89.315 208.315 ;
        RECT 18.100 207.055 89.400 207.225 ;
        RECT 18.185 205.965 19.395 207.055 ;
        RECT 18.185 205.255 18.705 205.795 ;
        RECT 18.875 205.425 19.395 205.965 ;
        RECT 20.485 206.335 20.945 206.885 ;
        RECT 21.135 206.335 21.465 207.055 ;
        RECT 18.185 204.505 19.395 205.255 ;
        RECT 20.485 204.965 20.735 206.335 ;
        RECT 21.665 206.165 21.965 206.715 ;
        RECT 22.135 206.385 22.415 207.055 ;
        RECT 21.025 205.995 21.965 206.165 ;
        RECT 21.025 205.745 21.195 205.995 ;
        RECT 22.335 205.745 22.600 206.105 ;
        RECT 22.790 205.905 23.050 207.055 ;
        RECT 23.225 205.980 23.480 206.885 ;
        RECT 23.650 206.295 23.980 207.055 ;
        RECT 24.195 206.125 24.365 206.885 ;
        RECT 24.825 206.385 25.105 207.055 ;
        RECT 20.905 205.415 21.195 205.745 ;
        RECT 21.365 205.495 21.705 205.745 ;
        RECT 21.925 205.495 22.600 205.745 ;
        RECT 21.025 205.325 21.195 205.415 ;
        RECT 21.025 205.135 22.415 205.325 ;
        RECT 20.485 204.675 21.045 204.965 ;
        RECT 21.215 204.505 21.465 204.965 ;
        RECT 22.085 204.775 22.415 205.135 ;
        RECT 22.790 204.505 23.050 205.345 ;
        RECT 23.225 205.250 23.395 205.980 ;
        RECT 23.650 205.955 24.365 206.125 ;
        RECT 25.275 206.165 25.575 206.715 ;
        RECT 25.775 206.335 26.105 207.055 ;
        RECT 26.295 206.335 26.755 206.885 ;
        RECT 23.650 205.745 23.820 205.955 ;
        RECT 23.565 205.415 23.820 205.745 ;
        RECT 23.225 204.675 23.480 205.250 ;
        RECT 23.650 205.225 23.820 205.415 ;
        RECT 24.100 205.405 24.455 205.775 ;
        RECT 24.640 205.745 24.905 206.105 ;
        RECT 25.275 205.995 26.215 206.165 ;
        RECT 26.045 205.745 26.215 205.995 ;
        RECT 24.640 205.495 25.315 205.745 ;
        RECT 25.535 205.495 25.875 205.745 ;
        RECT 26.045 205.415 26.335 205.745 ;
        RECT 26.045 205.325 26.215 205.415 ;
        RECT 23.650 205.055 24.365 205.225 ;
        RECT 23.650 204.505 23.980 204.885 ;
        RECT 24.195 204.675 24.365 205.055 ;
        RECT 24.825 205.135 26.215 205.325 ;
        RECT 24.825 204.775 25.155 205.135 ;
        RECT 26.505 204.965 26.755 206.335 ;
        RECT 26.925 205.995 27.240 207.055 ;
        RECT 27.870 206.550 28.485 207.055 ;
        RECT 26.985 205.165 27.250 205.745 ;
        RECT 27.420 205.665 27.695 206.325 ;
        RECT 27.890 206.015 28.125 206.380 ;
        RECT 28.295 206.375 28.485 206.550 ;
        RECT 28.655 206.545 29.130 206.885 ;
        RECT 28.295 206.185 28.625 206.375 ;
        RECT 28.850 206.015 29.040 206.310 ;
        RECT 29.300 206.210 29.515 207.055 ;
        RECT 29.715 206.215 30.000 206.885 ;
        RECT 27.890 205.845 29.660 206.015 ;
        RECT 27.420 205.435 28.255 205.665 ;
        RECT 25.775 204.505 26.025 204.965 ;
        RECT 26.195 204.675 26.755 204.965 ;
        RECT 26.925 204.505 27.195 204.995 ;
        RECT 27.420 204.725 27.695 205.435 ;
        RECT 28.425 204.990 28.680 205.845 ;
        RECT 27.895 204.725 28.680 204.990 ;
        RECT 28.850 205.185 29.260 205.665 ;
        RECT 29.430 205.415 29.660 205.845 ;
        RECT 29.830 205.865 30.000 206.215 ;
        RECT 30.170 206.045 30.435 207.055 ;
        RECT 31.065 205.890 31.355 207.055 ;
        RECT 31.990 205.910 32.285 207.055 ;
        RECT 29.830 205.345 30.435 205.865 ;
        RECT 28.850 204.725 29.060 205.185 ;
        RECT 29.830 205.135 30.000 205.345 ;
        RECT 29.250 204.505 29.580 205.000 ;
        RECT 29.755 204.675 30.000 205.135 ;
        RECT 30.170 204.505 30.435 205.165 ;
        RECT 31.065 204.505 31.355 205.230 ;
        RECT 31.990 204.505 32.285 205.325 ;
        RECT 32.455 205.055 32.685 206.755 ;
        RECT 32.900 206.250 33.155 207.055 ;
        RECT 33.355 206.440 33.685 206.885 ;
        RECT 33.855 206.610 34.130 207.055 ;
        RECT 34.365 206.440 34.695 206.885 ;
        RECT 33.355 206.260 34.695 206.440 ;
        RECT 35.155 206.080 35.485 206.745 ;
        RECT 35.685 206.255 36.015 207.055 ;
        RECT 32.900 205.910 35.485 206.080 ;
        RECT 36.190 205.915 36.525 206.885 ;
        RECT 36.695 206.255 37.025 207.055 ;
        RECT 37.425 206.085 37.675 206.885 ;
        RECT 37.860 206.335 38.190 207.055 ;
        RECT 38.410 206.085 38.660 206.885 ;
        RECT 38.835 206.675 39.165 207.055 ;
        RECT 36.705 205.915 38.760 206.085 ;
        RECT 32.900 205.295 33.210 205.910 ;
        RECT 36.190 205.695 36.365 205.915 ;
        RECT 36.705 205.735 36.930 205.915 ;
        RECT 33.380 205.465 33.710 205.695 ;
        RECT 33.880 205.465 34.350 205.695 ;
        RECT 34.520 205.525 34.975 205.695 ;
        RECT 34.520 205.465 34.970 205.525 ;
        RECT 35.160 205.465 35.495 205.695 ;
        RECT 36.185 205.525 36.365 205.695 ;
        RECT 32.900 205.115 35.485 205.295 ;
        RECT 32.455 204.675 32.675 205.055 ;
        RECT 32.845 204.505 33.695 204.865 ;
        RECT 34.175 204.695 34.505 205.115 ;
        RECT 34.710 204.505 34.985 204.945 ;
        RECT 35.155 204.695 35.485 205.115 ;
        RECT 35.675 204.505 36.005 205.230 ;
        RECT 36.190 205.225 36.365 205.525 ;
        RECT 36.535 205.495 36.930 205.735 ;
        RECT 36.190 204.760 36.525 205.225 ;
        RECT 36.195 204.715 36.525 204.760 ;
        RECT 36.695 204.505 36.930 205.310 ;
        RECT 37.100 204.835 37.360 205.745 ;
        RECT 37.670 205.725 37.840 205.745 ;
        RECT 37.540 204.835 37.840 205.725 ;
        RECT 38.015 204.840 38.370 205.745 ;
        RECT 38.590 205.005 38.760 205.915 ;
        RECT 38.930 205.175 39.135 206.495 ;
        RECT 39.435 206.310 39.705 207.055 ;
        RECT 40.335 207.050 46.610 207.055 ;
        RECT 39.875 206.140 40.165 206.880 ;
        RECT 40.335 206.325 40.590 207.050 ;
        RECT 40.775 206.155 41.035 206.880 ;
        RECT 41.205 206.325 41.450 207.050 ;
        RECT 41.635 206.155 41.895 206.880 ;
        RECT 42.065 206.325 42.310 207.050 ;
        RECT 42.495 206.155 42.755 206.880 ;
        RECT 42.925 206.325 43.170 207.050 ;
        RECT 43.340 206.155 43.600 206.880 ;
        RECT 43.770 206.325 44.030 207.050 ;
        RECT 44.200 206.155 44.460 206.880 ;
        RECT 44.630 206.325 44.890 207.050 ;
        RECT 45.060 206.155 45.320 206.880 ;
        RECT 45.490 206.325 45.750 207.050 ;
        RECT 45.920 206.155 46.180 206.880 ;
        RECT 46.350 206.255 46.610 207.050 ;
        RECT 40.775 206.140 46.180 206.155 ;
        RECT 39.435 205.915 46.180 206.140 ;
        RECT 39.435 205.325 40.600 205.915 ;
        RECT 46.780 205.745 47.030 206.880 ;
        RECT 47.210 206.245 47.470 207.055 ;
        RECT 47.645 205.745 47.890 206.885 ;
        RECT 48.070 206.245 48.365 207.055 ;
        RECT 48.635 206.045 48.805 206.885 ;
        RECT 48.975 206.715 50.145 206.885 ;
        RECT 48.975 206.215 49.305 206.715 ;
        RECT 49.815 206.675 50.145 206.715 ;
        RECT 50.335 206.635 50.690 207.055 ;
        RECT 49.475 206.455 49.705 206.545 ;
        RECT 50.860 206.455 51.110 206.885 ;
        RECT 49.475 206.215 51.110 206.455 ;
        RECT 51.280 206.295 51.610 207.055 ;
        RECT 51.780 206.215 52.035 206.885 ;
        RECT 48.635 205.875 51.695 206.045 ;
        RECT 40.770 205.495 47.890 205.745 ;
        RECT 39.435 205.155 46.180 205.325 ;
        RECT 38.590 204.675 39.085 205.005 ;
        RECT 39.435 204.505 39.735 204.985 ;
        RECT 39.905 204.700 40.165 205.155 ;
        RECT 40.335 204.505 40.595 204.985 ;
        RECT 40.775 204.700 41.035 205.155 ;
        RECT 41.205 204.505 41.455 204.985 ;
        RECT 41.635 204.700 41.895 205.155 ;
        RECT 42.065 204.505 42.315 204.985 ;
        RECT 42.495 204.700 42.755 205.155 ;
        RECT 42.925 204.505 43.170 204.985 ;
        RECT 43.340 204.700 43.615 205.155 ;
        RECT 43.785 204.505 44.030 204.985 ;
        RECT 44.200 204.700 44.460 205.155 ;
        RECT 44.630 204.505 44.890 204.985 ;
        RECT 45.060 204.700 45.320 205.155 ;
        RECT 45.490 204.505 45.750 204.985 ;
        RECT 45.920 204.700 46.180 205.155 ;
        RECT 46.350 204.505 46.610 205.065 ;
        RECT 46.780 204.685 47.030 205.495 ;
        RECT 47.210 204.505 47.470 205.030 ;
        RECT 47.640 204.685 47.890 205.495 ;
        RECT 48.060 205.185 48.375 205.745 ;
        RECT 48.545 205.495 48.900 205.705 ;
        RECT 49.070 205.495 49.515 205.695 ;
        RECT 49.685 205.495 50.160 205.695 ;
        RECT 48.635 205.155 49.700 205.325 ;
        RECT 48.070 204.505 48.375 205.015 ;
        RECT 48.635 204.675 48.805 205.155 ;
        RECT 48.975 204.505 49.305 204.985 ;
        RECT 49.530 204.925 49.700 205.155 ;
        RECT 49.880 205.095 50.160 205.495 ;
        RECT 50.430 205.495 50.760 205.695 ;
        RECT 50.930 205.495 51.295 205.695 ;
        RECT 50.430 205.095 50.715 205.495 ;
        RECT 51.525 205.325 51.695 205.875 ;
        RECT 50.895 205.155 51.695 205.325 ;
        RECT 50.895 204.925 51.065 205.155 ;
        RECT 51.865 205.085 52.035 206.215 ;
        RECT 52.205 205.865 52.375 207.055 ;
        RECT 52.695 206.080 53.025 206.745 ;
        RECT 53.485 206.440 53.815 206.885 ;
        RECT 54.050 206.610 54.325 207.055 ;
        RECT 54.495 206.440 54.825 206.885 ;
        RECT 53.485 206.260 54.825 206.440 ;
        RECT 55.025 206.250 55.280 207.055 ;
        RECT 52.695 205.910 55.280 206.080 ;
        RECT 52.685 205.465 53.020 205.695 ;
        RECT 53.205 205.525 53.660 205.695 ;
        RECT 53.210 205.465 53.660 205.525 ;
        RECT 53.830 205.465 54.300 205.695 ;
        RECT 54.470 205.465 54.800 205.695 ;
        RECT 51.850 205.015 52.035 205.085 ;
        RECT 51.825 205.005 52.035 205.015 ;
        RECT 49.530 204.675 51.065 204.925 ;
        RECT 51.235 204.505 51.565 204.985 ;
        RECT 51.780 204.675 52.035 205.005 ;
        RECT 52.205 204.505 52.375 205.400 ;
        RECT 54.970 205.295 55.280 205.910 ;
        RECT 52.695 205.115 55.280 205.295 ;
        RECT 52.695 204.695 53.025 205.115 ;
        RECT 53.195 204.505 53.470 204.945 ;
        RECT 53.675 204.695 54.005 205.115 ;
        RECT 55.495 205.055 55.725 206.755 ;
        RECT 55.895 205.910 56.190 207.055 ;
        RECT 56.825 205.890 57.115 207.055 ;
        RECT 57.285 206.085 57.595 206.885 ;
        RECT 57.765 206.255 58.075 207.055 ;
        RECT 58.245 206.425 58.505 206.885 ;
        RECT 58.675 206.595 58.930 207.055 ;
        RECT 59.105 206.425 59.365 206.885 ;
        RECT 58.245 206.255 59.365 206.425 ;
        RECT 57.285 205.915 58.315 206.085 ;
        RECT 54.485 204.505 55.335 204.865 ;
        RECT 55.505 204.675 55.725 205.055 ;
        RECT 55.895 204.505 56.190 205.325 ;
        RECT 56.825 204.505 57.115 205.230 ;
        RECT 57.285 205.005 57.455 205.915 ;
        RECT 57.625 205.175 57.975 205.745 ;
        RECT 58.145 205.665 58.315 205.915 ;
        RECT 59.105 206.005 59.365 206.255 ;
        RECT 59.535 206.185 59.820 207.055 ;
        RECT 60.045 206.460 60.480 206.885 ;
        RECT 60.650 206.630 61.035 207.055 ;
        RECT 60.045 206.290 61.035 206.460 ;
        RECT 59.105 205.835 59.860 206.005 ;
        RECT 58.145 205.495 59.285 205.665 ;
        RECT 59.455 205.325 59.860 205.835 ;
        RECT 60.045 205.415 60.530 206.120 ;
        RECT 60.700 205.745 61.035 206.290 ;
        RECT 61.205 206.095 61.630 206.885 ;
        RECT 61.800 206.460 62.075 206.885 ;
        RECT 62.245 206.630 62.630 207.055 ;
        RECT 61.800 206.265 62.630 206.460 ;
        RECT 61.205 205.915 62.110 206.095 ;
        RECT 60.700 205.415 61.110 205.745 ;
        RECT 61.280 205.415 62.110 205.915 ;
        RECT 62.280 205.745 62.630 206.265 ;
        RECT 62.800 206.095 63.045 206.885 ;
        RECT 63.235 206.460 63.490 206.885 ;
        RECT 63.660 206.630 64.045 207.055 ;
        RECT 63.235 206.265 64.045 206.460 ;
        RECT 62.800 205.915 63.525 206.095 ;
        RECT 62.280 205.415 62.705 205.745 ;
        RECT 62.875 205.415 63.525 205.915 ;
        RECT 63.695 205.745 64.045 206.265 ;
        RECT 64.215 205.915 64.475 206.885 ;
        RECT 64.655 206.245 64.950 207.055 ;
        RECT 63.695 205.415 64.120 205.745 ;
        RECT 58.210 205.155 59.860 205.325 ;
        RECT 60.700 205.245 61.035 205.415 ;
        RECT 61.280 205.245 61.630 205.415 ;
        RECT 62.280 205.245 62.630 205.415 ;
        RECT 62.875 205.245 63.045 205.415 ;
        RECT 63.695 205.245 64.045 205.415 ;
        RECT 64.290 205.245 64.475 205.915 ;
        RECT 65.130 205.745 65.375 206.885 ;
        RECT 65.550 206.245 65.810 207.055 ;
        RECT 66.410 207.050 72.685 207.055 ;
        RECT 65.990 205.745 66.240 206.880 ;
        RECT 66.410 206.255 66.670 207.050 ;
        RECT 66.840 206.155 67.100 206.880 ;
        RECT 67.270 206.325 67.530 207.050 ;
        RECT 67.700 206.155 67.960 206.880 ;
        RECT 68.130 206.325 68.390 207.050 ;
        RECT 68.560 206.155 68.820 206.880 ;
        RECT 68.990 206.325 69.250 207.050 ;
        RECT 69.420 206.155 69.680 206.880 ;
        RECT 69.850 206.325 70.095 207.050 ;
        RECT 70.265 206.155 70.525 206.880 ;
        RECT 70.710 206.325 70.955 207.050 ;
        RECT 71.125 206.155 71.385 206.880 ;
        RECT 71.570 206.325 71.815 207.050 ;
        RECT 71.985 206.155 72.245 206.880 ;
        RECT 72.430 206.325 72.685 207.050 ;
        RECT 66.840 206.140 72.245 206.155 ;
        RECT 72.855 206.140 73.145 206.880 ;
        RECT 73.315 206.310 73.585 207.055 ;
        RECT 73.865 206.465 74.105 206.855 ;
        RECT 74.275 206.645 74.625 207.055 ;
        RECT 73.865 206.265 74.615 206.465 ;
        RECT 66.840 205.915 73.585 206.140 ;
        RECT 57.285 204.675 57.585 205.005 ;
        RECT 57.755 204.505 58.030 204.985 ;
        RECT 58.210 204.765 58.505 205.155 ;
        RECT 58.675 204.505 58.930 204.985 ;
        RECT 59.105 204.765 59.365 205.155 ;
        RECT 60.045 205.075 61.035 205.245 ;
        RECT 59.535 204.505 59.815 204.985 ;
        RECT 60.045 204.675 60.480 205.075 ;
        RECT 60.650 204.505 61.035 204.905 ;
        RECT 61.205 204.675 61.630 205.245 ;
        RECT 61.820 205.075 62.630 205.245 ;
        RECT 61.820 204.675 62.075 205.075 ;
        RECT 62.245 204.505 62.630 204.905 ;
        RECT 62.800 204.675 63.045 205.245 ;
        RECT 63.235 205.075 64.045 205.245 ;
        RECT 63.235 204.675 63.490 205.075 ;
        RECT 63.660 204.505 64.045 204.905 ;
        RECT 64.215 204.675 64.475 205.245 ;
        RECT 64.645 205.185 64.960 205.745 ;
        RECT 65.130 205.495 72.250 205.745 ;
        RECT 64.645 204.505 64.950 205.015 ;
        RECT 65.130 204.685 65.380 205.495 ;
        RECT 65.550 204.505 65.810 205.030 ;
        RECT 65.990 204.685 66.240 205.495 ;
        RECT 72.420 205.325 73.585 205.915 ;
        RECT 66.840 205.155 73.585 205.325 ;
        RECT 66.410 204.505 66.670 205.065 ;
        RECT 66.840 204.700 67.100 205.155 ;
        RECT 67.270 204.505 67.530 204.985 ;
        RECT 67.700 204.700 67.960 205.155 ;
        RECT 68.130 204.505 68.390 204.985 ;
        RECT 68.560 204.700 68.820 205.155 ;
        RECT 68.990 204.505 69.235 204.985 ;
        RECT 69.405 204.700 69.680 205.155 ;
        RECT 69.850 204.505 70.095 204.985 ;
        RECT 70.265 204.700 70.525 205.155 ;
        RECT 70.705 204.505 70.955 204.985 ;
        RECT 71.125 204.700 71.385 205.155 ;
        RECT 71.565 204.505 71.815 204.985 ;
        RECT 71.985 204.700 72.245 205.155 ;
        RECT 72.425 204.505 72.685 204.985 ;
        RECT 72.855 204.700 73.115 205.155 ;
        RECT 73.285 204.505 73.585 204.985 ;
        RECT 73.865 204.745 74.095 206.085 ;
        RECT 74.275 205.585 74.615 206.265 ;
        RECT 74.795 205.765 75.125 206.875 ;
        RECT 75.295 206.405 75.475 206.875 ;
        RECT 75.645 206.575 75.975 207.055 ;
        RECT 76.150 206.405 76.320 206.875 ;
        RECT 75.295 206.205 76.320 206.405 ;
        RECT 74.275 204.685 74.505 205.585 ;
        RECT 74.795 205.465 75.340 205.765 ;
        RECT 74.705 204.505 74.950 205.285 ;
        RECT 75.120 205.235 75.340 205.465 ;
        RECT 75.510 205.415 75.935 206.035 ;
        RECT 76.130 205.415 76.390 206.035 ;
        RECT 76.585 205.915 76.870 207.055 ;
        RECT 76.600 205.235 76.860 205.745 ;
        RECT 75.120 205.045 76.860 205.235 ;
        RECT 75.120 204.685 75.550 205.045 ;
        RECT 76.130 204.505 76.860 204.875 ;
        RECT 77.060 204.685 77.340 206.875 ;
        RECT 77.545 206.465 77.785 206.855 ;
        RECT 77.955 206.645 78.305 207.055 ;
        RECT 77.545 206.265 78.295 206.465 ;
        RECT 77.545 204.745 77.775 206.085 ;
        RECT 77.955 205.585 78.295 206.265 ;
        RECT 78.475 205.765 78.805 206.875 ;
        RECT 78.975 206.405 79.155 206.875 ;
        RECT 79.325 206.575 79.655 207.055 ;
        RECT 79.830 206.405 80.000 206.875 ;
        RECT 78.975 206.205 80.000 206.405 ;
        RECT 77.955 204.685 78.185 205.585 ;
        RECT 78.475 205.465 79.020 205.765 ;
        RECT 78.385 204.505 78.630 205.285 ;
        RECT 78.800 205.235 79.020 205.465 ;
        RECT 79.190 205.415 79.615 206.035 ;
        RECT 79.810 205.415 80.070 206.035 ;
        RECT 80.265 205.915 80.550 207.055 ;
        RECT 80.280 205.235 80.540 205.745 ;
        RECT 78.800 205.045 80.540 205.235 ;
        RECT 78.800 204.685 79.230 205.045 ;
        RECT 79.810 204.505 80.540 204.875 ;
        RECT 80.740 204.685 81.020 206.875 ;
        RECT 81.265 205.915 81.475 207.055 ;
        RECT 81.645 205.905 81.975 206.885 ;
        RECT 82.145 205.915 82.375 207.055 ;
        RECT 81.265 204.505 81.475 205.325 ;
        RECT 81.645 205.305 81.895 205.905 ;
        RECT 82.585 205.890 82.875 207.055 ;
        RECT 83.065 206.465 83.305 206.855 ;
        RECT 83.475 206.645 83.825 207.055 ;
        RECT 83.065 206.265 83.815 206.465 ;
        RECT 82.065 205.495 82.395 205.745 ;
        RECT 81.645 204.675 81.975 205.305 ;
        RECT 82.145 204.505 82.375 205.325 ;
        RECT 82.585 204.505 82.875 205.230 ;
        RECT 83.065 204.745 83.295 206.085 ;
        RECT 83.475 205.585 83.815 206.265 ;
        RECT 83.995 205.765 84.325 206.875 ;
        RECT 84.495 206.405 84.675 206.875 ;
        RECT 84.845 206.575 85.175 207.055 ;
        RECT 85.350 206.405 85.520 206.875 ;
        RECT 84.495 206.205 85.520 206.405 ;
        RECT 83.475 204.685 83.705 205.585 ;
        RECT 83.995 205.465 84.540 205.765 ;
        RECT 83.905 204.505 84.150 205.285 ;
        RECT 84.320 205.235 84.540 205.465 ;
        RECT 84.710 205.415 85.135 206.035 ;
        RECT 85.330 205.415 85.590 206.035 ;
        RECT 85.785 205.915 86.070 207.055 ;
        RECT 85.800 205.235 86.060 205.745 ;
        RECT 84.320 205.045 86.060 205.235 ;
        RECT 84.320 204.685 84.750 205.045 ;
        RECT 85.330 204.505 86.060 204.875 ;
        RECT 86.260 204.685 86.540 206.875 ;
        RECT 86.725 205.980 86.995 206.885 ;
        RECT 87.165 206.295 87.495 207.055 ;
        RECT 87.675 206.125 87.845 206.885 ;
        RECT 86.725 205.180 86.895 205.980 ;
        RECT 87.180 205.955 87.845 206.125 ;
        RECT 88.105 205.965 89.315 207.055 ;
        RECT 87.180 205.810 87.350 205.955 ;
        RECT 87.065 205.480 87.350 205.810 ;
        RECT 87.180 205.225 87.350 205.480 ;
        RECT 87.585 205.405 87.915 205.775 ;
        RECT 88.105 205.425 88.625 205.965 ;
        RECT 88.795 205.255 89.315 205.795 ;
        RECT 86.725 204.675 86.985 205.180 ;
        RECT 87.180 205.055 87.845 205.225 ;
        RECT 87.165 204.505 87.495 204.885 ;
        RECT 87.675 204.675 87.845 205.055 ;
        RECT 88.105 204.505 89.315 205.255 ;
        RECT 18.100 204.335 89.400 204.505 ;
        RECT 18.185 203.585 19.395 204.335 ;
        RECT 18.185 203.045 18.705 203.585 ;
        RECT 19.570 203.495 19.830 204.335 ;
        RECT 20.005 203.590 20.260 204.165 ;
        RECT 20.430 203.955 20.760 204.335 ;
        RECT 20.975 203.785 21.145 204.165 ;
        RECT 20.430 203.615 21.145 203.785 ;
        RECT 18.875 202.875 19.395 203.415 ;
        RECT 18.185 201.785 19.395 202.875 ;
        RECT 19.570 201.785 19.830 202.935 ;
        RECT 20.005 202.860 20.175 203.590 ;
        RECT 20.430 203.425 20.600 203.615 ;
        RECT 21.405 203.535 21.715 204.335 ;
        RECT 21.920 203.535 22.615 204.165 ;
        RECT 22.785 203.535 23.095 204.335 ;
        RECT 23.300 203.535 23.995 204.165 ;
        RECT 24.210 203.875 24.960 204.165 ;
        RECT 25.470 203.875 25.800 204.335 ;
        RECT 20.345 203.095 20.600 203.425 ;
        RECT 20.430 202.885 20.600 203.095 ;
        RECT 20.880 203.065 21.235 203.435 ;
        RECT 21.415 203.095 21.750 203.365 ;
        RECT 21.920 202.935 22.090 203.535 ;
        RECT 23.300 203.485 23.475 203.535 ;
        RECT 22.260 203.095 22.595 203.345 ;
        RECT 22.795 203.095 23.130 203.365 ;
        RECT 23.300 202.935 23.470 203.485 ;
        RECT 23.640 203.095 23.975 203.345 ;
        RECT 20.005 201.955 20.260 202.860 ;
        RECT 20.430 202.715 21.145 202.885 ;
        RECT 20.430 201.785 20.760 202.545 ;
        RECT 20.975 201.955 21.145 202.715 ;
        RECT 21.405 201.785 21.685 202.925 ;
        RECT 21.855 201.955 22.185 202.935 ;
        RECT 22.355 201.785 22.615 202.925 ;
        RECT 22.785 201.785 23.065 202.925 ;
        RECT 23.235 201.955 23.565 202.935 ;
        RECT 23.735 201.785 23.995 202.925 ;
        RECT 24.210 202.585 24.580 203.875 ;
        RECT 26.020 203.685 26.290 203.895 ;
        RECT 24.955 203.515 26.290 203.685 ;
        RECT 26.465 203.675 26.740 204.335 ;
        RECT 26.910 203.705 27.160 204.165 ;
        RECT 27.335 203.840 27.665 204.335 ;
        RECT 24.955 203.345 25.125 203.515 ;
        RECT 26.910 203.495 27.080 203.705 ;
        RECT 27.845 203.670 28.075 204.115 ;
        RECT 24.750 203.095 25.125 203.345 ;
        RECT 25.295 203.105 25.770 203.345 ;
        RECT 25.940 203.105 26.290 203.345 ;
        RECT 24.955 202.925 25.125 203.095 ;
        RECT 26.465 202.975 27.080 203.495 ;
        RECT 27.250 202.995 27.480 203.425 ;
        RECT 27.665 203.175 28.075 203.670 ;
        RECT 28.245 203.850 29.035 204.115 ;
        RECT 28.245 202.995 28.500 203.850 ;
        RECT 29.425 203.705 29.755 204.065 ;
        RECT 30.385 203.875 30.635 204.335 ;
        RECT 30.805 203.875 31.355 204.165 ;
        RECT 28.670 203.175 29.055 203.655 ;
        RECT 29.425 203.515 30.815 203.705 ;
        RECT 30.645 203.425 30.815 203.515 ;
        RECT 29.225 203.095 29.915 203.345 ;
        RECT 30.145 203.095 30.475 203.345 ;
        RECT 30.645 203.095 30.935 203.425 ;
        RECT 24.955 202.755 26.290 202.925 ;
        RECT 26.010 202.595 26.290 202.755 ;
        RECT 24.210 202.415 25.380 202.585 ;
        RECT 24.665 201.785 24.880 202.245 ;
        RECT 25.050 201.955 25.380 202.415 ;
        RECT 25.550 201.785 25.800 202.585 ;
        RECT 26.465 201.785 26.725 202.795 ;
        RECT 26.895 202.625 27.065 202.975 ;
        RECT 27.250 202.825 29.040 202.995 ;
        RECT 26.895 201.955 27.170 202.625 ;
        RECT 27.370 201.785 27.585 202.630 ;
        RECT 27.810 202.530 28.060 202.825 ;
        RECT 28.285 202.465 28.615 202.655 ;
        RECT 27.770 201.955 28.245 202.295 ;
        RECT 28.425 202.290 28.615 202.465 ;
        RECT 28.785 202.460 29.040 202.825 ;
        RECT 29.225 202.655 29.540 203.095 ;
        RECT 30.645 202.845 30.815 203.095 ;
        RECT 29.875 202.675 30.815 202.845 ;
        RECT 28.425 201.785 29.055 202.290 ;
        RECT 29.425 201.785 29.705 202.455 ;
        RECT 29.875 202.125 30.175 202.675 ;
        RECT 31.105 202.505 31.355 203.875 ;
        RECT 31.525 203.535 31.815 204.335 ;
        RECT 32.045 203.855 32.325 204.335 ;
        RECT 32.495 203.685 32.755 204.075 ;
        RECT 32.930 203.855 33.185 204.335 ;
        RECT 33.355 203.685 33.650 204.075 ;
        RECT 33.830 203.855 34.105 204.335 ;
        RECT 34.275 203.835 34.575 204.165 ;
        RECT 34.835 203.855 35.135 204.335 ;
        RECT 32.000 203.515 33.650 203.685 ;
        RECT 32.000 203.005 32.405 203.515 ;
        RECT 32.575 203.175 33.715 203.345 ;
        RECT 30.385 201.785 30.715 202.505 ;
        RECT 30.905 201.955 31.355 202.505 ;
        RECT 31.525 201.785 31.815 202.925 ;
        RECT 32.000 202.835 32.755 203.005 ;
        RECT 32.040 201.785 32.325 202.655 ;
        RECT 32.495 202.585 32.755 202.835 ;
        RECT 33.545 202.925 33.715 203.175 ;
        RECT 33.885 203.095 34.235 203.665 ;
        RECT 34.405 202.925 34.575 203.835 ;
        RECT 35.305 203.685 35.565 204.140 ;
        RECT 35.735 203.855 35.995 204.335 ;
        RECT 36.175 203.685 36.435 204.140 ;
        RECT 36.605 203.855 36.855 204.335 ;
        RECT 37.035 203.685 37.295 204.140 ;
        RECT 37.465 203.855 37.715 204.335 ;
        RECT 37.895 203.685 38.155 204.140 ;
        RECT 38.325 203.855 38.570 204.335 ;
        RECT 38.740 203.685 39.015 204.140 ;
        RECT 39.185 203.855 39.430 204.335 ;
        RECT 39.600 203.685 39.860 204.140 ;
        RECT 40.030 203.855 40.290 204.335 ;
        RECT 40.460 203.685 40.720 204.140 ;
        RECT 40.890 203.855 41.150 204.335 ;
        RECT 41.320 203.685 41.580 204.140 ;
        RECT 41.750 203.775 42.010 204.335 ;
        RECT 33.545 202.755 34.575 202.925 ;
        RECT 32.495 202.415 33.615 202.585 ;
        RECT 32.495 201.955 32.755 202.415 ;
        RECT 32.930 201.785 33.185 202.245 ;
        RECT 33.355 201.955 33.615 202.415 ;
        RECT 33.785 201.785 34.095 202.585 ;
        RECT 34.265 201.955 34.575 202.755 ;
        RECT 34.835 203.515 41.580 203.685 ;
        RECT 34.835 202.925 36.000 203.515 ;
        RECT 42.180 203.345 42.430 204.155 ;
        RECT 42.610 203.810 42.870 204.335 ;
        RECT 43.040 203.345 43.290 204.155 ;
        RECT 43.470 203.825 43.775 204.335 ;
        RECT 36.170 203.095 43.290 203.345 ;
        RECT 43.460 203.095 43.775 203.655 ;
        RECT 43.945 203.610 44.235 204.335 ;
        RECT 45.325 203.825 45.630 204.335 ;
        RECT 45.325 203.095 45.640 203.655 ;
        RECT 45.810 203.345 46.060 204.155 ;
        RECT 46.230 203.810 46.490 204.335 ;
        RECT 46.670 203.345 46.920 204.155 ;
        RECT 47.090 203.775 47.350 204.335 ;
        RECT 47.520 203.685 47.780 204.140 ;
        RECT 47.950 203.855 48.210 204.335 ;
        RECT 48.380 203.685 48.640 204.140 ;
        RECT 48.810 203.855 49.070 204.335 ;
        RECT 49.240 203.685 49.500 204.140 ;
        RECT 49.670 203.855 49.915 204.335 ;
        RECT 50.085 203.685 50.360 204.140 ;
        RECT 50.530 203.855 50.775 204.335 ;
        RECT 50.945 203.685 51.205 204.140 ;
        RECT 51.385 203.855 51.635 204.335 ;
        RECT 51.805 203.685 52.065 204.140 ;
        RECT 52.245 203.855 52.495 204.335 ;
        RECT 52.665 203.685 52.925 204.140 ;
        RECT 53.105 203.855 53.365 204.335 ;
        RECT 53.535 203.685 53.795 204.140 ;
        RECT 53.965 203.855 54.265 204.335 ;
        RECT 54.615 203.855 54.915 204.335 ;
        RECT 55.085 203.685 55.345 204.140 ;
        RECT 55.515 203.855 55.775 204.335 ;
        RECT 55.955 203.685 56.215 204.140 ;
        RECT 56.385 203.855 56.635 204.335 ;
        RECT 56.815 203.685 57.075 204.140 ;
        RECT 57.245 203.855 57.495 204.335 ;
        RECT 57.675 203.685 57.935 204.140 ;
        RECT 58.105 203.855 58.350 204.335 ;
        RECT 58.520 203.685 58.795 204.140 ;
        RECT 58.965 203.855 59.210 204.335 ;
        RECT 59.380 203.685 59.640 204.140 ;
        RECT 59.810 203.855 60.070 204.335 ;
        RECT 60.240 203.685 60.500 204.140 ;
        RECT 60.670 203.855 60.930 204.335 ;
        RECT 61.100 203.685 61.360 204.140 ;
        RECT 61.530 203.775 61.790 204.335 ;
        RECT 47.520 203.515 54.265 203.685 ;
        RECT 45.810 203.095 52.930 203.345 ;
        RECT 34.835 202.700 41.580 202.925 ;
        RECT 34.835 201.785 35.105 202.530 ;
        RECT 35.275 201.960 35.565 202.700 ;
        RECT 36.175 202.685 41.580 202.700 ;
        RECT 35.735 201.790 35.990 202.515 ;
        RECT 36.175 201.960 36.435 202.685 ;
        RECT 36.605 201.790 36.850 202.515 ;
        RECT 37.035 201.960 37.295 202.685 ;
        RECT 37.465 201.790 37.710 202.515 ;
        RECT 37.895 201.960 38.155 202.685 ;
        RECT 38.325 201.790 38.570 202.515 ;
        RECT 38.740 201.960 39.000 202.685 ;
        RECT 39.170 201.790 39.430 202.515 ;
        RECT 39.600 201.960 39.860 202.685 ;
        RECT 40.030 201.790 40.290 202.515 ;
        RECT 40.460 201.960 40.720 202.685 ;
        RECT 40.890 201.790 41.150 202.515 ;
        RECT 41.320 201.960 41.580 202.685 ;
        RECT 41.750 201.790 42.010 202.585 ;
        RECT 42.180 201.960 42.430 203.095 ;
        RECT 35.735 201.785 42.010 201.790 ;
        RECT 42.610 201.785 42.870 202.595 ;
        RECT 43.045 201.955 43.290 203.095 ;
        RECT 43.470 201.785 43.765 202.595 ;
        RECT 43.945 201.785 44.235 202.950 ;
        RECT 45.335 201.785 45.630 202.595 ;
        RECT 45.810 201.955 46.055 203.095 ;
        RECT 46.230 201.785 46.490 202.595 ;
        RECT 46.670 201.960 46.920 203.095 ;
        RECT 53.100 202.925 54.265 203.515 ;
        RECT 47.520 202.700 54.265 202.925 ;
        RECT 54.615 203.515 61.360 203.685 ;
        RECT 54.615 202.925 55.780 203.515 ;
        RECT 61.960 203.345 62.210 204.155 ;
        RECT 62.390 203.810 62.650 204.335 ;
        RECT 62.820 203.345 63.070 204.155 ;
        RECT 63.250 203.825 63.555 204.335 ;
        RECT 55.950 203.095 63.070 203.345 ;
        RECT 63.240 203.095 63.555 203.655 ;
        RECT 63.735 203.525 64.005 204.335 ;
        RECT 64.175 203.525 64.505 204.165 ;
        RECT 64.675 203.525 64.915 204.335 ;
        RECT 65.110 203.955 67.125 204.125 ;
        RECT 67.315 203.955 67.645 204.335 ;
        RECT 65.110 203.635 65.365 203.955 ;
        RECT 63.725 203.095 64.075 203.345 ;
        RECT 54.615 202.700 61.360 202.925 ;
        RECT 47.520 202.685 52.925 202.700 ;
        RECT 47.090 201.790 47.350 202.585 ;
        RECT 47.520 201.960 47.780 202.685 ;
        RECT 47.950 201.790 48.210 202.515 ;
        RECT 48.380 201.960 48.640 202.685 ;
        RECT 48.810 201.790 49.070 202.515 ;
        RECT 49.240 201.960 49.500 202.685 ;
        RECT 49.670 201.790 49.930 202.515 ;
        RECT 50.100 201.960 50.360 202.685 ;
        RECT 50.530 201.790 50.775 202.515 ;
        RECT 50.945 201.960 51.205 202.685 ;
        RECT 51.390 201.790 51.635 202.515 ;
        RECT 51.805 201.960 52.065 202.685 ;
        RECT 52.250 201.790 52.495 202.515 ;
        RECT 52.665 201.960 52.925 202.685 ;
        RECT 53.110 201.790 53.365 202.515 ;
        RECT 53.535 201.960 53.825 202.700 ;
        RECT 47.090 201.785 53.365 201.790 ;
        RECT 53.995 201.785 54.265 202.530 ;
        RECT 54.615 201.785 54.885 202.530 ;
        RECT 55.055 201.960 55.345 202.700 ;
        RECT 55.955 202.685 61.360 202.700 ;
        RECT 55.515 201.790 55.770 202.515 ;
        RECT 55.955 201.960 56.215 202.685 ;
        RECT 56.385 201.790 56.630 202.515 ;
        RECT 56.815 201.960 57.075 202.685 ;
        RECT 57.245 201.790 57.490 202.515 ;
        RECT 57.675 201.960 57.935 202.685 ;
        RECT 58.105 201.790 58.350 202.515 ;
        RECT 58.520 201.960 58.780 202.685 ;
        RECT 58.950 201.790 59.210 202.515 ;
        RECT 59.380 201.960 59.640 202.685 ;
        RECT 59.810 201.790 60.070 202.515 ;
        RECT 60.240 201.960 60.500 202.685 ;
        RECT 60.670 201.790 60.930 202.515 ;
        RECT 61.100 201.960 61.360 202.685 ;
        RECT 61.530 201.790 61.790 202.585 ;
        RECT 61.960 201.960 62.210 203.095 ;
        RECT 55.515 201.785 61.790 201.790 ;
        RECT 62.390 201.785 62.650 202.595 ;
        RECT 62.825 201.955 63.070 203.095 ;
        RECT 64.245 202.925 64.415 203.525 ;
        RECT 64.585 203.095 64.935 203.345 ;
        RECT 65.110 203.095 65.350 203.425 ;
        RECT 65.535 202.975 65.865 203.785 ;
        RECT 66.375 203.515 68.065 203.785 ;
        RECT 68.235 203.535 68.615 204.335 ;
        RECT 69.705 203.610 69.995 204.335 ;
        RECT 66.090 203.145 67.180 203.345 ;
        RECT 67.490 203.145 68.615 203.345 ;
        RECT 63.250 201.785 63.545 202.595 ;
        RECT 63.735 201.785 64.065 202.925 ;
        RECT 64.245 202.755 64.925 202.925 ;
        RECT 64.595 201.970 64.925 202.755 ;
        RECT 65.110 201.785 65.365 202.925 ;
        RECT 65.535 202.755 68.065 202.975 ;
        RECT 65.535 201.955 65.865 202.755 ;
        RECT 66.035 201.785 66.205 202.585 ;
        RECT 66.375 201.955 66.705 202.755 ;
        RECT 66.875 201.785 67.565 202.585 ;
        RECT 67.735 201.955 68.065 202.755 ;
        RECT 68.235 201.785 68.615 202.975 ;
        RECT 69.705 201.785 69.995 202.950 ;
        RECT 70.180 201.965 70.460 204.155 ;
        RECT 70.660 203.965 71.390 204.335 ;
        RECT 71.970 203.795 72.400 204.155 ;
        RECT 70.660 203.605 72.400 203.795 ;
        RECT 70.660 203.095 70.920 203.605 ;
        RECT 70.650 201.785 70.935 202.925 ;
        RECT 71.130 202.805 71.390 203.425 ;
        RECT 71.585 202.805 72.010 203.425 ;
        RECT 72.180 203.375 72.400 203.605 ;
        RECT 72.570 203.555 72.815 204.335 ;
        RECT 72.180 203.075 72.725 203.375 ;
        RECT 73.015 203.255 73.245 204.155 ;
        RECT 71.200 202.435 72.225 202.635 ;
        RECT 71.200 201.965 71.370 202.435 ;
        RECT 71.545 201.785 71.875 202.265 ;
        RECT 72.045 201.965 72.225 202.435 ;
        RECT 72.395 201.965 72.725 203.075 ;
        RECT 72.905 202.575 73.245 203.255 ;
        RECT 73.425 202.755 73.655 204.095 ;
        RECT 73.885 203.515 74.115 204.335 ;
        RECT 74.285 203.535 74.615 204.165 ;
        RECT 73.865 203.095 74.195 203.345 ;
        RECT 74.365 202.935 74.615 203.535 ;
        RECT 74.785 203.515 74.995 204.335 ;
        RECT 75.315 203.855 75.615 204.335 ;
        RECT 75.785 203.685 76.045 204.140 ;
        RECT 76.215 203.855 76.475 204.335 ;
        RECT 76.655 203.685 76.915 204.140 ;
        RECT 77.085 203.855 77.335 204.335 ;
        RECT 77.515 203.685 77.775 204.140 ;
        RECT 77.945 203.855 78.195 204.335 ;
        RECT 78.375 203.685 78.635 204.140 ;
        RECT 78.805 203.855 79.050 204.335 ;
        RECT 79.220 203.685 79.495 204.140 ;
        RECT 79.665 203.855 79.910 204.335 ;
        RECT 80.080 203.685 80.340 204.140 ;
        RECT 80.510 203.855 80.770 204.335 ;
        RECT 80.940 203.685 81.200 204.140 ;
        RECT 81.370 203.855 81.630 204.335 ;
        RECT 81.800 203.685 82.060 204.140 ;
        RECT 82.230 203.775 82.490 204.335 ;
        RECT 75.315 203.515 82.060 203.685 ;
        RECT 72.905 202.375 73.655 202.575 ;
        RECT 72.895 201.785 73.245 202.195 ;
        RECT 73.415 201.985 73.655 202.375 ;
        RECT 73.885 201.785 74.115 202.925 ;
        RECT 74.285 201.955 74.615 202.935 ;
        RECT 75.315 202.925 76.480 203.515 ;
        RECT 82.660 203.345 82.910 204.155 ;
        RECT 83.090 203.810 83.350 204.335 ;
        RECT 83.520 203.345 83.770 204.155 ;
        RECT 83.950 203.825 84.255 204.335 ;
        RECT 84.425 203.855 84.685 204.335 ;
        RECT 84.855 204.085 85.100 204.165 ;
        RECT 84.855 203.915 85.185 204.085 ;
        RECT 76.650 203.095 83.770 203.345 ;
        RECT 83.940 203.095 84.255 203.655 ;
        RECT 84.470 203.095 84.665 203.665 ;
        RECT 74.785 201.785 74.995 202.925 ;
        RECT 75.315 202.700 82.060 202.925 ;
        RECT 75.315 201.785 75.585 202.530 ;
        RECT 75.755 201.960 76.045 202.700 ;
        RECT 76.655 202.685 82.060 202.700 ;
        RECT 76.215 201.790 76.470 202.515 ;
        RECT 76.655 201.960 76.915 202.685 ;
        RECT 77.085 201.790 77.330 202.515 ;
        RECT 77.515 201.960 77.775 202.685 ;
        RECT 77.945 201.790 78.190 202.515 ;
        RECT 78.375 201.960 78.635 202.685 ;
        RECT 78.805 201.790 79.050 202.515 ;
        RECT 79.220 201.960 79.480 202.685 ;
        RECT 79.650 201.790 79.910 202.515 ;
        RECT 80.080 201.960 80.340 202.685 ;
        RECT 80.510 201.790 80.770 202.515 ;
        RECT 80.940 201.960 81.200 202.685 ;
        RECT 81.370 201.790 81.630 202.515 ;
        RECT 81.800 201.960 82.060 202.685 ;
        RECT 82.230 201.790 82.490 202.585 ;
        RECT 82.660 201.960 82.910 203.095 ;
        RECT 76.215 201.785 82.490 201.790 ;
        RECT 83.090 201.785 83.350 202.595 ;
        RECT 83.525 201.955 83.770 203.095 ;
        RECT 84.855 202.925 85.025 203.915 ;
        RECT 85.385 203.720 85.595 204.005 ;
        RECT 85.860 203.995 86.030 204.020 ;
        RECT 85.860 203.825 86.035 203.995 ;
        RECT 86.275 203.955 86.605 204.335 ;
        RECT 86.795 203.995 86.965 204.165 ;
        RECT 86.375 203.875 86.545 203.955 ;
        RECT 86.785 203.825 86.965 203.995 ;
        RECT 87.215 203.875 87.470 204.335 ;
        RECT 85.860 203.725 86.030 203.825 ;
        RECT 85.205 203.550 85.595 203.720 ;
        RECT 85.765 203.555 86.030 203.725 ;
        RECT 86.795 203.705 86.965 203.825 ;
        RECT 85.205 203.485 85.485 203.550 ;
        RECT 85.205 203.095 85.375 203.485 ;
        RECT 85.765 203.345 85.935 203.555 ;
        RECT 86.290 203.425 86.495 203.660 ;
        RECT 86.795 203.535 87.470 203.705 ;
        RECT 88.105 203.585 89.315 204.335 ;
        RECT 85.605 203.175 85.935 203.345 ;
        RECT 85.765 203.160 85.935 203.175 ;
        RECT 86.165 203.095 86.495 203.425 ;
        RECT 86.675 203.175 87.005 203.345 ;
        RECT 86.835 202.925 87.005 203.175 ;
        RECT 84.515 202.755 87.005 202.925 ;
        RECT 83.950 201.785 84.245 202.595 ;
        RECT 84.515 201.955 84.685 202.755 ;
        RECT 87.215 202.585 87.470 203.535 ;
        RECT 84.915 202.415 86.205 202.585 ;
        RECT 84.975 201.995 85.225 202.415 ;
        RECT 85.415 201.785 85.745 202.245 ;
        RECT 85.955 201.995 86.205 202.415 ;
        RECT 86.375 201.785 86.625 202.585 ;
        RECT 86.795 202.415 87.470 202.585 ;
        RECT 88.105 202.875 88.625 203.415 ;
        RECT 88.795 203.045 89.315 203.585 ;
        RECT 86.795 201.955 86.965 202.415 ;
        RECT 87.175 201.785 87.425 202.245 ;
        RECT 88.105 201.785 89.315 202.875 ;
        RECT 18.100 201.615 89.400 201.785 ;
        RECT 18.185 200.525 19.395 201.615 ;
        RECT 18.185 199.815 18.705 200.355 ;
        RECT 18.875 199.985 19.395 200.525 ;
        RECT 20.575 200.685 20.745 201.445 ;
        RECT 20.960 200.855 21.290 201.615 ;
        RECT 20.575 200.515 21.290 200.685 ;
        RECT 21.460 200.540 21.715 201.445 ;
        RECT 20.485 199.965 20.840 200.335 ;
        RECT 21.120 200.305 21.290 200.515 ;
        RECT 21.120 199.975 21.375 200.305 ;
        RECT 18.185 199.065 19.395 199.815 ;
        RECT 21.120 199.785 21.290 199.975 ;
        RECT 21.545 199.810 21.715 200.540 ;
        RECT 21.890 200.465 22.150 201.615 ;
        RECT 22.330 200.465 22.590 201.615 ;
        RECT 22.765 200.540 23.020 201.445 ;
        RECT 23.190 200.855 23.520 201.615 ;
        RECT 23.735 200.685 23.905 201.445 ;
        RECT 20.575 199.615 21.290 199.785 ;
        RECT 20.575 199.235 20.745 199.615 ;
        RECT 20.960 199.065 21.290 199.445 ;
        RECT 21.460 199.235 21.715 199.810 ;
        RECT 21.890 199.065 22.150 199.905 ;
        RECT 22.330 199.065 22.590 199.905 ;
        RECT 22.765 199.810 22.935 200.540 ;
        RECT 23.190 200.515 23.905 200.685 ;
        RECT 23.190 200.305 23.360 200.515 ;
        RECT 25.085 200.475 25.365 201.615 ;
        RECT 25.535 200.465 25.865 201.445 ;
        RECT 26.035 200.475 26.295 201.615 ;
        RECT 26.665 200.945 26.945 201.615 ;
        RECT 27.115 200.725 27.415 201.275 ;
        RECT 27.615 200.895 27.945 201.615 ;
        RECT 28.135 200.895 28.595 201.445 ;
        RECT 23.105 199.975 23.360 200.305 ;
        RECT 22.765 199.235 23.020 199.810 ;
        RECT 23.190 199.785 23.360 199.975 ;
        RECT 23.640 199.965 23.995 200.335 ;
        RECT 25.095 200.035 25.430 200.305 ;
        RECT 25.600 199.865 25.770 200.465 ;
        RECT 26.480 200.305 26.745 200.665 ;
        RECT 27.115 200.555 28.055 200.725 ;
        RECT 27.885 200.305 28.055 200.555 ;
        RECT 25.940 200.055 26.275 200.305 ;
        RECT 26.480 200.055 27.155 200.305 ;
        RECT 27.375 200.055 27.715 200.305 ;
        RECT 27.885 199.975 28.175 200.305 ;
        RECT 27.885 199.885 28.055 199.975 ;
        RECT 23.190 199.615 23.905 199.785 ;
        RECT 23.190 199.065 23.520 199.445 ;
        RECT 23.735 199.235 23.905 199.615 ;
        RECT 25.085 199.065 25.395 199.865 ;
        RECT 25.600 199.235 26.295 199.865 ;
        RECT 26.665 199.695 28.055 199.885 ;
        RECT 26.665 199.335 26.995 199.695 ;
        RECT 28.345 199.525 28.595 200.895 ;
        RECT 28.785 200.815 29.065 201.615 ;
        RECT 29.265 200.645 29.595 201.445 ;
        RECT 29.795 200.815 29.965 201.615 ;
        RECT 30.135 200.645 30.465 201.445 ;
        RECT 28.765 199.975 29.005 200.645 ;
        RECT 29.185 200.475 30.465 200.645 ;
        RECT 30.635 200.475 30.895 201.615 ;
        RECT 29.185 199.805 29.355 200.475 ;
        RECT 31.065 200.450 31.355 201.615 ;
        RECT 31.525 200.540 31.795 201.445 ;
        RECT 31.965 200.855 32.295 201.615 ;
        RECT 32.475 200.685 32.645 201.445 ;
        RECT 29.525 199.975 29.835 200.305 ;
        RECT 30.005 199.975 30.385 200.305 ;
        RECT 30.585 199.975 30.870 200.305 ;
        RECT 29.630 199.805 29.835 199.975 ;
        RECT 27.615 199.065 27.865 199.525 ;
        RECT 28.035 199.235 28.595 199.525 ;
        RECT 28.765 199.235 29.460 199.805 ;
        RECT 29.630 199.280 29.980 199.805 ;
        RECT 30.170 199.280 30.385 199.975 ;
        RECT 30.555 199.065 30.890 199.805 ;
        RECT 31.065 199.065 31.355 199.790 ;
        RECT 31.525 199.740 31.695 200.540 ;
        RECT 31.980 200.515 32.645 200.685 ;
        RECT 32.925 200.725 33.185 201.435 ;
        RECT 33.355 200.905 33.685 201.615 ;
        RECT 33.855 200.725 34.085 201.435 ;
        RECT 31.980 200.370 32.150 200.515 ;
        RECT 32.925 200.485 34.085 200.725 ;
        RECT 34.265 200.705 34.535 201.435 ;
        RECT 34.715 200.885 35.055 201.615 ;
        RECT 34.265 200.485 35.035 200.705 ;
        RECT 31.865 200.040 32.150 200.370 ;
        RECT 31.980 199.785 32.150 200.040 ;
        RECT 32.385 199.965 32.715 200.335 ;
        RECT 32.915 199.975 33.215 200.305 ;
        RECT 33.395 199.995 33.920 200.305 ;
        RECT 34.100 199.995 34.565 200.305 ;
        RECT 31.525 199.235 31.785 199.740 ;
        RECT 31.980 199.615 32.645 199.785 ;
        RECT 31.965 199.065 32.295 199.445 ;
        RECT 32.475 199.235 32.645 199.615 ;
        RECT 32.925 199.065 33.215 199.795 ;
        RECT 33.395 199.355 33.625 199.995 ;
        RECT 34.745 199.815 35.035 200.485 ;
        RECT 33.805 199.615 35.035 199.815 ;
        RECT 33.805 199.245 34.115 199.615 ;
        RECT 34.295 199.065 34.965 199.435 ;
        RECT 35.225 199.245 35.485 201.435 ;
        RECT 35.665 200.645 35.975 201.445 ;
        RECT 36.145 200.815 36.455 201.615 ;
        RECT 36.625 200.985 36.885 201.445 ;
        RECT 37.055 201.155 37.310 201.615 ;
        RECT 37.485 200.985 37.745 201.445 ;
        RECT 36.625 200.815 37.745 200.985 ;
        RECT 35.665 200.475 36.695 200.645 ;
        RECT 35.665 199.565 35.835 200.475 ;
        RECT 36.005 199.735 36.355 200.305 ;
        RECT 36.525 200.225 36.695 200.475 ;
        RECT 37.485 200.565 37.745 200.815 ;
        RECT 37.915 200.745 38.200 201.615 ;
        RECT 38.515 200.870 38.785 201.615 ;
        RECT 39.415 201.610 45.690 201.615 ;
        RECT 38.955 200.700 39.245 201.440 ;
        RECT 39.415 200.885 39.670 201.610 ;
        RECT 39.855 200.715 40.115 201.440 ;
        RECT 40.285 200.885 40.530 201.610 ;
        RECT 40.715 200.715 40.975 201.440 ;
        RECT 41.145 200.885 41.390 201.610 ;
        RECT 41.575 200.715 41.835 201.440 ;
        RECT 42.005 200.885 42.250 201.610 ;
        RECT 42.420 200.715 42.680 201.440 ;
        RECT 42.850 200.885 43.110 201.610 ;
        RECT 43.280 200.715 43.540 201.440 ;
        RECT 43.710 200.885 43.970 201.610 ;
        RECT 44.140 200.715 44.400 201.440 ;
        RECT 44.570 200.885 44.830 201.610 ;
        RECT 45.000 200.715 45.260 201.440 ;
        RECT 45.430 200.815 45.690 201.610 ;
        RECT 39.855 200.700 45.260 200.715 ;
        RECT 37.485 200.395 38.240 200.565 ;
        RECT 36.525 200.055 37.665 200.225 ;
        RECT 37.835 199.885 38.240 200.395 ;
        RECT 36.590 199.715 38.240 199.885 ;
        RECT 38.515 200.475 45.260 200.700 ;
        RECT 38.515 199.885 39.680 200.475 ;
        RECT 45.860 200.305 46.110 201.440 ;
        RECT 46.290 200.805 46.550 201.615 ;
        RECT 46.725 200.305 46.970 201.445 ;
        RECT 47.150 200.805 47.445 201.615 ;
        RECT 47.715 200.870 47.985 201.615 ;
        RECT 48.615 201.610 54.890 201.615 ;
        RECT 48.155 200.700 48.445 201.440 ;
        RECT 48.615 200.885 48.870 201.610 ;
        RECT 49.055 200.715 49.315 201.440 ;
        RECT 49.485 200.885 49.730 201.610 ;
        RECT 49.915 200.715 50.175 201.440 ;
        RECT 50.345 200.885 50.590 201.610 ;
        RECT 50.775 200.715 51.035 201.440 ;
        RECT 51.205 200.885 51.450 201.610 ;
        RECT 51.620 200.715 51.880 201.440 ;
        RECT 52.050 200.885 52.310 201.610 ;
        RECT 52.480 200.715 52.740 201.440 ;
        RECT 52.910 200.885 53.170 201.610 ;
        RECT 53.340 200.715 53.600 201.440 ;
        RECT 53.770 200.885 54.030 201.610 ;
        RECT 54.200 200.715 54.460 201.440 ;
        RECT 54.630 200.815 54.890 201.610 ;
        RECT 49.055 200.700 54.460 200.715 ;
        RECT 47.715 200.475 54.460 200.700 ;
        RECT 39.850 200.055 46.970 200.305 ;
        RECT 38.515 199.715 45.260 199.885 ;
        RECT 35.665 199.235 35.965 199.565 ;
        RECT 36.135 199.065 36.410 199.545 ;
        RECT 36.590 199.325 36.885 199.715 ;
        RECT 37.055 199.065 37.310 199.545 ;
        RECT 37.485 199.325 37.745 199.715 ;
        RECT 37.915 199.065 38.195 199.545 ;
        RECT 38.515 199.065 38.815 199.545 ;
        RECT 38.985 199.260 39.245 199.715 ;
        RECT 39.415 199.065 39.675 199.545 ;
        RECT 39.855 199.260 40.115 199.715 ;
        RECT 40.285 199.065 40.535 199.545 ;
        RECT 40.715 199.260 40.975 199.715 ;
        RECT 41.145 199.065 41.395 199.545 ;
        RECT 41.575 199.260 41.835 199.715 ;
        RECT 42.005 199.065 42.250 199.545 ;
        RECT 42.420 199.260 42.695 199.715 ;
        RECT 42.865 199.065 43.110 199.545 ;
        RECT 43.280 199.260 43.540 199.715 ;
        RECT 43.710 199.065 43.970 199.545 ;
        RECT 44.140 199.260 44.400 199.715 ;
        RECT 44.570 199.065 44.830 199.545 ;
        RECT 45.000 199.260 45.260 199.715 ;
        RECT 45.430 199.065 45.690 199.625 ;
        RECT 45.860 199.245 46.110 200.055 ;
        RECT 46.290 199.065 46.550 199.590 ;
        RECT 46.720 199.245 46.970 200.055 ;
        RECT 47.140 199.745 47.455 200.305 ;
        RECT 47.715 199.885 48.880 200.475 ;
        RECT 55.060 200.305 55.310 201.440 ;
        RECT 55.490 200.805 55.750 201.615 ;
        RECT 55.925 200.305 56.170 201.445 ;
        RECT 56.350 200.805 56.645 201.615 ;
        RECT 56.825 200.450 57.115 201.615 ;
        RECT 57.285 200.645 57.575 201.445 ;
        RECT 57.745 200.815 57.980 201.615 ;
        RECT 58.165 201.275 59.700 201.445 ;
        RECT 58.165 200.645 58.495 201.275 ;
        RECT 57.285 200.475 58.495 200.645 ;
        RECT 49.050 200.055 56.170 200.305 ;
        RECT 47.715 199.715 54.460 199.885 ;
        RECT 47.150 199.065 47.455 199.575 ;
        RECT 47.715 199.065 48.015 199.545 ;
        RECT 48.185 199.260 48.445 199.715 ;
        RECT 48.615 199.065 48.875 199.545 ;
        RECT 49.055 199.260 49.315 199.715 ;
        RECT 49.485 199.065 49.735 199.545 ;
        RECT 49.915 199.260 50.175 199.715 ;
        RECT 50.345 199.065 50.595 199.545 ;
        RECT 50.775 199.260 51.035 199.715 ;
        RECT 51.205 199.065 51.450 199.545 ;
        RECT 51.620 199.260 51.895 199.715 ;
        RECT 52.065 199.065 52.310 199.545 ;
        RECT 52.480 199.260 52.740 199.715 ;
        RECT 52.910 199.065 53.170 199.545 ;
        RECT 53.340 199.260 53.600 199.715 ;
        RECT 53.770 199.065 54.030 199.545 ;
        RECT 54.200 199.260 54.460 199.715 ;
        RECT 54.630 199.065 54.890 199.625 ;
        RECT 55.060 199.245 55.310 200.055 ;
        RECT 55.490 199.065 55.750 199.590 ;
        RECT 55.920 199.245 56.170 200.055 ;
        RECT 56.340 199.745 56.655 200.305 ;
        RECT 57.285 199.975 57.530 200.305 ;
        RECT 57.700 199.805 57.870 200.475 ;
        RECT 58.665 200.305 58.900 201.050 ;
        RECT 58.040 199.975 58.440 200.305 ;
        RECT 58.610 199.975 58.900 200.305 ;
        RECT 59.090 200.305 59.360 201.050 ;
        RECT 59.530 200.645 59.700 201.275 ;
        RECT 59.870 200.815 60.265 201.615 ;
        RECT 59.530 200.475 60.265 200.645 ;
        RECT 59.090 199.975 59.420 200.305 ;
        RECT 59.590 199.975 59.925 200.305 ;
        RECT 60.095 199.975 60.265 200.475 ;
        RECT 60.435 200.295 60.790 201.445 ;
        RECT 60.960 200.465 61.255 201.615 ;
        RECT 61.435 200.475 61.765 201.615 ;
        RECT 62.295 200.645 62.625 201.430 ;
        RECT 62.815 200.805 63.110 201.615 ;
        RECT 61.945 200.475 62.625 200.645 ;
        RECT 60.435 200.035 61.255 200.295 ;
        RECT 61.425 200.055 61.775 200.305 ;
        RECT 60.435 199.975 60.790 200.035 ;
        RECT 56.350 199.065 56.655 199.575 ;
        RECT 56.825 199.065 57.115 199.790 ;
        RECT 57.285 199.235 57.870 199.805 ;
        RECT 58.120 199.635 59.505 199.805 ;
        RECT 58.120 199.290 58.450 199.635 ;
        RECT 58.665 199.065 59.040 199.465 ;
        RECT 59.220 199.290 59.505 199.635 ;
        RECT 59.675 199.065 60.345 199.805 ;
        RECT 60.515 199.235 60.790 199.975 ;
        RECT 61.945 199.875 62.115 200.475 ;
        RECT 63.290 200.305 63.535 201.445 ;
        RECT 63.710 200.805 63.970 201.615 ;
        RECT 64.570 201.610 70.845 201.615 ;
        RECT 64.150 200.305 64.400 201.440 ;
        RECT 64.570 200.815 64.830 201.610 ;
        RECT 65.000 200.715 65.260 201.440 ;
        RECT 65.430 200.885 65.690 201.610 ;
        RECT 65.860 200.715 66.120 201.440 ;
        RECT 66.290 200.885 66.550 201.610 ;
        RECT 66.720 200.715 66.980 201.440 ;
        RECT 67.150 200.885 67.410 201.610 ;
        RECT 67.580 200.715 67.840 201.440 ;
        RECT 68.010 200.885 68.255 201.610 ;
        RECT 68.425 200.715 68.685 201.440 ;
        RECT 68.870 200.885 69.115 201.610 ;
        RECT 69.285 200.715 69.545 201.440 ;
        RECT 69.730 200.885 69.975 201.610 ;
        RECT 70.145 200.715 70.405 201.440 ;
        RECT 70.590 200.885 70.845 201.610 ;
        RECT 65.000 200.700 70.405 200.715 ;
        RECT 71.015 200.700 71.305 201.440 ;
        RECT 71.475 200.870 71.745 201.615 ;
        RECT 72.015 200.805 72.310 201.615 ;
        RECT 65.000 200.475 71.745 200.700 ;
        RECT 62.285 200.055 62.635 200.305 ;
        RECT 60.960 199.065 61.255 199.865 ;
        RECT 61.435 199.065 61.705 199.875 ;
        RECT 61.875 199.235 62.205 199.875 ;
        RECT 62.375 199.065 62.615 199.875 ;
        RECT 62.805 199.745 63.120 200.305 ;
        RECT 63.290 200.055 70.410 200.305 ;
        RECT 62.805 199.065 63.110 199.575 ;
        RECT 63.290 199.245 63.540 200.055 ;
        RECT 63.710 199.065 63.970 199.590 ;
        RECT 64.150 199.245 64.400 200.055 ;
        RECT 70.580 199.885 71.745 200.475 ;
        RECT 72.490 200.305 72.735 201.445 ;
        RECT 72.910 200.805 73.170 201.615 ;
        RECT 73.770 201.610 80.045 201.615 ;
        RECT 73.350 200.305 73.600 201.440 ;
        RECT 73.770 200.815 74.030 201.610 ;
        RECT 74.200 200.715 74.460 201.440 ;
        RECT 74.630 200.885 74.890 201.610 ;
        RECT 75.060 200.715 75.320 201.440 ;
        RECT 75.490 200.885 75.750 201.610 ;
        RECT 75.920 200.715 76.180 201.440 ;
        RECT 76.350 200.885 76.610 201.610 ;
        RECT 76.780 200.715 77.040 201.440 ;
        RECT 77.210 200.885 77.455 201.610 ;
        RECT 77.625 200.715 77.885 201.440 ;
        RECT 78.070 200.885 78.315 201.610 ;
        RECT 78.485 200.715 78.745 201.440 ;
        RECT 78.930 200.885 79.175 201.610 ;
        RECT 79.345 200.715 79.605 201.440 ;
        RECT 79.790 200.885 80.045 201.610 ;
        RECT 74.200 200.700 79.605 200.715 ;
        RECT 80.215 200.700 80.505 201.440 ;
        RECT 80.675 200.870 80.945 201.615 ;
        RECT 74.200 200.475 80.945 200.700 ;
        RECT 81.295 200.685 81.465 201.445 ;
        RECT 81.645 200.855 81.975 201.615 ;
        RECT 81.295 200.515 81.960 200.685 ;
        RECT 82.145 200.540 82.415 201.445 ;
        RECT 65.000 199.715 71.745 199.885 ;
        RECT 72.005 199.745 72.320 200.305 ;
        RECT 72.490 200.055 79.610 200.305 ;
        RECT 64.570 199.065 64.830 199.625 ;
        RECT 65.000 199.260 65.260 199.715 ;
        RECT 65.430 199.065 65.690 199.545 ;
        RECT 65.860 199.260 66.120 199.715 ;
        RECT 66.290 199.065 66.550 199.545 ;
        RECT 66.720 199.260 66.980 199.715 ;
        RECT 67.150 199.065 67.395 199.545 ;
        RECT 67.565 199.260 67.840 199.715 ;
        RECT 68.010 199.065 68.255 199.545 ;
        RECT 68.425 199.260 68.685 199.715 ;
        RECT 68.865 199.065 69.115 199.545 ;
        RECT 69.285 199.260 69.545 199.715 ;
        RECT 69.725 199.065 69.975 199.545 ;
        RECT 70.145 199.260 70.405 199.715 ;
        RECT 70.585 199.065 70.845 199.545 ;
        RECT 71.015 199.260 71.275 199.715 ;
        RECT 71.445 199.065 71.745 199.545 ;
        RECT 72.005 199.065 72.310 199.575 ;
        RECT 72.490 199.245 72.740 200.055 ;
        RECT 72.910 199.065 73.170 199.590 ;
        RECT 73.350 199.245 73.600 200.055 ;
        RECT 79.780 199.885 80.945 200.475 ;
        RECT 81.790 200.370 81.960 200.515 ;
        RECT 81.225 199.965 81.555 200.335 ;
        RECT 81.790 200.040 82.075 200.370 ;
        RECT 74.200 199.715 80.945 199.885 ;
        RECT 81.790 199.785 81.960 200.040 ;
        RECT 73.770 199.065 74.030 199.625 ;
        RECT 74.200 199.260 74.460 199.715 ;
        RECT 74.630 199.065 74.890 199.545 ;
        RECT 75.060 199.260 75.320 199.715 ;
        RECT 75.490 199.065 75.750 199.545 ;
        RECT 75.920 199.260 76.180 199.715 ;
        RECT 76.350 199.065 76.595 199.545 ;
        RECT 76.765 199.260 77.040 199.715 ;
        RECT 77.210 199.065 77.455 199.545 ;
        RECT 77.625 199.260 77.885 199.715 ;
        RECT 78.065 199.065 78.315 199.545 ;
        RECT 78.485 199.260 78.745 199.715 ;
        RECT 78.925 199.065 79.175 199.545 ;
        RECT 79.345 199.260 79.605 199.715 ;
        RECT 79.785 199.065 80.045 199.545 ;
        RECT 80.215 199.260 80.475 199.715 ;
        RECT 81.295 199.615 81.960 199.785 ;
        RECT 82.245 199.740 82.415 200.540 ;
        RECT 82.585 200.450 82.875 201.615 ;
        RECT 83.045 200.475 83.375 201.615 ;
        RECT 83.545 200.985 83.900 201.445 ;
        RECT 84.070 201.155 84.645 201.615 ;
        RECT 84.815 200.985 85.145 201.445 ;
        RECT 83.545 200.815 85.145 200.985 ;
        RECT 85.345 200.815 85.600 201.615 ;
        RECT 83.545 200.475 83.820 200.815 ;
        RECT 84.000 200.255 84.190 200.635 ;
        RECT 83.045 200.055 84.190 200.255 ;
        RECT 84.370 199.915 84.650 200.815 ;
        RECT 85.770 200.645 86.070 200.840 ;
        RECT 84.820 200.475 86.070 200.645 ;
        RECT 86.355 200.685 86.525 201.445 ;
        RECT 86.740 200.855 87.070 201.615 ;
        RECT 86.355 200.515 87.070 200.685 ;
        RECT 87.240 200.540 87.495 201.445 ;
        RECT 84.820 200.055 85.150 200.475 ;
        RECT 85.380 199.975 85.725 200.305 ;
        RECT 84.370 199.885 84.655 199.915 ;
        RECT 80.645 199.065 80.945 199.545 ;
        RECT 81.295 199.235 81.465 199.615 ;
        RECT 81.645 199.065 81.975 199.445 ;
        RECT 82.155 199.235 82.415 199.740 ;
        RECT 82.585 199.065 82.875 199.790 ;
        RECT 83.045 199.675 84.155 199.885 ;
        RECT 83.045 199.235 83.395 199.675 ;
        RECT 83.565 199.065 83.735 199.505 ;
        RECT 83.905 199.445 84.155 199.675 ;
        RECT 84.325 199.615 84.655 199.885 ;
        RECT 84.825 199.445 85.100 199.885 ;
        RECT 85.900 199.820 86.070 200.475 ;
        RECT 86.265 199.965 86.620 200.335 ;
        RECT 86.900 200.305 87.070 200.515 ;
        RECT 86.900 199.975 87.155 200.305 ;
        RECT 83.905 199.235 85.100 199.445 ;
        RECT 85.335 199.065 85.665 199.805 ;
        RECT 85.835 199.490 86.070 199.820 ;
        RECT 86.900 199.785 87.070 199.975 ;
        RECT 87.325 199.810 87.495 200.540 ;
        RECT 87.670 200.465 87.930 201.615 ;
        RECT 88.105 200.525 89.315 201.615 ;
        RECT 88.105 199.985 88.625 200.525 ;
        RECT 86.355 199.615 87.070 199.785 ;
        RECT 86.355 199.235 86.525 199.615 ;
        RECT 86.740 199.065 87.070 199.445 ;
        RECT 87.240 199.235 87.495 199.810 ;
        RECT 87.670 199.065 87.930 199.905 ;
        RECT 88.795 199.815 89.315 200.355 ;
        RECT 88.105 199.065 89.315 199.815 ;
        RECT 18.100 198.895 89.400 199.065 ;
        RECT 18.185 198.145 19.395 198.895 ;
        RECT 18.185 197.605 18.705 198.145 ;
        RECT 19.570 198.055 19.830 198.895 ;
        RECT 20.005 198.150 20.260 198.725 ;
        RECT 20.430 198.515 20.760 198.895 ;
        RECT 20.975 198.345 21.145 198.725 ;
        RECT 20.430 198.175 21.145 198.345 ;
        RECT 18.875 197.435 19.395 197.975 ;
        RECT 18.185 196.345 19.395 197.435 ;
        RECT 19.570 196.345 19.830 197.495 ;
        RECT 20.005 197.420 20.175 198.150 ;
        RECT 20.430 197.985 20.600 198.175 ;
        RECT 20.345 197.655 20.600 197.985 ;
        RECT 20.430 197.445 20.600 197.655 ;
        RECT 20.880 197.625 21.235 197.995 ;
        RECT 20.005 196.515 20.260 197.420 ;
        RECT 20.430 197.275 21.145 197.445 ;
        RECT 20.430 196.345 20.760 197.105 ;
        RECT 20.975 196.515 21.145 197.275 ;
        RECT 21.865 196.515 22.615 198.725 ;
        RECT 22.875 198.345 23.045 198.725 ;
        RECT 23.225 198.515 23.555 198.895 ;
        RECT 22.875 198.175 23.540 198.345 ;
        RECT 23.735 198.220 23.995 198.725 ;
        RECT 22.805 197.625 23.145 197.995 ;
        RECT 23.370 197.920 23.540 198.175 ;
        RECT 23.370 197.590 23.645 197.920 ;
        RECT 23.370 197.445 23.540 197.590 ;
        RECT 22.865 197.275 23.540 197.445 ;
        RECT 23.815 197.420 23.995 198.220 ;
        RECT 22.865 196.515 23.045 197.275 ;
        RECT 23.225 196.345 23.555 197.105 ;
        RECT 23.725 196.515 23.995 197.420 ;
        RECT 24.170 198.420 24.505 198.680 ;
        RECT 24.675 198.495 25.005 198.895 ;
        RECT 25.175 198.495 26.790 198.665 ;
        RECT 24.170 197.065 24.425 198.420 ;
        RECT 25.175 198.325 25.345 198.495 ;
        RECT 24.785 198.155 25.345 198.325 ;
        RECT 24.785 197.985 24.955 198.155 ;
        RECT 24.650 197.655 24.955 197.985 ;
        RECT 25.150 197.875 25.400 197.985 ;
        RECT 25.610 197.875 25.880 198.315 ;
        RECT 26.070 198.215 26.360 198.315 ;
        RECT 26.065 198.045 26.360 198.215 ;
        RECT 25.145 197.705 25.400 197.875 ;
        RECT 25.605 197.705 25.880 197.875 ;
        RECT 25.150 197.655 25.400 197.705 ;
        RECT 25.610 197.655 25.880 197.705 ;
        RECT 26.070 197.655 26.360 198.045 ;
        RECT 26.530 197.655 26.950 198.320 ;
        RECT 27.335 198.175 27.665 198.895 ;
        RECT 27.260 197.655 27.610 197.985 ;
        RECT 24.785 197.485 24.955 197.655 ;
        RECT 27.405 197.535 27.610 197.655 ;
        RECT 27.845 197.950 28.185 198.725 ;
        RECT 28.355 198.435 28.525 198.895 ;
        RECT 28.765 198.460 29.125 198.725 ;
        RECT 28.765 198.455 29.120 198.460 ;
        RECT 28.765 198.445 29.115 198.455 ;
        RECT 28.765 198.440 29.110 198.445 ;
        RECT 28.765 198.430 29.105 198.440 ;
        RECT 29.755 198.435 29.925 198.895 ;
        RECT 28.765 198.425 29.100 198.430 ;
        RECT 28.765 198.415 29.090 198.425 ;
        RECT 28.765 198.405 29.080 198.415 ;
        RECT 28.765 198.265 29.065 198.405 ;
        RECT 28.355 198.075 29.065 198.265 ;
        RECT 29.255 198.265 29.585 198.345 ;
        RECT 30.095 198.265 30.435 198.725 ;
        RECT 29.255 198.075 30.435 198.265 ;
        RECT 30.640 198.155 31.255 198.725 ;
        RECT 31.425 198.385 31.640 198.895 ;
        RECT 31.870 198.385 32.150 198.715 ;
        RECT 32.330 198.385 32.570 198.895 ;
        RECT 24.785 197.315 27.155 197.485 ;
        RECT 27.405 197.365 27.615 197.535 ;
        RECT 24.170 196.555 24.505 197.065 ;
        RECT 24.755 196.345 25.085 197.145 ;
        RECT 25.330 196.935 26.755 197.105 ;
        RECT 25.330 196.515 25.615 196.935 ;
        RECT 25.870 196.345 26.200 196.765 ;
        RECT 26.425 196.685 26.755 196.935 ;
        RECT 26.985 196.855 27.155 197.315 ;
        RECT 27.415 196.685 27.585 197.185 ;
        RECT 26.425 196.515 27.585 196.685 ;
        RECT 27.845 196.515 28.125 197.950 ;
        RECT 28.355 197.505 28.640 198.075 ;
        RECT 28.825 197.675 29.295 197.905 ;
        RECT 29.465 197.885 29.795 197.905 ;
        RECT 29.465 197.705 29.915 197.885 ;
        RECT 30.105 197.705 30.435 197.905 ;
        RECT 28.355 197.290 29.505 197.505 ;
        RECT 28.295 196.345 29.005 197.120 ;
        RECT 29.175 196.515 29.505 197.290 ;
        RECT 29.700 196.590 29.915 197.705 ;
        RECT 30.205 197.365 30.435 197.705 ;
        RECT 30.640 197.135 30.955 198.155 ;
        RECT 31.125 197.485 31.295 197.985 ;
        RECT 31.545 197.655 31.810 198.215 ;
        RECT 31.980 197.485 32.150 198.385 ;
        RECT 32.320 197.655 32.675 198.215 ;
        RECT 32.910 198.130 33.365 198.895 ;
        RECT 33.640 198.515 34.940 198.725 ;
        RECT 35.195 198.535 35.525 198.895 ;
        RECT 34.770 198.365 34.940 198.515 ;
        RECT 35.695 198.395 35.955 198.725 ;
        RECT 33.840 197.905 34.060 198.305 ;
        RECT 32.905 197.705 33.395 197.905 ;
        RECT 33.585 197.695 34.060 197.905 ;
        RECT 34.305 197.905 34.515 198.305 ;
        RECT 34.770 198.240 35.525 198.365 ;
        RECT 34.770 198.195 35.615 198.240 ;
        RECT 35.345 198.075 35.615 198.195 ;
        RECT 34.305 197.695 34.635 197.905 ;
        RECT 34.805 197.635 35.215 197.940 ;
        RECT 31.125 197.315 32.550 197.485 ;
        RECT 30.095 196.345 30.425 197.065 ;
        RECT 30.640 196.515 31.175 197.135 ;
        RECT 31.345 196.345 31.675 197.145 ;
        RECT 32.160 197.140 32.550 197.315 ;
        RECT 32.910 197.465 34.085 197.525 ;
        RECT 35.445 197.500 35.615 198.075 ;
        RECT 35.415 197.465 35.615 197.500 ;
        RECT 32.910 197.355 35.615 197.465 ;
        RECT 32.910 196.735 33.165 197.355 ;
        RECT 33.755 197.295 35.555 197.355 ;
        RECT 33.755 197.265 34.085 197.295 ;
        RECT 35.785 197.195 35.955 198.395 ;
        RECT 33.415 197.095 33.600 197.185 ;
        RECT 34.190 197.095 35.025 197.105 ;
        RECT 33.415 196.895 35.025 197.095 ;
        RECT 33.415 196.855 33.645 196.895 ;
        RECT 32.910 196.515 33.245 196.735 ;
        RECT 34.250 196.345 34.605 196.725 ;
        RECT 34.775 196.515 35.025 196.895 ;
        RECT 35.275 196.345 35.525 197.125 ;
        RECT 35.695 196.515 35.955 197.195 ;
        RECT 36.125 198.395 36.385 198.725 ;
        RECT 36.555 198.535 36.885 198.895 ;
        RECT 37.140 198.515 38.440 198.725 ;
        RECT 36.125 197.195 36.295 198.395 ;
        RECT 37.140 198.365 37.310 198.515 ;
        RECT 36.555 198.240 37.310 198.365 ;
        RECT 36.465 198.195 37.310 198.240 ;
        RECT 36.465 198.075 36.735 198.195 ;
        RECT 36.465 197.500 36.635 198.075 ;
        RECT 36.865 197.635 37.275 197.940 ;
        RECT 37.565 197.905 37.775 198.305 ;
        RECT 37.445 197.695 37.775 197.905 ;
        RECT 38.020 197.905 38.240 198.305 ;
        RECT 38.715 198.130 39.170 198.895 ;
        RECT 39.345 198.095 40.040 198.725 ;
        RECT 40.245 198.095 40.555 198.895 ;
        RECT 40.735 198.170 41.065 198.680 ;
        RECT 41.235 198.495 41.565 198.895 ;
        RECT 42.615 198.325 42.945 198.665 ;
        RECT 43.115 198.495 43.445 198.895 ;
        RECT 38.020 197.695 38.495 197.905 ;
        RECT 38.685 197.705 39.175 197.905 ;
        RECT 39.365 197.655 39.700 197.905 ;
        RECT 36.465 197.465 36.665 197.500 ;
        RECT 37.995 197.465 39.170 197.525 ;
        RECT 39.870 197.495 40.040 198.095 ;
        RECT 40.210 197.655 40.545 197.925 ;
        RECT 36.465 197.355 39.170 197.465 ;
        RECT 36.525 197.295 38.325 197.355 ;
        RECT 37.995 197.265 38.325 197.295 ;
        RECT 36.125 196.515 36.385 197.195 ;
        RECT 36.555 196.345 36.805 197.125 ;
        RECT 37.055 197.095 37.890 197.105 ;
        RECT 38.480 197.095 38.665 197.185 ;
        RECT 37.055 196.895 38.665 197.095 ;
        RECT 37.055 196.515 37.305 196.895 ;
        RECT 38.435 196.855 38.665 196.895 ;
        RECT 38.915 196.735 39.170 197.355 ;
        RECT 37.475 196.345 37.830 196.725 ;
        RECT 38.835 196.515 39.170 196.735 ;
        RECT 39.345 196.345 39.605 197.485 ;
        RECT 39.775 196.515 40.105 197.495 ;
        RECT 40.275 196.345 40.555 197.485 ;
        RECT 40.735 197.405 40.925 198.170 ;
        RECT 41.235 198.155 43.600 198.325 ;
        RECT 43.945 198.170 44.235 198.895 ;
        RECT 41.235 197.985 41.405 198.155 ;
        RECT 41.095 197.655 41.405 197.985 ;
        RECT 41.575 197.655 41.880 197.985 ;
        RECT 40.735 196.555 41.065 197.405 ;
        RECT 41.235 196.345 41.485 197.485 ;
        RECT 41.665 197.325 41.880 197.655 ;
        RECT 42.055 197.325 42.340 197.985 ;
        RECT 42.535 197.325 42.800 197.985 ;
        RECT 43.015 197.325 43.260 197.985 ;
        RECT 43.430 197.155 43.600 198.155 ;
        RECT 44.405 198.155 44.725 198.530 ;
        RECT 44.980 198.155 45.150 198.895 ;
        RECT 45.400 198.325 45.570 198.530 ;
        RECT 45.815 198.495 46.170 198.895 ;
        RECT 46.345 198.325 46.515 198.675 ;
        RECT 46.715 198.495 47.045 198.895 ;
        RECT 47.215 198.325 47.385 198.675 ;
        RECT 47.555 198.495 47.935 198.895 ;
        RECT 45.400 198.155 45.920 198.325 ;
        RECT 46.345 198.155 47.955 198.325 ;
        RECT 48.125 198.220 48.400 198.565 ;
        RECT 41.675 196.985 42.965 197.155 ;
        RECT 41.675 196.565 41.925 196.985 ;
        RECT 42.155 196.345 42.485 196.815 ;
        RECT 42.715 196.565 42.965 196.985 ;
        RECT 43.145 196.985 43.600 197.155 ;
        RECT 43.145 196.555 43.475 196.985 ;
        RECT 43.945 196.345 44.235 197.510 ;
        RECT 44.405 197.115 44.580 198.155 ;
        RECT 44.750 197.285 45.100 197.985 ;
        RECT 45.270 197.655 45.560 197.985 ;
        RECT 45.730 197.905 45.920 198.155 ;
        RECT 47.785 197.985 47.955 198.155 ;
        RECT 45.730 197.735 46.175 197.905 ;
        RECT 45.730 197.455 45.920 197.735 ;
        RECT 46.570 197.565 46.740 197.985 ;
        RECT 46.960 197.655 47.615 197.985 ;
        RECT 47.785 197.655 48.060 197.985 ;
        RECT 45.315 197.285 45.920 197.455 ;
        RECT 46.090 197.395 46.740 197.565 ;
        RECT 47.785 197.485 47.955 197.655 ;
        RECT 48.230 197.485 48.400 198.220 ;
        RECT 48.570 197.955 48.740 198.895 ;
        RECT 49.015 198.555 49.350 198.725 ;
        RECT 49.015 198.155 49.630 198.555 ;
        RECT 50.310 198.515 50.645 198.895 ;
        RECT 51.235 198.455 51.470 198.895 ;
        RECT 51.640 198.365 51.970 198.725 ;
        RECT 52.140 198.535 52.470 198.895 ;
        RECT 52.685 198.385 52.990 198.895 ;
        RECT 49.800 198.155 51.070 198.345 ;
        RECT 51.640 198.195 52.460 198.365 ;
        RECT 49.005 197.655 49.280 197.985 ;
        RECT 46.090 197.115 46.260 197.395 ;
        RECT 47.295 197.315 47.955 197.485 ;
        RECT 47.295 197.195 47.465 197.315 ;
        RECT 44.405 196.945 46.260 197.115 ;
        RECT 46.430 197.025 47.465 197.195 ;
        RECT 44.405 196.525 44.665 196.945 ;
        RECT 46.430 196.775 46.600 197.025 ;
        RECT 44.835 196.345 45.165 196.775 ;
        RECT 45.855 196.605 46.600 196.775 ;
        RECT 46.825 196.525 47.465 196.855 ;
        RECT 47.635 196.345 47.915 197.145 ;
        RECT 48.125 196.515 48.400 197.485 ;
        RECT 48.570 196.345 48.740 197.540 ;
        RECT 49.450 197.470 49.630 198.155 ;
        RECT 49.800 197.655 50.160 197.985 ;
        RECT 50.450 197.875 50.740 197.985 ;
        RECT 50.445 197.705 50.740 197.875 ;
        RECT 50.450 197.655 50.740 197.705 ;
        RECT 50.910 197.655 51.245 197.985 ;
        RECT 51.415 197.655 52.095 197.985 ;
        RECT 51.415 197.470 51.585 197.655 ;
        RECT 49.010 197.215 51.585 197.470 ;
        RECT 49.010 196.515 49.275 197.215 ;
        RECT 49.445 196.345 49.775 197.045 ;
        RECT 49.945 196.515 50.615 197.215 ;
        RECT 52.265 197.075 52.460 198.195 ;
        RECT 52.685 197.655 53.000 198.215 ;
        RECT 53.170 197.905 53.420 198.715 ;
        RECT 53.590 198.370 53.850 198.895 ;
        RECT 54.030 197.905 54.280 198.715 ;
        RECT 54.450 198.335 54.710 198.895 ;
        RECT 54.880 198.245 55.140 198.700 ;
        RECT 55.310 198.415 55.570 198.895 ;
        RECT 55.740 198.245 56.000 198.700 ;
        RECT 56.170 198.415 56.430 198.895 ;
        RECT 56.600 198.245 56.860 198.700 ;
        RECT 57.030 198.415 57.275 198.895 ;
        RECT 57.445 198.245 57.720 198.700 ;
        RECT 57.890 198.415 58.135 198.895 ;
        RECT 58.305 198.245 58.565 198.700 ;
        RECT 58.745 198.415 58.995 198.895 ;
        RECT 59.165 198.245 59.425 198.700 ;
        RECT 59.605 198.415 59.855 198.895 ;
        RECT 60.025 198.245 60.285 198.700 ;
        RECT 60.465 198.415 60.725 198.895 ;
        RECT 60.895 198.245 61.155 198.700 ;
        RECT 61.325 198.415 61.625 198.895 ;
        RECT 61.885 198.555 63.245 198.725 ;
        RECT 54.880 198.075 61.625 198.245 ;
        RECT 61.885 198.075 62.245 198.555 ;
        RECT 62.415 198.155 62.745 198.385 ;
        RECT 62.915 198.325 63.245 198.555 ;
        RECT 63.415 198.495 63.745 198.895 ;
        RECT 63.915 198.325 64.245 198.725 ;
        RECT 62.915 198.155 64.245 198.325 ;
        RECT 64.515 198.155 64.845 198.895 ;
        RECT 53.170 197.655 60.290 197.905 ;
        RECT 51.120 196.345 51.550 197.045 ;
        RECT 51.730 196.905 52.460 197.075 ;
        RECT 51.730 196.515 51.920 196.905 ;
        RECT 52.090 196.345 52.420 196.725 ;
        RECT 52.695 196.345 52.990 197.155 ;
        RECT 53.170 196.515 53.415 197.655 ;
        RECT 53.590 196.345 53.850 197.155 ;
        RECT 54.030 196.520 54.280 197.655 ;
        RECT 60.460 197.485 61.625 198.075 ;
        RECT 61.885 197.735 62.245 197.905 ;
        RECT 61.885 197.655 62.215 197.735 ;
        RECT 54.880 197.260 61.625 197.485 ;
        RECT 54.880 197.245 60.285 197.260 ;
        RECT 54.450 196.350 54.710 197.145 ;
        RECT 54.880 196.520 55.140 197.245 ;
        RECT 55.310 196.350 55.570 197.075 ;
        RECT 55.740 196.520 56.000 197.245 ;
        RECT 56.170 196.350 56.430 197.075 ;
        RECT 56.600 196.520 56.860 197.245 ;
        RECT 57.030 196.350 57.290 197.075 ;
        RECT 57.460 196.520 57.720 197.245 ;
        RECT 57.890 196.350 58.135 197.075 ;
        RECT 58.305 196.520 58.565 197.245 ;
        RECT 58.750 196.350 58.995 197.075 ;
        RECT 59.165 196.520 59.425 197.245 ;
        RECT 59.610 196.350 59.855 197.075 ;
        RECT 60.025 196.520 60.285 197.245 ;
        RECT 60.470 196.350 60.725 197.075 ;
        RECT 60.895 196.520 61.185 197.260 ;
        RECT 54.450 196.345 60.725 196.350 ;
        RECT 61.355 196.345 61.625 197.090 ;
        RECT 61.885 196.345 62.245 197.485 ;
        RECT 62.415 197.195 62.615 198.155 ;
        RECT 62.785 197.875 63.030 197.985 ;
        RECT 62.785 197.705 63.035 197.875 ;
        RECT 62.785 197.365 63.030 197.705 ;
        RECT 63.305 197.365 63.525 197.985 ;
        RECT 63.780 197.365 63.955 197.985 ;
        RECT 64.225 197.365 64.445 197.985 ;
        RECT 64.615 197.195 64.925 197.985 ;
        RECT 62.415 197.025 64.925 197.195 ;
        RECT 62.915 196.515 63.245 197.025 ;
        RECT 64.415 196.345 64.925 196.855 ;
        RECT 65.095 196.515 65.425 198.725 ;
        RECT 65.595 198.095 65.855 198.895 ;
        RECT 66.205 198.515 66.535 198.895 ;
        RECT 66.705 198.345 66.895 198.725 ;
        RECT 67.065 198.535 67.395 198.895 ;
        RECT 66.495 198.155 66.895 198.345 ;
        RECT 67.615 198.325 67.805 198.725 ;
        RECT 67.065 198.155 67.805 198.325 ;
        RECT 65.595 196.345 65.855 197.485 ;
        RECT 66.035 196.345 66.325 197.315 ;
        RECT 66.495 196.515 66.725 198.155 ;
        RECT 67.065 197.985 67.235 198.155 ;
        RECT 66.895 197.290 67.235 197.985 ;
        RECT 67.405 197.570 67.730 197.985 ;
        RECT 68.180 197.655 68.560 198.615 ;
        RECT 68.745 198.415 69.075 198.895 ;
        RECT 68.750 197.655 69.065 198.230 ;
        RECT 69.705 198.170 69.995 198.895 ;
        RECT 70.165 198.385 70.470 198.895 ;
        RECT 70.165 197.655 70.480 198.215 ;
        RECT 70.650 197.905 70.900 198.715 ;
        RECT 71.070 198.370 71.330 198.895 ;
        RECT 71.510 197.905 71.760 198.715 ;
        RECT 71.930 198.335 72.190 198.895 ;
        RECT 72.360 198.245 72.620 198.700 ;
        RECT 72.790 198.415 73.050 198.895 ;
        RECT 73.220 198.245 73.480 198.700 ;
        RECT 73.650 198.415 73.910 198.895 ;
        RECT 74.080 198.245 74.340 198.700 ;
        RECT 74.510 198.415 74.755 198.895 ;
        RECT 74.925 198.245 75.200 198.700 ;
        RECT 75.370 198.415 75.615 198.895 ;
        RECT 75.785 198.245 76.045 198.700 ;
        RECT 76.225 198.415 76.475 198.895 ;
        RECT 76.645 198.245 76.905 198.700 ;
        RECT 77.085 198.415 77.335 198.895 ;
        RECT 77.505 198.245 77.765 198.700 ;
        RECT 77.945 198.415 78.205 198.895 ;
        RECT 78.375 198.245 78.635 198.700 ;
        RECT 78.805 198.415 79.105 198.895 ;
        RECT 72.360 198.075 79.105 198.245 ;
        RECT 79.365 198.075 79.660 198.895 ;
        RECT 79.830 198.155 80.270 198.715 ;
        RECT 80.440 198.155 80.890 198.895 ;
        RECT 81.060 198.325 81.230 198.725 ;
        RECT 81.400 198.495 81.820 198.895 ;
        RECT 81.990 198.325 82.220 198.725 ;
        RECT 81.060 198.155 82.220 198.325 ;
        RECT 82.390 198.155 82.875 198.725 ;
        RECT 70.650 197.655 77.770 197.905 ;
        RECT 66.895 197.060 67.730 197.290 ;
        RECT 66.895 196.345 67.225 196.760 ;
        RECT 67.415 196.515 67.730 197.060 ;
        RECT 67.900 197.045 69.015 197.310 ;
        RECT 67.900 196.515 68.125 197.045 ;
        RECT 68.295 196.345 68.625 196.855 ;
        RECT 68.795 196.515 69.015 197.045 ;
        RECT 69.705 196.345 69.995 197.510 ;
        RECT 70.175 196.345 70.470 197.155 ;
        RECT 70.650 196.515 70.895 197.655 ;
        RECT 71.070 196.345 71.330 197.155 ;
        RECT 71.510 196.520 71.760 197.655 ;
        RECT 77.940 197.485 79.105 198.075 ;
        RECT 79.830 197.905 80.140 198.155 ;
        RECT 79.365 197.685 80.140 197.905 ;
        RECT 72.360 197.260 79.105 197.485 ;
        RECT 72.360 197.245 77.765 197.260 ;
        RECT 71.930 196.350 72.190 197.145 ;
        RECT 72.360 196.520 72.620 197.245 ;
        RECT 72.790 196.350 73.050 197.075 ;
        RECT 73.220 196.520 73.480 197.245 ;
        RECT 73.650 196.350 73.910 197.075 ;
        RECT 74.080 196.520 74.340 197.245 ;
        RECT 74.510 196.350 74.770 197.075 ;
        RECT 74.940 196.520 75.200 197.245 ;
        RECT 75.370 196.350 75.615 197.075 ;
        RECT 75.785 196.520 76.045 197.245 ;
        RECT 76.230 196.350 76.475 197.075 ;
        RECT 76.645 196.520 76.905 197.245 ;
        RECT 77.090 196.350 77.335 197.075 ;
        RECT 77.505 196.520 77.765 197.245 ;
        RECT 77.950 196.350 78.205 197.075 ;
        RECT 78.375 196.520 78.665 197.260 ;
        RECT 71.930 196.345 78.205 196.350 ;
        RECT 78.835 196.345 79.105 197.090 ;
        RECT 79.365 196.345 79.660 197.515 ;
        RECT 79.830 197.145 80.140 197.685 ;
        RECT 80.310 197.535 80.480 197.985 ;
        RECT 80.650 197.705 81.040 197.985 ;
        RECT 81.225 197.655 81.470 197.985 ;
        RECT 80.310 197.365 81.100 197.535 ;
        RECT 79.830 196.515 80.270 197.145 ;
        RECT 80.445 196.345 80.760 197.195 ;
        RECT 80.930 196.685 81.100 197.365 ;
        RECT 81.270 196.855 81.470 197.655 ;
        RECT 81.670 196.855 81.920 197.985 ;
        RECT 82.135 197.655 82.535 197.985 ;
        RECT 82.705 197.485 82.875 198.155 ;
        RECT 83.045 198.075 83.340 198.895 ;
        RECT 83.510 198.155 83.950 198.715 ;
        RECT 84.120 198.155 84.570 198.895 ;
        RECT 84.740 198.325 84.910 198.725 ;
        RECT 85.080 198.495 85.500 198.895 ;
        RECT 85.670 198.325 85.900 198.725 ;
        RECT 84.740 198.155 85.900 198.325 ;
        RECT 86.070 198.155 86.555 198.725 ;
        RECT 83.510 197.905 83.820 198.155 ;
        RECT 83.045 197.685 83.820 197.905 ;
        RECT 82.110 197.315 82.875 197.485 ;
        RECT 82.110 196.685 82.360 197.315 ;
        RECT 80.930 196.515 82.360 196.685 ;
        RECT 82.535 196.345 82.870 197.145 ;
        RECT 83.045 196.345 83.340 197.515 ;
        RECT 83.510 197.145 83.820 197.685 ;
        RECT 83.990 197.535 84.160 197.985 ;
        RECT 84.330 197.705 84.720 197.985 ;
        RECT 84.905 197.655 85.150 197.985 ;
        RECT 83.990 197.365 84.780 197.535 ;
        RECT 83.510 196.515 83.950 197.145 ;
        RECT 84.125 196.345 84.440 197.195 ;
        RECT 84.610 196.685 84.780 197.365 ;
        RECT 84.950 196.855 85.150 197.655 ;
        RECT 85.350 196.855 85.600 197.985 ;
        RECT 85.815 197.655 86.215 197.985 ;
        RECT 86.385 197.485 86.555 198.155 ;
        RECT 85.790 197.315 86.555 197.485 ;
        RECT 86.725 198.220 86.985 198.725 ;
        RECT 87.165 198.515 87.495 198.895 ;
        RECT 87.675 198.345 87.845 198.725 ;
        RECT 86.725 197.420 86.905 198.220 ;
        RECT 87.180 198.175 87.845 198.345 ;
        RECT 87.180 197.920 87.350 198.175 ;
        RECT 88.105 198.145 89.315 198.895 ;
        RECT 87.075 197.590 87.350 197.920 ;
        RECT 87.575 197.625 87.915 197.995 ;
        RECT 87.180 197.445 87.350 197.590 ;
        RECT 85.790 196.685 86.040 197.315 ;
        RECT 84.610 196.515 86.040 196.685 ;
        RECT 86.215 196.345 86.550 197.145 ;
        RECT 86.725 196.515 86.995 197.420 ;
        RECT 87.180 197.275 87.855 197.445 ;
        RECT 87.165 196.345 87.495 197.105 ;
        RECT 87.675 196.515 87.855 197.275 ;
        RECT 88.105 197.435 88.625 197.975 ;
        RECT 88.795 197.605 89.315 198.145 ;
        RECT 88.105 196.345 89.315 197.435 ;
        RECT 18.100 196.175 89.400 196.345 ;
        RECT 18.185 195.085 19.395 196.175 ;
        RECT 18.185 194.375 18.705 194.915 ;
        RECT 18.875 194.545 19.395 195.085 ;
        RECT 20.025 195.035 20.315 196.175 ;
        RECT 20.485 195.455 20.935 196.005 ;
        RECT 21.125 195.455 21.455 196.175 ;
        RECT 18.185 193.625 19.395 194.375 ;
        RECT 20.025 193.625 20.315 194.425 ;
        RECT 20.485 194.085 20.735 195.455 ;
        RECT 21.665 195.285 21.965 195.835 ;
        RECT 22.135 195.505 22.415 196.175 ;
        RECT 21.025 195.115 21.965 195.285 ;
        RECT 21.025 194.865 21.195 195.115 ;
        RECT 22.300 194.865 22.615 195.305 ;
        RECT 22.970 195.205 23.360 195.380 ;
        RECT 23.845 195.375 24.175 196.175 ;
        RECT 24.345 195.385 24.880 196.005 ;
        RECT 22.970 195.035 24.395 195.205 ;
        RECT 20.905 194.535 21.195 194.865 ;
        RECT 21.365 194.615 21.695 194.865 ;
        RECT 21.925 194.615 22.615 194.865 ;
        RECT 21.025 194.445 21.195 194.535 ;
        RECT 21.025 194.255 22.415 194.445 ;
        RECT 22.845 194.305 23.200 194.865 ;
        RECT 20.485 193.795 21.035 194.085 ;
        RECT 21.205 193.625 21.455 194.085 ;
        RECT 22.085 193.895 22.415 194.255 ;
        RECT 23.370 194.135 23.540 195.035 ;
        RECT 23.710 194.305 23.975 194.865 ;
        RECT 24.225 194.535 24.395 195.035 ;
        RECT 24.565 194.365 24.880 195.385 ;
        RECT 25.175 195.835 26.335 196.005 ;
        RECT 25.175 195.335 25.345 195.835 ;
        RECT 25.605 195.205 25.775 195.665 ;
        RECT 26.005 195.585 26.335 195.835 ;
        RECT 26.560 195.755 26.890 196.175 ;
        RECT 27.145 195.585 27.430 196.005 ;
        RECT 26.005 195.415 27.430 195.585 ;
        RECT 27.675 195.375 28.005 196.175 ;
        RECT 28.255 195.455 28.590 195.965 ;
        RECT 25.150 194.865 25.355 195.155 ;
        RECT 25.605 195.035 27.975 195.205 ;
        RECT 27.805 194.865 27.975 195.035 ;
        RECT 25.150 194.815 25.500 194.865 ;
        RECT 25.145 194.645 25.500 194.815 ;
        RECT 25.150 194.535 25.500 194.645 ;
        RECT 22.950 193.625 23.190 194.135 ;
        RECT 23.370 193.805 23.650 194.135 ;
        RECT 23.880 193.625 24.095 194.135 ;
        RECT 24.265 193.795 24.880 194.365 ;
        RECT 25.095 193.625 25.425 194.345 ;
        RECT 25.810 194.200 26.230 194.865 ;
        RECT 26.400 194.205 26.690 194.865 ;
        RECT 26.880 194.815 27.150 194.865 ;
        RECT 27.360 194.815 27.610 194.865 ;
        RECT 26.880 194.645 27.155 194.815 ;
        RECT 27.360 194.645 27.615 194.815 ;
        RECT 26.880 194.205 27.150 194.645 ;
        RECT 27.360 194.535 27.610 194.645 ;
        RECT 27.805 194.535 28.110 194.865 ;
        RECT 27.805 194.365 27.975 194.535 ;
        RECT 27.415 194.195 27.975 194.365 ;
        RECT 27.415 194.025 27.585 194.195 ;
        RECT 28.335 194.100 28.590 195.455 ;
        RECT 25.970 193.855 27.585 194.025 ;
        RECT 27.755 193.625 28.085 194.025 ;
        RECT 28.255 193.840 28.590 194.100 ;
        RECT 29.685 195.100 29.955 196.005 ;
        RECT 30.125 195.415 30.455 196.175 ;
        RECT 30.635 195.245 30.805 196.005 ;
        RECT 29.685 194.300 29.855 195.100 ;
        RECT 30.140 195.075 30.805 195.245 ;
        RECT 30.140 194.930 30.310 195.075 ;
        RECT 31.065 195.010 31.355 196.175 ;
        RECT 31.525 195.035 31.785 196.175 ;
        RECT 31.955 195.025 32.285 196.005 ;
        RECT 32.455 195.035 32.735 196.175 ;
        RECT 32.910 195.035 33.230 196.175 ;
        RECT 30.025 194.600 30.310 194.930 ;
        RECT 30.140 194.345 30.310 194.600 ;
        RECT 30.545 194.525 30.875 194.895 ;
        RECT 31.545 194.615 31.880 194.865 ;
        RECT 32.050 194.425 32.220 195.025 ;
        RECT 33.410 194.865 33.605 195.915 ;
        RECT 33.785 195.325 34.115 196.005 ;
        RECT 34.315 195.375 34.570 196.175 ;
        RECT 33.785 195.045 34.135 195.325 ;
        RECT 32.390 194.595 32.725 194.865 ;
        RECT 32.970 194.815 33.230 194.865 ;
        RECT 32.965 194.645 33.230 194.815 ;
        RECT 32.970 194.535 33.230 194.645 ;
        RECT 33.410 194.535 33.795 194.865 ;
        RECT 33.965 194.665 34.135 195.045 ;
        RECT 34.325 194.835 34.570 195.195 ;
        RECT 34.900 195.165 35.200 196.005 ;
        RECT 35.395 195.335 35.645 196.175 ;
        RECT 36.235 195.585 37.040 196.005 ;
        RECT 35.815 195.415 37.380 195.585 ;
        RECT 35.815 195.165 35.985 195.415 ;
        RECT 34.900 194.995 35.985 195.165 ;
        RECT 33.965 194.495 34.485 194.665 ;
        RECT 34.745 194.535 35.075 194.825 ;
        RECT 29.685 193.795 29.945 194.300 ;
        RECT 30.140 194.175 30.805 194.345 ;
        RECT 30.125 193.625 30.455 194.005 ;
        RECT 30.635 193.795 30.805 194.175 ;
        RECT 31.065 193.625 31.355 194.350 ;
        RECT 31.525 193.795 32.220 194.425 ;
        RECT 32.425 193.625 32.735 194.425 ;
        RECT 32.910 194.155 34.125 194.325 ;
        RECT 32.910 193.805 33.200 194.155 ;
        RECT 33.395 193.625 33.725 193.985 ;
        RECT 33.895 193.850 34.125 194.155 ;
        RECT 34.315 193.930 34.485 194.495 ;
        RECT 35.245 194.365 35.415 194.995 ;
        RECT 36.155 194.865 36.475 195.245 ;
        RECT 35.585 194.615 35.915 194.825 ;
        RECT 36.095 194.615 36.475 194.865 ;
        RECT 36.665 194.825 37.040 195.245 ;
        RECT 37.210 195.165 37.380 195.415 ;
        RECT 37.550 195.335 37.880 196.175 ;
        RECT 38.050 195.415 38.715 196.005 ;
        RECT 37.210 194.995 38.130 195.165 ;
        RECT 37.960 194.825 38.130 194.995 ;
        RECT 36.665 194.815 37.150 194.825 ;
        RECT 36.645 194.645 37.150 194.815 ;
        RECT 36.665 194.615 37.150 194.645 ;
        RECT 37.340 194.615 37.790 194.825 ;
        RECT 37.960 194.615 38.295 194.825 ;
        RECT 38.465 194.445 38.715 195.415 ;
        RECT 39.350 195.785 39.685 196.005 ;
        RECT 40.690 195.795 41.045 196.175 ;
        RECT 39.350 195.165 39.605 195.785 ;
        RECT 39.855 195.625 40.085 195.665 ;
        RECT 41.215 195.625 41.465 196.005 ;
        RECT 39.855 195.425 41.465 195.625 ;
        RECT 39.855 195.335 40.040 195.425 ;
        RECT 40.630 195.415 41.465 195.425 ;
        RECT 41.715 195.395 41.965 196.175 ;
        RECT 42.135 195.325 42.395 196.005 ;
        RECT 42.655 195.430 42.925 196.175 ;
        RECT 43.555 196.170 49.830 196.175 ;
        RECT 40.195 195.225 40.525 195.255 ;
        RECT 40.195 195.165 41.995 195.225 ;
        RECT 39.350 195.055 42.055 195.165 ;
        RECT 39.350 194.995 40.525 195.055 ;
        RECT 41.855 195.020 42.055 195.055 ;
        RECT 39.345 194.615 39.835 194.815 ;
        RECT 40.025 194.615 40.500 194.825 ;
        RECT 34.905 194.185 35.415 194.365 ;
        RECT 35.820 194.275 37.520 194.445 ;
        RECT 35.820 194.185 36.205 194.275 ;
        RECT 34.905 193.795 35.235 194.185 ;
        RECT 35.405 193.845 36.590 194.015 ;
        RECT 36.850 193.625 37.020 194.095 ;
        RECT 37.190 193.810 37.520 194.275 ;
        RECT 37.690 193.625 37.860 194.445 ;
        RECT 38.030 193.805 38.715 194.445 ;
        RECT 39.350 193.625 39.805 194.390 ;
        RECT 40.280 194.215 40.500 194.615 ;
        RECT 40.745 194.615 41.075 194.825 ;
        RECT 40.745 194.215 40.955 194.615 ;
        RECT 41.245 194.580 41.655 194.885 ;
        RECT 41.885 194.445 42.055 195.020 ;
        RECT 41.785 194.325 42.055 194.445 ;
        RECT 41.210 194.280 42.055 194.325 ;
        RECT 41.210 194.155 41.965 194.280 ;
        RECT 41.210 194.005 41.380 194.155 ;
        RECT 42.225 194.125 42.395 195.325 ;
        RECT 43.095 195.260 43.385 196.000 ;
        RECT 43.555 195.445 43.810 196.170 ;
        RECT 43.995 195.275 44.255 196.000 ;
        RECT 44.425 195.445 44.670 196.170 ;
        RECT 44.855 195.275 45.115 196.000 ;
        RECT 45.285 195.445 45.530 196.170 ;
        RECT 45.715 195.275 45.975 196.000 ;
        RECT 46.145 195.445 46.390 196.170 ;
        RECT 46.560 195.275 46.820 196.000 ;
        RECT 46.990 195.445 47.250 196.170 ;
        RECT 47.420 195.275 47.680 196.000 ;
        RECT 47.850 195.445 48.110 196.170 ;
        RECT 48.280 195.275 48.540 196.000 ;
        RECT 48.710 195.445 48.970 196.170 ;
        RECT 49.140 195.275 49.400 196.000 ;
        RECT 49.570 195.375 49.830 196.170 ;
        RECT 43.995 195.260 49.400 195.275 ;
        RECT 42.655 195.035 49.400 195.260 ;
        RECT 42.655 194.445 43.820 195.035 ;
        RECT 50.000 194.865 50.250 196.000 ;
        RECT 50.430 195.365 50.690 196.175 ;
        RECT 50.865 194.865 51.110 196.005 ;
        RECT 51.290 195.365 51.585 196.175 ;
        RECT 51.765 195.035 52.025 196.175 ;
        RECT 43.990 194.615 51.110 194.865 ;
        RECT 42.655 194.275 49.400 194.445 ;
        RECT 40.080 193.795 41.380 194.005 ;
        RECT 41.635 193.625 41.965 193.985 ;
        RECT 42.135 193.795 42.395 194.125 ;
        RECT 42.655 193.625 42.955 194.105 ;
        RECT 43.125 193.820 43.385 194.275 ;
        RECT 43.555 193.625 43.815 194.105 ;
        RECT 43.995 193.820 44.255 194.275 ;
        RECT 44.425 193.625 44.675 194.105 ;
        RECT 44.855 193.820 45.115 194.275 ;
        RECT 45.285 193.625 45.535 194.105 ;
        RECT 45.715 193.820 45.975 194.275 ;
        RECT 46.145 193.625 46.390 194.105 ;
        RECT 46.560 193.820 46.835 194.275 ;
        RECT 47.005 193.625 47.250 194.105 ;
        RECT 47.420 193.820 47.680 194.275 ;
        RECT 47.850 193.625 48.110 194.105 ;
        RECT 48.280 193.820 48.540 194.275 ;
        RECT 48.710 193.625 48.970 194.105 ;
        RECT 49.140 193.820 49.400 194.275 ;
        RECT 49.570 193.625 49.830 194.185 ;
        RECT 50.000 193.805 50.250 194.615 ;
        RECT 50.430 193.625 50.690 194.150 ;
        RECT 50.860 193.805 51.110 194.615 ;
        RECT 51.280 194.305 51.595 194.865 ;
        RECT 51.290 193.625 51.595 194.135 ;
        RECT 51.765 193.625 52.025 194.425 ;
        RECT 52.195 193.795 52.525 196.005 ;
        RECT 52.695 195.665 53.205 196.175 ;
        RECT 54.375 195.495 54.705 196.005 ;
        RECT 52.695 195.325 55.205 195.495 ;
        RECT 52.695 194.535 53.005 195.325 ;
        RECT 53.175 194.535 53.395 195.155 ;
        RECT 53.665 194.535 53.840 195.155 ;
        RECT 54.095 194.535 54.315 195.155 ;
        RECT 54.585 194.985 54.835 195.155 ;
        RECT 54.590 194.535 54.835 194.985 ;
        RECT 55.005 194.365 55.205 195.325 ;
        RECT 55.375 195.035 55.735 196.175 ;
        RECT 56.825 195.010 57.115 196.175 ;
        RECT 57.375 195.430 57.645 196.175 ;
        RECT 58.275 196.170 64.550 196.175 ;
        RECT 57.815 195.260 58.105 196.000 ;
        RECT 58.275 195.445 58.530 196.170 ;
        RECT 58.715 195.275 58.975 196.000 ;
        RECT 59.145 195.445 59.390 196.170 ;
        RECT 59.575 195.275 59.835 196.000 ;
        RECT 60.005 195.445 60.250 196.170 ;
        RECT 60.435 195.275 60.695 196.000 ;
        RECT 60.865 195.445 61.110 196.170 ;
        RECT 61.280 195.275 61.540 196.000 ;
        RECT 61.710 195.445 61.970 196.170 ;
        RECT 62.140 195.275 62.400 196.000 ;
        RECT 62.570 195.445 62.830 196.170 ;
        RECT 63.000 195.275 63.260 196.000 ;
        RECT 63.430 195.445 63.690 196.170 ;
        RECT 63.860 195.275 64.120 196.000 ;
        RECT 64.290 195.375 64.550 196.170 ;
        RECT 58.715 195.260 64.120 195.275 ;
        RECT 57.375 195.035 64.120 195.260 ;
        RECT 55.405 194.785 55.735 194.865 ;
        RECT 55.375 194.615 55.735 194.785 ;
        RECT 57.375 194.475 58.540 195.035 ;
        RECT 64.720 194.865 64.970 196.000 ;
        RECT 65.150 195.365 65.410 196.175 ;
        RECT 65.585 194.865 65.830 196.005 ;
        RECT 66.010 195.365 66.305 196.175 ;
        RECT 66.575 195.205 66.745 196.005 ;
        RECT 67.035 195.545 67.285 195.965 ;
        RECT 67.475 195.715 67.805 196.175 ;
        RECT 68.015 195.545 68.265 195.965 ;
        RECT 66.975 195.375 68.265 195.545 ;
        RECT 68.435 195.375 68.685 196.175 ;
        RECT 68.855 195.545 69.025 196.005 ;
        RECT 69.235 195.715 69.485 196.175 ;
        RECT 68.855 195.375 69.530 195.545 ;
        RECT 66.575 195.035 69.065 195.205 ;
        RECT 58.710 194.615 65.830 194.865 ;
        RECT 57.345 194.445 58.540 194.475 ;
        RECT 52.775 193.625 53.105 194.365 ;
        RECT 53.375 194.195 54.705 194.365 ;
        RECT 53.375 193.795 53.705 194.195 ;
        RECT 53.875 193.625 54.205 194.025 ;
        RECT 54.375 193.965 54.705 194.195 ;
        RECT 54.875 194.135 55.205 194.365 ;
        RECT 55.375 193.965 55.735 194.445 ;
        RECT 54.375 193.795 55.735 193.965 ;
        RECT 56.825 193.625 57.115 194.350 ;
        RECT 57.345 194.305 64.120 194.445 ;
        RECT 57.375 194.275 64.120 194.305 ;
        RECT 57.375 193.625 57.675 194.105 ;
        RECT 57.845 193.820 58.105 194.275 ;
        RECT 58.275 193.625 58.535 194.105 ;
        RECT 58.715 193.820 58.975 194.275 ;
        RECT 59.145 193.625 59.395 194.105 ;
        RECT 59.575 193.820 59.835 194.275 ;
        RECT 60.005 193.625 60.255 194.105 ;
        RECT 60.435 193.820 60.695 194.275 ;
        RECT 60.865 193.625 61.110 194.105 ;
        RECT 61.280 193.820 61.555 194.275 ;
        RECT 61.725 193.625 61.970 194.105 ;
        RECT 62.140 193.820 62.400 194.275 ;
        RECT 62.570 193.625 62.830 194.105 ;
        RECT 63.000 193.820 63.260 194.275 ;
        RECT 63.430 193.625 63.690 194.105 ;
        RECT 63.860 193.820 64.120 194.275 ;
        RECT 64.290 193.625 64.550 194.185 ;
        RECT 64.720 193.805 64.970 194.615 ;
        RECT 65.150 193.625 65.410 194.150 ;
        RECT 65.580 193.805 65.830 194.615 ;
        RECT 66.000 194.305 66.315 194.865 ;
        RECT 66.530 194.295 66.725 194.865 ;
        RECT 66.010 193.625 66.315 194.135 ;
        RECT 66.485 193.625 66.745 194.105 ;
        RECT 66.915 194.045 67.085 195.035 ;
        RECT 67.265 194.410 67.435 194.865 ;
        RECT 67.825 194.785 67.995 194.800 ;
        RECT 67.665 194.615 67.995 194.785 ;
        RECT 67.265 194.240 67.655 194.410 ;
        RECT 66.915 193.875 67.245 194.045 ;
        RECT 67.445 193.955 67.655 194.240 ;
        RECT 67.825 194.405 67.995 194.615 ;
        RECT 68.225 194.535 68.555 194.865 ;
        RECT 68.895 194.785 69.065 195.035 ;
        RECT 68.735 194.615 69.065 194.785 ;
        RECT 67.825 194.235 68.090 194.405 ;
        RECT 68.350 194.300 68.555 194.535 ;
        RECT 69.275 194.425 69.530 195.375 ;
        RECT 69.710 195.030 70.005 196.175 ;
        RECT 67.920 194.135 68.090 194.235 ;
        RECT 68.855 194.255 69.530 194.425 ;
        RECT 67.920 193.965 68.095 194.135 ;
        RECT 68.435 194.005 68.605 194.085 ;
        RECT 67.920 193.940 68.090 193.965 ;
        RECT 66.915 193.795 67.160 193.875 ;
        RECT 68.335 193.625 68.665 194.005 ;
        RECT 68.855 193.795 69.025 194.255 ;
        RECT 69.275 193.625 69.530 194.085 ;
        RECT 69.710 193.625 70.005 194.445 ;
        RECT 70.175 194.175 70.405 195.875 ;
        RECT 70.620 195.370 70.875 196.175 ;
        RECT 71.075 195.560 71.405 196.005 ;
        RECT 71.575 195.730 71.850 196.175 ;
        RECT 72.085 195.560 72.415 196.005 ;
        RECT 71.075 195.380 72.415 195.560 ;
        RECT 72.875 195.200 73.205 195.865 ;
        RECT 73.475 195.430 73.745 196.175 ;
        RECT 74.375 196.170 80.650 196.175 ;
        RECT 73.915 195.260 74.205 196.000 ;
        RECT 74.375 195.445 74.630 196.170 ;
        RECT 74.815 195.275 75.075 196.000 ;
        RECT 75.245 195.445 75.490 196.170 ;
        RECT 75.675 195.275 75.935 196.000 ;
        RECT 76.105 195.445 76.350 196.170 ;
        RECT 76.535 195.275 76.795 196.000 ;
        RECT 76.965 195.445 77.210 196.170 ;
        RECT 77.380 195.275 77.640 196.000 ;
        RECT 77.810 195.445 78.070 196.170 ;
        RECT 78.240 195.275 78.500 196.000 ;
        RECT 78.670 195.445 78.930 196.170 ;
        RECT 79.100 195.275 79.360 196.000 ;
        RECT 79.530 195.445 79.790 196.170 ;
        RECT 79.960 195.275 80.220 196.000 ;
        RECT 80.390 195.375 80.650 196.170 ;
        RECT 74.815 195.260 80.220 195.275 ;
        RECT 70.620 195.030 73.205 195.200 ;
        RECT 73.475 195.035 80.220 195.260 ;
        RECT 70.620 194.415 70.930 195.030 ;
        RECT 71.100 194.585 71.430 194.815 ;
        RECT 71.600 194.585 72.070 194.815 ;
        RECT 72.240 194.645 72.695 194.815 ;
        RECT 72.240 194.585 72.690 194.645 ;
        RECT 72.880 194.585 73.215 194.815 ;
        RECT 73.475 194.445 74.640 195.035 ;
        RECT 80.820 194.865 81.070 196.000 ;
        RECT 81.250 195.365 81.510 196.175 ;
        RECT 81.685 194.865 81.930 196.005 ;
        RECT 82.110 195.365 82.405 196.175 ;
        RECT 82.585 195.010 82.875 196.175 ;
        RECT 83.065 195.585 83.305 195.975 ;
        RECT 83.475 195.765 83.825 196.175 ;
        RECT 83.065 195.385 83.815 195.585 ;
        RECT 74.810 194.615 81.930 194.865 ;
        RECT 70.620 194.235 73.205 194.415 ;
        RECT 73.475 194.275 80.220 194.445 ;
        RECT 70.175 193.795 70.395 194.175 ;
        RECT 70.565 193.625 71.415 193.985 ;
        RECT 71.895 193.815 72.225 194.235 ;
        RECT 72.430 193.625 72.705 194.065 ;
        RECT 72.875 193.815 73.205 194.235 ;
        RECT 73.475 193.625 73.775 194.105 ;
        RECT 73.945 193.820 74.205 194.275 ;
        RECT 74.375 193.625 74.635 194.105 ;
        RECT 74.815 193.820 75.075 194.275 ;
        RECT 75.245 193.625 75.495 194.105 ;
        RECT 75.675 193.820 75.935 194.275 ;
        RECT 76.105 193.625 76.355 194.105 ;
        RECT 76.535 193.820 76.795 194.275 ;
        RECT 76.965 193.625 77.210 194.105 ;
        RECT 77.380 193.820 77.655 194.275 ;
        RECT 77.825 193.625 78.070 194.105 ;
        RECT 78.240 193.820 78.500 194.275 ;
        RECT 78.670 193.625 78.930 194.105 ;
        RECT 79.100 193.820 79.360 194.275 ;
        RECT 79.530 193.625 79.790 194.105 ;
        RECT 79.960 193.820 80.220 194.275 ;
        RECT 80.390 193.625 80.650 194.185 ;
        RECT 80.820 193.805 81.070 194.615 ;
        RECT 81.250 193.625 81.510 194.150 ;
        RECT 81.680 193.805 81.930 194.615 ;
        RECT 82.100 194.305 82.415 194.865 ;
        RECT 82.110 193.625 82.415 194.135 ;
        RECT 82.585 193.625 82.875 194.350 ;
        RECT 83.065 193.865 83.295 195.205 ;
        RECT 83.475 194.705 83.815 195.385 ;
        RECT 83.995 194.885 84.325 195.995 ;
        RECT 84.495 195.525 84.675 195.995 ;
        RECT 84.845 195.695 85.175 196.175 ;
        RECT 85.350 195.525 85.520 195.995 ;
        RECT 84.495 195.325 85.520 195.525 ;
        RECT 83.475 193.805 83.705 194.705 ;
        RECT 83.995 194.585 84.540 194.885 ;
        RECT 83.905 193.625 84.150 194.405 ;
        RECT 84.320 194.355 84.540 194.585 ;
        RECT 84.710 194.535 85.135 195.155 ;
        RECT 85.330 194.535 85.590 195.155 ;
        RECT 85.785 195.035 86.070 196.175 ;
        RECT 85.800 194.355 86.060 194.865 ;
        RECT 84.320 194.165 86.060 194.355 ;
        RECT 84.320 193.805 84.750 194.165 ;
        RECT 85.330 193.625 86.060 193.995 ;
        RECT 86.260 193.805 86.540 195.995 ;
        RECT 86.765 195.035 86.995 196.175 ;
        RECT 87.165 195.025 87.495 196.005 ;
        RECT 87.665 195.035 87.875 196.175 ;
        RECT 88.105 195.085 89.315 196.175 ;
        RECT 86.745 194.615 87.075 194.865 ;
        RECT 86.765 193.625 86.995 194.445 ;
        RECT 87.245 194.425 87.495 195.025 ;
        RECT 88.105 194.545 88.625 195.085 ;
        RECT 87.165 193.795 87.495 194.425 ;
        RECT 87.665 193.625 87.875 194.445 ;
        RECT 88.795 194.375 89.315 194.915 ;
        RECT 88.105 193.625 89.315 194.375 ;
        RECT 18.100 193.455 89.400 193.625 ;
        RECT 18.185 192.705 19.395 193.455 ;
        RECT 18.185 192.165 18.705 192.705 ;
        RECT 19.570 192.615 19.830 193.455 ;
        RECT 20.005 192.710 20.260 193.285 ;
        RECT 20.430 193.075 20.760 193.455 ;
        RECT 20.975 192.905 21.145 193.285 ;
        RECT 20.430 192.735 21.145 192.905 ;
        RECT 21.495 192.905 21.665 193.285 ;
        RECT 21.845 193.075 22.175 193.455 ;
        RECT 21.495 192.735 22.160 192.905 ;
        RECT 22.355 192.780 22.615 193.285 ;
        RECT 18.875 191.995 19.395 192.535 ;
        RECT 18.185 190.905 19.395 191.995 ;
        RECT 19.570 190.905 19.830 192.055 ;
        RECT 20.005 191.980 20.175 192.710 ;
        RECT 20.430 192.545 20.600 192.735 ;
        RECT 20.345 192.215 20.600 192.545 ;
        RECT 20.430 192.005 20.600 192.215 ;
        RECT 20.880 192.185 21.235 192.555 ;
        RECT 21.425 192.185 21.765 192.555 ;
        RECT 21.990 192.480 22.160 192.735 ;
        RECT 21.990 192.150 22.265 192.480 ;
        RECT 21.990 192.005 22.160 192.150 ;
        RECT 20.005 191.075 20.260 191.980 ;
        RECT 20.430 191.835 21.145 192.005 ;
        RECT 20.430 190.905 20.760 191.665 ;
        RECT 20.975 191.075 21.145 191.835 ;
        RECT 21.485 191.835 22.160 192.005 ;
        RECT 22.435 191.980 22.615 192.780 ;
        RECT 21.485 191.075 21.665 191.835 ;
        RECT 21.845 190.905 22.175 191.665 ;
        RECT 22.345 191.075 22.615 191.980 ;
        RECT 22.785 192.780 23.045 193.285 ;
        RECT 23.225 193.075 23.555 193.455 ;
        RECT 23.735 192.905 23.905 193.285 ;
        RECT 22.785 191.980 22.955 192.780 ;
        RECT 23.240 192.735 23.905 192.905 ;
        RECT 23.240 192.480 23.410 192.735 ;
        RECT 24.225 192.635 24.435 193.455 ;
        RECT 24.605 192.655 24.935 193.285 ;
        RECT 23.125 192.150 23.410 192.480 ;
        RECT 23.645 192.185 23.975 192.555 ;
        RECT 23.240 192.005 23.410 192.150 ;
        RECT 24.605 192.055 24.855 192.655 ;
        RECT 25.105 192.635 25.335 193.455 ;
        RECT 25.025 192.215 25.355 192.465 ;
        RECT 22.785 191.075 23.055 191.980 ;
        RECT 23.240 191.835 23.905 192.005 ;
        RECT 23.225 190.905 23.555 191.665 ;
        RECT 23.735 191.075 23.905 191.835 ;
        RECT 24.225 190.905 24.435 192.045 ;
        RECT 24.605 191.075 24.935 192.055 ;
        RECT 25.105 190.905 25.335 192.045 ;
        RECT 26.015 191.085 26.275 193.275 ;
        RECT 26.535 193.085 27.205 193.455 ;
        RECT 27.385 192.905 27.695 193.275 ;
        RECT 26.465 192.705 27.695 192.905 ;
        RECT 26.465 192.035 26.755 192.705 ;
        RECT 27.875 192.525 28.105 193.165 ;
        RECT 28.285 192.725 28.575 193.455 ;
        RECT 28.800 192.715 29.415 193.285 ;
        RECT 29.585 192.945 29.800 193.455 ;
        RECT 30.030 192.945 30.310 193.275 ;
        RECT 30.490 192.945 30.730 193.455 ;
        RECT 26.935 192.215 27.400 192.525 ;
        RECT 27.580 192.215 28.105 192.525 ;
        RECT 28.285 192.215 28.585 192.545 ;
        RECT 26.465 191.815 27.235 192.035 ;
        RECT 26.445 190.905 26.785 191.635 ;
        RECT 26.965 191.085 27.235 191.815 ;
        RECT 27.415 191.795 28.575 192.035 ;
        RECT 27.415 191.085 27.645 191.795 ;
        RECT 27.815 190.905 28.145 191.615 ;
        RECT 28.315 191.085 28.575 191.795 ;
        RECT 28.800 191.695 29.115 192.715 ;
        RECT 29.285 192.045 29.455 192.545 ;
        RECT 29.705 192.215 29.970 192.775 ;
        RECT 30.140 192.045 30.310 192.945 ;
        RECT 31.615 192.905 31.785 193.285 ;
        RECT 31.965 193.075 32.295 193.455 ;
        RECT 30.480 192.215 30.835 192.775 ;
        RECT 31.615 192.735 32.280 192.905 ;
        RECT 32.475 192.780 32.735 193.285 ;
        RECT 31.545 192.185 31.885 192.555 ;
        RECT 32.110 192.480 32.280 192.735 ;
        RECT 32.110 192.150 32.385 192.480 ;
        RECT 29.285 191.875 30.710 192.045 ;
        RECT 32.110 192.005 32.280 192.150 ;
        RECT 28.800 191.075 29.335 191.695 ;
        RECT 29.505 190.905 29.835 191.705 ;
        RECT 30.320 191.700 30.710 191.875 ;
        RECT 31.605 191.835 32.280 192.005 ;
        RECT 32.555 191.980 32.735 192.780 ;
        RECT 32.915 192.725 33.215 193.455 ;
        RECT 33.395 192.545 33.625 193.165 ;
        RECT 33.825 192.895 34.050 193.275 ;
        RECT 34.220 193.065 34.550 193.455 ;
        RECT 35.665 192.995 36.225 193.285 ;
        RECT 36.395 192.995 36.645 193.455 ;
        RECT 33.825 192.715 34.155 192.895 ;
        RECT 32.920 192.215 33.215 192.545 ;
        RECT 33.395 192.215 33.810 192.545 ;
        RECT 33.980 192.045 34.155 192.715 ;
        RECT 34.325 192.215 34.565 192.865 ;
        RECT 31.605 191.075 31.785 191.835 ;
        RECT 31.965 190.905 32.295 191.665 ;
        RECT 32.465 191.075 32.735 191.980 ;
        RECT 32.915 191.685 33.810 192.015 ;
        RECT 33.980 191.855 34.565 192.045 ;
        RECT 32.915 191.515 34.120 191.685 ;
        RECT 32.915 191.085 33.245 191.515 ;
        RECT 33.425 190.905 33.620 191.345 ;
        RECT 33.790 191.085 34.120 191.515 ;
        RECT 34.290 191.085 34.565 191.855 ;
        RECT 35.665 191.625 35.915 192.995 ;
        RECT 37.265 192.825 37.595 193.185 ;
        RECT 37.970 192.950 38.305 193.455 ;
        RECT 38.475 192.885 38.715 193.260 ;
        RECT 38.995 193.125 39.165 193.270 ;
        RECT 38.995 192.930 39.370 193.125 ;
        RECT 39.730 192.960 40.125 193.455 ;
        RECT 36.205 192.635 37.595 192.825 ;
        RECT 36.205 192.545 36.375 192.635 ;
        RECT 36.085 192.215 36.375 192.545 ;
        RECT 36.545 192.215 36.885 192.465 ;
        RECT 37.105 192.215 37.780 192.465 ;
        RECT 36.205 191.965 36.375 192.215 ;
        RECT 36.205 191.795 37.145 191.965 ;
        RECT 37.515 191.855 37.780 192.215 ;
        RECT 38.025 191.925 38.325 192.775 ;
        RECT 38.495 192.735 38.715 192.885 ;
        RECT 38.495 192.405 39.030 192.735 ;
        RECT 39.200 192.595 39.370 192.930 ;
        RECT 40.295 192.765 40.535 193.285 ;
        RECT 41.185 193.075 41.515 193.455 ;
        RECT 35.665 191.075 36.125 191.625 ;
        RECT 36.315 190.905 36.645 191.625 ;
        RECT 36.845 191.245 37.145 191.795 ;
        RECT 38.495 191.755 38.730 192.405 ;
        RECT 39.200 192.235 40.185 192.595 ;
        RECT 37.315 190.905 37.595 191.575 ;
        RECT 38.055 191.525 38.730 191.755 ;
        RECT 38.900 192.215 40.185 192.235 ;
        RECT 38.900 192.065 39.760 192.215 ;
        RECT 38.055 191.095 38.225 191.525 ;
        RECT 38.395 190.905 38.725 191.355 ;
        RECT 38.900 191.120 39.185 192.065 ;
        RECT 40.360 191.960 40.535 192.765 ;
        RECT 40.740 192.905 41.015 193.045 ;
        RECT 41.685 192.905 41.895 193.075 ;
        RECT 40.740 192.715 41.895 192.905 ;
        RECT 42.065 192.905 42.395 193.285 ;
        RECT 42.585 193.075 42.915 193.455 ;
        RECT 42.065 192.700 42.915 192.905 ;
        RECT 40.735 192.090 40.995 192.545 ;
        RECT 41.250 192.140 41.835 192.515 ;
        RECT 39.360 191.585 40.055 191.895 ;
        RECT 39.365 190.905 40.050 191.375 ;
        RECT 40.230 191.175 40.535 191.960 ;
        RECT 40.740 190.905 41.065 191.890 ;
        RECT 41.250 191.755 41.455 192.140 ;
        RECT 42.005 191.925 42.415 192.530 ;
        RECT 42.585 192.210 42.915 192.700 ;
        RECT 42.585 191.755 42.755 192.210 ;
        RECT 41.245 191.585 41.455 191.755 ;
        RECT 41.250 191.555 41.455 191.585 ;
        RECT 41.635 191.535 42.755 191.755 ;
        RECT 41.635 191.075 41.895 191.535 ;
        RECT 42.065 190.905 42.915 191.355 ;
        RECT 43.085 191.075 43.330 193.285 ;
        RECT 43.515 192.655 43.755 193.455 ;
        RECT 43.945 192.730 44.235 193.455 ;
        RECT 44.405 192.955 44.665 193.285 ;
        RECT 44.835 193.095 45.165 193.455 ;
        RECT 45.420 193.075 46.720 193.285 ;
        RECT 43.515 190.905 43.770 191.905 ;
        RECT 43.945 190.905 44.235 192.070 ;
        RECT 44.405 191.755 44.575 192.955 ;
        RECT 45.420 192.925 45.590 193.075 ;
        RECT 44.835 192.800 45.590 192.925 ;
        RECT 44.745 192.755 45.590 192.800 ;
        RECT 44.745 192.635 45.015 192.755 ;
        RECT 44.745 192.060 44.915 192.635 ;
        RECT 45.145 192.195 45.555 192.500 ;
        RECT 45.845 192.465 46.055 192.865 ;
        RECT 45.725 192.255 46.055 192.465 ;
        RECT 46.300 192.465 46.520 192.865 ;
        RECT 46.995 192.690 47.450 193.455 ;
        RECT 46.300 192.255 46.775 192.465 ;
        RECT 46.965 192.265 47.455 192.465 ;
        RECT 44.745 192.025 44.945 192.060 ;
        RECT 46.275 192.025 47.450 192.085 ;
        RECT 44.745 191.915 47.450 192.025 ;
        RECT 44.805 191.855 46.605 191.915 ;
        RECT 46.275 191.825 46.605 191.855 ;
        RECT 44.405 191.075 44.665 191.755 ;
        RECT 44.835 190.905 45.085 191.685 ;
        RECT 45.335 191.655 46.170 191.665 ;
        RECT 46.760 191.655 46.945 191.745 ;
        RECT 45.335 191.455 46.945 191.655 ;
        RECT 45.335 191.075 45.585 191.455 ;
        RECT 46.715 191.415 46.945 191.455 ;
        RECT 47.195 191.295 47.450 191.915 ;
        RECT 45.755 190.905 46.110 191.285 ;
        RECT 47.115 191.075 47.450 191.295 ;
        RECT 47.625 191.075 47.905 193.175 ;
        RECT 48.135 192.995 48.305 193.455 ;
        RECT 48.575 193.065 49.825 193.245 ;
        RECT 48.960 192.825 49.325 192.895 ;
        RECT 48.075 192.645 49.325 192.825 ;
        RECT 49.495 192.845 49.825 193.065 ;
        RECT 49.995 193.015 50.165 193.455 ;
        RECT 50.335 192.845 50.675 193.260 ;
        RECT 50.935 192.975 51.235 193.455 ;
        RECT 49.495 192.675 50.675 192.845 ;
        RECT 51.405 192.805 51.665 193.260 ;
        RECT 51.835 192.975 52.095 193.455 ;
        RECT 52.275 192.805 52.535 193.260 ;
        RECT 52.705 192.975 52.955 193.455 ;
        RECT 53.135 192.805 53.395 193.260 ;
        RECT 53.565 192.975 53.815 193.455 ;
        RECT 53.995 192.805 54.255 193.260 ;
        RECT 54.425 192.975 54.670 193.455 ;
        RECT 54.840 192.805 55.115 193.260 ;
        RECT 55.285 192.975 55.530 193.455 ;
        RECT 55.700 192.805 55.960 193.260 ;
        RECT 56.130 192.975 56.390 193.455 ;
        RECT 56.560 192.805 56.820 193.260 ;
        RECT 56.990 192.975 57.250 193.455 ;
        RECT 57.420 192.805 57.680 193.260 ;
        RECT 57.850 192.895 58.110 193.455 ;
        RECT 48.075 192.045 48.350 192.645 ;
        RECT 50.935 192.635 57.680 192.805 ;
        RECT 48.520 192.215 48.875 192.465 ;
        RECT 49.070 192.435 49.535 192.465 ;
        RECT 49.065 192.265 49.535 192.435 ;
        RECT 49.070 192.215 49.535 192.265 ;
        RECT 49.705 192.215 50.035 192.465 ;
        RECT 50.210 192.265 50.675 192.465 ;
        RECT 49.855 192.095 50.035 192.215 ;
        RECT 48.075 191.835 49.685 192.045 ;
        RECT 49.855 191.925 50.185 192.095 ;
        RECT 49.275 191.735 49.685 191.835 ;
        RECT 48.095 190.905 48.880 191.665 ;
        RECT 49.275 191.075 49.660 191.735 ;
        RECT 49.985 191.135 50.185 191.925 ;
        RECT 50.355 190.905 50.675 192.085 ;
        RECT 50.935 192.045 52.100 192.635 ;
        RECT 58.280 192.465 58.530 193.275 ;
        RECT 58.710 192.930 58.970 193.455 ;
        RECT 59.140 192.465 59.390 193.275 ;
        RECT 59.570 192.945 59.875 193.455 ;
        RECT 60.595 192.975 60.895 193.455 ;
        RECT 61.065 192.805 61.325 193.260 ;
        RECT 61.495 192.975 61.755 193.455 ;
        RECT 61.935 192.805 62.195 193.260 ;
        RECT 62.365 192.975 62.615 193.455 ;
        RECT 62.795 192.805 63.055 193.260 ;
        RECT 63.225 192.975 63.475 193.455 ;
        RECT 63.655 192.805 63.915 193.260 ;
        RECT 64.085 192.975 64.330 193.455 ;
        RECT 64.500 192.805 64.775 193.260 ;
        RECT 64.945 192.975 65.190 193.455 ;
        RECT 65.360 192.805 65.620 193.260 ;
        RECT 65.790 192.975 66.050 193.455 ;
        RECT 66.220 192.805 66.480 193.260 ;
        RECT 66.650 192.975 66.910 193.455 ;
        RECT 67.080 192.805 67.340 193.260 ;
        RECT 67.510 192.895 67.770 193.455 ;
        RECT 52.270 192.215 59.390 192.465 ;
        RECT 59.560 192.215 59.875 192.775 ;
        RECT 60.595 192.635 67.340 192.805 ;
        RECT 50.935 191.820 57.680 192.045 ;
        RECT 50.935 190.905 51.205 191.650 ;
        RECT 51.375 191.080 51.665 191.820 ;
        RECT 52.275 191.805 57.680 191.820 ;
        RECT 51.835 190.910 52.090 191.635 ;
        RECT 52.275 191.080 52.535 191.805 ;
        RECT 52.705 190.910 52.950 191.635 ;
        RECT 53.135 191.080 53.395 191.805 ;
        RECT 53.565 190.910 53.810 191.635 ;
        RECT 53.995 191.080 54.255 191.805 ;
        RECT 54.425 190.910 54.670 191.635 ;
        RECT 54.840 191.080 55.100 191.805 ;
        RECT 55.270 190.910 55.530 191.635 ;
        RECT 55.700 191.080 55.960 191.805 ;
        RECT 56.130 190.910 56.390 191.635 ;
        RECT 56.560 191.080 56.820 191.805 ;
        RECT 56.990 190.910 57.250 191.635 ;
        RECT 57.420 191.080 57.680 191.805 ;
        RECT 57.850 190.910 58.110 191.705 ;
        RECT 58.280 191.080 58.530 192.215 ;
        RECT 51.835 190.905 58.110 190.910 ;
        RECT 58.710 190.905 58.970 191.715 ;
        RECT 59.145 191.075 59.390 192.215 ;
        RECT 60.595 192.045 61.760 192.635 ;
        RECT 67.940 192.465 68.190 193.275 ;
        RECT 68.370 192.930 68.630 193.455 ;
        RECT 68.800 192.465 69.050 193.275 ;
        RECT 69.230 192.945 69.535 193.455 ;
        RECT 61.930 192.215 69.050 192.465 ;
        RECT 69.220 192.215 69.535 192.775 ;
        RECT 69.705 192.730 69.995 193.455 ;
        RECT 70.165 192.805 70.425 193.250 ;
        RECT 70.675 192.975 70.845 193.455 ;
        RECT 71.015 192.945 71.365 193.275 ;
        RECT 71.600 192.975 71.770 193.455 ;
        RECT 70.165 192.635 70.845 192.805 ;
        RECT 60.595 191.820 67.340 192.045 ;
        RECT 59.570 190.905 59.865 191.715 ;
        RECT 60.595 190.905 60.865 191.650 ;
        RECT 61.035 191.080 61.325 191.820 ;
        RECT 61.935 191.805 67.340 191.820 ;
        RECT 61.495 190.910 61.750 191.635 ;
        RECT 61.935 191.080 62.195 191.805 ;
        RECT 62.365 190.910 62.610 191.635 ;
        RECT 62.795 191.080 63.055 191.805 ;
        RECT 63.225 190.910 63.470 191.635 ;
        RECT 63.655 191.080 63.915 191.805 ;
        RECT 64.085 190.910 64.330 191.635 ;
        RECT 64.500 191.080 64.760 191.805 ;
        RECT 64.930 190.910 65.190 191.635 ;
        RECT 65.360 191.080 65.620 191.805 ;
        RECT 65.790 190.910 66.050 191.635 ;
        RECT 66.220 191.080 66.480 191.805 ;
        RECT 66.650 190.910 66.910 191.635 ;
        RECT 67.080 191.080 67.340 191.805 ;
        RECT 67.510 190.910 67.770 191.705 ;
        RECT 67.940 191.080 68.190 192.215 ;
        RECT 61.495 190.905 67.770 190.910 ;
        RECT 68.370 190.905 68.630 191.715 ;
        RECT 68.805 191.075 69.050 192.215 ;
        RECT 69.230 190.905 69.525 191.715 ;
        RECT 69.705 190.905 69.995 192.070 ;
        RECT 70.165 191.900 70.505 192.465 ;
        RECT 70.675 191.730 70.845 192.635 ;
        RECT 71.015 192.045 71.185 192.945 ;
        RECT 72.070 192.885 72.240 193.235 ;
        RECT 72.410 193.055 72.740 193.455 ;
        RECT 72.910 192.935 73.165 193.235 ;
        RECT 72.910 192.885 73.215 192.935 ;
        RECT 72.070 192.805 73.215 192.885 ;
        RECT 71.505 192.775 73.215 192.805 ;
        RECT 71.355 192.715 73.215 192.775 ;
        RECT 71.355 192.635 72.240 192.715 ;
        RECT 71.355 192.605 71.675 192.635 ;
        RECT 71.355 192.215 71.525 192.605 ;
        RECT 71.015 191.840 71.410 192.045 ;
        RECT 71.775 191.925 72.310 192.465 ;
        RECT 72.570 192.215 72.870 192.545 ;
        RECT 72.570 191.755 72.740 192.215 ;
        RECT 73.045 192.045 73.215 192.715 ;
        RECT 73.845 192.655 74.105 193.455 ;
        RECT 70.165 191.670 70.845 191.730 ;
        RECT 71.630 191.670 72.740 191.755 ;
        RECT 70.165 191.585 72.740 191.670 ;
        RECT 72.910 191.615 73.215 192.045 ;
        RECT 70.165 191.500 71.800 191.585 ;
        RECT 70.165 191.320 70.425 191.500 ;
        RECT 70.630 190.905 70.990 191.330 ;
        RECT 71.505 190.905 71.835 191.330 ;
        RECT 72.015 191.175 73.215 191.415 ;
        RECT 73.845 190.905 74.105 192.045 ;
        RECT 74.275 191.075 74.605 193.285 ;
        RECT 74.855 192.715 75.185 193.455 ;
        RECT 75.455 192.885 75.785 193.285 ;
        RECT 75.955 193.055 76.285 193.455 ;
        RECT 76.455 193.115 77.815 193.285 ;
        RECT 76.455 192.885 76.785 193.115 ;
        RECT 75.455 192.715 76.785 192.885 ;
        RECT 76.955 192.715 77.285 192.945 ;
        RECT 74.775 191.755 75.085 192.545 ;
        RECT 75.255 191.925 75.475 192.545 ;
        RECT 75.745 191.925 75.920 192.545 ;
        RECT 76.175 191.925 76.395 192.545 ;
        RECT 76.670 192.435 76.915 192.545 ;
        RECT 76.665 192.265 76.915 192.435 ;
        RECT 76.670 191.925 76.915 192.265 ;
        RECT 77.085 191.755 77.285 192.715 ;
        RECT 77.455 192.635 77.815 193.115 ;
        RECT 78.995 192.975 79.295 193.455 ;
        RECT 79.465 192.805 79.725 193.260 ;
        RECT 79.895 192.975 80.155 193.455 ;
        RECT 80.335 192.805 80.595 193.260 ;
        RECT 80.765 192.975 81.015 193.455 ;
        RECT 81.195 192.805 81.455 193.260 ;
        RECT 81.625 192.975 81.875 193.455 ;
        RECT 82.055 192.805 82.315 193.260 ;
        RECT 82.485 192.975 82.730 193.455 ;
        RECT 82.900 192.805 83.175 193.260 ;
        RECT 83.345 192.975 83.590 193.455 ;
        RECT 83.760 192.805 84.020 193.260 ;
        RECT 84.190 192.975 84.450 193.455 ;
        RECT 84.620 192.805 84.880 193.260 ;
        RECT 85.050 192.975 85.310 193.455 ;
        RECT 85.480 192.805 85.740 193.260 ;
        RECT 85.910 192.895 86.170 193.455 ;
        RECT 78.995 192.635 85.740 192.805 ;
        RECT 77.455 192.295 77.815 192.465 ;
        RECT 77.485 192.215 77.815 192.295 ;
        RECT 78.995 192.045 80.160 192.635 ;
        RECT 86.340 192.465 86.590 193.275 ;
        RECT 86.770 192.930 87.030 193.455 ;
        RECT 87.200 192.465 87.450 193.275 ;
        RECT 87.630 192.945 87.935 193.455 ;
        RECT 80.330 192.215 87.450 192.465 ;
        RECT 87.620 192.215 87.935 192.775 ;
        RECT 88.105 192.705 89.315 193.455 ;
        RECT 74.775 191.585 77.285 191.755 ;
        RECT 74.775 190.905 75.285 191.415 ;
        RECT 76.455 191.075 76.785 191.585 ;
        RECT 77.455 190.905 77.815 192.045 ;
        RECT 78.995 191.820 85.740 192.045 ;
        RECT 78.995 190.905 79.265 191.650 ;
        RECT 79.435 191.080 79.725 191.820 ;
        RECT 80.335 191.805 85.740 191.820 ;
        RECT 79.895 190.910 80.150 191.635 ;
        RECT 80.335 191.080 80.595 191.805 ;
        RECT 80.765 190.910 81.010 191.635 ;
        RECT 81.195 191.080 81.455 191.805 ;
        RECT 81.625 190.910 81.870 191.635 ;
        RECT 82.055 191.080 82.315 191.805 ;
        RECT 82.485 190.910 82.730 191.635 ;
        RECT 82.900 191.080 83.160 191.805 ;
        RECT 83.330 190.910 83.590 191.635 ;
        RECT 83.760 191.080 84.020 191.805 ;
        RECT 84.190 190.910 84.450 191.635 ;
        RECT 84.620 191.080 84.880 191.805 ;
        RECT 85.050 190.910 85.310 191.635 ;
        RECT 85.480 191.080 85.740 191.805 ;
        RECT 85.910 190.910 86.170 191.705 ;
        RECT 86.340 191.080 86.590 192.215 ;
        RECT 79.895 190.905 86.170 190.910 ;
        RECT 86.770 190.905 87.030 191.715 ;
        RECT 87.205 191.075 87.450 192.215 ;
        RECT 88.105 191.995 88.625 192.535 ;
        RECT 88.795 192.165 89.315 192.705 ;
        RECT 87.630 190.905 87.925 191.715 ;
        RECT 88.105 190.905 89.315 191.995 ;
        RECT 18.100 190.735 89.400 190.905 ;
        RECT 18.185 189.645 19.395 190.735 ;
        RECT 18.185 188.935 18.705 189.475 ;
        RECT 18.875 189.105 19.395 189.645 ;
        RECT 20.485 189.660 20.755 190.565 ;
        RECT 20.925 189.975 21.255 190.735 ;
        RECT 21.435 189.805 21.605 190.565 ;
        RECT 18.185 188.185 19.395 188.935 ;
        RECT 20.485 188.860 20.655 189.660 ;
        RECT 20.940 189.635 21.605 189.805 ;
        RECT 21.865 189.660 22.135 190.565 ;
        RECT 22.305 189.975 22.635 190.735 ;
        RECT 22.815 189.805 22.985 190.565 ;
        RECT 20.940 189.490 21.110 189.635 ;
        RECT 20.825 189.160 21.110 189.490 ;
        RECT 20.940 188.905 21.110 189.160 ;
        RECT 21.345 189.085 21.675 189.455 ;
        RECT 20.485 188.355 20.745 188.860 ;
        RECT 20.940 188.735 21.605 188.905 ;
        RECT 20.925 188.185 21.255 188.565 ;
        RECT 21.435 188.355 21.605 188.735 ;
        RECT 21.865 188.860 22.035 189.660 ;
        RECT 22.320 189.635 22.985 189.805 ;
        RECT 23.245 189.660 23.515 190.565 ;
        RECT 23.685 189.975 24.015 190.735 ;
        RECT 24.195 189.805 24.365 190.565 ;
        RECT 24.815 190.010 25.145 190.735 ;
        RECT 22.320 189.490 22.490 189.635 ;
        RECT 22.205 189.160 22.490 189.490 ;
        RECT 22.320 188.905 22.490 189.160 ;
        RECT 22.725 189.085 23.055 189.455 ;
        RECT 21.865 188.355 22.125 188.860 ;
        RECT 22.320 188.735 22.985 188.905 ;
        RECT 22.305 188.185 22.635 188.565 ;
        RECT 22.815 188.355 22.985 188.735 ;
        RECT 23.245 188.860 23.415 189.660 ;
        RECT 23.700 189.635 24.365 189.805 ;
        RECT 23.700 189.490 23.870 189.635 ;
        RECT 23.585 189.160 23.870 189.490 ;
        RECT 23.700 188.905 23.870 189.160 ;
        RECT 24.105 189.085 24.435 189.455 ;
        RECT 23.245 188.355 23.505 188.860 ;
        RECT 23.700 188.735 24.365 188.905 ;
        RECT 23.685 188.185 24.015 188.565 ;
        RECT 24.195 188.355 24.365 188.735 ;
        RECT 24.625 188.355 25.145 189.840 ;
        RECT 25.315 189.015 25.835 190.565 ;
        RECT 26.190 189.765 26.580 189.940 ;
        RECT 27.065 189.935 27.395 190.735 ;
        RECT 27.565 189.945 28.100 190.565 ;
        RECT 26.190 189.595 27.615 189.765 ;
        RECT 26.065 188.865 26.420 189.425 ;
        RECT 25.315 188.185 25.655 188.845 ;
        RECT 26.590 188.695 26.760 189.595 ;
        RECT 26.930 188.865 27.195 189.425 ;
        RECT 27.445 189.095 27.615 189.595 ;
        RECT 27.785 188.925 28.100 189.945 ;
        RECT 28.310 189.585 28.570 190.735 ;
        RECT 28.745 189.660 29.000 190.565 ;
        RECT 29.170 189.975 29.500 190.735 ;
        RECT 29.715 189.805 29.885 190.565 ;
        RECT 26.170 188.185 26.410 188.695 ;
        RECT 26.590 188.365 26.870 188.695 ;
        RECT 27.100 188.185 27.315 188.695 ;
        RECT 27.485 188.355 28.100 188.925 ;
        RECT 28.310 188.185 28.570 189.025 ;
        RECT 28.745 188.930 28.915 189.660 ;
        RECT 29.170 189.635 29.885 189.805 ;
        RECT 29.170 189.425 29.340 189.635 ;
        RECT 31.065 189.570 31.355 190.735 ;
        RECT 32.450 189.595 32.785 190.565 ;
        RECT 32.955 189.595 33.125 190.735 ;
        RECT 33.295 190.395 35.325 190.565 ;
        RECT 29.085 189.095 29.340 189.425 ;
        RECT 28.745 188.355 29.000 188.930 ;
        RECT 29.170 188.905 29.340 189.095 ;
        RECT 29.620 189.085 29.975 189.455 ;
        RECT 32.450 188.925 32.620 189.595 ;
        RECT 33.295 189.425 33.465 190.395 ;
        RECT 32.790 189.095 33.045 189.425 ;
        RECT 33.270 189.095 33.465 189.425 ;
        RECT 33.635 190.055 34.760 190.225 ;
        RECT 32.875 188.925 33.045 189.095 ;
        RECT 33.635 188.925 33.805 190.055 ;
        RECT 29.170 188.735 29.885 188.905 ;
        RECT 29.170 188.185 29.500 188.565 ;
        RECT 29.715 188.355 29.885 188.735 ;
        RECT 31.065 188.185 31.355 188.910 ;
        RECT 32.450 188.355 32.705 188.925 ;
        RECT 32.875 188.755 33.805 188.925 ;
        RECT 33.975 189.715 34.985 189.885 ;
        RECT 33.975 188.915 34.145 189.715 ;
        RECT 33.630 188.720 33.805 188.755 ;
        RECT 32.875 188.185 33.205 188.585 ;
        RECT 33.630 188.355 34.160 188.720 ;
        RECT 34.350 188.695 34.625 189.515 ;
        RECT 34.345 188.525 34.625 188.695 ;
        RECT 34.350 188.355 34.625 188.525 ;
        RECT 34.795 188.355 34.985 189.715 ;
        RECT 35.155 189.730 35.325 190.395 ;
        RECT 35.495 189.975 35.665 190.735 ;
        RECT 35.900 189.975 36.415 190.385 ;
        RECT 35.155 189.540 35.905 189.730 ;
        RECT 36.075 189.165 36.415 189.975 ;
        RECT 37.135 189.805 37.305 190.565 ;
        RECT 37.485 189.975 37.815 190.735 ;
        RECT 37.135 189.635 37.800 189.805 ;
        RECT 37.985 189.660 38.255 190.565 ;
        RECT 37.630 189.490 37.800 189.635 ;
        RECT 35.185 188.995 36.415 189.165 ;
        RECT 37.065 189.085 37.395 189.455 ;
        RECT 37.630 189.160 37.915 189.490 ;
        RECT 35.165 188.185 35.675 188.720 ;
        RECT 35.895 188.390 36.140 188.995 ;
        RECT 37.630 188.905 37.800 189.160 ;
        RECT 37.135 188.735 37.800 188.905 ;
        RECT 38.085 188.860 38.255 189.660 ;
        RECT 38.435 190.125 38.765 190.555 ;
        RECT 38.945 190.295 39.140 190.735 ;
        RECT 39.310 190.125 39.640 190.555 ;
        RECT 38.435 189.955 39.640 190.125 ;
        RECT 38.435 189.625 39.330 189.955 ;
        RECT 39.810 189.785 40.085 190.555 ;
        RECT 40.355 189.990 40.625 190.735 ;
        RECT 41.255 190.730 47.530 190.735 ;
        RECT 40.795 189.820 41.085 190.560 ;
        RECT 41.255 190.005 41.510 190.730 ;
        RECT 41.695 189.835 41.955 190.560 ;
        RECT 42.125 190.005 42.370 190.730 ;
        RECT 42.555 189.835 42.815 190.560 ;
        RECT 42.985 190.005 43.230 190.730 ;
        RECT 43.415 189.835 43.675 190.560 ;
        RECT 43.845 190.005 44.090 190.730 ;
        RECT 44.260 189.835 44.520 190.560 ;
        RECT 44.690 190.005 44.950 190.730 ;
        RECT 45.120 189.835 45.380 190.560 ;
        RECT 45.550 190.005 45.810 190.730 ;
        RECT 45.980 189.835 46.240 190.560 ;
        RECT 46.410 190.005 46.670 190.730 ;
        RECT 46.840 189.835 47.100 190.560 ;
        RECT 47.270 189.935 47.530 190.730 ;
        RECT 41.695 189.820 47.100 189.835 ;
        RECT 39.500 189.595 40.085 189.785 ;
        RECT 40.355 189.595 47.100 189.820 ;
        RECT 38.440 189.095 38.735 189.425 ;
        RECT 38.915 189.095 39.330 189.425 ;
        RECT 37.135 188.355 37.305 188.735 ;
        RECT 37.485 188.185 37.815 188.565 ;
        RECT 37.995 188.355 38.255 188.860 ;
        RECT 38.435 188.185 38.735 188.915 ;
        RECT 38.915 188.475 39.145 189.095 ;
        RECT 39.500 188.925 39.675 189.595 ;
        RECT 39.345 188.745 39.675 188.925 ;
        RECT 39.845 188.775 40.085 189.425 ;
        RECT 40.355 189.005 41.520 189.595 ;
        RECT 47.700 189.425 47.950 190.560 ;
        RECT 48.130 189.925 48.390 190.735 ;
        RECT 48.565 189.425 48.810 190.565 ;
        RECT 48.990 189.925 49.285 190.735 ;
        RECT 49.470 189.865 49.735 190.565 ;
        RECT 49.905 190.035 50.235 190.735 ;
        RECT 50.405 189.865 51.075 190.565 ;
        RECT 51.580 190.035 52.010 190.735 ;
        RECT 52.190 190.175 52.380 190.565 ;
        RECT 52.550 190.355 52.880 190.735 ;
        RECT 53.235 190.395 54.395 190.565 ;
        RECT 52.190 190.005 52.920 190.175 ;
        RECT 49.470 189.610 52.045 189.865 ;
        RECT 41.690 189.175 48.810 189.425 ;
        RECT 40.355 188.835 47.100 189.005 ;
        RECT 39.345 188.365 39.570 188.745 ;
        RECT 39.740 188.185 40.070 188.575 ;
        RECT 40.355 188.185 40.655 188.665 ;
        RECT 40.825 188.380 41.085 188.835 ;
        RECT 41.255 188.185 41.515 188.665 ;
        RECT 41.695 188.380 41.955 188.835 ;
        RECT 42.125 188.185 42.375 188.665 ;
        RECT 42.555 188.380 42.815 188.835 ;
        RECT 42.985 188.185 43.235 188.665 ;
        RECT 43.415 188.380 43.675 188.835 ;
        RECT 43.845 188.185 44.090 188.665 ;
        RECT 44.260 188.380 44.535 188.835 ;
        RECT 44.705 188.185 44.950 188.665 ;
        RECT 45.120 188.380 45.380 188.835 ;
        RECT 45.550 188.185 45.810 188.665 ;
        RECT 45.980 188.380 46.240 188.835 ;
        RECT 46.410 188.185 46.670 188.665 ;
        RECT 46.840 188.380 47.100 188.835 ;
        RECT 47.270 188.185 47.530 188.745 ;
        RECT 47.700 188.365 47.950 189.175 ;
        RECT 48.130 188.185 48.390 188.710 ;
        RECT 48.560 188.365 48.810 189.175 ;
        RECT 48.980 188.865 49.295 189.425 ;
        RECT 49.465 189.095 49.740 189.425 ;
        RECT 49.910 188.925 50.090 189.610 ;
        RECT 51.875 189.425 52.045 189.610 ;
        RECT 50.260 189.095 50.620 189.425 ;
        RECT 50.910 189.375 51.200 189.425 ;
        RECT 50.905 189.205 51.200 189.375 ;
        RECT 50.910 189.095 51.200 189.205 ;
        RECT 51.370 189.095 51.705 189.425 ;
        RECT 51.875 189.095 52.555 189.425 ;
        RECT 48.990 188.185 49.295 188.695 ;
        RECT 49.475 188.525 50.090 188.925 ;
        RECT 50.260 188.735 51.530 188.925 ;
        RECT 52.725 188.885 52.920 190.005 ;
        RECT 53.235 189.895 53.405 190.395 ;
        RECT 53.665 189.765 53.835 190.225 ;
        RECT 54.065 190.145 54.395 190.395 ;
        RECT 54.620 190.315 54.950 190.735 ;
        RECT 55.205 190.145 55.490 190.565 ;
        RECT 54.065 189.975 55.490 190.145 ;
        RECT 55.735 189.935 56.065 190.735 ;
        RECT 56.315 190.015 56.650 190.525 ;
        RECT 53.210 189.425 53.415 189.715 ;
        RECT 53.665 189.595 56.035 189.765 ;
        RECT 55.865 189.425 56.035 189.595 ;
        RECT 53.210 189.375 53.560 189.425 ;
        RECT 53.205 189.205 53.560 189.375 ;
        RECT 53.210 189.095 53.560 189.205 ;
        RECT 52.100 188.715 52.920 188.885 ;
        RECT 49.475 188.355 49.810 188.525 ;
        RECT 50.770 188.185 51.105 188.565 ;
        RECT 51.695 188.185 51.930 188.625 ;
        RECT 52.100 188.355 52.430 188.715 ;
        RECT 52.600 188.185 52.930 188.545 ;
        RECT 53.155 188.185 53.485 188.905 ;
        RECT 53.870 188.760 54.290 189.425 ;
        RECT 54.460 189.035 54.750 189.425 ;
        RECT 54.940 189.375 55.210 189.425 ;
        RECT 55.420 189.375 55.670 189.425 ;
        RECT 54.940 189.205 55.215 189.375 ;
        RECT 55.420 189.205 55.675 189.375 ;
        RECT 54.460 188.865 54.755 189.035 ;
        RECT 54.460 188.765 54.750 188.865 ;
        RECT 54.940 188.765 55.210 189.205 ;
        RECT 55.420 189.095 55.670 189.205 ;
        RECT 55.865 189.095 56.170 189.425 ;
        RECT 55.865 188.925 56.035 189.095 ;
        RECT 55.475 188.755 56.035 188.925 ;
        RECT 55.475 188.585 55.645 188.755 ;
        RECT 56.395 188.660 56.650 190.015 ;
        RECT 56.825 189.570 57.115 190.735 ;
        RECT 57.340 189.865 57.625 190.735 ;
        RECT 57.795 190.105 58.055 190.565 ;
        RECT 58.230 190.275 58.485 190.735 ;
        RECT 58.655 190.105 58.915 190.565 ;
        RECT 57.795 189.935 58.915 190.105 ;
        RECT 59.085 189.935 59.395 190.735 ;
        RECT 57.795 189.685 58.055 189.935 ;
        RECT 59.565 189.765 59.875 190.565 ;
        RECT 60.045 190.315 60.385 190.735 ;
        RECT 60.555 190.145 60.805 190.565 ;
        RECT 57.300 189.515 58.055 189.685 ;
        RECT 58.845 189.595 59.875 189.765 ;
        RECT 57.300 189.005 57.705 189.515 ;
        RECT 58.845 189.345 59.015 189.595 ;
        RECT 57.875 189.175 59.015 189.345 ;
        RECT 54.030 188.415 55.645 188.585 ;
        RECT 55.815 188.185 56.145 188.585 ;
        RECT 56.315 188.400 56.650 188.660 ;
        RECT 56.825 188.185 57.115 188.910 ;
        RECT 57.300 188.835 58.950 189.005 ;
        RECT 59.185 188.855 59.535 189.425 ;
        RECT 57.345 188.185 57.625 188.665 ;
        RECT 57.795 188.445 58.055 188.835 ;
        RECT 58.230 188.185 58.485 188.665 ;
        RECT 58.655 188.445 58.950 188.835 ;
        RECT 59.705 188.685 59.875 189.595 ;
        RECT 60.045 189.975 60.805 190.145 ;
        RECT 60.045 189.005 60.355 189.975 ;
        RECT 60.975 189.895 61.305 190.735 ;
        RECT 61.795 190.145 62.550 190.565 ;
        RECT 61.475 189.975 62.940 190.145 ;
        RECT 61.475 189.725 61.645 189.975 ;
        RECT 60.685 189.555 61.645 189.725 ;
        RECT 60.685 189.385 60.855 189.555 ;
        RECT 61.815 189.385 62.120 189.805 ;
        RECT 60.525 189.175 60.855 189.385 ;
        RECT 61.025 189.175 61.465 189.385 ;
        RECT 61.635 189.175 62.120 189.385 ;
        RECT 62.310 189.375 62.600 189.805 ;
        RECT 62.770 189.770 62.940 189.975 ;
        RECT 63.110 189.950 63.350 190.735 ;
        RECT 63.520 189.770 63.850 190.565 ;
        RECT 64.195 189.925 64.490 190.735 ;
        RECT 62.770 189.595 63.850 189.770 ;
        RECT 62.770 189.545 63.555 189.595 ;
        RECT 62.310 189.175 62.700 189.375 ;
        RECT 62.870 189.175 63.215 189.375 ;
        RECT 60.045 188.835 60.805 189.005 ;
        RECT 59.130 188.185 59.405 188.665 ;
        RECT 59.575 188.355 59.875 188.685 ;
        RECT 60.135 188.185 60.305 188.665 ;
        RECT 60.475 188.365 60.805 188.835 ;
        RECT 60.975 188.185 61.145 189.005 ;
        RECT 61.315 188.835 63.015 189.005 ;
        RECT 61.315 188.370 61.645 188.835 ;
        RECT 62.630 188.745 63.015 188.835 ;
        RECT 63.385 188.905 63.555 189.545 ;
        RECT 64.670 189.425 64.915 190.565 ;
        RECT 65.090 189.925 65.350 190.735 ;
        RECT 65.950 190.730 72.225 190.735 ;
        RECT 65.530 189.425 65.780 190.560 ;
        RECT 65.950 189.935 66.210 190.730 ;
        RECT 66.380 189.835 66.640 190.560 ;
        RECT 66.810 190.005 67.070 190.730 ;
        RECT 67.240 189.835 67.500 190.560 ;
        RECT 67.670 190.005 67.930 190.730 ;
        RECT 68.100 189.835 68.360 190.560 ;
        RECT 68.530 190.005 68.790 190.730 ;
        RECT 68.960 189.835 69.220 190.560 ;
        RECT 69.390 190.005 69.635 190.730 ;
        RECT 69.805 189.835 70.065 190.560 ;
        RECT 70.250 190.005 70.495 190.730 ;
        RECT 70.665 189.835 70.925 190.560 ;
        RECT 71.110 190.005 71.355 190.730 ;
        RECT 71.525 189.835 71.785 190.560 ;
        RECT 71.970 190.005 72.225 190.730 ;
        RECT 66.380 189.820 71.785 189.835 ;
        RECT 72.395 189.820 72.685 190.560 ;
        RECT 72.855 189.990 73.125 190.735 ;
        RECT 73.475 189.990 73.745 190.735 ;
        RECT 74.375 190.730 80.650 190.735 ;
        RECT 73.915 189.820 74.205 190.560 ;
        RECT 74.375 190.005 74.630 190.730 ;
        RECT 74.815 189.835 75.075 190.560 ;
        RECT 75.245 190.005 75.490 190.730 ;
        RECT 75.675 189.835 75.935 190.560 ;
        RECT 76.105 190.005 76.350 190.730 ;
        RECT 76.535 189.835 76.795 190.560 ;
        RECT 76.965 190.005 77.210 190.730 ;
        RECT 77.380 189.835 77.640 190.560 ;
        RECT 77.810 190.005 78.070 190.730 ;
        RECT 78.240 189.835 78.500 190.560 ;
        RECT 78.670 190.005 78.930 190.730 ;
        RECT 79.100 189.835 79.360 190.560 ;
        RECT 79.530 190.005 79.790 190.730 ;
        RECT 79.960 189.835 80.220 190.560 ;
        RECT 80.390 189.935 80.650 190.730 ;
        RECT 74.815 189.820 80.220 189.835 ;
        RECT 66.380 189.595 73.125 189.820 ;
        RECT 63.755 189.075 64.015 189.425 ;
        RECT 63.385 188.735 63.930 188.905 ;
        RECT 64.185 188.865 64.500 189.425 ;
        RECT 64.670 189.175 71.790 189.425 ;
        RECT 71.960 189.375 73.125 189.595 ;
        RECT 73.475 189.595 80.220 189.820 ;
        RECT 71.960 189.205 73.155 189.375 ;
        RECT 61.815 188.185 61.985 188.655 ;
        RECT 62.245 188.395 63.430 188.565 ;
        RECT 63.600 188.355 63.930 188.735 ;
        RECT 64.185 188.185 64.490 188.695 ;
        RECT 64.670 188.365 64.920 189.175 ;
        RECT 65.090 188.185 65.350 188.710 ;
        RECT 65.530 188.365 65.780 189.175 ;
        RECT 71.960 189.005 73.125 189.205 ;
        RECT 66.380 188.835 73.125 189.005 ;
        RECT 73.475 189.005 74.640 189.595 ;
        RECT 80.820 189.425 81.070 190.560 ;
        RECT 81.250 189.925 81.510 190.735 ;
        RECT 81.685 189.425 81.930 190.565 ;
        RECT 82.110 189.925 82.405 190.735 ;
        RECT 82.585 189.570 82.875 190.735 ;
        RECT 83.105 190.035 83.325 190.565 ;
        RECT 83.495 190.225 83.825 190.735 ;
        RECT 83.995 190.035 84.220 190.565 ;
        RECT 83.105 189.770 84.220 190.035 ;
        RECT 84.390 190.020 84.705 190.565 ;
        RECT 84.895 190.320 85.225 190.735 ;
        RECT 84.390 189.790 85.225 190.020 ;
        RECT 74.810 189.175 81.930 189.425 ;
        RECT 73.475 188.835 80.220 189.005 ;
        RECT 65.950 188.185 66.210 188.745 ;
        RECT 66.380 188.380 66.640 188.835 ;
        RECT 66.810 188.185 67.070 188.665 ;
        RECT 67.240 188.380 67.500 188.835 ;
        RECT 67.670 188.185 67.930 188.665 ;
        RECT 68.100 188.380 68.360 188.835 ;
        RECT 68.530 188.185 68.775 188.665 ;
        RECT 68.945 188.380 69.220 188.835 ;
        RECT 69.390 188.185 69.635 188.665 ;
        RECT 69.805 188.380 70.065 188.835 ;
        RECT 70.245 188.185 70.495 188.665 ;
        RECT 70.665 188.380 70.925 188.835 ;
        RECT 71.105 188.185 71.355 188.665 ;
        RECT 71.525 188.380 71.785 188.835 ;
        RECT 71.965 188.185 72.225 188.665 ;
        RECT 72.395 188.380 72.655 188.835 ;
        RECT 72.825 188.185 73.125 188.665 ;
        RECT 73.475 188.185 73.775 188.665 ;
        RECT 73.945 188.380 74.205 188.835 ;
        RECT 74.375 188.185 74.635 188.665 ;
        RECT 74.815 188.380 75.075 188.835 ;
        RECT 75.245 188.185 75.495 188.665 ;
        RECT 75.675 188.380 75.935 188.835 ;
        RECT 76.105 188.185 76.355 188.665 ;
        RECT 76.535 188.380 76.795 188.835 ;
        RECT 76.965 188.185 77.210 188.665 ;
        RECT 77.380 188.380 77.655 188.835 ;
        RECT 77.825 188.185 78.070 188.665 ;
        RECT 78.240 188.380 78.500 188.835 ;
        RECT 78.670 188.185 78.930 188.665 ;
        RECT 79.100 188.380 79.360 188.835 ;
        RECT 79.530 188.185 79.790 188.665 ;
        RECT 79.960 188.380 80.220 188.835 ;
        RECT 80.390 188.185 80.650 188.745 ;
        RECT 80.820 188.365 81.070 189.175 ;
        RECT 81.250 188.185 81.510 188.710 ;
        RECT 81.680 188.365 81.930 189.175 ;
        RECT 82.100 188.865 82.415 189.425 ;
        RECT 82.110 188.185 82.415 188.695 ;
        RECT 82.585 188.185 82.875 188.910 ;
        RECT 83.055 188.850 83.370 189.425 ;
        RECT 83.045 188.185 83.375 188.665 ;
        RECT 83.560 188.465 83.940 189.425 ;
        RECT 84.390 189.095 84.715 189.510 ;
        RECT 84.885 189.095 85.225 189.790 ;
        RECT 84.885 188.925 85.055 189.095 ;
        RECT 85.395 188.925 85.625 190.565 ;
        RECT 85.795 189.765 86.085 190.735 ;
        RECT 86.270 189.935 86.525 190.735 ;
        RECT 86.725 189.885 87.055 190.565 ;
        RECT 86.270 189.395 86.515 189.755 ;
        RECT 86.705 189.605 87.055 189.885 ;
        RECT 86.705 189.225 86.875 189.605 ;
        RECT 87.235 189.425 87.430 190.475 ;
        RECT 87.610 189.595 87.930 190.735 ;
        RECT 88.105 189.645 89.315 190.735 ;
        RECT 84.315 188.755 85.055 188.925 ;
        RECT 84.315 188.355 84.505 188.755 ;
        RECT 85.225 188.735 85.625 188.925 ;
        RECT 86.355 189.055 86.875 189.225 ;
        RECT 87.045 189.095 87.430 189.425 ;
        RECT 87.610 189.375 87.870 189.425 ;
        RECT 87.610 189.205 87.875 189.375 ;
        RECT 87.610 189.095 87.870 189.205 ;
        RECT 88.105 189.105 88.625 189.645 ;
        RECT 84.725 188.185 85.055 188.545 ;
        RECT 85.225 188.355 85.415 188.735 ;
        RECT 85.585 188.185 85.915 188.565 ;
        RECT 86.355 188.490 86.525 189.055 ;
        RECT 88.795 188.935 89.315 189.475 ;
        RECT 86.715 188.715 87.930 188.885 ;
        RECT 86.715 188.410 86.945 188.715 ;
        RECT 87.115 188.185 87.445 188.545 ;
        RECT 87.640 188.365 87.930 188.715 ;
        RECT 88.105 188.185 89.315 188.935 ;
        RECT 18.100 188.015 89.400 188.185 ;
        RECT 18.185 187.265 19.395 188.015 ;
        RECT 18.185 186.725 18.705 187.265 ;
        RECT 19.570 187.175 19.830 188.015 ;
        RECT 20.005 187.270 20.260 187.845 ;
        RECT 20.430 187.635 20.760 188.015 ;
        RECT 20.975 187.465 21.145 187.845 ;
        RECT 20.430 187.295 21.145 187.465 ;
        RECT 18.875 186.555 19.395 187.095 ;
        RECT 18.185 185.465 19.395 186.555 ;
        RECT 19.570 185.465 19.830 186.615 ;
        RECT 20.005 186.540 20.175 187.270 ;
        RECT 20.430 187.105 20.600 187.295 ;
        RECT 21.405 187.215 21.715 188.015 ;
        RECT 21.920 187.215 22.615 187.845 ;
        RECT 22.785 187.275 23.275 187.845 ;
        RECT 23.445 187.445 23.675 187.845 ;
        RECT 23.845 187.615 24.265 188.015 ;
        RECT 24.435 187.445 24.605 187.845 ;
        RECT 23.445 187.275 24.605 187.445 ;
        RECT 24.775 187.275 25.225 188.015 ;
        RECT 25.395 187.275 25.835 187.835 ;
        RECT 21.920 187.165 22.095 187.215 ;
        RECT 20.345 186.775 20.600 187.105 ;
        RECT 20.430 186.565 20.600 186.775 ;
        RECT 20.880 186.745 21.235 187.115 ;
        RECT 21.415 186.775 21.750 187.045 ;
        RECT 21.920 186.615 22.090 187.165 ;
        RECT 22.260 186.775 22.595 187.025 ;
        RECT 20.005 185.635 20.260 186.540 ;
        RECT 20.430 186.395 21.145 186.565 ;
        RECT 20.430 185.465 20.760 186.225 ;
        RECT 20.975 185.635 21.145 186.395 ;
        RECT 21.405 185.465 21.685 186.605 ;
        RECT 21.855 185.635 22.185 186.615 ;
        RECT 22.785 186.605 22.955 187.275 ;
        RECT 23.125 186.775 23.530 187.105 ;
        RECT 22.355 185.465 22.615 186.605 ;
        RECT 22.785 186.435 23.555 186.605 ;
        RECT 22.795 185.465 23.125 186.265 ;
        RECT 23.305 185.805 23.555 186.435 ;
        RECT 23.745 185.975 23.995 187.105 ;
        RECT 24.195 186.775 24.440 187.105 ;
        RECT 24.625 186.825 25.015 187.105 ;
        RECT 24.195 185.975 24.395 186.775 ;
        RECT 25.185 186.655 25.355 187.105 ;
        RECT 24.565 186.485 25.355 186.655 ;
        RECT 24.565 185.805 24.735 186.485 ;
        RECT 23.305 185.635 24.735 185.805 ;
        RECT 24.905 185.465 25.220 186.315 ;
        RECT 25.525 186.265 25.835 187.275 ;
        RECT 25.395 185.635 25.835 186.265 ;
        RECT 26.925 187.275 27.265 187.845 ;
        RECT 27.460 187.350 27.630 188.015 ;
        RECT 27.910 187.675 28.130 187.720 ;
        RECT 27.905 187.505 28.130 187.675 ;
        RECT 28.300 187.535 28.745 187.705 ;
        RECT 27.910 187.365 28.130 187.505 ;
        RECT 26.925 186.305 27.100 187.275 ;
        RECT 27.910 187.195 28.405 187.365 ;
        RECT 27.270 186.655 27.440 187.105 ;
        RECT 27.610 186.825 28.060 187.025 ;
        RECT 28.230 187.000 28.405 187.195 ;
        RECT 28.575 186.745 28.745 187.535 ;
        RECT 28.915 187.410 29.165 187.780 ;
        RECT 28.995 187.025 29.165 187.410 ;
        RECT 29.335 187.375 29.585 187.780 ;
        RECT 29.755 187.545 29.925 188.015 ;
        RECT 30.095 187.375 30.435 187.780 ;
        RECT 29.335 187.195 30.435 187.375 ;
        RECT 30.625 187.205 30.865 188.015 ;
        RECT 31.035 187.205 31.365 187.845 ;
        RECT 31.535 187.205 31.805 188.015 ;
        RECT 28.995 186.855 29.190 187.025 ;
        RECT 27.270 186.485 27.665 186.655 ;
        RECT 28.575 186.605 28.850 186.745 ;
        RECT 26.925 185.635 27.185 186.305 ;
        RECT 27.495 186.215 27.665 186.485 ;
        RECT 27.835 186.385 28.850 186.605 ;
        RECT 29.020 186.605 29.190 186.855 ;
        RECT 29.360 186.775 29.920 187.025 ;
        RECT 29.020 186.215 29.575 186.605 ;
        RECT 27.495 186.045 29.575 186.215 ;
        RECT 27.355 185.465 27.685 185.865 ;
        RECT 28.555 185.465 28.955 185.865 ;
        RECT 29.245 185.810 29.575 186.045 ;
        RECT 29.745 185.675 29.920 186.775 ;
        RECT 30.090 186.455 30.435 187.025 ;
        RECT 30.605 186.775 30.955 187.025 ;
        RECT 31.125 186.605 31.295 187.205 ;
        RECT 32.025 187.195 32.255 188.015 ;
        RECT 32.425 187.215 32.755 187.845 ;
        RECT 31.465 186.775 31.815 187.025 ;
        RECT 32.005 186.775 32.335 187.025 ;
        RECT 32.505 186.615 32.755 187.215 ;
        RECT 32.925 187.195 33.135 188.015 ;
        RECT 33.370 187.275 33.625 187.845 ;
        RECT 33.795 187.615 34.125 188.015 ;
        RECT 34.550 187.480 35.080 187.845 ;
        RECT 34.550 187.445 34.725 187.480 ;
        RECT 33.795 187.275 34.725 187.445 ;
        RECT 35.270 187.335 35.545 187.845 ;
        RECT 30.615 186.435 31.295 186.605 ;
        RECT 30.090 185.465 30.435 186.285 ;
        RECT 30.615 185.650 30.945 186.435 ;
        RECT 31.475 185.465 31.805 186.605 ;
        RECT 32.025 185.465 32.255 186.605 ;
        RECT 32.425 185.635 32.755 186.615 ;
        RECT 33.370 186.605 33.540 187.275 ;
        RECT 33.795 187.105 33.965 187.275 ;
        RECT 33.710 186.775 33.965 187.105 ;
        RECT 34.190 186.775 34.385 187.105 ;
        RECT 32.925 185.465 33.135 186.605 ;
        RECT 33.370 185.635 33.705 186.605 ;
        RECT 33.875 185.465 34.045 186.605 ;
        RECT 34.215 185.805 34.385 186.775 ;
        RECT 34.555 186.145 34.725 187.275 ;
        RECT 34.895 186.485 35.065 187.285 ;
        RECT 35.265 187.165 35.545 187.335 ;
        RECT 35.270 186.685 35.545 187.165 ;
        RECT 35.715 186.485 35.905 187.845 ;
        RECT 36.085 187.480 36.595 188.015 ;
        RECT 36.815 187.205 37.060 187.810 ;
        RECT 37.510 187.275 37.765 187.845 ;
        RECT 37.935 187.615 38.265 188.015 ;
        RECT 38.690 187.480 39.220 187.845 ;
        RECT 38.690 187.445 38.865 187.480 ;
        RECT 37.935 187.275 38.865 187.445 ;
        RECT 36.105 187.035 37.335 187.205 ;
        RECT 34.895 186.315 35.905 186.485 ;
        RECT 36.075 186.470 36.825 186.660 ;
        RECT 34.555 185.975 35.680 186.145 ;
        RECT 36.075 185.805 36.245 186.470 ;
        RECT 36.995 186.225 37.335 187.035 ;
        RECT 34.215 185.635 36.245 185.805 ;
        RECT 36.415 185.465 36.585 186.225 ;
        RECT 36.820 185.815 37.335 186.225 ;
        RECT 37.510 186.605 37.680 187.275 ;
        RECT 37.935 187.105 38.105 187.275 ;
        RECT 37.850 186.775 38.105 187.105 ;
        RECT 38.330 186.775 38.525 187.105 ;
        RECT 37.510 185.635 37.845 186.605 ;
        RECT 38.015 185.465 38.185 186.605 ;
        RECT 38.355 185.805 38.525 186.775 ;
        RECT 38.695 186.145 38.865 187.275 ;
        RECT 39.035 186.485 39.205 187.285 ;
        RECT 39.410 186.995 39.685 187.845 ;
        RECT 39.405 186.825 39.685 186.995 ;
        RECT 39.410 186.685 39.685 186.825 ;
        RECT 39.855 186.485 40.045 187.845 ;
        RECT 40.225 187.480 40.735 188.015 ;
        RECT 40.955 187.205 41.200 187.810 ;
        RECT 42.195 187.465 42.365 187.845 ;
        RECT 42.580 187.635 42.910 188.015 ;
        RECT 42.195 187.295 42.910 187.465 ;
        RECT 40.245 187.035 41.475 187.205 ;
        RECT 39.035 186.315 40.045 186.485 ;
        RECT 40.215 186.470 40.965 186.660 ;
        RECT 38.695 185.975 39.820 186.145 ;
        RECT 40.215 185.805 40.385 186.470 ;
        RECT 41.135 186.225 41.475 187.035 ;
        RECT 42.105 186.745 42.460 187.115 ;
        RECT 42.740 187.105 42.910 187.295 ;
        RECT 43.080 187.270 43.335 187.845 ;
        RECT 42.740 186.775 42.995 187.105 ;
        RECT 42.740 186.565 42.910 186.775 ;
        RECT 38.355 185.635 40.385 185.805 ;
        RECT 40.555 185.465 40.725 186.225 ;
        RECT 40.960 185.815 41.475 186.225 ;
        RECT 42.195 186.395 42.910 186.565 ;
        RECT 43.165 186.540 43.335 187.270 ;
        RECT 43.510 187.175 43.770 188.015 ;
        RECT 43.945 187.290 44.235 188.015 ;
        RECT 44.455 187.215 44.665 188.015 ;
        RECT 42.195 185.635 42.365 186.395 ;
        RECT 42.580 185.465 42.910 186.225 ;
        RECT 43.080 185.635 43.335 186.540 ;
        RECT 43.510 185.465 43.770 186.615 ;
        RECT 43.945 185.465 44.235 186.630 ;
        RECT 44.455 185.465 44.665 186.605 ;
        RECT 44.835 185.635 45.175 187.845 ;
        RECT 45.355 187.555 45.605 188.015 ;
        RECT 45.795 187.385 46.125 187.845 ;
        RECT 46.325 187.675 46.710 187.845 ;
        RECT 46.305 187.505 46.710 187.675 ;
        RECT 45.350 187.215 46.125 187.385 ;
        RECT 45.350 186.315 45.625 187.215 ;
        RECT 45.825 186.485 46.155 187.025 ;
        RECT 46.325 186.485 46.710 187.505 ;
        RECT 47.185 187.475 47.515 187.845 ;
        RECT 47.705 187.645 48.035 188.015 ;
        RECT 48.205 187.475 48.535 187.845 ;
        RECT 47.185 187.275 48.535 187.475 ;
        RECT 49.005 187.215 49.700 187.845 ;
        RECT 49.905 187.215 50.215 188.015 ;
        RECT 50.470 187.465 50.800 187.845 ;
        RECT 50.970 187.635 52.155 187.805 ;
        RECT 52.415 187.545 52.585 188.015 ;
        RECT 50.470 187.295 51.015 187.465 ;
        RECT 47.000 186.485 47.420 187.025 ;
        RECT 47.620 186.775 47.980 187.105 ;
        RECT 48.150 186.785 48.835 187.095 ;
        RECT 45.350 186.075 47.515 186.315 ;
        RECT 45.355 185.465 45.975 185.905 ;
        RECT 46.180 185.635 46.460 186.075 ;
        RECT 46.645 185.465 46.975 185.845 ;
        RECT 47.185 185.635 47.515 186.075 ;
        RECT 47.690 185.975 47.980 186.775 ;
        RECT 47.685 185.805 47.980 185.975 ;
        RECT 47.690 185.730 47.980 185.805 ;
        RECT 48.205 185.465 48.460 186.605 ;
        RECT 48.630 185.745 48.835 186.785 ;
        RECT 49.025 186.775 49.360 187.025 ;
        RECT 49.530 186.615 49.700 187.215 ;
        RECT 49.870 186.775 50.205 187.045 ;
        RECT 50.385 186.775 50.645 187.125 ;
        RECT 50.845 186.655 51.015 187.295 ;
        RECT 51.385 187.365 51.770 187.455 ;
        RECT 52.755 187.365 53.085 187.830 ;
        RECT 51.385 187.195 53.085 187.365 ;
        RECT 53.255 187.195 53.425 188.015 ;
        RECT 53.595 187.365 53.925 187.835 ;
        RECT 54.095 187.535 54.265 188.015 ;
        RECT 54.535 187.675 55.725 187.845 ;
        RECT 54.535 187.505 54.845 187.675 ;
        RECT 53.595 187.195 54.355 187.365 ;
        RECT 51.185 186.825 51.530 187.025 ;
        RECT 51.700 186.825 52.090 187.025 ;
        RECT 49.005 185.465 49.265 186.605 ;
        RECT 49.435 185.635 49.765 186.615 ;
        RECT 50.845 186.605 51.630 186.655 ;
        RECT 49.935 185.465 50.215 186.605 ;
        RECT 50.550 186.430 51.630 186.605 ;
        RECT 50.550 185.635 50.880 186.430 ;
        RECT 51.050 185.465 51.290 186.250 ;
        RECT 51.460 186.225 51.630 186.430 ;
        RECT 51.800 186.395 52.090 186.825 ;
        RECT 52.280 186.815 52.765 187.025 ;
        RECT 52.935 186.815 53.375 187.025 ;
        RECT 53.545 186.815 53.875 187.025 ;
        RECT 52.280 186.395 52.585 186.815 ;
        RECT 53.545 186.645 53.715 186.815 ;
        RECT 52.755 186.475 53.715 186.645 ;
        RECT 52.755 186.225 52.925 186.475 ;
        RECT 51.460 186.055 52.925 186.225 ;
        RECT 51.850 185.635 52.605 186.055 ;
        RECT 53.095 185.465 53.425 186.305 ;
        RECT 54.045 186.225 54.355 187.195 ;
        RECT 54.530 186.700 54.845 187.335 ;
        RECT 53.595 186.055 54.355 186.225 ;
        RECT 53.595 185.635 53.845 186.055 ;
        RECT 54.015 185.465 54.355 185.885 ;
        RECT 54.535 185.465 54.845 186.530 ;
        RECT 55.015 186.315 55.225 187.505 ;
        RECT 55.395 187.385 55.725 187.675 ;
        RECT 55.965 187.555 56.135 188.015 ;
        RECT 56.365 187.385 56.695 187.845 ;
        RECT 56.875 187.555 57.045 188.015 ;
        RECT 57.225 187.385 57.555 187.845 ;
        RECT 57.805 187.535 58.085 188.015 ;
        RECT 55.395 187.215 57.555 187.385 ;
        RECT 58.255 187.365 58.515 187.755 ;
        RECT 58.690 187.535 58.945 188.015 ;
        RECT 59.115 187.365 59.410 187.755 ;
        RECT 59.590 187.535 59.865 188.015 ;
        RECT 60.035 187.515 60.335 187.845 ;
        RECT 60.595 187.535 60.895 188.015 ;
        RECT 57.760 187.195 59.410 187.365 ;
        RECT 55.565 186.655 56.060 187.025 ;
        RECT 56.240 186.825 57.040 187.025 ;
        RECT 57.210 186.655 57.540 187.045 ;
        RECT 55.505 186.485 57.540 186.655 ;
        RECT 57.760 186.685 58.165 187.195 ;
        RECT 58.335 186.855 59.475 187.025 ;
        RECT 57.760 186.515 58.515 186.685 ;
        RECT 55.015 186.135 56.665 186.315 ;
        RECT 55.015 185.635 55.250 186.135 ;
        RECT 56.365 185.975 56.665 186.135 ;
        RECT 55.420 185.465 55.750 185.925 ;
        RECT 55.945 185.805 56.135 185.965 ;
        RECT 56.835 185.805 57.055 186.315 ;
        RECT 55.945 185.635 57.055 185.805 ;
        RECT 57.225 185.465 57.555 186.315 ;
        RECT 57.800 185.465 58.085 186.335 ;
        RECT 58.255 186.265 58.515 186.515 ;
        RECT 59.305 186.605 59.475 186.855 ;
        RECT 59.645 186.775 59.995 187.345 ;
        RECT 60.165 186.605 60.335 187.515 ;
        RECT 61.065 187.365 61.325 187.820 ;
        RECT 61.495 187.535 61.755 188.015 ;
        RECT 61.935 187.365 62.195 187.820 ;
        RECT 62.365 187.535 62.615 188.015 ;
        RECT 62.795 187.365 63.055 187.820 ;
        RECT 63.225 187.535 63.475 188.015 ;
        RECT 63.655 187.365 63.915 187.820 ;
        RECT 64.085 187.535 64.330 188.015 ;
        RECT 64.500 187.365 64.775 187.820 ;
        RECT 64.945 187.535 65.190 188.015 ;
        RECT 65.360 187.365 65.620 187.820 ;
        RECT 65.790 187.535 66.050 188.015 ;
        RECT 66.220 187.365 66.480 187.820 ;
        RECT 66.650 187.535 66.910 188.015 ;
        RECT 67.080 187.365 67.340 187.820 ;
        RECT 67.510 187.455 67.770 188.015 ;
        RECT 59.305 186.435 60.335 186.605 ;
        RECT 58.255 186.095 59.375 186.265 ;
        RECT 58.255 185.635 58.515 186.095 ;
        RECT 58.690 185.465 58.945 185.925 ;
        RECT 59.115 185.635 59.375 186.095 ;
        RECT 59.545 185.465 59.855 186.265 ;
        RECT 60.025 185.635 60.335 186.435 ;
        RECT 60.595 187.195 67.340 187.365 ;
        RECT 60.595 186.605 61.760 187.195 ;
        RECT 67.940 187.025 68.190 187.835 ;
        RECT 68.370 187.490 68.630 188.015 ;
        RECT 68.800 187.025 69.050 187.835 ;
        RECT 69.230 187.505 69.535 188.015 ;
        RECT 61.930 186.775 69.050 187.025 ;
        RECT 69.220 186.775 69.535 187.335 ;
        RECT 69.705 187.290 69.995 188.015 ;
        RECT 70.190 187.190 70.445 188.015 ;
        RECT 70.615 187.275 70.950 187.845 ;
        RECT 71.145 187.350 71.315 188.015 ;
        RECT 71.595 187.365 71.815 187.720 ;
        RECT 71.985 187.535 72.445 187.705 ;
        RECT 71.595 187.330 72.100 187.365 ;
        RECT 60.595 186.380 67.340 186.605 ;
        RECT 60.595 185.465 60.865 186.210 ;
        RECT 61.035 185.640 61.325 186.380 ;
        RECT 61.935 186.365 67.340 186.380 ;
        RECT 61.495 185.470 61.750 186.195 ;
        RECT 61.935 185.640 62.195 186.365 ;
        RECT 62.365 185.470 62.610 186.195 ;
        RECT 62.795 185.640 63.055 186.365 ;
        RECT 63.225 185.470 63.470 186.195 ;
        RECT 63.655 185.640 63.915 186.365 ;
        RECT 64.085 185.470 64.330 186.195 ;
        RECT 64.500 185.640 64.760 186.365 ;
        RECT 64.930 185.470 65.190 186.195 ;
        RECT 65.360 185.640 65.620 186.365 ;
        RECT 65.790 185.470 66.050 186.195 ;
        RECT 66.220 185.640 66.480 186.365 ;
        RECT 66.650 185.470 66.910 186.195 ;
        RECT 67.080 185.640 67.340 186.365 ;
        RECT 67.510 185.470 67.770 186.265 ;
        RECT 67.940 185.640 68.190 186.775 ;
        RECT 61.495 185.465 67.770 185.470 ;
        RECT 68.370 185.465 68.630 186.275 ;
        RECT 68.805 185.635 69.050 186.775 ;
        RECT 69.230 185.465 69.525 186.275 ;
        RECT 69.705 185.465 69.995 186.630 ;
        RECT 70.190 185.465 70.445 186.690 ;
        RECT 70.615 186.315 70.785 187.275 ;
        RECT 71.595 187.195 72.105 187.330 ;
        RECT 70.955 186.655 71.125 187.105 ;
        RECT 71.295 186.825 71.765 187.025 ;
        RECT 71.935 187.000 72.105 187.195 ;
        RECT 72.275 186.745 72.445 187.535 ;
        RECT 72.615 187.410 72.860 187.780 ;
        RECT 72.690 187.025 72.860 187.410 ;
        RECT 73.035 187.375 73.265 187.780 ;
        RECT 73.455 187.545 73.625 188.015 ;
        RECT 73.795 187.375 74.125 187.780 ;
        RECT 73.035 187.195 74.125 187.375 ;
        RECT 74.305 187.215 74.595 188.015 ;
        RECT 74.765 187.555 75.315 187.845 ;
        RECT 75.485 187.555 75.735 188.015 ;
        RECT 72.690 186.855 72.880 187.025 ;
        RECT 70.955 186.485 71.350 186.655 ;
        RECT 72.275 186.605 72.540 186.745 ;
        RECT 70.615 186.305 70.855 186.315 ;
        RECT 70.615 185.635 70.870 186.305 ;
        RECT 71.180 186.215 71.350 186.485 ;
        RECT 71.520 186.385 72.540 186.605 ;
        RECT 72.710 186.605 72.880 186.855 ;
        RECT 73.050 186.775 73.605 187.025 ;
        RECT 72.710 186.215 73.265 186.605 ;
        RECT 71.180 186.045 73.265 186.215 ;
        RECT 71.040 185.465 71.370 185.865 ;
        RECT 72.240 185.465 72.645 185.865 ;
        RECT 72.915 185.675 73.265 186.045 ;
        RECT 73.435 185.975 73.605 186.775 ;
        RECT 73.780 186.455 74.125 187.025 ;
        RECT 73.435 185.805 73.615 185.975 ;
        RECT 73.435 185.675 73.605 185.805 ;
        RECT 73.810 185.465 74.125 186.285 ;
        RECT 74.305 185.465 74.595 186.605 ;
        RECT 74.765 186.185 75.015 187.555 ;
        RECT 76.365 187.385 76.695 187.745 ;
        RECT 77.155 187.535 77.455 188.015 ;
        RECT 75.305 187.195 76.695 187.385 ;
        RECT 77.625 187.365 77.885 187.820 ;
        RECT 78.055 187.535 78.315 188.015 ;
        RECT 78.495 187.365 78.755 187.820 ;
        RECT 78.925 187.535 79.175 188.015 ;
        RECT 79.355 187.365 79.615 187.820 ;
        RECT 79.785 187.535 80.035 188.015 ;
        RECT 80.215 187.365 80.475 187.820 ;
        RECT 80.645 187.535 80.890 188.015 ;
        RECT 81.060 187.365 81.335 187.820 ;
        RECT 81.505 187.535 81.750 188.015 ;
        RECT 81.920 187.365 82.180 187.820 ;
        RECT 82.350 187.535 82.610 188.015 ;
        RECT 82.780 187.365 83.040 187.820 ;
        RECT 83.210 187.535 83.470 188.015 ;
        RECT 83.640 187.365 83.900 187.820 ;
        RECT 84.070 187.455 84.330 188.015 ;
        RECT 77.155 187.195 83.900 187.365 ;
        RECT 75.305 187.105 75.475 187.195 ;
        RECT 75.185 186.775 75.475 187.105 ;
        RECT 75.645 186.775 75.975 187.025 ;
        RECT 76.205 186.775 76.895 187.025 ;
        RECT 75.305 186.525 75.475 186.775 ;
        RECT 75.305 186.355 76.245 186.525 ;
        RECT 74.765 185.635 75.215 186.185 ;
        RECT 75.405 185.465 75.735 186.185 ;
        RECT 75.945 185.805 76.245 186.355 ;
        RECT 76.580 186.335 76.895 186.775 ;
        RECT 77.155 186.605 78.320 187.195 ;
        RECT 84.500 187.025 84.750 187.835 ;
        RECT 84.930 187.490 85.190 188.015 ;
        RECT 85.360 187.025 85.610 187.835 ;
        RECT 85.790 187.505 86.095 188.015 ;
        RECT 86.270 187.615 86.605 188.015 ;
        RECT 86.775 187.445 86.980 187.845 ;
        RECT 87.190 187.535 87.465 188.015 ;
        RECT 87.675 187.515 87.935 187.845 ;
        RECT 78.490 186.775 85.610 187.025 ;
        RECT 85.780 186.775 86.095 187.335 ;
        RECT 86.295 187.275 86.980 187.445 ;
        RECT 77.155 186.380 83.900 186.605 ;
        RECT 76.415 185.465 76.695 186.135 ;
        RECT 77.155 185.465 77.425 186.210 ;
        RECT 77.595 185.640 77.885 186.380 ;
        RECT 78.495 186.365 83.900 186.380 ;
        RECT 78.055 185.470 78.310 186.195 ;
        RECT 78.495 185.640 78.755 186.365 ;
        RECT 78.925 185.470 79.170 186.195 ;
        RECT 79.355 185.640 79.615 186.365 ;
        RECT 79.785 185.470 80.030 186.195 ;
        RECT 80.215 185.640 80.475 186.365 ;
        RECT 80.645 185.470 80.890 186.195 ;
        RECT 81.060 185.640 81.320 186.365 ;
        RECT 81.490 185.470 81.750 186.195 ;
        RECT 81.920 185.640 82.180 186.365 ;
        RECT 82.350 185.470 82.610 186.195 ;
        RECT 82.780 185.640 83.040 186.365 ;
        RECT 83.210 185.470 83.470 186.195 ;
        RECT 83.640 185.640 83.900 186.365 ;
        RECT 84.070 185.470 84.330 186.265 ;
        RECT 84.500 185.640 84.750 186.775 ;
        RECT 78.055 185.465 84.330 185.470 ;
        RECT 84.930 185.465 85.190 186.275 ;
        RECT 85.365 185.635 85.610 186.775 ;
        RECT 85.790 185.465 86.085 186.275 ;
        RECT 86.295 186.245 86.635 187.275 ;
        RECT 86.805 186.605 87.055 187.105 ;
        RECT 87.235 186.775 87.595 187.355 ;
        RECT 87.765 186.605 87.935 187.515 ;
        RECT 88.105 187.265 89.315 188.015 ;
        RECT 86.805 186.435 87.935 186.605 ;
        RECT 86.295 186.070 86.960 186.245 ;
        RECT 86.270 185.465 86.605 185.890 ;
        RECT 86.775 185.665 86.960 186.070 ;
        RECT 87.165 185.465 87.495 186.245 ;
        RECT 87.665 185.665 87.935 186.435 ;
        RECT 88.105 186.555 88.625 187.095 ;
        RECT 88.795 186.725 89.315 187.265 ;
        RECT 88.105 185.465 89.315 186.555 ;
        RECT 18.100 185.295 89.400 185.465 ;
        RECT 18.185 184.205 19.395 185.295 ;
        RECT 18.185 183.495 18.705 184.035 ;
        RECT 18.875 183.665 19.395 184.205 ;
        RECT 19.645 184.365 19.825 185.125 ;
        RECT 20.005 184.535 20.335 185.295 ;
        RECT 19.645 184.195 20.320 184.365 ;
        RECT 20.505 184.220 20.775 185.125 ;
        RECT 20.150 184.050 20.320 184.195 ;
        RECT 19.585 183.645 19.925 184.015 ;
        RECT 20.150 183.720 20.425 184.050 ;
        RECT 18.185 182.745 19.395 183.495 ;
        RECT 20.150 183.465 20.320 183.720 ;
        RECT 19.655 183.295 20.320 183.465 ;
        RECT 20.595 183.420 20.775 184.220 ;
        RECT 21.405 184.155 21.685 185.295 ;
        RECT 21.855 184.145 22.185 185.125 ;
        RECT 22.355 184.155 22.615 185.295 ;
        RECT 22.795 184.495 23.125 185.295 ;
        RECT 23.305 184.955 24.735 185.125 ;
        RECT 23.305 184.325 23.555 184.955 ;
        RECT 22.785 184.155 23.555 184.325 ;
        RECT 21.920 184.105 22.095 184.145 ;
        RECT 21.415 183.715 21.750 183.985 ;
        RECT 21.920 183.545 22.090 184.105 ;
        RECT 22.260 183.735 22.595 183.985 ;
        RECT 19.655 182.915 19.825 183.295 ;
        RECT 20.005 182.745 20.335 183.125 ;
        RECT 20.515 182.915 20.775 183.420 ;
        RECT 21.405 182.745 21.715 183.545 ;
        RECT 21.920 182.915 22.615 183.545 ;
        RECT 22.785 183.485 22.955 184.155 ;
        RECT 23.125 183.655 23.530 183.985 ;
        RECT 23.745 183.655 23.995 184.785 ;
        RECT 24.195 183.985 24.395 184.785 ;
        RECT 24.565 184.275 24.735 184.955 ;
        RECT 24.905 184.445 25.220 185.295 ;
        RECT 25.395 184.495 25.835 185.125 ;
        RECT 24.565 184.105 25.355 184.275 ;
        RECT 24.195 183.655 24.440 183.985 ;
        RECT 24.625 183.655 25.015 183.935 ;
        RECT 25.185 183.655 25.355 184.105 ;
        RECT 25.525 183.485 25.835 184.495 ;
        RECT 22.785 182.915 23.275 183.485 ;
        RECT 23.445 183.315 24.605 183.485 ;
        RECT 23.445 182.915 23.675 183.315 ;
        RECT 23.845 182.745 24.265 183.145 ;
        RECT 24.435 182.915 24.605 183.315 ;
        RECT 24.775 182.745 25.225 183.485 ;
        RECT 25.395 182.925 25.835 183.485 ;
        RECT 26.465 184.455 26.725 185.125 ;
        RECT 26.895 184.895 27.225 185.295 ;
        RECT 28.095 184.895 28.495 185.295 ;
        RECT 28.785 184.715 29.115 184.950 ;
        RECT 27.035 184.545 29.115 184.715 ;
        RECT 26.465 184.445 26.695 184.455 ;
        RECT 26.465 183.485 26.640 184.445 ;
        RECT 27.035 184.275 27.205 184.545 ;
        RECT 26.810 184.105 27.205 184.275 ;
        RECT 27.375 184.155 28.390 184.375 ;
        RECT 26.810 183.655 26.980 184.105 ;
        RECT 28.115 184.015 28.390 184.155 ;
        RECT 28.560 184.155 29.115 184.545 ;
        RECT 27.150 183.735 27.600 183.935 ;
        RECT 27.770 183.565 27.945 183.760 ;
        RECT 26.465 182.915 26.805 183.485 ;
        RECT 27.000 182.745 27.170 183.410 ;
        RECT 27.450 183.395 27.945 183.565 ;
        RECT 27.450 183.255 27.670 183.395 ;
        RECT 27.445 183.085 27.670 183.255 ;
        RECT 28.115 183.225 28.285 184.015 ;
        RECT 28.560 183.905 28.730 184.155 ;
        RECT 29.285 183.985 29.460 185.085 ;
        RECT 29.630 184.475 29.975 185.295 ;
        RECT 28.535 183.735 28.730 183.905 ;
        RECT 28.900 183.735 29.460 183.985 ;
        RECT 29.630 183.735 29.975 184.305 ;
        RECT 31.065 184.130 31.355 185.295 ;
        RECT 31.525 184.220 31.795 185.125 ;
        RECT 31.965 184.535 32.295 185.295 ;
        RECT 32.475 184.365 32.655 185.125 ;
        RECT 28.535 183.350 28.705 183.735 ;
        RECT 27.450 183.040 27.670 183.085 ;
        RECT 27.840 183.055 28.285 183.225 ;
        RECT 28.455 182.980 28.705 183.350 ;
        RECT 28.875 183.385 29.975 183.565 ;
        RECT 28.875 182.980 29.125 183.385 ;
        RECT 29.295 182.745 29.465 183.215 ;
        RECT 29.635 182.980 29.975 183.385 ;
        RECT 31.065 182.745 31.355 183.470 ;
        RECT 31.525 183.420 31.705 184.220 ;
        RECT 31.980 184.195 32.655 184.365 ;
        RECT 31.980 184.050 32.150 184.195 ;
        RECT 31.875 183.720 32.150 184.050 ;
        RECT 32.910 184.155 33.245 185.125 ;
        RECT 33.415 184.155 33.585 185.295 ;
        RECT 33.755 184.955 35.785 185.125 ;
        RECT 31.980 183.465 32.150 183.720 ;
        RECT 32.375 183.645 32.715 184.015 ;
        RECT 32.910 183.485 33.080 184.155 ;
        RECT 33.755 183.985 33.925 184.955 ;
        RECT 33.250 183.655 33.505 183.985 ;
        RECT 33.730 183.655 33.925 183.985 ;
        RECT 34.095 184.615 35.220 184.785 ;
        RECT 33.335 183.485 33.505 183.655 ;
        RECT 34.095 183.485 34.265 184.615 ;
        RECT 31.525 182.915 31.785 183.420 ;
        RECT 31.980 183.295 32.645 183.465 ;
        RECT 31.965 182.745 32.295 183.125 ;
        RECT 32.475 182.915 32.645 183.295 ;
        RECT 32.910 182.915 33.165 183.485 ;
        RECT 33.335 183.315 34.265 183.485 ;
        RECT 34.435 184.275 35.445 184.445 ;
        RECT 34.435 183.475 34.605 184.275 ;
        RECT 34.810 183.595 35.085 184.075 ;
        RECT 34.805 183.425 35.085 183.595 ;
        RECT 34.090 183.280 34.265 183.315 ;
        RECT 33.335 182.745 33.665 183.145 ;
        RECT 34.090 182.915 34.620 183.280 ;
        RECT 34.810 182.915 35.085 183.425 ;
        RECT 35.255 182.915 35.445 184.275 ;
        RECT 35.615 184.290 35.785 184.955 ;
        RECT 35.955 184.535 36.125 185.295 ;
        RECT 36.360 184.535 36.875 184.945 ;
        RECT 35.615 184.100 36.365 184.290 ;
        RECT 36.535 183.725 36.875 184.535 ;
        RECT 37.135 184.365 37.305 185.125 ;
        RECT 37.485 184.535 37.815 185.295 ;
        RECT 37.135 184.195 37.800 184.365 ;
        RECT 37.985 184.220 38.255 185.125 ;
        RECT 37.630 184.050 37.800 184.195 ;
        RECT 35.645 183.555 36.875 183.725 ;
        RECT 37.065 183.645 37.395 184.015 ;
        RECT 37.630 183.720 37.915 184.050 ;
        RECT 35.625 182.745 36.135 183.280 ;
        RECT 36.355 182.950 36.600 183.555 ;
        RECT 37.630 183.465 37.800 183.720 ;
        RECT 37.135 183.295 37.800 183.465 ;
        RECT 38.085 183.420 38.255 184.220 ;
        RECT 37.135 182.915 37.305 183.295 ;
        RECT 37.485 182.745 37.815 183.125 ;
        RECT 37.995 182.915 38.255 183.420 ;
        RECT 38.885 184.220 39.155 185.125 ;
        RECT 39.325 184.535 39.655 185.295 ;
        RECT 39.835 184.365 40.015 185.125 ;
        RECT 38.885 183.420 39.065 184.220 ;
        RECT 39.340 184.195 40.015 184.365 ;
        RECT 41.205 184.405 41.465 185.115 ;
        RECT 41.635 184.585 41.965 185.295 ;
        RECT 42.135 184.405 42.365 185.115 ;
        RECT 39.340 184.050 39.510 184.195 ;
        RECT 41.205 184.165 42.365 184.405 ;
        RECT 42.545 184.385 42.815 185.115 ;
        RECT 42.995 184.565 43.335 185.295 ;
        RECT 42.545 184.165 43.315 184.385 ;
        RECT 39.235 183.720 39.510 184.050 ;
        RECT 39.340 183.465 39.510 183.720 ;
        RECT 39.735 183.645 40.075 184.015 ;
        RECT 41.195 183.655 41.495 183.985 ;
        RECT 41.675 183.675 42.200 183.985 ;
        RECT 42.380 183.675 42.845 183.985 ;
        RECT 38.885 182.915 39.145 183.420 ;
        RECT 39.340 183.295 40.005 183.465 ;
        RECT 39.325 182.745 39.655 183.125 ;
        RECT 39.835 182.915 40.005 183.295 ;
        RECT 41.205 182.745 41.495 183.475 ;
        RECT 41.675 183.035 41.905 183.675 ;
        RECT 43.025 183.495 43.315 184.165 ;
        RECT 42.085 183.295 43.315 183.495 ;
        RECT 42.085 182.925 42.395 183.295 ;
        RECT 42.575 182.745 43.245 183.115 ;
        RECT 43.505 182.925 43.765 185.115 ;
        RECT 44.405 184.875 44.745 185.295 ;
        RECT 44.915 184.705 45.165 185.125 ;
        RECT 44.405 184.535 45.165 184.705 ;
        RECT 44.405 183.565 44.715 184.535 ;
        RECT 45.335 184.455 45.665 185.295 ;
        RECT 46.155 184.705 46.910 185.125 ;
        RECT 45.835 184.535 47.300 184.705 ;
        RECT 45.835 184.285 46.005 184.535 ;
        RECT 45.045 184.115 46.005 184.285 ;
        RECT 45.045 183.945 45.215 184.115 ;
        RECT 46.175 183.945 46.480 184.365 ;
        RECT 44.885 183.735 45.215 183.945 ;
        RECT 45.385 183.735 45.825 183.945 ;
        RECT 45.995 183.735 46.480 183.945 ;
        RECT 46.670 183.935 46.960 184.365 ;
        RECT 47.130 184.330 47.300 184.535 ;
        RECT 47.470 184.510 47.710 185.295 ;
        RECT 47.880 184.330 48.210 185.125 ;
        RECT 47.130 184.155 48.210 184.330 ;
        RECT 47.130 184.105 47.915 184.155 ;
        RECT 46.670 183.735 47.060 183.935 ;
        RECT 47.230 183.735 47.575 183.935 ;
        RECT 44.405 183.395 45.165 183.565 ;
        RECT 44.495 182.745 44.665 183.225 ;
        RECT 44.835 182.925 45.165 183.395 ;
        RECT 45.335 182.745 45.505 183.565 ;
        RECT 45.675 183.395 47.375 183.565 ;
        RECT 45.675 182.930 46.005 183.395 ;
        RECT 46.990 183.305 47.375 183.395 ;
        RECT 47.745 183.465 47.915 184.105 ;
        RECT 48.115 183.635 48.375 183.985 ;
        RECT 47.745 183.295 48.290 183.465 ;
        RECT 46.175 182.745 46.345 183.215 ;
        RECT 46.605 182.955 47.790 183.125 ;
        RECT 47.960 182.915 48.290 183.295 ;
        RECT 49.465 183.025 49.745 185.125 ;
        RECT 49.935 184.535 50.720 185.295 ;
        RECT 51.115 184.465 51.500 185.125 ;
        RECT 51.115 184.365 51.525 184.465 ;
        RECT 49.915 184.155 51.525 184.365 ;
        RECT 51.825 184.275 52.025 185.065 ;
        RECT 49.915 183.555 50.190 184.155 ;
        RECT 51.695 184.105 52.025 184.275 ;
        RECT 52.195 184.115 52.515 185.295 ;
        RECT 52.695 184.685 53.025 185.115 ;
        RECT 53.205 184.855 53.400 185.295 ;
        RECT 53.570 184.685 53.900 185.115 ;
        RECT 52.695 184.515 53.900 184.685 ;
        RECT 52.695 184.185 53.590 184.515 ;
        RECT 54.070 184.345 54.345 185.115 ;
        RECT 54.630 184.495 54.885 185.295 ;
        RECT 53.760 184.155 54.345 184.345 ;
        RECT 55.055 184.325 55.385 185.125 ;
        RECT 55.555 184.495 55.725 185.295 ;
        RECT 55.895 184.325 56.225 185.125 ;
        RECT 54.525 184.155 56.225 184.325 ;
        RECT 56.395 184.155 56.655 185.295 ;
        RECT 51.695 183.985 51.875 184.105 ;
        RECT 50.360 183.735 50.715 183.985 ;
        RECT 50.910 183.935 51.375 183.985 ;
        RECT 50.905 183.765 51.375 183.935 ;
        RECT 50.910 183.735 51.375 183.765 ;
        RECT 51.545 183.735 51.875 183.985 ;
        RECT 52.050 183.735 52.515 183.935 ;
        RECT 52.700 183.655 52.995 183.985 ;
        RECT 53.175 183.655 53.590 183.985 ;
        RECT 49.915 183.375 51.165 183.555 ;
        RECT 50.800 183.305 51.165 183.375 ;
        RECT 51.335 183.355 52.515 183.525 ;
        RECT 49.975 182.745 50.145 183.205 ;
        RECT 51.335 183.135 51.665 183.355 ;
        RECT 50.415 182.955 51.665 183.135 ;
        RECT 51.835 182.745 52.005 183.185 ;
        RECT 52.175 182.940 52.515 183.355 ;
        RECT 52.695 182.745 52.995 183.475 ;
        RECT 53.175 183.035 53.405 183.655 ;
        RECT 53.760 183.485 53.935 184.155 ;
        RECT 53.605 183.305 53.935 183.485 ;
        RECT 54.105 183.335 54.345 183.985 ;
        RECT 54.525 183.565 54.805 184.155 ;
        RECT 56.825 184.130 57.115 185.295 ;
        RECT 57.375 184.550 57.645 185.295 ;
        RECT 58.275 185.290 64.550 185.295 ;
        RECT 57.815 184.380 58.105 185.120 ;
        RECT 58.275 184.565 58.530 185.290 ;
        RECT 58.715 184.395 58.975 185.120 ;
        RECT 59.145 184.565 59.390 185.290 ;
        RECT 59.575 184.395 59.835 185.120 ;
        RECT 60.005 184.565 60.250 185.290 ;
        RECT 60.435 184.395 60.695 185.120 ;
        RECT 60.865 184.565 61.110 185.290 ;
        RECT 61.280 184.395 61.540 185.120 ;
        RECT 61.710 184.565 61.970 185.290 ;
        RECT 62.140 184.395 62.400 185.120 ;
        RECT 62.570 184.565 62.830 185.290 ;
        RECT 63.000 184.395 63.260 185.120 ;
        RECT 63.430 184.565 63.690 185.290 ;
        RECT 63.860 184.395 64.120 185.120 ;
        RECT 64.290 184.495 64.550 185.290 ;
        RECT 58.715 184.380 64.120 184.395 ;
        RECT 57.375 184.155 64.120 184.380 ;
        RECT 54.975 183.735 55.725 183.985 ;
        RECT 55.895 183.735 56.655 183.985 ;
        RECT 57.375 183.565 58.540 184.155 ;
        RECT 64.720 183.985 64.970 185.120 ;
        RECT 65.150 184.485 65.410 185.295 ;
        RECT 65.585 183.985 65.830 185.125 ;
        RECT 66.010 184.485 66.305 185.295 ;
        RECT 66.540 184.425 66.825 185.295 ;
        RECT 66.995 184.665 67.255 185.125 ;
        RECT 67.430 184.835 67.685 185.295 ;
        RECT 67.855 184.665 68.115 185.125 ;
        RECT 66.995 184.495 68.115 184.665 ;
        RECT 68.285 184.495 68.595 185.295 ;
        RECT 66.995 184.245 67.255 184.495 ;
        RECT 68.765 184.325 69.075 185.125 ;
        RECT 69.255 184.485 69.550 185.295 ;
        RECT 66.500 184.075 67.255 184.245 ;
        RECT 68.045 184.155 69.075 184.325 ;
        RECT 58.710 183.735 65.830 183.985 ;
        RECT 54.525 183.315 55.385 183.565 ;
        RECT 55.555 183.375 56.655 183.545 ;
        RECT 53.605 182.925 53.830 183.305 ;
        RECT 54.000 182.745 54.330 183.135 ;
        RECT 54.635 183.125 54.965 183.145 ;
        RECT 55.555 183.125 55.805 183.375 ;
        RECT 54.635 182.915 55.805 183.125 ;
        RECT 55.975 182.745 56.145 183.205 ;
        RECT 56.315 182.915 56.655 183.375 ;
        RECT 56.825 182.745 57.115 183.470 ;
        RECT 57.375 183.395 64.120 183.565 ;
        RECT 57.375 182.745 57.675 183.225 ;
        RECT 57.845 182.940 58.105 183.395 ;
        RECT 58.275 182.745 58.535 183.225 ;
        RECT 58.715 182.940 58.975 183.395 ;
        RECT 59.145 182.745 59.395 183.225 ;
        RECT 59.575 182.940 59.835 183.395 ;
        RECT 60.005 182.745 60.255 183.225 ;
        RECT 60.435 182.940 60.695 183.395 ;
        RECT 60.865 182.745 61.110 183.225 ;
        RECT 61.280 182.940 61.555 183.395 ;
        RECT 61.725 182.745 61.970 183.225 ;
        RECT 62.140 182.940 62.400 183.395 ;
        RECT 62.570 182.745 62.830 183.225 ;
        RECT 63.000 182.940 63.260 183.395 ;
        RECT 63.430 182.745 63.690 183.225 ;
        RECT 63.860 182.940 64.120 183.395 ;
        RECT 64.290 182.745 64.550 183.305 ;
        RECT 64.720 182.925 64.970 183.735 ;
        RECT 65.150 182.745 65.410 183.270 ;
        RECT 65.580 182.925 65.830 183.735 ;
        RECT 66.000 183.425 66.315 183.985 ;
        RECT 66.500 183.565 66.905 184.075 ;
        RECT 68.045 183.905 68.215 184.155 ;
        RECT 67.075 183.735 68.215 183.905 ;
        RECT 66.500 183.395 68.150 183.565 ;
        RECT 68.385 183.415 68.735 183.985 ;
        RECT 66.010 182.745 66.315 183.255 ;
        RECT 66.545 182.745 66.825 183.225 ;
        RECT 66.995 183.005 67.255 183.395 ;
        RECT 67.430 182.745 67.685 183.225 ;
        RECT 67.855 183.005 68.150 183.395 ;
        RECT 68.905 183.245 69.075 184.155 ;
        RECT 69.730 183.985 69.975 185.125 ;
        RECT 70.150 184.485 70.410 185.295 ;
        RECT 71.010 185.290 77.285 185.295 ;
        RECT 70.590 183.985 70.840 185.120 ;
        RECT 71.010 184.495 71.270 185.290 ;
        RECT 71.440 184.395 71.700 185.120 ;
        RECT 71.870 184.565 72.130 185.290 ;
        RECT 72.300 184.395 72.560 185.120 ;
        RECT 72.730 184.565 72.990 185.290 ;
        RECT 73.160 184.395 73.420 185.120 ;
        RECT 73.590 184.565 73.850 185.290 ;
        RECT 74.020 184.395 74.280 185.120 ;
        RECT 74.450 184.565 74.695 185.290 ;
        RECT 74.865 184.395 75.125 185.120 ;
        RECT 75.310 184.565 75.555 185.290 ;
        RECT 75.725 184.395 75.985 185.120 ;
        RECT 76.170 184.565 76.415 185.290 ;
        RECT 76.585 184.395 76.845 185.120 ;
        RECT 77.030 184.565 77.285 185.290 ;
        RECT 71.440 184.380 76.845 184.395 ;
        RECT 77.455 184.380 77.745 185.120 ;
        RECT 77.915 184.550 78.185 185.295 ;
        RECT 78.450 184.425 78.715 185.125 ;
        RECT 78.885 184.595 79.215 185.295 ;
        RECT 79.385 184.425 80.055 185.125 ;
        RECT 80.560 184.595 80.990 185.295 ;
        RECT 81.170 184.735 81.360 185.125 ;
        RECT 81.530 184.915 81.860 185.295 ;
        RECT 81.170 184.565 81.900 184.735 ;
        RECT 71.440 184.155 78.185 184.380 ;
        RECT 78.450 184.170 81.025 184.425 ;
        RECT 69.245 183.425 69.560 183.985 ;
        RECT 69.730 183.735 76.850 183.985 ;
        RECT 68.330 182.745 68.605 183.225 ;
        RECT 68.775 182.915 69.075 183.245 ;
        RECT 69.245 182.745 69.550 183.255 ;
        RECT 69.730 182.925 69.980 183.735 ;
        RECT 70.150 182.745 70.410 183.270 ;
        RECT 70.590 182.925 70.840 183.735 ;
        RECT 77.020 183.565 78.185 184.155 ;
        RECT 78.445 183.655 78.720 183.985 ;
        RECT 71.440 183.395 78.185 183.565 ;
        RECT 78.890 183.485 79.070 184.170 ;
        RECT 80.855 183.985 81.025 184.170 ;
        RECT 79.240 183.655 79.600 183.985 ;
        RECT 79.890 183.935 80.180 183.985 ;
        RECT 79.885 183.765 80.180 183.935 ;
        RECT 79.890 183.655 80.180 183.765 ;
        RECT 80.350 183.655 80.685 183.985 ;
        RECT 80.855 183.655 81.535 183.985 ;
        RECT 71.010 182.745 71.270 183.305 ;
        RECT 71.440 182.940 71.700 183.395 ;
        RECT 71.870 182.745 72.130 183.225 ;
        RECT 72.300 182.940 72.560 183.395 ;
        RECT 72.730 182.745 72.990 183.225 ;
        RECT 73.160 182.940 73.420 183.395 ;
        RECT 73.590 182.745 73.835 183.225 ;
        RECT 74.005 182.940 74.280 183.395 ;
        RECT 74.450 182.745 74.695 183.225 ;
        RECT 74.865 182.940 75.125 183.395 ;
        RECT 75.305 182.745 75.555 183.225 ;
        RECT 75.725 182.940 75.985 183.395 ;
        RECT 76.165 182.745 76.415 183.225 ;
        RECT 76.585 182.940 76.845 183.395 ;
        RECT 77.025 182.745 77.285 183.225 ;
        RECT 77.455 182.940 77.715 183.395 ;
        RECT 77.885 182.745 78.185 183.225 ;
        RECT 78.455 183.085 79.070 183.485 ;
        RECT 79.240 183.295 80.510 183.485 ;
        RECT 81.705 183.445 81.900 184.565 ;
        RECT 82.585 184.130 82.875 185.295 ;
        RECT 83.070 184.325 83.370 184.520 ;
        RECT 83.540 184.495 83.795 185.295 ;
        RECT 83.995 184.665 84.325 185.125 ;
        RECT 84.495 184.835 85.070 185.295 ;
        RECT 85.240 184.665 85.595 185.125 ;
        RECT 83.995 184.495 85.595 184.665 ;
        RECT 83.070 184.155 84.320 184.325 ;
        RECT 83.070 183.500 83.240 184.155 ;
        RECT 83.415 183.655 83.760 183.985 ;
        RECT 83.990 183.735 84.320 184.155 ;
        RECT 84.490 183.565 84.770 184.495 ;
        RECT 84.950 183.935 85.140 184.315 ;
        RECT 85.320 184.155 85.595 184.495 ;
        RECT 85.765 184.155 86.095 185.295 ;
        RECT 86.275 184.325 86.605 185.110 ;
        RECT 86.275 184.155 86.955 184.325 ;
        RECT 87.135 184.155 87.465 185.295 ;
        RECT 88.105 184.205 89.315 185.295 ;
        RECT 84.950 183.735 86.095 183.935 ;
        RECT 86.265 183.735 86.615 183.985 ;
        RECT 81.080 183.275 81.900 183.445 ;
        RECT 78.455 182.915 78.790 183.085 ;
        RECT 79.750 182.745 80.085 183.125 ;
        RECT 80.675 182.745 80.910 183.185 ;
        RECT 81.080 182.915 81.410 183.275 ;
        RECT 81.580 182.745 81.910 183.105 ;
        RECT 82.585 182.745 82.875 183.470 ;
        RECT 83.070 183.170 83.305 183.500 ;
        RECT 83.475 182.745 83.805 183.485 ;
        RECT 84.040 183.125 84.315 183.565 ;
        RECT 84.490 183.465 84.815 183.565 ;
        RECT 84.485 183.295 84.815 183.465 ;
        RECT 84.985 183.355 86.095 183.565 ;
        RECT 86.785 183.555 86.955 184.155 ;
        RECT 87.125 183.735 87.475 183.985 ;
        RECT 88.105 183.665 88.625 184.205 ;
        RECT 84.985 183.125 85.235 183.355 ;
        RECT 84.040 182.915 85.235 183.125 ;
        RECT 85.405 182.745 85.575 183.185 ;
        RECT 85.745 182.915 86.095 183.355 ;
        RECT 86.285 182.745 86.525 183.555 ;
        RECT 86.695 182.915 87.025 183.555 ;
        RECT 87.195 182.745 87.465 183.555 ;
        RECT 88.795 183.495 89.315 184.035 ;
        RECT 88.105 182.745 89.315 183.495 ;
        RECT 18.100 182.575 89.400 182.745 ;
        RECT 18.185 181.825 19.395 182.575 ;
        RECT 20.485 181.900 20.745 182.405 ;
        RECT 20.925 182.195 21.255 182.575 ;
        RECT 21.435 182.025 21.605 182.405 ;
        RECT 18.185 181.285 18.705 181.825 ;
        RECT 18.875 181.115 19.395 181.655 ;
        RECT 18.185 180.025 19.395 181.115 ;
        RECT 20.485 181.100 20.655 181.900 ;
        RECT 20.940 181.855 21.605 182.025 ;
        RECT 21.865 181.900 22.125 182.405 ;
        RECT 22.305 182.195 22.635 182.575 ;
        RECT 22.815 182.025 22.985 182.405 ;
        RECT 20.940 181.600 21.110 181.855 ;
        RECT 20.825 181.270 21.110 181.600 ;
        RECT 21.345 181.305 21.675 181.675 ;
        RECT 20.940 181.125 21.110 181.270 ;
        RECT 20.485 180.195 20.755 181.100 ;
        RECT 20.940 180.955 21.605 181.125 ;
        RECT 20.925 180.025 21.255 180.785 ;
        RECT 21.435 180.195 21.605 180.955 ;
        RECT 21.865 181.100 22.045 181.900 ;
        RECT 22.320 181.855 22.985 182.025 ;
        RECT 23.245 182.075 23.505 182.405 ;
        RECT 23.715 182.095 23.990 182.575 ;
        RECT 22.320 181.600 22.490 181.855 ;
        RECT 22.215 181.270 22.490 181.600 ;
        RECT 22.715 181.305 23.055 181.675 ;
        RECT 22.320 181.125 22.490 181.270 ;
        RECT 23.245 181.165 23.415 182.075 ;
        RECT 24.200 182.005 24.405 182.405 ;
        RECT 24.575 182.175 24.910 182.575 ;
        RECT 23.585 181.335 23.945 181.915 ;
        RECT 24.200 181.835 24.885 182.005 ;
        RECT 24.125 181.165 24.375 181.665 ;
        RECT 21.865 180.195 22.135 181.100 ;
        RECT 22.320 180.955 22.995 181.125 ;
        RECT 22.305 180.025 22.635 180.785 ;
        RECT 22.815 180.195 22.995 180.955 ;
        RECT 23.245 180.995 24.375 181.165 ;
        RECT 23.245 180.225 23.515 180.995 ;
        RECT 24.545 180.805 24.885 181.835 ;
        RECT 25.105 181.765 25.345 182.575 ;
        RECT 25.515 181.765 25.845 182.405 ;
        RECT 26.015 181.765 26.285 182.575 ;
        RECT 26.465 181.900 26.725 182.405 ;
        RECT 26.905 182.195 27.235 182.575 ;
        RECT 27.415 182.025 27.585 182.405 ;
        RECT 25.085 181.335 25.435 181.585 ;
        RECT 25.605 181.165 25.775 181.765 ;
        RECT 25.945 181.335 26.295 181.585 ;
        RECT 23.685 180.025 24.015 180.805 ;
        RECT 24.220 180.630 24.885 180.805 ;
        RECT 25.095 180.995 25.775 181.165 ;
        RECT 24.220 180.225 24.405 180.630 ;
        RECT 24.575 180.025 24.910 180.450 ;
        RECT 25.095 180.210 25.425 180.995 ;
        RECT 25.955 180.025 26.285 181.165 ;
        RECT 26.465 181.100 26.645 181.900 ;
        RECT 26.920 181.855 27.585 182.025 ;
        RECT 27.935 182.025 28.105 182.405 ;
        RECT 28.285 182.195 28.615 182.575 ;
        RECT 27.935 181.855 28.600 182.025 ;
        RECT 28.795 181.900 29.055 182.405 ;
        RECT 26.920 181.600 27.090 181.855 ;
        RECT 26.815 181.270 27.090 181.600 ;
        RECT 27.315 181.305 27.655 181.675 ;
        RECT 27.865 181.305 28.205 181.675 ;
        RECT 28.430 181.600 28.600 181.855 ;
        RECT 26.920 181.125 27.090 181.270 ;
        RECT 28.430 181.270 28.705 181.600 ;
        RECT 28.430 181.125 28.600 181.270 ;
        RECT 26.465 180.195 26.735 181.100 ;
        RECT 26.920 180.955 27.595 181.125 ;
        RECT 26.905 180.025 27.235 180.785 ;
        RECT 27.415 180.195 27.595 180.955 ;
        RECT 27.925 180.955 28.600 181.125 ;
        RECT 28.875 181.100 29.055 181.900 ;
        RECT 29.315 182.025 29.485 182.405 ;
        RECT 29.665 182.195 29.995 182.575 ;
        RECT 29.315 181.855 29.980 182.025 ;
        RECT 30.175 181.900 30.435 182.405 ;
        RECT 29.245 181.305 29.585 181.675 ;
        RECT 29.810 181.600 29.980 181.855 ;
        RECT 29.810 181.270 30.085 181.600 ;
        RECT 29.810 181.125 29.980 181.270 ;
        RECT 27.925 180.195 28.105 180.955 ;
        RECT 28.285 180.025 28.615 180.785 ;
        RECT 28.785 180.195 29.055 181.100 ;
        RECT 29.305 180.955 29.980 181.125 ;
        RECT 30.255 181.100 30.435 181.900 ;
        RECT 30.645 181.755 30.875 182.575 ;
        RECT 31.045 181.775 31.375 182.405 ;
        RECT 30.625 181.335 30.955 181.585 ;
        RECT 31.125 181.175 31.375 181.775 ;
        RECT 31.545 181.755 31.755 182.575 ;
        RECT 31.985 181.900 32.245 182.405 ;
        RECT 32.425 182.195 32.755 182.575 ;
        RECT 32.935 182.025 33.105 182.405 ;
        RECT 29.305 180.195 29.485 180.955 ;
        RECT 29.665 180.025 29.995 180.785 ;
        RECT 30.165 180.195 30.435 181.100 ;
        RECT 30.645 180.025 30.875 181.165 ;
        RECT 31.045 180.195 31.375 181.175 ;
        RECT 31.545 180.025 31.755 181.165 ;
        RECT 31.985 181.100 32.165 181.900 ;
        RECT 32.440 181.855 33.105 182.025 ;
        RECT 32.440 181.600 32.610 181.855 ;
        RECT 34.285 181.775 34.595 182.575 ;
        RECT 34.800 181.775 35.495 182.405 ;
        RECT 35.665 182.030 41.010 182.575 ;
        RECT 32.335 181.270 32.610 181.600 ;
        RECT 32.835 181.305 33.175 181.675 ;
        RECT 34.295 181.335 34.630 181.605 ;
        RECT 32.440 181.125 32.610 181.270 ;
        RECT 34.800 181.175 34.970 181.775 ;
        RECT 35.140 181.335 35.475 181.585 ;
        RECT 37.250 181.200 37.590 182.030 ;
        RECT 41.185 181.805 43.775 182.575 ;
        RECT 43.945 181.850 44.235 182.575 ;
        RECT 44.405 181.815 45.115 182.405 ;
        RECT 45.625 182.045 45.955 182.405 ;
        RECT 46.155 182.215 46.485 182.575 ;
        RECT 46.655 182.045 46.985 182.405 ;
        RECT 45.625 181.835 46.985 182.045 ;
        RECT 47.165 181.900 47.425 182.405 ;
        RECT 47.605 182.195 47.935 182.575 ;
        RECT 48.115 182.025 48.285 182.405 ;
        RECT 31.985 180.195 32.255 181.100 ;
        RECT 32.440 180.955 33.115 181.125 ;
        RECT 32.425 180.025 32.755 180.785 ;
        RECT 32.935 180.195 33.115 180.955 ;
        RECT 34.285 180.025 34.565 181.165 ;
        RECT 34.735 180.195 35.065 181.175 ;
        RECT 35.235 180.025 35.495 181.165 ;
        RECT 39.070 180.460 39.420 181.710 ;
        RECT 41.185 181.285 42.395 181.805 ;
        RECT 42.565 181.115 43.775 181.635 ;
        RECT 35.665 180.025 41.010 180.460 ;
        RECT 41.185 180.025 43.775 181.115 ;
        RECT 43.945 180.025 44.235 181.190 ;
        RECT 44.405 180.845 44.610 181.815 ;
        RECT 44.780 181.045 45.110 181.585 ;
        RECT 45.285 181.335 45.780 181.665 ;
        RECT 46.100 181.335 46.475 181.665 ;
        RECT 46.685 181.335 46.995 181.665 ;
        RECT 45.285 181.045 45.610 181.335 ;
        RECT 45.805 180.845 46.135 181.065 ;
        RECT 44.405 180.615 46.135 180.845 ;
        RECT 44.405 180.195 45.105 180.615 ;
        RECT 45.305 180.025 45.635 180.385 ;
        RECT 45.805 180.215 46.135 180.615 ;
        RECT 46.305 180.365 46.475 181.335 ;
        RECT 47.165 181.100 47.345 181.900 ;
        RECT 47.620 181.855 48.285 182.025 ;
        RECT 48.545 181.900 48.805 182.405 ;
        RECT 48.985 182.195 49.315 182.575 ;
        RECT 49.495 182.025 49.665 182.405 ;
        RECT 47.620 181.600 47.790 181.855 ;
        RECT 47.515 181.270 47.790 181.600 ;
        RECT 48.015 181.305 48.355 181.675 ;
        RECT 47.620 181.125 47.790 181.270 ;
        RECT 46.655 180.025 46.985 181.085 ;
        RECT 47.165 180.195 47.435 181.100 ;
        RECT 47.620 180.955 48.295 181.125 ;
        RECT 47.605 180.025 47.935 180.785 ;
        RECT 48.115 180.195 48.295 180.955 ;
        RECT 48.545 181.100 48.725 181.900 ;
        RECT 49.000 181.855 49.665 182.025 ;
        RECT 50.015 182.025 50.185 182.405 ;
        RECT 50.365 182.195 50.695 182.575 ;
        RECT 50.015 181.855 50.680 182.025 ;
        RECT 50.875 181.900 51.135 182.405 ;
        RECT 49.000 181.600 49.170 181.855 ;
        RECT 48.895 181.270 49.170 181.600 ;
        RECT 49.395 181.305 49.735 181.675 ;
        RECT 49.945 181.305 50.285 181.675 ;
        RECT 50.510 181.600 50.680 181.855 ;
        RECT 49.000 181.125 49.170 181.270 ;
        RECT 50.510 181.270 50.785 181.600 ;
        RECT 50.510 181.125 50.680 181.270 ;
        RECT 48.545 180.195 48.815 181.100 ;
        RECT 49.000 180.955 49.675 181.125 ;
        RECT 48.985 180.025 49.315 180.785 ;
        RECT 49.495 180.195 49.675 180.955 ;
        RECT 50.005 180.955 50.680 181.125 ;
        RECT 50.955 181.100 51.135 181.900 ;
        RECT 50.005 180.195 50.185 180.955 ;
        RECT 50.365 180.025 50.695 180.785 ;
        RECT 50.865 180.195 51.135 181.100 ;
        RECT 51.305 181.900 51.565 182.405 ;
        RECT 51.745 182.195 52.075 182.575 ;
        RECT 52.255 182.025 52.425 182.405 ;
        RECT 51.305 181.100 51.485 181.900 ;
        RECT 51.760 181.855 52.425 182.025 ;
        RECT 52.685 181.900 52.945 182.405 ;
        RECT 53.125 182.195 53.455 182.575 ;
        RECT 53.635 182.025 53.805 182.405 ;
        RECT 51.760 181.600 51.930 181.855 ;
        RECT 51.655 181.270 51.930 181.600 ;
        RECT 52.155 181.305 52.495 181.675 ;
        RECT 51.760 181.125 51.930 181.270 ;
        RECT 51.305 180.195 51.575 181.100 ;
        RECT 51.760 180.955 52.435 181.125 ;
        RECT 51.745 180.025 52.075 180.785 ;
        RECT 52.255 180.195 52.435 180.955 ;
        RECT 52.685 181.100 52.865 181.900 ;
        RECT 53.140 181.855 53.805 182.025 ;
        RECT 53.140 181.600 53.310 181.855 ;
        RECT 54.070 181.810 54.525 182.575 ;
        RECT 54.800 182.195 56.100 182.405 ;
        RECT 56.355 182.215 56.685 182.575 ;
        RECT 55.930 182.045 56.100 182.195 ;
        RECT 56.855 182.075 57.115 182.405 ;
        RECT 53.035 181.270 53.310 181.600 ;
        RECT 53.535 181.305 53.875 181.675 ;
        RECT 55.000 181.585 55.220 181.985 ;
        RECT 54.065 181.385 54.555 181.585 ;
        RECT 54.745 181.375 55.220 181.585 ;
        RECT 55.465 181.585 55.675 181.985 ;
        RECT 55.930 181.920 56.685 182.045 ;
        RECT 55.930 181.875 56.775 181.920 ;
        RECT 56.505 181.755 56.775 181.875 ;
        RECT 55.465 181.375 55.795 181.585 ;
        RECT 55.965 181.315 56.375 181.620 ;
        RECT 53.140 181.125 53.310 181.270 ;
        RECT 54.070 181.145 55.245 181.205 ;
        RECT 56.605 181.180 56.775 181.755 ;
        RECT 56.575 181.145 56.775 181.180 ;
        RECT 52.685 180.195 52.955 181.100 ;
        RECT 53.140 180.955 53.815 181.125 ;
        RECT 53.125 180.025 53.455 180.785 ;
        RECT 53.635 180.195 53.815 180.955 ;
        RECT 54.070 181.035 56.775 181.145 ;
        RECT 54.070 180.415 54.325 181.035 ;
        RECT 54.915 180.975 56.715 181.035 ;
        RECT 54.915 180.945 55.245 180.975 ;
        RECT 56.945 180.875 57.115 182.075 ;
        RECT 54.575 180.775 54.760 180.865 ;
        RECT 55.350 180.775 56.185 180.785 ;
        RECT 54.575 180.575 56.185 180.775 ;
        RECT 54.575 180.535 54.805 180.575 ;
        RECT 54.070 180.195 54.405 180.415 ;
        RECT 55.410 180.025 55.765 180.405 ;
        RECT 55.935 180.195 56.185 180.575 ;
        RECT 56.435 180.025 56.685 180.805 ;
        RECT 56.855 180.195 57.115 180.875 ;
        RECT 57.285 181.755 57.970 182.395 ;
        RECT 58.140 181.755 58.310 182.575 ;
        RECT 58.480 181.925 58.810 182.390 ;
        RECT 58.980 182.105 59.150 182.575 ;
        RECT 59.410 182.185 60.595 182.355 ;
        RECT 60.765 182.015 61.095 182.405 ;
        RECT 59.795 181.925 60.180 182.015 ;
        RECT 58.480 181.755 60.180 181.925 ;
        RECT 60.585 181.835 61.095 182.015 ;
        RECT 61.425 182.075 61.685 182.405 ;
        RECT 61.855 182.215 62.185 182.575 ;
        RECT 62.440 182.195 63.740 182.405 ;
        RECT 57.285 180.785 57.535 181.755 ;
        RECT 57.705 181.375 58.040 181.585 ;
        RECT 58.210 181.375 58.660 181.585 ;
        RECT 58.850 181.375 59.335 181.585 ;
        RECT 57.870 181.205 58.040 181.375 ;
        RECT 58.960 181.215 59.335 181.375 ;
        RECT 59.525 181.335 59.905 181.585 ;
        RECT 60.085 181.375 60.415 181.585 ;
        RECT 57.870 181.035 58.790 181.205 ;
        RECT 57.285 180.195 57.950 180.785 ;
        RECT 58.120 180.025 58.450 180.865 ;
        RECT 58.620 180.785 58.790 181.035 ;
        RECT 58.960 181.045 59.355 181.215 ;
        RECT 58.960 180.955 59.335 181.045 ;
        RECT 59.525 180.955 59.845 181.335 ;
        RECT 60.585 181.205 60.755 181.835 ;
        RECT 60.925 181.375 61.255 181.665 ;
        RECT 60.015 181.035 61.100 181.205 ;
        RECT 60.015 180.785 60.185 181.035 ;
        RECT 58.620 180.615 60.185 180.785 ;
        RECT 58.960 180.195 59.765 180.615 ;
        RECT 60.355 180.025 60.605 180.865 ;
        RECT 60.800 180.195 61.100 181.035 ;
        RECT 61.425 180.875 61.595 182.075 ;
        RECT 62.440 182.045 62.610 182.195 ;
        RECT 61.855 181.920 62.610 182.045 ;
        RECT 61.765 181.875 62.610 181.920 ;
        RECT 61.765 181.755 62.035 181.875 ;
        RECT 61.765 181.180 61.935 181.755 ;
        RECT 62.165 181.315 62.575 181.620 ;
        RECT 62.865 181.585 63.075 181.985 ;
        RECT 62.745 181.375 63.075 181.585 ;
        RECT 63.320 181.585 63.540 181.985 ;
        RECT 64.015 181.810 64.470 182.575 ;
        RECT 63.320 181.375 63.795 181.585 ;
        RECT 63.985 181.385 64.475 181.585 ;
        RECT 61.765 181.145 61.965 181.180 ;
        RECT 63.295 181.145 64.470 181.205 ;
        RECT 61.765 181.035 64.470 181.145 ;
        RECT 61.825 180.975 63.625 181.035 ;
        RECT 63.295 180.945 63.625 180.975 ;
        RECT 61.425 180.195 61.685 180.875 ;
        RECT 61.855 180.025 62.105 180.805 ;
        RECT 62.355 180.775 63.190 180.785 ;
        RECT 63.780 180.775 63.965 180.865 ;
        RECT 62.355 180.575 63.965 180.775 ;
        RECT 62.355 180.195 62.605 180.575 ;
        RECT 63.735 180.535 63.965 180.575 ;
        RECT 64.215 180.415 64.470 181.035 ;
        RECT 62.775 180.025 63.130 180.405 ;
        RECT 64.135 180.195 64.470 180.415 ;
        RECT 65.580 180.205 65.860 182.395 ;
        RECT 66.060 182.205 66.790 182.575 ;
        RECT 67.370 182.035 67.800 182.395 ;
        RECT 66.060 181.845 67.800 182.035 ;
        RECT 66.060 181.335 66.320 181.845 ;
        RECT 66.050 180.025 66.335 181.165 ;
        RECT 66.530 181.045 66.790 181.665 ;
        RECT 66.985 181.045 67.410 181.665 ;
        RECT 67.580 181.615 67.800 181.845 ;
        RECT 67.970 181.795 68.215 182.575 ;
        RECT 67.580 181.315 68.125 181.615 ;
        RECT 68.415 181.495 68.645 182.395 ;
        RECT 66.600 180.675 67.625 180.875 ;
        RECT 66.600 180.205 66.770 180.675 ;
        RECT 66.945 180.025 67.275 180.505 ;
        RECT 67.445 180.205 67.625 180.675 ;
        RECT 67.795 180.205 68.125 181.315 ;
        RECT 68.305 180.815 68.645 181.495 ;
        RECT 68.825 180.995 69.055 182.335 ;
        RECT 69.705 181.850 69.995 182.575 ;
        RECT 70.615 182.095 70.785 182.575 ;
        RECT 70.955 181.925 71.285 182.400 ;
        RECT 71.455 182.095 71.625 182.575 ;
        RECT 71.795 181.925 72.125 182.400 ;
        RECT 72.295 182.095 72.465 182.575 ;
        RECT 72.635 181.925 72.965 182.400 ;
        RECT 73.135 182.095 73.305 182.575 ;
        RECT 73.475 181.925 73.805 182.400 ;
        RECT 73.975 182.095 74.145 182.575 ;
        RECT 74.315 181.925 74.645 182.400 ;
        RECT 74.815 182.095 74.985 182.575 ;
        RECT 75.155 181.925 75.485 182.400 ;
        RECT 70.165 181.755 73.805 181.925 ;
        RECT 73.975 181.755 75.485 181.925 ;
        RECT 75.675 181.755 76.005 182.400 ;
        RECT 76.175 181.755 76.345 182.575 ;
        RECT 76.610 181.925 76.880 182.135 ;
        RECT 77.100 182.115 77.430 182.575 ;
        RECT 77.940 182.115 78.690 182.405 ;
        RECT 76.610 181.755 77.945 181.925 ;
        RECT 70.165 181.215 70.550 181.755 ;
        RECT 73.975 181.585 74.145 181.755 ;
        RECT 75.675 181.585 75.845 181.755 ;
        RECT 77.775 181.585 77.945 181.755 ;
        RECT 70.760 181.385 74.145 181.585 ;
        RECT 74.315 181.385 75.845 181.585 ;
        RECT 76.015 181.385 76.435 181.585 ;
        RECT 73.975 181.215 74.145 181.385 ;
        RECT 68.305 180.615 69.055 180.815 ;
        RECT 68.295 180.025 68.645 180.435 ;
        RECT 68.815 180.225 69.055 180.615 ;
        RECT 69.705 180.025 69.995 181.190 ;
        RECT 70.165 181.045 73.805 181.215 ;
        RECT 73.975 181.045 75.485 181.215 ;
        RECT 70.615 180.025 70.785 180.825 ;
        RECT 70.955 180.195 71.285 181.045 ;
        RECT 71.455 180.025 71.625 180.825 ;
        RECT 71.795 180.195 72.125 181.045 ;
        RECT 72.295 180.025 72.465 180.825 ;
        RECT 72.635 180.195 72.965 181.045 ;
        RECT 73.135 180.025 73.305 180.825 ;
        RECT 73.475 180.195 73.805 181.045 ;
        RECT 73.975 180.025 74.145 180.875 ;
        RECT 74.315 180.195 74.645 181.045 ;
        RECT 74.815 180.025 74.985 180.875 ;
        RECT 75.155 180.195 75.485 181.045 ;
        RECT 75.675 181.115 75.845 181.385 ;
        RECT 76.610 181.345 76.960 181.585 ;
        RECT 77.130 181.345 77.605 181.585 ;
        RECT 77.775 181.335 78.150 181.585 ;
        RECT 75.675 180.195 76.005 181.115 ;
        RECT 76.175 180.025 76.345 181.215 ;
        RECT 77.775 181.165 77.945 181.335 ;
        RECT 76.610 180.995 77.945 181.165 ;
        RECT 76.610 180.835 76.890 180.995 ;
        RECT 78.320 180.825 78.690 182.115 ;
        RECT 78.995 182.095 79.295 182.575 ;
        RECT 79.465 181.925 79.725 182.380 ;
        RECT 79.895 182.095 80.155 182.575 ;
        RECT 80.335 181.925 80.595 182.380 ;
        RECT 80.765 182.095 81.015 182.575 ;
        RECT 81.195 181.925 81.455 182.380 ;
        RECT 81.625 182.095 81.875 182.575 ;
        RECT 82.055 181.925 82.315 182.380 ;
        RECT 82.485 182.095 82.730 182.575 ;
        RECT 82.900 181.925 83.175 182.380 ;
        RECT 83.345 182.095 83.590 182.575 ;
        RECT 83.760 181.925 84.020 182.380 ;
        RECT 84.190 182.095 84.450 182.575 ;
        RECT 84.620 181.925 84.880 182.380 ;
        RECT 85.050 182.095 85.310 182.575 ;
        RECT 85.480 181.925 85.740 182.380 ;
        RECT 85.910 182.015 86.170 182.575 ;
        RECT 78.995 181.755 85.740 181.925 ;
        RECT 78.995 181.165 80.160 181.755 ;
        RECT 86.340 181.585 86.590 182.395 ;
        RECT 86.770 182.050 87.030 182.575 ;
        RECT 87.200 181.585 87.450 182.395 ;
        RECT 87.630 182.065 87.935 182.575 ;
        RECT 80.330 181.335 87.450 181.585 ;
        RECT 87.620 181.335 87.935 181.895 ;
        RECT 88.105 181.825 89.315 182.575 ;
        RECT 78.995 180.940 85.740 181.165 ;
        RECT 77.100 180.025 77.350 180.825 ;
        RECT 77.520 180.655 78.690 180.825 ;
        RECT 77.520 180.195 77.850 180.655 ;
        RECT 78.020 180.025 78.235 180.485 ;
        RECT 78.995 180.025 79.265 180.770 ;
        RECT 79.435 180.200 79.725 180.940 ;
        RECT 80.335 180.925 85.740 180.940 ;
        RECT 79.895 180.030 80.150 180.755 ;
        RECT 80.335 180.200 80.595 180.925 ;
        RECT 80.765 180.030 81.010 180.755 ;
        RECT 81.195 180.200 81.455 180.925 ;
        RECT 81.625 180.030 81.870 180.755 ;
        RECT 82.055 180.200 82.315 180.925 ;
        RECT 82.485 180.030 82.730 180.755 ;
        RECT 82.900 180.200 83.160 180.925 ;
        RECT 83.330 180.030 83.590 180.755 ;
        RECT 83.760 180.200 84.020 180.925 ;
        RECT 84.190 180.030 84.450 180.755 ;
        RECT 84.620 180.200 84.880 180.925 ;
        RECT 85.050 180.030 85.310 180.755 ;
        RECT 85.480 180.200 85.740 180.925 ;
        RECT 85.910 180.030 86.170 180.825 ;
        RECT 86.340 180.200 86.590 181.335 ;
        RECT 79.895 180.025 86.170 180.030 ;
        RECT 86.770 180.025 87.030 180.835 ;
        RECT 87.205 180.195 87.450 181.335 ;
        RECT 88.105 181.115 88.625 181.655 ;
        RECT 88.795 181.285 89.315 181.825 ;
        RECT 87.630 180.025 87.925 180.835 ;
        RECT 88.105 180.025 89.315 181.115 ;
        RECT 18.100 179.855 89.400 180.025 ;
        RECT 18.185 178.765 19.395 179.855 ;
        RECT 18.185 178.055 18.705 178.595 ;
        RECT 18.875 178.225 19.395 178.765 ;
        RECT 20.670 178.885 21.060 179.060 ;
        RECT 21.545 179.055 21.875 179.855 ;
        RECT 22.045 179.065 22.580 179.685 ;
        RECT 20.670 178.715 22.095 178.885 ;
        RECT 18.185 177.305 19.395 178.055 ;
        RECT 20.545 177.985 20.900 178.545 ;
        RECT 21.070 177.815 21.240 178.715 ;
        RECT 21.410 177.985 21.675 178.545 ;
        RECT 21.925 178.215 22.095 178.715 ;
        RECT 22.265 178.045 22.580 179.065 ;
        RECT 22.785 178.900 23.055 179.855 ;
        RECT 20.650 177.305 20.890 177.815 ;
        RECT 21.070 177.485 21.350 177.815 ;
        RECT 21.580 177.305 21.795 177.815 ;
        RECT 21.965 177.475 22.580 178.045 ;
        RECT 23.240 178.800 23.545 179.585 ;
        RECT 23.725 179.385 24.410 179.855 ;
        RECT 23.720 178.865 24.415 179.175 ;
        RECT 23.240 177.995 23.415 178.800 ;
        RECT 24.590 178.695 24.875 179.640 ;
        RECT 25.075 179.405 25.405 179.855 ;
        RECT 25.575 179.235 25.745 179.665 ;
        RECT 24.015 178.545 24.875 178.695 ;
        RECT 23.585 178.525 24.875 178.545 ;
        RECT 25.065 179.005 25.745 179.235 ;
        RECT 26.095 179.235 26.265 179.665 ;
        RECT 26.435 179.405 26.765 179.855 ;
        RECT 26.095 179.005 26.770 179.235 ;
        RECT 23.585 178.165 24.575 178.525 ;
        RECT 25.065 178.355 25.300 179.005 ;
        RECT 22.785 177.305 23.055 177.940 ;
        RECT 23.240 177.475 23.475 177.995 ;
        RECT 24.405 177.830 24.575 178.165 ;
        RECT 24.745 178.025 25.300 178.355 ;
        RECT 25.085 177.875 25.300 178.025 ;
        RECT 25.470 178.665 25.775 178.835 ;
        RECT 25.470 177.985 25.770 178.665 ;
        RECT 26.065 177.985 26.365 178.835 ;
        RECT 26.535 178.355 26.770 179.005 ;
        RECT 26.940 178.695 27.225 179.640 ;
        RECT 27.405 179.385 28.090 179.855 ;
        RECT 27.400 178.865 28.095 179.175 ;
        RECT 28.270 178.800 28.575 179.585 ;
        RECT 26.940 178.545 27.800 178.695 ;
        RECT 26.940 178.525 28.225 178.545 ;
        RECT 26.535 178.025 27.070 178.355 ;
        RECT 27.240 178.165 28.225 178.525 ;
        RECT 26.535 177.875 26.755 178.025 ;
        RECT 23.645 177.305 24.045 177.800 ;
        RECT 24.405 177.635 24.805 177.830 ;
        RECT 24.635 177.490 24.805 177.635 ;
        RECT 25.085 177.500 25.325 177.875 ;
        RECT 25.495 177.305 25.825 177.810 ;
        RECT 26.010 177.305 26.345 177.810 ;
        RECT 26.515 177.500 26.755 177.875 ;
        RECT 27.240 177.830 27.410 178.165 ;
        RECT 28.400 177.995 28.575 178.800 ;
        RECT 29.235 179.245 29.565 179.675 ;
        RECT 29.745 179.415 29.940 179.855 ;
        RECT 30.110 179.245 30.440 179.675 ;
        RECT 29.235 179.075 30.440 179.245 ;
        RECT 29.235 178.745 30.130 179.075 ;
        RECT 30.610 178.905 30.885 179.675 ;
        RECT 30.300 178.715 30.885 178.905 ;
        RECT 29.240 178.215 29.535 178.545 ;
        RECT 29.715 178.215 30.130 178.545 ;
        RECT 27.035 177.635 27.410 177.830 ;
        RECT 27.035 177.490 27.205 177.635 ;
        RECT 27.770 177.305 28.165 177.800 ;
        RECT 28.335 177.475 28.575 177.995 ;
        RECT 29.235 177.305 29.535 178.035 ;
        RECT 29.715 177.595 29.945 178.215 ;
        RECT 30.300 178.045 30.475 178.715 ;
        RECT 31.065 178.690 31.355 179.855 ;
        RECT 32.455 178.795 32.785 179.645 ;
        RECT 32.455 178.665 32.675 178.795 ;
        RECT 32.955 178.715 33.205 179.855 ;
        RECT 33.395 179.215 33.645 179.635 ;
        RECT 33.875 179.385 34.205 179.855 ;
        RECT 34.435 179.215 34.685 179.635 ;
        RECT 33.395 179.045 34.685 179.215 ;
        RECT 34.865 179.215 35.195 179.645 ;
        RECT 34.865 179.045 35.320 179.215 ;
        RECT 30.145 177.865 30.475 178.045 ;
        RECT 30.645 177.895 30.885 178.545 ;
        RECT 32.455 178.030 32.645 178.665 ;
        RECT 33.385 178.545 33.600 178.875 ;
        RECT 32.815 178.215 33.125 178.545 ;
        RECT 33.295 178.215 33.600 178.545 ;
        RECT 33.775 178.215 34.060 178.875 ;
        RECT 34.255 178.215 34.520 178.875 ;
        RECT 34.735 178.215 34.980 178.875 ;
        RECT 32.955 178.045 33.125 178.215 ;
        RECT 35.150 178.045 35.320 179.045 ;
        RECT 35.670 178.715 35.990 179.855 ;
        RECT 36.170 178.545 36.365 179.595 ;
        RECT 36.545 179.005 36.875 179.685 ;
        RECT 37.075 179.055 37.330 179.855 ;
        RECT 37.525 179.015 37.780 179.685 ;
        RECT 37.950 179.095 38.280 179.855 ;
        RECT 38.450 179.255 38.700 179.685 ;
        RECT 38.870 179.435 39.225 179.855 ;
        RECT 39.415 179.515 40.585 179.685 ;
        RECT 39.415 179.475 39.745 179.515 ;
        RECT 39.855 179.255 40.085 179.345 ;
        RECT 38.450 179.015 40.085 179.255 ;
        RECT 40.255 179.015 40.585 179.515 ;
        RECT 37.525 179.005 37.735 179.015 ;
        RECT 36.545 178.725 36.895 179.005 ;
        RECT 35.730 178.495 35.990 178.545 ;
        RECT 35.725 178.325 35.990 178.495 ;
        RECT 35.730 178.215 35.990 178.325 ;
        RECT 36.170 178.215 36.555 178.545 ;
        RECT 36.725 178.345 36.895 178.725 ;
        RECT 37.085 178.515 37.330 178.875 ;
        RECT 36.725 178.175 37.245 178.345 ;
        RECT 30.145 177.485 30.370 177.865 ;
        RECT 30.540 177.305 30.870 177.695 ;
        RECT 31.065 177.305 31.355 178.030 ;
        RECT 32.455 177.520 32.785 178.030 ;
        RECT 32.955 177.875 35.320 178.045 ;
        RECT 32.955 177.305 33.285 177.705 ;
        RECT 34.335 177.535 34.665 177.875 ;
        RECT 35.670 177.835 36.885 178.005 ;
        RECT 34.835 177.305 35.165 177.705 ;
        RECT 35.670 177.485 35.960 177.835 ;
        RECT 36.155 177.305 36.485 177.665 ;
        RECT 36.655 177.530 36.885 177.835 ;
        RECT 37.075 177.610 37.245 178.175 ;
        RECT 37.525 177.885 37.695 179.005 ;
        RECT 40.755 178.845 40.925 179.685 ;
        RECT 37.865 178.675 40.925 178.845 ;
        RECT 41.190 179.135 41.525 179.645 ;
        RECT 37.865 178.125 38.035 178.675 ;
        RECT 38.265 178.295 38.630 178.495 ;
        RECT 38.800 178.295 39.130 178.495 ;
        RECT 37.865 177.955 38.665 178.125 ;
        RECT 37.525 177.805 37.710 177.885 ;
        RECT 37.525 177.475 37.780 177.805 ;
        RECT 37.995 177.305 38.325 177.785 ;
        RECT 38.495 177.725 38.665 177.955 ;
        RECT 38.845 177.895 39.130 178.295 ;
        RECT 39.400 178.295 39.875 178.495 ;
        RECT 40.045 178.295 40.490 178.495 ;
        RECT 40.660 178.295 41.010 178.505 ;
        RECT 39.400 177.895 39.680 178.295 ;
        RECT 39.860 177.955 40.925 178.125 ;
        RECT 39.860 177.725 40.030 177.955 ;
        RECT 38.495 177.475 40.030 177.725 ;
        RECT 40.255 177.305 40.585 177.785 ;
        RECT 40.755 177.475 40.925 177.955 ;
        RECT 41.190 177.780 41.445 179.135 ;
        RECT 41.775 179.055 42.105 179.855 ;
        RECT 42.350 179.265 42.635 179.685 ;
        RECT 42.890 179.435 43.220 179.855 ;
        RECT 43.445 179.515 44.605 179.685 ;
        RECT 43.445 179.265 43.775 179.515 ;
        RECT 42.350 179.095 43.775 179.265 ;
        RECT 44.005 178.885 44.175 179.345 ;
        RECT 44.435 179.015 44.605 179.515 ;
        RECT 41.805 178.715 44.175 178.885 ;
        RECT 41.805 178.545 41.975 178.715 ;
        RECT 44.425 178.665 44.635 178.835 ;
        RECT 44.865 178.745 45.125 179.685 ;
        RECT 45.295 179.455 45.625 179.855 ;
        RECT 46.770 179.590 47.025 179.685 ;
        RECT 45.885 179.420 47.025 179.590 ;
        RECT 47.195 179.475 47.525 179.645 ;
        RECT 45.885 179.195 46.055 179.420 ;
        RECT 45.295 179.025 46.055 179.195 ;
        RECT 46.770 179.285 47.025 179.420 ;
        RECT 44.425 178.545 44.630 178.665 ;
        RECT 41.670 178.215 41.975 178.545 ;
        RECT 42.170 178.495 42.420 178.545 ;
        RECT 42.165 178.325 42.420 178.495 ;
        RECT 42.170 178.215 42.420 178.325 ;
        RECT 41.805 178.045 41.975 178.215 ;
        RECT 42.630 178.155 42.900 178.545 ;
        RECT 43.090 178.495 43.380 178.545 ;
        RECT 43.085 178.325 43.380 178.495 ;
        RECT 41.805 177.875 42.365 178.045 ;
        RECT 42.625 177.985 42.900 178.155 ;
        RECT 42.630 177.885 42.900 177.985 ;
        RECT 43.090 177.885 43.380 178.325 ;
        RECT 43.550 177.880 43.970 178.545 ;
        RECT 44.280 178.215 44.630 178.545 ;
        RECT 44.865 178.030 45.040 178.745 ;
        RECT 45.295 178.545 45.465 179.025 ;
        RECT 46.320 178.935 46.490 179.125 ;
        RECT 46.770 179.115 47.180 179.285 ;
        RECT 45.210 178.215 45.465 178.545 ;
        RECT 45.690 178.215 46.020 178.835 ;
        RECT 46.320 178.765 46.840 178.935 ;
        RECT 46.190 178.215 46.480 178.595 ;
        RECT 46.670 178.045 46.840 178.765 ;
        RECT 41.190 177.520 41.525 177.780 ;
        RECT 42.195 177.705 42.365 177.875 ;
        RECT 41.695 177.305 42.025 177.705 ;
        RECT 42.195 177.535 43.810 177.705 ;
        RECT 44.355 177.305 44.685 178.025 ;
        RECT 44.865 177.475 45.125 178.030 ;
        RECT 45.960 177.875 46.840 178.045 ;
        RECT 47.010 178.090 47.180 179.115 ;
        RECT 47.355 179.225 47.525 179.475 ;
        RECT 47.695 179.395 47.945 179.855 ;
        RECT 48.115 179.225 48.295 179.685 ;
        RECT 47.355 179.055 48.295 179.225 ;
        RECT 49.010 179.055 49.265 179.855 ;
        RECT 49.465 179.005 49.795 179.685 ;
        RECT 47.380 178.575 47.860 178.875 ;
        RECT 47.010 177.920 47.360 178.090 ;
        RECT 47.600 177.985 47.860 178.575 ;
        RECT 48.060 177.985 48.320 178.875 ;
        RECT 49.010 178.515 49.255 178.875 ;
        RECT 49.445 178.725 49.795 179.005 ;
        RECT 49.445 178.345 49.615 178.725 ;
        RECT 49.975 178.545 50.170 179.595 ;
        RECT 50.350 178.715 50.670 179.855 ;
        RECT 50.865 178.800 51.170 179.585 ;
        RECT 51.350 179.385 52.035 179.855 ;
        RECT 51.345 178.865 52.040 179.175 ;
        RECT 49.095 178.175 49.615 178.345 ;
        RECT 49.785 178.215 50.170 178.545 ;
        RECT 50.350 178.495 50.610 178.545 ;
        RECT 50.350 178.325 50.615 178.495 ;
        RECT 50.350 178.215 50.610 178.325 ;
        RECT 49.095 178.155 49.265 178.175 ;
        RECT 49.065 177.985 49.265 178.155 ;
        RECT 45.295 177.305 45.725 177.750 ;
        RECT 45.960 177.475 46.130 177.875 ;
        RECT 46.300 177.305 47.020 177.705 ;
        RECT 47.190 177.475 47.360 177.920 ;
        RECT 47.935 177.305 48.335 177.815 ;
        RECT 49.095 177.610 49.265 177.985 ;
        RECT 49.455 177.835 50.670 178.005 ;
        RECT 49.455 177.530 49.685 177.835 ;
        RECT 49.855 177.305 50.185 177.665 ;
        RECT 50.380 177.485 50.670 177.835 ;
        RECT 50.865 177.995 51.040 178.800 ;
        RECT 52.215 178.695 52.500 179.640 ;
        RECT 52.675 179.405 53.005 179.855 ;
        RECT 53.175 179.235 53.345 179.665 ;
        RECT 51.640 178.545 52.500 178.695 ;
        RECT 51.215 178.525 52.500 178.545 ;
        RECT 52.670 179.005 53.345 179.235 ;
        RECT 53.695 179.235 53.865 179.665 ;
        RECT 54.035 179.405 54.365 179.855 ;
        RECT 53.695 179.005 54.370 179.235 ;
        RECT 51.215 178.165 52.200 178.525 ;
        RECT 52.670 178.355 52.905 179.005 ;
        RECT 50.865 177.475 51.105 177.995 ;
        RECT 52.030 177.830 52.200 178.165 ;
        RECT 52.370 178.025 52.905 178.355 ;
        RECT 52.685 177.875 52.905 178.025 ;
        RECT 53.075 177.985 53.375 178.835 ;
        RECT 53.665 177.985 53.965 178.835 ;
        RECT 54.135 178.355 54.370 179.005 ;
        RECT 54.540 178.695 54.825 179.640 ;
        RECT 55.005 179.385 55.690 179.855 ;
        RECT 55.000 178.865 55.695 179.175 ;
        RECT 55.870 178.800 56.175 179.585 ;
        RECT 54.540 178.545 55.400 178.695 ;
        RECT 54.540 178.525 55.825 178.545 ;
        RECT 54.135 178.025 54.670 178.355 ;
        RECT 54.840 178.165 55.825 178.525 ;
        RECT 54.135 177.875 54.355 178.025 ;
        RECT 51.275 177.305 51.670 177.800 ;
        RECT 52.030 177.635 52.405 177.830 ;
        RECT 52.235 177.490 52.405 177.635 ;
        RECT 52.685 177.500 52.925 177.875 ;
        RECT 53.095 177.305 53.430 177.810 ;
        RECT 53.610 177.305 53.945 177.810 ;
        RECT 54.115 177.500 54.355 177.875 ;
        RECT 54.840 177.830 55.010 178.165 ;
        RECT 56.000 177.995 56.175 178.800 ;
        RECT 56.825 178.690 57.115 179.855 ;
        RECT 57.290 179.465 57.625 179.685 ;
        RECT 58.630 179.475 58.985 179.855 ;
        RECT 57.290 178.845 57.545 179.465 ;
        RECT 57.795 179.305 58.025 179.345 ;
        RECT 59.155 179.305 59.405 179.685 ;
        RECT 57.795 179.105 59.405 179.305 ;
        RECT 57.795 179.015 57.980 179.105 ;
        RECT 58.570 179.095 59.405 179.105 ;
        RECT 59.655 179.075 59.905 179.855 ;
        RECT 60.075 179.005 60.335 179.685 ;
        RECT 58.135 178.905 58.465 178.935 ;
        RECT 58.135 178.845 59.935 178.905 ;
        RECT 57.290 178.735 59.995 178.845 ;
        RECT 57.290 178.675 58.465 178.735 ;
        RECT 59.795 178.700 59.995 178.735 ;
        RECT 57.285 178.295 57.775 178.495 ;
        RECT 57.965 178.295 58.440 178.505 ;
        RECT 54.635 177.635 55.010 177.830 ;
        RECT 54.635 177.490 54.805 177.635 ;
        RECT 55.370 177.305 55.765 177.800 ;
        RECT 55.935 177.475 56.175 177.995 ;
        RECT 56.825 177.305 57.115 178.030 ;
        RECT 57.290 177.305 57.745 178.070 ;
        RECT 58.220 177.895 58.440 178.295 ;
        RECT 58.685 178.295 59.015 178.505 ;
        RECT 58.685 177.895 58.895 178.295 ;
        RECT 59.185 178.260 59.595 178.565 ;
        RECT 59.825 178.125 59.995 178.700 ;
        RECT 59.725 178.005 59.995 178.125 ;
        RECT 59.150 177.960 59.995 178.005 ;
        RECT 59.150 177.835 59.905 177.960 ;
        RECT 59.150 177.685 59.320 177.835 ;
        RECT 60.165 177.805 60.335 179.005 ;
        RECT 61.435 179.515 62.605 179.685 ;
        RECT 61.435 178.845 61.765 179.515 ;
        RECT 62.275 179.475 62.605 179.515 ;
        RECT 62.775 179.475 63.150 179.855 ;
        RECT 61.935 179.305 62.165 179.345 ;
        RECT 61.935 179.255 62.550 179.305 ;
        RECT 63.295 179.255 63.465 179.385 ;
        RECT 61.935 179.055 63.465 179.255 ;
        RECT 63.700 179.075 63.965 179.855 ;
        RECT 61.935 179.015 62.815 179.055 ;
        RECT 64.275 178.925 64.445 179.685 ;
        RECT 64.660 179.095 64.990 179.855 ;
        RECT 62.955 178.845 64.015 178.885 ;
        RECT 61.435 178.715 64.015 178.845 ;
        RECT 64.275 178.755 64.990 178.925 ;
        RECT 65.160 178.780 65.415 179.685 ;
        RECT 61.435 178.665 63.180 178.715 ;
        RECT 61.465 177.985 61.915 178.495 ;
        RECT 62.105 178.295 62.580 178.495 ;
        RECT 62.330 177.895 62.580 178.295 ;
        RECT 62.830 178.295 63.180 178.495 ;
        RECT 62.830 177.895 63.040 178.295 ;
        RECT 63.350 178.215 63.675 178.545 ;
        RECT 63.845 178.045 64.015 178.715 ;
        RECT 64.185 178.205 64.540 178.575 ;
        RECT 64.820 178.545 64.990 178.755 ;
        RECT 64.820 178.215 65.075 178.545 ;
        RECT 63.285 177.875 64.015 178.045 ;
        RECT 64.820 178.025 64.990 178.215 ;
        RECT 65.245 178.050 65.415 178.780 ;
        RECT 65.590 178.705 65.850 179.855 ;
        RECT 66.025 178.715 66.365 179.685 ;
        RECT 66.535 178.715 66.705 179.855 ;
        RECT 66.975 179.055 67.225 179.855 ;
        RECT 67.870 178.885 68.200 179.685 ;
        RECT 68.500 179.055 68.830 179.855 ;
        RECT 69.000 178.885 69.330 179.685 ;
        RECT 66.895 178.715 69.330 178.885 ;
        RECT 69.745 178.715 69.975 179.855 ;
        RECT 58.020 177.475 59.320 177.685 ;
        RECT 59.575 177.305 59.905 177.665 ;
        RECT 60.075 177.475 60.335 177.805 ;
        RECT 61.435 177.305 61.885 177.815 ;
        RECT 63.285 177.725 63.465 177.875 ;
        RECT 62.160 177.475 63.465 177.725 ;
        RECT 64.275 177.855 64.990 178.025 ;
        RECT 63.645 177.305 63.975 177.705 ;
        RECT 64.275 177.475 64.445 177.855 ;
        RECT 64.660 177.305 64.990 177.685 ;
        RECT 65.160 177.475 65.415 178.050 ;
        RECT 65.590 177.305 65.850 178.145 ;
        RECT 66.025 178.105 66.200 178.715 ;
        RECT 66.895 178.465 67.065 178.715 ;
        RECT 66.370 178.295 67.065 178.465 ;
        RECT 67.240 178.295 67.660 178.495 ;
        RECT 67.830 178.295 68.160 178.495 ;
        RECT 68.330 178.295 68.660 178.495 ;
        RECT 66.025 177.475 66.365 178.105 ;
        RECT 66.535 177.305 66.785 178.105 ;
        RECT 66.975 177.955 68.200 178.125 ;
        RECT 66.975 177.475 67.305 177.955 ;
        RECT 67.475 177.305 67.700 177.765 ;
        RECT 67.870 177.475 68.200 177.955 ;
        RECT 68.830 178.085 69.000 178.715 ;
        RECT 70.145 178.705 70.475 179.685 ;
        RECT 70.645 178.715 70.855 179.855 ;
        RECT 71.095 179.045 71.390 179.855 ;
        RECT 69.185 178.295 69.535 178.545 ;
        RECT 69.725 178.295 70.055 178.545 ;
        RECT 68.830 177.475 69.330 178.085 ;
        RECT 69.745 177.305 69.975 178.125 ;
        RECT 70.225 178.105 70.475 178.705 ;
        RECT 71.570 178.545 71.815 179.685 ;
        RECT 71.990 179.045 72.250 179.855 ;
        RECT 72.850 179.850 79.125 179.855 ;
        RECT 72.430 178.545 72.680 179.680 ;
        RECT 72.850 179.055 73.110 179.850 ;
        RECT 73.280 178.955 73.540 179.680 ;
        RECT 73.710 179.125 73.970 179.850 ;
        RECT 74.140 178.955 74.400 179.680 ;
        RECT 74.570 179.125 74.830 179.850 ;
        RECT 75.000 178.955 75.260 179.680 ;
        RECT 75.430 179.125 75.690 179.850 ;
        RECT 75.860 178.955 76.120 179.680 ;
        RECT 76.290 179.125 76.535 179.850 ;
        RECT 76.705 178.955 76.965 179.680 ;
        RECT 77.150 179.125 77.395 179.850 ;
        RECT 77.565 178.955 77.825 179.680 ;
        RECT 78.010 179.125 78.255 179.850 ;
        RECT 78.425 178.955 78.685 179.680 ;
        RECT 78.870 179.125 79.125 179.850 ;
        RECT 73.280 178.940 78.685 178.955 ;
        RECT 79.295 178.940 79.585 179.680 ;
        RECT 79.755 179.110 80.025 179.855 ;
        RECT 73.280 178.715 80.025 178.940 ;
        RECT 70.145 177.475 70.475 178.105 ;
        RECT 70.645 177.305 70.855 178.125 ;
        RECT 71.085 177.985 71.400 178.545 ;
        RECT 71.570 178.295 78.690 178.545 ;
        RECT 71.085 177.305 71.390 177.815 ;
        RECT 71.570 177.485 71.820 178.295 ;
        RECT 71.990 177.305 72.250 177.830 ;
        RECT 72.430 177.485 72.680 178.295 ;
        RECT 78.860 178.125 80.025 178.715 ;
        RECT 80.290 178.885 80.565 179.685 ;
        RECT 80.735 179.055 81.065 179.855 ;
        RECT 81.235 179.515 82.375 179.685 ;
        RECT 81.235 178.885 81.405 179.515 ;
        RECT 80.290 178.675 81.405 178.885 ;
        RECT 81.575 178.885 81.905 179.345 ;
        RECT 82.075 179.055 82.375 179.515 ;
        RECT 81.575 178.665 82.335 178.885 ;
        RECT 82.585 178.690 82.875 179.855 ;
        RECT 83.050 178.855 83.305 179.855 ;
        RECT 80.290 178.295 81.010 178.495 ;
        RECT 81.180 178.295 81.950 178.495 ;
        RECT 82.120 178.125 82.335 178.665 ;
        RECT 73.280 177.955 80.025 178.125 ;
        RECT 72.850 177.305 73.110 177.865 ;
        RECT 73.280 177.500 73.540 177.955 ;
        RECT 73.710 177.305 73.970 177.785 ;
        RECT 74.140 177.500 74.400 177.955 ;
        RECT 74.570 177.305 74.830 177.785 ;
        RECT 75.000 177.500 75.260 177.955 ;
        RECT 75.430 177.305 75.675 177.785 ;
        RECT 75.845 177.500 76.120 177.955 ;
        RECT 76.290 177.305 76.535 177.785 ;
        RECT 76.705 177.500 76.965 177.955 ;
        RECT 77.145 177.305 77.395 177.785 ;
        RECT 77.565 177.500 77.825 177.955 ;
        RECT 78.005 177.305 78.255 177.785 ;
        RECT 78.425 177.500 78.685 177.955 ;
        RECT 78.865 177.305 79.125 177.785 ;
        RECT 79.295 177.500 79.555 177.955 ;
        RECT 79.725 177.305 80.025 177.785 ;
        RECT 80.290 177.305 80.565 178.125 ;
        RECT 80.735 177.955 82.335 178.125 ;
        RECT 80.735 177.945 81.905 177.955 ;
        RECT 80.735 177.475 81.065 177.945 ;
        RECT 81.235 177.305 81.405 177.775 ;
        RECT 81.575 177.475 81.905 177.945 ;
        RECT 82.075 177.305 82.365 177.775 ;
        RECT 82.585 177.305 82.875 178.030 ;
        RECT 83.065 177.305 83.305 178.105 ;
        RECT 83.490 177.475 83.735 179.685 ;
        RECT 83.905 179.405 84.755 179.855 ;
        RECT 84.925 179.225 85.185 179.685 ;
        RECT 84.065 179.005 85.185 179.225 ;
        RECT 85.365 179.175 85.570 179.205 ;
        RECT 85.365 179.005 85.575 179.175 ;
        RECT 84.065 178.550 84.235 179.005 ;
        RECT 83.905 178.060 84.235 178.550 ;
        RECT 84.405 178.230 84.815 178.835 ;
        RECT 85.365 178.620 85.570 179.005 ;
        RECT 85.755 178.870 86.080 179.855 ;
        RECT 86.355 178.925 86.525 179.685 ;
        RECT 86.740 179.095 87.070 179.855 ;
        RECT 86.355 178.755 87.070 178.925 ;
        RECT 87.240 178.780 87.495 179.685 ;
        RECT 84.985 178.245 85.570 178.620 ;
        RECT 85.825 178.215 86.085 178.670 ;
        RECT 86.265 178.205 86.620 178.575 ;
        RECT 86.900 178.545 87.070 178.755 ;
        RECT 86.900 178.215 87.155 178.545 ;
        RECT 83.905 177.855 84.755 178.060 ;
        RECT 83.905 177.305 84.235 177.685 ;
        RECT 84.425 177.475 84.755 177.855 ;
        RECT 84.925 177.855 86.080 178.045 ;
        RECT 86.900 178.025 87.070 178.215 ;
        RECT 87.325 178.050 87.495 178.780 ;
        RECT 87.670 178.705 87.930 179.855 ;
        RECT 88.105 178.765 89.315 179.855 ;
        RECT 88.105 178.225 88.625 178.765 ;
        RECT 84.925 177.685 85.135 177.855 ;
        RECT 85.805 177.715 86.080 177.855 ;
        RECT 86.355 177.855 87.070 178.025 ;
        RECT 85.305 177.305 85.635 177.685 ;
        RECT 86.355 177.475 86.525 177.855 ;
        RECT 86.740 177.305 87.070 177.685 ;
        RECT 87.240 177.475 87.495 178.050 ;
        RECT 87.670 177.305 87.930 178.145 ;
        RECT 88.795 178.055 89.315 178.595 ;
        RECT 88.105 177.305 89.315 178.055 ;
        RECT 18.100 177.135 89.400 177.305 ;
        RECT 18.185 176.385 19.395 177.135 ;
        RECT 19.655 176.585 19.825 176.965 ;
        RECT 20.005 176.755 20.335 177.135 ;
        RECT 19.655 176.415 20.320 176.585 ;
        RECT 20.515 176.460 20.775 176.965 ;
        RECT 18.185 175.845 18.705 176.385 ;
        RECT 18.875 175.675 19.395 176.215 ;
        RECT 19.585 175.865 19.925 176.235 ;
        RECT 20.150 176.160 20.320 176.415 ;
        RECT 20.150 175.830 20.425 176.160 ;
        RECT 20.150 175.685 20.320 175.830 ;
        RECT 18.185 174.585 19.395 175.675 ;
        RECT 19.645 175.515 20.320 175.685 ;
        RECT 20.595 175.660 20.775 176.460 ;
        RECT 21.870 176.485 22.140 176.695 ;
        RECT 22.360 176.675 22.690 177.135 ;
        RECT 23.200 176.675 23.950 176.965 ;
        RECT 21.870 176.315 23.205 176.485 ;
        RECT 23.035 176.145 23.205 176.315 ;
        RECT 21.870 175.905 22.220 176.145 ;
        RECT 22.390 175.905 22.865 176.145 ;
        RECT 23.035 175.895 23.410 176.145 ;
        RECT 23.035 175.725 23.205 175.895 ;
        RECT 19.645 174.755 19.825 175.515 ;
        RECT 20.005 174.585 20.335 175.345 ;
        RECT 20.505 174.755 20.775 175.660 ;
        RECT 21.870 175.555 23.205 175.725 ;
        RECT 21.870 175.395 22.150 175.555 ;
        RECT 23.580 175.385 23.950 176.675 ;
        RECT 24.170 176.295 24.430 177.135 ;
        RECT 24.605 176.390 24.860 176.965 ;
        RECT 25.030 176.755 25.360 177.135 ;
        RECT 25.575 176.585 25.745 176.965 ;
        RECT 25.030 176.415 25.745 176.585 ;
        RECT 26.005 176.460 26.265 176.965 ;
        RECT 26.445 176.755 26.775 177.135 ;
        RECT 26.955 176.585 27.125 176.965 ;
        RECT 22.360 174.585 22.610 175.385 ;
        RECT 22.780 175.215 23.950 175.385 ;
        RECT 22.780 174.755 23.110 175.215 ;
        RECT 23.280 174.585 23.495 175.045 ;
        RECT 24.170 174.585 24.430 175.735 ;
        RECT 24.605 175.660 24.775 176.390 ;
        RECT 25.030 176.225 25.200 176.415 ;
        RECT 24.945 175.895 25.200 176.225 ;
        RECT 25.030 175.685 25.200 175.895 ;
        RECT 25.480 175.865 25.835 176.235 ;
        RECT 24.605 174.755 24.860 175.660 ;
        RECT 25.030 175.515 25.745 175.685 ;
        RECT 25.030 174.585 25.360 175.345 ;
        RECT 25.575 174.755 25.745 175.515 ;
        RECT 26.005 175.660 26.175 176.460 ;
        RECT 26.460 176.415 27.125 176.585 ;
        RECT 27.475 176.585 27.645 176.965 ;
        RECT 27.825 176.755 28.155 177.135 ;
        RECT 27.475 176.415 28.140 176.585 ;
        RECT 28.335 176.460 28.595 176.965 ;
        RECT 26.460 176.160 26.630 176.415 ;
        RECT 26.345 175.830 26.630 176.160 ;
        RECT 26.865 175.865 27.195 176.235 ;
        RECT 27.405 175.865 27.735 176.235 ;
        RECT 27.970 176.160 28.140 176.415 ;
        RECT 26.460 175.685 26.630 175.830 ;
        RECT 27.970 175.830 28.255 176.160 ;
        RECT 27.970 175.685 28.140 175.830 ;
        RECT 26.005 174.755 26.275 175.660 ;
        RECT 26.460 175.515 27.125 175.685 ;
        RECT 26.445 174.585 26.775 175.345 ;
        RECT 26.955 174.755 27.125 175.515 ;
        RECT 27.475 175.515 28.140 175.685 ;
        RECT 28.425 175.660 28.595 176.460 ;
        RECT 28.765 176.365 32.275 177.135 ;
        RECT 28.765 175.845 30.415 176.365 ;
        RECT 33.365 176.335 33.675 177.135 ;
        RECT 33.880 176.335 34.575 176.965 ;
        RECT 34.745 176.590 40.090 177.135 ;
        RECT 33.880 176.285 34.055 176.335 ;
        RECT 30.585 175.675 32.275 176.195 ;
        RECT 33.375 175.895 33.710 176.165 ;
        RECT 33.880 175.735 34.050 176.285 ;
        RECT 34.220 175.895 34.555 176.145 ;
        RECT 36.330 175.760 36.670 176.590 ;
        RECT 40.265 176.365 43.775 177.135 ;
        RECT 43.945 176.410 44.235 177.135 ;
        RECT 44.490 176.635 44.985 176.965 ;
        RECT 27.475 174.755 27.645 175.515 ;
        RECT 27.825 174.585 28.155 175.345 ;
        RECT 28.325 174.755 28.595 175.660 ;
        RECT 28.765 174.585 32.275 175.675 ;
        RECT 33.365 174.585 33.645 175.725 ;
        RECT 33.815 174.755 34.145 175.735 ;
        RECT 34.315 174.585 34.575 175.725 ;
        RECT 38.150 175.020 38.500 176.270 ;
        RECT 40.265 175.845 41.915 176.365 ;
        RECT 42.085 175.675 43.775 176.195 ;
        RECT 34.745 174.585 40.090 175.020 ;
        RECT 40.265 174.585 43.775 175.675 ;
        RECT 43.945 174.585 44.235 175.750 ;
        RECT 44.405 175.145 44.645 176.455 ;
        RECT 44.815 175.725 44.985 176.635 ;
        RECT 45.205 175.895 45.555 176.860 ;
        RECT 45.735 175.895 46.035 176.865 ;
        RECT 46.215 175.895 46.495 176.865 ;
        RECT 46.675 176.335 46.945 177.135 ;
        RECT 47.115 176.415 47.455 176.925 ;
        RECT 47.650 176.745 47.980 177.135 ;
        RECT 48.150 176.575 48.375 176.955 ;
        RECT 46.690 175.895 47.020 176.145 ;
        RECT 46.690 175.725 47.005 175.895 ;
        RECT 44.815 175.555 47.005 175.725 ;
        RECT 44.410 174.585 44.745 174.965 ;
        RECT 44.915 174.755 45.165 175.555 ;
        RECT 45.385 174.585 45.715 175.305 ;
        RECT 45.900 174.755 46.150 175.555 ;
        RECT 46.615 174.585 46.945 175.385 ;
        RECT 47.195 175.015 47.455 176.415 ;
        RECT 47.635 175.895 47.875 176.545 ;
        RECT 48.045 176.395 48.375 176.575 ;
        RECT 48.045 175.725 48.220 176.395 ;
        RECT 48.575 176.225 48.805 176.845 ;
        RECT 48.985 176.405 49.285 177.135 ;
        RECT 49.925 176.335 50.620 176.965 ;
        RECT 50.825 176.335 51.135 177.135 ;
        RECT 51.305 176.460 51.565 176.965 ;
        RECT 51.745 176.755 52.075 177.135 ;
        RECT 52.255 176.585 52.425 176.965 ;
        RECT 48.390 175.895 48.805 176.225 ;
        RECT 48.985 175.895 49.280 176.225 ;
        RECT 49.945 175.895 50.280 176.145 ;
        RECT 50.450 175.735 50.620 176.335 ;
        RECT 50.790 175.895 51.125 176.165 ;
        RECT 47.115 174.755 47.455 175.015 ;
        RECT 47.635 175.535 48.220 175.725 ;
        RECT 47.635 174.765 47.910 175.535 ;
        RECT 48.390 175.365 49.285 175.695 ;
        RECT 48.080 175.195 49.285 175.365 ;
        RECT 48.080 174.765 48.410 175.195 ;
        RECT 48.580 174.585 48.775 175.025 ;
        RECT 48.955 174.765 49.285 175.195 ;
        RECT 49.925 174.585 50.185 175.725 ;
        RECT 50.355 174.755 50.685 175.735 ;
        RECT 50.855 174.585 51.135 175.725 ;
        RECT 51.305 175.660 51.475 176.460 ;
        RECT 51.760 176.415 52.425 176.585 ;
        RECT 52.685 176.460 52.945 176.965 ;
        RECT 53.125 176.755 53.455 177.135 ;
        RECT 53.635 176.585 53.805 176.965 ;
        RECT 51.760 176.160 51.930 176.415 ;
        RECT 51.645 175.830 51.930 176.160 ;
        RECT 52.165 175.865 52.495 176.235 ;
        RECT 51.760 175.685 51.930 175.830 ;
        RECT 51.305 174.755 51.575 175.660 ;
        RECT 51.760 175.515 52.425 175.685 ;
        RECT 51.745 174.585 52.075 175.345 ;
        RECT 52.255 174.755 52.425 175.515 ;
        RECT 52.685 175.660 52.865 176.460 ;
        RECT 53.140 176.415 53.805 176.585 ;
        RECT 53.140 176.160 53.310 176.415 ;
        RECT 54.065 176.335 54.760 176.965 ;
        RECT 54.965 176.335 55.275 177.135 ;
        RECT 55.445 176.460 55.705 176.965 ;
        RECT 55.885 176.755 56.215 177.135 ;
        RECT 56.395 176.585 56.565 176.965 ;
        RECT 53.035 175.830 53.310 176.160 ;
        RECT 53.535 175.865 53.875 176.235 ;
        RECT 54.085 175.895 54.420 176.145 ;
        RECT 53.140 175.685 53.310 175.830 ;
        RECT 54.590 175.775 54.760 176.335 ;
        RECT 54.930 175.895 55.265 176.165 ;
        RECT 54.585 175.735 54.760 175.775 ;
        RECT 52.685 174.755 52.955 175.660 ;
        RECT 53.140 175.515 53.815 175.685 ;
        RECT 53.125 174.585 53.455 175.345 ;
        RECT 53.635 174.755 53.815 175.515 ;
        RECT 54.065 174.585 54.325 175.725 ;
        RECT 54.495 174.755 54.825 175.735 ;
        RECT 54.995 174.585 55.275 175.725 ;
        RECT 55.445 175.660 55.625 176.460 ;
        RECT 55.900 176.415 56.565 176.585 ;
        RECT 55.900 176.160 56.070 176.415 ;
        RECT 55.795 175.830 56.070 176.160 ;
        RECT 56.295 175.865 56.635 176.235 ;
        RECT 55.900 175.685 56.070 175.830 ;
        RECT 55.445 174.755 55.715 175.660 ;
        RECT 55.900 175.515 56.575 175.685 ;
        RECT 55.885 174.585 56.215 175.345 ;
        RECT 56.395 174.755 56.575 175.515 ;
        RECT 56.840 174.765 57.120 176.955 ;
        RECT 57.320 176.765 58.050 177.135 ;
        RECT 58.630 176.595 59.060 176.955 ;
        RECT 57.320 176.405 59.060 176.595 ;
        RECT 57.320 175.895 57.580 176.405 ;
        RECT 57.310 174.585 57.595 175.725 ;
        RECT 57.790 175.605 58.050 176.225 ;
        RECT 58.245 175.605 58.670 176.225 ;
        RECT 58.840 176.175 59.060 176.405 ;
        RECT 59.230 176.355 59.475 177.135 ;
        RECT 58.840 175.875 59.385 176.175 ;
        RECT 59.675 176.055 59.905 176.955 ;
        RECT 57.860 175.235 58.885 175.435 ;
        RECT 57.860 174.765 58.030 175.235 ;
        RECT 58.205 174.585 58.535 175.065 ;
        RECT 58.705 174.765 58.885 175.235 ;
        RECT 59.055 174.765 59.385 175.875 ;
        RECT 59.565 175.375 59.905 176.055 ;
        RECT 60.085 175.555 60.315 176.895 ;
        RECT 60.505 176.335 61.200 176.965 ;
        RECT 61.405 176.335 61.715 177.135 ;
        RECT 61.895 176.625 62.345 177.135 ;
        RECT 62.620 176.715 63.925 176.965 ;
        RECT 64.105 176.735 64.435 177.135 ;
        RECT 63.745 176.565 63.925 176.715 ;
        RECT 60.525 175.895 60.860 176.145 ;
        RECT 61.030 175.735 61.200 176.335 ;
        RECT 61.370 175.895 61.705 176.165 ;
        RECT 61.925 175.945 62.375 176.455 ;
        RECT 62.790 176.145 63.040 176.545 ;
        RECT 62.565 175.945 63.040 176.145 ;
        RECT 63.290 176.145 63.500 176.545 ;
        RECT 63.745 176.395 64.475 176.565 ;
        RECT 63.290 175.945 63.640 176.145 ;
        RECT 63.810 175.895 64.135 176.225 ;
        RECT 59.565 175.175 60.315 175.375 ;
        RECT 59.555 174.585 59.905 174.995 ;
        RECT 60.075 174.785 60.315 175.175 ;
        RECT 60.505 174.585 60.765 175.725 ;
        RECT 60.935 174.755 61.265 175.735 ;
        RECT 61.895 175.725 63.640 175.775 ;
        RECT 64.305 175.725 64.475 176.395 ;
        RECT 61.435 174.585 61.715 175.725 ;
        RECT 61.895 175.595 64.475 175.725 ;
        RECT 61.895 174.925 62.225 175.595 ;
        RECT 63.415 175.555 64.475 175.595 ;
        RECT 65.105 176.410 65.365 176.965 ;
        RECT 65.535 176.690 65.965 177.135 ;
        RECT 66.200 176.565 66.370 176.965 ;
        RECT 66.540 176.735 67.260 177.135 ;
        RECT 65.105 175.695 65.280 176.410 ;
        RECT 66.200 176.395 67.080 176.565 ;
        RECT 67.430 176.520 67.600 176.965 ;
        RECT 68.175 176.625 68.575 177.135 ;
        RECT 65.450 175.895 65.705 176.225 ;
        RECT 62.395 175.385 63.275 175.425 ;
        RECT 62.395 175.185 63.925 175.385 ;
        RECT 62.395 175.135 63.010 175.185 ;
        RECT 62.395 175.095 62.625 175.135 ;
        RECT 63.755 175.055 63.925 175.185 ;
        RECT 62.735 174.925 63.065 174.965 ;
        RECT 61.895 174.755 63.065 174.925 ;
        RECT 63.235 174.585 63.610 174.965 ;
        RECT 64.160 174.585 64.425 175.365 ;
        RECT 65.105 174.755 65.365 175.695 ;
        RECT 65.535 175.415 65.705 175.895 ;
        RECT 65.930 175.605 66.260 176.225 ;
        RECT 66.430 175.845 66.720 176.225 ;
        RECT 66.910 175.675 67.080 176.395 ;
        RECT 66.560 175.505 67.080 175.675 ;
        RECT 67.250 176.350 67.600 176.520 ;
        RECT 65.535 175.245 66.295 175.415 ;
        RECT 66.560 175.315 66.730 175.505 ;
        RECT 67.250 175.325 67.420 176.350 ;
        RECT 67.840 175.865 68.100 176.455 ;
        RECT 67.620 175.565 68.100 175.865 ;
        RECT 68.300 175.565 68.560 176.455 ;
        RECT 69.705 176.410 69.995 177.135 ;
        RECT 70.165 176.635 70.425 176.965 ;
        RECT 70.595 176.775 70.925 177.135 ;
        RECT 71.180 176.755 72.480 176.965 ;
        RECT 66.125 175.020 66.295 175.245 ;
        RECT 67.010 175.155 67.420 175.325 ;
        RECT 67.595 175.215 68.535 175.385 ;
        RECT 67.010 175.020 67.265 175.155 ;
        RECT 65.535 174.585 65.865 174.985 ;
        RECT 66.125 174.850 67.265 175.020 ;
        RECT 67.595 174.965 67.765 175.215 ;
        RECT 67.010 174.755 67.265 174.850 ;
        RECT 67.435 174.795 67.765 174.965 ;
        RECT 67.935 174.585 68.185 175.045 ;
        RECT 68.355 174.755 68.535 175.215 ;
        RECT 69.705 174.585 69.995 175.750 ;
        RECT 70.165 175.435 70.335 176.635 ;
        RECT 71.180 176.605 71.350 176.755 ;
        RECT 70.595 176.480 71.350 176.605 ;
        RECT 70.505 176.435 71.350 176.480 ;
        RECT 70.505 176.315 70.775 176.435 ;
        RECT 70.505 175.740 70.675 176.315 ;
        RECT 70.905 175.875 71.315 176.180 ;
        RECT 71.605 176.145 71.815 176.545 ;
        RECT 71.485 175.935 71.815 176.145 ;
        RECT 72.060 176.145 72.280 176.545 ;
        RECT 72.755 176.370 73.210 177.135 ;
        RECT 73.870 176.380 74.105 176.710 ;
        RECT 74.275 176.395 74.605 177.135 ;
        RECT 74.840 176.755 76.035 176.965 ;
        RECT 72.060 175.935 72.535 176.145 ;
        RECT 72.725 175.945 73.215 176.145 ;
        RECT 70.505 175.705 70.705 175.740 ;
        RECT 72.035 175.705 73.210 175.765 ;
        RECT 70.505 175.595 73.210 175.705 ;
        RECT 70.565 175.535 72.365 175.595 ;
        RECT 72.035 175.505 72.365 175.535 ;
        RECT 70.165 174.755 70.425 175.435 ;
        RECT 70.595 174.585 70.845 175.365 ;
        RECT 71.095 175.335 71.930 175.345 ;
        RECT 72.520 175.335 72.705 175.425 ;
        RECT 71.095 175.135 72.705 175.335 ;
        RECT 71.095 174.755 71.345 175.135 ;
        RECT 72.475 175.095 72.705 175.135 ;
        RECT 72.955 174.975 73.210 175.595 ;
        RECT 73.870 175.725 74.040 176.380 ;
        RECT 74.840 176.315 75.115 176.755 ;
        RECT 75.285 176.415 75.615 176.585 ;
        RECT 75.290 176.315 75.615 176.415 ;
        RECT 75.785 176.525 76.035 176.755 ;
        RECT 76.205 176.695 76.375 177.135 ;
        RECT 76.545 176.525 76.895 176.965 ;
        RECT 77.985 176.625 78.290 177.135 ;
        RECT 75.785 176.315 76.895 176.525 ;
        RECT 74.215 175.895 74.560 176.225 ;
        RECT 74.790 175.725 75.120 176.145 ;
        RECT 73.870 175.555 75.120 175.725 ;
        RECT 73.870 175.360 74.170 175.555 ;
        RECT 75.290 175.385 75.570 176.315 ;
        RECT 75.750 175.945 76.895 176.145 ;
        RECT 75.750 175.775 75.940 175.945 ;
        RECT 77.985 175.895 78.300 176.455 ;
        RECT 78.470 176.145 78.720 176.955 ;
        RECT 78.890 176.610 79.150 177.135 ;
        RECT 79.330 176.145 79.580 176.955 ;
        RECT 79.750 176.575 80.010 177.135 ;
        RECT 80.180 176.485 80.440 176.940 ;
        RECT 80.610 176.655 80.870 177.135 ;
        RECT 81.040 176.485 81.300 176.940 ;
        RECT 81.470 176.655 81.730 177.135 ;
        RECT 81.900 176.485 82.160 176.940 ;
        RECT 82.330 176.655 82.575 177.135 ;
        RECT 82.745 176.485 83.020 176.940 ;
        RECT 83.190 176.655 83.435 177.135 ;
        RECT 83.605 176.485 83.865 176.940 ;
        RECT 84.045 176.655 84.295 177.135 ;
        RECT 84.465 176.485 84.725 176.940 ;
        RECT 84.905 176.655 85.155 177.135 ;
        RECT 85.325 176.485 85.585 176.940 ;
        RECT 85.765 176.655 86.025 177.135 ;
        RECT 86.195 176.485 86.455 176.940 ;
        RECT 86.625 176.655 86.925 177.135 ;
        RECT 80.180 176.315 86.925 176.485 ;
        RECT 88.105 176.385 89.315 177.135 ;
        RECT 78.470 175.895 85.590 176.145 ;
        RECT 75.745 175.605 75.940 175.775 ;
        RECT 76.205 175.725 76.375 175.775 ;
        RECT 75.750 175.565 75.940 175.605 ;
        RECT 76.120 175.385 76.395 175.725 ;
        RECT 71.515 174.585 71.870 174.965 ;
        RECT 72.875 174.755 73.210 174.975 ;
        RECT 74.340 174.585 74.595 175.385 ;
        RECT 74.795 175.215 76.395 175.385 ;
        RECT 74.795 174.755 75.125 175.215 ;
        RECT 75.295 174.585 75.870 175.045 ;
        RECT 76.040 174.755 76.395 175.215 ;
        RECT 76.565 174.585 76.895 175.725 ;
        RECT 77.995 174.585 78.290 175.395 ;
        RECT 78.470 174.755 78.715 175.895 ;
        RECT 78.890 174.585 79.150 175.395 ;
        RECT 79.330 174.760 79.580 175.895 ;
        RECT 85.760 175.725 86.925 176.315 ;
        RECT 80.180 175.500 86.925 175.725 ;
        RECT 88.105 175.675 88.625 176.215 ;
        RECT 88.795 175.845 89.315 176.385 ;
        RECT 80.180 175.485 85.585 175.500 ;
        RECT 79.750 174.590 80.010 175.385 ;
        RECT 80.180 174.760 80.440 175.485 ;
        RECT 80.610 174.590 80.870 175.315 ;
        RECT 81.040 174.760 81.300 175.485 ;
        RECT 81.470 174.590 81.730 175.315 ;
        RECT 81.900 174.760 82.160 175.485 ;
        RECT 82.330 174.590 82.590 175.315 ;
        RECT 82.760 174.760 83.020 175.485 ;
        RECT 83.190 174.590 83.435 175.315 ;
        RECT 83.605 174.760 83.865 175.485 ;
        RECT 84.050 174.590 84.295 175.315 ;
        RECT 84.465 174.760 84.725 175.485 ;
        RECT 84.910 174.590 85.155 175.315 ;
        RECT 85.325 174.760 85.585 175.485 ;
        RECT 85.770 174.590 86.025 175.315 ;
        RECT 86.195 174.760 86.485 175.500 ;
        RECT 79.750 174.585 86.025 174.590 ;
        RECT 86.655 174.585 86.925 175.330 ;
        RECT 88.105 174.585 89.315 175.675 ;
        RECT 18.100 174.415 89.400 174.585 ;
        RECT 18.185 173.325 19.395 174.415 ;
        RECT 18.185 172.615 18.705 173.155 ;
        RECT 18.875 172.785 19.395 173.325 ;
        RECT 18.185 171.865 19.395 172.615 ;
        RECT 20.485 172.145 20.765 174.245 ;
        RECT 20.955 173.655 21.740 174.415 ;
        RECT 22.135 173.585 22.520 174.245 ;
        RECT 22.135 173.485 22.545 173.585 ;
        RECT 20.935 173.275 22.545 173.485 ;
        RECT 22.845 173.395 23.045 174.185 ;
        RECT 20.935 172.675 21.210 173.275 ;
        RECT 22.715 173.225 23.045 173.395 ;
        RECT 23.215 173.235 23.535 174.415 ;
        RECT 23.705 173.980 29.050 174.415 ;
        RECT 22.715 173.105 22.895 173.225 ;
        RECT 21.380 172.855 21.735 173.105 ;
        RECT 21.930 173.055 22.395 173.105 ;
        RECT 21.925 172.885 22.395 173.055 ;
        RECT 21.930 172.855 22.395 172.885 ;
        RECT 22.565 172.855 22.895 173.105 ;
        RECT 23.070 172.855 23.535 173.055 ;
        RECT 20.935 172.495 22.185 172.675 ;
        RECT 21.820 172.425 22.185 172.495 ;
        RECT 22.355 172.475 23.535 172.645 ;
        RECT 20.995 171.865 21.165 172.325 ;
        RECT 22.355 172.255 22.685 172.475 ;
        RECT 21.435 172.075 22.685 172.255 ;
        RECT 22.855 171.865 23.025 172.305 ;
        RECT 23.195 172.060 23.535 172.475 ;
        RECT 25.290 172.410 25.630 173.240 ;
        RECT 27.110 172.730 27.460 173.980 ;
        RECT 29.225 173.325 30.895 174.415 ;
        RECT 29.225 172.635 29.975 173.155 ;
        RECT 30.145 172.805 30.895 173.325 ;
        RECT 31.065 173.250 31.355 174.415 ;
        RECT 31.545 173.525 31.805 174.235 ;
        RECT 31.975 173.705 32.305 174.415 ;
        RECT 32.475 173.525 32.705 174.235 ;
        RECT 31.545 173.285 32.705 173.525 ;
        RECT 32.885 173.505 33.155 174.235 ;
        RECT 33.335 173.685 33.675 174.415 ;
        RECT 32.885 173.285 33.655 173.505 ;
        RECT 31.535 172.775 31.835 173.105 ;
        RECT 32.015 172.795 32.540 173.105 ;
        RECT 32.720 172.795 33.185 173.105 ;
        RECT 23.705 171.865 29.050 172.410 ;
        RECT 29.225 171.865 30.895 172.635 ;
        RECT 31.065 171.865 31.355 172.590 ;
        RECT 31.545 171.865 31.835 172.595 ;
        RECT 32.015 172.155 32.245 172.795 ;
        RECT 33.365 172.615 33.655 173.285 ;
        RECT 32.425 172.415 33.655 172.615 ;
        RECT 32.425 172.045 32.735 172.415 ;
        RECT 32.915 171.865 33.585 172.235 ;
        RECT 33.845 172.045 34.105 174.235 ;
        RECT 34.285 173.325 37.795 174.415 ;
        RECT 34.285 172.635 35.935 173.155 ;
        RECT 36.105 172.805 37.795 173.325 ;
        RECT 38.425 173.275 38.685 174.415 ;
        RECT 38.855 173.265 39.185 174.245 ;
        RECT 39.355 173.275 39.635 174.415 ;
        RECT 39.805 173.980 45.150 174.415 ;
        RECT 45.325 173.980 50.670 174.415 ;
        RECT 38.445 172.855 38.780 173.105 ;
        RECT 38.950 172.665 39.120 173.265 ;
        RECT 39.290 172.835 39.625 173.105 ;
        RECT 34.285 171.865 37.795 172.635 ;
        RECT 38.425 172.035 39.120 172.665 ;
        RECT 39.325 171.865 39.635 172.665 ;
        RECT 41.390 172.410 41.730 173.240 ;
        RECT 43.210 172.730 43.560 173.980 ;
        RECT 46.910 172.410 47.250 173.240 ;
        RECT 48.730 172.730 49.080 173.980 ;
        RECT 51.775 173.465 52.050 174.235 ;
        RECT 52.220 173.805 52.550 174.235 ;
        RECT 52.720 173.975 52.915 174.415 ;
        RECT 53.095 173.805 53.425 174.235 ;
        RECT 52.220 173.635 53.425 173.805 ;
        RECT 51.775 173.275 52.360 173.465 ;
        RECT 52.530 173.305 53.425 173.635 ;
        RECT 54.535 173.465 54.810 174.235 ;
        RECT 54.980 173.805 55.310 174.235 ;
        RECT 55.480 173.975 55.675 174.415 ;
        RECT 55.855 173.805 56.185 174.235 ;
        RECT 54.980 173.635 56.185 173.805 ;
        RECT 54.535 173.275 55.120 173.465 ;
        RECT 55.290 173.305 56.185 173.635 ;
        RECT 51.775 172.455 52.015 173.105 ;
        RECT 52.185 172.605 52.360 173.275 ;
        RECT 52.530 172.775 52.945 173.105 ;
        RECT 53.125 172.775 53.420 173.105 ;
        RECT 52.185 172.425 52.515 172.605 ;
        RECT 39.805 171.865 45.150 172.410 ;
        RECT 45.325 171.865 50.670 172.410 ;
        RECT 51.790 171.865 52.120 172.255 ;
        RECT 52.290 172.045 52.515 172.425 ;
        RECT 52.715 172.155 52.945 172.775 ;
        RECT 53.125 171.865 53.425 172.595 ;
        RECT 54.535 172.455 54.775 173.105 ;
        RECT 54.945 172.605 55.120 173.275 ;
        RECT 56.825 173.250 57.115 174.415 ;
        RECT 57.745 173.340 58.015 174.245 ;
        RECT 58.185 173.655 58.515 174.415 ;
        RECT 58.695 173.485 58.875 174.245 ;
        RECT 55.290 172.775 55.705 173.105 ;
        RECT 55.885 172.775 56.180 173.105 ;
        RECT 54.945 172.425 55.275 172.605 ;
        RECT 54.550 171.865 54.880 172.255 ;
        RECT 55.050 172.045 55.275 172.425 ;
        RECT 55.475 172.155 55.705 172.775 ;
        RECT 55.885 171.865 56.185 172.595 ;
        RECT 56.825 171.865 57.115 172.590 ;
        RECT 57.745 172.540 57.925 173.340 ;
        RECT 58.200 173.315 58.875 173.485 ;
        RECT 58.200 173.170 58.370 173.315 ;
        RECT 59.165 173.275 59.395 174.415 ;
        RECT 59.565 173.265 59.895 174.245 ;
        RECT 60.065 173.275 60.275 174.415 ;
        RECT 60.505 173.275 60.785 174.415 ;
        RECT 60.955 173.265 61.285 174.245 ;
        RECT 61.455 173.275 61.715 174.415 ;
        RECT 61.885 173.565 62.145 174.245 ;
        RECT 62.315 173.635 62.565 174.415 ;
        RECT 62.815 173.865 63.065 174.245 ;
        RECT 63.235 174.035 63.590 174.415 ;
        RECT 64.595 174.025 64.930 174.245 ;
        RECT 64.195 173.865 64.425 173.905 ;
        RECT 62.815 173.665 64.425 173.865 ;
        RECT 62.815 173.655 63.650 173.665 ;
        RECT 64.240 173.575 64.425 173.665 ;
        RECT 58.095 172.840 58.370 173.170 ;
        RECT 58.200 172.585 58.370 172.840 ;
        RECT 58.595 172.765 58.935 173.135 ;
        RECT 59.145 172.855 59.475 173.105 ;
        RECT 57.745 172.035 58.005 172.540 ;
        RECT 58.200 172.415 58.865 172.585 ;
        RECT 58.185 171.865 58.515 172.245 ;
        RECT 58.695 172.035 58.865 172.415 ;
        RECT 59.165 171.865 59.395 172.685 ;
        RECT 59.645 172.665 59.895 173.265 ;
        RECT 60.515 172.835 60.850 173.105 ;
        RECT 59.565 172.035 59.895 172.665 ;
        RECT 60.065 171.865 60.275 172.685 ;
        RECT 61.020 172.665 61.190 173.265 ;
        RECT 61.360 172.855 61.695 173.105 ;
        RECT 60.505 171.865 60.815 172.665 ;
        RECT 61.020 172.035 61.715 172.665 ;
        RECT 61.885 172.365 62.055 173.565 ;
        RECT 63.755 173.465 64.085 173.495 ;
        RECT 62.285 173.405 64.085 173.465 ;
        RECT 64.675 173.405 64.930 174.025 ;
        RECT 62.225 173.295 64.930 173.405 ;
        RECT 62.225 173.260 62.425 173.295 ;
        RECT 62.225 172.685 62.395 173.260 ;
        RECT 63.755 173.235 64.930 173.295 ;
        RECT 65.565 173.340 65.835 174.245 ;
        RECT 66.005 173.655 66.335 174.415 ;
        RECT 66.515 173.485 66.695 174.245 ;
        RECT 62.625 172.820 63.035 173.125 ;
        RECT 63.205 172.855 63.535 173.065 ;
        RECT 62.225 172.565 62.495 172.685 ;
        RECT 62.225 172.520 63.070 172.565 ;
        RECT 62.315 172.395 63.070 172.520 ;
        RECT 63.325 172.455 63.535 172.855 ;
        RECT 63.780 172.855 64.255 173.065 ;
        RECT 64.445 172.855 64.935 173.055 ;
        RECT 63.780 172.455 64.000 172.855 ;
        RECT 61.885 172.035 62.145 172.365 ;
        RECT 62.900 172.245 63.070 172.395 ;
        RECT 62.315 171.865 62.645 172.225 ;
        RECT 62.900 172.035 64.200 172.245 ;
        RECT 64.475 171.865 64.930 172.630 ;
        RECT 65.565 172.540 65.745 173.340 ;
        RECT 66.020 173.315 66.695 173.485 ;
        RECT 66.020 173.170 66.190 173.315 ;
        RECT 66.955 173.275 67.285 174.415 ;
        RECT 67.815 173.445 68.145 174.230 ;
        RECT 67.465 173.275 68.145 173.445 ;
        RECT 68.365 173.275 68.595 174.415 ;
        RECT 65.915 172.840 66.190 173.170 ;
        RECT 66.020 172.585 66.190 172.840 ;
        RECT 66.415 172.765 66.755 173.135 ;
        RECT 66.945 172.855 67.295 173.105 ;
        RECT 67.465 172.675 67.635 173.275 ;
        RECT 68.765 173.265 69.095 174.245 ;
        RECT 69.265 173.275 69.475 174.415 ;
        RECT 69.810 173.615 70.065 174.415 ;
        RECT 70.235 173.445 70.565 174.245 ;
        RECT 70.735 173.615 70.905 174.415 ;
        RECT 71.075 173.445 71.405 174.245 ;
        RECT 69.705 173.275 71.405 173.445 ;
        RECT 71.575 173.275 71.835 174.415 ;
        RECT 72.210 173.975 72.540 174.415 ;
        RECT 72.710 173.805 72.945 174.245 ;
        RECT 73.130 174.035 73.460 174.415 ;
        RECT 73.670 173.805 74.015 174.245 ;
        RECT 72.005 173.565 74.015 173.805 ;
        RECT 67.805 172.855 68.155 173.105 ;
        RECT 68.345 172.855 68.675 173.105 ;
        RECT 65.565 172.035 65.825 172.540 ;
        RECT 66.020 172.415 66.685 172.585 ;
        RECT 66.005 171.865 66.335 172.245 ;
        RECT 66.515 172.035 66.685 172.415 ;
        RECT 66.955 171.865 67.225 172.675 ;
        RECT 67.395 172.035 67.725 172.675 ;
        RECT 67.895 171.865 68.135 172.675 ;
        RECT 68.365 171.865 68.595 172.685 ;
        RECT 68.845 172.665 69.095 173.265 ;
        RECT 69.705 172.685 69.985 173.275 ;
        RECT 70.155 172.855 70.905 173.105 ;
        RECT 71.075 172.855 71.835 173.105 ;
        RECT 68.765 172.035 69.095 172.665 ;
        RECT 69.265 171.865 69.475 172.685 ;
        RECT 69.705 172.435 70.565 172.685 ;
        RECT 72.005 172.665 72.235 173.565 ;
        RECT 74.190 173.395 74.535 174.150 ;
        RECT 74.705 173.575 75.035 174.415 ;
        RECT 75.245 173.575 75.575 174.415 ;
        RECT 75.745 173.395 76.090 174.150 ;
        RECT 76.265 173.805 76.610 174.245 ;
        RECT 76.820 174.035 77.150 174.415 ;
        RECT 77.335 173.805 77.570 174.245 ;
        RECT 77.740 173.975 78.070 174.415 ;
        RECT 76.265 173.565 78.275 173.805 ;
        RECT 72.405 172.855 72.735 173.395 ;
        RECT 70.735 172.495 71.835 172.665 ;
        RECT 69.815 172.245 70.145 172.265 ;
        RECT 70.735 172.245 70.985 172.495 ;
        RECT 69.815 172.035 70.985 172.245 ;
        RECT 71.155 171.865 71.325 172.325 ;
        RECT 71.495 172.035 71.835 172.495 ;
        RECT 72.005 172.035 72.610 172.665 ;
        RECT 72.945 172.035 73.275 173.395 ;
        RECT 73.445 172.775 73.735 173.395 ;
        RECT 73.905 172.775 74.535 173.395 ;
        RECT 74.705 172.785 75.035 173.395 ;
        RECT 75.245 172.785 75.575 173.395 ;
        RECT 75.745 172.775 76.375 173.395 ;
        RECT 76.545 172.775 76.835 173.395 ;
        RECT 73.670 172.405 75.035 172.605 ;
        RECT 73.670 172.035 74.015 172.405 ;
        RECT 74.205 171.865 74.535 172.235 ;
        RECT 74.705 172.035 75.035 172.405 ;
        RECT 75.245 172.405 76.610 172.605 ;
        RECT 75.245 172.035 75.575 172.405 ;
        RECT 75.745 171.865 76.075 172.235 ;
        RECT 76.265 172.035 76.610 172.405 ;
        RECT 77.005 172.035 77.335 173.395 ;
        RECT 77.545 172.855 77.875 173.395 ;
        RECT 78.045 172.665 78.275 173.565 ;
        RECT 78.905 173.275 79.235 174.415 ;
        RECT 79.405 173.785 79.760 174.245 ;
        RECT 79.930 173.955 80.505 174.415 ;
        RECT 80.675 173.785 81.005 174.245 ;
        RECT 79.405 173.615 81.005 173.785 ;
        RECT 81.205 173.615 81.460 174.415 ;
        RECT 79.405 173.275 79.680 173.615 ;
        RECT 79.860 173.055 80.050 173.435 ;
        RECT 78.905 172.855 80.050 173.055 ;
        RECT 80.230 172.685 80.510 173.615 ;
        RECT 81.630 173.445 81.930 173.640 ;
        RECT 80.680 173.275 81.930 173.445 ;
        RECT 80.680 172.855 81.010 173.275 ;
        RECT 81.240 172.775 81.585 173.105 ;
        RECT 77.670 172.035 78.275 172.665 ;
        RECT 78.905 172.475 80.015 172.685 ;
        RECT 78.905 172.035 79.255 172.475 ;
        RECT 79.425 171.865 79.595 172.305 ;
        RECT 79.765 172.245 80.015 172.475 ;
        RECT 80.185 172.585 80.510 172.685 ;
        RECT 80.185 172.415 80.515 172.585 ;
        RECT 80.685 172.245 80.960 172.685 ;
        RECT 81.760 172.620 81.930 173.275 ;
        RECT 82.585 173.250 82.875 174.415 ;
        RECT 83.045 173.275 83.375 174.415 ;
        RECT 83.545 173.785 83.900 174.245 ;
        RECT 84.070 173.955 84.645 174.415 ;
        RECT 84.815 173.785 85.145 174.245 ;
        RECT 83.545 173.615 85.145 173.785 ;
        RECT 85.345 173.615 85.600 174.415 ;
        RECT 83.545 173.275 83.820 173.615 ;
        RECT 84.000 173.055 84.190 173.435 ;
        RECT 83.045 172.885 84.195 173.055 ;
        RECT 83.045 172.855 84.190 172.885 ;
        RECT 84.370 172.685 84.650 173.615 ;
        RECT 85.770 173.445 86.070 173.640 ;
        RECT 84.820 173.275 86.070 173.445 ;
        RECT 86.355 173.485 86.525 174.245 ;
        RECT 86.740 173.655 87.070 174.415 ;
        RECT 86.355 173.315 87.070 173.485 ;
        RECT 87.240 173.340 87.495 174.245 ;
        RECT 84.820 172.855 85.150 173.275 ;
        RECT 85.380 172.775 85.725 173.105 ;
        RECT 79.765 172.035 80.960 172.245 ;
        RECT 81.195 171.865 81.525 172.605 ;
        RECT 81.695 172.290 81.930 172.620 ;
        RECT 82.585 171.865 82.875 172.590 ;
        RECT 83.045 172.475 84.155 172.685 ;
        RECT 83.045 172.035 83.395 172.475 ;
        RECT 83.565 171.865 83.735 172.305 ;
        RECT 83.905 172.245 84.155 172.475 ;
        RECT 84.325 172.585 84.650 172.685 ;
        RECT 84.325 172.415 84.655 172.585 ;
        RECT 84.825 172.245 85.100 172.685 ;
        RECT 85.900 172.620 86.070 173.275 ;
        RECT 86.265 172.765 86.620 173.135 ;
        RECT 86.900 173.105 87.070 173.315 ;
        RECT 86.900 172.775 87.155 173.105 ;
        RECT 83.905 172.035 85.100 172.245 ;
        RECT 85.335 171.865 85.665 172.605 ;
        RECT 85.835 172.290 86.070 172.620 ;
        RECT 86.900 172.585 87.070 172.775 ;
        RECT 87.325 172.610 87.495 173.340 ;
        RECT 87.670 173.265 87.930 174.415 ;
        RECT 88.105 173.325 89.315 174.415 ;
        RECT 88.105 172.785 88.625 173.325 ;
        RECT 86.355 172.415 87.070 172.585 ;
        RECT 86.355 172.035 86.525 172.415 ;
        RECT 86.740 171.865 87.070 172.245 ;
        RECT 87.240 172.035 87.495 172.610 ;
        RECT 87.670 171.865 87.930 172.705 ;
        RECT 88.795 172.615 89.315 173.155 ;
        RECT 88.105 171.865 89.315 172.615 ;
        RECT 18.100 171.695 89.400 171.865 ;
        RECT 18.185 170.945 19.395 171.695 ;
        RECT 18.185 170.405 18.705 170.945 ;
        RECT 19.565 170.925 21.235 171.695 ;
        RECT 21.870 170.955 22.125 171.525 ;
        RECT 22.295 171.295 22.625 171.695 ;
        RECT 23.050 171.160 23.580 171.525 ;
        RECT 23.770 171.355 24.045 171.525 ;
        RECT 23.765 171.185 24.045 171.355 ;
        RECT 23.050 171.125 23.225 171.160 ;
        RECT 22.295 170.955 23.225 171.125 ;
        RECT 18.875 170.235 19.395 170.775 ;
        RECT 19.565 170.405 20.315 170.925 ;
        RECT 20.485 170.235 21.235 170.755 ;
        RECT 18.185 169.145 19.395 170.235 ;
        RECT 19.565 169.145 21.235 170.235 ;
        RECT 21.870 170.285 22.040 170.955 ;
        RECT 22.295 170.785 22.465 170.955 ;
        RECT 22.210 170.455 22.465 170.785 ;
        RECT 22.690 170.455 22.885 170.785 ;
        RECT 21.870 169.315 22.205 170.285 ;
        RECT 22.375 169.145 22.545 170.285 ;
        RECT 22.715 169.485 22.885 170.455 ;
        RECT 23.055 169.825 23.225 170.955 ;
        RECT 23.395 170.165 23.565 170.965 ;
        RECT 23.770 170.365 24.045 171.185 ;
        RECT 24.215 170.165 24.405 171.525 ;
        RECT 24.585 171.160 25.095 171.695 ;
        RECT 25.315 170.885 25.560 171.490 ;
        RECT 26.005 170.925 28.595 171.695 ;
        RECT 28.775 170.965 29.075 171.695 ;
        RECT 24.605 170.715 25.835 170.885 ;
        RECT 23.395 169.995 24.405 170.165 ;
        RECT 24.575 170.150 25.325 170.340 ;
        RECT 23.055 169.655 24.180 169.825 ;
        RECT 24.575 169.485 24.745 170.150 ;
        RECT 25.495 169.905 25.835 170.715 ;
        RECT 26.005 170.405 27.215 170.925 ;
        RECT 29.255 170.785 29.485 171.405 ;
        RECT 29.685 171.135 29.910 171.515 ;
        RECT 30.080 171.305 30.410 171.695 ;
        RECT 29.685 170.955 30.015 171.135 ;
        RECT 27.385 170.235 28.595 170.755 ;
        RECT 28.780 170.455 29.075 170.785 ;
        RECT 29.255 170.455 29.670 170.785 ;
        RECT 29.840 170.285 30.015 170.955 ;
        RECT 30.185 170.455 30.425 171.105 ;
        RECT 30.640 170.955 31.255 171.525 ;
        RECT 31.425 171.185 31.640 171.695 ;
        RECT 31.870 171.185 32.150 171.515 ;
        RECT 32.330 171.185 32.570 171.695 ;
        RECT 22.715 169.315 24.745 169.485 ;
        RECT 24.915 169.145 25.085 169.905 ;
        RECT 25.320 169.495 25.835 169.905 ;
        RECT 26.005 169.145 28.595 170.235 ;
        RECT 28.775 169.925 29.670 170.255 ;
        RECT 29.840 170.095 30.425 170.285 ;
        RECT 28.775 169.755 29.980 169.925 ;
        RECT 28.775 169.325 29.105 169.755 ;
        RECT 29.285 169.145 29.480 169.585 ;
        RECT 29.650 169.325 29.980 169.755 ;
        RECT 30.150 169.325 30.425 170.095 ;
        RECT 30.640 169.935 30.955 170.955 ;
        RECT 31.125 170.285 31.295 170.785 ;
        RECT 31.545 170.455 31.810 171.015 ;
        RECT 31.980 170.285 32.150 171.185 ;
        RECT 32.905 171.085 33.245 171.500 ;
        RECT 33.415 171.255 33.585 171.695 ;
        RECT 33.755 171.305 35.005 171.485 ;
        RECT 33.755 171.085 34.085 171.305 ;
        RECT 35.275 171.235 35.445 171.695 ;
        RECT 32.320 170.455 32.675 171.015 ;
        RECT 32.905 170.915 34.085 171.085 ;
        RECT 34.255 171.065 34.620 171.135 ;
        RECT 34.255 170.885 35.505 171.065 ;
        RECT 32.905 170.505 33.370 170.705 ;
        RECT 33.545 170.455 33.875 170.705 ;
        RECT 34.045 170.675 34.510 170.705 ;
        RECT 34.045 170.505 34.515 170.675 ;
        RECT 34.045 170.455 34.510 170.505 ;
        RECT 34.705 170.455 35.060 170.705 ;
        RECT 33.545 170.335 33.725 170.455 ;
        RECT 31.125 170.115 32.550 170.285 ;
        RECT 30.640 169.315 31.175 169.935 ;
        RECT 31.345 169.145 31.675 169.945 ;
        RECT 32.160 169.940 32.550 170.115 ;
        RECT 32.905 169.145 33.225 170.325 ;
        RECT 33.395 170.165 33.725 170.335 ;
        RECT 35.230 170.285 35.505 170.885 ;
        RECT 33.395 169.375 33.595 170.165 ;
        RECT 33.895 170.075 35.505 170.285 ;
        RECT 33.895 169.975 34.305 170.075 ;
        RECT 33.920 169.315 34.305 169.975 ;
        RECT 34.700 169.145 35.485 169.905 ;
        RECT 35.675 169.315 35.955 171.415 ;
        RECT 37.050 170.955 37.305 171.525 ;
        RECT 37.475 171.295 37.805 171.695 ;
        RECT 38.230 171.160 38.760 171.525 ;
        RECT 38.230 171.125 38.405 171.160 ;
        RECT 37.475 170.955 38.405 171.125 ;
        RECT 37.050 170.285 37.220 170.955 ;
        RECT 37.475 170.785 37.645 170.955 ;
        RECT 37.390 170.455 37.645 170.785 ;
        RECT 37.870 170.455 38.065 170.785 ;
        RECT 37.050 169.315 37.385 170.285 ;
        RECT 37.555 169.145 37.725 170.285 ;
        RECT 37.895 169.485 38.065 170.455 ;
        RECT 38.235 169.825 38.405 170.955 ;
        RECT 38.575 170.165 38.745 170.965 ;
        RECT 38.950 170.675 39.225 171.525 ;
        RECT 38.945 170.505 39.225 170.675 ;
        RECT 38.950 170.365 39.225 170.505 ;
        RECT 39.395 170.165 39.585 171.525 ;
        RECT 39.765 171.160 40.275 171.695 ;
        RECT 40.495 170.885 40.740 171.490 ;
        RECT 41.185 170.925 43.775 171.695 ;
        RECT 43.945 170.970 44.235 171.695 ;
        RECT 44.415 170.965 44.715 171.695 ;
        RECT 39.785 170.715 41.015 170.885 ;
        RECT 38.575 169.995 39.585 170.165 ;
        RECT 39.755 170.150 40.505 170.340 ;
        RECT 38.235 169.655 39.360 169.825 ;
        RECT 39.755 169.485 39.925 170.150 ;
        RECT 40.675 169.905 41.015 170.715 ;
        RECT 41.185 170.405 42.395 170.925 ;
        RECT 44.895 170.785 45.125 171.405 ;
        RECT 45.325 171.135 45.550 171.515 ;
        RECT 45.720 171.305 46.050 171.695 ;
        RECT 45.325 170.955 45.655 171.135 ;
        RECT 42.565 170.235 43.775 170.755 ;
        RECT 44.420 170.455 44.715 170.785 ;
        RECT 44.895 170.455 45.310 170.785 ;
        RECT 37.895 169.315 39.925 169.485 ;
        RECT 40.095 169.145 40.265 169.905 ;
        RECT 40.500 169.495 41.015 169.905 ;
        RECT 41.185 169.145 43.775 170.235 ;
        RECT 43.945 169.145 44.235 170.310 ;
        RECT 45.480 170.285 45.655 170.955 ;
        RECT 45.825 170.455 46.065 171.105 ;
        RECT 44.415 169.925 45.310 170.255 ;
        RECT 45.480 170.095 46.065 170.285 ;
        RECT 44.415 169.755 45.620 169.925 ;
        RECT 44.415 169.325 44.745 169.755 ;
        RECT 44.925 169.145 45.120 169.585 ;
        RECT 45.290 169.325 45.620 169.755 ;
        RECT 45.790 169.325 46.065 170.095 ;
        RECT 46.715 169.325 46.975 171.515 ;
        RECT 47.235 171.325 47.905 171.695 ;
        RECT 48.085 171.145 48.395 171.515 ;
        RECT 47.165 170.945 48.395 171.145 ;
        RECT 47.165 170.275 47.455 170.945 ;
        RECT 48.575 170.765 48.805 171.405 ;
        RECT 48.985 170.965 49.275 171.695 ;
        RECT 49.465 170.925 52.055 171.695 ;
        RECT 52.250 171.305 52.580 171.695 ;
        RECT 52.750 171.135 52.975 171.515 ;
        RECT 47.635 170.455 48.100 170.765 ;
        RECT 48.280 170.455 48.805 170.765 ;
        RECT 48.985 170.455 49.285 170.785 ;
        RECT 49.465 170.405 50.675 170.925 ;
        RECT 47.165 170.055 47.935 170.275 ;
        RECT 47.145 169.145 47.485 169.875 ;
        RECT 47.665 169.325 47.935 170.055 ;
        RECT 48.115 170.035 49.275 170.275 ;
        RECT 50.845 170.235 52.055 170.755 ;
        RECT 52.235 170.455 52.475 171.105 ;
        RECT 52.645 170.955 52.975 171.135 ;
        RECT 52.645 170.285 52.820 170.955 ;
        RECT 53.175 170.785 53.405 171.405 ;
        RECT 53.585 170.965 53.885 171.695 ;
        RECT 55.010 171.305 55.340 171.695 ;
        RECT 55.510 171.135 55.735 171.515 ;
        RECT 52.990 170.455 53.405 170.785 ;
        RECT 53.585 170.455 53.880 170.785 ;
        RECT 54.995 170.455 55.235 171.105 ;
        RECT 55.405 170.955 55.735 171.135 ;
        RECT 55.405 170.285 55.580 170.955 ;
        RECT 55.935 170.785 56.165 171.405 ;
        RECT 56.345 170.965 56.645 171.695 ;
        RECT 57.745 171.020 58.005 171.525 ;
        RECT 58.185 171.315 58.515 171.695 ;
        RECT 58.695 171.145 58.865 171.525 ;
        RECT 55.750 170.455 56.165 170.785 ;
        RECT 56.345 170.455 56.640 170.785 ;
        RECT 48.115 169.325 48.345 170.035 ;
        RECT 48.515 169.145 48.845 169.855 ;
        RECT 49.015 169.325 49.275 170.035 ;
        RECT 49.465 169.145 52.055 170.235 ;
        RECT 52.235 170.095 52.820 170.285 ;
        RECT 52.235 169.325 52.510 170.095 ;
        RECT 52.990 169.925 53.885 170.255 ;
        RECT 52.680 169.755 53.885 169.925 ;
        RECT 52.680 169.325 53.010 169.755 ;
        RECT 53.180 169.145 53.375 169.585 ;
        RECT 53.555 169.325 53.885 169.755 ;
        RECT 54.995 170.095 55.580 170.285 ;
        RECT 54.995 169.325 55.270 170.095 ;
        RECT 55.750 169.925 56.645 170.255 ;
        RECT 55.440 169.755 56.645 169.925 ;
        RECT 55.440 169.325 55.770 169.755 ;
        RECT 55.940 169.145 56.135 169.585 ;
        RECT 56.315 169.325 56.645 169.755 ;
        RECT 57.745 170.220 57.925 171.020 ;
        RECT 58.200 170.975 58.865 171.145 ;
        RECT 58.200 170.720 58.370 170.975 ;
        RECT 58.095 170.390 58.370 170.720 ;
        RECT 58.595 170.425 58.935 170.795 ;
        RECT 58.200 170.245 58.370 170.390 ;
        RECT 57.745 169.315 58.015 170.220 ;
        RECT 58.200 170.075 58.875 170.245 ;
        RECT 58.185 169.145 58.515 169.905 ;
        RECT 58.695 169.315 58.875 170.075 ;
        RECT 59.140 169.325 59.420 171.515 ;
        RECT 59.620 171.325 60.350 171.695 ;
        RECT 60.930 171.155 61.360 171.515 ;
        RECT 59.620 170.965 61.360 171.155 ;
        RECT 59.620 170.455 59.880 170.965 ;
        RECT 59.610 169.145 59.895 170.285 ;
        RECT 60.090 170.165 60.350 170.785 ;
        RECT 60.545 170.165 60.970 170.785 ;
        RECT 61.140 170.735 61.360 170.965 ;
        RECT 61.530 170.915 61.775 171.695 ;
        RECT 61.140 170.435 61.685 170.735 ;
        RECT 61.975 170.615 62.205 171.515 ;
        RECT 60.160 169.795 61.185 169.995 ;
        RECT 60.160 169.325 60.330 169.795 ;
        RECT 60.505 169.145 60.835 169.625 ;
        RECT 61.005 169.325 61.185 169.795 ;
        RECT 61.355 169.325 61.685 170.435 ;
        RECT 61.865 169.935 62.205 170.615 ;
        RECT 62.385 170.115 62.615 171.455 ;
        RECT 62.895 171.145 63.065 171.525 ;
        RECT 63.245 171.315 63.575 171.695 ;
        RECT 62.895 170.975 63.560 171.145 ;
        RECT 63.755 171.020 64.015 171.525 ;
        RECT 62.825 170.425 63.155 170.795 ;
        RECT 63.390 170.720 63.560 170.975 ;
        RECT 63.390 170.390 63.675 170.720 ;
        RECT 63.390 170.245 63.560 170.390 ;
        RECT 62.895 170.075 63.560 170.245 ;
        RECT 63.845 170.220 64.015 171.020 ;
        RECT 61.865 169.735 62.615 169.935 ;
        RECT 61.855 169.145 62.205 169.555 ;
        RECT 62.375 169.345 62.615 169.735 ;
        RECT 62.895 169.315 63.065 170.075 ;
        RECT 63.245 169.145 63.575 169.905 ;
        RECT 63.745 169.315 64.015 170.220 ;
        RECT 64.185 171.020 64.445 171.525 ;
        RECT 64.625 171.315 64.955 171.695 ;
        RECT 65.135 171.145 65.305 171.525 ;
        RECT 64.185 170.220 64.355 171.020 ;
        RECT 64.640 170.975 65.305 171.145 ;
        RECT 65.655 171.145 65.825 171.525 ;
        RECT 66.005 171.315 66.335 171.695 ;
        RECT 65.655 170.975 66.320 171.145 ;
        RECT 66.515 171.020 66.775 171.525 ;
        RECT 64.640 170.720 64.810 170.975 ;
        RECT 64.525 170.390 64.810 170.720 ;
        RECT 65.045 170.425 65.375 170.795 ;
        RECT 65.585 170.425 65.925 170.795 ;
        RECT 66.150 170.720 66.320 170.975 ;
        RECT 64.640 170.245 64.810 170.390 ;
        RECT 66.150 170.390 66.425 170.720 ;
        RECT 66.150 170.245 66.320 170.390 ;
        RECT 64.185 169.315 64.455 170.220 ;
        RECT 64.640 170.075 65.305 170.245 ;
        RECT 64.625 169.145 64.955 169.905 ;
        RECT 65.135 169.315 65.305 170.075 ;
        RECT 65.645 170.075 66.320 170.245 ;
        RECT 66.595 170.220 66.775 171.020 ;
        RECT 65.645 169.315 65.825 170.075 ;
        RECT 66.005 169.145 66.335 169.905 ;
        RECT 66.505 169.315 66.775 170.220 ;
        RECT 66.945 171.020 67.205 171.525 ;
        RECT 67.385 171.315 67.715 171.695 ;
        RECT 67.895 171.145 68.065 171.525 ;
        RECT 66.945 170.220 67.125 171.020 ;
        RECT 67.400 170.975 68.065 171.145 ;
        RECT 68.415 171.145 68.585 171.525 ;
        RECT 68.765 171.315 69.095 171.695 ;
        RECT 68.415 170.975 69.080 171.145 ;
        RECT 69.275 171.020 69.535 171.525 ;
        RECT 67.400 170.720 67.570 170.975 ;
        RECT 67.295 170.390 67.570 170.720 ;
        RECT 67.795 170.425 68.135 170.795 ;
        RECT 68.345 170.425 68.675 170.795 ;
        RECT 68.910 170.720 69.080 170.975 ;
        RECT 67.400 170.245 67.570 170.390 ;
        RECT 68.910 170.390 69.195 170.720 ;
        RECT 68.910 170.245 69.080 170.390 ;
        RECT 66.945 169.315 67.215 170.220 ;
        RECT 67.400 170.075 68.075 170.245 ;
        RECT 67.385 169.145 67.715 169.905 ;
        RECT 67.895 169.315 68.075 170.075 ;
        RECT 68.415 170.075 69.080 170.245 ;
        RECT 69.365 170.220 69.535 171.020 ;
        RECT 69.705 170.970 69.995 171.695 ;
        RECT 70.715 171.145 70.885 171.525 ;
        RECT 71.065 171.315 71.395 171.695 ;
        RECT 70.715 170.975 71.380 171.145 ;
        RECT 71.575 171.020 71.835 171.525 ;
        RECT 70.645 170.425 70.985 170.795 ;
        RECT 71.210 170.720 71.380 170.975 ;
        RECT 71.210 170.390 71.485 170.720 ;
        RECT 68.415 169.315 68.585 170.075 ;
        RECT 68.765 169.145 69.095 169.905 ;
        RECT 69.265 169.315 69.535 170.220 ;
        RECT 69.705 169.145 69.995 170.310 ;
        RECT 71.210 170.245 71.380 170.390 ;
        RECT 70.705 170.075 71.380 170.245 ;
        RECT 71.655 170.220 71.835 171.020 ;
        RECT 72.065 170.875 72.275 171.695 ;
        RECT 72.445 170.895 72.775 171.525 ;
        RECT 72.445 170.295 72.695 170.895 ;
        RECT 72.945 170.875 73.175 171.695 ;
        RECT 73.540 171.045 73.870 171.510 ;
        RECT 74.040 171.225 74.210 171.695 ;
        RECT 74.380 171.045 74.710 171.525 ;
        RECT 73.540 170.875 74.710 171.045 ;
        RECT 72.865 170.455 73.195 170.705 ;
        RECT 73.385 170.495 74.030 170.705 ;
        RECT 74.200 170.495 74.770 170.705 ;
        RECT 74.940 170.325 75.110 171.525 ;
        RECT 75.650 171.125 75.820 171.330 ;
        RECT 70.705 169.315 70.885 170.075 ;
        RECT 71.065 169.145 71.395 169.905 ;
        RECT 71.565 169.315 71.835 170.220 ;
        RECT 72.065 169.145 72.275 170.285 ;
        RECT 72.445 169.315 72.775 170.295 ;
        RECT 72.945 169.145 73.175 170.285 ;
        RECT 73.600 169.145 73.930 170.245 ;
        RECT 74.405 169.915 75.110 170.325 ;
        RECT 75.280 170.955 75.820 171.125 ;
        RECT 76.100 170.955 76.270 171.695 ;
        RECT 76.535 170.955 76.895 171.330 ;
        RECT 77.155 171.145 77.325 171.525 ;
        RECT 77.540 171.315 77.870 171.695 ;
        RECT 77.155 170.975 77.870 171.145 ;
        RECT 75.280 170.255 75.450 170.955 ;
        RECT 75.620 170.455 75.950 170.785 ;
        RECT 76.120 170.455 76.470 170.785 ;
        RECT 75.280 170.085 75.905 170.255 ;
        RECT 76.120 169.915 76.385 170.455 ;
        RECT 76.640 170.300 76.895 170.955 ;
        RECT 77.065 170.425 77.420 170.795 ;
        RECT 77.700 170.785 77.870 170.975 ;
        RECT 78.040 170.950 78.295 171.525 ;
        RECT 77.700 170.455 77.955 170.785 ;
        RECT 74.405 169.745 76.385 169.915 ;
        RECT 74.405 169.315 74.730 169.745 ;
        RECT 74.900 169.145 75.230 169.565 ;
        RECT 75.975 169.145 76.385 169.575 ;
        RECT 76.555 169.315 76.895 170.300 ;
        RECT 77.700 170.245 77.870 170.455 ;
        RECT 77.155 170.075 77.870 170.245 ;
        RECT 78.125 170.220 78.295 170.950 ;
        RECT 78.470 170.855 78.730 171.695 ;
        RECT 78.905 171.185 79.210 171.695 ;
        RECT 78.905 170.455 79.220 171.015 ;
        RECT 79.390 170.705 79.640 171.515 ;
        RECT 79.810 171.170 80.070 171.695 ;
        RECT 80.250 170.705 80.500 171.515 ;
        RECT 80.670 171.135 80.930 171.695 ;
        RECT 81.100 171.045 81.360 171.500 ;
        RECT 81.530 171.215 81.790 171.695 ;
        RECT 81.960 171.045 82.220 171.500 ;
        RECT 82.390 171.215 82.650 171.695 ;
        RECT 82.820 171.045 83.080 171.500 ;
        RECT 83.250 171.215 83.495 171.695 ;
        RECT 83.665 171.045 83.940 171.500 ;
        RECT 84.110 171.215 84.355 171.695 ;
        RECT 84.525 171.045 84.785 171.500 ;
        RECT 84.965 171.215 85.215 171.695 ;
        RECT 85.385 171.045 85.645 171.500 ;
        RECT 85.825 171.215 86.075 171.695 ;
        RECT 86.245 171.045 86.505 171.500 ;
        RECT 86.685 171.215 86.945 171.695 ;
        RECT 87.115 171.045 87.375 171.500 ;
        RECT 87.545 171.215 87.845 171.695 ;
        RECT 81.100 170.875 87.845 171.045 ;
        RECT 88.105 170.945 89.315 171.695 ;
        RECT 79.390 170.455 86.510 170.705 ;
        RECT 77.155 169.315 77.325 170.075 ;
        RECT 77.540 169.145 77.870 169.905 ;
        RECT 78.040 169.315 78.295 170.220 ;
        RECT 78.470 169.145 78.730 170.295 ;
        RECT 78.915 169.145 79.210 169.955 ;
        RECT 79.390 169.315 79.635 170.455 ;
        RECT 79.810 169.145 80.070 169.955 ;
        RECT 80.250 169.320 80.500 170.455 ;
        RECT 86.680 170.285 87.845 170.875 ;
        RECT 81.100 170.060 87.845 170.285 ;
        RECT 88.105 170.235 88.625 170.775 ;
        RECT 88.795 170.405 89.315 170.945 ;
        RECT 81.100 170.045 86.505 170.060 ;
        RECT 80.670 169.150 80.930 169.945 ;
        RECT 81.100 169.320 81.360 170.045 ;
        RECT 81.530 169.150 81.790 169.875 ;
        RECT 81.960 169.320 82.220 170.045 ;
        RECT 82.390 169.150 82.650 169.875 ;
        RECT 82.820 169.320 83.080 170.045 ;
        RECT 83.250 169.150 83.510 169.875 ;
        RECT 83.680 169.320 83.940 170.045 ;
        RECT 84.110 169.150 84.355 169.875 ;
        RECT 84.525 169.320 84.785 170.045 ;
        RECT 84.970 169.150 85.215 169.875 ;
        RECT 85.385 169.320 85.645 170.045 ;
        RECT 85.830 169.150 86.075 169.875 ;
        RECT 86.245 169.320 86.505 170.045 ;
        RECT 86.690 169.150 86.945 169.875 ;
        RECT 87.115 169.320 87.405 170.060 ;
        RECT 80.670 169.145 86.945 169.150 ;
        RECT 87.575 169.145 87.845 169.890 ;
        RECT 88.105 169.145 89.315 170.235 ;
        RECT 18.100 168.975 89.400 169.145 ;
        RECT 18.185 167.885 19.395 168.975 ;
        RECT 19.565 167.885 21.235 168.975 ;
        RECT 18.185 167.175 18.705 167.715 ;
        RECT 18.875 167.345 19.395 167.885 ;
        RECT 19.565 167.195 20.315 167.715 ;
        RECT 20.485 167.365 21.235 167.885 ;
        RECT 21.410 167.835 21.745 168.805 ;
        RECT 21.915 167.835 22.085 168.975 ;
        RECT 22.255 168.635 24.285 168.805 ;
        RECT 18.185 166.425 19.395 167.175 ;
        RECT 19.565 166.425 21.235 167.195 ;
        RECT 21.410 167.165 21.580 167.835 ;
        RECT 22.255 167.665 22.425 168.635 ;
        RECT 21.750 167.335 22.005 167.665 ;
        RECT 22.230 167.335 22.425 167.665 ;
        RECT 22.595 168.295 23.720 168.465 ;
        RECT 21.835 167.165 22.005 167.335 ;
        RECT 22.595 167.165 22.765 168.295 ;
        RECT 21.410 166.595 21.665 167.165 ;
        RECT 21.835 166.995 22.765 167.165 ;
        RECT 22.935 167.955 23.945 168.125 ;
        RECT 22.935 167.155 23.105 167.955 ;
        RECT 22.590 166.960 22.765 166.995 ;
        RECT 21.835 166.425 22.165 166.825 ;
        RECT 22.590 166.595 23.120 166.960 ;
        RECT 23.310 166.935 23.585 167.755 ;
        RECT 23.305 166.765 23.585 166.935 ;
        RECT 23.310 166.595 23.585 166.765 ;
        RECT 23.755 166.595 23.945 167.955 ;
        RECT 24.115 167.970 24.285 168.635 ;
        RECT 24.455 168.215 24.625 168.975 ;
        RECT 24.860 168.215 25.375 168.625 ;
        RECT 24.115 167.780 24.865 167.970 ;
        RECT 25.035 167.405 25.375 168.215 ;
        RECT 25.545 167.885 28.135 168.975 ;
        RECT 24.145 167.235 25.375 167.405 ;
        RECT 24.125 166.425 24.635 166.960 ;
        RECT 24.855 166.630 25.100 167.235 ;
        RECT 25.545 167.195 26.755 167.715 ;
        RECT 26.925 167.365 28.135 167.885 ;
        RECT 28.315 168.365 28.645 168.795 ;
        RECT 28.825 168.535 29.020 168.975 ;
        RECT 29.190 168.365 29.520 168.795 ;
        RECT 28.315 168.195 29.520 168.365 ;
        RECT 28.315 167.865 29.210 168.195 ;
        RECT 29.690 168.025 29.965 168.795 ;
        RECT 29.380 167.835 29.965 168.025 ;
        RECT 28.320 167.335 28.615 167.665 ;
        RECT 28.795 167.335 29.210 167.665 ;
        RECT 25.545 166.425 28.135 167.195 ;
        RECT 28.315 166.425 28.615 167.155 ;
        RECT 28.795 166.715 29.025 167.335 ;
        RECT 29.380 167.165 29.555 167.835 ;
        RECT 31.065 167.810 31.355 168.975 ;
        RECT 31.560 168.185 32.095 168.805 ;
        RECT 29.225 166.985 29.555 167.165 ;
        RECT 29.725 167.015 29.965 167.665 ;
        RECT 31.560 167.165 31.875 168.185 ;
        RECT 32.265 168.175 32.595 168.975 ;
        RECT 33.835 168.365 34.165 168.795 ;
        RECT 34.345 168.535 34.540 168.975 ;
        RECT 34.710 168.365 35.040 168.795 ;
        RECT 33.835 168.195 35.040 168.365 ;
        RECT 33.080 168.005 33.470 168.180 ;
        RECT 32.045 167.835 33.470 168.005 ;
        RECT 33.835 167.865 34.730 168.195 ;
        RECT 35.210 168.025 35.485 168.795 ;
        RECT 34.900 167.835 35.485 168.025 ;
        RECT 36.590 167.835 36.925 168.805 ;
        RECT 37.095 167.835 37.265 168.975 ;
        RECT 37.435 168.635 39.465 168.805 ;
        RECT 32.045 167.335 32.215 167.835 ;
        RECT 29.225 166.605 29.450 166.985 ;
        RECT 29.620 166.425 29.950 166.815 ;
        RECT 31.065 166.425 31.355 167.150 ;
        RECT 31.560 166.595 32.175 167.165 ;
        RECT 32.465 167.105 32.730 167.665 ;
        RECT 32.900 166.935 33.070 167.835 ;
        RECT 33.240 167.105 33.595 167.665 ;
        RECT 33.840 167.335 34.135 167.665 ;
        RECT 34.315 167.335 34.730 167.665 ;
        RECT 32.345 166.425 32.560 166.935 ;
        RECT 32.790 166.605 33.070 166.935 ;
        RECT 33.250 166.425 33.490 166.935 ;
        RECT 33.835 166.425 34.135 167.155 ;
        RECT 34.315 166.715 34.545 167.335 ;
        RECT 34.900 167.165 35.075 167.835 ;
        RECT 34.745 166.985 35.075 167.165 ;
        RECT 35.245 167.015 35.485 167.665 ;
        RECT 36.590 167.165 36.760 167.835 ;
        RECT 37.435 167.665 37.605 168.635 ;
        RECT 36.930 167.335 37.185 167.665 ;
        RECT 37.410 167.335 37.605 167.665 ;
        RECT 37.775 168.295 38.900 168.465 ;
        RECT 37.015 167.165 37.185 167.335 ;
        RECT 37.775 167.165 37.945 168.295 ;
        RECT 34.745 166.605 34.970 166.985 ;
        RECT 35.140 166.425 35.470 166.815 ;
        RECT 36.590 166.595 36.845 167.165 ;
        RECT 37.015 166.995 37.945 167.165 ;
        RECT 38.115 167.955 39.125 168.125 ;
        RECT 38.115 167.155 38.285 167.955 ;
        RECT 37.770 166.960 37.945 166.995 ;
        RECT 37.015 166.425 37.345 166.825 ;
        RECT 37.770 166.595 38.300 166.960 ;
        RECT 38.490 166.935 38.765 167.755 ;
        RECT 38.485 166.765 38.765 166.935 ;
        RECT 38.490 166.595 38.765 166.765 ;
        RECT 38.935 166.595 39.125 167.955 ;
        RECT 39.295 167.970 39.465 168.635 ;
        RECT 39.635 168.215 39.805 168.975 ;
        RECT 40.040 168.215 40.555 168.625 ;
        RECT 39.295 167.780 40.045 167.970 ;
        RECT 40.215 167.405 40.555 168.215 ;
        RECT 40.765 167.835 40.995 168.975 ;
        RECT 41.165 167.825 41.495 168.805 ;
        RECT 41.665 167.835 41.875 168.975 ;
        RECT 42.105 167.835 42.365 168.975 ;
        RECT 42.535 167.825 42.865 168.805 ;
        RECT 43.035 167.835 43.315 168.975 ;
        RECT 44.415 168.365 44.745 168.795 ;
        RECT 44.925 168.535 45.120 168.975 ;
        RECT 45.290 168.365 45.620 168.795 ;
        RECT 44.415 168.195 45.620 168.365 ;
        RECT 44.415 167.865 45.310 168.195 ;
        RECT 45.790 168.025 46.065 168.795 ;
        RECT 45.480 167.835 46.065 168.025 ;
        RECT 46.285 167.835 46.515 168.975 ;
        RECT 40.745 167.415 41.075 167.665 ;
        RECT 39.325 167.235 40.555 167.405 ;
        RECT 39.305 166.425 39.815 166.960 ;
        RECT 40.035 166.630 40.280 167.235 ;
        RECT 40.765 166.425 40.995 167.245 ;
        RECT 41.245 167.225 41.495 167.825 ;
        RECT 42.125 167.415 42.460 167.665 ;
        RECT 41.165 166.595 41.495 167.225 ;
        RECT 41.665 166.425 41.875 167.245 ;
        RECT 42.630 167.225 42.800 167.825 ;
        RECT 42.970 167.395 43.305 167.665 ;
        RECT 44.420 167.335 44.715 167.665 ;
        RECT 44.895 167.335 45.310 167.665 ;
        RECT 42.105 166.595 42.800 167.225 ;
        RECT 43.005 166.425 43.315 167.225 ;
        RECT 44.415 166.425 44.715 167.155 ;
        RECT 44.895 166.715 45.125 167.335 ;
        RECT 45.480 167.165 45.655 167.835 ;
        RECT 46.685 167.825 47.015 168.805 ;
        RECT 47.185 167.835 47.395 168.975 ;
        RECT 47.625 167.885 48.835 168.975 ;
        RECT 45.325 166.985 45.655 167.165 ;
        RECT 45.825 167.015 46.065 167.665 ;
        RECT 46.265 167.415 46.595 167.665 ;
        RECT 45.325 166.605 45.550 166.985 ;
        RECT 45.720 166.425 46.050 166.815 ;
        RECT 46.285 166.425 46.515 167.245 ;
        RECT 46.765 167.225 47.015 167.825 ;
        RECT 46.685 166.595 47.015 167.225 ;
        RECT 47.185 166.425 47.395 167.245 ;
        RECT 47.625 167.175 48.145 167.715 ;
        RECT 48.315 167.345 48.835 167.885 ;
        RECT 49.005 167.835 49.265 168.975 ;
        RECT 49.435 167.825 49.765 168.805 ;
        RECT 49.935 167.835 50.215 168.975 ;
        RECT 50.385 168.540 55.730 168.975 ;
        RECT 49.025 167.415 49.360 167.665 ;
        RECT 49.530 167.225 49.700 167.825 ;
        RECT 49.870 167.395 50.205 167.665 ;
        RECT 47.625 166.425 48.835 167.175 ;
        RECT 49.005 166.595 49.700 167.225 ;
        RECT 49.905 166.425 50.215 167.225 ;
        RECT 51.970 166.970 52.310 167.800 ;
        RECT 53.790 167.290 54.140 168.540 ;
        RECT 56.825 167.810 57.115 168.975 ;
        RECT 57.285 167.835 57.560 168.805 ;
        RECT 57.770 168.175 58.050 168.975 ;
        RECT 58.220 168.465 59.835 168.795 ;
        RECT 58.220 168.125 59.395 168.295 ;
        RECT 58.220 168.005 58.390 168.125 ;
        RECT 57.730 167.835 58.390 168.005 ;
        RECT 50.385 166.425 55.730 166.970 ;
        RECT 56.825 166.425 57.115 167.150 ;
        RECT 57.285 167.100 57.455 167.835 ;
        RECT 57.730 167.665 57.900 167.835 ;
        RECT 58.650 167.665 58.895 167.955 ;
        RECT 59.065 167.835 59.395 168.125 ;
        RECT 59.655 167.665 59.825 168.225 ;
        RECT 60.075 167.835 60.335 168.975 ;
        RECT 60.505 167.885 62.175 168.975 ;
        RECT 57.625 167.335 57.900 167.665 ;
        RECT 58.070 167.335 58.895 167.665 ;
        RECT 59.110 167.335 59.825 167.665 ;
        RECT 59.995 167.415 60.330 167.665 ;
        RECT 57.730 167.165 57.900 167.335 ;
        RECT 59.575 167.245 59.825 167.335 ;
        RECT 57.285 166.755 57.560 167.100 ;
        RECT 57.730 166.995 59.395 167.165 ;
        RECT 57.750 166.425 58.125 166.825 ;
        RECT 58.295 166.645 58.465 166.995 ;
        RECT 58.635 166.425 58.965 166.825 ;
        RECT 59.135 166.595 59.395 166.995 ;
        RECT 59.575 166.825 59.905 167.245 ;
        RECT 60.075 166.425 60.335 167.245 ;
        RECT 60.505 167.195 61.255 167.715 ;
        RECT 61.425 167.365 62.175 167.885 ;
        RECT 62.810 168.025 63.075 168.795 ;
        RECT 63.245 168.255 63.575 168.975 ;
        RECT 63.765 168.435 64.025 168.795 ;
        RECT 64.195 168.605 64.525 168.975 ;
        RECT 64.695 168.435 64.955 168.795 ;
        RECT 63.765 168.205 64.955 168.435 ;
        RECT 65.525 168.025 65.815 168.795 ;
        RECT 60.505 166.425 62.175 167.195 ;
        RECT 62.810 166.605 63.145 168.025 ;
        RECT 63.320 167.845 65.815 168.025 ;
        RECT 66.045 168.135 66.300 168.805 ;
        RECT 66.470 168.215 66.800 168.975 ;
        RECT 66.970 168.375 67.220 168.805 ;
        RECT 67.390 168.555 67.745 168.975 ;
        RECT 67.935 168.635 69.105 168.805 ;
        RECT 67.935 168.595 68.265 168.635 ;
        RECT 68.375 168.375 68.605 168.465 ;
        RECT 66.970 168.135 68.605 168.375 ;
        RECT 68.775 168.135 69.105 168.635 ;
        RECT 66.045 168.125 66.255 168.135 ;
        RECT 63.320 167.155 63.545 167.845 ;
        RECT 63.745 167.335 64.025 167.665 ;
        RECT 64.205 167.335 64.780 167.665 ;
        RECT 64.960 167.335 65.395 167.665 ;
        RECT 65.575 167.335 65.845 167.665 ;
        RECT 63.320 166.965 65.805 167.155 ;
        RECT 63.325 166.425 64.070 166.795 ;
        RECT 64.635 166.605 64.890 166.965 ;
        RECT 65.070 166.425 65.400 166.795 ;
        RECT 65.580 166.605 65.805 166.965 ;
        RECT 66.045 167.005 66.215 168.125 ;
        RECT 69.275 167.965 69.445 168.805 ;
        RECT 66.385 167.795 69.445 167.965 ;
        RECT 69.715 168.365 70.045 168.795 ;
        RECT 70.225 168.535 70.420 168.975 ;
        RECT 70.590 168.365 70.920 168.795 ;
        RECT 69.715 168.195 70.920 168.365 ;
        RECT 69.715 167.865 70.610 168.195 ;
        RECT 71.090 168.025 71.365 168.795 ;
        RECT 72.475 168.175 72.805 168.975 ;
        RECT 72.985 168.635 74.415 168.805 ;
        RECT 70.780 167.835 71.365 168.025 ;
        RECT 72.985 168.005 73.235 168.635 ;
        RECT 72.465 167.835 73.235 168.005 ;
        RECT 66.385 167.245 66.555 167.795 ;
        RECT 66.785 167.415 67.150 167.615 ;
        RECT 67.320 167.415 67.650 167.615 ;
        RECT 66.385 167.075 67.185 167.245 ;
        RECT 66.045 166.925 66.230 167.005 ;
        RECT 66.045 166.595 66.300 166.925 ;
        RECT 66.515 166.425 66.845 166.905 ;
        RECT 67.015 166.845 67.185 167.075 ;
        RECT 67.365 167.015 67.650 167.415 ;
        RECT 67.920 167.415 68.395 167.615 ;
        RECT 68.565 167.415 69.010 167.615 ;
        RECT 69.180 167.415 69.530 167.625 ;
        RECT 67.920 167.015 68.200 167.415 ;
        RECT 69.720 167.335 70.015 167.665 ;
        RECT 70.195 167.335 70.610 167.665 ;
        RECT 68.380 167.075 69.445 167.245 ;
        RECT 68.380 166.845 68.550 167.075 ;
        RECT 67.015 166.595 68.550 166.845 ;
        RECT 68.775 166.425 69.105 166.905 ;
        RECT 69.275 166.595 69.445 167.075 ;
        RECT 69.715 166.425 70.015 167.155 ;
        RECT 70.195 166.715 70.425 167.335 ;
        RECT 70.780 167.165 70.955 167.835 ;
        RECT 70.625 166.985 70.955 167.165 ;
        RECT 71.125 167.015 71.365 167.665 ;
        RECT 72.465 167.165 72.635 167.835 ;
        RECT 72.805 167.335 73.210 167.665 ;
        RECT 73.425 167.335 73.675 168.465 ;
        RECT 73.875 167.665 74.075 168.465 ;
        RECT 74.245 167.955 74.415 168.635 ;
        RECT 74.585 168.125 74.900 168.975 ;
        RECT 75.075 168.175 75.515 168.805 ;
        RECT 74.245 167.785 75.035 167.955 ;
        RECT 73.875 167.335 74.120 167.665 ;
        RECT 74.305 167.335 74.695 167.615 ;
        RECT 74.865 167.335 75.035 167.785 ;
        RECT 75.205 167.165 75.515 168.175 ;
        RECT 76.675 168.005 77.035 168.180 ;
        RECT 77.620 168.175 77.790 168.975 ;
        RECT 77.960 168.345 78.290 168.805 ;
        RECT 78.460 168.515 78.630 168.975 ;
        RECT 77.960 168.175 78.735 168.345 ;
        RECT 76.675 167.835 78.135 168.005 ;
        RECT 76.670 167.615 76.865 167.665 ;
        RECT 76.665 167.445 76.865 167.615 ;
        RECT 70.625 166.605 70.850 166.985 ;
        RECT 71.020 166.425 71.350 166.815 ;
        RECT 72.465 166.595 72.955 167.165 ;
        RECT 73.125 166.995 74.285 167.165 ;
        RECT 73.125 166.595 73.355 166.995 ;
        RECT 73.525 166.425 73.945 166.825 ;
        RECT 74.115 166.595 74.285 166.995 ;
        RECT 74.455 166.425 74.905 167.165 ;
        RECT 75.075 166.605 75.515 167.165 ;
        RECT 76.670 167.105 76.865 167.445 ;
        RECT 77.035 166.935 77.215 167.835 ;
        RECT 77.385 167.105 77.795 167.665 ;
        RECT 77.965 167.335 78.135 167.835 ;
        RECT 78.305 167.165 78.735 168.175 ;
        RECT 78.960 168.105 79.245 168.975 ;
        RECT 79.415 168.345 79.675 168.805 ;
        RECT 79.850 168.515 80.105 168.975 ;
        RECT 80.275 168.345 80.535 168.805 ;
        RECT 79.415 168.175 80.535 168.345 ;
        RECT 80.705 168.175 81.015 168.975 ;
        RECT 79.415 167.925 79.675 168.175 ;
        RECT 81.185 168.005 81.495 168.805 ;
        RECT 78.040 166.995 78.735 167.165 ;
        RECT 78.920 167.755 79.675 167.925 ;
        RECT 80.465 167.835 81.495 168.005 ;
        RECT 78.920 167.245 79.325 167.755 ;
        RECT 80.465 167.585 80.635 167.835 ;
        RECT 79.495 167.415 80.635 167.585 ;
        RECT 78.920 167.075 80.570 167.245 ;
        RECT 80.805 167.095 81.155 167.665 ;
        RECT 76.625 166.425 76.865 166.935 ;
        RECT 77.035 166.595 77.325 166.935 ;
        RECT 77.555 166.425 77.870 166.935 ;
        RECT 78.040 166.725 78.210 166.995 ;
        RECT 78.380 166.425 78.710 166.825 ;
        RECT 78.965 166.425 79.245 166.905 ;
        RECT 79.415 166.685 79.675 167.075 ;
        RECT 79.850 166.425 80.105 166.905 ;
        RECT 80.275 166.685 80.570 167.075 ;
        RECT 81.325 166.925 81.495 167.835 ;
        RECT 82.585 167.810 82.875 168.975 ;
        RECT 83.085 168.635 84.225 168.805 ;
        RECT 83.085 168.175 83.385 168.635 ;
        RECT 83.555 168.005 83.885 168.465 ;
        RECT 83.125 167.955 83.885 168.005 ;
        RECT 83.105 167.785 83.885 167.955 ;
        RECT 84.055 168.005 84.225 168.635 ;
        RECT 84.395 168.175 84.725 168.975 ;
        RECT 84.895 168.005 85.170 168.805 ;
        RECT 84.055 167.795 85.170 168.005 ;
        RECT 85.345 168.005 85.655 168.805 ;
        RECT 85.825 168.175 86.135 168.975 ;
        RECT 86.305 168.345 86.565 168.805 ;
        RECT 86.735 168.515 86.990 168.975 ;
        RECT 87.165 168.345 87.425 168.805 ;
        RECT 86.305 168.175 87.425 168.345 ;
        RECT 85.345 167.835 86.375 168.005 ;
        RECT 83.125 167.245 83.340 167.785 ;
        RECT 83.510 167.415 84.280 167.615 ;
        RECT 84.450 167.415 85.170 167.615 ;
        RECT 80.750 166.425 81.025 166.905 ;
        RECT 81.195 166.595 81.495 166.925 ;
        RECT 82.585 166.425 82.875 167.150 ;
        RECT 83.125 167.075 84.725 167.245 ;
        RECT 83.555 167.065 84.725 167.075 ;
        RECT 83.095 166.425 83.385 166.895 ;
        RECT 83.555 166.595 83.885 167.065 ;
        RECT 84.055 166.425 84.225 166.895 ;
        RECT 84.395 166.595 84.725 167.065 ;
        RECT 84.895 166.425 85.170 167.245 ;
        RECT 85.345 166.925 85.515 167.835 ;
        RECT 85.685 167.095 86.035 167.665 ;
        RECT 86.205 167.585 86.375 167.835 ;
        RECT 87.165 167.925 87.425 168.175 ;
        RECT 87.595 168.105 87.880 168.975 ;
        RECT 87.165 167.755 87.920 167.925 ;
        RECT 86.205 167.415 87.345 167.585 ;
        RECT 87.515 167.245 87.920 167.755 ;
        RECT 88.105 167.885 89.315 168.975 ;
        RECT 88.105 167.345 88.625 167.885 ;
        RECT 86.270 167.075 87.920 167.245 ;
        RECT 88.795 167.175 89.315 167.715 ;
        RECT 85.345 166.595 85.645 166.925 ;
        RECT 85.815 166.425 86.090 166.905 ;
        RECT 86.270 166.685 86.565 167.075 ;
        RECT 86.735 166.425 86.990 166.905 ;
        RECT 87.165 166.685 87.425 167.075 ;
        RECT 87.595 166.425 87.875 166.905 ;
        RECT 88.105 166.425 89.315 167.175 ;
        RECT 18.100 166.255 89.400 166.425 ;
        RECT 18.185 165.505 19.395 166.255 ;
        RECT 18.185 164.965 18.705 165.505 ;
        RECT 19.565 165.485 22.155 166.255 ;
        RECT 18.875 164.795 19.395 165.335 ;
        RECT 19.565 164.965 20.775 165.485 ;
        RECT 22.600 165.445 22.845 166.050 ;
        RECT 23.065 165.720 23.575 166.255 ;
        RECT 20.945 164.795 22.155 165.315 ;
        RECT 18.185 163.705 19.395 164.795 ;
        RECT 19.565 163.705 22.155 164.795 ;
        RECT 22.325 165.275 23.555 165.445 ;
        RECT 22.325 164.465 22.665 165.275 ;
        RECT 22.835 164.710 23.585 164.900 ;
        RECT 22.325 164.055 22.840 164.465 ;
        RECT 23.075 163.705 23.245 164.465 ;
        RECT 23.415 164.045 23.585 164.710 ;
        RECT 23.755 164.725 23.945 166.085 ;
        RECT 24.115 165.235 24.390 166.085 ;
        RECT 24.580 165.720 25.110 166.085 ;
        RECT 25.535 165.855 25.865 166.255 ;
        RECT 24.935 165.685 25.110 165.720 ;
        RECT 24.115 165.065 24.395 165.235 ;
        RECT 24.115 164.925 24.390 165.065 ;
        RECT 24.595 164.725 24.765 165.525 ;
        RECT 23.755 164.555 24.765 164.725 ;
        RECT 24.935 165.515 25.865 165.685 ;
        RECT 26.035 165.515 26.290 166.085 ;
        RECT 24.935 164.385 25.105 165.515 ;
        RECT 25.695 165.345 25.865 165.515 ;
        RECT 23.980 164.215 25.105 164.385 ;
        RECT 25.275 165.015 25.470 165.345 ;
        RECT 25.695 165.015 25.950 165.345 ;
        RECT 25.275 164.045 25.445 165.015 ;
        RECT 26.120 164.845 26.290 165.515 ;
        RECT 26.465 165.645 26.805 166.060 ;
        RECT 26.975 165.815 27.145 166.255 ;
        RECT 27.315 165.865 28.565 166.045 ;
        RECT 27.315 165.645 27.645 165.865 ;
        RECT 28.835 165.795 29.005 166.255 ;
        RECT 26.465 165.475 27.645 165.645 ;
        RECT 27.815 165.625 28.180 165.695 ;
        RECT 27.815 165.445 29.065 165.625 ;
        RECT 26.465 165.065 26.930 165.265 ;
        RECT 27.105 165.015 27.435 165.265 ;
        RECT 27.605 165.235 28.070 165.265 ;
        RECT 27.605 165.065 28.075 165.235 ;
        RECT 27.605 165.015 28.070 165.065 ;
        RECT 28.265 165.015 28.620 165.265 ;
        RECT 27.105 164.895 27.285 165.015 ;
        RECT 23.415 163.875 25.445 164.045 ;
        RECT 25.615 163.705 25.785 164.845 ;
        RECT 25.955 163.875 26.290 164.845 ;
        RECT 26.465 163.705 26.785 164.885 ;
        RECT 26.955 164.725 27.285 164.895 ;
        RECT 28.790 164.845 29.065 165.445 ;
        RECT 26.955 163.935 27.155 164.725 ;
        RECT 27.455 164.635 29.065 164.845 ;
        RECT 27.455 164.535 27.865 164.635 ;
        RECT 27.480 163.875 27.865 164.535 ;
        RECT 28.260 163.705 29.045 164.465 ;
        RECT 29.235 163.875 29.515 165.975 ;
        RECT 29.685 165.710 35.030 166.255 ;
        RECT 35.205 165.710 40.550 166.255 ;
        RECT 31.270 164.880 31.610 165.710 ;
        RECT 33.090 164.140 33.440 165.390 ;
        RECT 36.790 164.880 37.130 165.710 ;
        RECT 40.725 165.485 43.315 166.255 ;
        RECT 43.945 165.530 44.235 166.255 ;
        RECT 44.405 165.485 46.995 166.255 ;
        RECT 47.625 165.515 47.965 166.085 ;
        RECT 48.160 165.590 48.330 166.255 ;
        RECT 48.610 165.915 48.830 165.960 ;
        RECT 48.605 165.745 48.830 165.915 ;
        RECT 49.000 165.775 49.445 165.945 ;
        RECT 48.610 165.605 48.830 165.745 ;
        RECT 38.610 164.140 38.960 165.390 ;
        RECT 40.725 164.965 41.935 165.485 ;
        RECT 42.105 164.795 43.315 165.315 ;
        RECT 44.405 164.965 45.615 165.485 ;
        RECT 29.685 163.705 35.030 164.140 ;
        RECT 35.205 163.705 40.550 164.140 ;
        RECT 40.725 163.705 43.315 164.795 ;
        RECT 43.945 163.705 44.235 164.870 ;
        RECT 45.785 164.795 46.995 165.315 ;
        RECT 44.405 163.705 46.995 164.795 ;
        RECT 47.625 164.545 47.800 165.515 ;
        RECT 48.610 165.435 49.105 165.605 ;
        RECT 47.970 164.895 48.140 165.345 ;
        RECT 48.310 165.065 48.760 165.265 ;
        RECT 48.930 165.240 49.105 165.435 ;
        RECT 49.275 164.985 49.445 165.775 ;
        RECT 49.615 165.650 49.865 166.020 ;
        RECT 49.695 165.265 49.865 165.650 ;
        RECT 50.035 165.615 50.285 166.020 ;
        RECT 50.455 165.785 50.625 166.255 ;
        RECT 50.795 165.615 51.135 166.020 ;
        RECT 50.035 165.435 51.135 165.615 ;
        RECT 51.305 165.485 52.975 166.255 ;
        RECT 53.155 165.530 53.485 166.040 ;
        RECT 53.655 165.855 53.985 166.255 ;
        RECT 55.035 165.685 55.365 166.025 ;
        RECT 55.535 165.855 55.865 166.255 ;
        RECT 49.695 165.095 49.890 165.265 ;
        RECT 47.970 164.725 48.365 164.895 ;
        RECT 49.275 164.845 49.550 164.985 ;
        RECT 47.625 163.875 47.885 164.545 ;
        RECT 48.195 164.455 48.365 164.725 ;
        RECT 48.535 164.625 49.550 164.845 ;
        RECT 49.720 164.845 49.890 165.095 ;
        RECT 50.060 165.015 50.620 165.265 ;
        RECT 49.720 164.455 50.275 164.845 ;
        RECT 48.195 164.285 50.275 164.455 ;
        RECT 48.055 163.705 48.385 164.105 ;
        RECT 49.255 163.705 49.655 164.105 ;
        RECT 49.945 164.050 50.275 164.285 ;
        RECT 50.445 163.915 50.620 165.015 ;
        RECT 50.790 164.695 51.135 165.265 ;
        RECT 51.305 164.965 52.055 165.485 ;
        RECT 52.225 164.795 52.975 165.315 ;
        RECT 50.790 163.705 51.135 164.525 ;
        RECT 51.305 163.705 52.975 164.795 ;
        RECT 53.155 164.765 53.345 165.530 ;
        RECT 53.655 165.515 56.020 165.685 ;
        RECT 53.655 165.345 53.825 165.515 ;
        RECT 53.515 165.015 53.825 165.345 ;
        RECT 53.995 165.015 54.300 165.345 ;
        RECT 53.155 163.915 53.485 164.765 ;
        RECT 53.655 163.705 53.905 164.845 ;
        RECT 54.085 164.685 54.300 165.015 ;
        RECT 54.475 164.685 54.760 165.345 ;
        RECT 54.955 164.685 55.220 165.345 ;
        RECT 55.435 164.685 55.680 165.345 ;
        RECT 55.850 164.515 56.020 165.515 ;
        RECT 56.570 165.475 57.070 166.085 ;
        RECT 56.365 165.015 56.715 165.265 ;
        RECT 56.900 164.845 57.070 165.475 ;
        RECT 57.700 165.605 58.030 166.085 ;
        RECT 58.200 165.795 58.425 166.255 ;
        RECT 58.595 165.605 58.925 166.085 ;
        RECT 57.700 165.435 58.925 165.605 ;
        RECT 59.115 165.455 59.365 166.255 ;
        RECT 59.535 165.455 59.875 166.085 ;
        RECT 60.210 165.745 60.450 166.255 ;
        RECT 60.630 165.745 60.910 166.075 ;
        RECT 61.140 165.745 61.355 166.255 ;
        RECT 57.240 165.065 57.570 165.265 ;
        RECT 57.740 165.065 58.070 165.265 ;
        RECT 58.240 165.065 58.660 165.265 ;
        RECT 58.835 165.095 59.530 165.265 ;
        RECT 58.835 164.845 59.005 165.095 ;
        RECT 59.700 164.845 59.875 165.455 ;
        RECT 60.105 165.015 60.460 165.575 ;
        RECT 60.630 164.845 60.800 165.745 ;
        RECT 60.970 165.015 61.235 165.575 ;
        RECT 61.525 165.515 62.140 166.085 ;
        RECT 61.485 164.845 61.655 165.345 ;
        RECT 54.095 164.345 55.385 164.515 ;
        RECT 54.095 163.925 54.345 164.345 ;
        RECT 54.575 163.705 54.905 164.175 ;
        RECT 55.135 163.925 55.385 164.345 ;
        RECT 55.565 164.345 56.020 164.515 ;
        RECT 56.570 164.675 59.005 164.845 ;
        RECT 55.565 163.915 55.895 164.345 ;
        RECT 56.570 163.875 56.900 164.675 ;
        RECT 57.070 163.705 57.400 164.505 ;
        RECT 57.700 163.875 58.030 164.675 ;
        RECT 58.675 163.705 58.925 164.505 ;
        RECT 59.195 163.705 59.365 164.845 ;
        RECT 59.535 163.875 59.875 164.845 ;
        RECT 60.230 164.675 61.655 164.845 ;
        RECT 60.230 164.500 60.620 164.675 ;
        RECT 61.105 163.705 61.435 164.505 ;
        RECT 61.825 164.495 62.140 165.515 ;
        RECT 62.345 165.455 63.040 166.085 ;
        RECT 63.245 165.455 63.555 166.255 ;
        RECT 63.725 165.485 66.315 166.255 ;
        RECT 66.510 165.865 66.840 166.255 ;
        RECT 67.010 165.695 67.235 166.075 ;
        RECT 62.365 165.015 62.700 165.265 ;
        RECT 62.870 164.895 63.040 165.455 ;
        RECT 63.210 165.015 63.545 165.285 ;
        RECT 63.725 164.965 64.935 165.485 ;
        RECT 62.865 164.855 63.040 164.895 ;
        RECT 61.605 163.875 62.140 164.495 ;
        RECT 62.345 163.705 62.605 164.845 ;
        RECT 62.775 163.875 63.105 164.855 ;
        RECT 63.275 163.705 63.555 164.845 ;
        RECT 65.105 164.795 66.315 165.315 ;
        RECT 66.495 165.015 66.735 165.665 ;
        RECT 66.905 165.515 67.235 165.695 ;
        RECT 66.905 164.845 67.080 165.515 ;
        RECT 67.435 165.345 67.665 165.965 ;
        RECT 67.845 165.525 68.145 166.255 ;
        RECT 68.415 165.705 68.585 166.085 ;
        RECT 68.765 165.875 69.095 166.255 ;
        RECT 68.415 165.535 69.080 165.705 ;
        RECT 69.275 165.580 69.535 166.085 ;
        RECT 67.250 165.015 67.665 165.345 ;
        RECT 67.845 165.015 68.140 165.345 ;
        RECT 68.345 164.985 68.685 165.355 ;
        RECT 68.910 165.280 69.080 165.535 ;
        RECT 63.725 163.705 66.315 164.795 ;
        RECT 66.495 164.655 67.080 164.845 ;
        RECT 68.910 164.950 69.185 165.280 ;
        RECT 66.495 163.885 66.770 164.655 ;
        RECT 67.250 164.485 68.145 164.815 ;
        RECT 68.910 164.805 69.080 164.950 ;
        RECT 66.940 164.315 68.145 164.485 ;
        RECT 66.940 163.885 67.270 164.315 ;
        RECT 67.440 163.705 67.635 164.145 ;
        RECT 67.815 163.885 68.145 164.315 ;
        RECT 68.405 164.635 69.080 164.805 ;
        RECT 69.355 164.780 69.535 165.580 ;
        RECT 69.705 165.530 69.995 166.255 ;
        RECT 71.175 165.705 71.345 166.085 ;
        RECT 71.525 165.875 71.855 166.255 ;
        RECT 71.175 165.535 71.840 165.705 ;
        RECT 72.035 165.580 72.295 166.085 ;
        RECT 71.105 164.985 71.435 165.355 ;
        RECT 71.670 165.280 71.840 165.535 ;
        RECT 71.670 164.950 71.955 165.280 ;
        RECT 68.405 163.875 68.585 164.635 ;
        RECT 68.765 163.705 69.095 164.465 ;
        RECT 69.265 163.875 69.535 164.780 ;
        RECT 69.705 163.705 69.995 164.870 ;
        RECT 71.670 164.805 71.840 164.950 ;
        RECT 71.175 164.635 71.840 164.805 ;
        RECT 72.125 164.780 72.295 165.580 ;
        RECT 72.555 165.705 72.725 166.085 ;
        RECT 72.905 165.875 73.235 166.255 ;
        RECT 72.555 165.535 73.220 165.705 ;
        RECT 73.415 165.580 73.675 166.085 ;
        RECT 72.485 164.985 72.815 165.355 ;
        RECT 73.050 165.280 73.220 165.535 ;
        RECT 73.050 164.950 73.335 165.280 ;
        RECT 73.050 164.805 73.220 164.950 ;
        RECT 71.175 163.875 71.345 164.635 ;
        RECT 71.525 163.705 71.855 164.465 ;
        RECT 72.025 163.875 72.295 164.780 ;
        RECT 72.555 164.635 73.220 164.805 ;
        RECT 73.505 164.780 73.675 165.580 ;
        RECT 72.555 163.875 72.725 164.635 ;
        RECT 72.905 163.705 73.235 164.465 ;
        RECT 73.405 163.875 73.675 164.780 ;
        RECT 73.845 165.515 74.205 165.890 ;
        RECT 74.470 165.515 74.640 166.255 ;
        RECT 74.920 165.685 75.090 165.890 ;
        RECT 74.920 165.515 75.460 165.685 ;
        RECT 73.845 164.860 74.100 165.515 ;
        RECT 74.270 165.015 74.620 165.345 ;
        RECT 74.790 165.015 75.120 165.345 ;
        RECT 73.845 163.875 74.185 164.860 ;
        RECT 74.355 164.475 74.620 165.015 ;
        RECT 75.290 164.815 75.460 165.515 ;
        RECT 74.835 164.645 75.460 164.815 ;
        RECT 75.630 164.885 75.800 166.085 ;
        RECT 76.030 165.605 76.360 166.085 ;
        RECT 76.530 165.785 76.700 166.255 ;
        RECT 76.870 165.605 77.200 166.070 ;
        RECT 76.030 165.435 77.200 165.605 ;
        RECT 77.540 165.685 77.795 166.035 ;
        RECT 77.965 165.855 78.295 166.255 ;
        RECT 78.465 165.685 78.635 166.035 ;
        RECT 78.805 165.855 79.185 166.255 ;
        RECT 77.540 165.515 79.205 165.685 ;
        RECT 79.375 165.580 79.650 165.925 ;
        RECT 80.750 165.750 81.085 166.255 ;
        RECT 81.255 165.685 81.495 166.060 ;
        RECT 81.775 165.925 81.945 166.070 ;
        RECT 81.775 165.730 82.150 165.925 ;
        RECT 82.510 165.760 82.905 166.255 ;
        RECT 79.035 165.345 79.205 165.515 ;
        RECT 75.970 165.055 76.540 165.265 ;
        RECT 76.710 165.055 77.355 165.265 ;
        RECT 77.525 165.015 77.870 165.345 ;
        RECT 78.040 165.015 78.865 165.345 ;
        RECT 79.035 165.015 79.310 165.345 ;
        RECT 75.630 164.475 76.335 164.885 ;
        RECT 74.355 164.305 76.335 164.475 ;
        RECT 74.355 163.705 74.765 164.135 ;
        RECT 75.510 163.705 75.840 164.125 ;
        RECT 76.010 163.875 76.335 164.305 ;
        RECT 76.810 163.705 77.140 164.805 ;
        RECT 77.545 164.555 77.870 164.845 ;
        RECT 78.040 164.725 78.235 165.015 ;
        RECT 79.035 164.845 79.205 165.015 ;
        RECT 79.480 164.845 79.650 165.580 ;
        RECT 78.545 164.675 79.205 164.845 ;
        RECT 78.545 164.555 78.715 164.675 ;
        RECT 77.545 164.385 78.715 164.555 ;
        RECT 77.525 163.925 78.715 164.215 ;
        RECT 78.885 163.705 79.165 164.505 ;
        RECT 79.375 163.875 79.650 164.845 ;
        RECT 80.805 164.725 81.105 165.575 ;
        RECT 81.275 165.535 81.495 165.685 ;
        RECT 81.275 165.205 81.810 165.535 ;
        RECT 81.980 165.395 82.150 165.730 ;
        RECT 83.075 165.565 83.315 166.085 ;
        RECT 83.505 165.595 83.780 166.255 ;
        RECT 83.950 165.625 84.200 166.085 ;
        RECT 84.375 165.760 84.705 166.255 ;
        RECT 81.275 164.555 81.510 165.205 ;
        RECT 81.980 165.035 82.965 165.395 ;
        RECT 80.835 164.325 81.510 164.555 ;
        RECT 81.680 165.015 82.965 165.035 ;
        RECT 81.680 164.865 82.540 165.015 ;
        RECT 80.835 163.895 81.005 164.325 ;
        RECT 81.175 163.705 81.505 164.155 ;
        RECT 81.680 163.920 81.965 164.865 ;
        RECT 83.140 164.760 83.315 165.565 ;
        RECT 83.950 165.415 84.120 165.625 ;
        RECT 84.885 165.590 85.115 166.035 ;
        RECT 83.505 164.895 84.120 165.415 ;
        RECT 84.290 164.915 84.520 165.345 ;
        RECT 84.705 165.095 85.115 165.590 ;
        RECT 85.285 165.770 86.075 166.035 ;
        RECT 85.285 164.915 85.540 165.770 ;
        RECT 86.355 165.705 86.525 166.085 ;
        RECT 86.740 165.875 87.070 166.255 ;
        RECT 85.710 165.095 86.095 165.575 ;
        RECT 86.355 165.535 87.070 165.705 ;
        RECT 86.265 164.985 86.620 165.355 ;
        RECT 86.900 165.345 87.070 165.535 ;
        RECT 87.240 165.510 87.495 166.085 ;
        RECT 86.900 165.015 87.155 165.345 ;
        RECT 82.140 164.385 82.835 164.695 ;
        RECT 82.145 163.705 82.830 164.175 ;
        RECT 83.010 163.975 83.315 164.760 ;
        RECT 83.505 163.705 83.765 164.715 ;
        RECT 83.935 164.545 84.105 164.895 ;
        RECT 84.290 164.745 86.080 164.915 ;
        RECT 86.900 164.805 87.070 165.015 ;
        RECT 83.935 163.875 84.210 164.545 ;
        RECT 84.410 163.705 84.625 164.550 ;
        RECT 84.850 164.450 85.100 164.745 ;
        RECT 85.325 164.385 85.655 164.575 ;
        RECT 84.810 163.875 85.285 164.215 ;
        RECT 85.465 164.210 85.655 164.385 ;
        RECT 85.825 164.380 86.080 164.745 ;
        RECT 86.355 164.635 87.070 164.805 ;
        RECT 87.325 164.780 87.495 165.510 ;
        RECT 87.670 165.415 87.930 166.255 ;
        RECT 88.105 165.505 89.315 166.255 ;
        RECT 85.465 163.705 86.095 164.210 ;
        RECT 86.355 163.875 86.525 164.635 ;
        RECT 86.740 163.705 87.070 164.465 ;
        RECT 87.240 163.875 87.495 164.780 ;
        RECT 87.670 163.705 87.930 164.855 ;
        RECT 88.105 164.795 88.625 165.335 ;
        RECT 88.795 164.965 89.315 165.505 ;
        RECT 88.105 163.705 89.315 164.795 ;
        RECT 18.100 163.535 89.400 163.705 ;
        RECT 18.185 162.445 19.395 163.535 ;
        RECT 19.565 162.445 22.155 163.535 ;
        RECT 18.185 161.735 18.705 162.275 ;
        RECT 18.875 161.905 19.395 162.445 ;
        RECT 19.565 161.755 20.775 162.275 ;
        RECT 20.945 161.925 22.155 162.445 ;
        RECT 22.325 162.775 22.840 163.185 ;
        RECT 23.075 162.775 23.245 163.535 ;
        RECT 23.415 163.195 25.445 163.365 ;
        RECT 22.325 161.965 22.665 162.775 ;
        RECT 23.415 162.530 23.585 163.195 ;
        RECT 23.980 162.855 25.105 163.025 ;
        RECT 22.835 162.340 23.585 162.530 ;
        RECT 23.755 162.515 24.765 162.685 ;
        RECT 22.325 161.795 23.555 161.965 ;
        RECT 18.185 160.985 19.395 161.735 ;
        RECT 19.565 160.985 22.155 161.755 ;
        RECT 22.600 161.190 22.845 161.795 ;
        RECT 23.065 160.985 23.575 161.520 ;
        RECT 23.755 161.155 23.945 162.515 ;
        RECT 24.115 162.175 24.390 162.315 ;
        RECT 24.115 162.005 24.395 162.175 ;
        RECT 24.115 161.155 24.390 162.005 ;
        RECT 24.595 161.715 24.765 162.515 ;
        RECT 24.935 161.725 25.105 162.855 ;
        RECT 25.275 162.225 25.445 163.195 ;
        RECT 25.615 162.395 25.785 163.535 ;
        RECT 25.955 162.395 26.290 163.365 ;
        RECT 26.465 162.445 29.055 163.535 ;
        RECT 25.275 161.895 25.470 162.225 ;
        RECT 25.695 161.895 25.950 162.225 ;
        RECT 25.695 161.725 25.865 161.895 ;
        RECT 26.120 161.725 26.290 162.395 ;
        RECT 24.935 161.555 25.865 161.725 ;
        RECT 24.935 161.520 25.110 161.555 ;
        RECT 24.580 161.155 25.110 161.520 ;
        RECT 25.535 160.985 25.865 161.385 ;
        RECT 26.035 161.155 26.290 161.725 ;
        RECT 26.465 161.755 27.675 162.275 ;
        RECT 27.845 161.925 29.055 162.445 ;
        RECT 29.685 162.395 29.945 163.535 ;
        RECT 30.115 162.385 30.445 163.365 ;
        RECT 30.615 162.395 30.895 163.535 ;
        RECT 29.705 161.975 30.040 162.225 ;
        RECT 30.210 161.785 30.380 162.385 ;
        RECT 31.065 162.370 31.355 163.535 ;
        RECT 31.525 162.355 31.845 163.535 ;
        RECT 32.015 162.515 32.215 163.305 ;
        RECT 32.540 162.705 32.925 163.365 ;
        RECT 33.320 162.775 34.105 163.535 ;
        RECT 32.515 162.605 32.925 162.705 ;
        RECT 32.015 162.345 32.345 162.515 ;
        RECT 32.515 162.395 34.125 162.605 ;
        RECT 32.165 162.225 32.345 162.345 ;
        RECT 30.550 161.955 30.885 162.225 ;
        RECT 31.525 161.975 31.990 162.175 ;
        RECT 32.165 161.975 32.495 162.225 ;
        RECT 32.665 162.175 33.130 162.225 ;
        RECT 32.665 162.005 33.135 162.175 ;
        RECT 32.665 161.975 33.130 162.005 ;
        RECT 33.325 161.975 33.680 162.225 ;
        RECT 33.850 161.795 34.125 162.395 ;
        RECT 26.465 160.985 29.055 161.755 ;
        RECT 29.685 161.155 30.380 161.785 ;
        RECT 30.585 160.985 30.895 161.785 ;
        RECT 31.065 160.985 31.355 161.710 ;
        RECT 31.525 161.595 32.705 161.765 ;
        RECT 31.525 161.180 31.865 161.595 ;
        RECT 32.035 160.985 32.205 161.425 ;
        RECT 32.375 161.375 32.705 161.595 ;
        RECT 32.875 161.615 34.125 161.795 ;
        RECT 32.875 161.545 33.240 161.615 ;
        RECT 32.375 161.195 33.625 161.375 ;
        RECT 33.895 160.985 34.065 161.445 ;
        RECT 34.295 161.265 34.575 163.365 ;
        RECT 35.210 162.395 35.545 163.365 ;
        RECT 35.715 162.395 35.885 163.535 ;
        RECT 36.055 163.195 38.085 163.365 ;
        RECT 35.210 161.725 35.380 162.395 ;
        RECT 36.055 162.225 36.225 163.195 ;
        RECT 35.550 161.895 35.805 162.225 ;
        RECT 36.030 161.895 36.225 162.225 ;
        RECT 36.395 162.855 37.520 163.025 ;
        RECT 35.635 161.725 35.805 161.895 ;
        RECT 36.395 161.725 36.565 162.855 ;
        RECT 35.210 161.155 35.465 161.725 ;
        RECT 35.635 161.555 36.565 161.725 ;
        RECT 36.735 162.515 37.745 162.685 ;
        RECT 36.735 161.715 36.905 162.515 ;
        RECT 36.390 161.520 36.565 161.555 ;
        RECT 35.635 160.985 35.965 161.385 ;
        RECT 36.390 161.155 36.920 161.520 ;
        RECT 37.110 161.495 37.385 162.315 ;
        RECT 37.105 161.325 37.385 161.495 ;
        RECT 37.110 161.155 37.385 161.325 ;
        RECT 37.555 161.155 37.745 162.515 ;
        RECT 37.915 162.530 38.085 163.195 ;
        RECT 38.255 162.775 38.425 163.535 ;
        RECT 38.660 162.775 39.175 163.185 ;
        RECT 37.915 162.340 38.665 162.530 ;
        RECT 38.835 161.965 39.175 162.775 ;
        RECT 39.345 162.395 39.605 163.535 ;
        RECT 39.775 162.385 40.105 163.365 ;
        RECT 40.275 162.395 40.555 163.535 ;
        RECT 40.725 162.445 43.315 163.535 ;
        RECT 39.365 161.975 39.700 162.225 ;
        RECT 37.945 161.795 39.175 161.965 ;
        RECT 37.925 160.985 38.435 161.520 ;
        RECT 38.655 161.190 38.900 161.795 ;
        RECT 39.870 161.785 40.040 162.385 ;
        RECT 40.210 161.955 40.545 162.225 ;
        RECT 39.345 161.155 40.040 161.785 ;
        RECT 40.245 160.985 40.555 161.785 ;
        RECT 40.725 161.755 41.935 162.275 ;
        RECT 42.105 161.925 43.315 162.445 ;
        RECT 43.490 162.585 43.755 163.355 ;
        RECT 43.925 162.815 44.255 163.535 ;
        RECT 44.445 162.995 44.705 163.355 ;
        RECT 44.875 163.165 45.205 163.535 ;
        RECT 45.375 162.995 45.635 163.355 ;
        RECT 44.445 162.765 45.635 162.995 ;
        RECT 46.205 162.585 46.495 163.355 ;
        RECT 46.705 163.100 52.050 163.535 ;
        RECT 40.725 160.985 43.315 161.755 ;
        RECT 43.490 161.165 43.825 162.585 ;
        RECT 44.000 162.405 46.495 162.585 ;
        RECT 44.000 161.715 44.225 162.405 ;
        RECT 44.425 161.895 44.705 162.225 ;
        RECT 44.885 161.895 45.460 162.225 ;
        RECT 45.640 161.895 46.075 162.225 ;
        RECT 46.255 161.895 46.525 162.225 ;
        RECT 44.000 161.525 46.485 161.715 ;
        RECT 48.290 161.530 48.630 162.360 ;
        RECT 50.110 161.850 50.460 163.100 ;
        RECT 52.225 162.445 55.735 163.535 ;
        RECT 52.225 161.755 53.875 162.275 ;
        RECT 54.045 161.925 55.735 162.445 ;
        RECT 56.825 162.370 57.115 163.535 ;
        RECT 57.285 162.395 57.560 163.365 ;
        RECT 57.770 162.735 58.050 163.535 ;
        RECT 58.220 163.025 59.835 163.355 ;
        RECT 58.220 162.685 59.395 162.855 ;
        RECT 58.220 162.565 58.390 162.685 ;
        RECT 57.730 162.395 58.390 162.565 ;
        RECT 44.005 160.985 44.750 161.355 ;
        RECT 45.315 161.165 45.570 161.525 ;
        RECT 45.750 160.985 46.080 161.355 ;
        RECT 46.260 161.165 46.485 161.525 ;
        RECT 46.705 160.985 52.050 161.530 ;
        RECT 52.225 160.985 55.735 161.755 ;
        RECT 56.825 160.985 57.115 161.710 ;
        RECT 57.285 161.660 57.455 162.395 ;
        RECT 57.730 162.225 57.900 162.395 ;
        RECT 58.650 162.225 58.895 162.515 ;
        RECT 59.065 162.395 59.395 162.685 ;
        RECT 59.655 162.225 59.825 162.785 ;
        RECT 60.075 162.395 60.335 163.535 ;
        RECT 60.505 163.100 65.850 163.535 ;
        RECT 57.625 161.895 57.900 162.225 ;
        RECT 58.070 161.895 58.895 162.225 ;
        RECT 59.110 161.895 59.825 162.225 ;
        RECT 59.995 161.975 60.330 162.225 ;
        RECT 57.730 161.725 57.900 161.895 ;
        RECT 59.575 161.805 59.825 161.895 ;
        RECT 57.285 161.315 57.560 161.660 ;
        RECT 57.730 161.555 59.395 161.725 ;
        RECT 57.750 160.985 58.125 161.385 ;
        RECT 58.295 161.205 58.465 161.555 ;
        RECT 58.635 160.985 58.965 161.385 ;
        RECT 59.135 161.155 59.395 161.555 ;
        RECT 59.575 161.385 59.905 161.805 ;
        RECT 60.075 160.985 60.335 161.805 ;
        RECT 62.090 161.530 62.430 162.360 ;
        RECT 63.910 161.850 64.260 163.100 ;
        RECT 66.025 162.445 69.535 163.535 ;
        RECT 69.705 162.445 70.915 163.535 ;
        RECT 66.025 161.755 67.675 162.275 ;
        RECT 67.845 161.925 69.535 162.445 ;
        RECT 60.505 160.985 65.850 161.530 ;
        RECT 66.025 160.985 69.535 161.755 ;
        RECT 69.705 161.735 70.225 162.275 ;
        RECT 70.395 161.905 70.915 162.445 ;
        RECT 69.705 160.985 70.915 161.735 ;
        RECT 71.085 161.155 71.835 163.365 ;
        RECT 72.005 162.980 72.610 163.535 ;
        RECT 72.785 163.025 73.265 163.365 ;
        RECT 73.435 162.990 73.690 163.535 ;
        RECT 72.005 162.880 72.620 162.980 ;
        RECT 72.435 162.855 72.620 162.880 ;
        RECT 72.005 162.260 72.265 162.710 ;
        RECT 72.435 162.610 72.765 162.855 ;
        RECT 72.935 162.535 73.690 162.785 ;
        RECT 73.860 162.665 74.135 163.365 ;
        RECT 72.920 162.500 73.690 162.535 ;
        RECT 72.905 162.490 73.690 162.500 ;
        RECT 72.900 162.475 73.795 162.490 ;
        RECT 72.880 162.460 73.795 162.475 ;
        RECT 72.860 162.450 73.795 162.460 ;
        RECT 72.835 162.440 73.795 162.450 ;
        RECT 72.765 162.410 73.795 162.440 ;
        RECT 72.745 162.380 73.795 162.410 ;
        RECT 72.725 162.350 73.795 162.380 ;
        RECT 72.695 162.325 73.795 162.350 ;
        RECT 72.660 162.290 73.795 162.325 ;
        RECT 72.630 162.285 73.795 162.290 ;
        RECT 72.630 162.280 73.020 162.285 ;
        RECT 72.630 162.270 72.995 162.280 ;
        RECT 72.630 162.265 72.980 162.270 ;
        RECT 72.630 162.260 72.965 162.265 ;
        RECT 72.005 162.255 72.965 162.260 ;
        RECT 72.005 162.245 72.955 162.255 ;
        RECT 72.005 162.240 72.945 162.245 ;
        RECT 72.005 162.230 72.935 162.240 ;
        RECT 72.005 162.220 72.930 162.230 ;
        RECT 72.005 162.215 72.925 162.220 ;
        RECT 72.005 162.200 72.915 162.215 ;
        RECT 72.005 162.185 72.910 162.200 ;
        RECT 72.005 162.160 72.900 162.185 ;
        RECT 72.005 162.090 72.895 162.160 ;
        RECT 72.005 161.535 72.555 161.920 ;
        RECT 72.725 161.365 72.895 162.090 ;
        RECT 72.005 161.195 72.895 161.365 ;
        RECT 73.065 161.690 73.395 162.115 ;
        RECT 73.565 161.890 73.795 162.285 ;
        RECT 73.065 161.205 73.285 161.690 ;
        RECT 73.965 161.635 74.135 162.665 ;
        RECT 74.315 162.395 74.645 163.535 ;
        RECT 75.175 162.565 75.505 163.350 ;
        RECT 74.825 162.395 75.505 162.565 ;
        RECT 76.225 162.605 76.405 163.365 ;
        RECT 76.585 162.775 76.915 163.535 ;
        RECT 76.225 162.435 76.900 162.605 ;
        RECT 77.085 162.460 77.355 163.365 ;
        RECT 77.525 163.025 78.715 163.315 ;
        RECT 74.305 161.975 74.655 162.225 ;
        RECT 74.825 161.795 74.995 162.395 ;
        RECT 76.730 162.290 76.900 162.435 ;
        RECT 75.165 161.975 75.515 162.225 ;
        RECT 76.165 161.885 76.505 162.255 ;
        RECT 76.730 161.960 77.005 162.290 ;
        RECT 73.455 160.985 73.705 161.525 ;
        RECT 73.875 161.155 74.135 161.635 ;
        RECT 74.315 160.985 74.585 161.795 ;
        RECT 74.755 161.155 75.085 161.795 ;
        RECT 75.255 160.985 75.495 161.795 ;
        RECT 76.730 161.705 76.900 161.960 ;
        RECT 76.235 161.535 76.900 161.705 ;
        RECT 77.175 161.660 77.355 162.460 ;
        RECT 77.545 162.685 78.715 162.855 ;
        RECT 78.885 162.735 79.165 163.535 ;
        RECT 77.545 162.395 77.870 162.685 ;
        RECT 78.545 162.565 78.715 162.685 ;
        RECT 78.040 162.225 78.235 162.515 ;
        RECT 78.545 162.395 79.205 162.565 ;
        RECT 79.375 162.395 79.650 163.365 ;
        RECT 80.325 163.195 81.465 163.365 ;
        RECT 80.325 162.735 80.625 163.195 ;
        RECT 80.795 162.565 81.125 163.025 ;
        RECT 80.365 162.515 81.125 162.565 ;
        RECT 79.035 162.225 79.205 162.395 ;
        RECT 77.525 161.895 77.870 162.225 ;
        RECT 78.040 161.895 78.865 162.225 ;
        RECT 79.035 161.895 79.310 162.225 ;
        RECT 79.035 161.725 79.205 161.895 ;
        RECT 76.235 161.155 76.405 161.535 ;
        RECT 76.585 160.985 76.915 161.365 ;
        RECT 77.095 161.155 77.355 161.660 ;
        RECT 77.540 161.555 79.205 161.725 ;
        RECT 79.480 161.660 79.650 162.395 ;
        RECT 80.345 162.345 81.125 162.515 ;
        RECT 81.295 162.565 81.465 163.195 ;
        RECT 81.635 162.735 81.965 163.535 ;
        RECT 82.135 162.565 82.410 163.365 ;
        RECT 81.295 162.355 82.410 162.565 ;
        RECT 82.585 162.370 82.875 163.535 ;
        RECT 83.085 162.395 83.315 163.535 ;
        RECT 83.485 162.385 83.815 163.365 ;
        RECT 83.985 162.395 84.195 163.535 ;
        RECT 84.555 163.195 86.605 163.365 ;
        RECT 84.555 162.695 84.805 163.195 ;
        RECT 84.975 162.525 85.185 163.025 ;
        RECT 85.395 162.695 85.605 163.195 ;
        RECT 85.935 162.525 86.185 163.025 ;
        RECT 86.355 162.695 86.605 163.195 ;
        RECT 86.775 162.525 87.025 163.365 ;
        RECT 87.195 162.695 87.445 163.535 ;
        RECT 87.615 162.525 87.870 163.365 ;
        RECT 77.540 161.205 77.795 161.555 ;
        RECT 77.965 160.985 78.295 161.385 ;
        RECT 78.465 161.205 78.635 161.555 ;
        RECT 78.805 160.985 79.185 161.385 ;
        RECT 79.375 161.315 79.650 161.660 ;
        RECT 80.365 161.805 80.580 162.345 ;
        RECT 80.750 161.975 81.520 162.175 ;
        RECT 81.690 161.975 82.410 162.175 ;
        RECT 83.065 161.975 83.395 162.225 ;
        RECT 80.365 161.635 81.965 161.805 ;
        RECT 80.795 161.625 81.965 161.635 ;
        RECT 80.335 160.985 80.625 161.455 ;
        RECT 80.795 161.155 81.125 161.625 ;
        RECT 81.295 160.985 81.465 161.455 ;
        RECT 81.635 161.155 81.965 161.625 ;
        RECT 82.135 160.985 82.410 161.805 ;
        RECT 82.585 160.985 82.875 161.710 ;
        RECT 83.085 160.985 83.315 161.805 ;
        RECT 83.565 161.785 83.815 162.385 ;
        RECT 84.425 162.355 85.185 162.525 ;
        RECT 84.425 161.805 84.885 162.355 ;
        RECT 85.380 162.185 85.645 162.525 ;
        RECT 85.935 162.355 87.870 162.525 ;
        RECT 88.105 162.445 89.315 163.535 ;
        RECT 85.055 161.975 85.645 162.185 ;
        RECT 85.835 161.975 86.885 162.185 ;
        RECT 87.055 161.975 87.885 162.185 ;
        RECT 88.105 161.905 88.625 162.445 ;
        RECT 83.485 161.155 83.815 161.785 ;
        RECT 83.985 160.985 84.195 161.805 ;
        RECT 84.425 161.625 87.485 161.805 ;
        RECT 84.475 160.985 84.765 161.455 ;
        RECT 84.935 161.155 85.265 161.625 ;
        RECT 85.435 160.985 86.145 161.455 ;
        RECT 86.315 161.155 86.645 161.625 ;
        RECT 86.815 160.985 86.985 161.455 ;
        RECT 87.155 161.155 87.485 161.625 ;
        RECT 87.655 160.985 87.930 161.805 ;
        RECT 88.795 161.735 89.315 162.275 ;
        RECT 88.105 160.985 89.315 161.735 ;
        RECT 18.100 160.815 89.400 160.985 ;
        RECT 18.185 160.065 19.395 160.815 ;
        RECT 18.185 159.525 18.705 160.065 ;
        RECT 19.570 159.975 19.830 160.815 ;
        RECT 20.005 160.070 20.260 160.645 ;
        RECT 20.430 160.435 20.760 160.815 ;
        RECT 20.975 160.265 21.145 160.645 ;
        RECT 20.430 160.095 21.145 160.265 ;
        RECT 21.405 160.315 21.665 160.645 ;
        RECT 21.875 160.335 22.150 160.815 ;
        RECT 18.875 159.355 19.395 159.895 ;
        RECT 18.185 158.265 19.395 159.355 ;
        RECT 19.570 158.265 19.830 159.415 ;
        RECT 20.005 159.340 20.175 160.070 ;
        RECT 20.430 159.905 20.600 160.095 ;
        RECT 20.345 159.575 20.600 159.905 ;
        RECT 20.430 159.365 20.600 159.575 ;
        RECT 20.880 159.545 21.235 159.915 ;
        RECT 21.405 159.405 21.575 160.315 ;
        RECT 22.360 160.245 22.565 160.645 ;
        RECT 22.735 160.415 23.070 160.815 ;
        RECT 21.745 159.575 22.105 160.155 ;
        RECT 22.360 160.075 23.045 160.245 ;
        RECT 22.285 159.405 22.535 159.905 ;
        RECT 20.005 158.435 20.260 159.340 ;
        RECT 20.430 159.195 21.145 159.365 ;
        RECT 20.430 158.265 20.760 159.025 ;
        RECT 20.975 158.435 21.145 159.195 ;
        RECT 21.405 159.235 22.535 159.405 ;
        RECT 21.405 158.465 21.675 159.235 ;
        RECT 22.705 159.045 23.045 160.075 ;
        RECT 21.845 158.265 22.175 159.045 ;
        RECT 22.380 158.870 23.045 159.045 ;
        RECT 23.245 160.140 23.505 160.645 ;
        RECT 23.685 160.435 24.015 160.815 ;
        RECT 24.195 160.265 24.365 160.645 ;
        RECT 24.625 160.270 29.970 160.815 ;
        RECT 23.245 159.340 23.415 160.140 ;
        RECT 23.700 160.095 24.365 160.265 ;
        RECT 23.700 159.840 23.870 160.095 ;
        RECT 23.585 159.510 23.870 159.840 ;
        RECT 24.105 159.545 24.435 159.915 ;
        RECT 23.700 159.365 23.870 159.510 ;
        RECT 26.210 159.440 26.550 160.270 ;
        RECT 30.665 159.995 30.875 160.815 ;
        RECT 31.045 160.015 31.375 160.645 ;
        RECT 22.380 158.465 22.565 158.870 ;
        RECT 22.735 158.265 23.070 158.690 ;
        RECT 23.245 158.435 23.515 159.340 ;
        RECT 23.700 159.195 24.365 159.365 ;
        RECT 23.685 158.265 24.015 159.025 ;
        RECT 24.195 158.435 24.365 159.195 ;
        RECT 28.030 158.700 28.380 159.950 ;
        RECT 31.045 159.415 31.295 160.015 ;
        RECT 31.545 159.995 31.775 160.815 ;
        RECT 32.185 160.185 32.515 160.545 ;
        RECT 33.145 160.355 33.395 160.815 ;
        RECT 33.565 160.355 34.115 160.645 ;
        RECT 32.185 159.995 33.575 160.185 ;
        RECT 33.405 159.905 33.575 159.995 ;
        RECT 31.465 159.575 31.795 159.825 ;
        RECT 31.985 159.575 32.675 159.825 ;
        RECT 32.905 159.575 33.235 159.825 ;
        RECT 33.405 159.575 33.695 159.905 ;
        RECT 24.625 158.265 29.970 158.700 ;
        RECT 30.665 158.265 30.875 159.405 ;
        RECT 31.045 158.435 31.375 159.415 ;
        RECT 31.545 158.265 31.775 159.405 ;
        RECT 31.985 159.135 32.300 159.575 ;
        RECT 33.405 159.325 33.575 159.575 ;
        RECT 32.635 159.155 33.575 159.325 ;
        RECT 32.185 158.265 32.465 158.935 ;
        RECT 32.635 158.605 32.935 159.155 ;
        RECT 33.865 158.985 34.115 160.355 ;
        RECT 34.285 160.015 34.575 160.815 ;
        RECT 34.750 160.075 35.005 160.645 ;
        RECT 35.175 160.415 35.505 160.815 ;
        RECT 35.930 160.280 36.460 160.645 ;
        RECT 35.930 160.245 36.105 160.280 ;
        RECT 35.175 160.075 36.105 160.245 ;
        RECT 34.750 159.405 34.920 160.075 ;
        RECT 35.175 159.905 35.345 160.075 ;
        RECT 35.090 159.575 35.345 159.905 ;
        RECT 35.570 159.575 35.765 159.905 ;
        RECT 33.145 158.265 33.475 158.985 ;
        RECT 33.665 158.435 34.115 158.985 ;
        RECT 34.285 158.265 34.575 159.405 ;
        RECT 34.750 158.435 35.085 159.405 ;
        RECT 35.255 158.265 35.425 159.405 ;
        RECT 35.595 158.605 35.765 159.575 ;
        RECT 35.935 158.945 36.105 160.075 ;
        RECT 36.275 159.285 36.445 160.085 ;
        RECT 36.650 159.795 36.925 160.645 ;
        RECT 36.645 159.625 36.925 159.795 ;
        RECT 36.650 159.485 36.925 159.625 ;
        RECT 37.095 159.285 37.285 160.645 ;
        RECT 37.465 160.280 37.975 160.815 ;
        RECT 38.195 160.005 38.440 160.610 ;
        RECT 38.885 160.045 40.555 160.815 ;
        RECT 40.890 160.305 41.130 160.815 ;
        RECT 41.310 160.305 41.590 160.635 ;
        RECT 41.820 160.305 42.035 160.815 ;
        RECT 37.485 159.835 38.715 160.005 ;
        RECT 36.275 159.115 37.285 159.285 ;
        RECT 37.455 159.270 38.205 159.460 ;
        RECT 35.935 158.775 37.060 158.945 ;
        RECT 37.455 158.605 37.625 159.270 ;
        RECT 38.375 159.025 38.715 159.835 ;
        RECT 38.885 159.525 39.635 160.045 ;
        RECT 39.805 159.355 40.555 159.875 ;
        RECT 40.785 159.575 41.140 160.135 ;
        RECT 41.310 159.405 41.480 160.305 ;
        RECT 41.650 159.575 41.915 160.135 ;
        RECT 42.205 160.075 42.820 160.645 ;
        RECT 43.945 160.090 44.235 160.815 ;
        RECT 42.165 159.405 42.335 159.905 ;
        RECT 35.595 158.435 37.625 158.605 ;
        RECT 37.795 158.265 37.965 159.025 ;
        RECT 38.200 158.615 38.715 159.025 ;
        RECT 38.885 158.265 40.555 159.355 ;
        RECT 40.910 159.235 42.335 159.405 ;
        RECT 40.910 159.060 41.300 159.235 ;
        RECT 41.785 158.265 42.115 159.065 ;
        RECT 42.505 159.055 42.820 160.075 ;
        RECT 44.405 159.995 45.090 160.635 ;
        RECT 45.260 159.995 45.430 160.815 ;
        RECT 45.600 160.165 45.930 160.630 ;
        RECT 46.100 160.345 46.270 160.815 ;
        RECT 46.530 160.425 47.715 160.595 ;
        RECT 47.885 160.255 48.215 160.645 ;
        RECT 46.915 160.165 47.300 160.255 ;
        RECT 45.600 159.995 47.300 160.165 ;
        RECT 47.705 160.075 48.215 160.255 ;
        RECT 48.555 160.095 48.885 160.815 ;
        RECT 49.430 160.415 51.045 160.585 ;
        RECT 51.215 160.415 51.545 160.815 ;
        RECT 50.875 160.245 51.045 160.415 ;
        RECT 51.715 160.340 52.050 160.600 ;
        RECT 42.285 158.435 42.820 159.055 ;
        RECT 43.945 158.265 44.235 159.430 ;
        RECT 44.405 159.025 44.655 159.995 ;
        RECT 44.825 159.615 45.160 159.825 ;
        RECT 45.330 159.615 45.780 159.825 ;
        RECT 45.970 159.615 46.455 159.825 ;
        RECT 44.990 159.445 45.160 159.615 ;
        RECT 46.080 159.455 46.455 159.615 ;
        RECT 46.645 159.575 47.025 159.825 ;
        RECT 47.205 159.615 47.535 159.825 ;
        RECT 44.990 159.275 45.910 159.445 ;
        RECT 44.405 158.435 45.070 159.025 ;
        RECT 45.240 158.265 45.570 159.105 ;
        RECT 45.740 159.025 45.910 159.275 ;
        RECT 46.080 159.285 46.475 159.455 ;
        RECT 46.080 159.195 46.455 159.285 ;
        RECT 46.645 159.195 46.965 159.575 ;
        RECT 47.705 159.445 47.875 160.075 ;
        RECT 48.045 159.615 48.375 159.905 ;
        RECT 48.610 159.795 48.960 159.905 ;
        RECT 48.605 159.625 48.960 159.795 ;
        RECT 48.610 159.575 48.960 159.625 ;
        RECT 49.270 159.575 49.690 160.240 ;
        RECT 49.860 160.135 50.150 160.235 ;
        RECT 50.340 160.135 50.610 160.235 ;
        RECT 49.860 159.965 50.155 160.135 ;
        RECT 50.340 159.965 50.615 160.135 ;
        RECT 50.875 160.075 51.435 160.245 ;
        RECT 49.860 159.575 50.150 159.965 ;
        RECT 50.340 159.575 50.610 159.965 ;
        RECT 51.265 159.905 51.435 160.075 ;
        RECT 50.820 159.795 51.070 159.905 ;
        RECT 50.820 159.625 51.075 159.795 ;
        RECT 50.820 159.575 51.070 159.625 ;
        RECT 51.265 159.575 51.570 159.905 ;
        RECT 47.135 159.275 48.220 159.445 ;
        RECT 48.610 159.285 48.815 159.575 ;
        RECT 51.265 159.405 51.435 159.575 ;
        RECT 47.135 159.025 47.305 159.275 ;
        RECT 45.740 158.855 47.305 159.025 ;
        RECT 46.080 158.435 46.885 158.855 ;
        RECT 47.475 158.265 47.725 159.105 ;
        RECT 47.920 158.435 48.220 159.275 ;
        RECT 49.065 159.235 51.435 159.405 ;
        RECT 48.635 158.605 48.805 159.105 ;
        RECT 49.065 158.775 49.235 159.235 ;
        RECT 49.465 158.855 50.890 159.025 ;
        RECT 49.465 158.605 49.795 158.855 ;
        RECT 48.635 158.435 49.795 158.605 ;
        RECT 50.020 158.265 50.350 158.685 ;
        RECT 50.605 158.435 50.890 158.855 ;
        RECT 51.135 158.265 51.465 159.065 ;
        RECT 51.795 158.985 52.050 160.340 ;
        RECT 52.230 160.050 52.685 160.815 ;
        RECT 52.960 160.435 54.260 160.645 ;
        RECT 54.515 160.455 54.845 160.815 ;
        RECT 54.090 160.285 54.260 160.435 ;
        RECT 55.015 160.315 55.275 160.645 ;
        RECT 55.045 160.305 55.275 160.315 ;
        RECT 53.160 159.825 53.380 160.225 ;
        RECT 52.225 159.625 52.715 159.825 ;
        RECT 52.905 159.615 53.380 159.825 ;
        RECT 53.625 159.825 53.835 160.225 ;
        RECT 54.090 160.160 54.845 160.285 ;
        RECT 54.090 160.115 54.935 160.160 ;
        RECT 54.665 159.995 54.935 160.115 ;
        RECT 53.625 159.615 53.955 159.825 ;
        RECT 54.125 159.555 54.535 159.860 ;
        RECT 51.715 158.475 52.050 158.985 ;
        RECT 52.230 159.385 53.405 159.445 ;
        RECT 54.765 159.420 54.935 159.995 ;
        RECT 54.735 159.385 54.935 159.420 ;
        RECT 52.230 159.275 54.935 159.385 ;
        RECT 52.230 158.655 52.485 159.275 ;
        RECT 53.075 159.215 54.875 159.275 ;
        RECT 53.075 159.185 53.405 159.215 ;
        RECT 55.105 159.115 55.275 160.305 ;
        RECT 55.445 160.270 60.790 160.815 ;
        RECT 57.030 159.440 57.370 160.270 ;
        RECT 60.975 160.220 61.225 160.645 ;
        RECT 61.395 160.390 61.725 160.815 ;
        RECT 61.895 160.395 62.985 160.645 ;
        RECT 63.175 160.395 64.265 160.645 ;
        RECT 61.895 160.220 62.065 160.395 ;
        RECT 60.975 160.050 62.065 160.220 ;
        RECT 62.235 160.055 63.925 160.225 ;
        RECT 64.095 160.220 64.265 160.395 ;
        RECT 64.435 160.390 64.765 160.815 ;
        RECT 64.935 160.220 65.255 160.645 ;
        RECT 52.735 159.015 52.920 159.105 ;
        RECT 53.510 159.015 54.345 159.025 ;
        RECT 52.735 158.815 54.345 159.015 ;
        RECT 52.735 158.775 52.965 158.815 ;
        RECT 52.230 158.435 52.565 158.655 ;
        RECT 53.570 158.265 53.925 158.645 ;
        RECT 54.095 158.435 54.345 158.815 ;
        RECT 54.595 158.265 54.845 159.045 ;
        RECT 55.015 158.435 55.275 159.115 ;
        RECT 58.850 158.700 59.200 159.950 ;
        RECT 61.030 159.795 61.660 159.825 ;
        RECT 61.950 159.795 62.580 159.825 ;
        RECT 61.025 159.625 61.660 159.795 ;
        RECT 61.945 159.625 62.580 159.795 ;
        RECT 62.750 159.415 63.040 160.055 ;
        RECT 64.095 160.050 65.255 160.220 ;
        RECT 65.585 160.085 65.875 160.815 ;
        RECT 63.325 159.625 63.980 159.825 ;
        RECT 64.270 159.795 65.380 159.825 ;
        RECT 64.245 159.625 65.380 159.795 ;
        RECT 65.575 159.575 65.875 159.905 ;
        RECT 66.055 159.885 66.285 160.525 ;
        RECT 66.465 160.265 66.775 160.635 ;
        RECT 66.955 160.445 67.625 160.815 ;
        RECT 66.465 160.065 67.695 160.265 ;
        RECT 66.055 159.575 66.580 159.885 ;
        RECT 66.760 159.575 67.225 159.885 ;
        RECT 60.975 159.245 63.040 159.415 ;
        RECT 55.445 158.265 60.790 158.700 ;
        RECT 60.975 158.435 61.225 159.245 ;
        RECT 61.395 158.605 61.645 159.075 ;
        RECT 61.815 158.775 62.145 159.245 ;
        RECT 62.315 158.605 62.485 159.075 ;
        RECT 62.655 158.775 63.040 159.245 ;
        RECT 63.255 159.245 65.185 159.415 ;
        RECT 67.405 159.395 67.695 160.065 ;
        RECT 63.255 158.605 63.505 159.245 ;
        RECT 61.395 158.435 63.505 158.605 ;
        RECT 63.675 158.265 63.845 159.075 ;
        RECT 64.015 158.435 64.345 159.245 ;
        RECT 64.515 158.265 64.685 159.075 ;
        RECT 64.855 158.435 65.185 159.245 ;
        RECT 65.585 159.155 66.745 159.395 ;
        RECT 65.585 158.445 65.845 159.155 ;
        RECT 66.015 158.265 66.345 158.975 ;
        RECT 66.515 158.445 66.745 159.155 ;
        RECT 66.925 159.175 67.695 159.395 ;
        RECT 66.925 158.445 67.195 159.175 ;
        RECT 67.375 158.265 67.715 158.995 ;
        RECT 67.885 158.445 68.145 160.635 ;
        RECT 68.325 160.065 69.535 160.815 ;
        RECT 69.705 160.090 69.995 160.815 ;
        RECT 68.325 159.525 68.845 160.065 ;
        RECT 69.015 159.355 69.535 159.895 ;
        RECT 68.325 158.265 69.535 159.355 ;
        RECT 69.705 158.265 69.995 159.430 ;
        RECT 70.165 158.435 70.445 160.535 ;
        RECT 70.675 160.355 70.845 160.815 ;
        RECT 71.115 160.425 72.365 160.605 ;
        RECT 71.500 160.185 71.865 160.255 ;
        RECT 70.615 160.005 71.865 160.185 ;
        RECT 72.035 160.205 72.365 160.425 ;
        RECT 72.535 160.375 72.705 160.815 ;
        RECT 72.875 160.205 73.215 160.620 ;
        RECT 73.385 160.435 74.275 160.605 ;
        RECT 72.035 160.035 73.215 160.205 ;
        RECT 70.615 159.405 70.890 160.005 ;
        RECT 73.385 159.880 73.935 160.265 ;
        RECT 71.060 159.575 71.415 159.825 ;
        RECT 71.610 159.795 72.075 159.825 ;
        RECT 71.605 159.625 72.075 159.795 ;
        RECT 71.610 159.575 72.075 159.625 ;
        RECT 72.245 159.575 72.575 159.825 ;
        RECT 72.750 159.625 73.215 159.825 ;
        RECT 74.105 159.710 74.275 160.435 ;
        RECT 73.385 159.640 74.275 159.710 ;
        RECT 74.445 160.110 74.665 160.595 ;
        RECT 74.835 160.275 75.085 160.815 ;
        RECT 75.255 160.165 75.515 160.645 ;
        RECT 75.685 160.435 76.575 160.605 ;
        RECT 74.445 159.685 74.775 160.110 ;
        RECT 72.395 159.455 72.575 159.575 ;
        RECT 73.385 159.615 74.280 159.640 ;
        RECT 73.385 159.600 74.290 159.615 ;
        RECT 73.385 159.585 74.295 159.600 ;
        RECT 73.385 159.580 74.305 159.585 ;
        RECT 73.385 159.570 74.310 159.580 ;
        RECT 73.385 159.560 74.315 159.570 ;
        RECT 73.385 159.555 74.325 159.560 ;
        RECT 73.385 159.545 74.335 159.555 ;
        RECT 73.385 159.540 74.345 159.545 ;
        RECT 70.615 159.195 72.225 159.405 ;
        RECT 72.395 159.285 72.725 159.455 ;
        RECT 71.815 159.095 72.225 159.195 ;
        RECT 70.635 158.265 71.420 159.025 ;
        RECT 71.815 158.435 72.200 159.095 ;
        RECT 72.525 158.495 72.725 159.285 ;
        RECT 72.895 158.265 73.215 159.445 ;
        RECT 73.385 159.090 73.645 159.540 ;
        RECT 74.010 159.535 74.345 159.540 ;
        RECT 74.010 159.530 74.360 159.535 ;
        RECT 74.010 159.520 74.375 159.530 ;
        RECT 74.010 159.515 74.400 159.520 ;
        RECT 74.945 159.515 75.175 159.910 ;
        RECT 74.010 159.510 75.175 159.515 ;
        RECT 74.040 159.475 75.175 159.510 ;
        RECT 74.075 159.450 75.175 159.475 ;
        RECT 74.105 159.420 75.175 159.450 ;
        RECT 74.125 159.390 75.175 159.420 ;
        RECT 74.145 159.360 75.175 159.390 ;
        RECT 74.215 159.350 75.175 159.360 ;
        RECT 74.240 159.340 75.175 159.350 ;
        RECT 74.260 159.325 75.175 159.340 ;
        RECT 74.280 159.310 75.175 159.325 ;
        RECT 74.285 159.300 75.070 159.310 ;
        RECT 74.300 159.265 75.070 159.300 ;
        RECT 73.815 158.945 74.145 159.190 ;
        RECT 74.315 159.015 75.070 159.265 ;
        RECT 75.345 159.135 75.515 160.165 ;
        RECT 75.685 159.880 76.235 160.265 ;
        RECT 76.405 159.710 76.575 160.435 ;
        RECT 73.815 158.920 74.000 158.945 ;
        RECT 73.385 158.820 74.000 158.920 ;
        RECT 73.385 158.265 73.990 158.820 ;
        RECT 74.165 158.435 74.645 158.775 ;
        RECT 74.815 158.265 75.070 158.810 ;
        RECT 75.240 158.435 75.515 159.135 ;
        RECT 75.685 159.640 76.575 159.710 ;
        RECT 76.745 160.110 76.965 160.595 ;
        RECT 77.135 160.275 77.385 160.815 ;
        RECT 77.555 160.165 77.815 160.645 ;
        RECT 78.905 160.305 79.210 160.815 ;
        RECT 76.745 159.685 77.075 160.110 ;
        RECT 75.685 159.615 76.580 159.640 ;
        RECT 75.685 159.600 76.590 159.615 ;
        RECT 75.685 159.585 76.595 159.600 ;
        RECT 75.685 159.580 76.605 159.585 ;
        RECT 75.685 159.570 76.610 159.580 ;
        RECT 75.685 159.560 76.615 159.570 ;
        RECT 75.685 159.555 76.625 159.560 ;
        RECT 75.685 159.545 76.635 159.555 ;
        RECT 75.685 159.540 76.645 159.545 ;
        RECT 75.685 159.090 75.945 159.540 ;
        RECT 76.310 159.535 76.645 159.540 ;
        RECT 76.310 159.530 76.660 159.535 ;
        RECT 76.310 159.520 76.675 159.530 ;
        RECT 76.310 159.515 76.700 159.520 ;
        RECT 77.245 159.515 77.475 159.910 ;
        RECT 76.310 159.510 77.475 159.515 ;
        RECT 76.340 159.475 77.475 159.510 ;
        RECT 76.375 159.450 77.475 159.475 ;
        RECT 76.405 159.420 77.475 159.450 ;
        RECT 76.425 159.390 77.475 159.420 ;
        RECT 76.445 159.360 77.475 159.390 ;
        RECT 76.515 159.350 77.475 159.360 ;
        RECT 76.540 159.340 77.475 159.350 ;
        RECT 76.560 159.325 77.475 159.340 ;
        RECT 76.580 159.310 77.475 159.325 ;
        RECT 76.585 159.300 77.370 159.310 ;
        RECT 76.600 159.265 77.370 159.300 ;
        RECT 76.115 158.945 76.445 159.190 ;
        RECT 76.615 159.015 77.370 159.265 ;
        RECT 77.645 159.135 77.815 160.165 ;
        RECT 78.905 159.575 79.220 160.135 ;
        RECT 79.390 159.825 79.640 160.635 ;
        RECT 79.810 160.290 80.070 160.815 ;
        RECT 80.250 159.825 80.500 160.635 ;
        RECT 80.670 160.255 80.930 160.815 ;
        RECT 81.100 160.165 81.360 160.620 ;
        RECT 81.530 160.335 81.790 160.815 ;
        RECT 81.960 160.165 82.220 160.620 ;
        RECT 82.390 160.335 82.650 160.815 ;
        RECT 82.820 160.165 83.080 160.620 ;
        RECT 83.250 160.335 83.495 160.815 ;
        RECT 83.665 160.165 83.940 160.620 ;
        RECT 84.110 160.335 84.355 160.815 ;
        RECT 84.525 160.165 84.785 160.620 ;
        RECT 84.965 160.335 85.215 160.815 ;
        RECT 85.385 160.165 85.645 160.620 ;
        RECT 85.825 160.335 86.075 160.815 ;
        RECT 86.245 160.165 86.505 160.620 ;
        RECT 86.685 160.335 86.945 160.815 ;
        RECT 87.115 160.165 87.375 160.620 ;
        RECT 87.545 160.335 87.845 160.815 ;
        RECT 81.100 159.995 87.845 160.165 ;
        RECT 88.105 160.065 89.315 160.815 ;
        RECT 79.390 159.575 86.510 159.825 ;
        RECT 76.115 158.920 76.300 158.945 ;
        RECT 75.685 158.820 76.300 158.920 ;
        RECT 75.685 158.265 76.290 158.820 ;
        RECT 76.465 158.435 76.945 158.775 ;
        RECT 77.115 158.265 77.370 158.810 ;
        RECT 77.540 158.435 77.815 159.135 ;
        RECT 78.915 158.265 79.210 159.075 ;
        RECT 79.390 158.435 79.635 159.575 ;
        RECT 79.810 158.265 80.070 159.075 ;
        RECT 80.250 158.440 80.500 159.575 ;
        RECT 86.680 159.405 87.845 159.995 ;
        RECT 81.100 159.180 87.845 159.405 ;
        RECT 88.105 159.355 88.625 159.895 ;
        RECT 88.795 159.525 89.315 160.065 ;
        RECT 81.100 159.165 86.505 159.180 ;
        RECT 80.670 158.270 80.930 159.065 ;
        RECT 81.100 158.440 81.360 159.165 ;
        RECT 81.530 158.270 81.790 158.995 ;
        RECT 81.960 158.440 82.220 159.165 ;
        RECT 82.390 158.270 82.650 158.995 ;
        RECT 82.820 158.440 83.080 159.165 ;
        RECT 83.250 158.270 83.510 158.995 ;
        RECT 83.680 158.440 83.940 159.165 ;
        RECT 84.110 158.270 84.355 158.995 ;
        RECT 84.525 158.440 84.785 159.165 ;
        RECT 84.970 158.270 85.215 158.995 ;
        RECT 85.385 158.440 85.645 159.165 ;
        RECT 85.830 158.270 86.075 158.995 ;
        RECT 86.245 158.440 86.505 159.165 ;
        RECT 86.690 158.270 86.945 158.995 ;
        RECT 87.115 158.440 87.405 159.180 ;
        RECT 80.670 158.265 86.945 158.270 ;
        RECT 87.575 158.265 87.845 159.010 ;
        RECT 88.105 158.265 89.315 159.355 ;
        RECT 18.100 158.095 89.400 158.265 ;
        RECT 18.185 157.005 19.395 158.095 ;
        RECT 18.185 156.295 18.705 156.835 ;
        RECT 18.875 156.465 19.395 157.005 ;
        RECT 20.490 156.955 20.810 158.095 ;
        RECT 20.990 156.785 21.185 157.835 ;
        RECT 21.365 157.245 21.695 157.925 ;
        RECT 21.895 157.295 22.150 158.095 ;
        RECT 22.415 157.475 22.585 157.905 ;
        RECT 22.755 157.645 23.085 158.095 ;
        RECT 22.415 157.245 23.095 157.475 ;
        RECT 21.365 156.965 21.715 157.245 ;
        RECT 20.550 156.735 20.810 156.785 ;
        RECT 20.545 156.565 20.810 156.735 ;
        RECT 20.550 156.455 20.810 156.565 ;
        RECT 20.990 156.455 21.375 156.785 ;
        RECT 21.545 156.585 21.715 156.965 ;
        RECT 21.905 156.755 22.150 157.115 ;
        RECT 21.545 156.415 22.065 156.585 ;
        RECT 18.185 155.545 19.395 156.295 ;
        RECT 20.490 156.075 21.705 156.245 ;
        RECT 20.490 155.725 20.780 156.075 ;
        RECT 20.975 155.545 21.305 155.905 ;
        RECT 21.475 155.770 21.705 156.075 ;
        RECT 21.895 155.850 22.065 156.415 ;
        RECT 22.390 156.395 22.690 157.075 ;
        RECT 22.385 156.225 22.690 156.395 ;
        RECT 22.860 156.595 23.095 157.245 ;
        RECT 23.285 156.935 23.570 157.880 ;
        RECT 23.750 157.625 24.435 158.095 ;
        RECT 23.745 157.105 24.440 157.415 ;
        RECT 24.615 157.040 24.920 157.825 ;
        RECT 25.105 157.140 25.375 158.095 ;
        RECT 25.550 157.295 25.805 158.095 ;
        RECT 26.005 157.245 26.335 157.925 ;
        RECT 23.285 156.785 24.145 156.935 ;
        RECT 23.285 156.765 24.575 156.785 ;
        RECT 22.860 156.265 23.415 156.595 ;
        RECT 23.585 156.405 24.575 156.765 ;
        RECT 22.860 156.115 23.075 156.265 ;
        RECT 22.335 155.545 22.665 156.050 ;
        RECT 22.835 155.740 23.075 156.115 ;
        RECT 23.585 156.070 23.755 156.405 ;
        RECT 24.745 156.235 24.920 157.040 ;
        RECT 25.550 156.755 25.795 157.115 ;
        RECT 25.985 156.965 26.335 157.245 ;
        RECT 25.985 156.585 26.155 156.965 ;
        RECT 26.515 156.785 26.710 157.835 ;
        RECT 26.890 156.955 27.210 158.095 ;
        RECT 27.385 157.005 30.895 158.095 ;
        RECT 23.355 155.875 23.755 156.070 ;
        RECT 23.355 155.730 23.525 155.875 ;
        RECT 24.115 155.545 24.515 156.040 ;
        RECT 24.685 155.715 24.920 156.235 ;
        RECT 25.635 156.415 26.155 156.585 ;
        RECT 26.325 156.455 26.710 156.785 ;
        RECT 26.890 156.735 27.150 156.785 ;
        RECT 26.890 156.565 27.155 156.735 ;
        RECT 26.890 156.455 27.150 156.565 ;
        RECT 25.105 155.545 25.375 156.180 ;
        RECT 25.635 155.850 25.805 156.415 ;
        RECT 27.385 156.315 29.035 156.835 ;
        RECT 29.205 156.485 30.895 157.005 ;
        RECT 31.065 156.930 31.355 158.095 ;
        RECT 31.530 156.945 31.790 158.095 ;
        RECT 31.965 157.020 32.220 157.925 ;
        RECT 32.390 157.335 32.720 158.095 ;
        RECT 32.935 157.165 33.105 157.925 ;
        RECT 25.995 156.075 27.210 156.245 ;
        RECT 25.995 155.770 26.225 156.075 ;
        RECT 26.395 155.545 26.725 155.905 ;
        RECT 26.920 155.725 27.210 156.075 ;
        RECT 27.385 155.545 30.895 156.315 ;
        RECT 31.065 155.545 31.355 156.270 ;
        RECT 31.530 155.545 31.790 156.385 ;
        RECT 31.965 156.290 32.135 157.020 ;
        RECT 32.390 156.995 33.105 157.165 ;
        RECT 33.365 157.005 36.875 158.095 ;
        RECT 38.165 157.425 38.445 158.095 ;
        RECT 38.615 157.205 38.915 157.755 ;
        RECT 39.115 157.375 39.445 158.095 ;
        RECT 39.635 157.375 40.095 157.925 ;
        RECT 40.265 157.660 45.610 158.095 ;
        RECT 32.390 156.785 32.560 156.995 ;
        RECT 32.305 156.455 32.560 156.785 ;
        RECT 31.965 155.715 32.220 156.290 ;
        RECT 32.390 156.265 32.560 156.455 ;
        RECT 32.840 156.445 33.195 156.815 ;
        RECT 33.365 156.315 35.015 156.835 ;
        RECT 35.185 156.485 36.875 157.005 ;
        RECT 37.980 156.785 38.245 157.145 ;
        RECT 38.615 157.035 39.555 157.205 ;
        RECT 39.385 156.785 39.555 157.035 ;
        RECT 37.980 156.535 38.655 156.785 ;
        RECT 38.875 156.535 39.215 156.785 ;
        RECT 39.385 156.455 39.675 156.785 ;
        RECT 39.385 156.365 39.555 156.455 ;
        RECT 32.390 156.095 33.105 156.265 ;
        RECT 32.390 155.545 32.720 155.925 ;
        RECT 32.935 155.715 33.105 156.095 ;
        RECT 33.365 155.545 36.875 156.315 ;
        RECT 38.165 156.175 39.555 156.365 ;
        RECT 38.165 155.815 38.495 156.175 ;
        RECT 39.845 156.005 40.095 157.375 ;
        RECT 41.850 156.090 42.190 156.920 ;
        RECT 43.670 156.410 44.020 157.660 ;
        RECT 45.785 157.005 47.455 158.095 ;
        RECT 45.785 156.315 46.535 156.835 ;
        RECT 46.705 156.485 47.455 157.005 ;
        RECT 47.625 156.490 47.905 157.925 ;
        RECT 48.075 157.320 48.785 158.095 ;
        RECT 48.955 157.150 49.285 157.925 ;
        RECT 48.135 156.935 49.285 157.150 ;
        RECT 39.115 155.545 39.365 156.005 ;
        RECT 39.535 155.715 40.095 156.005 ;
        RECT 40.265 155.545 45.610 156.090 ;
        RECT 45.785 155.545 47.455 156.315 ;
        RECT 47.625 155.715 47.965 156.490 ;
        RECT 48.135 156.365 48.420 156.935 ;
        RECT 48.605 156.535 49.075 156.765 ;
        RECT 49.480 156.735 49.695 157.850 ;
        RECT 49.875 157.375 50.205 158.095 ;
        RECT 49.985 156.735 50.215 157.075 ;
        RECT 50.385 157.005 52.055 158.095 ;
        RECT 52.315 157.475 52.485 157.905 ;
        RECT 52.655 157.645 52.985 158.095 ;
        RECT 52.315 157.245 52.995 157.475 ;
        RECT 49.245 156.555 49.695 156.735 ;
        RECT 49.245 156.535 49.575 156.555 ;
        RECT 49.885 156.535 50.215 156.735 ;
        RECT 48.135 156.175 48.845 156.365 ;
        RECT 48.545 156.035 48.845 156.175 ;
        RECT 49.035 156.175 50.215 156.365 ;
        RECT 49.035 156.095 49.365 156.175 ;
        RECT 48.545 156.025 48.860 156.035 ;
        RECT 48.545 156.015 48.870 156.025 ;
        RECT 48.545 156.010 48.880 156.015 ;
        RECT 48.135 155.545 48.305 156.005 ;
        RECT 48.545 156.000 48.885 156.010 ;
        RECT 48.545 155.995 48.890 156.000 ;
        RECT 48.545 155.985 48.895 155.995 ;
        RECT 48.545 155.980 48.900 155.985 ;
        RECT 48.545 155.715 48.905 155.980 ;
        RECT 49.535 155.545 49.705 156.005 ;
        RECT 49.875 155.715 50.215 156.175 ;
        RECT 50.385 156.315 51.135 156.835 ;
        RECT 51.305 156.485 52.055 157.005 ;
        RECT 52.290 156.735 52.590 157.075 ;
        RECT 52.285 156.565 52.590 156.735 ;
        RECT 50.385 155.545 52.055 156.315 ;
        RECT 52.290 156.225 52.590 156.565 ;
        RECT 52.760 156.595 52.995 157.245 ;
        RECT 53.185 156.935 53.470 157.880 ;
        RECT 53.650 157.625 54.335 158.095 ;
        RECT 53.645 157.105 54.340 157.415 ;
        RECT 54.515 157.040 54.820 157.825 ;
        RECT 55.005 157.140 55.275 158.095 ;
        RECT 53.185 156.785 54.045 156.935 ;
        RECT 53.185 156.765 54.475 156.785 ;
        RECT 52.760 156.265 53.315 156.595 ;
        RECT 53.485 156.405 54.475 156.765 ;
        RECT 52.760 156.115 52.975 156.265 ;
        RECT 52.235 155.545 52.565 156.050 ;
        RECT 52.735 155.740 52.975 156.115 ;
        RECT 53.485 156.070 53.655 156.405 ;
        RECT 54.645 156.235 54.820 157.040 ;
        RECT 55.445 157.005 56.655 158.095 ;
        RECT 53.255 155.875 53.655 156.070 ;
        RECT 53.255 155.730 53.425 155.875 ;
        RECT 54.015 155.545 54.415 156.040 ;
        RECT 54.585 155.715 54.820 156.235 ;
        RECT 55.445 156.295 55.965 156.835 ;
        RECT 56.135 156.465 56.655 157.005 ;
        RECT 56.825 156.930 57.115 158.095 ;
        RECT 57.725 156.955 58.065 158.095 ;
        RECT 58.235 157.415 58.405 157.925 ;
        RECT 58.615 157.595 58.865 158.095 ;
        RECT 59.075 157.715 60.335 157.925 ;
        RECT 59.075 157.415 59.325 157.715 ;
        RECT 58.235 157.245 59.325 157.415 ;
        RECT 59.555 157.245 59.905 157.545 ;
        RECT 60.075 157.295 60.335 157.715 ;
        RECT 58.235 157.205 58.405 157.245 ;
        RECT 59.165 156.885 59.565 157.075 ;
        RECT 57.670 156.475 58.085 156.785 ;
        RECT 58.255 156.455 58.615 156.785 ;
        RECT 58.825 156.535 59.190 156.715 ;
        RECT 55.005 155.545 55.275 156.180 ;
        RECT 55.445 155.545 56.655 156.295 ;
        RECT 56.825 155.545 57.115 156.270 ;
        RECT 57.725 155.545 58.065 156.265 ;
        RECT 58.255 155.875 58.455 156.455 ;
        RECT 58.825 156.225 59.015 156.535 ;
        RECT 59.395 156.455 59.565 156.885 ;
        RECT 59.735 156.265 59.905 157.245 ;
        RECT 60.505 157.005 62.175 158.095 ;
        RECT 60.075 156.455 60.335 156.785 ;
        RECT 58.715 155.805 59.015 156.225 ;
        RECT 59.255 156.095 59.905 156.265 ;
        RECT 60.505 156.315 61.255 156.835 ;
        RECT 61.425 156.485 62.175 157.005 ;
        RECT 62.815 157.485 63.145 157.915 ;
        RECT 63.325 157.655 63.520 158.095 ;
        RECT 63.690 157.485 64.020 157.915 ;
        RECT 62.815 157.315 64.020 157.485 ;
        RECT 62.815 156.985 63.710 157.315 ;
        RECT 64.190 157.145 64.465 157.915 ;
        RECT 65.110 157.585 66.765 157.875 ;
        RECT 63.880 156.955 64.465 157.145 ;
        RECT 65.110 157.245 66.700 157.415 ;
        RECT 66.935 157.295 67.215 158.095 ;
        RECT 65.110 156.955 65.430 157.245 ;
        RECT 66.530 157.125 66.700 157.245 ;
        RECT 62.820 156.455 63.115 156.785 ;
        RECT 63.295 156.455 63.710 156.785 ;
        RECT 59.255 156.055 59.505 156.095 ;
        RECT 59.185 155.885 59.505 156.055 ;
        RECT 59.255 155.755 59.505 155.885 ;
        RECT 59.995 155.545 60.325 155.925 ;
        RECT 60.505 155.545 62.175 156.315 ;
        RECT 62.815 155.545 63.115 156.275 ;
        RECT 63.295 155.835 63.525 156.455 ;
        RECT 63.880 156.285 64.055 156.955 ;
        RECT 65.625 156.905 66.340 157.075 ;
        RECT 66.530 156.955 67.255 157.125 ;
        RECT 67.425 156.955 67.695 157.925 ;
        RECT 67.865 157.005 70.455 158.095 ;
        RECT 71.085 157.540 71.690 158.095 ;
        RECT 71.865 157.585 72.345 157.925 ;
        RECT 72.515 157.550 72.770 158.095 ;
        RECT 71.085 157.440 71.700 157.540 ;
        RECT 71.515 157.415 71.700 157.440 ;
        RECT 63.725 156.105 64.055 156.285 ;
        RECT 64.225 156.135 64.465 156.785 ;
        RECT 65.110 156.215 65.460 156.785 ;
        RECT 65.630 156.455 66.340 156.905 ;
        RECT 67.085 156.785 67.255 156.955 ;
        RECT 66.510 156.455 66.915 156.785 ;
        RECT 67.085 156.455 67.355 156.785 ;
        RECT 67.085 156.285 67.255 156.455 ;
        RECT 65.645 156.115 67.255 156.285 ;
        RECT 67.525 156.220 67.695 156.955 ;
        RECT 63.725 155.725 63.950 156.105 ;
        RECT 64.120 155.545 64.450 155.935 ;
        RECT 65.115 155.545 65.445 156.045 ;
        RECT 65.645 155.765 65.815 156.115 ;
        RECT 66.015 155.545 66.345 155.945 ;
        RECT 66.515 155.765 66.685 156.115 ;
        RECT 66.855 155.545 67.235 155.945 ;
        RECT 67.425 155.875 67.695 156.220 ;
        RECT 67.865 156.315 69.075 156.835 ;
        RECT 69.245 156.485 70.455 157.005 ;
        RECT 71.085 156.820 71.345 157.270 ;
        RECT 71.515 157.170 71.845 157.415 ;
        RECT 72.015 157.095 72.770 157.345 ;
        RECT 72.940 157.225 73.215 157.925 ;
        RECT 72.000 157.060 72.770 157.095 ;
        RECT 71.985 157.050 72.770 157.060 ;
        RECT 71.980 157.035 72.875 157.050 ;
        RECT 71.960 157.020 72.875 157.035 ;
        RECT 71.940 157.010 72.875 157.020 ;
        RECT 71.915 157.000 72.875 157.010 ;
        RECT 71.845 156.970 72.875 157.000 ;
        RECT 71.825 156.940 72.875 156.970 ;
        RECT 71.805 156.910 72.875 156.940 ;
        RECT 71.775 156.885 72.875 156.910 ;
        RECT 71.740 156.850 72.875 156.885 ;
        RECT 71.710 156.845 72.875 156.850 ;
        RECT 71.710 156.840 72.100 156.845 ;
        RECT 71.710 156.830 72.075 156.840 ;
        RECT 71.710 156.825 72.060 156.830 ;
        RECT 71.710 156.820 72.045 156.825 ;
        RECT 71.085 156.815 72.045 156.820 ;
        RECT 71.085 156.805 72.035 156.815 ;
        RECT 71.085 156.800 72.025 156.805 ;
        RECT 71.085 156.790 72.015 156.800 ;
        RECT 71.085 156.780 72.010 156.790 ;
        RECT 71.085 156.775 72.005 156.780 ;
        RECT 71.085 156.760 71.995 156.775 ;
        RECT 71.085 156.745 71.990 156.760 ;
        RECT 71.085 156.720 71.980 156.745 ;
        RECT 71.085 156.650 71.975 156.720 ;
        RECT 67.865 155.545 70.455 156.315 ;
        RECT 71.085 156.095 71.635 156.480 ;
        RECT 71.805 155.925 71.975 156.650 ;
        RECT 71.085 155.755 71.975 155.925 ;
        RECT 72.145 156.250 72.475 156.675 ;
        RECT 72.645 156.450 72.875 156.845 ;
        RECT 72.145 155.765 72.365 156.250 ;
        RECT 73.045 156.195 73.215 157.225 ;
        RECT 73.395 156.955 73.725 158.095 ;
        RECT 74.255 157.125 74.585 157.910 ;
        RECT 73.905 156.955 74.585 157.125 ;
        RECT 74.765 157.005 78.275 158.095 ;
        RECT 73.385 156.535 73.735 156.785 ;
        RECT 73.905 156.355 74.075 156.955 ;
        RECT 74.245 156.535 74.595 156.785 ;
        RECT 72.535 155.545 72.785 156.085 ;
        RECT 72.955 155.715 73.215 156.195 ;
        RECT 73.395 155.545 73.665 156.355 ;
        RECT 73.835 155.715 74.165 156.355 ;
        RECT 74.335 155.545 74.575 156.355 ;
        RECT 74.765 156.315 76.415 156.835 ;
        RECT 76.585 156.485 78.275 157.005 ;
        RECT 79.445 157.165 79.625 157.925 ;
        RECT 79.805 157.335 80.135 158.095 ;
        RECT 79.445 156.995 80.120 157.165 ;
        RECT 80.305 157.020 80.575 157.925 ;
        RECT 80.750 157.670 81.085 158.095 ;
        RECT 81.255 157.490 81.440 157.895 ;
        RECT 79.950 156.850 80.120 156.995 ;
        RECT 79.385 156.445 79.725 156.815 ;
        RECT 79.950 156.520 80.225 156.850 ;
        RECT 74.765 155.545 78.275 156.315 ;
        RECT 79.950 156.265 80.120 156.520 ;
        RECT 79.455 156.095 80.120 156.265 ;
        RECT 80.395 156.220 80.575 157.020 ;
        RECT 79.455 155.715 79.625 156.095 ;
        RECT 79.805 155.545 80.135 155.925 ;
        RECT 80.315 155.715 80.575 156.220 ;
        RECT 80.775 157.315 81.440 157.490 ;
        RECT 81.645 157.315 81.975 158.095 ;
        RECT 80.775 156.285 81.115 157.315 ;
        RECT 82.145 157.125 82.415 157.895 ;
        RECT 81.285 156.955 82.415 157.125 ;
        RECT 81.285 156.455 81.535 156.955 ;
        RECT 80.775 156.115 81.460 156.285 ;
        RECT 81.715 156.205 82.075 156.785 ;
        RECT 80.750 155.545 81.085 155.945 ;
        RECT 81.255 155.715 81.460 156.115 ;
        RECT 82.245 156.045 82.415 156.955 ;
        RECT 82.585 156.930 82.875 158.095 ;
        RECT 83.595 157.515 83.765 157.925 ;
        RECT 83.935 157.715 84.265 158.095 ;
        RECT 84.910 157.715 85.580 158.095 ;
        RECT 85.815 157.545 85.985 157.925 ;
        RECT 86.155 157.715 86.495 158.095 ;
        RECT 86.665 157.545 86.835 157.925 ;
        RECT 87.175 157.715 87.505 158.095 ;
        RECT 87.675 157.545 87.935 157.925 ;
        RECT 83.595 157.345 85.345 157.515 ;
        RECT 83.570 156.735 83.750 157.095 ;
        RECT 83.565 156.565 83.750 156.735 ;
        RECT 83.570 156.455 83.750 156.565 ;
        RECT 81.670 155.545 81.945 156.025 ;
        RECT 82.155 155.715 82.415 156.045 ;
        RECT 82.585 155.545 82.875 156.270 ;
        RECT 83.920 156.265 84.090 157.345 ;
        RECT 84.410 157.005 84.740 157.175 ;
        RECT 83.595 156.095 84.090 156.265 ;
        RECT 83.595 155.715 83.765 156.095 ;
        RECT 83.935 155.545 84.265 155.925 ;
        RECT 84.435 155.715 84.660 157.005 ;
        RECT 85.175 156.785 85.345 157.345 ;
        RECT 85.655 157.375 86.835 157.545 ;
        RECT 87.005 157.375 87.935 157.545 ;
        RECT 84.835 156.265 85.005 156.785 ;
        RECT 85.175 156.455 85.485 156.785 ;
        RECT 85.655 156.265 85.825 157.375 ;
        RECT 87.005 157.205 87.175 157.375 ;
        RECT 85.995 157.035 87.175 157.205 ;
        RECT 85.995 156.860 86.165 157.035 ;
        RECT 86.325 156.565 86.595 156.735 ;
        RECT 84.835 156.095 85.825 156.265 ;
        RECT 84.830 155.545 85.160 155.925 ;
        RECT 85.430 155.715 85.600 156.095 ;
        RECT 86.330 155.880 86.595 156.565 ;
        RECT 86.770 155.885 87.075 156.865 ;
        RECT 87.245 156.225 87.595 156.765 ;
        RECT 87.765 156.045 87.935 157.375 ;
        RECT 88.105 157.005 89.315 158.095 ;
        RECT 88.105 156.465 88.625 157.005 ;
        RECT 88.795 156.295 89.315 156.835 ;
        RECT 87.255 155.545 87.505 156.045 ;
        RECT 87.675 155.715 87.935 156.045 ;
        RECT 88.105 155.545 89.315 156.295 ;
        RECT 18.100 155.375 89.400 155.545 ;
        RECT 18.185 154.625 19.395 155.375 ;
        RECT 19.565 154.805 20.000 155.205 ;
        RECT 20.170 154.975 20.555 155.375 ;
        RECT 19.565 154.635 20.555 154.805 ;
        RECT 20.725 154.635 21.150 155.205 ;
        RECT 21.340 154.805 21.595 155.205 ;
        RECT 21.765 154.975 22.150 155.375 ;
        RECT 21.340 154.635 22.150 154.805 ;
        RECT 22.320 154.635 22.565 155.205 ;
        RECT 22.755 154.805 23.010 155.205 ;
        RECT 23.180 154.975 23.565 155.375 ;
        RECT 22.755 154.635 23.565 154.805 ;
        RECT 23.735 154.635 23.995 155.205 ;
        RECT 25.170 154.805 25.345 155.205 ;
        RECT 25.515 154.995 25.845 155.375 ;
        RECT 26.090 154.875 26.320 155.205 ;
        RECT 25.170 154.635 25.800 154.805 ;
        RECT 18.185 154.085 18.705 154.625 ;
        RECT 20.220 154.465 20.555 154.635 ;
        RECT 20.800 154.465 21.150 154.635 ;
        RECT 21.800 154.465 22.150 154.635 ;
        RECT 22.395 154.465 22.565 154.635 ;
        RECT 23.215 154.465 23.565 154.635 ;
        RECT 18.875 153.915 19.395 154.455 ;
        RECT 18.185 152.825 19.395 153.915 ;
        RECT 19.565 153.760 20.050 154.465 ;
        RECT 20.220 154.135 20.630 154.465 ;
        RECT 20.220 153.590 20.555 154.135 ;
        RECT 20.800 153.965 21.630 154.465 ;
        RECT 19.565 153.420 20.555 153.590 ;
        RECT 20.725 153.785 21.630 153.965 ;
        RECT 21.800 154.135 22.225 154.465 ;
        RECT 19.565 152.995 20.000 153.420 ;
        RECT 20.170 152.825 20.555 153.250 ;
        RECT 20.725 152.995 21.150 153.785 ;
        RECT 21.800 153.615 22.150 154.135 ;
        RECT 22.395 153.965 23.045 154.465 ;
        RECT 21.320 153.420 22.150 153.615 ;
        RECT 22.320 153.785 23.045 153.965 ;
        RECT 23.215 154.135 23.640 154.465 ;
        RECT 21.320 152.995 21.595 153.420 ;
        RECT 21.765 152.825 22.150 153.250 ;
        RECT 22.320 152.995 22.565 153.785 ;
        RECT 23.215 153.615 23.565 154.135 ;
        RECT 23.810 153.965 23.995 154.635 ;
        RECT 25.630 154.465 25.800 154.635 ;
        RECT 22.755 153.420 23.565 153.615 ;
        RECT 22.755 152.995 23.010 153.420 ;
        RECT 23.180 152.825 23.565 153.250 ;
        RECT 23.735 152.995 23.995 153.965 ;
        RECT 25.085 153.785 25.450 154.465 ;
        RECT 25.630 154.135 25.980 154.465 ;
        RECT 25.630 153.615 25.800 154.135 ;
        RECT 25.170 153.445 25.800 153.615 ;
        RECT 26.150 153.585 26.320 154.875 ;
        RECT 26.520 153.765 26.800 155.040 ;
        RECT 27.025 154.015 27.295 155.040 ;
        RECT 27.755 154.995 28.085 155.375 ;
        RECT 28.255 155.120 28.590 155.165 ;
        RECT 26.985 153.845 27.295 154.015 ;
        RECT 27.025 153.765 27.295 153.845 ;
        RECT 27.485 153.765 27.825 154.795 ;
        RECT 28.255 154.655 28.595 155.120 ;
        RECT 27.995 154.135 28.255 154.465 ;
        RECT 27.995 153.585 28.165 154.135 ;
        RECT 28.425 153.965 28.595 154.655 ;
        RECT 25.170 152.995 25.345 153.445 ;
        RECT 26.150 153.415 28.165 153.585 ;
        RECT 25.515 152.825 25.845 153.265 ;
        RECT 26.150 152.995 26.320 153.415 ;
        RECT 26.555 152.825 27.225 153.235 ;
        RECT 27.440 152.995 27.610 153.415 ;
        RECT 27.810 152.825 28.140 153.235 ;
        RECT 28.335 152.995 28.595 153.965 ;
        RECT 28.765 154.875 29.025 155.205 ;
        RECT 29.335 154.995 29.665 155.375 ;
        RECT 29.845 155.035 31.325 155.205 ;
        RECT 28.765 154.175 28.935 154.875 ;
        RECT 29.845 154.705 30.245 155.035 ;
        RECT 29.285 154.515 29.495 154.695 ;
        RECT 29.285 154.345 29.905 154.515 ;
        RECT 30.075 154.225 30.245 154.705 ;
        RECT 30.435 154.535 30.985 154.865 ;
        RECT 28.765 154.005 29.895 154.175 ;
        RECT 30.075 154.055 30.645 154.225 ;
        RECT 28.765 153.325 28.935 154.005 ;
        RECT 29.725 153.885 29.895 154.005 ;
        RECT 29.105 153.505 29.455 153.835 ;
        RECT 29.725 153.715 30.305 153.885 ;
        RECT 30.475 153.545 30.645 154.055 ;
        RECT 29.905 153.375 30.645 153.545 ;
        RECT 30.815 153.545 30.985 154.535 ;
        RECT 31.155 154.135 31.325 155.035 ;
        RECT 31.575 154.465 31.760 155.045 ;
        RECT 32.030 154.465 32.225 155.040 ;
        RECT 32.435 154.995 32.765 155.375 ;
        RECT 31.575 154.135 31.805 154.465 ;
        RECT 32.030 154.135 32.285 154.465 ;
        RECT 31.575 153.825 31.760 154.135 ;
        RECT 32.030 153.825 32.225 154.135 ;
        RECT 32.595 153.545 32.765 154.465 ;
        RECT 30.815 153.375 32.765 153.545 ;
        RECT 28.765 152.995 29.025 153.325 ;
        RECT 29.335 152.825 29.665 153.205 ;
        RECT 29.905 152.995 30.095 153.375 ;
        RECT 30.345 152.825 30.675 153.205 ;
        RECT 30.885 152.995 31.055 153.375 ;
        RECT 31.250 152.825 31.580 153.205 ;
        RECT 31.840 152.995 32.010 153.375 ;
        RECT 32.435 152.825 32.765 153.205 ;
        RECT 32.935 152.995 33.195 155.205 ;
        RECT 33.365 154.605 35.955 155.375 ;
        RECT 36.280 154.725 36.610 155.190 ;
        RECT 36.780 154.905 36.950 155.375 ;
        RECT 37.120 154.725 37.450 155.205 ;
        RECT 33.365 154.085 34.575 154.605 ;
        RECT 36.280 154.555 37.450 154.725 ;
        RECT 34.745 153.915 35.955 154.435 ;
        RECT 36.125 154.175 36.770 154.385 ;
        RECT 36.940 154.175 37.510 154.385 ;
        RECT 37.680 154.005 37.850 155.205 ;
        RECT 38.390 154.805 38.560 155.010 ;
        RECT 33.365 152.825 35.955 153.915 ;
        RECT 36.340 152.825 36.670 153.925 ;
        RECT 37.145 153.595 37.850 154.005 ;
        RECT 38.020 154.635 38.560 154.805 ;
        RECT 38.840 154.635 39.010 155.375 ;
        RECT 39.275 154.635 39.635 155.010 ;
        RECT 38.020 153.935 38.190 154.635 ;
        RECT 38.360 154.135 38.690 154.465 ;
        RECT 38.860 154.135 39.210 154.465 ;
        RECT 38.020 153.765 38.645 153.935 ;
        RECT 38.860 153.595 39.125 154.135 ;
        RECT 39.380 153.980 39.635 154.635 ;
        RECT 39.805 154.605 43.315 155.375 ;
        RECT 43.945 154.650 44.235 155.375 ;
        RECT 39.805 154.085 41.455 154.605 ;
        RECT 37.145 153.425 39.125 153.595 ;
        RECT 37.145 152.995 37.470 153.425 ;
        RECT 37.640 152.825 37.970 153.245 ;
        RECT 38.715 152.825 39.125 153.255 ;
        RECT 39.295 152.995 39.635 153.980 ;
        RECT 41.625 153.915 43.315 154.435 ;
        RECT 39.805 152.825 43.315 153.915 ;
        RECT 43.945 152.825 44.235 153.990 ;
        RECT 44.410 153.775 44.745 155.195 ;
        RECT 44.925 155.005 45.670 155.375 ;
        RECT 46.235 154.835 46.490 155.195 ;
        RECT 46.670 155.005 47.000 155.375 ;
        RECT 47.180 154.835 47.405 155.195 ;
        RECT 44.920 154.645 47.405 154.835 ;
        RECT 44.920 153.955 45.145 154.645 ;
        RECT 45.345 154.135 45.625 154.465 ;
        RECT 45.805 154.135 46.380 154.465 ;
        RECT 46.560 154.135 46.995 154.465 ;
        RECT 47.175 154.135 47.445 154.465 ;
        RECT 44.920 153.775 47.415 153.955 ;
        RECT 44.410 153.005 44.675 153.775 ;
        RECT 44.845 152.825 45.175 153.545 ;
        RECT 45.365 153.365 46.555 153.595 ;
        RECT 45.365 153.005 45.625 153.365 ;
        RECT 45.795 152.825 46.125 153.195 ;
        RECT 46.295 153.005 46.555 153.365 ;
        RECT 47.125 153.005 47.415 153.775 ;
        RECT 47.635 153.005 47.895 155.195 ;
        RECT 48.155 155.005 48.825 155.375 ;
        RECT 49.005 154.825 49.315 155.195 ;
        RECT 48.085 154.625 49.315 154.825 ;
        RECT 48.085 153.955 48.375 154.625 ;
        RECT 49.495 154.445 49.725 155.085 ;
        RECT 49.905 154.645 50.195 155.375 ;
        RECT 50.385 154.605 52.055 155.375 ;
        RECT 48.555 154.135 49.020 154.445 ;
        RECT 49.200 154.135 49.725 154.445 ;
        RECT 49.905 154.135 50.205 154.465 ;
        RECT 50.385 154.085 51.135 154.605 ;
        RECT 52.235 154.565 52.505 155.375 ;
        RECT 52.675 154.565 53.005 155.205 ;
        RECT 53.175 154.565 53.415 155.375 ;
        RECT 53.605 154.830 58.950 155.375 ;
        RECT 48.085 153.735 48.855 153.955 ;
        RECT 48.065 152.825 48.405 153.555 ;
        RECT 48.585 153.005 48.855 153.735 ;
        RECT 49.035 153.715 50.195 153.955 ;
        RECT 51.305 153.915 52.055 154.435 ;
        RECT 52.225 154.135 52.575 154.385 ;
        RECT 52.745 153.965 52.915 154.565 ;
        RECT 53.085 154.135 53.435 154.385 ;
        RECT 55.190 154.000 55.530 154.830 ;
        RECT 59.125 154.605 62.635 155.375 ;
        RECT 62.805 154.625 64.015 155.375 ;
        RECT 49.035 153.005 49.265 153.715 ;
        RECT 49.435 152.825 49.765 153.535 ;
        RECT 49.935 153.005 50.195 153.715 ;
        RECT 50.385 152.825 52.055 153.915 ;
        RECT 52.235 152.825 52.565 153.965 ;
        RECT 52.745 153.795 53.425 153.965 ;
        RECT 53.095 153.010 53.425 153.795 ;
        RECT 57.010 153.260 57.360 154.510 ;
        RECT 59.125 154.085 60.775 154.605 ;
        RECT 60.945 153.915 62.635 154.435 ;
        RECT 62.805 154.085 63.325 154.625 ;
        RECT 64.245 154.555 64.455 155.375 ;
        RECT 64.625 154.575 64.955 155.205 ;
        RECT 63.495 153.915 64.015 154.455 ;
        RECT 64.625 153.975 64.875 154.575 ;
        RECT 65.125 154.555 65.355 155.375 ;
        RECT 65.565 154.605 69.075 155.375 ;
        RECT 69.705 154.650 69.995 155.375 ;
        RECT 70.185 154.645 70.475 155.375 ;
        RECT 65.045 154.135 65.375 154.385 ;
        RECT 65.565 154.085 67.215 154.605 ;
        RECT 53.605 152.825 58.950 153.260 ;
        RECT 59.125 152.825 62.635 153.915 ;
        RECT 62.805 152.825 64.015 153.915 ;
        RECT 64.245 152.825 64.455 153.965 ;
        RECT 64.625 152.995 64.955 153.975 ;
        RECT 65.125 152.825 65.355 153.965 ;
        RECT 67.385 153.915 69.075 154.435 ;
        RECT 70.175 154.135 70.475 154.465 ;
        RECT 70.655 154.445 70.885 155.085 ;
        RECT 71.065 154.825 71.375 155.195 ;
        RECT 71.555 155.005 72.225 155.375 ;
        RECT 71.065 154.625 72.295 154.825 ;
        RECT 70.655 154.135 71.180 154.445 ;
        RECT 71.360 154.135 71.825 154.445 ;
        RECT 65.565 152.825 69.075 153.915 ;
        RECT 69.705 152.825 69.995 153.990 ;
        RECT 72.005 153.955 72.295 154.625 ;
        RECT 70.185 153.715 71.345 153.955 ;
        RECT 70.185 153.005 70.445 153.715 ;
        RECT 70.615 152.825 70.945 153.535 ;
        RECT 71.115 153.005 71.345 153.715 ;
        RECT 71.525 153.735 72.295 153.955 ;
        RECT 71.525 153.005 71.795 153.735 ;
        RECT 71.975 152.825 72.315 153.555 ;
        RECT 72.485 153.005 72.745 155.195 ;
        RECT 72.925 154.915 73.485 155.205 ;
        RECT 73.655 154.915 73.905 155.375 ;
        RECT 72.925 153.545 73.175 154.915 ;
        RECT 74.525 154.745 74.855 155.105 ;
        RECT 75.225 154.830 80.570 155.375 ;
        RECT 73.465 154.555 74.855 154.745 ;
        RECT 73.465 154.465 73.635 154.555 ;
        RECT 73.345 154.135 73.635 154.465 ;
        RECT 73.805 154.135 74.145 154.385 ;
        RECT 74.365 154.135 75.040 154.385 ;
        RECT 73.465 153.885 73.635 154.135 ;
        RECT 73.465 153.715 74.405 153.885 ;
        RECT 74.775 153.775 75.040 154.135 ;
        RECT 76.810 154.000 77.150 154.830 ;
        RECT 81.665 154.700 81.925 155.205 ;
        RECT 82.105 154.995 82.435 155.375 ;
        RECT 82.615 154.825 82.785 155.205 ;
        RECT 72.925 152.995 73.385 153.545 ;
        RECT 73.575 152.825 73.905 153.545 ;
        RECT 74.105 153.165 74.405 153.715 ;
        RECT 74.575 152.825 74.855 153.495 ;
        RECT 78.630 153.260 78.980 154.510 ;
        RECT 81.665 153.900 81.845 154.700 ;
        RECT 82.120 154.655 82.785 154.825 ;
        RECT 83.135 154.825 83.305 155.205 ;
        RECT 83.485 154.995 83.815 155.375 ;
        RECT 83.135 154.655 83.800 154.825 ;
        RECT 83.995 154.700 84.255 155.205 ;
        RECT 82.120 154.400 82.290 154.655 ;
        RECT 82.015 154.070 82.290 154.400 ;
        RECT 82.515 154.105 82.855 154.475 ;
        RECT 83.065 154.105 83.405 154.475 ;
        RECT 83.630 154.400 83.800 154.655 ;
        RECT 82.120 153.925 82.290 154.070 ;
        RECT 83.630 154.070 83.905 154.400 ;
        RECT 83.630 153.925 83.800 154.070 ;
        RECT 75.225 152.825 80.570 153.260 ;
        RECT 81.665 152.995 81.935 153.900 ;
        RECT 82.120 153.755 82.795 153.925 ;
        RECT 82.105 152.825 82.435 153.585 ;
        RECT 82.615 152.995 82.795 153.755 ;
        RECT 83.125 153.755 83.800 153.925 ;
        RECT 84.075 153.900 84.255 154.700 ;
        RECT 84.430 154.535 84.690 155.375 ;
        RECT 84.865 154.630 85.120 155.205 ;
        RECT 85.290 154.995 85.620 155.375 ;
        RECT 85.835 154.825 86.005 155.205 ;
        RECT 85.290 154.655 86.005 154.825 ;
        RECT 86.355 154.825 86.525 155.205 ;
        RECT 86.740 154.995 87.070 155.375 ;
        RECT 86.355 154.655 87.070 154.825 ;
        RECT 83.125 152.995 83.305 153.755 ;
        RECT 83.485 152.825 83.815 153.585 ;
        RECT 83.985 152.995 84.255 153.900 ;
        RECT 84.430 152.825 84.690 153.975 ;
        RECT 84.865 153.900 85.035 154.630 ;
        RECT 85.290 154.465 85.460 154.655 ;
        RECT 85.205 154.135 85.460 154.465 ;
        RECT 85.290 153.925 85.460 154.135 ;
        RECT 85.740 154.105 86.095 154.475 ;
        RECT 86.265 154.105 86.620 154.475 ;
        RECT 86.900 154.465 87.070 154.655 ;
        RECT 87.240 154.630 87.495 155.205 ;
        RECT 86.900 154.135 87.155 154.465 ;
        RECT 86.900 153.925 87.070 154.135 ;
        RECT 84.865 152.995 85.120 153.900 ;
        RECT 85.290 153.755 86.005 153.925 ;
        RECT 85.290 152.825 85.620 153.585 ;
        RECT 85.835 152.995 86.005 153.755 ;
        RECT 86.355 153.755 87.070 153.925 ;
        RECT 87.325 153.900 87.495 154.630 ;
        RECT 87.670 154.535 87.930 155.375 ;
        RECT 88.105 154.625 89.315 155.375 ;
        RECT 86.355 152.995 86.525 153.755 ;
        RECT 86.740 152.825 87.070 153.585 ;
        RECT 87.240 152.995 87.495 153.900 ;
        RECT 87.670 152.825 87.930 153.975 ;
        RECT 88.105 153.915 88.625 154.455 ;
        RECT 88.795 154.085 89.315 154.625 ;
        RECT 88.105 152.825 89.315 153.915 ;
        RECT 18.100 152.655 89.400 152.825 ;
        RECT 18.185 151.565 19.395 152.655 ;
        RECT 18.185 150.855 18.705 151.395 ;
        RECT 18.875 151.025 19.395 151.565 ;
        RECT 19.565 151.515 19.855 152.655 ;
        RECT 20.025 151.935 20.475 152.485 ;
        RECT 20.665 151.935 20.995 152.655 ;
        RECT 18.185 150.105 19.395 150.855 ;
        RECT 19.565 150.105 19.855 150.905 ;
        RECT 20.025 150.565 20.275 151.935 ;
        RECT 21.205 151.765 21.505 152.315 ;
        RECT 21.675 151.985 21.955 152.655 ;
        RECT 22.415 152.035 22.585 152.465 ;
        RECT 22.755 152.205 23.085 152.655 ;
        RECT 22.415 151.805 23.090 152.035 ;
        RECT 20.565 151.595 21.505 151.765 ;
        RECT 20.565 151.345 20.735 151.595 ;
        RECT 21.840 151.345 22.155 151.785 ;
        RECT 20.445 151.015 20.735 151.345 ;
        RECT 20.905 151.095 21.235 151.345 ;
        RECT 21.465 151.095 22.155 151.345 ;
        RECT 20.565 150.925 20.735 151.015 ;
        RECT 20.565 150.735 21.955 150.925 ;
        RECT 22.385 150.785 22.685 151.635 ;
        RECT 22.855 151.155 23.090 151.805 ;
        RECT 23.260 151.495 23.545 152.440 ;
        RECT 23.725 152.185 24.410 152.655 ;
        RECT 23.720 151.665 24.415 151.975 ;
        RECT 24.590 151.600 24.895 152.385 ;
        RECT 23.260 151.345 24.120 151.495 ;
        RECT 23.260 151.325 24.545 151.345 ;
        RECT 22.855 150.825 23.390 151.155 ;
        RECT 23.560 150.965 24.545 151.325 ;
        RECT 20.025 150.275 20.575 150.565 ;
        RECT 20.745 150.105 20.995 150.565 ;
        RECT 21.625 150.375 21.955 150.735 ;
        RECT 22.855 150.675 23.075 150.825 ;
        RECT 22.330 150.105 22.665 150.610 ;
        RECT 22.835 150.300 23.075 150.675 ;
        RECT 23.560 150.630 23.730 150.965 ;
        RECT 24.720 150.795 24.895 151.600 ;
        RECT 25.085 151.565 26.755 152.655 ;
        RECT 27.385 152.145 27.645 152.655 ;
        RECT 23.355 150.435 23.730 150.630 ;
        RECT 23.355 150.290 23.525 150.435 ;
        RECT 24.090 150.105 24.485 150.600 ;
        RECT 24.655 150.275 24.895 150.795 ;
        RECT 25.085 150.875 25.835 151.395 ;
        RECT 26.005 151.045 26.755 151.565 ;
        RECT 27.385 151.095 27.725 151.975 ;
        RECT 27.895 151.265 28.065 152.485 ;
        RECT 28.305 152.150 28.920 152.655 ;
        RECT 28.305 151.615 28.555 151.980 ;
        RECT 28.725 151.975 28.920 152.150 ;
        RECT 29.090 152.145 29.565 152.485 ;
        RECT 29.735 152.110 29.950 152.655 ;
        RECT 28.725 151.785 29.055 151.975 ;
        RECT 29.275 151.615 29.990 151.910 ;
        RECT 30.160 151.785 30.435 152.485 ;
        RECT 28.305 151.445 30.095 151.615 ;
        RECT 27.895 151.015 28.690 151.265 ;
        RECT 27.895 150.925 28.145 151.015 ;
        RECT 25.085 150.105 26.755 150.875 ;
        RECT 27.385 150.105 27.645 150.925 ;
        RECT 27.815 150.505 28.145 150.925 ;
        RECT 28.860 150.590 29.115 151.445 ;
        RECT 28.325 150.325 29.115 150.590 ;
        RECT 29.285 150.745 29.695 151.265 ;
        RECT 29.865 151.015 30.095 151.445 ;
        RECT 30.265 150.755 30.435 151.785 ;
        RECT 31.065 151.490 31.355 152.655 ;
        RECT 31.525 152.145 31.785 152.655 ;
        RECT 31.525 151.095 31.865 151.975 ;
        RECT 32.035 151.265 32.205 152.485 ;
        RECT 32.445 152.150 33.060 152.655 ;
        RECT 32.445 151.615 32.695 151.980 ;
        RECT 32.865 151.975 33.060 152.150 ;
        RECT 33.230 152.145 33.705 152.485 ;
        RECT 33.875 152.110 34.090 152.655 ;
        RECT 32.865 151.785 33.195 151.975 ;
        RECT 33.415 151.615 34.130 151.910 ;
        RECT 34.300 151.785 34.575 152.485 ;
        RECT 32.445 151.445 34.235 151.615 ;
        RECT 32.035 151.015 32.830 151.265 ;
        RECT 32.035 150.925 32.285 151.015 ;
        RECT 29.285 150.325 29.485 150.745 ;
        RECT 29.675 150.105 30.005 150.565 ;
        RECT 30.175 150.275 30.435 150.755 ;
        RECT 31.065 150.105 31.355 150.830 ;
        RECT 31.525 150.105 31.785 150.925 ;
        RECT 31.955 150.505 32.285 150.925 ;
        RECT 33.000 150.590 33.255 151.445 ;
        RECT 32.465 150.325 33.255 150.590 ;
        RECT 33.425 150.745 33.835 151.265 ;
        RECT 34.005 151.015 34.235 151.445 ;
        RECT 34.405 150.755 34.575 151.785 ;
        RECT 35.730 151.685 36.000 152.480 ;
        RECT 36.180 151.855 36.395 152.655 ;
        RECT 36.575 151.685 36.860 152.480 ;
        RECT 35.730 151.515 36.860 151.685 ;
        RECT 35.710 151.045 36.210 151.310 ;
        RECT 36.430 151.015 36.815 151.345 ;
        RECT 37.040 151.015 37.320 152.485 ;
        RECT 37.500 151.070 37.830 152.485 ;
        RECT 38.000 151.310 38.205 152.485 ;
        RECT 38.375 151.665 38.585 152.480 ;
        RECT 38.825 151.835 39.155 152.655 ;
        RECT 38.375 151.485 39.025 151.665 ;
        RECT 39.330 151.640 39.585 152.480 ;
        RECT 39.810 152.230 40.145 152.655 ;
        RECT 40.315 152.050 40.500 152.455 ;
        RECT 38.000 151.070 38.430 151.310 ;
        RECT 36.430 150.865 36.735 151.015 ;
        RECT 33.425 150.325 33.625 150.745 ;
        RECT 33.815 150.105 34.145 150.565 ;
        RECT 34.315 150.275 34.575 150.755 ;
        RECT 35.765 150.105 36.005 150.780 ;
        RECT 36.180 150.305 36.735 150.865 ;
        RECT 38.805 150.845 39.025 151.485 ;
        RECT 36.915 150.675 39.025 150.845 ;
        RECT 36.915 150.280 37.120 150.675 ;
        RECT 37.805 150.670 39.025 150.675 ;
        RECT 37.290 150.105 37.635 150.505 ;
        RECT 37.805 150.280 38.135 150.670 ;
        RECT 38.410 150.105 39.085 150.490 ;
        RECT 39.255 150.275 39.585 151.640 ;
        RECT 39.835 151.875 40.500 152.050 ;
        RECT 40.705 151.875 41.035 152.655 ;
        RECT 39.835 150.845 40.175 151.875 ;
        RECT 41.205 151.685 41.475 152.455 ;
        RECT 40.345 151.515 41.475 151.685 ;
        RECT 41.655 151.515 41.985 152.655 ;
        RECT 42.515 151.685 42.845 152.470 ;
        RECT 43.685 151.985 43.965 152.655 ;
        RECT 44.135 151.765 44.435 152.315 ;
        RECT 44.635 151.935 44.965 152.655 ;
        RECT 45.155 151.935 45.615 152.485 ;
        RECT 42.165 151.515 42.845 151.685 ;
        RECT 40.345 151.015 40.595 151.515 ;
        RECT 39.835 150.675 40.520 150.845 ;
        RECT 40.775 150.765 41.135 151.345 ;
        RECT 39.810 150.105 40.145 150.505 ;
        RECT 40.315 150.275 40.520 150.675 ;
        RECT 41.305 150.605 41.475 151.515 ;
        RECT 41.645 151.095 41.995 151.345 ;
        RECT 42.165 150.915 42.335 151.515 ;
        RECT 43.500 151.345 43.765 151.705 ;
        RECT 44.135 151.595 45.075 151.765 ;
        RECT 44.905 151.345 45.075 151.595 ;
        RECT 42.505 151.095 42.855 151.345 ;
        RECT 43.500 151.095 44.175 151.345 ;
        RECT 44.395 151.095 44.735 151.345 ;
        RECT 44.905 151.015 45.195 151.345 ;
        RECT 44.905 150.925 45.075 151.015 ;
        RECT 40.730 150.105 41.005 150.585 ;
        RECT 41.215 150.275 41.475 150.605 ;
        RECT 41.655 150.105 41.925 150.915 ;
        RECT 42.095 150.275 42.425 150.915 ;
        RECT 42.595 150.105 42.835 150.915 ;
        RECT 43.685 150.735 45.075 150.925 ;
        RECT 43.685 150.375 44.015 150.735 ;
        RECT 45.365 150.565 45.615 151.935 ;
        RECT 46.280 151.855 46.530 152.655 ;
        RECT 46.700 152.025 47.030 152.485 ;
        RECT 47.200 152.195 47.415 152.655 ;
        RECT 46.700 151.855 47.870 152.025 ;
        RECT 45.790 151.685 46.070 151.845 ;
        RECT 45.790 151.515 47.125 151.685 ;
        RECT 46.955 151.345 47.125 151.515 ;
        RECT 45.790 151.095 46.140 151.335 ;
        RECT 46.310 151.095 46.785 151.335 ;
        RECT 46.955 151.095 47.330 151.345 ;
        RECT 46.955 150.925 47.125 151.095 ;
        RECT 44.635 150.105 44.885 150.565 ;
        RECT 45.055 150.275 45.615 150.565 ;
        RECT 45.790 150.755 47.125 150.925 ;
        RECT 45.790 150.545 46.060 150.755 ;
        RECT 47.500 150.565 47.870 151.855 ;
        RECT 48.085 151.565 49.755 152.655 ;
        RECT 46.280 150.105 46.610 150.565 ;
        RECT 47.120 150.275 47.870 150.565 ;
        RECT 48.085 150.875 48.835 151.395 ;
        RECT 49.005 151.045 49.755 151.565 ;
        RECT 50.385 151.805 50.725 152.445 ;
        RECT 50.895 152.195 51.140 152.655 ;
        RECT 51.315 152.025 51.565 152.485 ;
        RECT 51.755 152.275 52.425 152.655 ;
        RECT 52.625 152.025 52.875 152.485 ;
        RECT 51.315 151.855 52.875 152.025 ;
        RECT 48.085 150.105 49.755 150.875 ;
        RECT 50.385 150.690 50.555 151.805 ;
        RECT 53.635 151.685 53.805 152.485 ;
        RECT 50.865 151.515 53.805 151.685 ;
        RECT 54.155 151.725 54.325 152.485 ;
        RECT 54.540 151.895 54.870 152.655 ;
        RECT 54.155 151.555 54.870 151.725 ;
        RECT 55.040 151.580 55.295 152.485 ;
        RECT 50.865 151.345 51.035 151.515 ;
        RECT 50.725 151.015 51.035 151.345 ;
        RECT 51.205 151.015 51.540 151.345 ;
        RECT 50.865 150.845 51.035 151.015 ;
        RECT 50.385 150.275 50.695 150.690 ;
        RECT 50.865 150.675 51.560 150.845 ;
        RECT 51.810 150.770 52.005 151.345 ;
        RECT 52.265 151.015 52.610 151.345 ;
        RECT 52.920 151.015 53.395 151.345 ;
        RECT 53.650 151.015 53.835 151.345 ;
        RECT 52.265 150.785 52.455 151.015 ;
        RECT 54.065 151.005 54.420 151.375 ;
        RECT 54.700 151.345 54.870 151.555 ;
        RECT 54.700 151.015 54.955 151.345 ;
        RECT 50.890 150.105 51.220 150.485 ;
        RECT 51.390 150.445 51.560 150.675 ;
        RECT 52.625 150.675 53.805 150.845 ;
        RECT 54.700 150.825 54.870 151.015 ;
        RECT 55.125 150.850 55.295 151.580 ;
        RECT 55.470 151.505 55.730 152.655 ;
        RECT 56.825 151.490 57.115 152.655 ;
        RECT 52.625 150.445 52.795 150.675 ;
        RECT 51.390 150.275 52.795 150.445 ;
        RECT 53.065 150.105 53.395 150.505 ;
        RECT 53.635 150.275 53.805 150.675 ;
        RECT 54.155 150.655 54.870 150.825 ;
        RECT 54.155 150.275 54.325 150.655 ;
        RECT 54.540 150.105 54.870 150.485 ;
        RECT 55.040 150.275 55.295 150.850 ;
        RECT 55.470 150.105 55.730 150.945 ;
        RECT 56.825 150.105 57.115 150.830 ;
        RECT 57.285 150.385 57.565 152.485 ;
        RECT 57.755 151.895 58.540 152.655 ;
        RECT 58.935 151.825 59.320 152.485 ;
        RECT 58.935 151.725 59.345 151.825 ;
        RECT 57.735 151.515 59.345 151.725 ;
        RECT 59.645 151.635 59.845 152.425 ;
        RECT 57.735 150.915 58.010 151.515 ;
        RECT 59.515 151.465 59.845 151.635 ;
        RECT 60.015 151.475 60.335 152.655 ;
        RECT 60.505 152.055 60.765 152.475 ;
        RECT 60.935 152.225 61.265 152.655 ;
        RECT 61.955 152.225 62.700 152.395 ;
        RECT 60.505 151.885 62.360 152.055 ;
        RECT 59.515 151.345 59.695 151.465 ;
        RECT 58.180 151.095 58.535 151.345 ;
        RECT 58.730 151.295 59.195 151.345 ;
        RECT 58.725 151.125 59.195 151.295 ;
        RECT 58.730 151.095 59.195 151.125 ;
        RECT 59.365 151.095 59.695 151.345 ;
        RECT 59.870 151.095 60.335 151.295 ;
        RECT 57.735 150.735 58.985 150.915 ;
        RECT 58.620 150.665 58.985 150.735 ;
        RECT 59.155 150.715 60.335 150.885 ;
        RECT 57.795 150.105 57.965 150.565 ;
        RECT 59.155 150.495 59.485 150.715 ;
        RECT 58.235 150.315 59.485 150.495 ;
        RECT 59.655 150.105 59.825 150.545 ;
        RECT 59.995 150.300 60.335 150.715 ;
        RECT 60.505 150.845 60.680 151.885 ;
        RECT 60.850 151.015 61.200 151.715 ;
        RECT 61.415 151.545 62.020 151.715 ;
        RECT 61.370 151.015 61.660 151.345 ;
        RECT 61.830 151.265 62.020 151.545 ;
        RECT 62.190 151.605 62.360 151.885 ;
        RECT 62.530 151.975 62.700 152.225 ;
        RECT 62.925 152.145 63.565 152.475 ;
        RECT 62.530 151.805 63.565 151.975 ;
        RECT 63.735 151.855 64.015 152.655 ;
        RECT 63.395 151.685 63.565 151.805 ;
        RECT 62.190 151.435 62.840 151.605 ;
        RECT 63.395 151.515 64.055 151.685 ;
        RECT 64.225 151.515 64.500 152.485 ;
        RECT 61.830 151.095 62.275 151.265 ;
        RECT 61.830 150.845 62.020 151.095 ;
        RECT 62.670 151.015 62.840 151.435 ;
        RECT 63.885 151.345 64.055 151.515 ;
        RECT 63.060 151.015 63.715 151.345 ;
        RECT 63.885 151.015 64.160 151.345 ;
        RECT 63.885 150.845 64.055 151.015 ;
        RECT 60.505 150.470 60.825 150.845 ;
        RECT 61.080 150.105 61.250 150.845 ;
        RECT 61.500 150.675 62.020 150.845 ;
        RECT 62.445 150.675 64.055 150.845 ;
        RECT 64.330 150.780 64.500 151.515 ;
        RECT 64.670 151.460 64.840 152.655 ;
        RECT 65.105 151.515 65.365 152.655 ;
        RECT 65.535 151.505 65.865 152.485 ;
        RECT 66.035 151.515 66.315 152.655 ;
        RECT 66.485 151.565 67.695 152.655 ;
        RECT 65.125 151.095 65.460 151.345 ;
        RECT 61.500 150.470 61.670 150.675 ;
        RECT 61.915 150.105 62.270 150.505 ;
        RECT 62.445 150.325 62.615 150.675 ;
        RECT 62.815 150.105 63.145 150.505 ;
        RECT 63.315 150.325 63.485 150.675 ;
        RECT 63.655 150.105 64.035 150.505 ;
        RECT 64.225 150.435 64.500 150.780 ;
        RECT 64.670 150.105 64.840 151.045 ;
        RECT 65.630 150.905 65.800 151.505 ;
        RECT 65.970 151.075 66.305 151.345 ;
        RECT 65.105 150.275 65.800 150.905 ;
        RECT 66.005 150.105 66.315 150.905 ;
        RECT 66.485 150.855 67.005 151.395 ;
        RECT 67.175 151.025 67.695 151.565 ;
        RECT 67.885 151.765 68.145 152.475 ;
        RECT 68.315 151.945 68.645 152.655 ;
        RECT 68.815 151.765 69.045 152.475 ;
        RECT 67.885 151.525 69.045 151.765 ;
        RECT 69.225 151.745 69.495 152.475 ;
        RECT 69.675 151.925 70.015 152.655 ;
        RECT 69.225 151.525 69.995 151.745 ;
        RECT 67.875 151.015 68.175 151.345 ;
        RECT 68.355 151.035 68.880 151.345 ;
        RECT 69.060 151.035 69.525 151.345 ;
        RECT 66.485 150.105 67.695 150.855 ;
        RECT 67.885 150.105 68.175 150.835 ;
        RECT 68.355 150.395 68.585 151.035 ;
        RECT 69.705 150.855 69.995 151.525 ;
        RECT 68.765 150.655 69.995 150.855 ;
        RECT 68.765 150.285 69.075 150.655 ;
        RECT 69.255 150.105 69.925 150.475 ;
        RECT 70.185 150.285 70.445 152.475 ;
        RECT 70.635 152.045 70.965 152.475 ;
        RECT 71.145 152.215 71.340 152.655 ;
        RECT 71.510 152.045 71.840 152.475 ;
        RECT 70.635 151.875 71.840 152.045 ;
        RECT 70.635 151.545 71.530 151.875 ;
        RECT 72.010 151.705 72.285 152.475 ;
        RECT 72.465 152.220 77.810 152.655 ;
        RECT 71.700 151.515 72.285 151.705 ;
        RECT 70.640 151.015 70.935 151.345 ;
        RECT 71.115 151.015 71.530 151.345 ;
        RECT 70.635 150.105 70.935 150.835 ;
        RECT 71.115 150.395 71.345 151.015 ;
        RECT 71.700 150.845 71.875 151.515 ;
        RECT 71.545 150.665 71.875 150.845 ;
        RECT 72.045 150.695 72.285 151.345 ;
        RECT 71.545 150.285 71.770 150.665 ;
        RECT 74.050 150.650 74.390 151.480 ;
        RECT 75.870 150.970 76.220 152.220 ;
        RECT 77.985 151.565 81.495 152.655 ;
        RECT 77.985 150.875 79.635 151.395 ;
        RECT 79.805 151.045 81.495 151.565 ;
        RECT 82.585 151.490 82.875 152.655 ;
        RECT 83.045 151.565 84.715 152.655 ;
        RECT 83.045 150.875 83.795 151.395 ;
        RECT 83.965 151.045 84.715 151.565 ;
        RECT 84.965 151.725 85.145 152.485 ;
        RECT 85.325 151.895 85.655 152.655 ;
        RECT 84.965 151.555 85.640 151.725 ;
        RECT 85.825 151.580 86.095 152.485 ;
        RECT 85.470 151.410 85.640 151.555 ;
        RECT 84.905 151.005 85.245 151.375 ;
        RECT 85.470 151.080 85.745 151.410 ;
        RECT 71.940 150.105 72.270 150.495 ;
        RECT 72.465 150.105 77.810 150.650 ;
        RECT 77.985 150.105 81.495 150.875 ;
        RECT 82.585 150.105 82.875 150.830 ;
        RECT 83.045 150.105 84.715 150.875 ;
        RECT 85.470 150.825 85.640 151.080 ;
        RECT 84.975 150.655 85.640 150.825 ;
        RECT 85.915 150.780 86.095 151.580 ;
        RECT 84.975 150.275 85.145 150.655 ;
        RECT 85.325 150.105 85.655 150.485 ;
        RECT 85.835 150.275 86.095 150.780 ;
        RECT 86.265 151.685 86.535 152.455 ;
        RECT 86.705 151.875 87.035 152.655 ;
        RECT 87.240 152.050 87.425 152.455 ;
        RECT 87.595 152.230 87.930 152.655 ;
        RECT 87.240 151.875 87.905 152.050 ;
        RECT 86.265 151.515 87.395 151.685 ;
        RECT 86.265 150.605 86.435 151.515 ;
        RECT 86.605 150.765 86.965 151.345 ;
        RECT 87.145 151.015 87.395 151.515 ;
        RECT 87.565 150.845 87.905 151.875 ;
        RECT 88.105 151.565 89.315 152.655 ;
        RECT 88.105 151.025 88.625 151.565 ;
        RECT 88.795 150.855 89.315 151.395 ;
        RECT 87.220 150.675 87.905 150.845 ;
        RECT 86.265 150.275 86.525 150.605 ;
        RECT 86.735 150.105 87.010 150.585 ;
        RECT 87.220 150.275 87.425 150.675 ;
        RECT 87.595 150.105 87.930 150.505 ;
        RECT 88.105 150.105 89.315 150.855 ;
        RECT 18.100 149.935 89.400 150.105 ;
        RECT 18.185 149.185 19.395 149.935 ;
        RECT 18.185 148.645 18.705 149.185 ;
        RECT 19.570 149.095 19.830 149.935 ;
        RECT 20.005 149.190 20.260 149.765 ;
        RECT 20.430 149.555 20.760 149.935 ;
        RECT 20.975 149.385 21.145 149.765 ;
        RECT 20.430 149.215 21.145 149.385 ;
        RECT 18.875 148.475 19.395 149.015 ;
        RECT 18.185 147.385 19.395 148.475 ;
        RECT 19.570 147.385 19.830 148.535 ;
        RECT 20.005 148.460 20.175 149.190 ;
        RECT 20.430 149.025 20.600 149.215 ;
        RECT 21.445 149.115 21.675 149.935 ;
        RECT 21.845 149.135 22.175 149.765 ;
        RECT 20.345 148.695 20.600 149.025 ;
        RECT 20.430 148.485 20.600 148.695 ;
        RECT 20.880 148.665 21.235 149.035 ;
        RECT 21.425 148.695 21.755 148.945 ;
        RECT 21.925 148.535 22.175 149.135 ;
        RECT 22.345 149.115 22.555 149.935 ;
        RECT 22.785 149.260 23.045 149.765 ;
        RECT 23.225 149.555 23.555 149.935 ;
        RECT 23.735 149.385 23.905 149.765 ;
        RECT 24.165 149.390 29.510 149.935 ;
        RECT 29.685 149.390 35.030 149.935 ;
        RECT 35.230 149.545 35.560 149.935 ;
        RECT 20.005 147.555 20.260 148.460 ;
        RECT 20.430 148.315 21.145 148.485 ;
        RECT 20.430 147.385 20.760 148.145 ;
        RECT 20.975 147.555 21.145 148.315 ;
        RECT 21.445 147.385 21.675 148.525 ;
        RECT 21.845 147.555 22.175 148.535 ;
        RECT 22.345 147.385 22.555 148.525 ;
        RECT 22.785 148.460 22.955 149.260 ;
        RECT 23.240 149.215 23.905 149.385 ;
        RECT 23.240 148.960 23.410 149.215 ;
        RECT 23.125 148.630 23.410 148.960 ;
        RECT 23.645 148.665 23.975 149.035 ;
        RECT 23.240 148.485 23.410 148.630 ;
        RECT 25.750 148.560 26.090 149.390 ;
        RECT 22.785 147.555 23.055 148.460 ;
        RECT 23.240 148.315 23.905 148.485 ;
        RECT 23.225 147.385 23.555 148.145 ;
        RECT 23.735 147.555 23.905 148.315 ;
        RECT 27.570 147.820 27.920 149.070 ;
        RECT 31.270 148.560 31.610 149.390 ;
        RECT 35.730 149.375 35.955 149.755 ;
        RECT 33.090 147.820 33.440 149.070 ;
        RECT 35.215 148.695 35.455 149.345 ;
        RECT 35.625 149.195 35.955 149.375 ;
        RECT 35.625 148.525 35.800 149.195 ;
        RECT 36.155 149.025 36.385 149.645 ;
        RECT 36.565 149.205 36.865 149.935 ;
        RECT 37.135 149.385 37.305 149.765 ;
        RECT 37.520 149.555 37.850 149.935 ;
        RECT 37.135 149.215 37.850 149.385 ;
        RECT 35.970 148.695 36.385 149.025 ;
        RECT 36.565 148.695 36.860 149.025 ;
        RECT 37.045 148.665 37.400 149.035 ;
        RECT 37.680 149.025 37.850 149.215 ;
        RECT 38.020 149.190 38.275 149.765 ;
        RECT 37.680 148.695 37.935 149.025 ;
        RECT 35.215 148.335 35.800 148.525 ;
        RECT 24.165 147.385 29.510 147.820 ;
        RECT 29.685 147.385 35.030 147.820 ;
        RECT 35.215 147.565 35.490 148.335 ;
        RECT 35.970 148.165 36.865 148.495 ;
        RECT 37.680 148.485 37.850 148.695 ;
        RECT 35.660 147.995 36.865 148.165 ;
        RECT 35.660 147.565 35.990 147.995 ;
        RECT 36.160 147.385 36.355 147.825 ;
        RECT 36.535 147.565 36.865 147.995 ;
        RECT 37.135 148.315 37.850 148.485 ;
        RECT 38.105 148.460 38.275 149.190 ;
        RECT 38.450 149.095 38.710 149.935 ;
        RECT 38.885 149.165 42.395 149.935 ;
        RECT 42.565 149.185 43.775 149.935 ;
        RECT 43.945 149.210 44.235 149.935 ;
        RECT 44.405 149.390 49.750 149.935 ;
        RECT 38.885 148.645 40.535 149.165 ;
        RECT 37.135 147.555 37.305 148.315 ;
        RECT 37.520 147.385 37.850 148.145 ;
        RECT 38.020 147.555 38.275 148.460 ;
        RECT 38.450 147.385 38.710 148.535 ;
        RECT 40.705 148.475 42.395 148.995 ;
        RECT 42.565 148.645 43.085 149.185 ;
        RECT 43.255 148.475 43.775 149.015 ;
        RECT 45.990 148.560 46.330 149.390 ;
        RECT 50.385 149.350 50.695 149.765 ;
        RECT 50.890 149.555 51.220 149.935 ;
        RECT 51.390 149.595 52.795 149.765 ;
        RECT 51.390 149.365 51.560 149.595 ;
        RECT 38.885 147.385 42.395 148.475 ;
        RECT 42.565 147.385 43.775 148.475 ;
        RECT 43.945 147.385 44.235 148.550 ;
        RECT 47.810 147.820 48.160 149.070 ;
        RECT 50.385 148.235 50.555 149.350 ;
        RECT 50.865 149.195 51.560 149.365 ;
        RECT 52.625 149.365 52.795 149.595 ;
        RECT 53.065 149.535 53.395 149.935 ;
        RECT 53.635 149.365 53.805 149.765 ;
        RECT 50.865 149.025 51.035 149.195 ;
        RECT 50.725 148.695 51.035 149.025 ;
        RECT 51.205 148.695 51.540 149.025 ;
        RECT 51.810 148.695 52.005 149.270 ;
        RECT 52.265 149.025 52.455 149.255 ;
        RECT 52.625 149.195 53.805 149.365 ;
        RECT 54.100 149.195 54.715 149.765 ;
        RECT 54.885 149.425 55.100 149.935 ;
        RECT 55.330 149.425 55.610 149.755 ;
        RECT 55.790 149.425 56.030 149.935 ;
        RECT 52.265 148.695 52.610 149.025 ;
        RECT 52.920 148.695 53.395 149.025 ;
        RECT 53.650 148.695 53.835 149.025 ;
        RECT 50.865 148.525 51.035 148.695 ;
        RECT 50.865 148.355 53.805 148.525 ;
        RECT 44.405 147.385 49.750 147.820 ;
        RECT 50.385 147.595 50.725 148.235 ;
        RECT 51.315 148.015 52.875 148.185 ;
        RECT 50.895 147.385 51.140 147.845 ;
        RECT 51.315 147.555 51.565 148.015 ;
        RECT 51.755 147.385 52.425 147.765 ;
        RECT 52.625 147.555 52.875 148.015 ;
        RECT 53.635 147.555 53.805 148.355 ;
        RECT 54.100 148.175 54.415 149.195 ;
        RECT 54.585 148.525 54.755 149.025 ;
        RECT 55.005 148.695 55.270 149.255 ;
        RECT 55.440 148.525 55.610 149.425 ;
        RECT 55.780 148.695 56.135 149.255 ;
        RECT 56.385 149.125 56.625 149.935 ;
        RECT 56.795 149.125 57.125 149.765 ;
        RECT 57.295 149.125 57.565 149.935 ;
        RECT 56.365 148.695 56.715 148.945 ;
        RECT 56.885 148.525 57.055 149.125 ;
        RECT 57.225 148.695 57.575 148.945 ;
        RECT 54.585 148.355 56.010 148.525 ;
        RECT 54.100 147.555 54.635 148.175 ;
        RECT 54.805 147.385 55.135 148.185 ;
        RECT 55.620 148.180 56.010 148.355 ;
        RECT 56.375 148.355 57.055 148.525 ;
        RECT 56.375 147.570 56.705 148.355 ;
        RECT 57.235 147.385 57.565 148.525 ;
        RECT 57.745 147.555 58.025 149.655 ;
        RECT 58.255 149.475 58.425 149.935 ;
        RECT 58.695 149.545 59.945 149.725 ;
        RECT 59.080 149.305 59.445 149.375 ;
        RECT 58.195 149.125 59.445 149.305 ;
        RECT 59.615 149.325 59.945 149.545 ;
        RECT 60.115 149.495 60.285 149.935 ;
        RECT 60.455 149.325 60.795 149.740 ;
        RECT 59.615 149.155 60.795 149.325 ;
        RECT 60.965 149.135 61.275 149.935 ;
        RECT 61.480 149.135 62.175 149.765 ;
        RECT 62.345 149.390 67.690 149.935 ;
        RECT 58.195 148.525 58.470 149.125 ;
        RECT 58.640 148.695 58.995 148.945 ;
        RECT 59.190 148.915 59.655 148.945 ;
        RECT 59.185 148.745 59.655 148.915 ;
        RECT 59.190 148.695 59.655 148.745 ;
        RECT 59.825 148.695 60.155 148.945 ;
        RECT 60.330 148.745 60.795 148.945 ;
        RECT 60.975 148.695 61.310 148.965 ;
        RECT 59.975 148.575 60.155 148.695 ;
        RECT 58.195 148.315 59.805 148.525 ;
        RECT 59.975 148.405 60.305 148.575 ;
        RECT 59.395 148.215 59.805 148.315 ;
        RECT 58.215 147.385 59.000 148.145 ;
        RECT 59.395 147.555 59.780 148.215 ;
        RECT 60.105 147.615 60.305 148.405 ;
        RECT 60.475 147.385 60.795 148.565 ;
        RECT 61.480 148.535 61.650 149.135 ;
        RECT 61.820 148.695 62.155 148.945 ;
        RECT 63.930 148.560 64.270 149.390 ;
        RECT 67.875 149.205 68.175 149.935 ;
        RECT 60.965 147.385 61.245 148.525 ;
        RECT 61.415 147.555 61.745 148.535 ;
        RECT 61.915 147.385 62.175 148.525 ;
        RECT 65.750 147.820 66.100 149.070 ;
        RECT 68.355 149.025 68.585 149.645 ;
        RECT 68.785 149.375 69.010 149.755 ;
        RECT 69.180 149.545 69.510 149.935 ;
        RECT 68.785 149.195 69.115 149.375 ;
        RECT 67.880 148.695 68.175 149.025 ;
        RECT 68.355 148.695 68.770 149.025 ;
        RECT 68.940 148.525 69.115 149.195 ;
        RECT 69.285 148.695 69.525 149.345 ;
        RECT 69.705 149.210 69.995 149.935 ;
        RECT 70.165 149.390 75.510 149.935 ;
        RECT 75.685 149.390 81.030 149.935 ;
        RECT 81.205 149.390 86.550 149.935 ;
        RECT 71.750 148.560 72.090 149.390 ;
        RECT 67.875 148.165 68.770 148.495 ;
        RECT 68.940 148.335 69.525 148.525 ;
        RECT 67.875 147.995 69.080 148.165 ;
        RECT 62.345 147.385 67.690 147.820 ;
        RECT 67.875 147.565 68.205 147.995 ;
        RECT 68.385 147.385 68.580 147.825 ;
        RECT 68.750 147.565 69.080 147.995 ;
        RECT 69.250 147.565 69.525 148.335 ;
        RECT 69.705 147.385 69.995 148.550 ;
        RECT 73.570 147.820 73.920 149.070 ;
        RECT 77.270 148.560 77.610 149.390 ;
        RECT 79.090 147.820 79.440 149.070 ;
        RECT 82.790 148.560 83.130 149.390 ;
        RECT 86.725 149.260 86.985 149.765 ;
        RECT 87.165 149.555 87.495 149.935 ;
        RECT 87.675 149.385 87.845 149.765 ;
        RECT 84.610 147.820 84.960 149.070 ;
        RECT 86.725 148.460 86.895 149.260 ;
        RECT 87.180 149.215 87.845 149.385 ;
        RECT 87.180 148.960 87.350 149.215 ;
        RECT 88.105 149.185 89.315 149.935 ;
        RECT 87.065 148.630 87.350 148.960 ;
        RECT 87.585 148.665 87.915 149.035 ;
        RECT 87.180 148.485 87.350 148.630 ;
        RECT 70.165 147.385 75.510 147.820 ;
        RECT 75.685 147.385 81.030 147.820 ;
        RECT 81.205 147.385 86.550 147.820 ;
        RECT 86.725 147.555 86.995 148.460 ;
        RECT 87.180 148.315 87.845 148.485 ;
        RECT 87.165 147.385 87.495 148.145 ;
        RECT 87.675 147.555 87.845 148.315 ;
        RECT 88.105 148.475 88.625 149.015 ;
        RECT 88.795 148.645 89.315 149.185 ;
        RECT 88.105 147.385 89.315 148.475 ;
        RECT 18.100 147.215 89.400 147.385 ;
        RECT 18.185 146.125 19.395 147.215 ;
        RECT 19.565 146.780 24.910 147.215 ;
        RECT 25.085 146.780 30.430 147.215 ;
        RECT 18.185 145.415 18.705 145.955 ;
        RECT 18.875 145.585 19.395 146.125 ;
        RECT 18.185 144.665 19.395 145.415 ;
        RECT 21.150 145.210 21.490 146.040 ;
        RECT 22.970 145.530 23.320 146.780 ;
        RECT 26.670 145.210 27.010 146.040 ;
        RECT 28.490 145.530 28.840 146.780 ;
        RECT 31.065 146.050 31.355 147.215 ;
        RECT 31.525 146.125 33.195 147.215 ;
        RECT 31.525 145.435 32.275 145.955 ;
        RECT 32.445 145.605 33.195 146.125 ;
        RECT 33.825 146.075 34.105 147.215 ;
        RECT 34.275 146.065 34.605 147.045 ;
        RECT 34.775 146.075 35.035 147.215 ;
        RECT 35.210 146.375 35.530 147.215 ;
        RECT 35.700 146.195 35.900 146.985 ;
        RECT 36.225 146.285 36.610 147.045 ;
        RECT 37.005 146.455 37.805 147.215 ;
        RECT 34.340 146.025 34.515 146.065 ;
        RECT 33.835 145.635 34.170 145.905 ;
        RECT 34.340 145.465 34.510 146.025 ;
        RECT 34.680 145.655 35.015 145.905 ;
        RECT 35.210 145.855 35.530 146.195 ;
        RECT 35.700 146.025 36.055 146.195 ;
        RECT 36.225 146.075 37.825 146.285 ;
        RECT 35.875 145.905 36.055 146.025 ;
        RECT 35.210 145.655 35.705 145.855 ;
        RECT 35.875 145.655 36.205 145.905 ;
        RECT 36.375 145.655 36.840 145.905 ;
        RECT 37.010 145.655 37.365 145.905 ;
        RECT 37.545 145.475 37.825 146.075 ;
        RECT 19.565 144.665 24.910 145.210 ;
        RECT 25.085 144.665 30.430 145.210 ;
        RECT 31.065 144.665 31.355 145.390 ;
        RECT 31.525 144.665 33.195 145.435 ;
        RECT 33.825 144.665 34.135 145.465 ;
        RECT 34.340 144.835 35.035 145.465 ;
        RECT 35.210 145.405 36.240 145.445 ;
        RECT 35.210 145.275 36.410 145.405 ;
        RECT 35.210 144.860 35.545 145.275 ;
        RECT 35.715 144.665 35.885 145.105 ;
        RECT 36.070 145.055 36.410 145.275 ;
        RECT 36.585 145.295 37.825 145.475 ;
        RECT 36.585 145.225 36.950 145.295 ;
        RECT 36.070 144.875 37.335 145.055 ;
        RECT 37.595 144.665 37.775 145.125 ;
        RECT 37.995 144.945 38.210 147.045 ;
        RECT 38.435 146.025 38.685 147.215 ;
        RECT 38.885 146.075 39.270 147.035 ;
        RECT 39.485 146.415 39.775 147.215 ;
        RECT 39.945 146.875 41.310 147.045 ;
        RECT 39.945 146.245 40.115 146.875 ;
        RECT 39.440 146.075 40.115 146.245 ;
        RECT 38.445 144.665 38.615 145.465 ;
        RECT 38.885 145.405 39.060 146.075 ;
        RECT 39.440 145.905 39.610 146.075 ;
        RECT 40.285 145.905 40.610 146.705 ;
        RECT 40.980 146.665 41.310 146.875 ;
        RECT 40.980 146.415 41.935 146.665 ;
        RECT 39.245 145.655 39.610 145.905 ;
        RECT 39.805 145.655 40.055 145.905 ;
        RECT 39.245 145.575 39.435 145.655 ;
        RECT 39.805 145.575 39.975 145.655 ;
        RECT 40.265 145.575 40.610 145.905 ;
        RECT 40.780 145.575 41.055 146.240 ;
        RECT 41.240 145.575 41.595 146.240 ;
        RECT 41.765 145.405 41.935 146.415 ;
        RECT 42.105 146.075 42.395 147.215 ;
        RECT 42.565 146.125 45.155 147.215 ;
        RECT 42.120 145.575 42.395 145.905 ;
        RECT 38.885 144.835 39.395 145.405 ;
        RECT 39.940 145.235 41.340 145.405 ;
        RECT 39.565 144.665 39.735 145.225 ;
        RECT 39.940 144.835 40.270 145.235 ;
        RECT 40.445 144.665 40.775 145.065 ;
        RECT 41.010 145.045 41.340 145.235 ;
        RECT 41.510 145.215 41.935 145.405 ;
        RECT 42.565 145.435 43.775 145.955 ;
        RECT 43.945 145.605 45.155 146.125 ;
        RECT 45.325 146.075 45.655 147.215 ;
        RECT 45.825 146.585 46.180 147.045 ;
        RECT 46.350 146.755 46.925 147.215 ;
        RECT 47.095 146.585 47.425 147.045 ;
        RECT 45.825 146.415 47.425 146.585 ;
        RECT 47.625 146.415 47.880 147.215 ;
        RECT 48.545 146.780 53.890 147.215 ;
        RECT 45.825 146.075 46.100 146.415 ;
        RECT 46.280 145.855 46.470 146.235 ;
        RECT 45.325 145.655 46.470 145.855 ;
        RECT 46.650 145.485 46.930 146.415 ;
        RECT 48.050 146.245 48.350 146.440 ;
        RECT 47.100 146.075 48.350 146.245 ;
        RECT 47.100 145.655 47.430 146.075 ;
        RECT 47.660 145.575 48.005 145.905 ;
        RECT 42.105 145.045 42.395 145.315 ;
        RECT 41.010 144.835 42.395 145.045 ;
        RECT 42.565 144.665 45.155 145.435 ;
        RECT 45.325 145.275 46.435 145.485 ;
        RECT 45.325 144.835 45.675 145.275 ;
        RECT 45.845 144.665 46.015 145.105 ;
        RECT 46.185 145.045 46.435 145.275 ;
        RECT 46.605 145.385 46.930 145.485 ;
        RECT 46.605 145.215 46.935 145.385 ;
        RECT 47.105 145.045 47.380 145.485 ;
        RECT 48.180 145.420 48.350 146.075 ;
        RECT 46.185 144.835 47.380 145.045 ;
        RECT 47.615 144.665 47.945 145.405 ;
        RECT 48.115 145.090 48.350 145.420 ;
        RECT 50.130 145.210 50.470 146.040 ;
        RECT 51.950 145.530 52.300 146.780 ;
        RECT 54.065 146.125 56.655 147.215 ;
        RECT 54.065 145.435 55.275 145.955 ;
        RECT 55.445 145.605 56.655 146.125 ;
        RECT 56.825 146.050 57.115 147.215 ;
        RECT 57.745 146.615 58.005 147.035 ;
        RECT 58.175 146.785 58.505 147.215 ;
        RECT 59.170 146.785 59.915 146.955 ;
        RECT 60.140 146.875 60.780 147.035 ;
        RECT 57.745 146.445 59.575 146.615 ;
        RECT 48.545 144.665 53.890 145.210 ;
        RECT 54.065 144.665 56.655 145.435 ;
        RECT 57.745 145.405 57.915 146.445 ;
        RECT 58.085 145.575 58.435 146.275 ;
        RECT 58.650 146.105 59.235 146.275 ;
        RECT 58.605 145.575 58.895 145.905 ;
        RECT 59.065 145.825 59.235 146.105 ;
        RECT 59.405 146.165 59.575 146.445 ;
        RECT 59.745 146.535 59.915 146.785 ;
        RECT 60.105 146.705 60.780 146.875 ;
        RECT 59.745 146.365 60.780 146.535 ;
        RECT 60.950 146.415 61.230 147.215 ;
        RECT 60.610 146.245 60.780 146.365 ;
        RECT 59.405 145.995 60.055 146.165 ;
        RECT 60.610 146.075 61.270 146.245 ;
        RECT 61.440 146.075 61.715 147.045 ;
        RECT 61.975 146.285 62.145 147.045 ;
        RECT 62.360 146.455 62.690 147.215 ;
        RECT 61.975 146.115 62.690 146.285 ;
        RECT 62.860 146.140 63.115 147.045 ;
        RECT 59.065 145.655 59.490 145.825 ;
        RECT 59.065 145.405 59.235 145.655 ;
        RECT 59.885 145.575 60.055 145.995 ;
        RECT 61.100 145.905 61.270 146.075 ;
        RECT 60.275 145.575 60.930 145.905 ;
        RECT 61.100 145.575 61.375 145.905 ;
        RECT 61.100 145.405 61.270 145.575 ;
        RECT 56.825 144.665 57.115 145.390 ;
        RECT 57.745 145.030 58.060 145.405 ;
        RECT 58.315 144.665 58.485 145.405 ;
        RECT 58.735 145.235 59.235 145.405 ;
        RECT 59.675 145.235 61.270 145.405 ;
        RECT 61.545 145.340 61.715 146.075 ;
        RECT 61.885 145.565 62.240 145.935 ;
        RECT 62.520 145.905 62.690 146.115 ;
        RECT 62.520 145.575 62.775 145.905 ;
        RECT 62.520 145.385 62.690 145.575 ;
        RECT 62.945 145.410 63.115 146.140 ;
        RECT 63.290 146.065 63.550 147.215 ;
        RECT 63.730 146.645 64.050 147.045 ;
        RECT 63.730 146.195 63.900 146.645 ;
        RECT 64.220 146.415 64.530 147.215 ;
        RECT 64.700 146.585 65.030 147.045 ;
        RECT 65.200 146.755 65.370 147.215 ;
        RECT 65.540 146.585 65.870 147.045 ;
        RECT 66.040 146.755 66.290 147.215 ;
        RECT 66.480 146.755 66.730 147.215 ;
        RECT 64.700 146.535 65.870 146.585 ;
        RECT 66.900 146.585 67.150 147.045 ;
        RECT 67.400 146.755 67.690 147.215 ;
        RECT 67.865 146.780 73.210 147.215 ;
        RECT 73.385 146.780 78.730 147.215 ;
        RECT 66.900 146.535 67.690 146.585 ;
        RECT 64.700 146.365 67.690 146.535 ;
        RECT 63.730 146.025 67.290 146.195 ;
        RECT 58.735 145.030 58.905 145.235 ;
        RECT 59.130 144.665 59.505 145.065 ;
        RECT 59.675 144.885 59.845 145.235 ;
        RECT 60.030 144.665 60.360 145.065 ;
        RECT 60.530 144.885 60.700 145.235 ;
        RECT 60.870 144.665 61.250 145.065 ;
        RECT 61.440 144.995 61.715 145.340 ;
        RECT 61.975 145.215 62.690 145.385 ;
        RECT 61.975 144.835 62.145 145.215 ;
        RECT 62.360 144.665 62.690 145.045 ;
        RECT 62.860 144.835 63.115 145.410 ;
        RECT 63.290 144.665 63.550 145.505 ;
        RECT 63.730 145.235 63.900 146.025 ;
        RECT 64.070 145.655 64.420 145.855 ;
        RECT 64.700 145.655 65.380 145.855 ;
        RECT 65.590 145.655 66.780 145.855 ;
        RECT 66.960 145.655 67.290 146.025 ;
        RECT 67.490 145.485 67.690 146.365 ;
        RECT 63.730 144.835 64.050 145.235 ;
        RECT 64.220 144.665 64.530 145.485 ;
        RECT 64.700 145.295 66.390 145.485 ;
        RECT 64.700 144.835 65.030 145.295 ;
        RECT 65.640 145.215 66.390 145.295 ;
        RECT 65.200 144.665 65.450 145.125 ;
        RECT 66.560 145.045 66.730 145.485 ;
        RECT 66.900 145.215 67.690 145.485 ;
        RECT 69.450 145.210 69.790 146.040 ;
        RECT 71.270 145.530 71.620 146.780 ;
        RECT 74.970 145.210 75.310 146.040 ;
        RECT 76.790 145.530 77.140 146.780 ;
        RECT 78.905 146.125 82.415 147.215 ;
        RECT 78.905 145.435 80.555 145.955 ;
        RECT 80.725 145.605 82.415 146.125 ;
        RECT 82.585 146.050 82.875 147.215 ;
        RECT 83.045 146.125 85.635 147.215 ;
        RECT 86.270 146.790 86.605 147.215 ;
        RECT 86.775 146.610 86.960 147.015 ;
        RECT 83.045 145.435 84.255 145.955 ;
        RECT 84.425 145.605 85.635 146.125 ;
        RECT 86.295 146.435 86.960 146.610 ;
        RECT 87.165 146.435 87.495 147.215 ;
        RECT 65.640 144.835 67.690 145.045 ;
        RECT 67.865 144.665 73.210 145.210 ;
        RECT 73.385 144.665 78.730 145.210 ;
        RECT 78.905 144.665 82.415 145.435 ;
        RECT 82.585 144.665 82.875 145.390 ;
        RECT 83.045 144.665 85.635 145.435 ;
        RECT 86.295 145.405 86.635 146.435 ;
        RECT 87.665 146.245 87.935 147.015 ;
        RECT 86.805 146.075 87.935 146.245 ;
        RECT 86.805 145.575 87.055 146.075 ;
        RECT 86.295 145.235 86.980 145.405 ;
        RECT 87.235 145.325 87.595 145.905 ;
        RECT 86.270 144.665 86.605 145.065 ;
        RECT 86.775 144.835 86.980 145.235 ;
        RECT 87.765 145.165 87.935 146.075 ;
        RECT 88.105 146.125 89.315 147.215 ;
        RECT 88.105 145.585 88.625 146.125 ;
        RECT 88.795 145.415 89.315 145.955 ;
        RECT 87.190 144.665 87.465 145.145 ;
        RECT 87.675 144.835 87.935 145.165 ;
        RECT 88.105 144.665 89.315 145.415 ;
        RECT 18.100 144.495 89.400 144.665 ;
        RECT 18.185 143.745 19.395 144.495 ;
        RECT 19.565 143.950 24.910 144.495 ;
        RECT 25.085 143.950 30.430 144.495 ;
        RECT 30.605 143.950 35.950 144.495 ;
        RECT 36.215 144.155 36.385 144.190 ;
        RECT 36.185 143.985 36.385 144.155 ;
        RECT 18.185 143.205 18.705 143.745 ;
        RECT 18.875 143.035 19.395 143.575 ;
        RECT 21.150 143.120 21.490 143.950 ;
        RECT 18.185 141.945 19.395 143.035 ;
        RECT 22.970 142.380 23.320 143.630 ;
        RECT 26.670 143.120 27.010 143.950 ;
        RECT 28.490 142.380 28.840 143.630 ;
        RECT 32.190 143.120 32.530 143.950 ;
        RECT 34.010 142.380 34.360 143.630 ;
        RECT 36.215 143.625 36.385 143.985 ;
        RECT 36.575 143.965 36.805 144.270 ;
        RECT 36.975 144.135 37.305 144.495 ;
        RECT 37.500 143.965 37.790 144.315 ;
        RECT 36.575 143.795 37.790 143.965 ;
        RECT 37.965 144.035 38.525 144.325 ;
        RECT 38.695 144.035 38.945 144.495 ;
        RECT 36.215 143.455 36.735 143.625 ;
        RECT 36.130 142.925 36.375 143.285 ;
        RECT 36.565 143.075 36.735 143.455 ;
        RECT 36.905 143.255 37.290 143.585 ;
        RECT 37.470 143.475 37.730 143.585 ;
        RECT 37.470 143.305 37.735 143.475 ;
        RECT 37.470 143.255 37.730 143.305 ;
        RECT 36.565 142.795 36.915 143.075 ;
        RECT 19.565 141.945 24.910 142.380 ;
        RECT 25.085 141.945 30.430 142.380 ;
        RECT 30.605 141.945 35.950 142.380 ;
        RECT 36.130 141.945 36.385 142.745 ;
        RECT 36.585 142.115 36.915 142.795 ;
        RECT 37.095 142.205 37.290 143.255 ;
        RECT 37.470 141.945 37.790 143.085 ;
        RECT 37.965 142.665 38.215 144.035 ;
        RECT 39.565 143.865 39.895 144.225 ;
        RECT 41.205 143.985 41.445 144.495 ;
        RECT 41.615 143.985 41.905 144.325 ;
        RECT 42.135 143.985 42.450 144.495 ;
        RECT 38.505 143.675 39.895 143.865 ;
        RECT 38.505 143.585 38.675 143.675 ;
        RECT 38.385 143.255 38.675 143.585 ;
        RECT 38.845 143.255 39.185 143.505 ;
        RECT 39.405 143.255 40.080 143.505 ;
        RECT 41.250 143.475 41.445 143.815 ;
        RECT 41.245 143.305 41.445 143.475 ;
        RECT 41.250 143.255 41.445 143.305 ;
        RECT 38.505 143.005 38.675 143.255 ;
        RECT 38.505 142.835 39.445 143.005 ;
        RECT 39.815 142.895 40.080 143.255 ;
        RECT 41.615 143.085 41.795 143.985 ;
        RECT 42.620 143.925 42.790 144.195 ;
        RECT 42.960 144.095 43.290 144.495 ;
        RECT 41.965 143.255 42.375 143.815 ;
        RECT 42.620 143.755 43.315 143.925 ;
        RECT 43.945 143.770 44.235 144.495 ;
        RECT 44.410 144.095 44.745 144.495 ;
        RECT 44.915 143.925 45.120 144.325 ;
        RECT 45.330 144.015 45.605 144.495 ;
        RECT 45.815 143.995 46.075 144.325 ;
        RECT 42.545 143.085 42.715 143.585 ;
        RECT 41.255 142.915 42.715 143.085 ;
        RECT 37.965 142.115 38.425 142.665 ;
        RECT 38.615 141.945 38.945 142.665 ;
        RECT 39.145 142.285 39.445 142.835 ;
        RECT 41.255 142.740 41.615 142.915 ;
        RECT 42.885 142.745 43.315 143.755 ;
        RECT 44.435 143.755 45.120 143.925 ;
        RECT 39.615 141.945 39.895 142.615 ;
        RECT 42.200 141.945 42.370 142.745 ;
        RECT 42.540 142.575 43.315 142.745 ;
        RECT 42.540 142.115 42.870 142.575 ;
        RECT 43.040 141.945 43.210 142.405 ;
        RECT 43.945 141.945 44.235 143.110 ;
        RECT 44.435 142.725 44.775 143.755 ;
        RECT 44.945 143.085 45.195 143.585 ;
        RECT 45.375 143.255 45.735 143.835 ;
        RECT 45.905 143.085 46.075 143.995 ;
        RECT 46.335 143.945 46.505 144.325 ;
        RECT 46.685 144.115 47.015 144.495 ;
        RECT 46.335 143.775 47.000 143.945 ;
        RECT 47.195 143.820 47.455 144.325 ;
        RECT 47.625 143.950 52.970 144.495 ;
        RECT 53.145 143.950 58.490 144.495 ;
        RECT 46.265 143.225 46.595 143.595 ;
        RECT 46.830 143.520 47.000 143.775 ;
        RECT 44.945 142.915 46.075 143.085 ;
        RECT 46.830 143.190 47.115 143.520 ;
        RECT 46.830 143.045 47.000 143.190 ;
        RECT 44.435 142.550 45.100 142.725 ;
        RECT 44.410 141.945 44.745 142.370 ;
        RECT 44.915 142.145 45.100 142.550 ;
        RECT 45.305 141.945 45.635 142.725 ;
        RECT 45.805 142.145 46.075 142.915 ;
        RECT 46.335 142.875 47.000 143.045 ;
        RECT 47.285 143.020 47.455 143.820 ;
        RECT 49.210 143.120 49.550 143.950 ;
        RECT 46.335 142.115 46.505 142.875 ;
        RECT 46.685 141.945 47.015 142.705 ;
        RECT 47.185 142.115 47.455 143.020 ;
        RECT 51.030 142.380 51.380 143.630 ;
        RECT 54.730 143.120 55.070 143.950 ;
        RECT 58.665 143.725 62.175 144.495 ;
        RECT 62.810 144.115 64.860 144.325 ;
        RECT 56.550 142.380 56.900 143.630 ;
        RECT 58.665 143.205 60.315 143.725 ;
        RECT 62.810 143.675 63.600 143.945 ;
        RECT 63.770 143.675 63.940 144.115 ;
        RECT 65.050 144.035 65.300 144.495 ;
        RECT 64.110 143.865 64.860 143.945 ;
        RECT 65.470 143.865 65.800 144.325 ;
        RECT 64.110 143.675 65.800 143.865 ;
        RECT 65.970 143.675 66.280 144.495 ;
        RECT 66.450 143.925 66.770 144.325 ;
        RECT 62.810 143.645 63.035 143.675 ;
        RECT 60.485 143.035 62.175 143.555 ;
        RECT 47.625 141.945 52.970 142.380 ;
        RECT 53.145 141.945 58.490 142.380 ;
        RECT 58.665 141.945 62.175 143.035 ;
        RECT 62.810 142.795 63.010 143.645 ;
        RECT 63.210 143.135 63.540 143.505 ;
        RECT 63.720 143.305 64.910 143.505 ;
        RECT 65.120 143.305 65.800 143.505 ;
        RECT 66.080 143.305 66.430 143.505 ;
        RECT 66.600 143.135 66.770 143.925 ;
        RECT 66.945 143.725 69.535 144.495 ;
        RECT 69.705 143.770 69.995 144.495 ;
        RECT 70.165 143.950 75.510 144.495 ;
        RECT 75.685 143.950 81.030 144.495 ;
        RECT 81.205 143.950 86.550 144.495 ;
        RECT 66.945 143.205 68.155 143.725 ;
        RECT 63.210 142.965 66.770 143.135 ;
        RECT 68.325 143.035 69.535 143.555 ;
        RECT 71.750 143.120 72.090 143.950 ;
        RECT 62.810 142.625 65.800 142.795 ;
        RECT 62.810 142.575 63.600 142.625 ;
        RECT 62.810 141.945 63.100 142.405 ;
        RECT 63.350 142.115 63.600 142.575 ;
        RECT 64.630 142.575 65.800 142.625 ;
        RECT 63.770 141.945 64.020 142.405 ;
        RECT 64.210 141.945 64.460 142.405 ;
        RECT 64.630 142.115 64.960 142.575 ;
        RECT 65.130 141.945 65.300 142.405 ;
        RECT 65.470 142.115 65.800 142.575 ;
        RECT 65.970 141.945 66.280 142.745 ;
        RECT 66.600 142.515 66.770 142.965 ;
        RECT 66.450 142.115 66.770 142.515 ;
        RECT 66.945 141.945 69.535 143.035 ;
        RECT 69.705 141.945 69.995 143.110 ;
        RECT 73.570 142.380 73.920 143.630 ;
        RECT 77.270 143.120 77.610 143.950 ;
        RECT 79.090 142.380 79.440 143.630 ;
        RECT 82.790 143.120 83.130 143.950 ;
        RECT 86.905 143.835 87.245 144.495 ;
        RECT 84.610 142.380 84.960 143.630 ;
        RECT 70.165 141.945 75.510 142.380 ;
        RECT 75.685 141.945 81.030 142.380 ;
        RECT 81.205 141.945 86.550 142.380 ;
        RECT 86.725 142.115 87.245 143.665 ;
        RECT 87.415 142.840 87.935 144.325 ;
        RECT 88.105 143.745 89.315 144.495 ;
        RECT 88.105 143.035 88.625 143.575 ;
        RECT 88.795 143.205 89.315 143.745 ;
        RECT 87.415 141.945 87.745 142.670 ;
        RECT 88.105 141.945 89.315 143.035 ;
        RECT 18.100 141.775 89.400 141.945 ;
        RECT 18.185 140.685 19.395 141.775 ;
        RECT 19.565 141.340 24.910 141.775 ;
        RECT 18.185 139.975 18.705 140.515 ;
        RECT 18.875 140.145 19.395 140.685 ;
        RECT 18.185 139.225 19.395 139.975 ;
        RECT 21.150 139.770 21.490 140.600 ;
        RECT 22.970 140.090 23.320 141.340 ;
        RECT 26.005 140.055 26.525 141.605 ;
        RECT 26.695 141.050 27.025 141.775 ;
        RECT 19.565 139.225 24.910 139.770 ;
        RECT 26.185 139.225 26.525 139.885 ;
        RECT 26.695 139.395 27.215 140.880 ;
        RECT 27.385 140.685 30.895 141.775 ;
        RECT 27.385 139.995 29.035 140.515 ;
        RECT 29.205 140.165 30.895 140.685 ;
        RECT 31.065 140.610 31.355 141.775 ;
        RECT 31.525 140.685 35.035 141.775 ;
        RECT 31.525 139.995 33.175 140.515 ;
        RECT 33.345 140.165 35.035 140.685 ;
        RECT 35.665 140.700 35.935 141.605 ;
        RECT 36.105 141.015 36.435 141.775 ;
        RECT 36.615 140.845 36.785 141.605 ;
        RECT 27.385 139.225 30.895 139.995 ;
        RECT 31.065 139.225 31.355 139.950 ;
        RECT 31.525 139.225 35.035 139.995 ;
        RECT 35.665 139.900 35.835 140.700 ;
        RECT 36.120 140.675 36.785 140.845 ;
        RECT 37.045 140.685 38.715 141.775 ;
        RECT 36.120 140.530 36.290 140.675 ;
        RECT 36.005 140.200 36.290 140.530 ;
        RECT 36.120 139.945 36.290 140.200 ;
        RECT 36.525 140.125 36.855 140.495 ;
        RECT 37.045 139.995 37.795 140.515 ;
        RECT 37.965 140.165 38.715 140.685 ;
        RECT 38.975 140.845 39.145 141.605 ;
        RECT 39.360 141.015 39.690 141.775 ;
        RECT 38.975 140.675 39.690 140.845 ;
        RECT 39.860 140.700 40.115 141.605 ;
        RECT 38.885 140.125 39.240 140.495 ;
        RECT 39.520 140.465 39.690 140.675 ;
        RECT 39.520 140.135 39.775 140.465 ;
        RECT 35.665 139.395 35.925 139.900 ;
        RECT 36.120 139.775 36.785 139.945 ;
        RECT 36.105 139.225 36.435 139.605 ;
        RECT 36.615 139.395 36.785 139.775 ;
        RECT 37.045 139.225 38.715 139.995 ;
        RECT 39.520 139.945 39.690 140.135 ;
        RECT 39.945 139.970 40.115 140.700 ;
        RECT 40.290 140.625 40.550 141.775 ;
        RECT 40.725 140.635 40.985 141.775 ;
        RECT 41.155 140.625 41.485 141.605 ;
        RECT 41.655 140.635 41.935 141.775 ;
        RECT 42.185 140.845 42.365 141.605 ;
        RECT 42.545 141.015 42.875 141.775 ;
        RECT 42.185 140.675 42.860 140.845 ;
        RECT 43.045 140.700 43.315 141.605 ;
        RECT 40.745 140.215 41.080 140.465 ;
        RECT 38.975 139.775 39.690 139.945 ;
        RECT 38.975 139.395 39.145 139.775 ;
        RECT 39.360 139.225 39.690 139.605 ;
        RECT 39.860 139.395 40.115 139.970 ;
        RECT 40.290 139.225 40.550 140.065 ;
        RECT 41.250 140.025 41.420 140.625 ;
        RECT 42.690 140.530 42.860 140.675 ;
        RECT 41.590 140.195 41.925 140.465 ;
        RECT 42.125 140.125 42.465 140.495 ;
        RECT 42.690 140.200 42.965 140.530 ;
        RECT 40.725 139.395 41.420 140.025 ;
        RECT 41.625 139.225 41.935 140.025 ;
        RECT 42.690 139.945 42.860 140.200 ;
        RECT 42.195 139.775 42.860 139.945 ;
        RECT 43.135 139.900 43.315 140.700 ;
        RECT 43.945 140.610 44.235 141.775 ;
        RECT 45.325 140.805 45.595 141.575 ;
        RECT 45.765 140.995 46.095 141.775 ;
        RECT 46.300 141.170 46.485 141.575 ;
        RECT 46.655 141.350 46.990 141.775 ;
        RECT 46.300 140.995 46.965 141.170 ;
        RECT 45.325 140.635 46.455 140.805 ;
        RECT 42.195 139.395 42.365 139.775 ;
        RECT 42.545 139.225 42.875 139.605 ;
        RECT 43.055 139.395 43.315 139.900 ;
        RECT 43.945 139.225 44.235 139.950 ;
        RECT 45.325 139.725 45.495 140.635 ;
        RECT 45.665 139.885 46.025 140.465 ;
        RECT 46.205 140.135 46.455 140.635 ;
        RECT 46.625 139.965 46.965 140.995 ;
        RECT 47.165 140.685 48.375 141.775 ;
        RECT 46.280 139.795 46.965 139.965 ;
        RECT 47.165 139.975 47.685 140.515 ;
        RECT 47.855 140.145 48.375 140.685 ;
        RECT 48.635 140.845 48.805 141.605 ;
        RECT 49.020 141.015 49.350 141.775 ;
        RECT 48.635 140.675 49.350 140.845 ;
        RECT 49.520 140.700 49.775 141.605 ;
        RECT 48.545 140.125 48.900 140.495 ;
        RECT 49.180 140.465 49.350 140.675 ;
        RECT 49.180 140.135 49.435 140.465 ;
        RECT 45.325 139.395 45.585 139.725 ;
        RECT 45.795 139.225 46.070 139.705 ;
        RECT 46.280 139.395 46.485 139.795 ;
        RECT 46.655 139.225 46.990 139.625 ;
        RECT 47.165 139.225 48.375 139.975 ;
        RECT 49.180 139.945 49.350 140.135 ;
        RECT 49.605 139.970 49.775 140.700 ;
        RECT 49.950 140.625 50.210 141.775 ;
        RECT 50.385 141.340 55.730 141.775 ;
        RECT 48.635 139.775 49.350 139.945 ;
        RECT 48.635 139.395 48.805 139.775 ;
        RECT 49.020 139.225 49.350 139.605 ;
        RECT 49.520 139.395 49.775 139.970 ;
        RECT 49.950 139.225 50.210 140.065 ;
        RECT 51.970 139.770 52.310 140.600 ;
        RECT 53.790 140.090 54.140 141.340 ;
        RECT 56.825 140.610 57.115 141.775 ;
        RECT 57.285 141.340 62.630 141.775 ;
        RECT 62.805 141.340 68.150 141.775 ;
        RECT 50.385 139.225 55.730 139.770 ;
        RECT 56.825 139.225 57.115 139.950 ;
        RECT 58.870 139.770 59.210 140.600 ;
        RECT 60.690 140.090 61.040 141.340 ;
        RECT 64.390 139.770 64.730 140.600 ;
        RECT 66.210 140.090 66.560 141.340 ;
        RECT 68.325 140.685 69.535 141.775 ;
        RECT 68.325 139.975 68.845 140.515 ;
        RECT 69.015 140.145 69.535 140.685 ;
        RECT 69.705 140.610 69.995 141.775 ;
        RECT 70.165 141.340 75.510 141.775 ;
        RECT 75.685 141.340 81.030 141.775 ;
        RECT 57.285 139.225 62.630 139.770 ;
        RECT 62.805 139.225 68.150 139.770 ;
        RECT 68.325 139.225 69.535 139.975 ;
        RECT 69.705 139.225 69.995 139.950 ;
        RECT 71.750 139.770 72.090 140.600 ;
        RECT 73.570 140.090 73.920 141.340 ;
        RECT 77.270 139.770 77.610 140.600 ;
        RECT 79.090 140.090 79.440 141.340 ;
        RECT 81.205 140.685 82.415 141.775 ;
        RECT 81.205 139.975 81.725 140.515 ;
        RECT 81.895 140.145 82.415 140.685 ;
        RECT 82.585 140.610 82.875 141.775 ;
        RECT 83.045 140.685 86.555 141.775 ;
        RECT 86.725 140.685 87.935 141.775 ;
        RECT 83.045 139.995 84.695 140.515 ;
        RECT 84.865 140.165 86.555 140.685 ;
        RECT 70.165 139.225 75.510 139.770 ;
        RECT 75.685 139.225 81.030 139.770 ;
        RECT 81.205 139.225 82.415 139.975 ;
        RECT 82.585 139.225 82.875 139.950 ;
        RECT 83.045 139.225 86.555 139.995 ;
        RECT 86.725 139.975 87.245 140.515 ;
        RECT 87.415 140.145 87.935 140.685 ;
        RECT 88.105 140.685 89.315 141.775 ;
        RECT 88.105 140.145 88.625 140.685 ;
        RECT 88.795 139.975 89.315 140.515 ;
        RECT 86.725 139.225 87.935 139.975 ;
        RECT 88.105 139.225 89.315 139.975 ;
        RECT 18.100 139.055 89.400 139.225 ;
      LAYER met1 ;
        RECT 21.850 214.180 22.170 214.240 ;
        RECT 41.630 214.180 41.950 214.240 ;
        RECT 21.850 214.040 41.950 214.180 ;
        RECT 21.850 213.980 22.170 214.040 ;
        RECT 41.630 213.980 41.950 214.040 ;
        RECT 24.610 213.160 24.930 213.220 ;
        RECT 80.270 213.160 80.590 213.220 ;
        RECT 24.610 213.020 80.590 213.160 ;
        RECT 24.610 212.960 24.930 213.020 ;
        RECT 80.270 212.960 80.590 213.020 ;
        RECT 26.450 212.820 26.770 212.880 ;
        RECT 32.430 212.820 32.750 212.880 ;
        RECT 81.650 212.820 81.970 212.880 ;
        RECT 26.450 212.680 81.970 212.820 ;
        RECT 26.450 212.620 26.770 212.680 ;
        RECT 32.430 212.620 32.750 212.680 ;
        RECT 81.650 212.620 81.970 212.680 ;
        RECT 25.070 212.480 25.390 212.540 ;
        RECT 54.510 212.480 54.830 212.540 ;
        RECT 25.070 212.340 54.830 212.480 ;
        RECT 25.070 212.280 25.390 212.340 ;
        RECT 54.510 212.280 54.830 212.340 ;
        RECT 19.550 212.140 19.870 212.200 ;
        RECT 31.970 212.140 32.290 212.200 ;
        RECT 19.550 212.000 32.290 212.140 ;
        RECT 19.550 211.940 19.870 212.000 ;
        RECT 31.970 211.940 32.290 212.000 ;
        RECT 36.570 212.140 36.890 212.200 ;
        RECT 59.110 212.140 59.430 212.200 ;
        RECT 36.570 212.000 59.430 212.140 ;
        RECT 36.570 211.940 36.890 212.000 ;
        RECT 59.110 211.940 59.430 212.000 ;
        RECT 16.790 211.460 17.110 211.520 ;
        RECT 22.310 211.460 22.630 211.520 ;
        RECT 16.790 211.320 22.630 211.460 ;
        RECT 16.790 211.260 17.110 211.320 ;
        RECT 22.310 211.260 22.630 211.320 ;
        RECT 35.190 211.460 35.510 211.520 ;
        RECT 42.090 211.460 42.410 211.520 ;
        RECT 35.190 211.320 42.410 211.460 ;
        RECT 35.190 211.260 35.510 211.320 ;
        RECT 42.090 211.260 42.410 211.320 ;
        RECT 59.570 211.460 59.890 211.520 ;
        RECT 82.570 211.460 82.890 211.520 ;
        RECT 59.570 211.320 82.890 211.460 ;
        RECT 59.570 211.260 59.890 211.320 ;
        RECT 82.570 211.260 82.890 211.320 ;
        RECT 29.670 211.120 29.990 211.180 ;
        RECT 61.410 211.120 61.730 211.180 ;
        RECT 29.670 210.980 61.730 211.120 ;
        RECT 29.670 210.920 29.990 210.980 ;
        RECT 61.410 210.920 61.730 210.980 ;
        RECT 31.050 210.780 31.370 210.840 ;
        RECT 71.530 210.780 71.850 210.840 ;
        RECT 31.050 210.640 71.850 210.780 ;
        RECT 31.050 210.580 31.370 210.640 ;
        RECT 71.530 210.580 71.850 210.640 ;
        RECT 24.150 210.440 24.470 210.500 ;
        RECT 41.630 210.440 41.950 210.500 ;
        RECT 24.150 210.300 41.950 210.440 ;
        RECT 24.150 210.240 24.470 210.300 ;
        RECT 41.630 210.240 41.950 210.300 ;
        RECT 18.100 209.620 89.400 210.100 ;
        RECT 21.850 209.220 22.170 209.480 ;
        RECT 25.070 209.220 25.390 209.480 ;
        RECT 29.210 209.420 29.530 209.480 ;
        RECT 62.790 209.420 63.110 209.480 ;
        RECT 67.390 209.420 67.710 209.480 ;
        RECT 26.080 209.280 29.530 209.420 ;
        RECT 20.025 209.080 20.315 209.125 ;
        RECT 26.080 209.080 26.220 209.280 ;
        RECT 29.210 209.220 29.530 209.280 ;
        RECT 32.520 209.280 67.710 209.420 ;
        RECT 20.025 208.940 21.160 209.080 ;
        RECT 20.025 208.895 20.315 208.940 ;
        RECT 21.020 208.800 21.160 208.940 ;
        RECT 24.240 208.940 26.220 209.080 ;
        RECT 20.485 208.555 20.775 208.785 ;
        RECT 20.560 208.400 20.700 208.555 ;
        RECT 20.930 208.540 21.250 208.800 ;
        RECT 24.240 208.785 24.380 208.940 ;
        RECT 26.450 208.880 26.770 209.140 ;
        RECT 24.165 208.555 24.455 208.785 ;
        RECT 25.990 208.540 26.310 208.800 ;
        RECT 27.370 208.540 27.690 208.800 ;
        RECT 29.670 208.540 29.990 208.800 ;
        RECT 30.590 208.540 30.910 208.800 ;
        RECT 32.520 208.785 32.660 209.280 ;
        RECT 62.790 209.220 63.110 209.280 ;
        RECT 67.390 209.220 67.710 209.280 ;
        RECT 67.940 209.280 74.750 209.420 ;
        RECT 37.030 209.080 37.350 209.140 ;
        RECT 45.325 209.080 45.615 209.125 ;
        RECT 33.440 208.940 45.615 209.080 ;
        RECT 33.440 208.785 33.580 208.940 ;
        RECT 37.030 208.880 37.350 208.940 ;
        RECT 45.325 208.895 45.615 208.940 ;
        RECT 54.065 209.080 54.355 209.125 ;
        RECT 56.810 209.080 57.130 209.140 ;
        RECT 54.065 208.940 57.130 209.080 ;
        RECT 54.065 208.895 54.355 208.940 ;
        RECT 56.810 208.880 57.130 208.940 ;
        RECT 66.010 209.080 66.330 209.140 ;
        RECT 67.940 209.080 68.080 209.280 ;
        RECT 66.010 208.940 68.080 209.080 ;
        RECT 71.530 209.080 71.850 209.140 ;
        RECT 73.370 209.080 73.690 209.140 ;
        RECT 71.530 208.940 73.690 209.080 ;
        RECT 74.610 209.080 74.750 209.280 ;
        RECT 81.650 209.220 81.970 209.480 ;
        RECT 74.610 208.940 85.100 209.080 ;
        RECT 66.010 208.880 66.330 208.940 ;
        RECT 71.530 208.880 71.850 208.940 ;
        RECT 73.370 208.880 73.690 208.940 ;
        RECT 32.445 208.555 32.735 208.785 ;
        RECT 33.365 208.555 33.655 208.785 ;
        RECT 34.745 208.555 35.035 208.785 ;
        RECT 36.570 208.740 36.890 208.800 ;
        RECT 37.505 208.740 37.795 208.785 ;
        RECT 36.570 208.600 37.795 208.740 ;
        RECT 31.050 208.400 31.370 208.460 ;
        RECT 20.560 208.260 31.370 208.400 ;
        RECT 31.050 208.200 31.370 208.260 ;
        RECT 31.970 208.400 32.290 208.460 ;
        RECT 31.970 208.260 33.580 208.400 ;
        RECT 31.970 208.200 32.290 208.260 ;
        RECT 23.245 208.060 23.535 208.105 ;
        RECT 31.510 208.060 31.830 208.120 ;
        RECT 23.245 207.920 31.830 208.060 ;
        RECT 23.245 207.875 23.535 207.920 ;
        RECT 31.510 207.860 31.830 207.920 ;
        RECT 32.890 207.860 33.210 208.120 ;
        RECT 33.440 208.060 33.580 208.260 ;
        RECT 33.810 208.200 34.130 208.460 ;
        RECT 34.820 208.060 34.960 208.555 ;
        RECT 36.570 208.540 36.890 208.600 ;
        RECT 37.505 208.555 37.795 208.600 ;
        RECT 37.950 208.540 38.270 208.800 ;
        RECT 38.410 208.540 38.730 208.800 ;
        RECT 39.790 208.540 40.110 208.800 ;
        RECT 40.545 208.555 40.835 208.785 ;
        RECT 35.190 208.400 35.510 208.460 ;
        RECT 38.870 208.400 39.190 208.460 ;
        RECT 35.190 208.260 39.190 208.400 ;
        RECT 35.190 208.200 35.510 208.260 ;
        RECT 33.440 207.920 34.960 208.060 ;
        RECT 35.650 207.860 35.970 208.120 ;
        RECT 36.660 208.105 36.800 208.260 ;
        RECT 38.870 208.200 39.190 208.260 ;
        RECT 36.585 207.875 36.875 208.105 ;
        RECT 40.620 208.060 40.760 208.555 ;
        RECT 41.630 208.540 41.950 208.800 ;
        RECT 42.550 208.540 42.870 208.800 ;
        RECT 54.525 208.740 54.815 208.785 ;
        RECT 54.970 208.740 55.290 208.800 ;
        RECT 54.525 208.600 55.290 208.740 ;
        RECT 54.525 208.555 54.815 208.600 ;
        RECT 54.970 208.540 55.290 208.600 ;
        RECT 55.445 208.740 55.735 208.785 ;
        RECT 60.950 208.740 61.270 208.800 ;
        RECT 55.445 208.600 61.270 208.740 ;
        RECT 55.445 208.555 55.735 208.600 ;
        RECT 60.950 208.540 61.270 208.600 ;
        RECT 69.230 208.540 69.550 208.800 ;
        RECT 69.690 208.740 70.010 208.800 ;
        RECT 70.165 208.740 70.455 208.785 ;
        RECT 69.690 208.600 70.455 208.740 ;
        RECT 69.690 208.540 70.010 208.600 ;
        RECT 70.165 208.555 70.455 208.600 ;
        RECT 70.610 208.540 70.930 208.800 ;
        RECT 72.005 208.740 72.295 208.785 ;
        RECT 75.210 208.740 75.530 208.800 ;
        RECT 72.005 208.600 75.530 208.740 ;
        RECT 72.005 208.555 72.295 208.600 ;
        RECT 75.210 208.540 75.530 208.600 ;
        RECT 81.190 208.540 81.510 208.800 ;
        RECT 84.960 208.785 85.100 208.940 ;
        RECT 84.885 208.555 85.175 208.785 ;
        RECT 87.630 208.540 87.950 208.800 ;
        RECT 41.170 208.200 41.490 208.460 ;
        RECT 57.730 208.200 58.050 208.460 ;
        RECT 58.190 208.200 58.510 208.460 ;
        RECT 58.650 208.200 58.970 208.460 ;
        RECT 59.125 208.215 59.415 208.445 ;
        RECT 60.045 208.400 60.335 208.445 ;
        RECT 60.045 208.260 80.500 208.400 ;
        RECT 60.045 208.215 60.335 208.260 ;
        RECT 37.120 207.920 40.760 208.060 ;
        RECT 43.485 208.060 43.775 208.105 ;
        RECT 49.910 208.060 50.230 208.120 ;
        RECT 59.200 208.060 59.340 208.215 ;
        RECT 43.485 207.920 50.230 208.060 ;
        RECT 28.290 207.520 28.610 207.780 ;
        RECT 30.130 207.520 30.450 207.780 ;
        RECT 30.590 207.720 30.910 207.780 ;
        RECT 37.120 207.720 37.260 207.920 ;
        RECT 43.485 207.875 43.775 207.920 ;
        RECT 49.910 207.860 50.230 207.920 ;
        RECT 50.460 207.920 59.340 208.060 ;
        RECT 62.805 208.060 63.095 208.105 ;
        RECT 75.210 208.060 75.530 208.120 ;
        RECT 62.805 207.920 75.530 208.060 ;
        RECT 30.590 207.580 37.260 207.720 ;
        RECT 30.590 207.520 30.910 207.580 ;
        RECT 39.330 207.520 39.650 207.780 ;
        RECT 40.710 207.720 41.030 207.780 ;
        RECT 50.460 207.720 50.600 207.920 ;
        RECT 62.805 207.875 63.095 207.920 ;
        RECT 75.210 207.860 75.530 207.920 ;
        RECT 40.710 207.580 50.600 207.720 ;
        RECT 40.710 207.520 41.030 207.580 ;
        RECT 55.890 207.520 56.210 207.780 ;
        RECT 68.310 207.720 68.630 207.780 ;
        RECT 71.545 207.720 71.835 207.765 ;
        RECT 68.310 207.580 71.835 207.720 ;
        RECT 80.360 207.720 80.500 208.260 ;
        RECT 80.730 208.200 81.050 208.460 ;
        RECT 83.030 208.200 83.350 208.460 ;
        RECT 85.345 208.400 85.635 208.445 ;
        RECT 87.170 208.400 87.490 208.460 ;
        RECT 85.345 208.260 87.490 208.400 ;
        RECT 85.345 208.215 85.635 208.260 ;
        RECT 87.170 208.200 87.490 208.260 ;
        RECT 82.110 208.060 82.430 208.120 ;
        RECT 86.725 208.060 87.015 208.105 ;
        RECT 82.110 207.920 87.015 208.060 ;
        RECT 82.110 207.860 82.430 207.920 ;
        RECT 86.725 207.875 87.015 207.920 ;
        RECT 84.410 207.720 84.730 207.780 ;
        RECT 80.360 207.580 84.730 207.720 ;
        RECT 68.310 207.520 68.630 207.580 ;
        RECT 71.545 207.535 71.835 207.580 ;
        RECT 84.410 207.520 84.730 207.580 ;
        RECT 85.330 207.720 85.650 207.780 ;
        RECT 86.265 207.720 86.555 207.765 ;
        RECT 85.330 207.580 86.555 207.720 ;
        RECT 85.330 207.520 85.650 207.580 ;
        RECT 86.265 207.535 86.555 207.580 ;
        RECT 18.100 206.900 89.400 207.380 ;
        RECT 17.710 206.700 18.030 206.760 ;
        RECT 23.245 206.700 23.535 206.745 ;
        RECT 17.710 206.560 23.535 206.700 ;
        RECT 17.710 206.500 18.030 206.560 ;
        RECT 23.245 206.515 23.535 206.560 ;
        RECT 26.910 206.700 27.230 206.760 ;
        RECT 28.765 206.700 29.055 206.745 ;
        RECT 26.910 206.560 29.055 206.700 ;
        RECT 26.910 206.500 27.230 206.560 ;
        RECT 28.765 206.515 29.055 206.560 ;
        RECT 29.210 206.700 29.530 206.760 ;
        RECT 31.510 206.700 31.830 206.760 ;
        RECT 35.190 206.700 35.510 206.760 ;
        RECT 29.210 206.560 31.830 206.700 ;
        RECT 29.210 206.500 29.530 206.560 ;
        RECT 31.510 206.500 31.830 206.560 ;
        RECT 33.080 206.560 35.510 206.700 ;
        RECT 21.850 206.360 22.170 206.420 ;
        RECT 25.530 206.360 25.850 206.420 ;
        RECT 29.670 206.360 29.990 206.420 ;
        RECT 33.080 206.360 33.220 206.560 ;
        RECT 35.190 206.500 35.510 206.560 ;
        RECT 67.390 206.700 67.710 206.760 ;
        RECT 71.085 206.700 71.375 206.745 ;
        RECT 67.390 206.560 71.375 206.700 ;
        RECT 67.390 206.500 67.710 206.560 ;
        RECT 71.085 206.515 71.375 206.560 ;
        RECT 72.910 206.700 73.230 206.760 ;
        RECT 72.910 206.560 83.260 206.700 ;
        RECT 72.910 206.500 73.230 206.560 ;
        RECT 41.645 206.360 41.935 206.405 ;
        RECT 42.550 206.360 42.870 206.420 ;
        RECT 49.450 206.360 49.770 206.420 ;
        RECT 21.850 206.220 25.300 206.360 ;
        RECT 21.850 206.160 22.170 206.220 ;
        RECT 22.325 206.020 22.615 206.065 ;
        RECT 25.160 206.020 25.300 206.220 ;
        RECT 25.530 206.220 33.220 206.360 ;
        RECT 33.440 206.220 40.760 206.360 ;
        RECT 25.530 206.160 25.850 206.220 ;
        RECT 29.670 206.160 29.990 206.220 ;
        RECT 30.590 206.020 30.910 206.080 ;
        RECT 22.325 205.880 24.840 206.020 ;
        RECT 25.160 205.880 30.910 206.020 ;
        RECT 22.325 205.835 22.615 205.880 ;
        RECT 21.390 205.480 21.710 205.740 ;
        RECT 24.165 205.495 24.455 205.725 ;
        RECT 24.700 205.680 24.840 205.880 ;
        RECT 30.590 205.820 30.910 205.880 ;
        RECT 25.085 205.680 25.375 205.725 ;
        RECT 24.700 205.540 25.375 205.680 ;
        RECT 25.085 205.495 25.375 205.540 ;
        RECT 25.545 205.680 25.835 205.725 ;
        RECT 26.450 205.680 26.770 205.740 ;
        RECT 25.545 205.540 26.770 205.680 ;
        RECT 25.545 205.495 25.835 205.540 ;
        RECT 17.250 205.340 17.570 205.400 ;
        RECT 24.240 205.340 24.380 205.495 ;
        RECT 17.250 205.200 24.380 205.340 ;
        RECT 25.160 205.340 25.300 205.495 ;
        RECT 26.450 205.480 26.770 205.540 ;
        RECT 26.925 205.680 27.215 205.725 ;
        RECT 28.290 205.680 28.610 205.740 ;
        RECT 26.925 205.540 28.610 205.680 ;
        RECT 26.925 205.495 27.215 205.540 ;
        RECT 28.290 205.480 28.610 205.540 ;
        RECT 30.130 205.480 30.450 205.740 ;
        RECT 33.440 205.725 33.580 206.220 ;
        RECT 34.270 206.020 34.590 206.080 ;
        RECT 38.870 206.020 39.190 206.080 ;
        RECT 40.620 206.020 40.760 206.220 ;
        RECT 41.645 206.220 49.770 206.360 ;
        RECT 41.645 206.175 41.935 206.220 ;
        RECT 42.550 206.160 42.870 206.220 ;
        RECT 49.450 206.160 49.770 206.220 ;
        RECT 54.510 206.360 54.830 206.420 ;
        RECT 58.650 206.360 58.970 206.420 ;
        RECT 77.510 206.360 77.830 206.420 ;
        RECT 80.745 206.360 81.035 206.405 ;
        RECT 54.510 206.220 77.830 206.360 ;
        RECT 54.510 206.160 54.830 206.220 ;
        RECT 58.650 206.160 58.970 206.220 ;
        RECT 77.510 206.160 77.830 206.220 ;
        RECT 78.520 206.220 81.035 206.360 ;
        RECT 60.045 206.020 60.335 206.065 ;
        RECT 60.490 206.020 60.810 206.080 ;
        RECT 70.150 206.020 70.470 206.080 ;
        RECT 34.270 205.880 37.720 206.020 ;
        RECT 34.270 205.820 34.590 205.880 ;
        RECT 37.580 205.740 37.720 205.880 ;
        RECT 38.870 205.880 40.475 206.020 ;
        RECT 40.620 205.880 54.280 206.020 ;
        RECT 38.870 205.820 39.190 205.880 ;
        RECT 33.365 205.495 33.655 205.725 ;
        RECT 27.370 205.340 27.690 205.400 ;
        RECT 25.160 205.200 27.690 205.340 ;
        RECT 17.250 205.140 17.570 205.200 ;
        RECT 27.370 205.140 27.690 205.200 ;
        RECT 27.830 205.340 28.150 205.400 ;
        RECT 28.995 205.340 29.285 205.385 ;
        RECT 33.440 205.340 33.580 205.495 ;
        RECT 33.810 205.480 34.130 205.740 ;
        RECT 34.745 205.495 35.035 205.725 ;
        RECT 35.205 205.680 35.495 205.725 ;
        RECT 36.125 205.680 36.415 205.725 ;
        RECT 35.205 205.540 36.415 205.680 ;
        RECT 35.205 205.495 35.495 205.540 ;
        RECT 36.125 205.495 36.415 205.540 ;
        RECT 27.830 205.200 33.580 205.340 ;
        RECT 34.820 205.340 34.960 205.495 ;
        RECT 37.490 205.480 37.810 205.740 ;
        RECT 37.950 205.480 38.270 205.740 ;
        RECT 39.790 205.480 40.110 205.740 ;
        RECT 40.335 205.680 40.475 205.880 ;
        RECT 43.470 205.680 43.790 205.740 ;
        RECT 40.335 205.540 43.790 205.680 ;
        RECT 43.470 205.480 43.790 205.540 ;
        RECT 47.150 205.680 47.470 205.740 ;
        RECT 48.085 205.680 48.375 205.725 ;
        RECT 47.150 205.540 48.375 205.680 ;
        RECT 47.150 205.480 47.470 205.540 ;
        RECT 48.085 205.495 48.375 205.540 ;
        RECT 48.545 205.495 48.835 205.725 ;
        RECT 36.570 205.340 36.890 205.400 ;
        RECT 34.820 205.200 36.890 205.340 ;
        RECT 27.830 205.140 28.150 205.200 ;
        RECT 28.995 205.155 29.285 205.200 ;
        RECT 36.570 205.140 36.890 205.200 ;
        RECT 38.885 205.340 39.175 205.385 ;
        RECT 39.880 205.340 40.020 205.480 ;
        RECT 41.630 205.340 41.950 205.400 ;
        RECT 38.885 205.200 41.950 205.340 ;
        RECT 38.885 205.155 39.175 205.200 ;
        RECT 41.630 205.140 41.950 205.200 ;
        RECT 47.610 205.340 47.930 205.400 ;
        RECT 48.620 205.340 48.760 205.495 ;
        RECT 48.990 205.480 49.310 205.740 ;
        RECT 49.910 205.480 50.230 205.740 ;
        RECT 50.945 205.725 51.085 205.880 ;
        RECT 54.140 205.740 54.280 205.880 ;
        RECT 60.045 205.880 60.810 206.020 ;
        RECT 60.045 205.835 60.335 205.880 ;
        RECT 60.490 205.820 60.810 205.880 ;
        RECT 61.040 205.880 70.470 206.020 ;
        RECT 50.870 205.495 51.160 205.725 ;
        RECT 52.670 205.480 52.990 205.740 ;
        RECT 53.130 205.480 53.450 205.740 ;
        RECT 54.050 205.480 54.370 205.740 ;
        RECT 54.525 205.680 54.815 205.725 ;
        RECT 61.040 205.680 61.180 205.880 ;
        RECT 70.150 205.820 70.470 205.880 ;
        RECT 76.145 206.020 76.435 206.065 ;
        RECT 78.520 206.020 78.660 206.220 ;
        RECT 80.745 206.175 81.035 206.220 ;
        RECT 76.145 205.880 78.660 206.020 ;
        RECT 76.145 205.835 76.435 205.880 ;
        RECT 79.350 205.820 79.670 206.080 ;
        RECT 83.120 206.065 83.260 206.560 ;
        RECT 86.265 206.360 86.555 206.405 ;
        RECT 83.580 206.220 86.555 206.360 ;
        RECT 79.825 206.020 80.115 206.065 ;
        RECT 79.825 205.880 82.800 206.020 ;
        RECT 79.825 205.835 80.115 205.880 ;
        RECT 54.525 205.540 61.180 205.680 ;
        RECT 54.525 205.495 54.815 205.540 ;
        RECT 61.410 205.480 61.730 205.740 ;
        RECT 67.850 205.680 68.170 205.740 ;
        RECT 73.845 205.680 74.135 205.725 ;
        RECT 67.850 205.540 74.135 205.680 ;
        RECT 67.850 205.480 68.170 205.540 ;
        RECT 73.845 205.495 74.135 205.540 ;
        RECT 75.670 205.480 75.990 205.740 ;
        RECT 77.510 205.480 77.830 205.740 ;
        RECT 82.110 205.480 82.430 205.740 ;
        RECT 82.660 205.680 82.800 205.880 ;
        RECT 83.045 205.835 83.335 206.065 ;
        RECT 83.580 205.680 83.720 206.220 ;
        RECT 86.265 206.175 86.555 206.220 ;
        RECT 85.330 205.820 85.650 206.080 ;
        RECT 82.660 205.540 83.720 205.680 ;
        RECT 84.870 205.480 85.190 205.740 ;
        RECT 87.630 205.480 87.950 205.740 ;
        RECT 47.610 205.200 48.760 205.340 ;
        RECT 47.610 205.140 47.930 205.200 ;
        RECT 50.370 205.140 50.690 205.400 ;
        RECT 51.290 205.340 51.610 205.400 ;
        RECT 57.745 205.340 58.035 205.385 ;
        RECT 60.950 205.340 61.270 205.400 ;
        RECT 63.710 205.340 64.030 205.400 ;
        RECT 51.290 205.200 56.120 205.340 ;
        RECT 51.290 205.140 51.610 205.200 ;
        RECT 18.170 205.000 18.490 205.060 ;
        RECT 20.485 205.000 20.775 205.045 ;
        RECT 18.170 204.860 20.775 205.000 ;
        RECT 18.170 204.800 18.490 204.860 ;
        RECT 20.485 204.815 20.775 204.860 ;
        RECT 21.390 205.000 21.710 205.060 ;
        RECT 25.530 205.000 25.850 205.060 ;
        RECT 21.390 204.860 25.850 205.000 ;
        RECT 21.390 204.800 21.710 204.860 ;
        RECT 25.530 204.800 25.850 204.860 ;
        RECT 26.465 205.000 26.755 205.045 ;
        RECT 31.050 205.000 31.370 205.060 ;
        RECT 26.465 204.860 31.370 205.000 ;
        RECT 26.465 204.815 26.755 204.860 ;
        RECT 31.050 204.800 31.370 204.860 ;
        RECT 32.445 205.000 32.735 205.045 ;
        RECT 32.890 205.000 33.210 205.060 ;
        RECT 32.445 204.860 33.210 205.000 ;
        RECT 32.445 204.815 32.735 204.860 ;
        RECT 32.890 204.800 33.210 204.860 ;
        RECT 35.190 205.000 35.510 205.060 ;
        RECT 37.045 205.000 37.335 205.045 ;
        RECT 44.390 205.000 44.710 205.060 ;
        RECT 35.190 204.860 44.710 205.000 ;
        RECT 35.190 204.800 35.510 204.860 ;
        RECT 37.045 204.815 37.335 204.860 ;
        RECT 44.390 204.800 44.710 204.860 ;
        RECT 48.530 205.000 48.850 205.060 ;
        RECT 51.765 205.000 52.055 205.045 ;
        RECT 48.530 204.860 52.055 205.000 ;
        RECT 48.530 204.800 48.850 204.860 ;
        RECT 51.765 204.815 52.055 204.860 ;
        RECT 55.430 204.800 55.750 205.060 ;
        RECT 55.980 205.000 56.120 205.200 ;
        RECT 57.745 205.200 64.030 205.340 ;
        RECT 57.745 205.155 58.035 205.200 ;
        RECT 60.950 205.140 61.270 205.200 ;
        RECT 63.710 205.140 64.030 205.200 ;
        RECT 64.645 205.155 64.935 205.385 ;
        RECT 71.070 205.340 71.390 205.400 ;
        RECT 77.065 205.340 77.355 205.385 ;
        RECT 85.790 205.340 86.110 205.400 ;
        RECT 71.070 205.200 77.355 205.340 ;
        RECT 64.720 205.000 64.860 205.155 ;
        RECT 71.070 205.140 71.390 205.200 ;
        RECT 77.065 205.155 77.355 205.200 ;
        RECT 77.600 205.200 86.110 205.340 ;
        RECT 55.980 204.860 64.860 205.000 ;
        RECT 71.530 205.000 71.850 205.060 ;
        RECT 77.600 205.000 77.740 205.200 ;
        RECT 85.790 205.140 86.110 205.200 ;
        RECT 71.530 204.860 77.740 205.000 ;
        RECT 71.530 204.800 71.850 204.860 ;
        RECT 81.650 204.800 81.970 205.060 ;
        RECT 86.250 205.000 86.570 205.060 ;
        RECT 86.725 205.000 87.015 205.045 ;
        RECT 86.250 204.860 87.015 205.000 ;
        RECT 86.250 204.800 86.570 204.860 ;
        RECT 86.725 204.815 87.015 204.860 ;
        RECT 18.100 204.180 89.400 204.660 ;
        RECT 18.630 203.980 18.950 204.040 ;
        RECT 20.025 203.980 20.315 204.025 ;
        RECT 18.630 203.840 20.315 203.980 ;
        RECT 18.630 203.780 18.950 203.840 ;
        RECT 20.025 203.795 20.315 203.840 ;
        RECT 21.850 203.780 22.170 204.040 ;
        RECT 25.990 203.980 26.310 204.040 ;
        RECT 22.860 203.840 26.310 203.980 ;
        RECT 20.470 203.300 20.790 203.360 ;
        RECT 20.945 203.300 21.235 203.345 ;
        RECT 20.470 203.160 21.235 203.300 ;
        RECT 20.470 203.100 20.790 203.160 ;
        RECT 20.945 203.115 21.235 203.160 ;
        RECT 21.390 203.100 21.710 203.360 ;
        RECT 22.860 203.345 23.000 203.840 ;
        RECT 25.990 203.780 26.310 203.840 ;
        RECT 27.830 203.780 28.150 204.040 ;
        RECT 57.730 203.980 58.050 204.040 ;
        RECT 69.230 203.980 69.550 204.040 ;
        RECT 28.365 203.840 58.050 203.980 ;
        RECT 23.245 203.640 23.535 203.685 ;
        RECT 28.365 203.640 28.505 203.840 ;
        RECT 57.730 203.780 58.050 203.840 ;
        RECT 58.280 203.840 69.550 203.980 ;
        RECT 23.245 203.500 28.505 203.640 ;
        RECT 23.245 203.455 23.535 203.500 ;
        RECT 28.765 203.455 29.055 203.685 ;
        RECT 30.590 203.640 30.910 203.700 ;
        RECT 34.270 203.640 34.590 203.700 ;
        RECT 30.590 203.500 34.590 203.640 ;
        RECT 22.325 203.115 22.615 203.345 ;
        RECT 22.785 203.115 23.075 203.345 ;
        RECT 22.400 202.960 22.540 203.115 ;
        RECT 23.690 203.100 24.010 203.360 ;
        RECT 24.150 203.100 24.470 203.360 ;
        RECT 25.540 203.115 25.830 203.345 ;
        RECT 26.005 203.300 26.295 203.345 ;
        RECT 26.450 203.300 26.770 203.360 ;
        RECT 27.830 203.300 28.150 203.360 ;
        RECT 26.005 203.160 26.770 203.300 ;
        RECT 26.005 203.115 26.295 203.160 ;
        RECT 25.615 202.960 25.755 203.115 ;
        RECT 26.450 203.100 26.770 203.160 ;
        RECT 27.000 203.160 28.150 203.300 ;
        RECT 27.000 202.960 27.140 203.160 ;
        RECT 27.830 203.100 28.150 203.160 ;
        RECT 28.290 203.300 28.610 203.360 ;
        RECT 28.840 203.300 28.980 203.455 ;
        RECT 30.590 203.440 30.910 203.500 ;
        RECT 34.270 203.440 34.590 203.500 ;
        RECT 34.730 203.640 35.050 203.700 ;
        RECT 45.325 203.640 45.615 203.685 ;
        RECT 34.730 203.500 45.615 203.640 ;
        RECT 34.730 203.440 35.050 203.500 ;
        RECT 45.325 203.455 45.615 203.500 ;
        RECT 47.150 203.640 47.470 203.700 ;
        RECT 53.590 203.640 53.910 203.700 ;
        RECT 47.150 203.500 53.910 203.640 ;
        RECT 47.150 203.440 47.470 203.500 ;
        RECT 53.590 203.440 53.910 203.500 ;
        RECT 28.290 203.160 28.980 203.300 ;
        RECT 28.290 203.100 28.610 203.160 ;
        RECT 30.145 203.115 30.435 203.345 ;
        RECT 31.050 203.300 31.370 203.360 ;
        RECT 33.350 203.300 33.670 203.360 ;
        RECT 31.050 203.160 33.670 203.300 ;
        RECT 22.400 202.820 27.140 202.960 ;
        RECT 27.370 202.960 27.690 203.020 ;
        RECT 29.225 202.960 29.515 203.005 ;
        RECT 27.370 202.820 29.515 202.960 ;
        RECT 30.220 202.960 30.360 203.115 ;
        RECT 31.050 203.100 31.370 203.160 ;
        RECT 33.350 203.100 33.670 203.160 ;
        RECT 33.825 203.300 34.115 203.345 ;
        RECT 37.030 203.300 37.350 203.360 ;
        RECT 33.825 203.160 37.350 203.300 ;
        RECT 33.825 203.115 34.115 203.160 ;
        RECT 37.030 203.100 37.350 203.160 ;
        RECT 43.485 203.300 43.775 203.345 ;
        RECT 51.290 203.300 51.610 203.360 ;
        RECT 43.485 203.160 51.610 203.300 ;
        RECT 43.485 203.115 43.775 203.160 ;
        RECT 51.290 203.100 51.610 203.160 ;
        RECT 51.750 203.300 52.070 203.360 ;
        RECT 58.280 203.300 58.420 203.840 ;
        RECT 69.230 203.780 69.550 203.840 ;
        RECT 70.150 203.780 70.470 204.040 ;
        RECT 71.530 203.980 71.850 204.040 ;
        RECT 85.805 203.980 86.095 204.025 ;
        RECT 70.700 203.840 71.850 203.980 ;
        RECT 58.650 203.640 58.970 203.700 ;
        RECT 67.390 203.640 67.710 203.700 ;
        RECT 70.700 203.640 70.840 203.840 ;
        RECT 71.530 203.780 71.850 203.840 ;
        RECT 81.280 203.840 86.095 203.980 ;
        RECT 81.280 203.640 81.420 203.840 ;
        RECT 85.805 203.795 86.095 203.840 ;
        RECT 86.250 203.980 86.570 204.040 ;
        RECT 86.725 203.980 87.015 204.025 ;
        RECT 86.250 203.840 87.015 203.980 ;
        RECT 86.250 203.780 86.570 203.840 ;
        RECT 86.725 203.795 87.015 203.840 ;
        RECT 58.650 203.500 67.710 203.640 ;
        RECT 58.650 203.440 58.970 203.500 ;
        RECT 67.390 203.440 67.710 203.500 ;
        RECT 68.400 203.500 70.840 203.640 ;
        RECT 71.620 203.500 81.420 203.640 ;
        RECT 85.255 203.640 85.545 203.685 ;
        RECT 85.255 203.500 87.860 203.640 ;
        RECT 51.750 203.160 58.420 203.300 ;
        RECT 60.950 203.300 61.270 203.360 ;
        RECT 63.265 203.300 63.555 203.345 ;
        RECT 60.950 203.160 63.555 203.300 ;
        RECT 51.750 203.100 52.070 203.160 ;
        RECT 60.950 203.100 61.270 203.160 ;
        RECT 63.265 203.115 63.555 203.160 ;
        RECT 63.725 203.115 64.015 203.345 ;
        RECT 64.645 203.115 64.935 203.345 ;
        RECT 31.970 202.960 32.290 203.020 ;
        RECT 36.110 202.960 36.430 203.020 ;
        RECT 30.220 202.820 36.430 202.960 ;
        RECT 27.370 202.760 27.690 202.820 ;
        RECT 29.225 202.775 29.515 202.820 ;
        RECT 29.300 202.620 29.440 202.775 ;
        RECT 31.970 202.760 32.290 202.820 ;
        RECT 36.110 202.760 36.430 202.820 ;
        RECT 37.490 202.960 37.810 203.020 ;
        RECT 42.550 202.960 42.870 203.020 ;
        RECT 37.490 202.820 42.870 202.960 ;
        RECT 37.490 202.760 37.810 202.820 ;
        RECT 42.550 202.760 42.870 202.820 ;
        RECT 53.590 202.960 53.910 203.020 ;
        RECT 60.490 202.960 60.810 203.020 ;
        RECT 53.590 202.820 60.810 202.960 ;
        RECT 53.590 202.760 53.910 202.820 ;
        RECT 60.490 202.760 60.810 202.820 ;
        RECT 61.410 202.960 61.730 203.020 ;
        RECT 63.800 202.960 63.940 203.115 ;
        RECT 61.410 202.820 63.940 202.960 ;
        RECT 61.410 202.760 61.730 202.820 ;
        RECT 64.170 202.760 64.490 203.020 ;
        RECT 64.720 202.960 64.860 203.115 ;
        RECT 65.090 203.100 65.410 203.360 ;
        RECT 66.485 203.300 66.775 203.345 ;
        RECT 67.850 203.300 68.170 203.360 ;
        RECT 68.400 203.345 68.540 203.500 ;
        RECT 66.485 203.160 68.170 203.300 ;
        RECT 66.485 203.115 66.775 203.160 ;
        RECT 67.850 203.100 68.170 203.160 ;
        RECT 68.325 203.115 68.615 203.345 ;
        RECT 71.620 203.020 71.760 203.500 ;
        RECT 85.255 203.455 85.545 203.500 ;
        RECT 73.830 203.100 74.150 203.360 ;
        RECT 74.290 203.300 74.610 203.360 ;
        RECT 74.290 203.100 74.750 203.300 ;
        RECT 83.950 203.100 84.270 203.360 ;
        RECT 84.425 203.115 84.715 203.345 ;
        RECT 85.790 203.300 86.110 203.360 ;
        RECT 86.265 203.300 86.555 203.345 ;
        RECT 85.790 203.160 86.555 203.300 ;
        RECT 65.550 202.960 65.870 203.020 ;
        RECT 64.720 202.820 65.870 202.960 ;
        RECT 65.550 202.760 65.870 202.820 ;
        RECT 66.930 202.760 67.250 203.020 ;
        RECT 69.230 202.960 69.550 203.020 ;
        RECT 70.610 202.960 70.930 203.020 ;
        RECT 69.230 202.820 70.930 202.960 ;
        RECT 69.230 202.760 69.550 202.820 ;
        RECT 70.610 202.760 70.930 202.820 ;
        RECT 71.070 202.760 71.390 203.020 ;
        RECT 71.530 202.760 71.850 203.020 ;
        RECT 73.385 202.960 73.675 203.005 ;
        RECT 74.610 202.960 74.750 203.100 ;
        RECT 80.730 202.960 81.050 203.020 ;
        RECT 84.500 202.960 84.640 203.115 ;
        RECT 85.790 203.100 86.110 203.160 ;
        RECT 86.265 203.115 86.555 203.160 ;
        RECT 73.385 202.820 80.500 202.960 ;
        RECT 73.385 202.775 73.675 202.820 ;
        RECT 30.130 202.620 30.450 202.680 ;
        RECT 29.300 202.480 30.450 202.620 ;
        RECT 30.130 202.420 30.450 202.480 ;
        RECT 33.350 202.620 33.670 202.680 ;
        RECT 38.870 202.620 39.190 202.680 ;
        RECT 33.350 202.480 39.190 202.620 ;
        RECT 33.350 202.420 33.670 202.480 ;
        RECT 38.870 202.420 39.190 202.480 ;
        RECT 39.330 202.620 39.650 202.680 ;
        RECT 61.870 202.620 62.190 202.680 ;
        RECT 74.305 202.620 74.595 202.665 ;
        RECT 39.330 202.480 60.950 202.620 ;
        RECT 39.330 202.420 39.650 202.480 ;
        RECT 25.990 202.280 26.310 202.340 ;
        RECT 26.925 202.280 27.215 202.325 ;
        RECT 25.990 202.140 27.215 202.280 ;
        RECT 25.990 202.080 26.310 202.140 ;
        RECT 26.925 202.095 27.215 202.140 ;
        RECT 27.845 202.280 28.135 202.325 ;
        RECT 28.290 202.280 28.610 202.340 ;
        RECT 27.845 202.140 28.610 202.280 ;
        RECT 27.845 202.095 28.135 202.140 ;
        RECT 28.290 202.080 28.610 202.140 ;
        RECT 29.670 202.280 29.990 202.340 ;
        RECT 30.590 202.280 30.910 202.340 ;
        RECT 29.670 202.140 30.910 202.280 ;
        RECT 29.670 202.080 29.990 202.140 ;
        RECT 30.590 202.080 30.910 202.140 ;
        RECT 31.050 202.080 31.370 202.340 ;
        RECT 37.030 202.280 37.350 202.340 ;
        RECT 41.170 202.280 41.490 202.340 ;
        RECT 50.370 202.280 50.690 202.340 ;
        RECT 37.030 202.140 50.690 202.280 ;
        RECT 37.030 202.080 37.350 202.140 ;
        RECT 41.170 202.080 41.490 202.140 ;
        RECT 50.370 202.080 50.690 202.140 ;
        RECT 56.810 202.080 57.130 202.340 ;
        RECT 60.810 202.280 60.950 202.480 ;
        RECT 61.870 202.480 74.595 202.620 ;
        RECT 80.360 202.620 80.500 202.820 ;
        RECT 80.730 202.820 84.640 202.960 ;
        RECT 80.730 202.760 81.050 202.820 ;
        RECT 87.720 202.620 87.860 203.500 ;
        RECT 80.360 202.480 87.860 202.620 ;
        RECT 61.870 202.420 62.190 202.480 ;
        RECT 74.305 202.435 74.595 202.480 ;
        RECT 66.470 202.280 66.790 202.340 ;
        RECT 73.830 202.280 74.150 202.340 ;
        RECT 60.810 202.140 74.150 202.280 ;
        RECT 66.470 202.080 66.790 202.140 ;
        RECT 73.830 202.080 74.150 202.140 ;
        RECT 76.590 202.080 76.910 202.340 ;
        RECT 18.100 201.460 89.400 201.940 ;
        RECT 24.610 201.260 24.930 201.320 ;
        RECT 25.545 201.260 25.835 201.305 ;
        RECT 37.490 201.260 37.810 201.320 ;
        RECT 24.610 201.120 25.835 201.260 ;
        RECT 24.610 201.060 24.930 201.120 ;
        RECT 25.545 201.075 25.835 201.120 ;
        RECT 30.680 201.120 37.810 201.260 ;
        RECT 17.710 200.920 18.030 200.980 ;
        RECT 22.785 200.920 23.075 200.965 ;
        RECT 17.710 200.780 23.075 200.920 ;
        RECT 17.710 200.720 18.030 200.780 ;
        RECT 22.785 200.735 23.075 200.780 ;
        RECT 26.465 200.580 26.755 200.625 ;
        RECT 29.670 200.580 29.990 200.640 ;
        RECT 30.680 200.580 30.820 201.120 ;
        RECT 37.490 201.060 37.810 201.120 ;
        RECT 37.950 201.260 38.270 201.320 ;
        RECT 39.790 201.260 40.110 201.320 ;
        RECT 37.950 201.120 40.110 201.260 ;
        RECT 37.950 201.060 38.270 201.120 ;
        RECT 39.790 201.060 40.110 201.120 ;
        RECT 40.725 201.260 41.015 201.305 ;
        RECT 76.130 201.260 76.450 201.320 ;
        RECT 40.725 201.120 76.450 201.260 ;
        RECT 40.725 201.075 41.015 201.120 ;
        RECT 76.130 201.060 76.450 201.120 ;
        RECT 31.510 200.720 31.830 200.980 ;
        RECT 33.350 200.920 33.670 200.980 ;
        RECT 46.690 200.920 47.010 200.980 ;
        RECT 33.350 200.780 47.010 200.920 ;
        RECT 33.350 200.720 33.670 200.780 ;
        RECT 46.690 200.720 47.010 200.780 ;
        RECT 49.925 200.920 50.215 200.965 ;
        RECT 51.290 200.920 51.610 200.980 ;
        RECT 49.925 200.780 51.610 200.920 ;
        RECT 49.925 200.735 50.215 200.780 ;
        RECT 51.290 200.720 51.610 200.780 ;
        RECT 58.650 200.720 58.970 200.980 ;
        RECT 59.110 200.920 59.430 200.980 ;
        RECT 78.445 200.920 78.735 200.965 ;
        RECT 59.110 200.780 78.735 200.920 ;
        RECT 59.110 200.720 59.430 200.780 ;
        RECT 78.445 200.735 78.735 200.780 ;
        RECT 79.810 200.920 80.130 200.980 ;
        RECT 87.185 200.920 87.475 200.965 ;
        RECT 79.810 200.780 87.475 200.920 ;
        RECT 79.810 200.720 80.130 200.780 ;
        RECT 87.185 200.735 87.475 200.780 ;
        RECT 21.940 200.440 26.755 200.580 ;
        RECT 21.940 200.300 22.080 200.440 ;
        RECT 26.465 200.395 26.755 200.440 ;
        RECT 27.460 200.440 29.990 200.580 ;
        RECT 20.485 200.240 20.775 200.285 ;
        RECT 21.850 200.240 22.170 200.300 ;
        RECT 20.485 200.100 22.170 200.240 ;
        RECT 20.485 200.055 20.775 200.100 ;
        RECT 21.850 200.040 22.170 200.100 ;
        RECT 23.690 200.040 24.010 200.300 ;
        RECT 25.070 200.040 25.390 200.300 ;
        RECT 25.530 200.240 25.850 200.300 ;
        RECT 27.460 200.285 27.600 200.440 ;
        RECT 29.670 200.380 29.990 200.440 ;
        RECT 30.220 200.440 30.820 200.580 ;
        RECT 31.970 200.580 32.290 200.640 ;
        RECT 45.310 200.580 45.630 200.640 ;
        RECT 58.740 200.580 58.880 200.720 ;
        RECT 31.970 200.440 45.630 200.580 ;
        RECT 30.220 200.285 30.360 200.440 ;
        RECT 31.970 200.380 32.290 200.440 ;
        RECT 45.310 200.380 45.630 200.440 ;
        RECT 57.820 200.440 58.880 200.580 ;
        RECT 60.505 200.580 60.795 200.625 ;
        RECT 72.910 200.580 73.230 200.640 ;
        RECT 60.505 200.440 73.230 200.580 ;
        RECT 26.005 200.240 26.295 200.285 ;
        RECT 25.530 200.100 26.295 200.240 ;
        RECT 25.530 200.040 25.850 200.100 ;
        RECT 26.005 200.055 26.295 200.100 ;
        RECT 27.385 200.055 27.675 200.285 ;
        RECT 28.765 200.240 29.055 200.285 ;
        RECT 27.920 200.100 29.055 200.240 ;
        RECT 26.450 199.900 26.770 199.960 ;
        RECT 27.920 199.900 28.060 200.100 ;
        RECT 28.765 200.055 29.055 200.100 ;
        RECT 30.145 200.055 30.435 200.285 ;
        RECT 30.605 200.240 30.895 200.285 ;
        RECT 30.605 200.100 32.200 200.240 ;
        RECT 30.605 200.055 30.895 200.100 ;
        RECT 26.450 199.760 28.060 199.900 ;
        RECT 28.305 199.900 28.595 199.945 ;
        RECT 31.510 199.900 31.830 199.960 ;
        RECT 28.305 199.760 31.830 199.900 ;
        RECT 32.060 199.900 32.200 200.100 ;
        RECT 32.430 200.040 32.750 200.300 ;
        RECT 32.905 200.240 33.195 200.285 ;
        RECT 33.810 200.240 34.130 200.300 ;
        RECT 32.905 200.100 34.130 200.240 ;
        RECT 32.905 200.055 33.195 200.100 ;
        RECT 33.810 200.040 34.130 200.100 ;
        RECT 34.270 200.040 34.590 200.300 ;
        RECT 54.510 200.240 54.830 200.300 ;
        RECT 34.820 200.100 54.830 200.240 ;
        RECT 34.820 199.900 34.960 200.100 ;
        RECT 54.510 200.040 54.830 200.100 ;
        RECT 55.430 200.240 55.750 200.300 ;
        RECT 57.285 200.240 57.575 200.285 ;
        RECT 57.820 200.240 57.960 200.440 ;
        RECT 60.505 200.395 60.795 200.440 ;
        RECT 72.910 200.380 73.230 200.440 ;
        RECT 55.430 200.100 57.960 200.240 ;
        RECT 55.430 200.040 55.750 200.100 ;
        RECT 57.285 200.055 57.575 200.100 ;
        RECT 58.190 200.040 58.510 200.300 ;
        RECT 58.650 200.040 58.970 200.300 ;
        RECT 59.585 200.055 59.875 200.285 ;
        RECT 60.030 200.240 60.350 200.300 ;
        RECT 61.425 200.240 61.715 200.285 ;
        RECT 60.030 200.100 61.715 200.240 ;
        RECT 32.060 199.760 34.960 199.900 ;
        RECT 36.125 199.900 36.415 199.945 ;
        RECT 38.410 199.900 38.730 199.960 ;
        RECT 36.125 199.760 38.730 199.900 ;
        RECT 26.450 199.700 26.770 199.760 ;
        RECT 28.305 199.715 28.595 199.760 ;
        RECT 31.510 199.700 31.830 199.760 ;
        RECT 36.125 199.715 36.415 199.760 ;
        RECT 38.410 199.700 38.730 199.760 ;
        RECT 38.870 199.900 39.190 199.960 ;
        RECT 46.690 199.900 47.010 199.960 ;
        RECT 38.870 199.760 47.010 199.900 ;
        RECT 38.870 199.700 39.190 199.760 ;
        RECT 46.690 199.700 47.010 199.760 ;
        RECT 47.150 199.700 47.470 199.960 ;
        RECT 53.590 199.900 53.910 199.960 ;
        RECT 56.365 199.900 56.655 199.945 ;
        RECT 53.590 199.760 56.655 199.900 ;
        RECT 53.590 199.700 53.910 199.760 ;
        RECT 56.365 199.715 56.655 199.760 ;
        RECT 21.405 199.560 21.695 199.605 ;
        RECT 22.310 199.560 22.630 199.620 ;
        RECT 21.405 199.420 22.630 199.560 ;
        RECT 21.405 199.375 21.695 199.420 ;
        RECT 22.310 199.360 22.630 199.420 ;
        RECT 25.530 199.560 25.850 199.620 ;
        RECT 26.910 199.560 27.230 199.620 ;
        RECT 25.530 199.420 27.230 199.560 ;
        RECT 25.530 199.360 25.850 199.420 ;
        RECT 26.910 199.360 27.230 199.420 ;
        RECT 27.370 199.560 27.690 199.620 ;
        RECT 28.765 199.560 29.055 199.605 ;
        RECT 27.370 199.420 29.055 199.560 ;
        RECT 27.370 199.360 27.690 199.420 ;
        RECT 28.765 199.375 29.055 199.420 ;
        RECT 29.685 199.560 29.975 199.605 ;
        RECT 32.430 199.560 32.750 199.620 ;
        RECT 29.685 199.420 32.750 199.560 ;
        RECT 29.685 199.375 29.975 199.420 ;
        RECT 32.430 199.360 32.750 199.420 ;
        RECT 33.365 199.560 33.655 199.605 ;
        RECT 33.810 199.560 34.130 199.620 ;
        RECT 33.365 199.420 34.130 199.560 ;
        RECT 33.365 199.375 33.655 199.420 ;
        RECT 33.810 199.360 34.130 199.420 ;
        RECT 35.205 199.560 35.495 199.605 ;
        RECT 41.630 199.560 41.950 199.620 ;
        RECT 35.205 199.420 41.950 199.560 ;
        RECT 35.205 199.375 35.495 199.420 ;
        RECT 41.630 199.360 41.950 199.420 ;
        RECT 45.770 199.560 46.090 199.620 ;
        RECT 59.660 199.560 59.800 200.055 ;
        RECT 60.030 200.040 60.350 200.100 ;
        RECT 61.425 200.055 61.715 200.100 ;
        RECT 62.345 200.240 62.635 200.285 ;
        RECT 63.250 200.240 63.570 200.300 ;
        RECT 81.205 200.240 81.495 200.285 ;
        RECT 81.650 200.240 81.970 200.300 ;
        RECT 62.345 200.100 72.680 200.240 ;
        RECT 62.345 200.055 62.635 200.100 ;
        RECT 63.250 200.040 63.570 200.100 ;
        RECT 60.490 199.900 60.810 199.960 ;
        RECT 62.805 199.900 63.095 199.945 ;
        RECT 72.005 199.900 72.295 199.945 ;
        RECT 60.490 199.760 63.095 199.900 ;
        RECT 60.490 199.700 60.810 199.760 ;
        RECT 62.805 199.715 63.095 199.760 ;
        RECT 63.340 199.760 72.295 199.900 ;
        RECT 72.540 199.900 72.680 200.100 ;
        RECT 81.205 200.100 81.970 200.240 ;
        RECT 81.205 200.055 81.495 200.100 ;
        RECT 81.280 199.900 81.420 200.055 ;
        RECT 81.650 200.040 81.970 200.100 ;
        RECT 82.570 200.240 82.890 200.300 ;
        RECT 83.045 200.240 83.335 200.285 ;
        RECT 82.570 200.100 83.335 200.240 ;
        RECT 82.570 200.040 82.890 200.100 ;
        RECT 83.045 200.055 83.335 200.100 ;
        RECT 83.490 200.240 83.810 200.300 ;
        RECT 85.345 200.240 85.635 200.285 ;
        RECT 86.265 200.240 86.555 200.285 ;
        RECT 83.490 200.100 85.635 200.240 ;
        RECT 83.490 200.040 83.810 200.100 ;
        RECT 85.345 200.055 85.635 200.100 ;
        RECT 85.880 200.100 86.555 200.240 ;
        RECT 72.540 199.760 81.420 199.900 ;
        RECT 45.770 199.420 59.800 199.560 ;
        RECT 61.410 199.560 61.730 199.620 ;
        RECT 61.885 199.560 62.175 199.605 ;
        RECT 61.410 199.420 62.175 199.560 ;
        RECT 45.770 199.360 46.090 199.420 ;
        RECT 61.410 199.360 61.730 199.420 ;
        RECT 61.885 199.375 62.175 199.420 ;
        RECT 62.330 199.560 62.650 199.620 ;
        RECT 63.340 199.560 63.480 199.760 ;
        RECT 72.005 199.715 72.295 199.760 ;
        RECT 84.410 199.700 84.730 199.960 ;
        RECT 62.330 199.420 63.480 199.560 ;
        RECT 63.710 199.560 64.030 199.620 ;
        RECT 69.245 199.560 69.535 199.605 ;
        RECT 63.710 199.420 69.535 199.560 ;
        RECT 62.330 199.360 62.650 199.420 ;
        RECT 63.710 199.360 64.030 199.420 ;
        RECT 69.245 199.375 69.535 199.420 ;
        RECT 82.125 199.560 82.415 199.605 ;
        RECT 85.880 199.560 86.020 200.100 ;
        RECT 86.265 200.055 86.555 200.100 ;
        RECT 82.125 199.420 86.020 199.560 ;
        RECT 82.125 199.375 82.415 199.420 ;
        RECT 18.100 198.740 89.400 199.220 ;
        RECT 22.325 198.540 22.615 198.585 ;
        RECT 22.770 198.540 23.090 198.600 ;
        RECT 22.325 198.400 23.090 198.540 ;
        RECT 22.325 198.355 22.615 198.400 ;
        RECT 22.770 198.340 23.090 198.400 ;
        RECT 23.230 198.540 23.550 198.600 ;
        RECT 23.705 198.540 23.995 198.585 ;
        RECT 23.230 198.400 23.995 198.540 ;
        RECT 23.230 198.340 23.550 198.400 ;
        RECT 23.705 198.355 23.995 198.400 ;
        RECT 30.605 198.540 30.895 198.585 ;
        RECT 31.970 198.540 32.290 198.600 ;
        RECT 30.605 198.400 32.290 198.540 ;
        RECT 30.605 198.355 30.895 198.400 ;
        RECT 31.970 198.340 32.290 198.400 ;
        RECT 35.650 198.540 35.970 198.600 ;
        RECT 35.650 198.400 37.720 198.540 ;
        RECT 35.650 198.340 35.970 198.400 ;
        RECT 20.930 197.660 21.250 197.920 ;
        RECT 22.860 197.905 23.000 198.340 ;
        RECT 24.610 198.200 24.930 198.260 ;
        RECT 26.005 198.200 26.295 198.245 ;
        RECT 24.610 198.060 26.295 198.200 ;
        RECT 24.610 198.000 24.930 198.060 ;
        RECT 26.005 198.015 26.295 198.060 ;
        RECT 27.370 198.200 27.690 198.260 ;
        RECT 27.370 198.060 28.520 198.200 ;
        RECT 27.370 198.000 27.690 198.060 ;
        RECT 22.785 197.675 23.075 197.905 ;
        RECT 25.070 197.660 25.390 197.920 ;
        RECT 25.530 197.660 25.850 197.920 ;
        RECT 26.450 197.905 26.770 197.920 ;
        RECT 26.450 197.860 26.985 197.905 ;
        RECT 27.845 197.860 28.135 197.905 ;
        RECT 26.450 197.720 28.135 197.860 ;
        RECT 28.380 197.860 28.520 198.060 ;
        RECT 31.510 198.000 31.830 198.260 ;
        RECT 37.580 198.245 37.720 198.400 ;
        RECT 39.330 198.340 39.650 198.600 ;
        RECT 40.710 198.340 41.030 198.600 ;
        RECT 41.170 198.540 41.490 198.600 ;
        RECT 48.085 198.540 48.375 198.585 ;
        RECT 48.990 198.540 49.310 198.600 ;
        RECT 55.430 198.540 55.750 198.600 ;
        RECT 41.170 198.400 47.840 198.540 ;
        RECT 41.170 198.340 41.490 198.400 ;
        RECT 32.100 198.060 37.260 198.200 ;
        RECT 28.765 197.860 29.055 197.905 ;
        RECT 28.380 197.720 29.055 197.860 ;
        RECT 26.450 197.675 26.985 197.720 ;
        RECT 27.845 197.675 28.135 197.720 ;
        RECT 28.765 197.675 29.055 197.720 ;
        RECT 30.145 197.860 30.435 197.905 ;
        RECT 32.100 197.860 32.240 198.060 ;
        RECT 32.980 197.905 33.120 198.060 ;
        RECT 37.120 197.920 37.260 198.060 ;
        RECT 37.505 198.015 37.795 198.245 ;
        RECT 38.410 198.200 38.730 198.260 ;
        RECT 47.700 198.200 47.840 198.400 ;
        RECT 48.085 198.400 49.310 198.540 ;
        RECT 48.085 198.355 48.375 198.400 ;
        RECT 48.990 198.340 49.310 198.400 ;
        RECT 49.540 198.400 55.750 198.540 ;
        RECT 49.540 198.200 49.680 198.400 ;
        RECT 55.430 198.340 55.750 198.400 ;
        RECT 56.810 198.540 57.130 198.600 ;
        RECT 68.325 198.540 68.615 198.585 ;
        RECT 69.230 198.540 69.550 198.600 ;
        RECT 56.810 198.400 67.160 198.540 ;
        RECT 56.810 198.340 57.130 198.400 ;
        RECT 52.225 198.200 52.515 198.245 ;
        RECT 53.130 198.200 53.450 198.260 ;
        RECT 38.410 198.060 47.380 198.200 ;
        RECT 47.700 198.060 49.680 198.200 ;
        RECT 38.410 198.000 38.730 198.060 ;
        RECT 30.145 197.720 32.240 197.860 ;
        RECT 30.145 197.675 30.435 197.720 ;
        RECT 32.445 197.675 32.735 197.905 ;
        RECT 32.905 197.675 33.195 197.905 ;
        RECT 33.350 197.860 33.670 197.920 ;
        RECT 33.825 197.860 34.115 197.905 ;
        RECT 33.350 197.720 34.115 197.860 ;
        RECT 26.450 197.660 26.770 197.675 ;
        RECT 24.150 197.320 24.470 197.580 ;
        RECT 27.370 197.320 27.690 197.580 ;
        RECT 28.290 197.520 28.610 197.580 ;
        RECT 29.685 197.520 29.975 197.565 ;
        RECT 28.290 197.380 29.975 197.520 ;
        RECT 28.290 197.320 28.610 197.380 ;
        RECT 29.685 197.335 29.975 197.380 ;
        RECT 31.510 197.520 31.830 197.580 ;
        RECT 32.520 197.520 32.660 197.675 ;
        RECT 33.350 197.660 33.670 197.720 ;
        RECT 33.825 197.675 34.115 197.720 ;
        RECT 34.270 197.660 34.590 197.920 ;
        RECT 34.745 197.860 35.035 197.905 ;
        RECT 34.745 197.720 36.870 197.860 ;
        RECT 34.745 197.675 35.035 197.720 ;
        RECT 31.510 197.380 32.660 197.520 ;
        RECT 29.760 197.180 29.900 197.335 ;
        RECT 31.510 197.320 31.830 197.380 ;
        RECT 34.820 197.180 34.960 197.675 ;
        RECT 36.730 197.520 36.870 197.720 ;
        RECT 37.030 197.660 37.350 197.920 ;
        RECT 37.965 197.675 38.255 197.905 ;
        RECT 38.040 197.520 38.180 197.675 ;
        RECT 38.870 197.660 39.190 197.920 ;
        RECT 39.420 197.905 39.560 198.060 ;
        RECT 39.345 197.675 39.635 197.905 ;
        RECT 40.265 197.860 40.555 197.905 ;
        RECT 41.170 197.860 41.490 197.920 ;
        RECT 40.265 197.720 41.490 197.860 ;
        RECT 40.265 197.675 40.555 197.720 ;
        RECT 41.170 197.660 41.490 197.720 ;
        RECT 41.630 197.660 41.950 197.920 ;
        RECT 42.105 197.860 42.395 197.905 ;
        RECT 43.930 197.860 44.250 197.920 ;
        RECT 42.105 197.720 44.250 197.860 ;
        RECT 42.105 197.675 42.395 197.720 ;
        RECT 43.930 197.660 44.250 197.720 ;
        RECT 44.390 197.860 44.710 197.920 ;
        RECT 44.865 197.860 45.155 197.905 ;
        RECT 44.390 197.720 45.155 197.860 ;
        RECT 44.390 197.660 44.710 197.720 ;
        RECT 44.865 197.675 45.155 197.720 ;
        RECT 45.310 197.660 45.630 197.920 ;
        RECT 47.240 197.905 47.380 198.060 ;
        RECT 47.165 197.675 47.455 197.905 ;
        RECT 49.005 197.860 49.295 197.905 ;
        RECT 49.540 197.860 49.680 198.060 ;
        RECT 50.460 198.060 51.505 198.200 ;
        RECT 49.005 197.720 49.680 197.860 ;
        RECT 49.005 197.675 49.295 197.720 ;
        RECT 49.910 197.660 50.230 197.920 ;
        RECT 50.460 197.905 50.600 198.060 ;
        RECT 50.385 197.675 50.675 197.905 ;
        RECT 50.850 197.625 51.140 197.855 ;
        RECT 40.710 197.520 41.030 197.580 ;
        RECT 36.730 197.380 41.030 197.520 ;
        RECT 40.710 197.320 41.030 197.380 ;
        RECT 42.550 197.320 42.870 197.580 ;
        RECT 43.010 197.320 43.330 197.580 ;
        RECT 29.760 197.040 34.960 197.180 ;
        RECT 35.665 197.180 35.955 197.225 ;
        RECT 39.790 197.180 40.110 197.240 ;
        RECT 50.925 197.180 51.065 197.625 ;
        RECT 35.665 197.040 37.260 197.180 ;
        RECT 35.665 196.995 35.955 197.040 ;
        RECT 20.010 196.640 20.330 196.900 ;
        RECT 31.970 196.840 32.290 196.900 ;
        RECT 36.125 196.840 36.415 196.885 ;
        RECT 31.970 196.700 36.415 196.840 ;
        RECT 37.120 196.840 37.260 197.040 ;
        RECT 39.790 197.040 51.065 197.180 ;
        RECT 39.790 196.980 40.110 197.040 ;
        RECT 38.410 196.840 38.730 196.900 ;
        RECT 37.120 196.700 38.730 196.840 ;
        RECT 31.970 196.640 32.290 196.700 ;
        RECT 36.125 196.655 36.415 196.700 ;
        RECT 38.410 196.640 38.730 196.700 ;
        RECT 42.550 196.840 42.870 196.900 ;
        RECT 47.165 196.840 47.455 196.885 ;
        RECT 51.365 196.840 51.505 198.060 ;
        RECT 52.225 198.060 53.450 198.200 ;
        RECT 52.225 198.015 52.515 198.060 ;
        RECT 53.130 198.000 53.450 198.060 ;
        RECT 58.190 198.200 58.510 198.260 ;
        RECT 66.485 198.200 66.775 198.245 ;
        RECT 58.190 198.060 66.775 198.200 ;
        RECT 67.020 198.200 67.160 198.400 ;
        RECT 68.325 198.400 69.550 198.540 ;
        RECT 68.325 198.355 68.615 198.400 ;
        RECT 69.230 198.340 69.550 198.400 ;
        RECT 70.150 198.540 70.470 198.600 ;
        RECT 76.605 198.540 76.895 198.585 ;
        RECT 70.150 198.400 76.895 198.540 ;
        RECT 70.150 198.340 70.470 198.400 ;
        RECT 76.605 198.355 76.895 198.400 ;
        RECT 80.730 198.540 81.050 198.600 ;
        RECT 84.410 198.540 84.730 198.600 ;
        RECT 80.730 198.400 84.730 198.540 ;
        RECT 80.730 198.340 81.050 198.400 ;
        RECT 84.410 198.340 84.730 198.400 ;
        RECT 86.725 198.540 87.015 198.585 ;
        RECT 89.470 198.540 89.790 198.600 ;
        RECT 86.725 198.400 89.790 198.540 ;
        RECT 86.725 198.355 87.015 198.400 ;
        RECT 89.470 198.340 89.790 198.400 ;
        RECT 71.990 198.200 72.310 198.260 ;
        RECT 67.020 198.060 70.380 198.200 ;
        RECT 58.190 198.000 58.510 198.060 ;
        RECT 66.485 198.015 66.775 198.060 ;
        RECT 52.685 197.860 52.975 197.905 ;
        RECT 55.890 197.860 56.210 197.920 ;
        RECT 52.685 197.720 56.210 197.860 ;
        RECT 52.685 197.675 52.975 197.720 ;
        RECT 55.890 197.660 56.210 197.720 ;
        RECT 61.870 197.660 62.190 197.920 ;
        RECT 62.790 197.660 63.110 197.920 ;
        RECT 63.710 197.660 64.030 197.920 ;
        RECT 65.105 197.860 65.395 197.905 ;
        RECT 67.405 197.860 67.695 197.905 ;
        RECT 65.105 197.720 67.695 197.860 ;
        RECT 65.105 197.675 65.395 197.720 ;
        RECT 67.405 197.675 67.695 197.720 ;
        RECT 68.785 197.860 69.075 197.905 ;
        RECT 69.690 197.860 70.010 197.920 ;
        RECT 70.240 197.905 70.380 198.060 ;
        RECT 71.990 198.060 81.880 198.200 ;
        RECT 71.990 198.000 72.310 198.060 ;
        RECT 68.785 197.720 70.010 197.860 ;
        RECT 68.785 197.675 69.075 197.720 ;
        RECT 60.490 197.520 60.810 197.580 ;
        RECT 62.330 197.520 62.650 197.580 ;
        RECT 60.490 197.380 62.650 197.520 ;
        RECT 60.490 197.320 60.810 197.380 ;
        RECT 62.330 197.320 62.650 197.380 ;
        RECT 63.265 197.335 63.555 197.565 ;
        RECT 64.185 197.335 64.475 197.565 ;
        RECT 56.810 197.180 57.130 197.240 ;
        RECT 62.790 197.180 63.110 197.240 ;
        RECT 63.340 197.180 63.480 197.335 ;
        RECT 56.810 197.040 59.340 197.180 ;
        RECT 56.810 196.980 57.130 197.040 ;
        RECT 42.550 196.700 51.505 196.840 ;
        RECT 54.510 196.840 54.830 196.900 ;
        RECT 58.650 196.840 58.970 196.900 ;
        RECT 54.510 196.700 58.970 196.840 ;
        RECT 59.200 196.840 59.340 197.040 ;
        RECT 62.790 197.040 63.480 197.180 ;
        RECT 63.710 197.180 64.030 197.240 ;
        RECT 64.260 197.180 64.400 197.335 ;
        RECT 63.710 197.040 64.400 197.180 ;
        RECT 62.790 196.980 63.110 197.040 ;
        RECT 63.710 196.980 64.030 197.040 ;
        RECT 68.860 196.840 69.000 197.675 ;
        RECT 69.690 197.660 70.010 197.720 ;
        RECT 70.165 197.675 70.455 197.905 ;
        RECT 70.610 197.860 70.930 197.920 ;
        RECT 79.365 197.860 79.655 197.905 ;
        RECT 70.610 197.720 79.655 197.860 ;
        RECT 70.610 197.660 70.930 197.720 ;
        RECT 79.365 197.675 79.655 197.720 ;
        RECT 80.730 197.660 81.050 197.920 ;
        RECT 81.190 197.660 81.510 197.920 ;
        RECT 81.740 197.905 81.880 198.060 ;
        RECT 82.200 198.060 86.020 198.200 ;
        RECT 82.200 197.905 82.340 198.060 ;
        RECT 85.880 197.920 86.020 198.060 ;
        RECT 81.665 197.675 81.955 197.905 ;
        RECT 82.125 197.675 82.415 197.905 ;
        RECT 84.410 197.660 84.730 197.920 ;
        RECT 85.790 197.660 86.110 197.920 ;
        RECT 87.645 197.860 87.935 197.905 ;
        RECT 88.090 197.860 88.410 197.920 ;
        RECT 87.645 197.720 88.410 197.860 ;
        RECT 87.645 197.675 87.935 197.720 ;
        RECT 88.090 197.660 88.410 197.720 ;
        RECT 78.890 197.520 79.210 197.580 ;
        RECT 83.505 197.520 83.795 197.565 ;
        RECT 85.345 197.520 85.635 197.565 ;
        RECT 78.890 197.380 83.795 197.520 ;
        RECT 78.890 197.320 79.210 197.380 ;
        RECT 83.505 197.335 83.795 197.380 ;
        RECT 84.040 197.380 85.635 197.520 ;
        RECT 81.190 197.180 81.510 197.240 ;
        RECT 84.040 197.180 84.180 197.380 ;
        RECT 85.345 197.335 85.635 197.380 ;
        RECT 81.190 197.040 84.180 197.180 ;
        RECT 81.190 196.980 81.510 197.040 ;
        RECT 84.905 196.995 85.195 197.225 ;
        RECT 59.200 196.700 69.000 196.840 ;
        RECT 80.270 196.840 80.590 196.900 ;
        RECT 84.960 196.840 85.100 196.995 ;
        RECT 80.270 196.700 85.100 196.840 ;
        RECT 42.550 196.640 42.870 196.700 ;
        RECT 47.165 196.655 47.455 196.700 ;
        RECT 54.510 196.640 54.830 196.700 ;
        RECT 58.650 196.640 58.970 196.700 ;
        RECT 80.270 196.640 80.590 196.700 ;
        RECT 18.100 196.020 89.400 196.500 ;
        RECT 24.625 195.820 24.915 195.865 ;
        RECT 25.070 195.820 25.390 195.880 ;
        RECT 24.625 195.680 25.390 195.820 ;
        RECT 24.625 195.635 24.915 195.680 ;
        RECT 25.070 195.620 25.390 195.680 ;
        RECT 29.210 195.820 29.530 195.880 ;
        RECT 29.685 195.820 29.975 195.865 ;
        RECT 29.210 195.680 29.975 195.820 ;
        RECT 29.210 195.620 29.530 195.680 ;
        RECT 29.685 195.635 29.975 195.680 ;
        RECT 30.590 195.820 30.910 195.880 ;
        RECT 31.985 195.820 32.275 195.865 ;
        RECT 30.590 195.680 32.275 195.820 ;
        RECT 30.590 195.620 30.910 195.680 ;
        RECT 31.985 195.635 32.275 195.680 ;
        RECT 33.825 195.820 34.115 195.865 ;
        RECT 44.390 195.820 44.710 195.880 ;
        RECT 33.825 195.680 44.710 195.820 ;
        RECT 33.825 195.635 34.115 195.680 ;
        RECT 44.390 195.620 44.710 195.680 ;
        RECT 49.910 195.820 50.230 195.880 ;
        RECT 52.225 195.820 52.515 195.865 ;
        RECT 49.910 195.680 52.515 195.820 ;
        RECT 49.910 195.620 50.230 195.680 ;
        RECT 52.225 195.635 52.515 195.680 ;
        RECT 54.510 195.820 54.830 195.880 ;
        RECT 60.030 195.820 60.350 195.880 ;
        RECT 80.730 195.820 81.050 195.880 ;
        RECT 54.510 195.680 60.350 195.820 ;
        RECT 54.510 195.620 54.830 195.680 ;
        RECT 60.030 195.620 60.350 195.680 ;
        RECT 66.100 195.680 81.050 195.820 ;
        RECT 25.530 195.480 25.850 195.540 ;
        RECT 31.510 195.480 31.830 195.540 ;
        RECT 33.350 195.480 33.670 195.540 ;
        RECT 36.110 195.480 36.430 195.540 ;
        RECT 25.530 195.340 27.140 195.480 ;
        RECT 25.530 195.280 25.850 195.340 ;
        RECT 22.310 194.940 22.630 195.200 ;
        RECT 26.450 195.140 26.770 195.200 ;
        RECT 26.310 194.940 26.770 195.140 ;
        RECT 21.405 194.665 21.695 194.895 ;
        RECT 21.850 194.800 22.170 194.860 ;
        RECT 23.705 194.800 23.995 194.845 ;
        RECT 21.480 194.520 21.620 194.665 ;
        RECT 21.850 194.660 23.995 194.800 ;
        RECT 21.850 194.600 22.170 194.660 ;
        RECT 23.705 194.615 23.995 194.660 ;
        RECT 25.070 194.600 25.390 194.860 ;
        RECT 25.875 194.800 26.165 194.845 ;
        RECT 26.310 194.800 26.450 194.940 ;
        RECT 27.000 194.845 27.140 195.340 ;
        RECT 31.510 195.340 33.670 195.480 ;
        RECT 31.510 195.280 31.830 195.340 ;
        RECT 33.350 195.280 33.670 195.340 ;
        RECT 34.360 195.340 36.430 195.480 ;
        RECT 34.360 195.185 34.500 195.340 ;
        RECT 36.110 195.280 36.430 195.340 ;
        RECT 38.870 195.280 39.190 195.540 ;
        RECT 42.105 195.480 42.395 195.525 ;
        RECT 47.150 195.480 47.470 195.540 ;
        RECT 42.105 195.340 47.470 195.480 ;
        RECT 42.105 195.295 42.395 195.340 ;
        RECT 47.150 195.280 47.470 195.340 ;
        RECT 50.370 195.480 50.690 195.540 ;
        RECT 50.370 195.340 54.740 195.480 ;
        RECT 50.370 195.280 50.690 195.340 ;
        RECT 27.460 195.000 34.040 195.140 ;
        RECT 27.460 194.860 27.600 195.000 ;
        RECT 25.875 194.660 26.450 194.800 ;
        RECT 25.875 194.615 26.165 194.660 ;
        RECT 26.925 194.615 27.215 194.845 ;
        RECT 21.390 194.260 21.710 194.520 ;
        RECT 22.770 194.260 23.090 194.520 ;
        RECT 26.460 194.275 26.750 194.505 ;
        RECT 27.000 194.460 27.140 194.615 ;
        RECT 27.370 194.600 27.690 194.860 ;
        RECT 28.290 194.600 28.610 194.860 ;
        RECT 30.590 194.600 30.910 194.860 ;
        RECT 31.525 194.615 31.815 194.845 ;
        RECT 32.445 194.615 32.735 194.845 ;
        RECT 32.905 194.800 33.195 194.845 ;
        RECT 33.350 194.800 33.670 194.860 ;
        RECT 32.905 194.660 33.670 194.800 ;
        RECT 33.900 194.800 34.040 195.000 ;
        RECT 34.285 194.955 34.575 195.185 ;
        RECT 38.960 195.140 39.100 195.280 ;
        RECT 36.200 195.000 39.100 195.140 ;
        RECT 41.630 195.140 41.950 195.200 ;
        RECT 44.390 195.140 44.710 195.200 ;
        RECT 41.630 195.000 44.710 195.140 ;
        RECT 34.745 194.800 35.035 194.845 ;
        RECT 33.900 194.660 35.035 194.800 ;
        RECT 32.905 194.615 33.195 194.660 ;
        RECT 28.380 194.460 28.520 194.600 ;
        RECT 27.000 194.320 28.520 194.460 ;
        RECT 29.210 194.460 29.530 194.520 ;
        RECT 31.600 194.460 31.740 194.615 ;
        RECT 29.210 194.320 31.740 194.460 ;
        RECT 32.520 194.460 32.660 194.615 ;
        RECT 33.350 194.600 33.670 194.660 ;
        RECT 34.745 194.615 35.035 194.660 ;
        RECT 35.190 194.800 35.510 194.860 ;
        RECT 36.200 194.845 36.340 195.000 ;
        RECT 41.630 194.940 41.950 195.000 ;
        RECT 44.390 194.940 44.710 195.000 ;
        RECT 49.450 195.140 49.770 195.200 ;
        RECT 54.600 195.185 54.740 195.340 ;
        RECT 53.605 195.140 53.895 195.185 ;
        RECT 49.450 195.000 53.895 195.140 ;
        RECT 49.450 194.940 49.770 195.000 ;
        RECT 53.605 194.955 53.895 195.000 ;
        RECT 54.525 194.955 54.815 195.185 ;
        RECT 62.790 195.140 63.110 195.200 ;
        RECT 55.060 195.000 63.110 195.140 ;
        RECT 35.665 194.800 35.955 194.845 ;
        RECT 35.190 194.660 35.955 194.800 ;
        RECT 35.190 194.600 35.510 194.660 ;
        RECT 35.665 194.615 35.955 194.660 ;
        RECT 36.125 194.615 36.415 194.845 ;
        RECT 36.570 194.600 36.890 194.860 ;
        RECT 37.505 194.800 37.795 194.845 ;
        RECT 38.870 194.800 39.190 194.860 ;
        RECT 37.505 194.660 39.190 194.800 ;
        RECT 37.505 194.615 37.795 194.660 ;
        RECT 38.870 194.600 39.190 194.660 ;
        RECT 39.345 194.800 39.635 194.845 ;
        RECT 39.790 194.800 40.110 194.860 ;
        RECT 39.345 194.660 40.110 194.800 ;
        RECT 39.345 194.615 39.635 194.660 ;
        RECT 39.790 194.600 40.110 194.660 ;
        RECT 41.185 194.800 41.475 194.845 ;
        RECT 43.470 194.800 43.790 194.860 ;
        RECT 41.185 194.660 43.790 194.800 ;
        RECT 41.185 194.615 41.475 194.660 ;
        RECT 43.470 194.600 43.790 194.660 ;
        RECT 45.310 194.800 45.630 194.860 ;
        RECT 47.610 194.800 47.930 194.860 ;
        RECT 53.145 194.800 53.435 194.845 ;
        RECT 45.310 194.660 47.930 194.800 ;
        RECT 45.310 194.600 45.630 194.660 ;
        RECT 47.610 194.600 47.930 194.660 ;
        RECT 48.160 194.660 53.435 194.800 ;
        RECT 40.265 194.460 40.555 194.505 ;
        RECT 32.520 194.320 40.555 194.460 ;
        RECT 20.485 194.120 20.775 194.165 ;
        RECT 26.540 194.120 26.680 194.275 ;
        RECT 29.210 194.260 29.530 194.320 ;
        RECT 40.265 194.275 40.555 194.320 ;
        RECT 40.710 194.460 41.030 194.520 ;
        RECT 48.160 194.460 48.300 194.660 ;
        RECT 53.145 194.615 53.435 194.660 ;
        RECT 54.065 194.800 54.355 194.845 ;
        RECT 55.060 194.800 55.200 195.000 ;
        RECT 62.790 194.940 63.110 195.000 ;
        RECT 54.065 194.660 55.200 194.800 ;
        RECT 55.430 194.800 55.750 194.860 ;
        RECT 61.870 194.800 62.190 194.860 ;
        RECT 66.100 194.845 66.240 195.680 ;
        RECT 80.730 195.620 81.050 195.680 ;
        RECT 86.265 195.820 86.555 195.865 ;
        RECT 87.170 195.820 87.490 195.880 ;
        RECT 86.265 195.680 87.490 195.820 ;
        RECT 86.265 195.635 86.555 195.680 ;
        RECT 87.170 195.620 87.490 195.680 ;
        RECT 75.685 195.480 75.975 195.525 ;
        RECT 84.870 195.480 85.190 195.540 ;
        RECT 75.685 195.340 85.190 195.480 ;
        RECT 75.685 195.295 75.975 195.340 ;
        RECT 84.870 195.280 85.190 195.340 ;
        RECT 70.610 195.140 70.930 195.200 ;
        RECT 71.990 195.140 72.310 195.200 ;
        RECT 78.890 195.140 79.210 195.200 ;
        RECT 67.940 195.000 70.930 195.140 ;
        RECT 55.430 194.660 62.190 194.800 ;
        RECT 54.065 194.615 54.355 194.660 ;
        RECT 40.710 194.320 48.300 194.460 ;
        RECT 26.910 194.120 27.230 194.180 ;
        RECT 20.485 193.980 27.230 194.120 ;
        RECT 20.485 193.935 20.775 193.980 ;
        RECT 26.910 193.920 27.230 193.980 ;
        RECT 27.370 194.120 27.690 194.180 ;
        RECT 28.305 194.120 28.595 194.165 ;
        RECT 27.370 193.980 28.595 194.120 ;
        RECT 27.370 193.920 27.690 193.980 ;
        RECT 28.305 193.935 28.595 193.980 ;
        RECT 30.590 194.120 30.910 194.180 ;
        RECT 33.350 194.120 33.670 194.180 ;
        RECT 30.590 193.980 33.670 194.120 ;
        RECT 30.590 193.920 30.910 193.980 ;
        RECT 33.350 193.920 33.670 193.980 ;
        RECT 33.810 194.120 34.130 194.180 ;
        RECT 37.950 194.120 38.270 194.180 ;
        RECT 33.810 193.980 38.270 194.120 ;
        RECT 33.810 193.920 34.130 193.980 ;
        RECT 37.950 193.920 38.270 193.980 ;
        RECT 38.425 194.120 38.715 194.165 ;
        RECT 39.790 194.120 40.110 194.180 ;
        RECT 38.425 193.980 40.110 194.120 ;
        RECT 40.340 194.120 40.480 194.275 ;
        RECT 40.710 194.260 41.030 194.320 ;
        RECT 51.305 194.275 51.595 194.505 ;
        RECT 51.750 194.460 52.070 194.520 ;
        RECT 54.140 194.460 54.280 194.615 ;
        RECT 55.430 194.600 55.750 194.660 ;
        RECT 61.870 194.600 62.190 194.660 ;
        RECT 66.025 194.615 66.315 194.845 ;
        RECT 66.485 194.800 66.775 194.845 ;
        RECT 67.940 194.800 68.080 195.000 ;
        RECT 70.610 194.940 70.930 195.000 ;
        RECT 71.160 195.000 72.310 195.140 ;
        RECT 71.160 194.845 71.300 195.000 ;
        RECT 71.990 194.940 72.310 195.000 ;
        RECT 72.540 195.000 79.210 195.140 ;
        RECT 66.485 194.660 68.080 194.800 ;
        RECT 66.485 194.615 66.775 194.660 ;
        RECT 71.085 194.615 71.375 194.845 ;
        RECT 71.530 194.600 71.850 194.860 ;
        RECT 72.540 194.845 72.680 195.000 ;
        RECT 78.890 194.940 79.210 195.000 ;
        RECT 72.465 194.615 72.755 194.845 ;
        RECT 72.910 194.600 73.230 194.860 ;
        RECT 82.570 194.600 82.890 194.860 ;
        RECT 83.030 194.800 83.350 194.860 ;
        RECT 84.885 194.800 85.175 194.845 ;
        RECT 83.030 194.660 85.175 194.800 ;
        RECT 83.030 194.600 83.350 194.660 ;
        RECT 84.885 194.615 85.175 194.660 ;
        RECT 85.330 194.600 85.650 194.860 ;
        RECT 86.710 194.600 87.030 194.860 ;
        RECT 51.750 194.320 54.280 194.460 ;
        RECT 41.170 194.120 41.490 194.180 ;
        RECT 43.930 194.120 44.250 194.180 ;
        RECT 40.340 193.980 44.250 194.120 ;
        RECT 38.425 193.935 38.715 193.980 ;
        RECT 39.790 193.920 40.110 193.980 ;
        RECT 41.170 193.920 41.490 193.980 ;
        RECT 43.930 193.920 44.250 193.980 ;
        RECT 44.390 194.120 44.710 194.180 ;
        RECT 44.865 194.120 45.155 194.165 ;
        RECT 46.230 194.120 46.550 194.180 ;
        RECT 44.390 193.980 46.550 194.120 ;
        RECT 44.390 193.920 44.710 193.980 ;
        RECT 44.865 193.935 45.155 193.980 ;
        RECT 46.230 193.920 46.550 193.980 ;
        RECT 46.690 194.120 47.010 194.180 ;
        RECT 49.910 194.120 50.230 194.180 ;
        RECT 46.690 193.980 50.230 194.120 ;
        RECT 51.380 194.120 51.520 194.275 ;
        RECT 51.750 194.260 52.070 194.320 ;
        RECT 57.285 194.275 57.575 194.505 ;
        RECT 66.560 194.320 68.080 194.460 ;
        RECT 57.360 194.120 57.500 194.275 ;
        RECT 66.560 194.180 66.700 194.320 ;
        RECT 64.170 194.120 64.490 194.180 ;
        RECT 51.380 193.980 64.490 194.120 ;
        RECT 46.690 193.920 47.010 193.980 ;
        RECT 49.910 193.920 50.230 193.980 ;
        RECT 64.170 193.920 64.490 193.980 ;
        RECT 66.470 193.920 66.790 194.180 ;
        RECT 67.390 193.920 67.710 194.180 ;
        RECT 67.940 194.165 68.080 194.320 ;
        RECT 68.310 194.260 68.630 194.520 ;
        RECT 69.245 194.460 69.535 194.505 ;
        RECT 69.245 194.320 74.750 194.460 ;
        RECT 69.245 194.275 69.535 194.320 ;
        RECT 67.865 193.935 68.155 194.165 ;
        RECT 68.770 194.120 69.090 194.180 ;
        RECT 70.165 194.120 70.455 194.165 ;
        RECT 68.770 193.980 70.455 194.120 ;
        RECT 74.610 194.120 74.750 194.320 ;
        RECT 82.110 194.260 82.430 194.520 ;
        RECT 82.660 194.460 82.800 194.600 ;
        RECT 82.660 194.320 83.260 194.460 ;
        RECT 82.570 194.120 82.890 194.180 ;
        RECT 83.120 194.165 83.260 194.320 ;
        RECT 74.610 193.980 82.890 194.120 ;
        RECT 68.770 193.920 69.090 193.980 ;
        RECT 70.165 193.935 70.455 193.980 ;
        RECT 82.570 193.920 82.890 193.980 ;
        RECT 83.045 193.935 83.335 194.165 ;
        RECT 87.170 193.920 87.490 194.180 ;
        RECT 18.100 193.300 89.400 193.780 ;
        RECT 20.930 193.100 21.250 193.160 ;
        RECT 22.785 193.100 23.075 193.145 ;
        RECT 20.930 192.960 23.075 193.100 ;
        RECT 20.930 192.900 21.250 192.960 ;
        RECT 22.785 192.915 23.075 192.960 ;
        RECT 23.230 193.100 23.550 193.160 ;
        RECT 24.625 193.100 24.915 193.145 ;
        RECT 25.530 193.100 25.850 193.160 ;
        RECT 23.230 192.960 25.850 193.100 ;
        RECT 23.230 192.900 23.550 192.960 ;
        RECT 24.625 192.915 24.915 192.960 ;
        RECT 25.530 192.900 25.850 192.960 ;
        RECT 27.830 193.100 28.150 193.160 ;
        RECT 28.765 193.100 29.055 193.145 ;
        RECT 37.030 193.100 37.350 193.160 ;
        RECT 27.830 192.960 29.055 193.100 ;
        RECT 27.830 192.900 28.150 192.960 ;
        RECT 28.765 192.915 29.055 192.960 ;
        RECT 29.760 192.960 33.580 193.100 ;
        RECT 17.250 192.760 17.570 192.820 ;
        RECT 29.760 192.760 29.900 192.960 ;
        RECT 17.250 192.620 21.620 192.760 ;
        RECT 17.250 192.560 17.570 192.620 ;
        RECT 20.930 192.220 21.250 192.480 ;
        RECT 21.480 192.465 21.620 192.620 ;
        RECT 27.920 192.620 29.900 192.760 ;
        RECT 21.405 192.235 21.695 192.465 ;
        RECT 23.705 192.420 23.995 192.465 ;
        RECT 24.610 192.420 24.930 192.480 ;
        RECT 23.705 192.280 24.930 192.420 ;
        RECT 23.705 192.235 23.995 192.280 ;
        RECT 20.010 192.080 20.330 192.140 ;
        RECT 23.780 192.080 23.920 192.235 ;
        RECT 24.610 192.220 24.930 192.280 ;
        RECT 25.085 192.235 25.375 192.465 ;
        RECT 26.925 192.420 27.215 192.465 ;
        RECT 27.370 192.420 27.690 192.480 ;
        RECT 27.920 192.465 28.060 192.620 ;
        RECT 30.590 192.560 30.910 192.820 ;
        RECT 26.925 192.280 27.690 192.420 ;
        RECT 26.925 192.235 27.215 192.280 ;
        RECT 20.010 191.940 23.920 192.080 ;
        RECT 20.010 191.880 20.330 191.940 ;
        RECT 25.160 191.740 25.300 192.235 ;
        RECT 27.370 192.220 27.690 192.280 ;
        RECT 27.845 192.235 28.135 192.465 ;
        RECT 28.305 192.235 28.595 192.465 ;
        RECT 28.750 192.420 29.070 192.480 ;
        RECT 29.685 192.420 29.975 192.465 ;
        RECT 28.750 192.280 29.975 192.420 ;
        RECT 25.530 192.080 25.850 192.140 ;
        RECT 27.920 192.080 28.060 192.235 ;
        RECT 25.530 191.940 28.060 192.080 ;
        RECT 28.380 192.080 28.520 192.235 ;
        RECT 28.750 192.220 29.070 192.280 ;
        RECT 29.685 192.235 29.975 192.280 ;
        RECT 31.510 192.220 31.830 192.480 ;
        RECT 31.970 192.420 32.290 192.480 ;
        RECT 33.440 192.465 33.580 192.960 ;
        RECT 33.900 192.960 37.350 193.100 ;
        RECT 33.900 192.820 34.040 192.960 ;
        RECT 37.030 192.900 37.350 192.960 ;
        RECT 40.265 192.915 40.555 193.145 ;
        RECT 43.025 193.100 43.315 193.145 ;
        RECT 45.310 193.100 45.630 193.160 ;
        RECT 50.370 193.100 50.690 193.160 ;
        RECT 43.025 192.960 45.630 193.100 ;
        RECT 43.025 192.915 43.315 192.960 ;
        RECT 33.810 192.560 34.130 192.820 ;
        RECT 34.285 192.760 34.575 192.805 ;
        RECT 39.790 192.760 40.110 192.820 ;
        RECT 34.285 192.620 40.110 192.760 ;
        RECT 40.340 192.760 40.480 192.915 ;
        RECT 45.310 192.900 45.630 192.960 ;
        RECT 45.860 192.960 50.690 193.100 ;
        RECT 45.860 192.805 46.000 192.960 ;
        RECT 50.370 192.900 50.690 192.960 ;
        RECT 53.145 193.100 53.435 193.145 ;
        RECT 54.050 193.100 54.370 193.160 ;
        RECT 53.145 192.960 54.370 193.100 ;
        RECT 53.145 192.915 53.435 192.960 ;
        RECT 54.050 192.900 54.370 192.960 ;
        RECT 62.805 192.915 63.095 193.145 ;
        RECT 67.850 193.100 68.170 193.160 ;
        RECT 71.085 193.100 71.375 193.145 ;
        RECT 86.710 193.100 87.030 193.160 ;
        RECT 67.850 192.960 71.375 193.100 ;
        RECT 40.340 192.620 45.540 192.760 ;
        RECT 34.285 192.575 34.575 192.620 ;
        RECT 39.790 192.560 40.110 192.620 ;
        RECT 45.400 192.480 45.540 192.620 ;
        RECT 45.785 192.575 46.075 192.805 ;
        RECT 46.245 192.760 46.535 192.805 ;
        RECT 46.690 192.760 47.010 192.820 ;
        RECT 46.245 192.620 47.010 192.760 ;
        RECT 46.245 192.575 46.535 192.620 ;
        RECT 46.690 192.560 47.010 192.620 ;
        RECT 47.610 192.760 47.930 192.820 ;
        RECT 51.750 192.760 52.070 192.820 ;
        RECT 47.610 192.620 52.070 192.760 ;
        RECT 47.610 192.560 47.930 192.620 ;
        RECT 51.750 192.560 52.070 192.620 ;
        RECT 60.030 192.760 60.350 192.820 ;
        RECT 62.880 192.760 63.020 192.915 ;
        RECT 67.850 192.900 68.170 192.960 ;
        RECT 71.085 192.915 71.375 192.960 ;
        RECT 74.610 192.960 87.030 193.100 ;
        RECT 74.610 192.760 74.750 192.960 ;
        RECT 86.710 192.900 87.030 192.960 ;
        RECT 87.170 192.760 87.490 192.820 ;
        RECT 60.030 192.620 74.750 192.760 ;
        RECT 76.220 192.620 87.490 192.760 ;
        RECT 60.030 192.560 60.350 192.620 ;
        RECT 32.905 192.420 33.195 192.465 ;
        RECT 31.970 192.280 33.195 192.420 ;
        RECT 31.970 192.220 32.290 192.280 ;
        RECT 32.905 192.235 33.195 192.280 ;
        RECT 33.365 192.420 33.655 192.465 ;
        RECT 35.650 192.420 35.970 192.480 ;
        RECT 33.365 192.280 35.970 192.420 ;
        RECT 33.365 192.235 33.655 192.280 ;
        RECT 35.650 192.220 35.970 192.280 ;
        RECT 36.110 192.420 36.430 192.480 ;
        RECT 36.585 192.420 36.875 192.465 ;
        RECT 36.110 192.280 36.875 192.420 ;
        RECT 36.110 192.220 36.430 192.280 ;
        RECT 36.585 192.235 36.875 192.280 ;
        RECT 32.060 192.080 32.200 192.220 ;
        RECT 28.380 191.940 32.200 192.080 ;
        RECT 36.660 192.080 36.800 192.235 ;
        RECT 37.490 192.220 37.810 192.480 ;
        RECT 40.725 192.420 41.015 192.465 ;
        RECT 43.010 192.420 43.330 192.480 ;
        RECT 40.725 192.280 43.330 192.420 ;
        RECT 40.725 192.235 41.015 192.280 ;
        RECT 43.010 192.220 43.330 192.280 ;
        RECT 45.310 192.220 45.630 192.480 ;
        RECT 47.150 192.220 47.470 192.480 ;
        RECT 48.545 192.440 48.835 192.465 ;
        RECT 48.160 192.300 48.835 192.440 ;
        RECT 37.950 192.080 38.270 192.140 ;
        RECT 36.660 191.940 38.270 192.080 ;
        RECT 25.530 191.880 25.850 191.940 ;
        RECT 37.950 191.880 38.270 191.940 ;
        RECT 39.330 192.080 39.650 192.140 ;
        RECT 42.105 192.080 42.395 192.125 ;
        RECT 44.390 192.080 44.710 192.140 ;
        RECT 39.330 191.940 40.020 192.080 ;
        RECT 39.330 191.880 39.650 191.940 ;
        RECT 28.750 191.740 29.070 191.800 ;
        RECT 25.160 191.600 29.070 191.740 ;
        RECT 28.750 191.540 29.070 191.600 ;
        RECT 31.970 191.740 32.290 191.800 ;
        RECT 32.445 191.740 32.735 191.785 ;
        RECT 31.970 191.600 32.735 191.740 ;
        RECT 31.970 191.540 32.290 191.600 ;
        RECT 32.445 191.555 32.735 191.600 ;
        RECT 34.285 191.740 34.575 191.785 ;
        RECT 36.110 191.740 36.430 191.800 ;
        RECT 34.285 191.600 36.430 191.740 ;
        RECT 34.285 191.555 34.575 191.600 ;
        RECT 36.110 191.540 36.430 191.600 ;
        RECT 37.030 191.740 37.350 191.800 ;
        RECT 39.880 191.785 40.020 191.940 ;
        RECT 42.105 191.940 44.710 192.080 ;
        RECT 48.160 192.080 48.300 192.300 ;
        RECT 48.545 192.235 48.835 192.300 ;
        RECT 49.005 192.420 49.295 192.465 ;
        RECT 49.910 192.420 50.230 192.480 ;
        RECT 49.005 192.280 50.230 192.420 ;
        RECT 49.005 192.235 49.295 192.280 ;
        RECT 49.910 192.220 50.230 192.280 ;
        RECT 50.370 192.220 50.690 192.480 ;
        RECT 59.570 192.220 59.890 192.480 ;
        RECT 69.245 192.420 69.535 192.465 ;
        RECT 71.070 192.420 71.390 192.480 ;
        RECT 76.220 192.465 76.360 192.620 ;
        RECT 87.170 192.560 87.490 192.620 ;
        RECT 69.245 192.280 71.390 192.420 ;
        RECT 69.245 192.235 69.535 192.280 ;
        RECT 71.070 192.220 71.390 192.280 ;
        RECT 71.620 192.280 72.680 192.420 ;
        RECT 58.190 192.080 58.510 192.140 ;
        RECT 48.160 191.940 58.510 192.080 ;
        RECT 42.105 191.895 42.395 191.940 ;
        RECT 44.390 191.880 44.710 191.940 ;
        RECT 58.190 191.880 58.510 191.940 ;
        RECT 67.850 192.080 68.170 192.140 ;
        RECT 70.150 192.080 70.470 192.140 ;
        RECT 67.850 191.940 70.470 192.080 ;
        RECT 67.850 191.880 68.170 191.940 ;
        RECT 70.150 191.880 70.470 191.940 ;
        RECT 37.030 191.600 39.560 191.740 ;
        RECT 37.030 191.540 37.350 191.600 ;
        RECT 16.790 191.400 17.110 191.460 ;
        RECT 20.025 191.400 20.315 191.445 ;
        RECT 16.790 191.260 20.315 191.400 ;
        RECT 16.790 191.200 17.110 191.260 ;
        RECT 20.025 191.215 20.315 191.260 ;
        RECT 21.390 191.400 21.710 191.460 ;
        RECT 22.325 191.400 22.615 191.445 ;
        RECT 22.770 191.400 23.090 191.460 ;
        RECT 21.390 191.260 23.090 191.400 ;
        RECT 21.390 191.200 21.710 191.260 ;
        RECT 22.325 191.215 22.615 191.260 ;
        RECT 22.770 191.200 23.090 191.260 ;
        RECT 26.005 191.400 26.295 191.445 ;
        RECT 26.450 191.400 26.770 191.460 ;
        RECT 26.005 191.260 26.770 191.400 ;
        RECT 26.005 191.215 26.295 191.260 ;
        RECT 26.450 191.200 26.770 191.260 ;
        RECT 28.290 191.400 28.610 191.460 ;
        RECT 35.665 191.400 35.955 191.445 ;
        RECT 38.410 191.400 38.730 191.460 ;
        RECT 28.290 191.260 38.730 191.400 ;
        RECT 39.420 191.400 39.560 191.600 ;
        RECT 39.805 191.555 40.095 191.785 ;
        RECT 41.185 191.740 41.475 191.785 ;
        RECT 41.630 191.740 41.950 191.800 ;
        RECT 47.610 191.740 47.930 191.800 ;
        RECT 41.185 191.600 41.950 191.740 ;
        RECT 41.185 191.555 41.475 191.600 ;
        RECT 41.630 191.540 41.950 191.600 ;
        RECT 43.560 191.600 47.930 191.740 ;
        RECT 43.560 191.400 43.700 191.600 ;
        RECT 47.610 191.540 47.930 191.600 ;
        RECT 49.925 191.740 50.215 191.785 ;
        RECT 71.620 191.740 71.760 192.280 ;
        RECT 72.005 191.895 72.295 192.125 ;
        RECT 49.925 191.600 71.760 191.740 ;
        RECT 49.925 191.555 50.215 191.600 ;
        RECT 39.420 191.260 43.700 191.400 ;
        RECT 43.930 191.400 44.250 191.460 ;
        RECT 44.405 191.400 44.695 191.445 ;
        RECT 43.930 191.260 44.695 191.400 ;
        RECT 28.290 191.200 28.610 191.260 ;
        RECT 35.665 191.215 35.955 191.260 ;
        RECT 38.410 191.200 38.730 191.260 ;
        RECT 43.930 191.200 44.250 191.260 ;
        RECT 44.405 191.215 44.695 191.260 ;
        RECT 50.370 191.400 50.690 191.460 ;
        RECT 56.810 191.400 57.130 191.460 ;
        RECT 50.370 191.260 57.130 191.400 ;
        RECT 50.370 191.200 50.690 191.260 ;
        RECT 56.810 191.200 57.130 191.260 ;
        RECT 57.730 191.400 58.050 191.460 ;
        RECT 60.950 191.400 61.270 191.460 ;
        RECT 57.730 191.260 61.270 191.400 ;
        RECT 57.730 191.200 58.050 191.260 ;
        RECT 60.950 191.200 61.270 191.260 ;
        RECT 61.870 191.400 62.190 191.460 ;
        RECT 72.080 191.400 72.220 191.895 ;
        RECT 72.540 191.740 72.680 192.280 ;
        RECT 76.145 192.235 76.435 192.465 ;
        RECT 76.590 192.220 76.910 192.480 ;
        RECT 77.510 192.220 77.830 192.480 ;
        RECT 87.630 192.220 87.950 192.480 ;
        RECT 74.750 192.080 75.070 192.140 ;
        RECT 75.225 192.080 75.515 192.125 ;
        RECT 74.750 191.940 75.515 192.080 ;
        RECT 74.750 191.880 75.070 191.940 ;
        RECT 75.225 191.895 75.515 191.940 ;
        RECT 75.685 192.080 75.975 192.125 ;
        RECT 75.685 191.940 76.085 192.080 ;
        RECT 75.685 191.895 75.975 191.940 ;
        RECT 75.760 191.740 75.900 191.895 ;
        RECT 79.810 191.740 80.130 191.800 ;
        RECT 72.540 191.600 80.130 191.740 ;
        RECT 79.810 191.540 80.130 191.600 ;
        RECT 81.205 191.740 81.495 191.785 ;
        RECT 81.650 191.740 81.970 191.800 ;
        RECT 81.205 191.600 81.970 191.740 ;
        RECT 81.205 191.555 81.495 191.600 ;
        RECT 81.650 191.540 81.970 191.600 ;
        RECT 82.110 191.740 82.430 191.800 ;
        RECT 84.410 191.740 84.730 191.800 ;
        RECT 82.110 191.600 84.730 191.740 ;
        RECT 82.110 191.540 82.430 191.600 ;
        RECT 84.410 191.540 84.730 191.600 ;
        RECT 61.870 191.260 72.220 191.400 ;
        RECT 72.925 191.400 73.215 191.445 ;
        RECT 73.370 191.400 73.690 191.460 ;
        RECT 72.925 191.260 73.690 191.400 ;
        RECT 61.870 191.200 62.190 191.260 ;
        RECT 72.925 191.215 73.215 191.260 ;
        RECT 73.370 191.200 73.690 191.260 ;
        RECT 74.290 191.200 74.610 191.460 ;
        RECT 18.100 190.580 89.400 191.060 ;
        RECT 23.245 190.380 23.535 190.425 ;
        RECT 23.690 190.380 24.010 190.440 ;
        RECT 23.245 190.240 24.010 190.380 ;
        RECT 23.245 190.195 23.535 190.240 ;
        RECT 23.690 190.180 24.010 190.240 ;
        RECT 29.210 190.380 29.530 190.440 ;
        RECT 41.630 190.380 41.950 190.440 ;
        RECT 29.210 190.240 41.950 190.380 ;
        RECT 29.210 190.180 29.530 190.240 ;
        RECT 41.630 190.180 41.950 190.240 ;
        RECT 42.550 190.180 42.870 190.440 ;
        RECT 43.470 190.380 43.790 190.440 ;
        RECT 50.370 190.380 50.690 190.440 ;
        RECT 43.470 190.240 50.690 190.380 ;
        RECT 43.470 190.180 43.790 190.240 ;
        RECT 50.370 190.180 50.690 190.240 ;
        RECT 52.670 190.180 52.990 190.440 ;
        RECT 54.050 190.380 54.370 190.440 ;
        RECT 55.430 190.380 55.750 190.440 ;
        RECT 54.050 190.240 55.750 190.380 ;
        RECT 54.050 190.180 54.370 190.240 ;
        RECT 55.430 190.180 55.750 190.240 ;
        RECT 56.365 190.380 56.655 190.425 ;
        RECT 56.810 190.380 57.130 190.440 ;
        RECT 56.365 190.240 57.130 190.380 ;
        RECT 56.365 190.195 56.655 190.240 ;
        RECT 56.810 190.180 57.130 190.240 ;
        RECT 57.730 190.380 58.050 190.440 ;
        RECT 60.505 190.380 60.795 190.425 ;
        RECT 71.530 190.380 71.850 190.440 ;
        RECT 57.730 190.240 60.795 190.380 ;
        RECT 57.730 190.180 58.050 190.240 ;
        RECT 60.505 190.195 60.795 190.240 ;
        RECT 61.960 190.240 71.850 190.380 ;
        RECT 19.550 190.040 19.870 190.100 ;
        RECT 25.545 190.040 25.835 190.085 ;
        RECT 19.550 189.900 25.835 190.040 ;
        RECT 19.550 189.840 19.870 189.900 ;
        RECT 25.545 189.855 25.835 189.900 ;
        RECT 25.990 190.040 26.310 190.100 ;
        RECT 28.765 190.040 29.055 190.085 ;
        RECT 37.490 190.040 37.810 190.100 ;
        RECT 37.965 190.040 38.255 190.085 ;
        RECT 25.990 189.900 37.260 190.040 ;
        RECT 25.990 189.840 26.310 189.900 ;
        RECT 28.765 189.855 29.055 189.900 ;
        RECT 25.070 189.700 25.390 189.760 ;
        RECT 21.480 189.560 25.390 189.700 ;
        RECT 20.930 189.160 21.250 189.420 ;
        RECT 21.480 189.405 21.620 189.560 ;
        RECT 25.070 189.500 25.390 189.560 ;
        RECT 31.510 189.700 31.830 189.760 ;
        RECT 33.350 189.700 33.670 189.760 ;
        RECT 31.510 189.560 33.670 189.700 ;
        RECT 31.510 189.500 31.830 189.560 ;
        RECT 33.350 189.500 33.670 189.560 ;
        RECT 34.730 189.700 35.050 189.760 ;
        RECT 35.665 189.700 35.955 189.745 ;
        RECT 36.110 189.700 36.430 189.760 ;
        RECT 34.730 189.560 36.430 189.700 ;
        RECT 37.120 189.700 37.260 189.900 ;
        RECT 37.490 189.900 38.255 190.040 ;
        RECT 37.490 189.840 37.810 189.900 ;
        RECT 37.965 189.855 38.255 189.900 ;
        RECT 38.870 189.840 39.190 190.100 ;
        RECT 39.330 190.040 39.650 190.100 ;
        RECT 39.805 190.040 40.095 190.085 ;
        RECT 39.330 189.900 40.095 190.040 ;
        RECT 39.330 189.840 39.650 189.900 ;
        RECT 39.805 189.855 40.095 189.900 ;
        RECT 44.850 190.040 45.170 190.100 ;
        RECT 47.150 190.040 47.470 190.100 ;
        RECT 50.830 190.040 51.150 190.100 ;
        RECT 44.850 189.900 47.470 190.040 ;
        RECT 44.850 189.840 45.170 189.900 ;
        RECT 47.150 189.840 47.470 189.900 ;
        RECT 48.160 189.900 51.150 190.040 ;
        RECT 37.120 189.560 38.180 189.700 ;
        RECT 34.730 189.500 35.050 189.560 ;
        RECT 35.665 189.515 35.955 189.560 ;
        RECT 36.110 189.500 36.430 189.560 ;
        RECT 21.405 189.175 21.695 189.405 ;
        RECT 22.310 189.360 22.630 189.420 ;
        RECT 22.785 189.360 23.075 189.405 ;
        RECT 23.230 189.360 23.550 189.420 ;
        RECT 22.310 189.220 23.550 189.360 ;
        RECT 22.310 189.160 22.630 189.220 ;
        RECT 22.785 189.175 23.075 189.220 ;
        RECT 23.230 189.160 23.550 189.220 ;
        RECT 24.165 189.360 24.455 189.405 ;
        RECT 28.750 189.360 29.070 189.420 ;
        RECT 24.165 189.220 29.070 189.360 ;
        RECT 24.165 189.175 24.455 189.220 ;
        RECT 28.750 189.160 29.070 189.220 ;
        RECT 29.685 189.175 29.975 189.405 ;
        RECT 21.020 189.020 21.160 189.160 ;
        RECT 26.005 189.020 26.295 189.065 ;
        RECT 21.020 188.880 22.080 189.020 ;
        RECT 20.485 188.680 20.775 188.725 ;
        RECT 20.930 188.680 21.250 188.740 ;
        RECT 21.940 188.725 22.080 188.880 ;
        RECT 25.160 188.880 26.295 189.020 ;
        RECT 20.485 188.540 21.250 188.680 ;
        RECT 20.485 188.495 20.775 188.540 ;
        RECT 20.930 188.480 21.250 188.540 ;
        RECT 21.865 188.495 22.155 188.725 ;
        RECT 24.610 188.680 24.930 188.740 ;
        RECT 25.160 188.680 25.300 188.880 ;
        RECT 26.005 188.835 26.295 188.880 ;
        RECT 26.450 189.020 26.770 189.080 ;
        RECT 26.925 189.020 27.215 189.065 ;
        RECT 26.450 188.880 27.215 189.020 ;
        RECT 29.760 189.020 29.900 189.175 ;
        RECT 37.030 189.160 37.350 189.420 ;
        RECT 30.130 189.020 30.450 189.080 ;
        RECT 29.760 188.880 30.450 189.020 ;
        RECT 38.040 189.020 38.180 189.560 ;
        RECT 38.425 189.360 38.715 189.405 ;
        RECT 38.960 189.360 39.100 189.840 ;
        RECT 38.425 189.220 39.100 189.360 ;
        RECT 38.425 189.175 38.715 189.220 ;
        RECT 39.790 189.160 40.110 189.420 ;
        RECT 43.470 189.360 43.790 189.420 ;
        RECT 48.160 189.360 48.300 189.900 ;
        RECT 50.830 189.840 51.150 189.900 ;
        RECT 51.290 189.840 51.610 190.100 ;
        RECT 51.380 189.700 51.520 189.840 ;
        RECT 52.760 189.745 52.900 190.180 ;
        RECT 49.540 189.560 51.520 189.700 ;
        RECT 43.470 189.220 48.300 189.360 ;
        RECT 43.470 189.160 43.790 189.220 ;
        RECT 48.990 189.160 49.310 189.420 ;
        RECT 49.540 189.405 49.680 189.560 ;
        RECT 52.685 189.515 52.975 189.745 ;
        RECT 49.465 189.175 49.755 189.405 ;
        RECT 50.385 189.175 50.675 189.405 ;
        RECT 46.690 189.020 47.010 189.080 ;
        RECT 38.040 188.880 47.010 189.020 ;
        RECT 26.450 188.820 26.770 188.880 ;
        RECT 26.925 188.835 27.215 188.880 ;
        RECT 30.130 188.820 30.450 188.880 ;
        RECT 46.690 188.820 47.010 188.880 ;
        RECT 50.460 188.740 50.600 189.175 ;
        RECT 50.830 189.160 51.150 189.420 ;
        RECT 51.390 189.360 51.680 189.405 ;
        RECT 51.390 189.220 51.980 189.360 ;
        RECT 51.390 189.175 51.680 189.220 ;
        RECT 51.840 189.020 51.980 189.220 ;
        RECT 53.130 189.160 53.450 189.420 ;
        RECT 54.140 189.405 54.280 190.180 ;
        RECT 60.950 190.040 61.270 190.100 ;
        RECT 55.060 189.900 61.270 190.040 ;
        RECT 55.060 189.405 55.200 189.900 ;
        RECT 60.950 189.840 61.270 189.900 ;
        RECT 61.960 189.700 62.100 190.240 ;
        RECT 71.530 190.180 71.850 190.240 ;
        RECT 83.490 190.380 83.810 190.440 ;
        RECT 84.410 190.380 84.730 190.440 ;
        RECT 83.490 190.240 84.730 190.380 ;
        RECT 83.490 190.180 83.810 190.240 ;
        RECT 84.410 190.180 84.730 190.240 ;
        RECT 85.330 190.380 85.650 190.440 ;
        RECT 86.725 190.380 87.015 190.425 ;
        RECT 85.330 190.240 87.015 190.380 ;
        RECT 85.330 190.180 85.650 190.240 ;
        RECT 86.725 190.195 87.015 190.240 ;
        RECT 78.890 190.040 79.210 190.100 ;
        RECT 78.890 189.900 87.860 190.040 ;
        RECT 78.890 189.840 79.210 189.900 ;
        RECT 56.900 189.560 62.100 189.700 ;
        RECT 62.345 189.740 62.635 189.745 ;
        RECT 62.345 189.700 63.480 189.740 ;
        RECT 68.310 189.700 68.630 189.760 ;
        RECT 77.510 189.700 77.830 189.760 ;
        RECT 81.190 189.700 81.510 189.760 ;
        RECT 62.345 189.600 81.510 189.700 ;
        RECT 53.935 189.220 54.280 189.405 ;
        RECT 53.935 189.175 54.225 189.220 ;
        RECT 54.985 189.175 55.275 189.405 ;
        RECT 55.445 189.360 55.735 189.405 ;
        RECT 56.350 189.360 56.670 189.420 ;
        RECT 55.445 189.220 56.670 189.360 ;
        RECT 55.445 189.175 55.735 189.220 ;
        RECT 56.350 189.160 56.670 189.220 ;
        RECT 52.670 189.020 52.990 189.080 ;
        RECT 51.840 188.880 52.990 189.020 ;
        RECT 52.670 188.820 52.990 188.880 ;
        RECT 54.510 188.820 54.830 189.080 ;
        RECT 24.610 188.540 25.300 188.680 ;
        RECT 27.845 188.680 28.135 188.725 ;
        RECT 28.290 188.680 28.610 188.740 ;
        RECT 27.845 188.540 28.610 188.680 ;
        RECT 24.610 188.480 24.930 188.540 ;
        RECT 27.845 188.495 28.135 188.540 ;
        RECT 28.290 188.480 28.610 188.540 ;
        RECT 29.210 188.680 29.530 188.740 ;
        RECT 32.445 188.680 32.735 188.725 ;
        RECT 29.210 188.540 32.735 188.680 ;
        RECT 29.210 188.480 29.530 188.540 ;
        RECT 32.445 188.495 32.735 188.540 ;
        RECT 34.270 188.480 34.590 188.740 ;
        RECT 34.745 188.680 35.035 188.725 ;
        RECT 35.190 188.680 35.510 188.740 ;
        RECT 34.745 188.540 35.510 188.680 ;
        RECT 34.745 188.495 35.035 188.540 ;
        RECT 35.190 188.480 35.510 188.540 ;
        RECT 35.650 188.680 35.970 188.740 ;
        RECT 38.885 188.680 39.175 188.725 ;
        RECT 35.650 188.540 39.175 188.680 ;
        RECT 35.650 188.480 35.970 188.540 ;
        RECT 38.885 188.495 39.175 188.540 ;
        RECT 50.370 188.480 50.690 188.740 ;
        RECT 51.290 188.680 51.610 188.740 ;
        RECT 56.900 188.680 57.040 189.560 ;
        RECT 62.345 189.515 62.635 189.600 ;
        RECT 63.340 189.560 81.510 189.600 ;
        RECT 68.310 189.500 68.630 189.560 ;
        RECT 77.510 189.500 77.830 189.560 ;
        RECT 81.190 189.500 81.510 189.560 ;
        RECT 83.030 189.700 83.350 189.760 ;
        RECT 86.265 189.700 86.555 189.745 ;
        RECT 83.030 189.560 86.555 189.700 ;
        RECT 83.030 189.500 83.350 189.560 ;
        RECT 86.265 189.515 86.555 189.560 ;
        RECT 59.110 189.160 59.430 189.420 ;
        RECT 60.965 189.360 61.255 189.405 ;
        RECT 61.410 189.360 61.730 189.420 ;
        RECT 60.965 189.220 61.730 189.360 ;
        RECT 60.965 189.175 61.255 189.220 ;
        RECT 51.290 188.540 57.040 188.680 ;
        RECT 61.040 188.680 61.180 189.175 ;
        RECT 61.410 189.160 61.730 189.220 ;
        RECT 61.870 189.160 62.190 189.420 ;
        RECT 62.985 189.230 63.275 189.375 ;
        RECT 62.985 189.145 63.480 189.230 ;
        RECT 63.710 189.160 64.030 189.420 ;
        RECT 64.170 189.160 64.490 189.420 ;
        RECT 71.530 189.360 71.850 189.420 ;
        RECT 72.925 189.360 73.215 189.405 ;
        RECT 82.570 189.360 82.890 189.420 ;
        RECT 84.425 189.360 84.715 189.405 ;
        RECT 71.530 189.220 78.200 189.360 ;
        RECT 71.530 189.160 71.850 189.220 ;
        RECT 72.925 189.175 73.215 189.220 ;
        RECT 63.060 189.090 63.480 189.145 ;
        RECT 63.340 189.020 63.480 189.090 ;
        RECT 77.510 189.020 77.830 189.080 ;
        RECT 63.340 188.880 77.830 189.020 ;
        RECT 77.510 188.820 77.830 188.880 ;
        RECT 69.690 188.680 70.010 188.740 ;
        RECT 61.040 188.540 70.010 188.680 ;
        RECT 51.290 188.480 51.610 188.540 ;
        RECT 69.690 188.480 70.010 188.540 ;
        RECT 71.070 188.680 71.390 188.740 ;
        RECT 74.765 188.680 75.055 188.725 ;
        RECT 71.070 188.540 75.055 188.680 ;
        RECT 78.060 188.680 78.200 189.220 ;
        RECT 82.570 189.220 84.715 189.360 ;
        RECT 82.570 189.160 82.890 189.220 ;
        RECT 84.425 189.175 84.715 189.220 ;
        RECT 87.170 189.160 87.490 189.420 ;
        RECT 87.720 189.405 87.860 189.900 ;
        RECT 87.645 189.175 87.935 189.405 ;
        RECT 82.110 188.820 82.430 189.080 ;
        RECT 83.045 189.020 83.335 189.065 ;
        RECT 83.045 188.880 84.180 189.020 ;
        RECT 83.045 188.835 83.335 188.880 ;
        RECT 83.505 188.680 83.795 188.725 ;
        RECT 78.060 188.540 83.795 188.680 ;
        RECT 84.040 188.680 84.180 188.880 ;
        RECT 85.330 188.820 85.650 189.080 ;
        RECT 86.710 188.680 87.030 188.740 ;
        RECT 84.040 188.540 87.030 188.680 ;
        RECT 71.070 188.480 71.390 188.540 ;
        RECT 74.765 188.495 75.055 188.540 ;
        RECT 83.505 188.495 83.795 188.540 ;
        RECT 86.710 188.480 87.030 188.540 ;
        RECT 18.100 187.860 89.400 188.340 ;
        RECT 16.790 187.660 17.110 187.720 ;
        RECT 20.025 187.660 20.315 187.705 ;
        RECT 24.150 187.660 24.470 187.720 ;
        RECT 16.790 187.520 20.315 187.660 ;
        RECT 16.790 187.460 17.110 187.520 ;
        RECT 20.025 187.475 20.315 187.520 ;
        RECT 21.480 187.520 24.470 187.660 ;
        RECT 20.930 186.780 21.250 187.040 ;
        RECT 21.480 187.025 21.620 187.520 ;
        RECT 24.150 187.460 24.470 187.520 ;
        RECT 25.990 187.660 26.310 187.720 ;
        RECT 27.845 187.660 28.135 187.705 ;
        RECT 37.950 187.660 38.270 187.720 ;
        RECT 43.470 187.660 43.790 187.720 ;
        RECT 25.990 187.520 28.135 187.660 ;
        RECT 25.990 187.460 26.310 187.520 ;
        RECT 27.845 187.475 28.135 187.520 ;
        RECT 30.680 187.520 37.720 187.660 ;
        RECT 21.865 187.320 22.155 187.365 ;
        RECT 23.690 187.320 24.010 187.380 ;
        RECT 25.545 187.320 25.835 187.365 ;
        RECT 30.680 187.320 30.820 187.520 ;
        RECT 21.865 187.180 23.460 187.320 ;
        RECT 21.865 187.135 22.155 187.180 ;
        RECT 23.320 187.025 23.460 187.180 ;
        RECT 23.690 187.180 25.300 187.320 ;
        RECT 23.690 187.120 24.010 187.180 ;
        RECT 21.405 186.795 21.695 187.025 ;
        RECT 22.325 186.980 22.615 187.025 ;
        RECT 22.325 186.840 23.000 186.980 ;
        RECT 22.325 186.795 22.615 186.840 ;
        RECT 22.860 186.300 23.000 186.840 ;
        RECT 23.245 186.795 23.535 187.025 ;
        RECT 24.150 186.780 24.470 187.040 ;
        RECT 24.610 186.780 24.930 187.040 ;
        RECT 25.160 186.980 25.300 187.180 ;
        RECT 25.545 187.180 30.820 187.320 ;
        RECT 35.205 187.320 35.495 187.365 ;
        RECT 37.580 187.320 37.720 187.520 ;
        RECT 37.950 187.520 43.790 187.660 ;
        RECT 37.950 187.460 38.270 187.520 ;
        RECT 43.470 187.460 43.790 187.520 ;
        RECT 43.930 187.660 44.250 187.720 ;
        RECT 44.865 187.660 45.155 187.705 ;
        RECT 43.930 187.520 45.155 187.660 ;
        RECT 43.930 187.460 44.250 187.520 ;
        RECT 44.865 187.475 45.155 187.520 ;
        RECT 46.230 187.460 46.550 187.720 ;
        RECT 48.990 187.460 49.310 187.720 ;
        RECT 51.290 187.460 51.610 187.720 ;
        RECT 65.090 187.660 65.410 187.720 ;
        RECT 55.060 187.520 65.410 187.660 ;
        RECT 51.380 187.320 51.520 187.460 ;
        RECT 35.205 187.180 36.800 187.320 ;
        RECT 37.580 187.180 48.800 187.320 ;
        RECT 25.545 187.135 25.835 187.180 ;
        RECT 35.205 187.135 35.495 187.180 ;
        RECT 27.550 186.980 27.840 187.025 ;
        RECT 25.160 186.840 27.840 186.980 ;
        RECT 27.550 186.795 27.840 186.840 ;
        RECT 28.290 186.980 28.610 187.040 ;
        RECT 29.685 186.980 29.975 187.025 ;
        RECT 28.290 186.840 29.975 186.980 ;
        RECT 28.290 186.780 28.610 186.840 ;
        RECT 29.685 186.795 29.975 186.840 ;
        RECT 30.130 186.780 30.450 187.040 ;
        RECT 30.590 186.780 30.910 187.040 ;
        RECT 31.525 186.795 31.815 187.025 ;
        RECT 31.985 186.980 32.275 187.025 ;
        RECT 33.350 186.980 33.670 187.040 ;
        RECT 31.985 186.840 33.670 186.980 ;
        RECT 31.985 186.795 32.275 186.840 ;
        RECT 23.705 186.640 23.995 186.685 ;
        RECT 25.070 186.640 25.390 186.700 ;
        RECT 23.705 186.500 25.390 186.640 ;
        RECT 23.705 186.455 23.995 186.500 ;
        RECT 25.070 186.440 25.390 186.500 ;
        RECT 26.450 186.640 26.770 186.700 ;
        RECT 31.600 186.640 31.740 186.795 ;
        RECT 26.450 186.500 31.740 186.640 ;
        RECT 26.450 186.440 26.770 186.500 ;
        RECT 25.530 186.300 25.850 186.360 ;
        RECT 22.860 186.160 25.850 186.300 ;
        RECT 25.530 186.100 25.850 186.160 ;
        RECT 30.605 186.300 30.895 186.345 ;
        RECT 32.060 186.300 32.200 186.795 ;
        RECT 33.350 186.780 33.670 186.840 ;
        RECT 34.730 186.980 35.050 187.040 ;
        RECT 36.660 186.980 36.800 187.180 ;
        RECT 37.490 186.980 37.810 187.040 ;
        RECT 39.345 186.980 39.635 187.025 ;
        RECT 34.730 186.970 35.880 186.980 ;
        RECT 34.730 186.840 36.340 186.970 ;
        RECT 36.660 186.840 39.635 186.980 ;
        RECT 34.730 186.780 35.050 186.840 ;
        RECT 35.740 186.830 36.340 186.840 ;
        RECT 32.430 186.640 32.750 186.700 ;
        RECT 36.200 186.685 36.340 186.830 ;
        RECT 37.490 186.780 37.810 186.840 ;
        RECT 39.345 186.795 39.635 186.840 ;
        RECT 39.805 186.980 40.095 187.025 ;
        RECT 42.090 186.980 42.410 187.040 ;
        RECT 45.310 186.980 45.630 187.040 ;
        RECT 39.805 186.840 41.860 186.980 ;
        RECT 39.805 186.795 40.095 186.840 ;
        RECT 32.430 186.500 34.040 186.640 ;
        RECT 32.430 186.440 32.750 186.500 ;
        RECT 30.605 186.160 32.200 186.300 ;
        RECT 33.900 186.300 34.040 186.500 ;
        RECT 35.665 186.455 35.955 186.685 ;
        RECT 36.125 186.455 36.415 186.685 ;
        RECT 39.880 186.640 40.020 186.795 ;
        RECT 36.660 186.500 40.020 186.640 ;
        RECT 35.740 186.300 35.880 186.455 ;
        RECT 36.660 186.300 36.800 186.500 ;
        RECT 40.265 186.455 40.555 186.685 ;
        RECT 33.900 186.160 35.420 186.300 ;
        RECT 35.740 186.160 36.800 186.300 ;
        RECT 39.330 186.300 39.650 186.360 ;
        RECT 40.340 186.300 40.480 186.455 ;
        RECT 39.330 186.160 40.480 186.300 ;
        RECT 41.720 186.300 41.860 186.840 ;
        RECT 42.090 186.840 45.630 186.980 ;
        RECT 42.090 186.780 42.410 186.840 ;
        RECT 45.310 186.780 45.630 186.840 ;
        RECT 43.470 186.640 43.790 186.700 ;
        RECT 45.785 186.640 46.075 186.685 ;
        RECT 43.470 186.500 46.075 186.640 ;
        RECT 43.470 186.440 43.790 186.500 ;
        RECT 45.785 186.455 46.075 186.500 ;
        RECT 46.690 186.640 47.010 186.700 ;
        RECT 47.165 186.640 47.455 186.685 ;
        RECT 46.690 186.500 47.455 186.640 ;
        RECT 48.660 186.640 48.800 187.180 ;
        RECT 50.460 187.180 51.520 187.320 ;
        RECT 52.670 187.320 52.990 187.380 ;
        RECT 55.060 187.365 55.200 187.520 ;
        RECT 65.090 187.460 65.410 187.520 ;
        RECT 71.530 187.460 71.850 187.720 ;
        RECT 77.050 187.660 77.370 187.720 ;
        RECT 85.330 187.660 85.650 187.720 ;
        RECT 77.050 187.520 85.650 187.660 ;
        RECT 77.050 187.460 77.370 187.520 ;
        RECT 85.330 187.460 85.650 187.520 ;
        RECT 52.670 187.180 53.820 187.320 ;
        RECT 49.005 186.980 49.295 187.025 ;
        RECT 49.450 186.980 49.770 187.040 ;
        RECT 49.005 186.840 49.770 186.980 ;
        RECT 49.005 186.795 49.295 186.840 ;
        RECT 49.450 186.780 49.770 186.840 ;
        RECT 49.910 186.780 50.230 187.040 ;
        RECT 50.460 187.025 50.600 187.180 ;
        RECT 52.670 187.120 52.990 187.180 ;
        RECT 50.385 186.795 50.675 187.025 ;
        RECT 51.125 186.795 51.415 187.025 ;
        RECT 53.145 186.795 53.435 187.025 ;
        RECT 51.200 186.640 51.340 186.795 ;
        RECT 48.660 186.500 51.340 186.640 ;
        RECT 46.690 186.440 47.010 186.500 ;
        RECT 47.165 186.455 47.455 186.500 ;
        RECT 51.765 186.455 52.055 186.685 ;
        RECT 43.930 186.300 44.250 186.360 ;
        RECT 41.720 186.160 44.250 186.300 ;
        RECT 30.605 186.115 30.895 186.160 ;
        RECT 26.925 185.960 27.215 186.005 ;
        RECT 27.830 185.960 28.150 186.020 ;
        RECT 26.925 185.820 28.150 185.960 ;
        RECT 26.925 185.775 27.215 185.820 ;
        RECT 27.830 185.760 28.150 185.820 ;
        RECT 31.970 185.960 32.290 186.020 ;
        RECT 32.445 185.960 32.735 186.005 ;
        RECT 31.970 185.820 32.735 185.960 ;
        RECT 31.970 185.760 32.290 185.820 ;
        RECT 32.445 185.775 32.735 185.820 ;
        RECT 33.365 185.960 33.655 186.005 ;
        RECT 33.810 185.960 34.130 186.020 ;
        RECT 33.365 185.820 34.130 185.960 ;
        RECT 35.280 185.960 35.420 186.160 ;
        RECT 39.330 186.100 39.650 186.160 ;
        RECT 43.930 186.100 44.250 186.160 ;
        RECT 48.585 186.300 48.875 186.345 ;
        RECT 49.910 186.300 50.230 186.360 ;
        RECT 51.840 186.300 51.980 186.455 ;
        RECT 52.210 186.440 52.530 186.700 ;
        RECT 52.670 186.640 52.990 186.700 ;
        RECT 53.220 186.640 53.360 186.795 ;
        RECT 52.670 186.500 53.360 186.640 ;
        RECT 53.680 186.640 53.820 187.180 ;
        RECT 54.985 187.135 55.275 187.365 ;
        RECT 55.430 187.320 55.750 187.380 ;
        RECT 59.110 187.320 59.430 187.380 ;
        RECT 55.430 187.180 59.430 187.320 ;
        RECT 55.430 187.120 55.750 187.180 ;
        RECT 59.110 187.120 59.430 187.180 ;
        RECT 59.585 187.320 59.875 187.365 ;
        RECT 60.030 187.320 60.350 187.380 ;
        RECT 59.585 187.180 60.350 187.320 ;
        RECT 59.585 187.135 59.875 187.180 ;
        RECT 60.030 187.120 60.350 187.180 ;
        RECT 69.245 187.320 69.535 187.365 ;
        RECT 75.210 187.320 75.530 187.380 ;
        RECT 69.245 187.180 75.530 187.320 ;
        RECT 69.245 187.135 69.535 187.180 ;
        RECT 75.210 187.120 75.530 187.180 ;
        RECT 86.250 187.320 86.570 187.380 ;
        RECT 87.185 187.320 87.475 187.365 ;
        RECT 86.250 187.180 87.475 187.320 ;
        RECT 86.250 187.120 86.570 187.180 ;
        RECT 87.185 187.135 87.475 187.180 ;
        RECT 54.065 186.980 54.355 187.025 ;
        RECT 54.525 186.980 54.815 187.025 ;
        RECT 54.065 186.840 54.815 186.980 ;
        RECT 54.065 186.795 54.355 186.840 ;
        RECT 54.525 186.795 54.815 186.840 ;
        RECT 56.365 186.980 56.655 187.025 ;
        RECT 57.270 186.980 57.590 187.040 ;
        RECT 71.235 186.980 71.525 187.025 ;
        RECT 56.365 186.840 57.590 186.980 ;
        RECT 56.365 186.795 56.655 186.840 ;
        RECT 57.270 186.780 57.590 186.840 ;
        RECT 65.640 186.840 71.525 186.980 ;
        RECT 65.640 186.700 65.780 186.840 ;
        RECT 71.235 186.795 71.525 186.840 ;
        RECT 73.845 186.980 74.135 187.025 ;
        RECT 74.290 186.980 74.610 187.040 ;
        RECT 73.845 186.840 74.610 186.980 ;
        RECT 73.845 186.795 74.135 186.840 ;
        RECT 74.290 186.780 74.610 186.840 ;
        RECT 75.685 186.795 75.975 187.025 ;
        RECT 76.130 186.980 76.450 187.040 ;
        RECT 77.970 186.980 78.290 187.040 ;
        RECT 76.130 186.840 78.290 186.980 ;
        RECT 55.445 186.640 55.735 186.685 ;
        RECT 56.810 186.640 57.130 186.700 ;
        RECT 53.680 186.500 57.130 186.640 ;
        RECT 52.670 186.440 52.990 186.500 ;
        RECT 55.445 186.455 55.735 186.500 ;
        RECT 56.810 186.440 57.130 186.500 ;
        RECT 58.190 186.640 58.510 186.700 ;
        RECT 60.030 186.640 60.350 186.700 ;
        RECT 58.190 186.500 60.350 186.640 ;
        RECT 58.190 186.440 58.510 186.500 ;
        RECT 60.030 186.440 60.350 186.500 ;
        RECT 65.550 186.440 65.870 186.700 ;
        RECT 73.370 186.640 73.690 186.700 ;
        RECT 75.760 186.640 75.900 186.795 ;
        RECT 76.130 186.780 76.450 186.840 ;
        RECT 77.970 186.780 78.290 186.840 ;
        RECT 85.330 186.980 85.650 187.040 ;
        RECT 85.805 186.980 86.095 187.025 ;
        RECT 85.330 186.840 86.095 186.980 ;
        RECT 85.330 186.780 85.650 186.840 ;
        RECT 85.805 186.795 86.095 186.840 ;
        RECT 86.265 186.640 86.555 186.685 ;
        RECT 73.370 186.500 86.555 186.640 ;
        RECT 73.370 186.440 73.690 186.500 ;
        RECT 86.265 186.455 86.555 186.500 ;
        RECT 48.585 186.160 51.980 186.300 ;
        RECT 53.590 186.300 53.910 186.360 ;
        RECT 70.625 186.300 70.915 186.345 ;
        RECT 53.590 186.160 70.915 186.300 ;
        RECT 48.585 186.115 48.875 186.160 ;
        RECT 49.910 186.100 50.230 186.160 ;
        RECT 53.590 186.100 53.910 186.160 ;
        RECT 70.625 186.115 70.915 186.160 ;
        RECT 37.505 185.960 37.795 186.005 ;
        RECT 35.280 185.820 37.795 185.960 ;
        RECT 33.365 185.775 33.655 185.820 ;
        RECT 33.810 185.760 34.130 185.820 ;
        RECT 37.505 185.775 37.795 185.820 ;
        RECT 41.630 185.960 41.950 186.020 ;
        RECT 43.025 185.960 43.315 186.005 ;
        RECT 41.630 185.820 43.315 185.960 ;
        RECT 41.630 185.760 41.950 185.820 ;
        RECT 43.025 185.775 43.315 185.820 ;
        RECT 45.310 185.960 45.630 186.020 ;
        RECT 47.625 185.960 47.915 186.005 ;
        RECT 45.310 185.820 47.915 185.960 ;
        RECT 45.310 185.760 45.630 185.820 ;
        RECT 47.625 185.775 47.915 185.820 ;
        RECT 53.130 185.960 53.450 186.020 ;
        RECT 61.410 185.960 61.730 186.020 ;
        RECT 53.130 185.820 61.730 185.960 ;
        RECT 53.130 185.760 53.450 185.820 ;
        RECT 61.410 185.760 61.730 185.820 ;
        RECT 62.790 185.760 63.110 186.020 ;
        RECT 64.630 185.960 64.950 186.020 ;
        RECT 73.385 185.960 73.675 186.005 ;
        RECT 64.630 185.820 73.675 185.960 ;
        RECT 64.630 185.760 64.950 185.820 ;
        RECT 73.385 185.775 73.675 185.820 ;
        RECT 74.750 185.760 75.070 186.020 ;
        RECT 79.365 185.960 79.655 186.005 ;
        RECT 84.410 185.960 84.730 186.020 ;
        RECT 79.365 185.820 84.730 185.960 ;
        RECT 79.365 185.775 79.655 185.820 ;
        RECT 84.410 185.760 84.730 185.820 ;
        RECT 18.100 185.140 89.400 185.620 ;
        RECT 20.485 184.940 20.775 184.985 ;
        RECT 21.850 184.940 22.170 185.000 ;
        RECT 29.210 184.940 29.530 185.000 ;
        RECT 20.485 184.800 22.170 184.940 ;
        RECT 20.485 184.755 20.775 184.800 ;
        RECT 21.850 184.740 22.170 184.800 ;
        RECT 23.780 184.800 29.530 184.940 ;
        RECT 23.780 184.645 23.920 184.800 ;
        RECT 29.210 184.740 29.530 184.800 ;
        RECT 31.525 184.940 31.815 184.985 ;
        RECT 31.970 184.940 32.290 185.000 ;
        RECT 31.525 184.800 32.290 184.940 ;
        RECT 31.525 184.755 31.815 184.800 ;
        RECT 31.970 184.740 32.290 184.800 ;
        RECT 32.905 184.940 33.195 184.985 ;
        RECT 33.350 184.940 33.670 185.000 ;
        RECT 32.905 184.800 33.670 184.940 ;
        RECT 32.905 184.755 33.195 184.800 ;
        RECT 33.350 184.740 33.670 184.800 ;
        RECT 35.190 184.940 35.510 185.000 ;
        RECT 37.490 184.940 37.810 185.000 ;
        RECT 35.190 184.800 37.810 184.940 ;
        RECT 35.190 184.740 35.510 184.800 ;
        RECT 37.490 184.740 37.810 184.800 ;
        RECT 37.950 184.740 38.270 185.000 ;
        RECT 38.885 184.940 39.175 184.985 ;
        RECT 40.250 184.940 40.570 185.000 ;
        RECT 38.885 184.800 40.570 184.940 ;
        RECT 38.885 184.755 39.175 184.800 ;
        RECT 40.250 184.740 40.570 184.800 ;
        RECT 43.470 184.740 43.790 185.000 ;
        RECT 49.465 184.940 49.755 184.985 ;
        RECT 50.370 184.940 50.690 185.000 ;
        RECT 45.860 184.800 49.220 184.940 ;
        RECT 23.705 184.415 23.995 184.645 ;
        RECT 24.150 184.400 24.470 184.660 ;
        RECT 26.465 184.600 26.755 184.645 ;
        RECT 27.370 184.600 27.690 184.660 ;
        RECT 26.465 184.460 27.690 184.600 ;
        RECT 26.465 184.415 26.755 184.460 ;
        RECT 27.370 184.400 27.690 184.460 ;
        RECT 27.830 184.600 28.150 184.660 ;
        RECT 31.050 184.600 31.370 184.660 ;
        RECT 27.830 184.460 30.820 184.600 ;
        RECT 27.830 184.400 28.150 184.460 ;
        RECT 21.865 184.260 22.155 184.305 ;
        RECT 21.865 184.120 23.460 184.260 ;
        RECT 21.865 184.075 22.155 184.120 ;
        RECT 19.550 183.720 19.870 183.980 ;
        RECT 21.405 183.735 21.695 183.965 ;
        RECT 22.325 183.920 22.615 183.965 ;
        RECT 22.770 183.920 23.090 183.980 ;
        RECT 23.320 183.965 23.460 184.120 ;
        RECT 25.530 184.060 25.850 184.320 ;
        RECT 28.290 184.260 28.610 184.320 ;
        RECT 29.685 184.260 29.975 184.305 ;
        RECT 28.290 184.120 29.975 184.260 ;
        RECT 30.680 184.260 30.820 184.460 ;
        RECT 31.050 184.460 40.020 184.600 ;
        RECT 31.050 184.400 31.370 184.460 ;
        RECT 36.125 184.260 36.415 184.305 ;
        RECT 39.330 184.260 39.650 184.320 ;
        RECT 30.680 184.120 35.880 184.260 ;
        RECT 28.290 184.060 28.610 184.120 ;
        RECT 29.685 184.075 29.975 184.120 ;
        RECT 22.325 183.780 23.090 183.920 ;
        RECT 22.325 183.735 22.615 183.780 ;
        RECT 21.480 183.580 21.620 183.735 ;
        RECT 22.770 183.720 23.090 183.780 ;
        RECT 23.245 183.735 23.535 183.965 ;
        RECT 24.610 183.720 24.930 183.980 ;
        RECT 25.620 183.920 25.760 184.060 ;
        RECT 27.090 183.920 27.380 183.965 ;
        RECT 25.620 183.780 27.380 183.920 ;
        RECT 27.090 183.735 27.380 183.780 ;
        RECT 29.225 183.920 29.515 183.965 ;
        RECT 31.970 183.920 32.290 183.980 ;
        RECT 29.225 183.780 32.290 183.920 ;
        RECT 29.225 183.735 29.515 183.780 ;
        RECT 31.970 183.720 32.290 183.780 ;
        RECT 32.445 183.920 32.735 183.965 ;
        RECT 34.270 183.920 34.590 183.980 ;
        RECT 32.445 183.780 34.590 183.920 ;
        RECT 35.740 183.920 35.880 184.120 ;
        RECT 36.125 184.120 39.650 184.260 ;
        RECT 36.125 184.075 36.415 184.120 ;
        RECT 39.330 184.060 39.650 184.120 ;
        RECT 39.880 184.045 40.020 184.460 ;
        RECT 44.390 184.400 44.710 184.660 ;
        RECT 37.045 183.920 37.335 183.965 ;
        RECT 37.950 183.920 38.270 183.980 ;
        RECT 35.740 183.780 36.870 183.920 ;
        RECT 32.445 183.735 32.735 183.780 ;
        RECT 34.270 183.720 34.590 183.780 ;
        RECT 24.150 183.580 24.470 183.640 ;
        RECT 21.480 183.440 24.470 183.580 ;
        RECT 24.150 183.380 24.470 183.440 ;
        RECT 25.545 183.580 25.835 183.625 ;
        RECT 34.745 183.580 35.035 183.625 ;
        RECT 35.650 183.580 35.970 183.640 ;
        RECT 25.545 183.440 30.360 183.580 ;
        RECT 25.545 183.395 25.835 183.440 ;
        RECT 25.990 183.240 26.310 183.300 ;
        RECT 27.385 183.240 27.675 183.285 ;
        RECT 25.990 183.100 27.675 183.240 ;
        RECT 25.990 183.040 26.310 183.100 ;
        RECT 27.385 183.055 27.675 183.100 ;
        RECT 28.290 183.240 28.610 183.300 ;
        RECT 29.670 183.240 29.990 183.300 ;
        RECT 28.290 183.100 29.990 183.240 ;
        RECT 30.220 183.240 30.360 183.440 ;
        RECT 34.745 183.440 35.970 183.580 ;
        RECT 36.730 183.580 36.870 183.780 ;
        RECT 37.045 183.780 38.270 183.920 ;
        RECT 39.805 183.815 40.095 184.045 ;
        RECT 37.045 183.735 37.335 183.780 ;
        RECT 37.950 183.720 38.270 183.780 ;
        RECT 41.170 183.720 41.490 183.980 ;
        RECT 41.630 183.720 41.950 183.980 ;
        RECT 42.565 183.920 42.855 183.965 ;
        RECT 43.010 183.920 43.330 183.980 ;
        RECT 42.565 183.780 43.330 183.920 ;
        RECT 42.565 183.735 42.855 183.780 ;
        RECT 43.010 183.720 43.330 183.780 ;
        RECT 45.325 183.920 45.615 183.965 ;
        RECT 45.860 183.920 46.000 184.800 ;
        RECT 46.230 184.600 46.550 184.660 ;
        RECT 49.080 184.600 49.220 184.800 ;
        RECT 49.465 184.800 50.690 184.940 ;
        RECT 49.465 184.755 49.755 184.800 ;
        RECT 50.370 184.740 50.690 184.800 ;
        RECT 54.065 184.940 54.355 184.985 ;
        RECT 54.970 184.940 55.290 185.000 ;
        RECT 54.065 184.800 55.290 184.940 ;
        RECT 54.065 184.755 54.355 184.800 ;
        RECT 54.970 184.740 55.290 184.800 ;
        RECT 55.905 184.940 56.195 184.985 ;
        RECT 56.810 184.940 57.130 185.000 ;
        RECT 65.550 184.940 65.870 185.000 ;
        RECT 55.905 184.800 65.870 184.940 ;
        RECT 55.905 184.755 56.195 184.800 ;
        RECT 56.810 184.740 57.130 184.800 ;
        RECT 65.550 184.740 65.870 184.800 ;
        RECT 67.390 184.940 67.710 185.000 ;
        RECT 72.910 184.940 73.230 185.000 ;
        RECT 67.390 184.800 69.920 184.940 ;
        RECT 67.390 184.740 67.710 184.800 ;
        RECT 49.910 184.600 50.230 184.660 ;
        RECT 52.670 184.600 52.990 184.660 ;
        RECT 59.570 184.600 59.890 184.660 ;
        RECT 69.780 184.600 69.920 184.800 ;
        RECT 72.910 184.800 80.500 184.940 ;
        RECT 72.910 184.740 73.230 184.800 ;
        RECT 75.210 184.600 75.530 184.660 ;
        RECT 79.810 184.600 80.130 184.660 ;
        RECT 46.230 184.460 48.300 184.600 ;
        RECT 49.080 184.460 50.230 184.600 ;
        RECT 46.230 184.400 46.550 184.460 ;
        RECT 47.610 183.965 47.930 183.990 ;
        RECT 48.160 183.965 48.300 184.460 ;
        RECT 49.910 184.400 50.230 184.460 ;
        RECT 51.365 184.460 52.990 184.600 ;
        RECT 51.365 184.260 51.505 184.460 ;
        RECT 52.670 184.400 52.990 184.460 ;
        RECT 54.140 184.460 59.340 184.600 ;
        RECT 49.540 184.120 51.505 184.260 ;
        RECT 45.325 183.780 46.000 183.920 ;
        RECT 45.325 183.735 45.615 183.780 ;
        RECT 46.245 183.735 46.535 183.965 ;
        RECT 46.705 183.735 46.995 183.965 ;
        RECT 47.345 183.735 47.930 183.965 ;
        RECT 48.085 183.735 48.375 183.965 ;
        RECT 46.320 183.580 46.460 183.735 ;
        RECT 36.730 183.440 46.460 183.580 ;
        RECT 46.780 183.580 46.920 183.735 ;
        RECT 47.610 183.730 47.930 183.735 ;
        RECT 49.540 183.580 49.680 184.120 ;
        RECT 50.370 183.720 50.690 183.980 ;
        RECT 50.845 183.735 51.135 183.965 ;
        RECT 51.365 183.920 51.505 184.120 ;
        RECT 51.750 184.060 52.070 184.320 ;
        RECT 52.225 183.920 52.515 183.965 ;
        RECT 51.365 183.780 52.515 183.920 ;
        RECT 52.225 183.735 52.515 183.780 ;
        RECT 46.780 183.440 49.680 183.580 ;
        RECT 49.910 183.580 50.230 183.640 ;
        RECT 50.920 183.580 51.060 183.735 ;
        RECT 52.670 183.720 52.990 183.980 ;
        RECT 53.130 183.720 53.450 183.980 ;
        RECT 54.140 183.965 54.280 184.460 ;
        RECT 54.510 184.260 54.830 184.320 ;
        RECT 59.200 184.260 59.340 184.460 ;
        RECT 59.570 184.460 69.460 184.600 ;
        RECT 69.780 184.460 80.130 184.600 ;
        RECT 59.570 184.400 59.890 184.460 ;
        RECT 66.010 184.260 66.330 184.320 ;
        RECT 54.510 184.120 55.200 184.260 ;
        RECT 59.200 184.120 66.330 184.260 ;
        RECT 54.510 184.060 54.830 184.120 ;
        RECT 55.060 183.965 55.200 184.120 ;
        RECT 66.010 184.060 66.330 184.120 ;
        RECT 54.065 183.735 54.355 183.965 ;
        RECT 54.985 183.735 55.275 183.965 ;
        RECT 56.365 183.920 56.655 183.965 ;
        RECT 60.950 183.920 61.270 183.980 ;
        RECT 56.365 183.780 61.270 183.920 ;
        RECT 56.365 183.735 56.655 183.780 ;
        RECT 60.950 183.720 61.270 183.780 ;
        RECT 67.850 183.920 68.170 183.980 ;
        RECT 69.320 183.965 69.460 184.460 ;
        RECT 75.210 184.400 75.530 184.460 ;
        RECT 79.810 184.400 80.130 184.460 ;
        RECT 77.510 184.260 77.830 184.320 ;
        RECT 80.360 184.260 80.500 184.800 ;
        RECT 85.330 184.740 85.650 185.000 ;
        RECT 77.510 184.120 79.580 184.260 ;
        RECT 80.360 184.120 86.480 184.260 ;
        RECT 77.510 184.060 77.830 184.120 ;
        RECT 68.325 183.920 68.615 183.965 ;
        RECT 67.850 183.780 68.615 183.920 ;
        RECT 67.850 183.720 68.170 183.780 ;
        RECT 68.325 183.735 68.615 183.780 ;
        RECT 69.245 183.735 69.535 183.965 ;
        RECT 74.750 183.920 75.070 183.980 ;
        RECT 79.440 183.965 79.580 184.120 ;
        RECT 74.610 183.720 75.070 183.920 ;
        RECT 78.445 183.735 78.735 183.965 ;
        RECT 79.365 183.735 79.655 183.965 ;
        RECT 66.025 183.580 66.315 183.625 ;
        RECT 74.610 183.580 74.750 183.720 ;
        RECT 49.910 183.440 65.780 183.580 ;
        RECT 34.745 183.395 35.035 183.440 ;
        RECT 35.650 183.380 35.970 183.440 ;
        RECT 32.430 183.240 32.750 183.300 ;
        RECT 30.220 183.100 32.750 183.240 ;
        RECT 28.290 183.040 28.610 183.100 ;
        RECT 29.670 183.040 29.990 183.100 ;
        RECT 32.430 183.040 32.750 183.100 ;
        RECT 35.205 183.240 35.495 183.285 ;
        RECT 36.570 183.240 36.890 183.300 ;
        RECT 35.205 183.100 36.890 183.240 ;
        RECT 35.205 183.055 35.495 183.100 ;
        RECT 36.570 183.040 36.890 183.100 ;
        RECT 37.030 183.240 37.350 183.300 ;
        RECT 39.790 183.240 40.110 183.300 ;
        RECT 37.030 183.100 40.110 183.240 ;
        RECT 37.030 183.040 37.350 183.100 ;
        RECT 39.790 183.040 40.110 183.100 ;
        RECT 43.930 183.240 44.250 183.300 ;
        RECT 46.780 183.240 46.920 183.440 ;
        RECT 49.910 183.380 50.230 183.440 ;
        RECT 43.930 183.100 46.920 183.240 ;
        RECT 53.590 183.240 53.910 183.300 ;
        RECT 55.890 183.240 56.210 183.300 ;
        RECT 53.590 183.100 56.210 183.240 ;
        RECT 43.930 183.040 44.250 183.100 ;
        RECT 53.590 183.040 53.910 183.100 ;
        RECT 55.890 183.040 56.210 183.100 ;
        RECT 59.110 183.240 59.430 183.300 ;
        RECT 64.170 183.240 64.490 183.300 ;
        RECT 59.110 183.100 64.490 183.240 ;
        RECT 65.640 183.240 65.780 183.440 ;
        RECT 66.025 183.440 74.750 183.580 ;
        RECT 78.520 183.580 78.660 183.735 ;
        RECT 79.810 183.720 80.130 183.980 ;
        RECT 80.270 183.720 80.590 183.980 ;
        RECT 83.030 183.920 83.350 183.980 ;
        RECT 86.340 183.965 86.480 184.120 ;
        RECT 83.505 183.920 83.795 183.965 ;
        RECT 83.030 183.780 83.795 183.920 ;
        RECT 83.030 183.720 83.350 183.780 ;
        RECT 83.505 183.735 83.795 183.780 ;
        RECT 85.805 183.735 86.095 183.965 ;
        RECT 86.265 183.735 86.555 183.965 ;
        RECT 81.665 183.580 81.955 183.625 ;
        RECT 85.330 183.580 85.650 183.640 ;
        RECT 78.520 183.440 80.500 183.580 ;
        RECT 66.025 183.395 66.315 183.440 ;
        RECT 80.360 183.300 80.500 183.440 ;
        RECT 81.665 183.440 85.650 183.580 ;
        RECT 85.880 183.580 86.020 183.735 ;
        RECT 87.170 183.720 87.490 183.980 ;
        RECT 88.550 183.580 88.870 183.640 ;
        RECT 89.470 183.580 89.790 183.640 ;
        RECT 85.880 183.440 89.790 183.580 ;
        RECT 81.665 183.395 81.955 183.440 ;
        RECT 85.330 183.380 85.650 183.440 ;
        RECT 88.550 183.380 88.870 183.440 ;
        RECT 89.470 183.380 89.790 183.440 ;
        RECT 70.610 183.240 70.930 183.300 ;
        RECT 65.640 183.100 70.930 183.240 ;
        RECT 59.110 183.040 59.430 183.100 ;
        RECT 64.170 183.040 64.490 183.100 ;
        RECT 70.610 183.040 70.930 183.100 ;
        RECT 76.130 183.240 76.450 183.300 ;
        RECT 76.605 183.240 76.895 183.285 ;
        RECT 76.130 183.100 76.895 183.240 ;
        RECT 76.130 183.040 76.450 183.100 ;
        RECT 76.605 183.055 76.895 183.100 ;
        RECT 80.270 183.040 80.590 183.300 ;
        RECT 81.190 183.240 81.510 183.300 ;
        RECT 83.950 183.240 84.270 183.300 ;
        RECT 86.725 183.240 87.015 183.285 ;
        RECT 81.190 183.100 87.015 183.240 ;
        RECT 81.190 183.040 81.510 183.100 ;
        RECT 83.950 183.040 84.270 183.100 ;
        RECT 86.725 183.055 87.015 183.100 ;
        RECT 18.100 182.420 89.400 182.900 ;
        RECT 18.630 182.220 18.950 182.280 ;
        RECT 21.865 182.220 22.155 182.265 ;
        RECT 18.630 182.080 22.155 182.220 ;
        RECT 18.630 182.020 18.950 182.080 ;
        RECT 21.865 182.035 22.155 182.080 ;
        RECT 24.610 182.220 24.930 182.280 ;
        RECT 25.545 182.220 25.835 182.265 ;
        RECT 24.610 182.080 25.835 182.220 ;
        RECT 24.610 182.020 24.930 182.080 ;
        RECT 25.545 182.035 25.835 182.080 ;
        RECT 26.465 182.220 26.755 182.265 ;
        RECT 27.830 182.220 28.150 182.280 ;
        RECT 26.465 182.080 28.150 182.220 ;
        RECT 26.465 182.035 26.755 182.080 ;
        RECT 27.830 182.020 28.150 182.080 ;
        RECT 28.765 182.035 29.055 182.265 ;
        RECT 20.930 181.880 21.250 181.940 ;
        RECT 23.705 181.880 23.995 181.925 ;
        RECT 20.930 181.740 23.995 181.880 ;
        RECT 28.840 181.880 28.980 182.035 ;
        RECT 30.130 182.020 30.450 182.280 ;
        RECT 30.590 182.220 30.910 182.280 ;
        RECT 31.065 182.220 31.355 182.265 ;
        RECT 30.590 182.080 31.355 182.220 ;
        RECT 30.590 182.020 30.910 182.080 ;
        RECT 31.065 182.035 31.355 182.080 ;
        RECT 35.190 182.020 35.510 182.280 ;
        RECT 36.110 182.220 36.430 182.280 ;
        RECT 37.030 182.220 37.350 182.280 ;
        RECT 36.110 182.080 37.350 182.220 ;
        RECT 36.110 182.020 36.430 182.080 ;
        RECT 37.030 182.020 37.350 182.080 ;
        RECT 41.170 182.220 41.490 182.280 ;
        RECT 44.405 182.220 44.695 182.265 ;
        RECT 41.170 182.080 44.695 182.220 ;
        RECT 41.170 182.020 41.490 182.080 ;
        RECT 44.405 182.035 44.695 182.080 ;
        RECT 47.150 182.020 47.470 182.280 ;
        RECT 48.070 182.220 48.390 182.280 ;
        RECT 48.545 182.220 48.835 182.265 ;
        RECT 48.070 182.080 48.835 182.220 ;
        RECT 48.070 182.020 48.390 182.080 ;
        RECT 48.545 182.035 48.835 182.080 ;
        RECT 50.845 182.220 51.135 182.265 ;
        RECT 54.050 182.220 54.370 182.280 ;
        RECT 50.845 182.080 54.370 182.220 ;
        RECT 50.845 182.035 51.135 182.080 ;
        RECT 54.050 182.020 54.370 182.080 ;
        RECT 60.030 182.220 60.350 182.280 ;
        RECT 60.950 182.220 61.270 182.280 ;
        RECT 60.030 182.080 61.270 182.220 ;
        RECT 60.030 182.020 60.350 182.080 ;
        RECT 60.950 182.020 61.270 182.080 ;
        RECT 61.410 182.020 61.730 182.280 ;
        RECT 62.330 182.220 62.650 182.280 ;
        RECT 63.710 182.220 64.030 182.280 ;
        RECT 65.565 182.220 65.855 182.265 ;
        RECT 62.330 182.080 63.020 182.220 ;
        RECT 62.330 182.020 62.650 182.080 ;
        RECT 31.510 181.880 31.830 181.940 ;
        RECT 28.840 181.740 31.830 181.880 ;
        RECT 20.930 181.680 21.250 181.740 ;
        RECT 23.705 181.695 23.995 181.740 ;
        RECT 31.510 181.680 31.830 181.740 ;
        RECT 33.810 181.880 34.130 181.940 ;
        RECT 45.310 181.880 45.630 181.940 ;
        RECT 54.985 181.880 55.275 181.925 ;
        RECT 56.810 181.880 57.130 181.940 ;
        RECT 61.500 181.880 61.640 182.020 ;
        RECT 62.880 181.925 63.020 182.080 ;
        RECT 63.710 182.080 65.855 182.220 ;
        RECT 63.710 182.020 64.030 182.080 ;
        RECT 65.565 182.035 65.855 182.080 ;
        RECT 68.310 182.220 68.630 182.280 ;
        RECT 68.785 182.220 69.075 182.265 ;
        RECT 68.310 182.080 69.075 182.220 ;
        RECT 68.310 182.020 68.630 182.080 ;
        RECT 68.785 182.035 69.075 182.080 ;
        RECT 73.830 182.220 74.150 182.280 ;
        RECT 78.445 182.220 78.735 182.265 ;
        RECT 87.170 182.220 87.490 182.280 ;
        RECT 73.830 182.080 87.490 182.220 ;
        RECT 73.830 182.020 74.150 182.080 ;
        RECT 78.445 182.035 78.735 182.080 ;
        RECT 87.170 182.020 87.490 182.080 ;
        RECT 33.810 181.740 45.630 181.880 ;
        RECT 33.810 181.680 34.130 181.740 ;
        RECT 45.310 181.680 45.630 181.740 ;
        RECT 46.320 181.740 54.280 181.880 ;
        RECT 18.170 181.540 18.490 181.600 ;
        RECT 21.405 181.540 21.695 181.585 ;
        RECT 18.170 181.400 21.695 181.540 ;
        RECT 18.170 181.340 18.490 181.400 ;
        RECT 21.405 181.355 21.695 181.400 ;
        RECT 22.770 181.340 23.090 181.600 ;
        RECT 25.070 181.340 25.390 181.600 ;
        RECT 25.990 181.340 26.310 181.600 ;
        RECT 26.910 181.540 27.230 181.600 ;
        RECT 27.385 181.540 27.675 181.585 ;
        RECT 26.910 181.400 27.675 181.540 ;
        RECT 26.910 181.340 27.230 181.400 ;
        RECT 27.385 181.355 27.675 181.400 ;
        RECT 27.830 181.340 28.150 181.600 ;
        RECT 29.210 181.340 29.530 181.600 ;
        RECT 30.605 181.355 30.895 181.585 ;
        RECT 21.850 181.200 22.170 181.260 ;
        RECT 30.680 181.200 30.820 181.355 ;
        RECT 32.890 181.340 33.210 181.600 ;
        RECT 34.285 181.355 34.575 181.585 ;
        RECT 35.205 181.540 35.495 181.585 ;
        RECT 40.710 181.540 41.030 181.600 ;
        RECT 35.205 181.400 41.030 181.540 ;
        RECT 35.205 181.355 35.495 181.400 ;
        RECT 21.850 181.060 30.820 181.200 ;
        RECT 34.360 181.200 34.500 181.355 ;
        RECT 40.710 181.340 41.030 181.400 ;
        RECT 43.930 181.540 44.250 181.600 ;
        RECT 46.320 181.540 46.460 181.740 ;
        RECT 54.140 181.600 54.280 181.740 ;
        RECT 54.985 181.740 58.420 181.880 ;
        RECT 54.985 181.695 55.275 181.740 ;
        RECT 56.810 181.680 57.130 181.740 ;
        RECT 43.930 181.400 46.460 181.540 ;
        RECT 43.930 181.340 44.250 181.400 ;
        RECT 46.690 181.340 47.010 181.600 ;
        RECT 48.085 181.540 48.375 181.585 ;
        RECT 48.530 181.540 48.850 181.600 ;
        RECT 48.085 181.400 48.850 181.540 ;
        RECT 48.085 181.355 48.375 181.400 ;
        RECT 48.530 181.340 48.850 181.400 ;
        RECT 49.450 181.340 49.770 181.600 ;
        RECT 49.925 181.355 50.215 181.585 ;
        RECT 52.225 181.540 52.515 181.585 ;
        RECT 53.130 181.540 53.450 181.600 ;
        RECT 52.225 181.400 53.450 181.540 ;
        RECT 52.225 181.355 52.515 181.400 ;
        RECT 36.110 181.200 36.430 181.260 ;
        RECT 44.865 181.200 45.155 181.245 ;
        RECT 34.360 181.060 45.155 181.200 ;
        RECT 21.850 181.000 22.170 181.060 ;
        RECT 36.110 181.000 36.430 181.060 ;
        RECT 44.865 181.015 45.155 181.060 ;
        RECT 45.325 181.015 45.615 181.245 ;
        RECT 50.000 181.200 50.140 181.355 ;
        RECT 53.130 181.340 53.450 181.400 ;
        RECT 53.590 181.340 53.910 181.600 ;
        RECT 54.050 181.340 54.370 181.600 ;
        RECT 54.510 181.540 54.830 181.600 ;
        RECT 55.445 181.540 55.735 181.585 ;
        RECT 54.510 181.400 55.735 181.540 ;
        RECT 54.510 181.340 54.830 181.400 ;
        RECT 55.445 181.355 55.735 181.400 ;
        RECT 55.890 181.340 56.210 181.600 ;
        RECT 58.280 181.585 58.420 181.740 ;
        RECT 58.740 181.740 61.640 181.880 ;
        RECT 58.205 181.355 58.495 181.585 ;
        RECT 52.670 181.200 52.990 181.260 ;
        RECT 57.285 181.200 57.575 181.245 ;
        RECT 50.000 181.060 52.440 181.200 ;
        RECT 19.090 180.860 19.410 180.920 ;
        RECT 31.985 180.860 32.275 180.905 ;
        RECT 19.090 180.720 32.275 180.860 ;
        RECT 19.090 180.660 19.410 180.720 ;
        RECT 31.985 180.675 32.275 180.720 ;
        RECT 32.430 180.860 32.750 180.920 ;
        RECT 43.930 180.860 44.250 180.920 ;
        RECT 45.400 180.860 45.540 181.015 ;
        RECT 32.430 180.720 44.250 180.860 ;
        RECT 32.430 180.660 32.750 180.720 ;
        RECT 43.930 180.660 44.250 180.720 ;
        RECT 44.480 180.720 45.540 180.860 ;
        RECT 45.770 180.860 46.090 180.920 ;
        RECT 51.305 180.860 51.595 180.905 ;
        RECT 45.770 180.720 51.595 180.860 ;
        RECT 52.300 180.860 52.440 181.060 ;
        RECT 52.670 181.060 57.575 181.200 ;
        RECT 52.670 181.000 52.990 181.060 ;
        RECT 57.285 181.015 57.575 181.060 ;
        RECT 58.740 180.860 58.880 181.740 ;
        RECT 62.805 181.695 63.095 181.925 ;
        RECT 74.750 181.880 75.070 181.940 ;
        RECT 84.410 181.880 84.730 181.940 ;
        RECT 87.645 181.880 87.935 181.925 ;
        RECT 74.750 181.740 76.820 181.880 ;
        RECT 74.750 181.680 75.070 181.740 ;
        RECT 60.045 181.355 60.335 181.585 ;
        RECT 60.965 181.540 61.255 181.585 ;
        RECT 61.410 181.540 61.730 181.600 ;
        RECT 60.965 181.400 61.730 181.540 ;
        RECT 60.965 181.355 61.255 181.400 ;
        RECT 59.125 181.015 59.415 181.245 ;
        RECT 52.300 180.720 58.880 180.860 ;
        RECT 59.200 180.860 59.340 181.015 ;
        RECT 59.570 181.000 59.890 181.260 ;
        RECT 60.120 181.200 60.260 181.355 ;
        RECT 61.410 181.340 61.730 181.400 ;
        RECT 62.345 181.355 62.635 181.585 ;
        RECT 63.265 181.540 63.555 181.585 ;
        RECT 63.710 181.540 64.030 181.600 ;
        RECT 63.265 181.400 64.030 181.540 ;
        RECT 63.265 181.355 63.555 181.400 ;
        RECT 61.870 181.200 62.190 181.260 ;
        RECT 60.120 181.060 62.190 181.200 ;
        RECT 62.420 181.200 62.560 181.355 ;
        RECT 63.710 181.340 64.030 181.400 ;
        RECT 64.185 181.540 64.475 181.585 ;
        RECT 64.630 181.540 64.950 181.600 ;
        RECT 64.185 181.400 64.950 181.540 ;
        RECT 64.185 181.355 64.475 181.400 ;
        RECT 64.630 181.340 64.950 181.400 ;
        RECT 65.550 181.540 65.870 181.600 ;
        RECT 66.945 181.540 67.235 181.585 ;
        RECT 65.550 181.400 67.235 181.540 ;
        RECT 65.550 181.340 65.870 181.400 ;
        RECT 66.945 181.355 67.235 181.400 ;
        RECT 76.130 181.340 76.450 181.600 ;
        RECT 76.680 181.585 76.820 181.740 ;
        RECT 84.410 181.740 87.935 181.880 ;
        RECT 84.410 181.680 84.730 181.740 ;
        RECT 87.645 181.695 87.935 181.740 ;
        RECT 76.605 181.355 76.895 181.585 ;
        RECT 77.050 181.340 77.370 181.600 ;
        RECT 62.420 181.060 65.320 181.200 ;
        RECT 61.870 181.000 62.190 181.060 ;
        RECT 61.960 180.860 62.100 181.000 ;
        RECT 65.180 180.920 65.320 181.060 ;
        RECT 66.485 181.015 66.775 181.245 ;
        RECT 76.220 181.200 76.360 181.340 ;
        RECT 86.250 181.200 86.570 181.260 ;
        RECT 76.220 181.060 86.570 181.200 ;
        RECT 64.630 180.860 64.950 180.920 ;
        RECT 59.200 180.720 60.400 180.860 ;
        RECT 61.960 180.720 64.950 180.860 ;
        RECT 44.480 180.580 44.620 180.720 ;
        RECT 45.770 180.660 46.090 180.720 ;
        RECT 51.305 180.675 51.595 180.720 ;
        RECT 20.470 180.320 20.790 180.580 ;
        RECT 24.165 180.520 24.455 180.565 ;
        RECT 25.070 180.520 25.390 180.580 ;
        RECT 26.450 180.520 26.770 180.580 ;
        RECT 24.165 180.380 26.770 180.520 ;
        RECT 24.165 180.335 24.455 180.380 ;
        RECT 25.070 180.320 25.390 180.380 ;
        RECT 26.450 180.320 26.770 180.380 ;
        RECT 29.210 180.520 29.530 180.580 ;
        RECT 44.390 180.520 44.710 180.580 ;
        RECT 29.210 180.380 44.710 180.520 ;
        RECT 29.210 180.320 29.530 180.380 ;
        RECT 44.390 180.320 44.710 180.380 ;
        RECT 44.850 180.520 45.170 180.580 ;
        RECT 46.245 180.520 46.535 180.565 ;
        RECT 44.850 180.380 46.535 180.520 ;
        RECT 44.850 180.320 45.170 180.380 ;
        RECT 46.245 180.335 46.535 180.380 ;
        RECT 50.370 180.520 50.690 180.580 ;
        RECT 52.670 180.520 52.990 180.580 ;
        RECT 50.370 180.380 52.990 180.520 ;
        RECT 50.370 180.320 50.690 180.380 ;
        RECT 52.670 180.320 52.990 180.380 ;
        RECT 55.890 180.520 56.210 180.580 ;
        RECT 56.825 180.520 57.115 180.565 ;
        RECT 55.890 180.380 57.115 180.520 ;
        RECT 60.260 180.520 60.400 180.720 ;
        RECT 64.630 180.660 64.950 180.720 ;
        RECT 65.090 180.660 65.410 180.920 ;
        RECT 66.560 180.860 66.700 181.015 ;
        RECT 86.250 181.000 86.570 181.060 ;
        RECT 69.230 180.860 69.550 180.920 ;
        RECT 81.190 180.860 81.510 180.920 ;
        RECT 66.560 180.720 69.550 180.860 ;
        RECT 69.230 180.660 69.550 180.720 ;
        RECT 74.610 180.720 81.510 180.860 ;
        RECT 60.950 180.520 61.270 180.580 ;
        RECT 60.260 180.380 61.270 180.520 ;
        RECT 55.890 180.320 56.210 180.380 ;
        RECT 56.825 180.335 57.115 180.380 ;
        RECT 60.950 180.320 61.270 180.380 ;
        RECT 61.425 180.520 61.715 180.565 ;
        RECT 61.870 180.520 62.190 180.580 ;
        RECT 61.425 180.380 62.190 180.520 ;
        RECT 61.425 180.335 61.715 180.380 ;
        RECT 61.870 180.320 62.190 180.380 ;
        RECT 66.930 180.520 67.250 180.580 ;
        RECT 74.610 180.520 74.750 180.720 ;
        RECT 81.190 180.660 81.510 180.720 ;
        RECT 66.930 180.380 74.750 180.520 ;
        RECT 66.930 180.320 67.250 180.380 ;
        RECT 80.270 180.320 80.590 180.580 ;
        RECT 18.100 179.700 89.400 180.180 ;
        RECT 23.230 179.300 23.550 179.560 ;
        RECT 26.910 179.500 27.230 179.560 ;
        RECT 29.210 179.500 29.530 179.560 ;
        RECT 26.910 179.360 29.530 179.500 ;
        RECT 26.910 179.300 27.230 179.360 ;
        RECT 29.210 179.300 29.530 179.360 ;
        RECT 30.605 179.500 30.895 179.545 ;
        RECT 32.890 179.500 33.210 179.560 ;
        RECT 41.185 179.500 41.475 179.545 ;
        RECT 30.605 179.360 33.210 179.500 ;
        RECT 30.605 179.315 30.895 179.360 ;
        RECT 32.890 179.300 33.210 179.360 ;
        RECT 34.820 179.360 41.475 179.500 ;
        RECT 24.165 179.160 24.455 179.205 ;
        RECT 26.450 179.160 26.770 179.220 ;
        RECT 27.370 179.160 27.690 179.220 ;
        RECT 24.165 179.020 25.340 179.160 ;
        RECT 24.165 178.975 24.455 179.020 ;
        RECT 21.405 178.480 21.695 178.525 ;
        RECT 22.310 178.480 22.630 178.540 ;
        RECT 21.405 178.340 22.630 178.480 ;
        RECT 25.200 178.480 25.340 179.020 ;
        RECT 26.310 179.020 27.690 179.160 ;
        RECT 26.310 178.960 26.770 179.020 ;
        RECT 27.370 178.960 27.690 179.020 ;
        RECT 28.290 178.960 28.610 179.220 ;
        RECT 25.545 178.820 25.835 178.865 ;
        RECT 26.310 178.820 26.450 178.960 ;
        RECT 25.545 178.680 26.450 178.820 ;
        RECT 26.910 178.820 27.230 178.880 ;
        RECT 30.590 178.820 30.910 178.880 ;
        RECT 34.820 178.865 34.960 179.360 ;
        RECT 41.185 179.315 41.475 179.360 ;
        RECT 44.850 179.300 45.170 179.560 ;
        RECT 49.910 179.300 50.230 179.560 ;
        RECT 54.510 179.500 54.830 179.560 ;
        RECT 55.905 179.500 56.195 179.545 ;
        RECT 51.385 179.360 56.195 179.500 ;
        RECT 36.570 178.960 36.890 179.220 ;
        RECT 37.505 179.160 37.795 179.205 ;
        RECT 43.930 179.160 44.250 179.220 ;
        RECT 51.385 179.160 51.525 179.360 ;
        RECT 54.510 179.300 54.830 179.360 ;
        RECT 55.905 179.315 56.195 179.360 ;
        RECT 58.190 179.500 58.510 179.560 ;
        RECT 64.170 179.500 64.490 179.560 ;
        RECT 65.105 179.500 65.395 179.545 ;
        RECT 58.190 179.360 63.020 179.500 ;
        RECT 37.505 179.020 44.250 179.160 ;
        RECT 37.505 178.975 37.795 179.020 ;
        RECT 43.930 178.960 44.250 179.020 ;
        RECT 44.480 179.020 51.525 179.160 ;
        RECT 44.480 178.865 44.620 179.020 ;
        RECT 51.765 178.975 52.055 179.205 ;
        RECT 54.985 179.160 55.275 179.205 ;
        RECT 54.140 179.020 55.275 179.160 ;
        RECT 26.910 178.680 30.910 178.820 ;
        RECT 25.545 178.635 25.835 178.680 ;
        RECT 26.910 178.620 27.230 178.680 ;
        RECT 30.590 178.620 30.910 178.680 ;
        RECT 32.445 178.635 32.735 178.865 ;
        RECT 34.745 178.635 35.035 178.865 ;
        RECT 37.045 178.820 37.335 178.865 ;
        RECT 44.405 178.820 44.695 178.865 ;
        RECT 37.045 178.680 44.695 178.820 ;
        RECT 37.045 178.635 37.335 178.680 ;
        RECT 44.405 178.635 44.695 178.680 ;
        RECT 45.310 178.820 45.630 178.880 ;
        RECT 47.625 178.820 47.915 178.865 ;
        RECT 48.070 178.820 48.390 178.880 ;
        RECT 45.310 178.680 48.390 178.820 ;
        RECT 25.990 178.480 26.310 178.540 ;
        RECT 25.200 178.340 26.310 178.480 ;
        RECT 21.405 178.295 21.695 178.340 ;
        RECT 22.310 178.280 22.630 178.340 ;
        RECT 25.990 178.280 26.310 178.340 ;
        RECT 29.225 178.480 29.515 178.525 ;
        RECT 32.520 178.480 32.660 178.635 ;
        RECT 45.310 178.620 45.630 178.680 ;
        RECT 47.625 178.635 47.915 178.680 ;
        RECT 48.070 178.620 48.390 178.680 ;
        RECT 49.005 178.820 49.295 178.865 ;
        RECT 51.290 178.820 51.610 178.880 ;
        RECT 51.840 178.820 51.980 178.975 ;
        RECT 53.605 178.820 53.895 178.865 ;
        RECT 49.005 178.680 51.060 178.820 ;
        RECT 49.005 178.635 49.295 178.680 ;
        RECT 29.225 178.340 32.660 178.480 ;
        RECT 29.225 178.295 29.515 178.340 ;
        RECT 33.350 178.280 33.670 178.540 ;
        RECT 33.810 178.280 34.130 178.540 ;
        RECT 34.270 178.280 34.590 178.540 ;
        RECT 35.665 178.295 35.955 178.525 ;
        RECT 36.125 178.480 36.415 178.525 ;
        RECT 37.490 178.480 37.810 178.540 ;
        RECT 36.125 178.340 37.810 178.480 ;
        RECT 36.125 178.295 36.415 178.340 ;
        RECT 20.485 178.140 20.775 178.185 ;
        RECT 24.610 178.140 24.930 178.200 ;
        RECT 20.485 178.000 24.930 178.140 ;
        RECT 20.485 177.955 20.775 178.000 ;
        RECT 21.940 177.860 22.080 178.000 ;
        RECT 24.610 177.940 24.930 178.000 ;
        RECT 30.605 178.140 30.895 178.185 ;
        RECT 35.190 178.140 35.510 178.200 ;
        RECT 30.605 178.000 35.510 178.140 ;
        RECT 30.605 177.955 30.895 178.000 ;
        RECT 35.190 177.940 35.510 178.000 ;
        RECT 21.850 177.600 22.170 177.860 ;
        RECT 22.310 177.600 22.630 177.860 ;
        RECT 29.210 177.800 29.530 177.860 ;
        RECT 29.685 177.800 29.975 177.845 ;
        RECT 29.210 177.660 29.975 177.800 ;
        RECT 35.740 177.800 35.880 178.295 ;
        RECT 37.490 178.280 37.810 178.340 ;
        RECT 37.950 178.530 38.270 178.540 ;
        RECT 37.950 178.525 38.410 178.530 ;
        RECT 37.950 178.295 38.495 178.525 ;
        RECT 37.950 178.280 38.270 178.295 ;
        RECT 38.870 178.280 39.190 178.540 ;
        RECT 40.250 178.480 40.570 178.540 ;
        RECT 40.055 178.340 40.570 178.480 ;
        RECT 40.250 178.280 40.570 178.340 ;
        RECT 40.710 178.280 41.030 178.540 ;
        RECT 42.090 178.280 42.410 178.540 ;
        RECT 43.010 178.280 43.330 178.540 ;
        RECT 43.930 178.525 44.250 178.540 ;
        RECT 43.715 178.295 44.250 178.525 ;
        RECT 43.930 178.280 44.250 178.295 ;
        RECT 44.850 178.480 45.170 178.540 ;
        RECT 45.785 178.480 46.075 178.525 ;
        RECT 44.850 178.340 46.075 178.480 ;
        RECT 44.850 178.280 45.170 178.340 ;
        RECT 45.785 178.295 46.075 178.340 ;
        RECT 46.245 178.295 46.535 178.525 ;
        RECT 49.910 178.480 50.230 178.540 ;
        RECT 50.385 178.480 50.675 178.525 ;
        RECT 49.910 178.340 50.675 178.480 ;
        RECT 39.345 178.140 39.635 178.185 ;
        RECT 39.345 178.000 40.020 178.140 ;
        RECT 39.345 177.955 39.635 178.000 ;
        RECT 39.880 177.860 40.020 178.000 ;
        RECT 38.870 177.800 39.190 177.860 ;
        RECT 35.740 177.660 39.190 177.800 ;
        RECT 29.210 177.600 29.530 177.660 ;
        RECT 29.685 177.615 29.975 177.660 ;
        RECT 38.870 177.600 39.190 177.660 ;
        RECT 39.790 177.600 40.110 177.860 ;
        RECT 40.340 177.800 40.480 178.280 ;
        RECT 42.550 177.940 42.870 178.200 ;
        RECT 45.310 177.800 45.630 177.860 ;
        RECT 40.340 177.660 45.630 177.800 ;
        RECT 46.320 177.800 46.460 178.295 ;
        RECT 49.910 178.280 50.230 178.340 ;
        RECT 50.385 178.295 50.675 178.340 ;
        RECT 48.085 178.140 48.375 178.185 ;
        RECT 48.530 178.140 48.850 178.200 ;
        RECT 48.085 178.000 48.850 178.140 ;
        RECT 48.085 177.955 48.375 178.000 ;
        RECT 48.530 177.940 48.850 178.000 ;
        RECT 49.005 178.140 49.295 178.185 ;
        RECT 49.450 178.140 49.770 178.200 ;
        RECT 49.005 178.000 49.770 178.140 ;
        RECT 49.005 177.955 49.295 178.000 ;
        RECT 49.450 177.940 49.770 178.000 ;
        RECT 46.690 177.800 47.010 177.860 ;
        RECT 50.920 177.845 51.060 178.680 ;
        RECT 51.290 178.680 53.895 178.820 ;
        RECT 51.290 178.620 51.610 178.680 ;
        RECT 53.605 178.635 53.895 178.680 ;
        RECT 51.750 178.480 52.070 178.540 ;
        RECT 52.670 178.480 52.990 178.540 ;
        RECT 54.140 178.480 54.280 179.020 ;
        RECT 54.985 178.975 55.275 179.020 ;
        RECT 55.980 178.820 56.120 179.315 ;
        RECT 58.190 179.300 58.510 179.360 ;
        RECT 59.570 179.160 59.890 179.220 ;
        RECT 59.200 179.020 59.890 179.160 ;
        RECT 59.200 178.820 59.340 179.020 ;
        RECT 59.570 178.960 59.890 179.020 ;
        RECT 60.045 178.975 60.335 179.205 ;
        RECT 60.490 179.160 60.810 179.220 ;
        RECT 61.425 179.160 61.715 179.205 ;
        RECT 60.490 179.020 61.715 179.160 ;
        RECT 62.880 179.160 63.020 179.360 ;
        RECT 64.170 179.360 65.395 179.500 ;
        RECT 64.170 179.300 64.490 179.360 ;
        RECT 65.105 179.315 65.395 179.360 ;
        RECT 66.010 179.300 66.330 179.560 ;
        RECT 71.530 179.500 71.850 179.560 ;
        RECT 83.505 179.500 83.795 179.545 ;
        RECT 71.530 179.360 83.795 179.500 ;
        RECT 71.530 179.300 71.850 179.360 ;
        RECT 83.505 179.315 83.795 179.360 ;
        RECT 72.910 179.160 73.230 179.220 ;
        RECT 62.880 179.020 64.400 179.160 ;
        RECT 60.120 178.820 60.260 178.975 ;
        RECT 60.490 178.960 60.810 179.020 ;
        RECT 61.425 178.975 61.715 179.020 ;
        RECT 63.710 178.820 64.030 178.880 ;
        RECT 55.980 178.680 59.340 178.820 ;
        RECT 56.810 178.480 57.130 178.540 ;
        RECT 59.200 178.525 59.340 178.680 ;
        RECT 59.660 178.680 60.260 178.820 ;
        RECT 60.580 178.680 64.030 178.820 ;
        RECT 59.660 178.540 59.800 178.680 ;
        RECT 57.285 178.480 57.575 178.525 ;
        RECT 51.750 178.340 52.990 178.480 ;
        RECT 51.750 178.280 52.070 178.340 ;
        RECT 52.670 178.280 52.990 178.340 ;
        RECT 53.220 178.340 54.280 178.480 ;
        RECT 54.600 178.340 57.575 178.480 ;
        RECT 53.220 178.200 53.360 178.340 ;
        RECT 53.130 177.940 53.450 178.200 ;
        RECT 46.320 177.660 47.010 177.800 ;
        RECT 45.310 177.600 45.630 177.660 ;
        RECT 46.690 177.600 47.010 177.660 ;
        RECT 50.845 177.800 51.135 177.845 ;
        RECT 54.600 177.800 54.740 178.340 ;
        RECT 56.810 178.280 57.130 178.340 ;
        RECT 57.285 178.295 57.575 178.340 ;
        RECT 59.125 178.295 59.415 178.525 ;
        RECT 59.570 178.280 59.890 178.540 ;
        RECT 54.970 178.140 55.290 178.200 ;
        RECT 58.205 178.140 58.495 178.185 ;
        RECT 54.970 178.000 58.495 178.140 ;
        RECT 54.970 177.940 55.290 178.000 ;
        RECT 58.205 177.955 58.495 178.000 ;
        RECT 50.845 177.660 54.740 177.800 ;
        RECT 58.280 177.800 58.420 177.955 ;
        RECT 58.650 177.940 58.970 178.200 ;
        RECT 60.580 177.800 60.720 178.680 ;
        RECT 63.710 178.620 64.030 178.680 ;
        RECT 61.410 178.280 61.730 178.540 ;
        RECT 61.870 178.480 62.190 178.540 ;
        RECT 63.250 178.525 63.570 178.540 ;
        RECT 64.260 178.525 64.400 179.020 ;
        RECT 68.400 179.020 73.230 179.160 ;
        RECT 66.930 178.820 67.250 178.880 ;
        RECT 68.400 178.820 68.540 179.020 ;
        RECT 72.910 178.960 73.230 179.020 ;
        RECT 77.510 178.960 77.830 179.220 ;
        RECT 80.730 179.160 81.050 179.220 ;
        RECT 81.665 179.160 81.955 179.205 ;
        RECT 80.730 179.020 81.955 179.160 ;
        RECT 80.730 178.960 81.050 179.020 ;
        RECT 81.665 178.975 81.955 179.020 ;
        RECT 83.950 179.160 84.270 179.220 ;
        RECT 83.950 179.020 85.100 179.160 ;
        RECT 83.950 178.960 84.270 179.020 ;
        RECT 66.930 178.680 68.540 178.820 ;
        RECT 66.930 178.620 67.250 178.680 ;
        RECT 62.805 178.480 63.095 178.525 ;
        RECT 61.870 178.340 63.095 178.480 ;
        RECT 61.870 178.280 62.190 178.340 ;
        RECT 62.805 178.295 63.095 178.340 ;
        RECT 63.250 178.295 63.580 178.525 ;
        RECT 64.185 178.295 64.475 178.525 ;
        RECT 65.550 178.480 65.870 178.540 ;
        RECT 68.400 178.525 68.540 178.680 ;
        RECT 69.320 178.680 84.640 178.820 ;
        RECT 69.320 178.540 69.460 178.680 ;
        RECT 84.500 178.540 84.640 178.680 ;
        RECT 67.405 178.480 67.695 178.525 ;
        RECT 65.550 178.340 67.695 178.480 ;
        RECT 63.250 178.280 63.570 178.295 ;
        RECT 65.550 178.280 65.870 178.340 ;
        RECT 67.405 178.295 67.695 178.340 ;
        RECT 67.865 178.295 68.155 178.525 ;
        RECT 68.325 178.295 68.615 178.525 ;
        RECT 62.330 177.940 62.650 178.200 ;
        RECT 67.940 178.140 68.080 178.295 ;
        RECT 69.230 178.280 69.550 178.540 ;
        RECT 69.690 178.280 70.010 178.540 ;
        RECT 71.070 178.280 71.390 178.540 ;
        RECT 73.830 178.480 74.150 178.540 ;
        RECT 72.540 178.340 74.150 178.480 ;
        RECT 72.540 178.140 72.680 178.340 ;
        RECT 73.830 178.280 74.150 178.340 ;
        RECT 74.290 178.480 74.610 178.540 ;
        RECT 77.970 178.480 78.290 178.540 ;
        RECT 80.285 178.480 80.575 178.525 ;
        RECT 74.290 178.340 80.575 178.480 ;
        RECT 74.290 178.280 74.610 178.340 ;
        RECT 77.970 178.280 78.290 178.340 ;
        RECT 80.285 178.295 80.575 178.340 ;
        RECT 81.190 178.280 81.510 178.540 ;
        RECT 84.410 178.280 84.730 178.540 ;
        RECT 84.960 178.480 85.100 179.020 ;
        RECT 85.330 178.960 85.650 179.220 ;
        RECT 85.805 178.480 86.095 178.525 ;
        RECT 84.960 178.340 86.095 178.480 ;
        RECT 85.805 178.295 86.095 178.340 ;
        RECT 86.265 178.295 86.555 178.525 ;
        RECT 67.940 178.000 72.680 178.140 ;
        RECT 72.910 178.140 73.230 178.200 ;
        RECT 86.340 178.140 86.480 178.295 ;
        RECT 72.910 178.000 86.480 178.140 ;
        RECT 69.320 177.860 69.460 178.000 ;
        RECT 72.910 177.940 73.230 178.000 ;
        RECT 58.280 177.660 60.720 177.800 ;
        RECT 50.845 177.615 51.135 177.660 ;
        RECT 69.230 177.600 69.550 177.860 ;
        RECT 70.165 177.800 70.455 177.845 ;
        RECT 70.610 177.800 70.930 177.860 ;
        RECT 70.165 177.660 70.930 177.800 ;
        RECT 70.165 177.615 70.455 177.660 ;
        RECT 70.610 177.600 70.930 177.660 ;
        RECT 87.170 177.600 87.490 177.860 ;
        RECT 18.100 176.980 89.400 177.460 ;
        RECT 26.005 176.595 26.295 176.825 ;
        RECT 33.350 176.780 33.670 176.840 ;
        RECT 40.250 176.780 40.570 176.840 ;
        RECT 46.245 176.780 46.535 176.825 ;
        RECT 33.350 176.640 46.535 176.780 ;
        RECT 17.710 176.440 18.030 176.500 ;
        RECT 26.080 176.440 26.220 176.595 ;
        RECT 33.350 176.580 33.670 176.640 ;
        RECT 40.250 176.580 40.570 176.640 ;
        RECT 46.245 176.595 46.535 176.640 ;
        RECT 47.150 176.580 47.470 176.840 ;
        RECT 48.530 176.630 48.850 176.840 ;
        RECT 51.305 176.780 51.595 176.825 ;
        RECT 53.130 176.780 53.450 176.840 ;
        RECT 49.080 176.640 49.680 176.780 ;
        RECT 49.080 176.630 49.220 176.640 ;
        RECT 48.530 176.580 49.220 176.630 ;
        RECT 17.710 176.300 26.220 176.440 ;
        RECT 33.825 176.440 34.115 176.485 ;
        RECT 35.650 176.440 35.970 176.500 ;
        RECT 33.825 176.300 35.970 176.440 ;
        RECT 17.710 176.240 18.030 176.300 ;
        RECT 33.825 176.255 34.115 176.300 ;
        RECT 35.650 176.240 35.970 176.300 ;
        RECT 42.550 176.440 42.870 176.500 ;
        RECT 48.625 176.490 49.220 176.580 ;
        RECT 49.540 176.440 49.680 176.640 ;
        RECT 51.305 176.640 53.450 176.780 ;
        RECT 51.305 176.595 51.595 176.640 ;
        RECT 53.130 176.580 53.450 176.640 ;
        RECT 63.250 176.780 63.570 176.840 ;
        RECT 65.105 176.780 65.395 176.825 ;
        RECT 63.250 176.640 65.395 176.780 ;
        RECT 63.250 176.580 63.570 176.640 ;
        RECT 60.030 176.440 60.350 176.500 ;
        RECT 61.885 176.440 62.175 176.485 ;
        RECT 42.550 176.300 46.000 176.440 ;
        RECT 49.540 176.300 57.040 176.440 ;
        RECT 42.550 176.240 42.870 176.300 ;
        RECT 45.860 176.160 46.000 176.300 ;
        RECT 19.550 175.900 19.870 176.160 ;
        RECT 21.850 175.900 22.170 176.160 ;
        RECT 22.635 176.100 22.925 176.145 ;
        RECT 24.610 176.100 24.930 176.160 ;
        RECT 22.635 175.960 24.930 176.100 ;
        RECT 22.635 175.915 22.925 175.960 ;
        RECT 24.610 175.900 24.930 175.960 ;
        RECT 25.070 176.100 25.390 176.160 ;
        RECT 25.545 176.100 25.835 176.145 ;
        RECT 25.070 175.960 25.835 176.100 ;
        RECT 25.070 175.900 25.390 175.960 ;
        RECT 25.545 175.915 25.835 175.960 ;
        RECT 26.910 175.900 27.230 176.160 ;
        RECT 27.385 175.915 27.675 176.145 ;
        RECT 33.365 175.915 33.655 176.145 ;
        RECT 34.270 176.100 34.590 176.160 ;
        RECT 39.790 176.100 40.110 176.160 ;
        RECT 34.270 175.960 40.110 176.100 ;
        RECT 17.250 175.760 17.570 175.820 ;
        RECT 27.460 175.760 27.600 175.915 ;
        RECT 17.250 175.620 27.600 175.760 ;
        RECT 33.440 175.760 33.580 175.915 ;
        RECT 34.270 175.900 34.590 175.960 ;
        RECT 39.790 175.900 40.110 175.960 ;
        RECT 45.325 175.915 45.615 176.145 ;
        RECT 33.810 175.760 34.130 175.820 ;
        RECT 36.110 175.760 36.430 175.820 ;
        RECT 33.440 175.620 36.430 175.760 ;
        RECT 17.250 175.560 17.570 175.620 ;
        RECT 33.810 175.560 34.130 175.620 ;
        RECT 36.110 175.560 36.430 175.620 ;
        RECT 44.850 175.760 45.170 175.820 ;
        RECT 45.400 175.760 45.540 175.915 ;
        RECT 45.770 175.900 46.090 176.160 ;
        RECT 47.150 176.100 47.470 176.160 ;
        RECT 47.625 176.100 47.915 176.145 ;
        RECT 47.150 175.960 47.915 176.100 ;
        RECT 48.990 176.020 49.310 176.280 ;
        RECT 47.150 175.900 47.470 175.960 ;
        RECT 47.625 175.915 47.915 175.960 ;
        RECT 49.005 175.915 49.295 176.020 ;
        RECT 49.925 175.915 50.215 176.145 ;
        RECT 50.370 176.100 50.690 176.160 ;
        RECT 50.845 176.100 51.135 176.145 ;
        RECT 50.370 175.960 51.135 176.100 ;
        RECT 44.850 175.620 45.540 175.760 ;
        RECT 45.860 175.620 49.225 175.760 ;
        RECT 44.850 175.560 45.170 175.620 ;
        RECT 45.860 175.480 46.000 175.620 ;
        RECT 23.690 175.220 24.010 175.480 ;
        RECT 28.290 175.220 28.610 175.480 ;
        RECT 44.405 175.420 44.695 175.465 ;
        RECT 45.770 175.420 46.090 175.480 ;
        RECT 44.405 175.280 46.090 175.420 ;
        RECT 44.405 175.235 44.695 175.280 ;
        RECT 45.770 175.220 46.090 175.280 ;
        RECT 20.470 174.880 20.790 175.140 ;
        RECT 24.610 174.880 24.930 175.140 ;
        RECT 38.870 175.080 39.190 175.140 ;
        RECT 40.710 175.080 41.030 175.140 ;
        RECT 38.870 174.940 41.030 175.080 ;
        RECT 38.870 174.880 39.190 174.940 ;
        RECT 40.710 174.880 41.030 174.940 ;
        RECT 46.690 175.080 47.010 175.140 ;
        RECT 47.625 175.080 47.915 175.125 ;
        RECT 46.690 174.940 47.915 175.080 ;
        RECT 49.085 175.080 49.225 175.620 ;
        RECT 49.450 175.420 49.770 175.480 ;
        RECT 50.000 175.420 50.140 175.915 ;
        RECT 50.370 175.900 50.690 175.960 ;
        RECT 50.845 175.915 51.135 175.960 ;
        RECT 52.225 176.100 52.515 176.145 ;
        RECT 53.130 176.100 53.450 176.160 ;
        RECT 52.225 175.960 53.450 176.100 ;
        RECT 52.225 175.915 52.515 175.960 ;
        RECT 53.130 175.900 53.450 175.960 ;
        RECT 53.590 175.900 53.910 176.160 ;
        RECT 54.050 175.900 54.370 176.160 ;
        RECT 54.985 176.100 55.275 176.145 ;
        RECT 55.890 176.100 56.210 176.160 ;
        RECT 54.985 175.960 56.210 176.100 ;
        RECT 54.985 175.915 55.275 175.960 ;
        RECT 55.890 175.900 56.210 175.960 ;
        RECT 56.350 175.900 56.670 176.160 ;
        RECT 56.900 176.100 57.040 176.300 ;
        RECT 60.030 176.300 62.175 176.440 ;
        RECT 60.030 176.240 60.350 176.300 ;
        RECT 61.885 176.255 62.175 176.300 ;
        RECT 63.800 176.255 63.940 176.640 ;
        RECT 65.105 176.595 65.395 176.640 ;
        RECT 71.070 176.780 71.390 176.840 ;
        RECT 78.430 176.780 78.750 176.840 ;
        RECT 71.070 176.640 78.750 176.780 ;
        RECT 71.070 176.580 71.390 176.640 ;
        RECT 64.630 176.440 64.950 176.500 ;
        RECT 69.230 176.440 69.550 176.500 ;
        RECT 72.080 176.485 72.220 176.640 ;
        RECT 78.430 176.580 78.750 176.640 ;
        RECT 81.190 176.780 81.510 176.840 ;
        RECT 84.410 176.780 84.730 176.840 ;
        RECT 81.190 176.640 84.730 176.780 ;
        RECT 81.190 176.580 81.510 176.640 ;
        RECT 84.410 176.580 84.730 176.640 ;
        RECT 71.545 176.440 71.835 176.485 ;
        RECT 64.630 176.300 69.000 176.440 ;
        RECT 60.505 176.100 60.795 176.145 ;
        RECT 60.950 176.100 61.270 176.160 ;
        RECT 56.900 175.960 59.800 176.100 ;
        RECT 54.525 175.760 54.815 175.805 ;
        RECT 50.920 175.620 54.815 175.760 ;
        RECT 50.920 175.480 51.060 175.620 ;
        RECT 54.525 175.575 54.815 175.620 ;
        RECT 57.745 175.575 58.035 175.805 ;
        RECT 58.205 175.760 58.495 175.805 ;
        RECT 59.110 175.760 59.430 175.820 ;
        RECT 58.205 175.620 59.430 175.760 ;
        RECT 59.660 175.760 59.800 175.960 ;
        RECT 60.505 175.960 61.270 176.100 ;
        RECT 60.505 175.915 60.795 175.960 ;
        RECT 60.950 175.900 61.270 175.960 ;
        RECT 61.410 175.900 61.730 176.160 ;
        RECT 62.330 176.100 62.650 176.160 ;
        RECT 62.805 176.100 63.095 176.145 ;
        RECT 62.330 175.960 63.095 176.100 ;
        RECT 62.330 175.900 62.650 175.960 ;
        RECT 62.805 175.915 63.095 175.960 ;
        RECT 60.045 175.760 60.335 175.805 ;
        RECT 59.660 175.620 62.560 175.760 ;
        RECT 58.205 175.575 58.495 175.620 ;
        RECT 49.450 175.280 50.140 175.420 ;
        RECT 49.450 175.220 49.770 175.280 ;
        RECT 50.370 175.220 50.690 175.480 ;
        RECT 50.830 175.220 51.150 175.480 ;
        RECT 52.685 175.420 52.975 175.465 ;
        RECT 54.970 175.420 55.290 175.480 ;
        RECT 52.685 175.280 55.290 175.420 ;
        RECT 52.685 175.235 52.975 175.280 ;
        RECT 54.970 175.220 55.290 175.280 ;
        RECT 55.445 175.420 55.735 175.465 ;
        RECT 57.820 175.420 57.960 175.575 ;
        RECT 59.110 175.560 59.430 175.620 ;
        RECT 60.045 175.575 60.335 175.620 ;
        RECT 61.885 175.420 62.175 175.465 ;
        RECT 55.445 175.280 57.500 175.420 ;
        RECT 57.820 175.280 62.175 175.420 ;
        RECT 55.445 175.235 55.735 175.280 ;
        RECT 51.290 175.080 51.610 175.140 ;
        RECT 49.085 174.940 51.610 175.080 ;
        RECT 46.690 174.880 47.010 174.940 ;
        RECT 47.625 174.895 47.915 174.940 ;
        RECT 51.290 174.880 51.610 174.940 ;
        RECT 55.890 175.080 56.210 175.140 ;
        RECT 56.825 175.080 57.115 175.125 ;
        RECT 55.890 174.940 57.115 175.080 ;
        RECT 57.360 175.080 57.500 175.280 ;
        RECT 61.885 175.235 62.175 175.280 ;
        RECT 58.190 175.080 58.510 175.140 ;
        RECT 57.360 174.940 58.510 175.080 ;
        RECT 55.890 174.880 56.210 174.940 ;
        RECT 56.825 174.895 57.115 174.940 ;
        RECT 58.190 174.880 58.510 174.940 ;
        RECT 59.110 175.080 59.430 175.140 ;
        RECT 60.965 175.080 61.255 175.125 ;
        RECT 59.110 174.940 61.255 175.080 ;
        RECT 59.110 174.880 59.430 174.940 ;
        RECT 60.965 174.895 61.255 174.940 ;
        RECT 61.410 175.080 61.730 175.140 ;
        RECT 62.420 175.080 62.560 175.620 ;
        RECT 62.880 175.420 63.020 175.915 ;
        RECT 63.250 175.900 63.570 176.160 ;
        RECT 63.750 176.025 64.040 176.255 ;
        RECT 64.630 176.240 64.950 176.300 ;
        RECT 66.485 176.100 66.775 176.145 ;
        RECT 64.720 175.960 66.775 176.100 ;
        RECT 64.720 175.820 64.860 175.960 ;
        RECT 66.485 175.915 66.775 175.960 ;
        RECT 67.390 176.100 67.710 176.160 ;
        RECT 67.865 176.100 68.155 176.145 ;
        RECT 67.390 175.960 68.155 176.100 ;
        RECT 67.390 175.900 67.710 175.960 ;
        RECT 67.865 175.915 68.155 175.960 ;
        RECT 64.630 175.560 64.950 175.820 ;
        RECT 65.550 175.760 65.870 175.820 ;
        RECT 66.025 175.760 66.315 175.805 ;
        RECT 65.550 175.620 66.315 175.760 ;
        RECT 65.550 175.560 65.870 175.620 ;
        RECT 66.025 175.575 66.315 175.620 ;
        RECT 66.930 175.760 67.250 175.820 ;
        RECT 68.325 175.760 68.615 175.805 ;
        RECT 66.930 175.620 68.615 175.760 ;
        RECT 68.860 175.760 69.000 176.300 ;
        RECT 69.230 176.300 71.835 176.440 ;
        RECT 69.230 176.240 69.550 176.300 ;
        RECT 71.545 176.255 71.835 176.300 ;
        RECT 72.005 176.255 72.295 176.485 ;
        RECT 77.985 176.440 78.275 176.485 ;
        RECT 81.650 176.440 81.970 176.500 ;
        RECT 77.985 176.300 81.970 176.440 ;
        RECT 77.985 176.255 78.275 176.300 ;
        RECT 81.650 176.240 81.970 176.300 ;
        RECT 71.070 175.900 71.390 176.160 ;
        RECT 72.925 175.915 73.215 176.145 ;
        RECT 74.305 176.100 74.595 176.145 ;
        RECT 75.210 176.100 75.530 176.160 ;
        RECT 77.050 176.100 77.370 176.160 ;
        RECT 74.305 175.960 77.370 176.100 ;
        RECT 74.305 175.915 74.595 175.960 ;
        RECT 73.000 175.760 73.140 175.915 ;
        RECT 75.210 175.900 75.530 175.960 ;
        RECT 77.050 175.900 77.370 175.960 ;
        RECT 74.750 175.760 75.070 175.820 ;
        RECT 75.685 175.760 75.975 175.805 ;
        RECT 68.860 175.620 74.520 175.760 ;
        RECT 66.930 175.560 67.250 175.620 ;
        RECT 68.325 175.575 68.615 175.620 ;
        RECT 70.165 175.420 70.455 175.465 ;
        RECT 62.880 175.280 70.455 175.420 ;
        RECT 70.165 175.235 70.455 175.280 ;
        RECT 71.530 175.420 71.850 175.480 ;
        RECT 73.370 175.420 73.690 175.480 ;
        RECT 71.530 175.280 73.690 175.420 ;
        RECT 74.380 175.420 74.520 175.620 ;
        RECT 74.750 175.620 75.975 175.760 ;
        RECT 74.750 175.560 75.070 175.620 ;
        RECT 75.685 175.575 75.975 175.620 ;
        RECT 76.130 175.760 76.450 175.820 ;
        RECT 79.350 175.760 79.670 175.820 ;
        RECT 76.130 175.620 79.670 175.760 ;
        RECT 76.130 175.560 76.450 175.620 ;
        RECT 79.350 175.560 79.670 175.620 ;
        RECT 83.950 175.420 84.270 175.480 ;
        RECT 74.380 175.280 84.270 175.420 ;
        RECT 71.530 175.220 71.850 175.280 ;
        RECT 73.370 175.220 73.690 175.280 ;
        RECT 83.950 175.220 84.270 175.280 ;
        RECT 61.410 174.940 62.560 175.080 ;
        RECT 63.710 175.080 64.030 175.140 ;
        RECT 64.630 175.080 64.950 175.140 ;
        RECT 63.710 174.940 64.950 175.080 ;
        RECT 61.410 174.880 61.730 174.940 ;
        RECT 63.710 174.880 64.030 174.940 ;
        RECT 64.630 174.880 64.950 174.940 ;
        RECT 65.550 175.080 65.870 175.140 ;
        RECT 66.930 175.080 67.250 175.140 ;
        RECT 65.550 174.940 67.250 175.080 ;
        RECT 65.550 174.880 65.870 174.940 ;
        RECT 66.930 174.880 67.250 174.940 ;
        RECT 71.070 175.080 71.390 175.140 ;
        RECT 76.130 175.080 76.450 175.140 ;
        RECT 71.070 174.940 76.450 175.080 ;
        RECT 71.070 174.880 71.390 174.940 ;
        RECT 76.130 174.880 76.450 174.940 ;
        RECT 83.030 175.080 83.350 175.140 ;
        RECT 84.410 175.080 84.730 175.140 ;
        RECT 83.030 174.940 84.730 175.080 ;
        RECT 83.030 174.880 83.350 174.940 ;
        RECT 84.410 174.880 84.730 174.940 ;
        RECT 18.100 174.260 89.400 174.740 ;
        RECT 33.825 174.060 34.115 174.105 ;
        RECT 41.630 174.060 41.950 174.120 ;
        RECT 55.430 174.060 55.750 174.120 ;
        RECT 61.885 174.060 62.175 174.105 ;
        RECT 63.250 174.060 63.570 174.120 ;
        RECT 33.825 173.920 41.950 174.060 ;
        RECT 33.825 173.875 34.115 173.920 ;
        RECT 41.630 173.860 41.950 173.920 ;
        RECT 51.200 173.920 55.750 174.060 ;
        RECT 34.270 173.720 34.590 173.780 ;
        RECT 21.940 173.580 34.590 173.720 ;
        RECT 20.010 173.380 20.330 173.440 ;
        RECT 21.940 173.380 22.080 173.580 ;
        RECT 34.270 173.520 34.590 173.580 ;
        RECT 39.330 173.720 39.650 173.780 ;
        RECT 51.200 173.720 51.340 173.920 ;
        RECT 55.430 173.860 55.750 173.920 ;
        RECT 55.980 173.920 58.880 174.060 ;
        RECT 39.330 173.580 51.340 173.720 ;
        RECT 51.765 173.720 52.055 173.765 ;
        RECT 53.130 173.720 53.450 173.780 ;
        RECT 51.765 173.580 53.450 173.720 ;
        RECT 39.330 173.520 39.650 173.580 ;
        RECT 51.765 173.535 52.055 173.580 ;
        RECT 53.130 173.520 53.450 173.580 ;
        RECT 54.525 173.535 54.815 173.765 ;
        RECT 54.970 173.720 55.290 173.780 ;
        RECT 55.980 173.720 56.120 173.920 ;
        RECT 54.970 173.580 56.120 173.720 ;
        RECT 57.745 173.720 58.035 173.765 ;
        RECT 58.190 173.720 58.510 173.780 ;
        RECT 57.745 173.580 58.510 173.720 ;
        RECT 58.740 173.720 58.880 173.920 ;
        RECT 61.885 173.920 63.570 174.060 ;
        RECT 61.885 173.875 62.175 173.920 ;
        RECT 63.250 173.860 63.570 173.920 ;
        RECT 64.630 174.060 64.950 174.120 ;
        RECT 65.565 174.060 65.855 174.105 ;
        RECT 64.630 173.920 65.855 174.060 ;
        RECT 64.630 173.860 64.950 173.920 ;
        RECT 65.565 173.875 65.855 173.920 ;
        RECT 67.865 174.060 68.155 174.105 ;
        RECT 70.150 174.060 70.470 174.120 ;
        RECT 73.370 174.060 73.690 174.120 ;
        RECT 67.865 173.920 70.470 174.060 ;
        RECT 67.865 173.875 68.155 173.920 ;
        RECT 70.150 173.860 70.470 173.920 ;
        RECT 71.160 173.920 73.690 174.060 ;
        RECT 58.740 173.580 68.540 173.720 ;
        RECT 20.010 173.240 22.080 173.380 ;
        RECT 20.010 173.180 20.330 173.240 ;
        RECT 21.390 172.840 21.710 173.100 ;
        RECT 21.940 173.085 22.080 173.240 ;
        RECT 22.770 173.180 23.090 173.440 ;
        RECT 24.610 173.380 24.930 173.440 ;
        RECT 43.470 173.380 43.790 173.440 ;
        RECT 54.600 173.380 54.740 173.535 ;
        RECT 54.970 173.520 55.290 173.580 ;
        RECT 57.745 173.535 58.035 173.580 ;
        RECT 58.190 173.520 58.510 173.580 ;
        RECT 24.610 173.240 43.790 173.380 ;
        RECT 24.610 173.180 24.930 173.240 ;
        RECT 43.470 173.180 43.790 173.240 ;
        RECT 51.840 173.240 54.740 173.380 ;
        RECT 55.430 173.380 55.750 173.440 ;
        RECT 63.250 173.380 63.570 173.440 ;
        RECT 55.430 173.240 59.340 173.380 ;
        RECT 21.865 172.855 22.155 173.085 ;
        RECT 23.245 173.040 23.535 173.085 ;
        RECT 27.830 173.040 28.150 173.100 ;
        RECT 23.245 172.900 28.150 173.040 ;
        RECT 23.245 172.855 23.535 172.900 ;
        RECT 27.830 172.840 28.150 172.900 ;
        RECT 28.750 172.840 29.070 173.100 ;
        RECT 31.510 172.840 31.830 173.100 ;
        RECT 32.905 172.855 33.195 173.085 ;
        RECT 36.110 173.040 36.430 173.100 ;
        RECT 38.425 173.040 38.715 173.085 ;
        RECT 36.110 172.900 38.715 173.040 ;
        RECT 28.840 172.700 28.980 172.840 ;
        RECT 32.980 172.700 33.120 172.855 ;
        RECT 36.110 172.840 36.430 172.900 ;
        RECT 38.425 172.855 38.715 172.900 ;
        RECT 39.345 173.040 39.635 173.085 ;
        RECT 42.090 173.040 42.410 173.100 ;
        RECT 51.840 173.085 51.980 173.240 ;
        RECT 55.430 173.180 55.750 173.240 ;
        RECT 39.345 172.900 42.410 173.040 ;
        RECT 39.345 172.855 39.635 172.900 ;
        RECT 42.090 172.840 42.410 172.900 ;
        RECT 51.765 172.855 52.055 173.085 ;
        RECT 53.130 172.840 53.450 173.100 ;
        RECT 55.890 172.840 56.210 173.100 ;
        RECT 59.200 173.085 59.340 173.240 ;
        RECT 61.500 173.240 63.570 173.380 ;
        RECT 58.665 173.040 58.955 173.085 ;
        RECT 58.280 172.900 58.955 173.040 ;
        RECT 28.840 172.560 33.120 172.700 ;
        RECT 54.510 172.500 54.830 172.760 ;
        RECT 56.350 172.500 56.670 172.760 ;
        RECT 58.280 172.700 58.420 172.900 ;
        RECT 58.665 172.855 58.955 172.900 ;
        RECT 59.125 172.855 59.415 173.085 ;
        RECT 59.585 172.855 59.875 173.085 ;
        RECT 60.030 173.040 60.350 173.100 ;
        RECT 61.500 173.085 61.640 173.240 ;
        RECT 63.250 173.180 63.570 173.240 ;
        RECT 63.710 173.380 64.030 173.440 ;
        RECT 63.710 173.240 66.240 173.380 ;
        RECT 63.710 173.180 64.030 173.240 ;
        RECT 60.505 173.040 60.795 173.085 ;
        RECT 60.030 172.900 60.795 173.040 ;
        RECT 59.660 172.700 59.800 172.855 ;
        RECT 60.030 172.840 60.350 172.900 ;
        RECT 60.505 172.855 60.795 172.900 ;
        RECT 61.425 172.855 61.715 173.085 ;
        RECT 62.330 173.040 62.650 173.100 ;
        RECT 62.805 173.040 63.095 173.085 ;
        RECT 62.330 172.900 63.095 173.040 ;
        RECT 62.330 172.840 62.650 172.900 ;
        RECT 62.805 172.855 63.095 172.900 ;
        RECT 64.170 172.840 64.490 173.100 ;
        RECT 64.630 172.840 64.950 173.100 ;
        RECT 58.280 172.560 58.880 172.700 ;
        RECT 59.660 172.560 60.260 172.700 ;
        RECT 20.485 172.360 20.775 172.405 ;
        RECT 28.750 172.360 29.070 172.420 ;
        RECT 20.485 172.220 29.070 172.360 ;
        RECT 20.485 172.175 20.775 172.220 ;
        RECT 28.750 172.160 29.070 172.220 ;
        RECT 30.590 172.360 30.910 172.420 ;
        RECT 31.985 172.360 32.275 172.405 ;
        RECT 30.590 172.220 32.275 172.360 ;
        RECT 30.590 172.160 30.910 172.220 ;
        RECT 31.985 172.175 32.275 172.220 ;
        RECT 38.870 172.160 39.190 172.420 ;
        RECT 44.390 172.360 44.710 172.420 ;
        RECT 51.750 172.360 52.070 172.420 ;
        RECT 52.685 172.360 52.975 172.405 ;
        RECT 44.390 172.220 52.975 172.360 ;
        RECT 44.390 172.160 44.710 172.220 ;
        RECT 51.750 172.160 52.070 172.220 ;
        RECT 52.685 172.175 52.975 172.220 ;
        RECT 53.590 172.360 53.910 172.420 ;
        RECT 54.050 172.360 54.370 172.420 ;
        RECT 53.590 172.220 54.370 172.360 ;
        RECT 53.590 172.160 53.910 172.220 ;
        RECT 54.050 172.160 54.370 172.220 ;
        RECT 55.430 172.160 55.750 172.420 ;
        RECT 56.440 172.360 56.580 172.500 ;
        RECT 58.190 172.360 58.510 172.420 ;
        RECT 56.440 172.220 58.510 172.360 ;
        RECT 58.740 172.360 58.880 172.560 ;
        RECT 60.120 172.420 60.260 172.560 ;
        RECT 63.250 172.500 63.570 172.760 ;
        RECT 63.725 172.700 64.015 172.745 ;
        RECT 64.260 172.700 64.400 172.840 ;
        RECT 63.725 172.560 64.400 172.700 ;
        RECT 66.100 172.700 66.240 173.240 ;
        RECT 66.485 173.100 66.775 173.165 ;
        RECT 66.470 172.840 66.790 173.100 ;
        RECT 66.930 172.840 67.250 173.100 ;
        RECT 67.850 172.840 68.170 173.100 ;
        RECT 68.400 173.085 68.540 173.580 ;
        RECT 69.690 173.180 70.010 173.440 ;
        RECT 71.160 173.380 71.300 173.920 ;
        RECT 73.370 173.860 73.690 173.920 ;
        RECT 74.290 173.860 74.610 174.120 ;
        RECT 74.750 174.060 75.070 174.120 ;
        RECT 77.510 174.060 77.830 174.120 ;
        RECT 74.750 173.920 77.830 174.060 ;
        RECT 74.750 173.860 75.070 173.920 ;
        RECT 77.510 173.860 77.830 173.920 ;
        RECT 80.745 174.060 81.035 174.105 ;
        RECT 82.110 174.060 82.430 174.120 ;
        RECT 80.745 173.920 82.430 174.060 ;
        RECT 80.745 173.875 81.035 173.920 ;
        RECT 82.110 173.860 82.430 173.920 ;
        RECT 83.505 174.060 83.795 174.105 ;
        RECT 83.950 174.060 84.270 174.120 ;
        RECT 83.505 173.920 84.270 174.060 ;
        RECT 83.505 173.875 83.795 173.920 ;
        RECT 83.950 173.860 84.270 173.920 ;
        RECT 85.790 174.060 86.110 174.120 ;
        RECT 89.010 174.060 89.330 174.120 ;
        RECT 85.790 173.920 89.330 174.060 ;
        RECT 85.790 173.860 86.110 173.920 ;
        RECT 89.010 173.860 89.330 173.920 ;
        RECT 71.990 173.520 72.310 173.780 ;
        RECT 74.840 173.720 74.980 173.860 ;
        RECT 78.890 173.720 79.210 173.780 ;
        RECT 73.920 173.580 74.980 173.720 ;
        RECT 75.300 173.580 79.210 173.720 ;
        RECT 70.700 173.240 71.300 173.380 ;
        RECT 73.385 173.380 73.675 173.425 ;
        RECT 73.920 173.380 74.060 173.580 ;
        RECT 74.750 173.425 75.070 173.440 ;
        RECT 75.300 173.425 75.440 173.580 ;
        RECT 78.890 173.520 79.210 173.580 ;
        RECT 79.350 173.720 79.670 173.780 ;
        RECT 79.350 173.580 86.480 173.720 ;
        RECT 79.350 173.520 79.670 173.580 ;
        RECT 73.385 173.240 74.060 173.380 ;
        RECT 70.700 173.085 70.840 173.240 ;
        RECT 73.385 173.195 73.675 173.240 ;
        RECT 74.725 173.195 75.070 173.425 ;
        RECT 75.225 173.195 75.515 173.425 ;
        RECT 84.410 173.380 84.730 173.440 ;
        RECT 85.790 173.380 86.110 173.440 ;
        RECT 78.980 173.240 84.730 173.380 ;
        RECT 74.750 173.180 75.070 173.195 ;
        RECT 68.325 172.855 68.615 173.085 ;
        RECT 70.625 172.855 70.915 173.085 ;
        RECT 71.530 172.840 71.850 173.100 ;
        RECT 72.465 172.855 72.755 173.085 ;
        RECT 68.785 172.700 69.075 172.745 ;
        RECT 72.540 172.700 72.680 172.855 ;
        RECT 76.130 172.840 76.450 173.100 ;
        RECT 76.590 172.840 76.910 173.100 ;
        RECT 77.525 172.855 77.815 173.085 ;
        RECT 77.970 173.040 78.290 173.100 ;
        RECT 78.980 173.085 79.120 173.240 ;
        RECT 84.410 173.180 84.730 173.240 ;
        RECT 84.960 173.240 86.110 173.380 ;
        RECT 78.905 173.040 79.195 173.085 ;
        RECT 77.970 172.900 79.195 173.040 ;
        RECT 77.600 172.700 77.740 172.855 ;
        RECT 77.970 172.840 78.290 172.900 ;
        RECT 78.905 172.855 79.195 172.900 ;
        RECT 81.205 172.855 81.495 173.085 ;
        RECT 83.965 173.040 84.255 173.085 ;
        RECT 84.960 173.040 85.100 173.240 ;
        RECT 85.790 173.180 86.110 173.240 ;
        RECT 83.965 172.900 85.100 173.040 ;
        RECT 83.965 172.855 84.255 172.900 ;
        RECT 66.100 172.560 77.740 172.700 ;
        RECT 81.280 172.700 81.420 172.855 ;
        RECT 85.330 172.840 85.650 173.100 ;
        RECT 86.340 173.085 86.480 173.580 ;
        RECT 86.265 172.855 86.555 173.085 ;
        RECT 88.550 172.700 88.870 172.760 ;
        RECT 81.280 172.560 88.870 172.700 ;
        RECT 63.725 172.515 64.015 172.560 ;
        RECT 68.785 172.515 69.075 172.560 ;
        RECT 88.550 172.500 88.870 172.560 ;
        RECT 59.570 172.360 59.890 172.420 ;
        RECT 58.740 172.220 59.890 172.360 ;
        RECT 58.190 172.160 58.510 172.220 ;
        RECT 59.570 172.160 59.890 172.220 ;
        RECT 60.030 172.160 60.350 172.420 ;
        RECT 60.950 172.160 61.270 172.420 ;
        RECT 61.870 172.360 62.190 172.420 ;
        RECT 66.930 172.360 67.250 172.420 ;
        RECT 61.870 172.220 67.250 172.360 ;
        RECT 61.870 172.160 62.190 172.220 ;
        RECT 66.930 172.160 67.250 172.220 ;
        RECT 70.150 172.360 70.470 172.420 ;
        RECT 72.925 172.360 73.215 172.405 ;
        RECT 77.065 172.360 77.355 172.405 ;
        RECT 70.150 172.220 77.355 172.360 ;
        RECT 70.150 172.160 70.470 172.220 ;
        RECT 72.925 172.175 73.215 172.220 ;
        RECT 77.065 172.175 77.355 172.220 ;
        RECT 77.985 172.360 78.275 172.405 ;
        RECT 86.710 172.360 87.030 172.420 ;
        RECT 77.985 172.220 87.030 172.360 ;
        RECT 77.985 172.175 78.275 172.220 ;
        RECT 86.710 172.160 87.030 172.220 ;
        RECT 87.170 172.160 87.490 172.420 ;
        RECT 18.100 171.540 89.400 172.020 ;
        RECT 21.865 171.340 22.155 171.385 ;
        RECT 22.770 171.340 23.090 171.400 ;
        RECT 21.865 171.200 23.090 171.340 ;
        RECT 21.865 171.155 22.155 171.200 ;
        RECT 22.770 171.140 23.090 171.200 ;
        RECT 23.690 171.140 24.010 171.400 ;
        RECT 29.225 171.340 29.515 171.385 ;
        RECT 30.590 171.340 30.910 171.400 ;
        RECT 29.225 171.200 30.910 171.340 ;
        RECT 29.225 171.155 29.515 171.200 ;
        RECT 30.590 171.140 30.910 171.200 ;
        RECT 31.510 171.340 31.830 171.400 ;
        RECT 35.665 171.340 35.955 171.385 ;
        RECT 31.510 171.200 35.955 171.340 ;
        RECT 31.510 171.140 31.830 171.200 ;
        RECT 35.665 171.155 35.955 171.200 ;
        RECT 38.870 171.340 39.190 171.400 ;
        RECT 39.345 171.340 39.635 171.385 ;
        RECT 38.870 171.200 39.635 171.340 ;
        RECT 38.870 171.140 39.190 171.200 ;
        RECT 39.345 171.155 39.635 171.200 ;
        RECT 44.390 171.340 44.710 171.400 ;
        RECT 44.865 171.340 45.155 171.385 ;
        RECT 44.390 171.200 45.155 171.340 ;
        RECT 44.390 171.140 44.710 171.200 ;
        RECT 44.865 171.155 45.155 171.200 ;
        RECT 46.230 171.340 46.550 171.400 ;
        RECT 46.705 171.340 46.995 171.385 ;
        RECT 56.810 171.340 57.130 171.400 ;
        RECT 46.230 171.200 46.995 171.340 ;
        RECT 46.230 171.140 46.550 171.200 ;
        RECT 46.705 171.155 46.995 171.200 ;
        RECT 48.160 171.200 57.130 171.340 ;
        RECT 27.830 171.000 28.150 171.060 ;
        RECT 45.785 171.000 46.075 171.045 ;
        RECT 27.830 170.860 33.220 171.000 ;
        RECT 27.830 170.800 28.150 170.860 ;
        RECT 28.750 170.460 29.070 170.720 ;
        RECT 29.210 170.660 29.530 170.720 ;
        RECT 30.145 170.660 30.435 170.705 ;
        RECT 29.210 170.520 30.435 170.660 ;
        RECT 29.210 170.460 29.530 170.520 ;
        RECT 30.145 170.475 30.435 170.520 ;
        RECT 31.510 170.460 31.830 170.720 ;
        RECT 32.335 170.460 32.655 170.720 ;
        RECT 33.080 170.705 33.220 170.860 ;
        RECT 38.040 170.860 46.075 171.000 ;
        RECT 32.905 170.520 33.220 170.705 ;
        RECT 32.905 170.475 33.195 170.520 ;
        RECT 34.270 170.460 34.590 170.720 ;
        RECT 34.745 170.660 35.035 170.705 ;
        RECT 37.030 170.660 37.350 170.720 ;
        RECT 34.745 170.520 37.350 170.660 ;
        RECT 34.745 170.475 35.035 170.520 ;
        RECT 37.030 170.460 37.350 170.520 ;
        RECT 24.150 170.120 24.470 170.380 ;
        RECT 24.610 170.120 24.930 170.380 ;
        RECT 38.040 170.320 38.180 170.860 ;
        RECT 45.785 170.815 46.075 170.860 ;
        RECT 38.885 170.660 39.175 170.705 ;
        RECT 41.170 170.660 41.490 170.720 ;
        RECT 38.885 170.520 41.490 170.660 ;
        RECT 38.885 170.475 39.175 170.520 ;
        RECT 41.170 170.460 41.490 170.520 ;
        RECT 43.470 170.660 43.790 170.720 ;
        RECT 44.405 170.660 44.695 170.705 ;
        RECT 43.470 170.520 44.695 170.660 ;
        RECT 43.470 170.460 43.790 170.520 ;
        RECT 44.405 170.475 44.695 170.520 ;
        RECT 47.150 170.660 47.470 170.720 ;
        RECT 47.625 170.660 47.915 170.705 ;
        RECT 47.150 170.520 47.915 170.660 ;
        RECT 47.150 170.460 47.470 170.520 ;
        RECT 47.625 170.475 47.915 170.520 ;
        RECT 30.220 170.180 38.180 170.320 ;
        RECT 39.330 170.320 39.650 170.380 ;
        RECT 39.805 170.320 40.095 170.365 ;
        RECT 39.330 170.180 40.095 170.320 ;
        RECT 30.220 170.025 30.360 170.180 ;
        RECT 39.330 170.120 39.650 170.180 ;
        RECT 39.805 170.135 40.095 170.180 ;
        RECT 40.250 170.320 40.570 170.380 ;
        RECT 46.690 170.320 47.010 170.380 ;
        RECT 40.250 170.180 47.010 170.320 ;
        RECT 40.250 170.120 40.570 170.180 ;
        RECT 46.690 170.120 47.010 170.180 ;
        RECT 30.145 169.795 30.435 170.025 ;
        RECT 33.365 169.980 33.655 170.025 ;
        RECT 37.045 169.980 37.335 170.025 ;
        RECT 33.365 169.840 37.335 169.980 ;
        RECT 33.365 169.795 33.655 169.840 ;
        RECT 37.045 169.795 37.335 169.840 ;
        RECT 45.785 169.980 46.075 170.025 ;
        RECT 48.160 169.980 48.300 171.200 ;
        RECT 56.810 171.140 57.130 171.200 ;
        RECT 57.730 171.140 58.050 171.400 ;
        RECT 58.190 171.340 58.510 171.400 ;
        RECT 64.185 171.340 64.475 171.385 ;
        RECT 68.310 171.340 68.630 171.400 ;
        RECT 58.190 171.200 64.475 171.340 ;
        RECT 58.190 171.140 58.510 171.200 ;
        RECT 64.185 171.155 64.475 171.200 ;
        RECT 65.180 171.200 68.630 171.340 ;
        RECT 48.545 171.000 48.835 171.045 ;
        RECT 52.670 171.000 52.990 171.060 ;
        RECT 48.545 170.860 52.990 171.000 ;
        RECT 48.545 170.815 48.835 170.860 ;
        RECT 52.670 170.800 52.990 170.860 ;
        RECT 53.145 171.000 53.435 171.045 ;
        RECT 54.050 171.000 54.370 171.060 ;
        RECT 53.145 170.860 54.370 171.000 ;
        RECT 53.145 170.815 53.435 170.860 ;
        RECT 54.050 170.800 54.370 170.860 ;
        RECT 54.510 171.000 54.830 171.060 ;
        RECT 54.985 171.000 55.275 171.045 ;
        RECT 54.510 170.860 55.275 171.000 ;
        RECT 54.510 170.800 54.830 170.860 ;
        RECT 54.985 170.815 55.275 170.860 ;
        RECT 48.990 170.460 49.310 170.720 ;
        RECT 52.225 170.475 52.515 170.705 ;
        RECT 52.300 170.320 52.440 170.475 ;
        RECT 53.590 170.460 53.910 170.720 ;
        RECT 55.890 170.460 56.210 170.720 ;
        RECT 56.365 170.475 56.655 170.705 ;
        RECT 56.440 170.320 56.580 170.475 ;
        RECT 58.650 170.460 58.970 170.720 ;
        RECT 60.030 170.460 60.350 170.720 ;
        RECT 60.505 170.660 60.795 170.705 ;
        RECT 60.950 170.660 61.270 170.720 ;
        RECT 60.505 170.520 61.270 170.660 ;
        RECT 60.505 170.475 60.795 170.520 ;
        RECT 60.950 170.460 61.270 170.520 ;
        RECT 62.805 170.660 63.095 170.705 ;
        RECT 63.710 170.660 64.030 170.720 ;
        RECT 65.180 170.705 65.320 171.200 ;
        RECT 68.310 171.140 68.630 171.200 ;
        RECT 69.245 171.155 69.535 171.385 ;
        RECT 71.545 171.340 71.835 171.385 ;
        RECT 82.570 171.340 82.890 171.400 ;
        RECT 71.545 171.200 82.890 171.340 ;
        RECT 71.545 171.155 71.835 171.200 ;
        RECT 68.770 171.000 69.090 171.060 ;
        RECT 65.640 170.860 69.090 171.000 ;
        RECT 69.320 171.000 69.460 171.155 ;
        RECT 82.570 171.140 82.890 171.200 ;
        RECT 83.490 171.340 83.810 171.400 ;
        RECT 85.345 171.340 85.635 171.385 ;
        RECT 83.490 171.200 85.635 171.340 ;
        RECT 83.490 171.140 83.810 171.200 ;
        RECT 85.345 171.155 85.635 171.200 ;
        RECT 71.990 171.000 72.310 171.060 ;
        RECT 77.970 171.000 78.290 171.060 ;
        RECT 69.320 170.860 72.310 171.000 ;
        RECT 65.640 170.705 65.780 170.860 ;
        RECT 68.770 170.800 69.090 170.860 ;
        RECT 71.990 170.800 72.310 170.860 ;
        RECT 73.000 170.860 78.290 171.000 ;
        RECT 62.805 170.520 64.030 170.660 ;
        RECT 62.805 170.475 63.095 170.520 ;
        RECT 63.710 170.460 64.030 170.520 ;
        RECT 65.105 170.475 65.395 170.705 ;
        RECT 65.565 170.475 65.855 170.705 ;
        RECT 67.850 170.460 68.170 170.720 ;
        RECT 68.325 170.660 68.615 170.705 ;
        RECT 69.690 170.660 70.010 170.720 ;
        RECT 68.325 170.520 70.010 170.660 ;
        RECT 68.325 170.475 68.615 170.520 ;
        RECT 69.690 170.460 70.010 170.520 ;
        RECT 70.610 170.460 70.930 170.720 ;
        RECT 73.000 170.705 73.140 170.860 ;
        RECT 77.970 170.800 78.290 170.860 ;
        RECT 72.925 170.475 73.215 170.705 ;
        RECT 73.370 170.460 73.690 170.720 ;
        RECT 73.830 170.660 74.150 170.720 ;
        RECT 74.305 170.660 74.595 170.705 ;
        RECT 73.830 170.520 74.595 170.660 ;
        RECT 73.830 170.460 74.150 170.520 ;
        RECT 74.305 170.475 74.595 170.520 ;
        RECT 75.685 170.660 75.975 170.705 ;
        RECT 76.590 170.660 76.910 170.720 ;
        RECT 75.685 170.520 76.910 170.660 ;
        RECT 75.685 170.475 75.975 170.520 ;
        RECT 76.590 170.460 76.910 170.520 ;
        RECT 77.065 170.680 77.355 170.705 ;
        RECT 77.065 170.540 77.740 170.680 ;
        RECT 77.065 170.475 77.355 170.540 ;
        RECT 59.125 170.320 59.415 170.365 ;
        RECT 52.300 170.180 55.200 170.320 ;
        RECT 56.440 170.180 59.415 170.320 ;
        RECT 45.785 169.840 48.300 169.980 ;
        RECT 48.620 169.840 51.980 169.980 ;
        RECT 45.785 169.795 46.075 169.840 ;
        RECT 34.270 169.640 34.590 169.700 ;
        RECT 37.490 169.640 37.810 169.700 ;
        RECT 34.270 169.500 37.810 169.640 ;
        RECT 34.270 169.440 34.590 169.500 ;
        RECT 37.490 169.440 37.810 169.500 ;
        RECT 39.790 169.640 40.110 169.700 ;
        RECT 46.230 169.640 46.550 169.700 ;
        RECT 39.790 169.500 46.550 169.640 ;
        RECT 39.790 169.440 40.110 169.500 ;
        RECT 46.230 169.440 46.550 169.500 ;
        RECT 46.690 169.640 47.010 169.700 ;
        RECT 48.620 169.640 48.760 169.840 ;
        RECT 46.690 169.500 48.760 169.640 ;
        RECT 51.840 169.640 51.980 169.840 ;
        RECT 52.210 169.780 52.530 170.040 ;
        RECT 55.060 170.025 55.200 170.180 ;
        RECT 59.125 170.135 59.415 170.180 ;
        RECT 61.410 170.320 61.730 170.380 ;
        RECT 62.345 170.320 62.635 170.365 ;
        RECT 77.600 170.320 77.740 170.540 ;
        RECT 78.430 170.660 78.750 170.720 ;
        RECT 78.905 170.660 79.195 170.705 ;
        RECT 78.430 170.520 79.195 170.660 ;
        RECT 78.430 170.460 78.750 170.520 ;
        RECT 78.905 170.475 79.195 170.520 ;
        RECT 61.410 170.180 62.635 170.320 ;
        RECT 61.410 170.120 61.730 170.180 ;
        RECT 62.345 170.135 62.635 170.180 ;
        RECT 63.800 170.180 77.740 170.320 ;
        RECT 54.985 169.795 55.275 170.025 ;
        RECT 61.870 169.980 62.190 170.040 ;
        RECT 63.800 170.025 63.940 170.180 ;
        RECT 55.520 169.840 62.190 169.980 ;
        RECT 55.520 169.640 55.660 169.840 ;
        RECT 61.870 169.780 62.190 169.840 ;
        RECT 63.725 169.795 64.015 170.025 ;
        RECT 64.630 169.980 64.950 170.040 ;
        RECT 66.010 169.980 66.330 170.040 ;
        RECT 64.630 169.840 66.330 169.980 ;
        RECT 64.630 169.780 64.950 169.840 ;
        RECT 66.010 169.780 66.330 169.840 ;
        RECT 66.930 169.780 67.250 170.040 ;
        RECT 75.670 169.980 75.990 170.040 ;
        RECT 67.480 169.840 75.990 169.980 ;
        RECT 51.840 169.500 55.660 169.640 ;
        RECT 66.485 169.640 66.775 169.685 ;
        RECT 67.480 169.640 67.620 169.840 ;
        RECT 75.670 169.780 75.990 169.840 ;
        RECT 76.130 169.980 76.450 170.040 ;
        RECT 76.605 169.980 76.895 170.025 ;
        RECT 76.130 169.840 76.895 169.980 ;
        RECT 76.130 169.780 76.450 169.840 ;
        RECT 76.605 169.795 76.895 169.840 ;
        RECT 77.970 169.780 78.290 170.040 ;
        RECT 66.485 169.500 67.620 169.640 ;
        RECT 46.690 169.440 47.010 169.500 ;
        RECT 66.485 169.455 66.775 169.500 ;
        RECT 18.100 168.820 89.400 169.300 ;
        RECT 21.390 168.420 21.710 168.680 ;
        RECT 33.350 168.620 33.670 168.680 ;
        RECT 26.310 168.480 33.670 168.620 ;
        RECT 23.690 167.740 24.010 168.000 ;
        RECT 24.165 167.940 24.455 167.985 ;
        RECT 24.610 167.940 24.930 168.000 ;
        RECT 26.310 167.940 26.450 168.480 ;
        RECT 33.350 168.420 33.670 168.480 ;
        RECT 35.205 168.620 35.495 168.665 ;
        RECT 35.650 168.620 35.970 168.680 ;
        RECT 35.205 168.480 35.970 168.620 ;
        RECT 35.205 168.435 35.495 168.480 ;
        RECT 35.650 168.420 35.970 168.480 ;
        RECT 36.585 168.620 36.875 168.665 ;
        RECT 37.030 168.620 37.350 168.680 ;
        RECT 36.585 168.480 37.350 168.620 ;
        RECT 36.585 168.435 36.875 168.480 ;
        RECT 37.030 168.420 37.350 168.480 ;
        RECT 37.950 168.620 38.270 168.680 ;
        RECT 43.010 168.620 43.330 168.680 ;
        RECT 46.690 168.620 47.010 168.680 ;
        RECT 37.950 168.480 47.010 168.620 ;
        RECT 37.950 168.420 38.270 168.480 ;
        RECT 43.010 168.420 43.330 168.480 ;
        RECT 46.690 168.420 47.010 168.480 ;
        RECT 48.990 168.620 49.310 168.680 ;
        RECT 49.465 168.620 49.755 168.665 ;
        RECT 48.990 168.480 49.755 168.620 ;
        RECT 48.990 168.420 49.310 168.480 ;
        RECT 49.465 168.435 49.755 168.480 ;
        RECT 58.190 168.420 58.510 168.680 ;
        RECT 65.090 168.620 65.410 168.680 ;
        RECT 75.225 168.620 75.515 168.665 ;
        RECT 65.090 168.480 75.515 168.620 ;
        RECT 65.090 168.420 65.410 168.480 ;
        RECT 75.225 168.435 75.515 168.480 ;
        RECT 29.685 168.280 29.975 168.325 ;
        RECT 31.050 168.280 31.370 168.340 ;
        RECT 29.685 168.140 31.370 168.280 ;
        RECT 29.685 168.095 29.975 168.140 ;
        RECT 31.050 168.080 31.370 168.140 ;
        RECT 31.510 168.280 31.830 168.340 ;
        RECT 31.510 168.140 40.480 168.280 ;
        RECT 31.510 168.080 31.830 168.140 ;
        RECT 24.165 167.800 26.450 167.940 ;
        RECT 24.165 167.755 24.455 167.800 ;
        RECT 23.230 167.600 23.550 167.660 ;
        RECT 24.240 167.600 24.380 167.755 ;
        RECT 24.610 167.740 24.930 167.800 ;
        RECT 38.870 167.740 39.190 168.000 ;
        RECT 39.790 167.740 40.110 168.000 ;
        RECT 23.230 167.460 24.380 167.600 ;
        RECT 28.305 167.600 28.595 167.645 ;
        RECT 29.210 167.600 29.530 167.660 ;
        RECT 28.305 167.460 29.530 167.600 ;
        RECT 23.230 167.400 23.550 167.460 ;
        RECT 28.305 167.415 28.595 167.460 ;
        RECT 29.210 167.400 29.530 167.460 ;
        RECT 29.670 167.400 29.990 167.660 ;
        RECT 31.510 167.600 31.830 167.660 ;
        RECT 32.445 167.600 32.735 167.645 ;
        RECT 31.510 167.460 32.735 167.600 ;
        RECT 31.510 167.400 31.830 167.460 ;
        RECT 32.445 167.415 32.735 167.460 ;
        RECT 33.350 167.400 33.670 167.660 ;
        RECT 33.825 167.600 34.115 167.645 ;
        RECT 35.650 167.600 35.970 167.660 ;
        RECT 33.825 167.460 35.970 167.600 ;
        RECT 33.825 167.415 34.115 167.460 ;
        RECT 35.650 167.400 35.970 167.460 ;
        RECT 40.340 167.610 40.480 168.140 ;
        RECT 40.710 168.080 41.030 168.340 ;
        RECT 42.550 168.280 42.870 168.340 ;
        RECT 45.785 168.280 46.075 168.325 ;
        RECT 50.830 168.280 51.150 168.340 ;
        RECT 42.550 168.140 43.700 168.280 ;
        RECT 42.550 168.080 42.870 168.140 ;
        RECT 40.800 167.940 40.940 168.080 ;
        RECT 40.800 167.800 42.320 167.940 ;
        RECT 42.180 167.655 42.320 167.800 ;
        RECT 40.685 167.610 40.975 167.655 ;
        RECT 40.340 167.425 40.975 167.610 ;
        RECT 42.105 167.425 42.395 167.655 ;
        RECT 40.340 167.410 40.940 167.425 ;
        RECT 29.760 167.260 29.900 167.400 ;
        RECT 32.890 167.260 33.210 167.320 ;
        RECT 35.205 167.260 35.495 167.305 ;
        RECT 29.760 167.120 35.495 167.260 ;
        RECT 32.890 167.060 33.210 167.120 ;
        RECT 35.205 167.075 35.495 167.120 ;
        RECT 21.390 166.920 21.710 166.980 ;
        RECT 23.245 166.920 23.535 166.965 ;
        RECT 24.150 166.920 24.470 166.980 ;
        RECT 21.390 166.780 24.470 166.920 ;
        RECT 21.390 166.720 21.710 166.780 ;
        RECT 23.245 166.735 23.535 166.780 ;
        RECT 24.150 166.720 24.470 166.780 ;
        RECT 28.765 166.920 29.055 166.965 ;
        RECT 31.525 166.920 31.815 166.965 ;
        RECT 34.285 166.920 34.575 166.965 ;
        RECT 28.765 166.780 34.575 166.920 ;
        RECT 28.765 166.735 29.055 166.780 ;
        RECT 31.525 166.735 31.815 166.780 ;
        RECT 34.285 166.735 34.575 166.780 ;
        RECT 37.950 166.920 38.270 166.980 ;
        RECT 38.425 166.920 38.715 166.965 ;
        RECT 37.950 166.780 38.715 166.920 ;
        RECT 40.800 166.920 40.940 167.410 ;
        RECT 43.010 167.400 43.330 167.660 ;
        RECT 41.185 167.260 41.475 167.305 ;
        RECT 43.560 167.260 43.700 168.140 ;
        RECT 45.785 168.140 51.150 168.280 ;
        RECT 45.785 168.095 46.075 168.140 ;
        RECT 50.830 168.080 51.150 168.140 ;
        RECT 53.130 168.280 53.450 168.340 ;
        RECT 66.025 168.280 66.315 168.325 ;
        RECT 53.130 168.140 66.315 168.280 ;
        RECT 53.130 168.080 53.450 168.140 ;
        RECT 66.025 168.095 66.315 168.140 ;
        RECT 66.930 168.080 67.250 168.340 ;
        RECT 71.085 168.280 71.375 168.325 ;
        RECT 69.320 168.140 71.375 168.280 ;
        RECT 43.930 167.940 44.250 168.000 ;
        RECT 61.870 167.940 62.190 168.000 ;
        RECT 63.250 167.940 63.570 168.000 ;
        RECT 43.930 167.800 49.220 167.940 ;
        RECT 43.930 167.740 44.250 167.800 ;
        RECT 44.390 167.400 44.710 167.660 ;
        RECT 44.940 167.645 45.080 167.800 ;
        RECT 44.865 167.415 45.155 167.645 ;
        RECT 46.230 167.400 46.550 167.660 ;
        RECT 49.080 167.645 49.220 167.800 ;
        RECT 61.870 167.800 64.400 167.940 ;
        RECT 61.870 167.740 62.190 167.800 ;
        RECT 63.250 167.740 63.570 167.800 ;
        RECT 49.005 167.415 49.295 167.645 ;
        RECT 49.925 167.600 50.215 167.645 ;
        RECT 50.370 167.600 50.690 167.660 ;
        RECT 58.650 167.600 58.970 167.660 ;
        RECT 49.925 167.460 50.690 167.600 ;
        RECT 49.925 167.415 50.215 167.460 ;
        RECT 50.370 167.400 50.690 167.460 ;
        RECT 50.920 167.460 58.970 167.600 ;
        RECT 45.785 167.260 46.075 167.305 ;
        RECT 41.185 167.120 42.780 167.260 ;
        RECT 43.560 167.120 46.075 167.260 ;
        RECT 41.185 167.075 41.475 167.120 ;
        RECT 42.105 166.920 42.395 166.965 ;
        RECT 40.800 166.780 42.395 166.920 ;
        RECT 42.640 166.920 42.780 167.120 ;
        RECT 45.785 167.075 46.075 167.120 ;
        RECT 45.310 166.920 45.630 166.980 ;
        RECT 42.640 166.780 45.630 166.920 ;
        RECT 46.320 166.920 46.460 167.400 ;
        RECT 46.705 167.260 46.995 167.305 ;
        RECT 47.150 167.260 47.470 167.320 ;
        RECT 50.920 167.260 51.060 167.460 ;
        RECT 58.650 167.400 58.970 167.460 ;
        RECT 60.030 167.400 60.350 167.660 ;
        RECT 64.260 167.645 64.400 167.800 ;
        RECT 63.725 167.415 64.015 167.645 ;
        RECT 64.185 167.415 64.475 167.645 ;
        RECT 46.705 167.120 51.060 167.260 ;
        RECT 53.590 167.260 53.910 167.320 ;
        RECT 62.805 167.260 63.095 167.305 ;
        RECT 53.590 167.120 63.095 167.260 ;
        RECT 63.800 167.260 63.940 167.415 ;
        RECT 65.090 167.400 65.410 167.660 ;
        RECT 65.550 167.400 65.870 167.660 ;
        RECT 67.020 167.645 67.160 168.080 ;
        RECT 66.920 167.415 67.210 167.645 ;
        RECT 67.390 167.400 67.710 167.660 ;
        RECT 68.770 167.600 69.090 167.660 ;
        RECT 69.320 167.645 69.460 168.140 ;
        RECT 71.085 168.095 71.375 168.140 ;
        RECT 73.370 168.280 73.690 168.340 ;
        RECT 73.845 168.280 74.135 168.325 ;
        RECT 77.510 168.280 77.830 168.340 ;
        RECT 73.370 168.140 77.830 168.280 ;
        RECT 73.370 168.080 73.690 168.140 ;
        RECT 73.845 168.095 74.135 168.140 ;
        RECT 77.510 168.080 77.830 168.140 ;
        RECT 78.430 168.080 78.750 168.340 ;
        RECT 70.610 167.940 70.930 168.000 ;
        RECT 83.045 167.940 83.335 167.985 ;
        RECT 84.870 167.940 85.190 168.000 ;
        RECT 70.610 167.800 83.335 167.940 ;
        RECT 70.610 167.740 70.930 167.800 ;
        RECT 83.045 167.755 83.335 167.800 ;
        RECT 84.040 167.800 85.190 167.940 ;
        RECT 68.575 167.460 69.090 167.600 ;
        RECT 68.770 167.400 69.090 167.460 ;
        RECT 69.245 167.415 69.535 167.645 ;
        RECT 69.690 167.450 70.010 167.710 ;
        RECT 71.990 167.600 72.310 167.660 ;
        RECT 72.925 167.600 73.215 167.645 ;
        RECT 71.990 167.460 73.215 167.600 ;
        RECT 71.990 167.400 72.310 167.460 ;
        RECT 72.925 167.415 73.215 167.460 ;
        RECT 73.385 167.600 73.675 167.645 ;
        RECT 73.830 167.600 74.150 167.660 ;
        RECT 73.385 167.460 74.150 167.600 ;
        RECT 73.385 167.415 73.675 167.460 ;
        RECT 73.830 167.400 74.150 167.460 ;
        RECT 74.305 167.600 74.595 167.645 ;
        RECT 74.750 167.600 75.070 167.660 ;
        RECT 74.305 167.460 75.070 167.600 ;
        RECT 74.305 167.415 74.595 167.460 ;
        RECT 74.750 167.400 75.070 167.460 ;
        RECT 76.590 167.600 76.910 167.660 ;
        RECT 84.040 167.645 84.180 167.800 ;
        RECT 84.870 167.740 85.190 167.800 ;
        RECT 76.590 167.460 81.420 167.600 ;
        RECT 76.590 167.400 76.910 167.460 ;
        RECT 67.865 167.260 68.155 167.305 ;
        RECT 63.800 167.120 70.840 167.260 ;
        RECT 46.705 167.075 46.995 167.120 ;
        RECT 47.150 167.060 47.470 167.120 ;
        RECT 53.590 167.060 53.910 167.120 ;
        RECT 62.805 167.075 63.095 167.120 ;
        RECT 67.865 167.075 68.155 167.120 ;
        RECT 53.130 166.920 53.450 166.980 ;
        RECT 46.320 166.780 53.450 166.920 ;
        RECT 37.950 166.720 38.270 166.780 ;
        RECT 38.425 166.735 38.715 166.780 ;
        RECT 42.105 166.735 42.395 166.780 ;
        RECT 45.310 166.720 45.630 166.780 ;
        RECT 53.130 166.720 53.450 166.780 ;
        RECT 54.970 166.920 55.290 166.980 ;
        RECT 57.285 166.920 57.575 166.965 ;
        RECT 54.970 166.780 57.575 166.920 ;
        RECT 54.970 166.720 55.290 166.780 ;
        RECT 57.285 166.735 57.575 166.780 ;
        RECT 66.930 166.920 67.250 166.980 ;
        RECT 70.165 166.920 70.455 166.965 ;
        RECT 66.930 166.780 70.455 166.920 ;
        RECT 70.700 166.920 70.840 167.120 ;
        RECT 71.070 167.060 71.390 167.320 ;
        RECT 77.525 167.260 77.815 167.305 ;
        RECT 77.970 167.260 78.290 167.320 ;
        RECT 77.525 167.120 78.290 167.260 ;
        RECT 77.525 167.075 77.815 167.120 ;
        RECT 77.970 167.060 78.290 167.120 ;
        RECT 80.270 167.260 80.590 167.320 ;
        RECT 80.745 167.260 81.035 167.305 ;
        RECT 80.270 167.120 81.035 167.260 ;
        RECT 81.280 167.260 81.420 167.460 ;
        RECT 83.965 167.415 84.255 167.645 ;
        RECT 84.410 167.400 84.730 167.660 ;
        RECT 85.805 167.260 86.095 167.305 ;
        RECT 81.280 167.120 86.095 167.260 ;
        RECT 80.270 167.060 80.590 167.120 ;
        RECT 80.745 167.075 81.035 167.120 ;
        RECT 85.805 167.075 86.095 167.120 ;
        RECT 75.670 166.920 75.990 166.980 ;
        RECT 70.700 166.780 75.990 166.920 ;
        RECT 66.930 166.720 67.250 166.780 ;
        RECT 70.165 166.735 70.455 166.780 ;
        RECT 75.670 166.720 75.990 166.780 ;
        RECT 18.100 166.100 89.400 166.580 ;
        RECT 22.310 165.900 22.630 165.960 ;
        RECT 23.705 165.900 23.995 165.945 ;
        RECT 22.310 165.760 23.995 165.900 ;
        RECT 22.310 165.700 22.630 165.760 ;
        RECT 23.705 165.715 23.995 165.760 ;
        RECT 29.210 165.700 29.530 165.960 ;
        RECT 33.350 165.900 33.670 165.960 ;
        RECT 39.790 165.900 40.110 165.960 ;
        RECT 33.350 165.760 40.110 165.900 ;
        RECT 33.350 165.700 33.670 165.760 ;
        RECT 39.790 165.700 40.110 165.760 ;
        RECT 47.610 165.700 47.930 165.960 ;
        RECT 48.530 165.700 48.850 165.960 ;
        RECT 52.670 165.900 52.990 165.960 ;
        RECT 53.145 165.900 53.435 165.945 ;
        RECT 55.430 165.900 55.750 165.960 ;
        RECT 61.885 165.900 62.175 165.945 ;
        RECT 68.310 165.900 68.630 165.960 ;
        RECT 52.670 165.760 53.435 165.900 ;
        RECT 52.670 165.700 52.990 165.760 ;
        RECT 53.145 165.715 53.435 165.760 ;
        RECT 54.140 165.760 62.175 165.900 ;
        RECT 38.870 165.560 39.190 165.620 ;
        RECT 26.540 165.420 39.190 165.560 ;
        RECT 23.690 165.220 24.010 165.280 ;
        RECT 26.540 165.265 26.680 165.420 ;
        RECT 38.870 165.360 39.190 165.420 ;
        RECT 24.165 165.220 24.455 165.265 ;
        RECT 23.690 165.080 24.455 165.220 ;
        RECT 23.690 165.020 24.010 165.080 ;
        RECT 24.165 165.035 24.455 165.080 ;
        RECT 26.465 165.035 26.755 165.265 ;
        RECT 27.830 165.020 28.150 165.280 ;
        RECT 28.290 165.020 28.610 165.280 ;
        RECT 43.930 165.220 44.250 165.280 ;
        RECT 54.140 165.265 54.280 165.760 ;
        RECT 55.430 165.700 55.750 165.760 ;
        RECT 61.885 165.715 62.175 165.760 ;
        RECT 66.560 165.760 68.630 165.900 ;
        RECT 54.510 165.560 54.830 165.620 ;
        RECT 60.950 165.560 61.270 165.620 ;
        RECT 66.560 165.605 66.700 165.760 ;
        RECT 68.310 165.700 68.630 165.760 ;
        RECT 69.245 165.900 69.535 165.945 ;
        RECT 83.950 165.900 84.270 165.960 ;
        RECT 69.245 165.760 84.270 165.900 ;
        RECT 69.245 165.715 69.535 165.760 ;
        RECT 83.950 165.700 84.270 165.760 ;
        RECT 84.885 165.900 85.175 165.945 ;
        RECT 86.250 165.900 86.570 165.960 ;
        RECT 84.885 165.760 86.570 165.900 ;
        RECT 84.885 165.715 85.175 165.760 ;
        RECT 86.250 165.700 86.570 165.760 ;
        RECT 54.510 165.420 55.660 165.560 ;
        RECT 54.510 165.360 54.830 165.420 ;
        RECT 48.250 165.220 48.540 165.265 ;
        RECT 43.930 165.080 48.540 165.220 ;
        RECT 43.930 165.020 44.250 165.080 ;
        RECT 48.250 165.035 48.540 165.080 ;
        RECT 54.065 165.035 54.355 165.265 ;
        RECT 54.970 165.020 55.290 165.280 ;
        RECT 55.520 165.265 55.660 165.420 ;
        RECT 57.820 165.420 59.340 165.560 ;
        RECT 55.445 165.035 55.735 165.265 ;
        RECT 55.890 165.220 56.210 165.280 ;
        RECT 56.365 165.220 56.655 165.265 ;
        RECT 55.890 165.080 56.655 165.220 ;
        RECT 55.890 165.020 56.210 165.080 ;
        RECT 56.365 165.035 56.655 165.080 ;
        RECT 57.270 165.020 57.590 165.280 ;
        RECT 57.820 165.265 57.960 165.420 ;
        RECT 59.200 165.280 59.340 165.420 ;
        RECT 60.950 165.420 63.480 165.560 ;
        RECT 60.950 165.360 61.270 165.420 ;
        RECT 57.745 165.035 58.035 165.265 ;
        RECT 58.190 165.020 58.510 165.280 ;
        RECT 59.110 165.220 59.430 165.280 ;
        RECT 60.045 165.220 60.335 165.265 ;
        RECT 59.110 165.080 60.335 165.220 ;
        RECT 59.110 165.020 59.430 165.080 ;
        RECT 60.045 165.035 60.335 165.080 ;
        RECT 60.490 165.220 60.810 165.280 ;
        RECT 63.340 165.265 63.480 165.420 ;
        RECT 66.485 165.375 66.775 165.605 ;
        RECT 66.930 165.560 67.250 165.620 ;
        RECT 67.405 165.560 67.695 165.605 ;
        RECT 66.930 165.420 67.695 165.560 ;
        RECT 66.930 165.360 67.250 165.420 ;
        RECT 67.405 165.375 67.695 165.420 ;
        RECT 70.150 165.560 70.470 165.620 ;
        RECT 73.370 165.560 73.690 165.620 ;
        RECT 77.970 165.560 78.290 165.620 ;
        RECT 85.805 165.560 86.095 165.605 ;
        RECT 87.630 165.560 87.950 165.620 ;
        RECT 70.150 165.420 72.680 165.560 ;
        RECT 62.345 165.220 62.635 165.265 ;
        RECT 60.490 165.080 62.635 165.220 ;
        RECT 60.490 165.020 60.810 165.080 ;
        RECT 62.345 165.035 62.635 165.080 ;
        RECT 63.265 165.035 63.555 165.265 ;
        RECT 67.845 165.145 68.135 165.375 ;
        RECT 70.150 165.360 70.470 165.420 ;
        RECT 23.230 164.680 23.550 164.940 ;
        RECT 32.890 164.880 33.210 164.940 ;
        RECT 50.845 164.880 51.135 164.925 ;
        RECT 53.590 164.880 53.910 164.940 ;
        RECT 32.890 164.740 53.910 164.880 ;
        RECT 32.890 164.680 33.210 164.740 ;
        RECT 50.845 164.695 51.135 164.740 ;
        RECT 53.590 164.680 53.910 164.740 ;
        RECT 54.525 164.880 54.815 164.925 ;
        RECT 56.810 164.880 57.130 164.940 ;
        RECT 54.525 164.740 57.130 164.880 ;
        RECT 58.280 164.880 58.420 165.020 ;
        RECT 67.940 164.940 68.080 165.145 ;
        RECT 68.325 165.035 68.615 165.265 ;
        RECT 71.085 165.220 71.375 165.265 ;
        RECT 71.990 165.220 72.310 165.280 ;
        RECT 72.540 165.265 72.680 165.420 ;
        RECT 73.370 165.420 77.740 165.560 ;
        RECT 73.370 165.360 73.690 165.420 ;
        RECT 71.085 165.080 72.310 165.220 ;
        RECT 71.085 165.035 71.375 165.080 ;
        RECT 62.805 164.880 63.095 164.925 ;
        RECT 58.280 164.740 63.095 164.880 ;
        RECT 54.525 164.695 54.815 164.740 ;
        RECT 56.810 164.680 57.130 164.740 ;
        RECT 62.805 164.695 63.095 164.740 ;
        RECT 67.850 164.680 68.170 164.940 ;
        RECT 68.400 164.880 68.540 165.035 ;
        RECT 71.990 165.020 72.310 165.080 ;
        RECT 72.465 165.035 72.755 165.265 ;
        RECT 73.845 165.220 74.135 165.265 ;
        RECT 74.290 165.220 74.610 165.280 ;
        RECT 73.845 165.080 74.610 165.220 ;
        RECT 73.845 165.035 74.135 165.080 ;
        RECT 74.290 165.020 74.610 165.080 ;
        RECT 74.765 165.220 75.055 165.265 ;
        RECT 75.210 165.220 75.530 165.280 ;
        RECT 74.765 165.080 75.530 165.220 ;
        RECT 74.765 165.035 75.055 165.080 ;
        RECT 75.210 165.020 75.530 165.080 ;
        RECT 76.130 165.020 76.450 165.280 ;
        RECT 76.590 165.220 76.910 165.280 ;
        RECT 77.600 165.265 77.740 165.420 ;
        RECT 77.970 165.420 87.950 165.560 ;
        RECT 77.970 165.360 78.290 165.420 ;
        RECT 85.805 165.375 86.095 165.420 ;
        RECT 87.630 165.360 87.950 165.420 ;
        RECT 77.065 165.220 77.355 165.265 ;
        RECT 76.590 165.080 77.355 165.220 ;
        RECT 76.590 165.020 76.910 165.080 ;
        RECT 77.065 165.035 77.355 165.080 ;
        RECT 77.525 165.035 77.815 165.265 ;
        RECT 78.430 165.020 78.750 165.280 ;
        RECT 86.265 165.220 86.555 165.265 ;
        RECT 82.200 165.080 86.555 165.220 ;
        RECT 82.200 164.940 82.340 165.080 ;
        RECT 86.265 165.035 86.555 165.080 ;
        RECT 80.270 164.880 80.590 164.940 ;
        RECT 68.400 164.740 80.590 164.880 ;
        RECT 80.270 164.680 80.590 164.740 ;
        RECT 80.730 164.680 81.050 164.940 ;
        RECT 82.110 164.680 82.430 164.940 ;
        RECT 83.030 164.880 83.350 164.940 ;
        RECT 84.410 164.880 84.730 164.940 ;
        RECT 83.030 164.740 84.730 164.880 ;
        RECT 83.030 164.680 83.350 164.740 ;
        RECT 84.410 164.680 84.730 164.740 ;
        RECT 50.385 164.540 50.675 164.585 ;
        RECT 59.585 164.540 59.875 164.585 ;
        RECT 50.385 164.400 59.875 164.540 ;
        RECT 50.385 164.355 50.675 164.400 ;
        RECT 59.585 164.355 59.875 164.400 ;
        RECT 65.550 164.540 65.870 164.600 ;
        RECT 66.485 164.540 66.775 164.585 ;
        RECT 65.550 164.400 66.775 164.540 ;
        RECT 67.940 164.540 68.080 164.680 ;
        RECT 69.690 164.540 70.010 164.600 ;
        RECT 67.940 164.400 70.010 164.540 ;
        RECT 65.550 164.340 65.870 164.400 ;
        RECT 66.485 164.355 66.775 164.400 ;
        RECT 69.690 164.340 70.010 164.400 ;
        RECT 71.990 164.340 72.310 164.600 ;
        RECT 72.910 164.540 73.230 164.600 ;
        RECT 73.385 164.540 73.675 164.585 ;
        RECT 72.910 164.400 73.675 164.540 ;
        RECT 72.910 164.340 73.230 164.400 ;
        RECT 73.385 164.355 73.675 164.400 ;
        RECT 74.750 164.540 75.070 164.600 ;
        RECT 78.430 164.540 78.750 164.600 ;
        RECT 74.750 164.400 78.750 164.540 ;
        RECT 74.750 164.340 75.070 164.400 ;
        RECT 78.430 164.340 78.750 164.400 ;
        RECT 79.350 164.340 79.670 164.600 ;
        RECT 82.585 164.540 82.875 164.585 ;
        RECT 85.330 164.540 85.650 164.600 ;
        RECT 87.185 164.540 87.475 164.585 ;
        RECT 82.585 164.400 87.475 164.540 ;
        RECT 82.585 164.355 82.875 164.400 ;
        RECT 85.330 164.340 85.650 164.400 ;
        RECT 87.185 164.355 87.475 164.400 ;
        RECT 26.005 164.200 26.295 164.245 ;
        RECT 26.925 164.200 27.215 164.245 ;
        RECT 26.005 164.060 27.215 164.200 ;
        RECT 26.005 164.015 26.295 164.060 ;
        RECT 26.925 164.015 27.215 164.060 ;
        RECT 30.130 164.200 30.450 164.260 ;
        RECT 50.830 164.200 51.150 164.260 ;
        RECT 30.130 164.060 51.150 164.200 ;
        RECT 30.130 164.000 30.450 164.060 ;
        RECT 50.830 164.000 51.150 164.060 ;
        RECT 75.210 164.200 75.530 164.260 ;
        RECT 77.510 164.200 77.830 164.260 ;
        RECT 75.210 164.060 77.830 164.200 ;
        RECT 75.210 164.000 75.530 164.060 ;
        RECT 77.510 164.000 77.830 164.060 ;
        RECT 81.650 164.200 81.970 164.260 ;
        RECT 83.030 164.200 83.350 164.260 ;
        RECT 81.650 164.060 83.350 164.200 ;
        RECT 81.650 164.000 81.970 164.060 ;
        RECT 83.030 164.000 83.350 164.060 ;
        RECT 83.950 164.000 84.270 164.260 ;
        RECT 84.410 164.200 84.730 164.260 ;
        RECT 84.885 164.200 85.175 164.245 ;
        RECT 86.710 164.200 87.030 164.260 ;
        RECT 84.410 164.060 87.030 164.200 ;
        RECT 84.410 164.000 84.730 164.060 ;
        RECT 84.885 164.015 85.175 164.060 ;
        RECT 86.710 164.000 87.030 164.060 ;
        RECT 18.100 163.380 89.400 163.860 ;
        RECT 27.830 163.180 28.150 163.240 ;
        RECT 30.145 163.180 30.435 163.225 ;
        RECT 27.830 163.040 30.435 163.180 ;
        RECT 27.830 162.980 28.150 163.040 ;
        RECT 30.145 162.995 30.435 163.040 ;
        RECT 34.285 163.180 34.575 163.225 ;
        RECT 35.650 163.180 35.970 163.240 ;
        RECT 34.285 163.040 35.970 163.180 ;
        RECT 34.285 162.995 34.575 163.040 ;
        RECT 23.230 162.300 23.550 162.560 ;
        RECT 30.220 162.500 30.360 162.995 ;
        RECT 35.650 162.980 35.970 163.040 ;
        RECT 43.470 162.980 43.790 163.240 ;
        RECT 45.310 163.180 45.630 163.240 ;
        RECT 47.610 163.180 47.930 163.240 ;
        RECT 45.310 163.040 47.930 163.180 ;
        RECT 45.310 162.980 45.630 163.040 ;
        RECT 47.610 162.980 47.930 163.040 ;
        RECT 55.890 163.180 56.210 163.240 ;
        RECT 57.285 163.180 57.575 163.225 ;
        RECT 55.890 163.040 57.575 163.180 ;
        RECT 55.890 162.980 56.210 163.040 ;
        RECT 57.285 162.995 57.575 163.040 ;
        RECT 59.585 163.180 59.875 163.225 ;
        RECT 60.490 163.180 60.810 163.240 ;
        RECT 59.585 163.040 60.810 163.180 ;
        RECT 59.585 162.995 59.875 163.040 ;
        RECT 60.490 162.980 60.810 163.040 ;
        RECT 71.545 163.180 71.835 163.225 ;
        RECT 72.450 163.180 72.770 163.240 ;
        RECT 71.545 163.040 72.770 163.180 ;
        RECT 71.545 162.995 71.835 163.040 ;
        RECT 72.450 162.980 72.770 163.040 ;
        RECT 72.910 163.180 73.230 163.240 ;
        RECT 74.750 163.180 75.070 163.240 ;
        RECT 75.225 163.180 75.515 163.225 ;
        RECT 72.910 163.040 74.520 163.180 ;
        RECT 72.910 162.980 73.230 163.040 ;
        RECT 35.205 162.655 35.495 162.885 ;
        RECT 31.985 162.500 32.275 162.545 ;
        RECT 35.280 162.500 35.420 162.655 ;
        RECT 30.220 162.360 31.740 162.500 ;
        RECT 22.310 162.160 22.630 162.220 ;
        RECT 24.165 162.160 24.455 162.205 ;
        RECT 22.310 162.020 24.455 162.160 ;
        RECT 22.310 161.960 22.630 162.020 ;
        RECT 24.165 161.975 24.455 162.020 ;
        RECT 29.685 161.975 29.975 162.205 ;
        RECT 29.760 161.820 29.900 161.975 ;
        RECT 30.590 161.960 30.910 162.220 ;
        RECT 31.600 162.205 31.740 162.360 ;
        RECT 31.985 162.360 35.420 162.500 ;
        RECT 38.425 162.500 38.715 162.545 ;
        RECT 38.870 162.500 39.190 162.560 ;
        RECT 38.425 162.360 39.190 162.500 ;
        RECT 31.985 162.315 32.275 162.360 ;
        RECT 38.425 162.315 38.715 162.360 ;
        RECT 38.870 162.300 39.190 162.360 ;
        RECT 42.550 162.500 42.870 162.560 ;
        RECT 48.990 162.500 49.310 162.560 ;
        RECT 42.550 162.360 49.310 162.500 ;
        RECT 42.550 162.300 42.870 162.360 ;
        RECT 31.525 161.975 31.815 162.205 ;
        RECT 32.905 161.975 33.195 162.205 ;
        RECT 33.365 162.160 33.655 162.205 ;
        RECT 34.730 162.160 35.050 162.220 ;
        RECT 33.365 162.020 35.050 162.160 ;
        RECT 33.365 161.975 33.655 162.020 ;
        RECT 31.970 161.820 32.290 161.880 ;
        RECT 29.760 161.680 32.290 161.820 ;
        RECT 32.980 161.820 33.120 161.975 ;
        RECT 34.730 161.960 35.050 162.020 ;
        RECT 35.650 162.160 35.970 162.220 ;
        RECT 39.345 162.160 39.635 162.205 ;
        RECT 35.650 162.020 39.635 162.160 ;
        RECT 35.650 161.960 35.970 162.020 ;
        RECT 39.345 161.975 39.635 162.020 ;
        RECT 40.250 161.960 40.570 162.220 ;
        RECT 44.940 162.205 45.080 162.360 ;
        RECT 48.990 162.300 49.310 162.360 ;
        RECT 58.650 162.300 58.970 162.560 ;
        RECT 66.010 162.500 66.330 162.560 ;
        RECT 59.660 162.360 66.330 162.500 ;
        RECT 44.405 161.975 44.695 162.205 ;
        RECT 44.865 161.975 45.155 162.205 ;
        RECT 38.410 161.820 38.730 161.880 ;
        RECT 32.980 161.680 38.730 161.820 ;
        RECT 44.480 161.820 44.620 161.975 ;
        RECT 45.770 161.960 46.090 162.220 ;
        RECT 46.245 162.160 46.535 162.205 ;
        RECT 51.750 162.160 52.070 162.220 ;
        RECT 46.245 162.020 52.070 162.160 ;
        RECT 46.245 161.975 46.535 162.020 ;
        RECT 51.750 161.960 52.070 162.020 ;
        RECT 54.050 162.160 54.370 162.220 ;
        RECT 59.660 162.160 59.800 162.360 ;
        RECT 66.010 162.300 66.330 162.360 ;
        RECT 54.050 162.020 59.800 162.160 ;
        RECT 54.050 161.960 54.370 162.020 ;
        RECT 60.030 161.960 60.350 162.220 ;
        RECT 74.380 162.205 74.520 163.040 ;
        RECT 74.750 163.040 75.515 163.180 ;
        RECT 74.750 162.980 75.070 163.040 ;
        RECT 75.225 162.995 75.515 163.040 ;
        RECT 76.130 163.180 76.450 163.240 ;
        RECT 77.510 163.180 77.830 163.240 ;
        RECT 76.130 163.040 77.830 163.180 ;
        RECT 76.130 162.980 76.450 163.040 ;
        RECT 77.510 162.980 77.830 163.040 ;
        RECT 75.670 162.840 75.990 162.900 ;
        RECT 79.365 162.840 79.655 162.885 ;
        RECT 75.670 162.700 79.655 162.840 ;
        RECT 75.670 162.640 75.990 162.700 ;
        RECT 79.365 162.655 79.655 162.700 ;
        RECT 76.590 162.500 76.910 162.560 ;
        RECT 77.985 162.500 78.275 162.545 ;
        RECT 76.590 162.360 78.275 162.500 ;
        RECT 76.590 162.300 76.910 162.360 ;
        RECT 77.985 162.315 78.275 162.360 ;
        RECT 80.270 162.300 80.590 162.560 ;
        RECT 81.280 162.360 85.560 162.500 ;
        RECT 74.305 161.975 74.595 162.205 ;
        RECT 74.750 162.160 75.070 162.220 ;
        RECT 75.225 162.160 75.515 162.205 ;
        RECT 74.750 162.020 75.515 162.160 ;
        RECT 74.750 161.960 75.070 162.020 ;
        RECT 75.225 161.975 75.515 162.020 ;
        RECT 76.130 161.960 76.450 162.220 ;
        RECT 54.970 161.820 55.290 161.880 ;
        RECT 44.480 161.680 63.940 161.820 ;
        RECT 31.970 161.620 32.290 161.680 ;
        RECT 38.410 161.620 38.730 161.680 ;
        RECT 54.970 161.620 55.290 161.680 ;
        RECT 63.800 161.540 63.940 161.680 ;
        RECT 71.990 161.620 72.310 161.880 ;
        RECT 76.680 161.820 76.820 162.300 ;
        RECT 77.525 162.160 77.815 162.205 ;
        RECT 78.890 162.160 79.210 162.220 ;
        RECT 81.280 162.205 81.420 162.360 ;
        RECT 85.420 162.220 85.560 162.360 ;
        RECT 77.525 162.020 79.210 162.160 ;
        RECT 77.525 161.975 77.815 162.020 ;
        RECT 78.890 161.960 79.210 162.020 ;
        RECT 81.205 161.975 81.495 162.205 ;
        RECT 82.125 162.160 82.415 162.205 ;
        RECT 82.570 162.160 82.890 162.220 ;
        RECT 82.125 162.020 82.890 162.160 ;
        RECT 82.125 161.975 82.415 162.020 ;
        RECT 82.570 161.960 82.890 162.020 ;
        RECT 83.045 162.160 83.335 162.205 ;
        RECT 84.870 162.160 85.190 162.220 ;
        RECT 83.045 162.020 85.190 162.160 ;
        RECT 83.045 161.975 83.335 162.020 ;
        RECT 84.870 161.960 85.190 162.020 ;
        RECT 85.330 161.960 85.650 162.220 ;
        RECT 86.265 162.160 86.555 162.205 ;
        RECT 86.710 162.160 87.030 162.220 ;
        RECT 86.265 162.020 87.030 162.160 ;
        RECT 86.265 161.975 86.555 162.020 ;
        RECT 86.710 161.960 87.030 162.020 ;
        RECT 87.185 161.975 87.475 162.205 ;
        RECT 73.920 161.680 76.820 161.820 ;
        RECT 80.730 161.820 81.050 161.880 ;
        RECT 87.260 161.820 87.400 161.975 ;
        RECT 80.730 161.680 87.400 161.820 ;
        RECT 23.690 161.280 24.010 161.540 ;
        RECT 26.005 161.480 26.295 161.525 ;
        RECT 28.290 161.480 28.610 161.540 ;
        RECT 26.005 161.340 28.610 161.480 ;
        RECT 26.005 161.295 26.295 161.340 ;
        RECT 28.290 161.280 28.610 161.340 ;
        RECT 36.110 161.480 36.430 161.540 ;
        RECT 37.045 161.480 37.335 161.525 ;
        RECT 36.110 161.340 37.335 161.480 ;
        RECT 36.110 161.280 36.430 161.340 ;
        RECT 37.045 161.295 37.335 161.340 ;
        RECT 37.505 161.480 37.795 161.525 ;
        RECT 38.870 161.480 39.190 161.540 ;
        RECT 39.345 161.480 39.635 161.525 ;
        RECT 37.505 161.340 39.635 161.480 ;
        RECT 37.505 161.295 37.795 161.340 ;
        RECT 38.870 161.280 39.190 161.340 ;
        RECT 39.345 161.295 39.635 161.340 ;
        RECT 49.910 161.480 50.230 161.540 ;
        RECT 52.210 161.480 52.530 161.540 ;
        RECT 53.590 161.480 53.910 161.540 ;
        RECT 63.250 161.480 63.570 161.540 ;
        RECT 49.910 161.340 63.570 161.480 ;
        RECT 49.910 161.280 50.230 161.340 ;
        RECT 52.210 161.280 52.530 161.340 ;
        RECT 53.590 161.280 53.910 161.340 ;
        RECT 63.250 161.280 63.570 161.340 ;
        RECT 63.710 161.480 64.030 161.540 ;
        RECT 73.920 161.525 74.060 161.680 ;
        RECT 80.730 161.620 81.050 161.680 ;
        RECT 73.005 161.480 73.295 161.525 ;
        RECT 63.710 161.340 73.295 161.480 ;
        RECT 63.710 161.280 64.030 161.340 ;
        RECT 73.005 161.295 73.295 161.340 ;
        RECT 73.845 161.295 74.135 161.525 ;
        RECT 77.050 161.280 77.370 161.540 ;
        RECT 81.190 161.480 81.510 161.540 ;
        RECT 84.885 161.480 85.175 161.525 ;
        RECT 81.190 161.340 85.175 161.480 ;
        RECT 81.190 161.280 81.510 161.340 ;
        RECT 84.885 161.295 85.175 161.340 ;
        RECT 18.100 160.660 89.400 161.140 ;
        RECT 22.770 160.460 23.090 160.520 ;
        RECT 24.610 160.460 24.930 160.520 ;
        RECT 22.770 160.320 34.500 160.460 ;
        RECT 22.770 160.260 23.090 160.320 ;
        RECT 24.610 160.260 24.930 160.320 ;
        RECT 30.590 160.120 30.910 160.180 ;
        RECT 34.360 160.120 34.500 160.320 ;
        RECT 34.730 160.260 35.050 160.520 ;
        RECT 37.045 160.460 37.335 160.505 ;
        RECT 38.870 160.460 39.190 160.520 ;
        RECT 37.045 160.320 39.190 160.460 ;
        RECT 37.045 160.275 37.335 160.320 ;
        RECT 38.870 160.260 39.190 160.320 ;
        RECT 44.405 160.460 44.695 160.505 ;
        RECT 45.770 160.460 46.090 160.520 ;
        RECT 44.405 160.320 46.090 160.460 ;
        RECT 44.405 160.275 44.695 160.320 ;
        RECT 45.770 160.260 46.090 160.320 ;
        RECT 46.230 160.460 46.550 160.520 ;
        RECT 46.230 160.320 50.600 160.460 ;
        RECT 46.230 160.260 46.550 160.320 ;
        RECT 39.790 160.120 40.110 160.180 ;
        RECT 40.725 160.120 41.015 160.165 ;
        RECT 47.610 160.120 47.930 160.180 ;
        RECT 30.590 159.980 33.120 160.120 ;
        RECT 34.360 159.980 39.560 160.120 ;
        RECT 30.590 159.920 30.910 159.980 ;
        RECT 20.945 159.595 21.235 159.825 ;
        RECT 21.020 159.440 21.160 159.595 ;
        RECT 21.850 159.580 22.170 159.840 ;
        RECT 31.140 159.825 31.280 159.980 ;
        RECT 24.165 159.780 24.455 159.825 ;
        RECT 31.065 159.780 31.355 159.825 ;
        RECT 24.165 159.640 31.355 159.780 ;
        RECT 24.165 159.595 24.455 159.640 ;
        RECT 31.065 159.595 31.355 159.640 ;
        RECT 31.510 159.580 31.830 159.840 ;
        RECT 31.970 159.780 32.290 159.840 ;
        RECT 32.980 159.825 33.120 159.980 ;
        RECT 32.445 159.780 32.735 159.825 ;
        RECT 31.970 159.640 32.735 159.780 ;
        RECT 31.970 159.580 32.290 159.640 ;
        RECT 32.445 159.595 32.735 159.640 ;
        RECT 32.905 159.595 33.195 159.825 ;
        RECT 36.110 159.780 36.430 159.840 ;
        RECT 36.585 159.780 36.875 159.825 ;
        RECT 38.410 159.780 38.730 159.840 ;
        RECT 36.110 159.640 38.730 159.780 ;
        RECT 39.420 159.780 39.560 159.980 ;
        RECT 39.790 159.980 46.920 160.120 ;
        RECT 39.790 159.920 40.110 159.980 ;
        RECT 40.725 159.935 41.015 159.980 ;
        RECT 41.645 159.780 41.935 159.825 ;
        RECT 42.550 159.780 42.870 159.840 ;
        RECT 39.420 159.640 41.400 159.780 ;
        RECT 32.520 159.440 32.660 159.595 ;
        RECT 36.110 159.580 36.430 159.640 ;
        RECT 36.585 159.595 36.875 159.640 ;
        RECT 38.410 159.580 38.730 159.640 ;
        RECT 37.965 159.440 38.255 159.485 ;
        RECT 38.870 159.440 39.190 159.500 ;
        RECT 40.250 159.440 40.570 159.500 ;
        RECT 21.020 159.300 23.460 159.440 ;
        RECT 32.520 159.300 34.500 159.440 ;
        RECT 20.010 158.900 20.330 159.160 ;
        RECT 23.320 159.145 23.460 159.300 ;
        RECT 23.245 158.915 23.535 159.145 ;
        RECT 34.360 159.100 34.500 159.300 ;
        RECT 37.965 159.300 40.570 159.440 ;
        RECT 41.260 159.440 41.400 159.640 ;
        RECT 41.645 159.640 42.870 159.780 ;
        RECT 41.645 159.595 41.935 159.640 ;
        RECT 42.550 159.580 42.870 159.640 ;
        RECT 43.010 159.780 43.330 159.840 ;
        RECT 46.780 159.825 46.920 159.980 ;
        RECT 47.610 159.980 48.760 160.120 ;
        RECT 47.610 159.920 47.930 159.980 ;
        RECT 45.325 159.780 45.615 159.825 ;
        RECT 43.010 159.640 45.615 159.780 ;
        RECT 43.010 159.580 43.330 159.640 ;
        RECT 45.325 159.595 45.615 159.640 ;
        RECT 46.705 159.595 46.995 159.825 ;
        RECT 47.150 159.580 47.470 159.840 ;
        RECT 48.070 159.780 48.390 159.840 ;
        RECT 48.620 159.825 48.760 159.980 ;
        RECT 49.910 159.920 50.230 160.180 ;
        RECT 50.460 160.165 50.600 160.320 ;
        RECT 51.750 160.260 52.070 160.520 ;
        RECT 52.760 160.320 54.740 160.460 ;
        RECT 50.385 160.120 50.675 160.165 ;
        RECT 52.760 160.120 52.900 160.320 ;
        RECT 50.385 159.980 52.900 160.120 ;
        RECT 50.385 159.935 50.675 159.980 ;
        RECT 53.130 159.920 53.450 160.180 ;
        RECT 53.590 159.920 53.910 160.180 ;
        RECT 54.600 160.120 54.740 160.320 ;
        RECT 54.970 160.260 55.290 160.520 ;
        RECT 56.350 160.460 56.670 160.520 ;
        RECT 63.250 160.460 63.570 160.520 ;
        RECT 66.025 160.460 66.315 160.505 ;
        RECT 56.350 160.320 63.020 160.460 ;
        RECT 56.350 160.260 56.670 160.320 ;
        RECT 60.490 160.120 60.810 160.180 ;
        RECT 62.880 160.120 63.020 160.320 ;
        RECT 63.250 160.320 66.315 160.460 ;
        RECT 63.250 160.260 63.570 160.320 ;
        RECT 66.025 160.275 66.315 160.320 ;
        RECT 67.850 160.460 68.170 160.520 ;
        RECT 70.165 160.460 70.455 160.505 ;
        RECT 67.850 160.320 70.455 160.460 ;
        RECT 67.850 160.260 68.170 160.320 ;
        RECT 70.165 160.275 70.455 160.320 ;
        RECT 75.210 160.260 75.530 160.520 ;
        RECT 77.510 160.260 77.830 160.520 ;
        RECT 85.330 160.260 85.650 160.520 ;
        RECT 64.630 160.120 64.950 160.180 ;
        RECT 71.990 160.120 72.310 160.180 ;
        RECT 73.370 160.120 73.690 160.180 ;
        RECT 54.600 159.980 60.810 160.120 ;
        RECT 60.490 159.920 60.810 159.980 ;
        RECT 61.040 159.980 62.560 160.120 ;
        RECT 62.880 159.980 64.400 160.120 ;
        RECT 47.700 159.640 48.390 159.780 ;
        RECT 45.770 159.440 46.090 159.500 ;
        RECT 46.245 159.440 46.535 159.485 ;
        RECT 47.700 159.440 47.840 159.640 ;
        RECT 48.070 159.580 48.390 159.640 ;
        RECT 48.545 159.595 48.835 159.825 ;
        RECT 49.235 159.595 49.525 159.825 ;
        RECT 50.845 159.780 51.135 159.825 ;
        RECT 52.225 159.780 52.515 159.825 ;
        RECT 50.845 159.640 52.515 159.780 ;
        RECT 50.845 159.595 51.135 159.640 ;
        RECT 52.225 159.595 52.515 159.640 ;
        RECT 54.065 159.780 54.355 159.825 ;
        RECT 56.350 159.780 56.670 159.840 ;
        RECT 61.040 159.825 61.180 159.980 ;
        RECT 54.065 159.640 56.670 159.780 ;
        RECT 54.065 159.595 54.355 159.640 ;
        RECT 49.310 159.440 49.450 159.595 ;
        RECT 41.260 159.300 46.535 159.440 ;
        RECT 37.965 159.255 38.255 159.300 ;
        RECT 38.870 159.240 39.190 159.300 ;
        RECT 40.250 159.240 40.570 159.300 ;
        RECT 45.770 159.240 46.090 159.300 ;
        RECT 46.245 159.255 46.535 159.300 ;
        RECT 47.240 159.300 47.840 159.440 ;
        RECT 48.325 159.300 49.450 159.440 ;
        RECT 49.910 159.440 50.230 159.500 ;
        RECT 50.920 159.440 51.060 159.595 ;
        RECT 49.910 159.300 51.060 159.440 ;
        RECT 52.300 159.440 52.440 159.595 ;
        RECT 56.350 159.580 56.670 159.640 ;
        RECT 60.965 159.595 61.255 159.825 ;
        RECT 61.885 159.595 62.175 159.825 ;
        RECT 58.190 159.440 58.510 159.500 ;
        RECT 61.040 159.440 61.180 159.595 ;
        RECT 52.300 159.300 61.180 159.440 ;
        RECT 40.710 159.100 41.030 159.160 ;
        RECT 34.360 158.960 41.030 159.100 ;
        RECT 40.710 158.900 41.030 158.960 ;
        RECT 42.565 159.100 42.855 159.145 ;
        RECT 43.470 159.100 43.790 159.160 ;
        RECT 42.565 158.960 43.790 159.100 ;
        RECT 42.565 158.915 42.855 158.960 ;
        RECT 43.470 158.900 43.790 158.960 ;
        RECT 22.310 158.560 22.630 158.820 ;
        RECT 33.825 158.760 34.115 158.805 ;
        RECT 47.240 158.760 47.380 159.300 ;
        RECT 48.325 159.160 48.465 159.300 ;
        RECT 49.910 159.240 50.230 159.300 ;
        RECT 58.190 159.240 58.510 159.300 ;
        RECT 48.070 158.960 48.465 159.160 ;
        RECT 53.130 159.100 53.450 159.160 ;
        RECT 55.430 159.100 55.750 159.160 ;
        RECT 58.650 159.100 58.970 159.160 ;
        RECT 61.960 159.100 62.100 159.595 ;
        RECT 62.420 159.500 62.560 159.980 ;
        RECT 63.250 159.580 63.570 159.840 ;
        RECT 64.260 159.825 64.400 159.980 ;
        RECT 64.630 159.980 67.160 160.120 ;
        RECT 64.630 159.920 64.950 159.980 ;
        RECT 67.020 159.825 67.160 159.980 ;
        RECT 71.990 159.980 73.690 160.120 ;
        RECT 71.990 159.920 72.310 159.980 ;
        RECT 64.185 159.595 64.475 159.825 ;
        RECT 65.565 159.780 65.855 159.825 ;
        RECT 64.720 159.640 65.855 159.780 ;
        RECT 62.330 159.440 62.650 159.500 ;
        RECT 64.720 159.440 64.860 159.640 ;
        RECT 65.565 159.595 65.855 159.640 ;
        RECT 66.945 159.595 67.235 159.825 ;
        RECT 70.610 159.780 70.930 159.840 ;
        RECT 71.085 159.780 71.375 159.825 ;
        RECT 70.610 159.640 71.375 159.780 ;
        RECT 70.610 159.580 70.930 159.640 ;
        RECT 71.085 159.595 71.375 159.640 ;
        RECT 71.545 159.780 71.835 159.825 ;
        RECT 72.450 159.780 72.770 159.840 ;
        RECT 73.000 159.825 73.140 159.980 ;
        RECT 73.370 159.920 73.690 159.980 ;
        RECT 71.545 159.640 72.770 159.780 ;
        RECT 71.545 159.595 71.835 159.640 ;
        RECT 72.450 159.580 72.770 159.640 ;
        RECT 72.925 159.595 73.215 159.825 ;
        RECT 74.535 159.780 74.825 159.995 ;
        RECT 75.670 159.920 75.990 160.180 ;
        RECT 76.590 160.165 76.910 160.180 ;
        RECT 76.590 159.935 76.975 160.165 ;
        RECT 78.905 160.120 79.195 160.165 ;
        RECT 83.490 160.120 83.810 160.180 ;
        RECT 78.905 159.980 83.810 160.120 ;
        RECT 78.905 159.935 79.195 159.980 ;
        RECT 76.590 159.920 76.910 159.935 ;
        RECT 83.490 159.920 83.810 159.980 ;
        RECT 73.460 159.765 74.825 159.780 ;
        RECT 73.460 159.640 74.750 159.765 ;
        RECT 62.330 159.300 64.860 159.440 ;
        RECT 65.090 159.440 65.410 159.500 ;
        RECT 67.865 159.440 68.155 159.485 ;
        RECT 73.460 159.440 73.600 159.640 ;
        RECT 65.090 159.300 73.600 159.440 ;
        RECT 62.330 159.240 62.650 159.300 ;
        RECT 65.090 159.240 65.410 159.300 ;
        RECT 67.865 159.255 68.155 159.300 ;
        RECT 53.130 158.960 62.100 159.100 ;
        RECT 62.805 159.100 63.095 159.145 ;
        RECT 71.990 159.100 72.310 159.160 ;
        RECT 72.465 159.100 72.755 159.145 ;
        RECT 74.750 159.100 75.070 159.160 ;
        RECT 62.805 158.960 76.820 159.100 ;
        RECT 48.070 158.900 48.390 158.960 ;
        RECT 53.130 158.900 53.450 158.960 ;
        RECT 55.430 158.900 55.750 158.960 ;
        RECT 58.650 158.900 58.970 158.960 ;
        RECT 62.805 158.915 63.095 158.960 ;
        RECT 71.990 158.900 72.310 158.960 ;
        RECT 72.465 158.915 72.755 158.960 ;
        RECT 74.750 158.900 75.070 158.960 ;
        RECT 33.825 158.620 47.380 158.760 ;
        RECT 47.610 158.760 47.930 158.820 ;
        RECT 49.450 158.760 49.770 158.820 ;
        RECT 47.610 158.620 49.770 158.760 ;
        RECT 33.825 158.575 34.115 158.620 ;
        RECT 47.610 158.560 47.930 158.620 ;
        RECT 49.450 158.560 49.770 158.620 ;
        RECT 50.830 158.760 51.150 158.820 ;
        RECT 54.050 158.760 54.370 158.820 ;
        RECT 50.830 158.620 54.370 158.760 ;
        RECT 50.830 158.560 51.150 158.620 ;
        RECT 54.050 158.560 54.370 158.620 ;
        RECT 60.490 158.760 60.810 158.820 ;
        RECT 68.770 158.760 69.090 158.820 ;
        RECT 71.530 158.760 71.850 158.820 ;
        RECT 60.490 158.620 71.850 158.760 ;
        RECT 60.490 158.560 60.810 158.620 ;
        RECT 68.770 158.560 69.090 158.620 ;
        RECT 71.530 158.560 71.850 158.620 ;
        RECT 72.910 158.760 73.230 158.820 ;
        RECT 76.680 158.805 76.820 158.960 ;
        RECT 74.305 158.760 74.595 158.805 ;
        RECT 72.910 158.620 74.595 158.760 ;
        RECT 72.910 158.560 73.230 158.620 ;
        RECT 74.305 158.575 74.595 158.620 ;
        RECT 76.605 158.575 76.895 158.805 ;
        RECT 18.100 157.940 89.400 158.420 ;
        RECT 21.390 157.540 21.710 157.800 ;
        RECT 23.690 157.740 24.010 157.800 ;
        RECT 26.005 157.740 26.295 157.785 ;
        RECT 23.690 157.600 26.295 157.740 ;
        RECT 23.690 157.540 24.010 157.600 ;
        RECT 26.005 157.555 26.295 157.600 ;
        RECT 26.450 157.540 26.770 157.800 ;
        RECT 29.210 157.740 29.530 157.800 ;
        RECT 31.970 157.740 32.290 157.800 ;
        RECT 29.210 157.600 32.290 157.740 ;
        RECT 29.210 157.540 29.530 157.600 ;
        RECT 31.970 157.540 32.290 157.600 ;
        RECT 39.790 157.540 40.110 157.800 ;
        RECT 45.770 157.740 46.090 157.800 ;
        RECT 49.465 157.740 49.755 157.785 ;
        RECT 45.770 157.600 55.200 157.740 ;
        RECT 45.770 157.540 46.090 157.600 ;
        RECT 49.465 157.555 49.755 157.600 ;
        RECT 22.310 157.400 22.630 157.460 ;
        RECT 24.165 157.400 24.455 157.445 ;
        RECT 27.370 157.400 27.690 157.460 ;
        RECT 20.560 157.260 27.690 157.400 ;
        RECT 20.560 156.765 20.700 157.260 ;
        RECT 22.310 157.200 22.630 157.260 ;
        RECT 24.165 157.215 24.455 157.260 ;
        RECT 27.370 157.200 27.690 157.260 ;
        RECT 36.570 157.400 36.890 157.460 ;
        RECT 38.410 157.400 38.730 157.460 ;
        RECT 48.070 157.400 48.390 157.460 ;
        RECT 36.570 157.260 38.180 157.400 ;
        RECT 36.570 157.200 36.890 157.260 ;
        RECT 21.865 156.875 22.155 157.105 ;
        RECT 24.610 157.060 24.930 157.120 ;
        RECT 38.040 157.105 38.180 157.260 ;
        RECT 38.410 157.260 48.390 157.400 ;
        RECT 38.410 157.200 38.730 157.260 ;
        RECT 48.070 157.200 48.390 157.260 ;
        RECT 53.590 157.200 53.910 157.460 ;
        RECT 54.525 157.400 54.815 157.445 ;
        RECT 54.140 157.260 54.815 157.400 ;
        RECT 55.060 157.400 55.200 157.600 ;
        RECT 65.550 157.540 65.870 157.800 ;
        RECT 66.930 157.740 67.250 157.800 ;
        RECT 67.405 157.740 67.695 157.785 ;
        RECT 66.930 157.600 67.695 157.740 ;
        RECT 66.930 157.540 67.250 157.600 ;
        RECT 67.405 157.555 67.695 157.600 ;
        RECT 71.990 157.540 72.310 157.800 ;
        RECT 72.925 157.740 73.215 157.785 ;
        RECT 73.830 157.740 74.150 157.800 ;
        RECT 72.925 157.600 74.150 157.740 ;
        RECT 72.925 157.555 73.215 157.600 ;
        RECT 73.830 157.540 74.150 157.600 ;
        RECT 74.305 157.740 74.595 157.785 ;
        RECT 78.890 157.740 79.210 157.800 ;
        RECT 74.305 157.600 79.210 157.740 ;
        RECT 74.305 157.555 74.595 157.600 ;
        RECT 78.890 157.540 79.210 157.600 ;
        RECT 80.270 157.540 80.590 157.800 ;
        RECT 64.185 157.400 64.475 157.445 ;
        RECT 70.610 157.400 70.930 157.460 ;
        RECT 55.060 157.260 59.800 157.400 ;
        RECT 25.545 157.060 25.835 157.105 ;
        RECT 37.965 157.060 38.255 157.105 ;
        RECT 39.790 157.060 40.110 157.120 ;
        RECT 54.140 157.060 54.280 157.260 ;
        RECT 54.525 157.215 54.815 157.260 ;
        RECT 55.430 157.060 55.750 157.120 ;
        RECT 59.125 157.060 59.415 157.105 ;
        RECT 24.610 156.920 25.835 157.060 ;
        RECT 20.485 156.535 20.775 156.765 ;
        RECT 20.945 156.535 21.235 156.765 ;
        RECT 21.940 156.720 22.080 156.875 ;
        RECT 24.610 156.860 24.930 156.920 ;
        RECT 25.545 156.875 25.835 156.920 ;
        RECT 26.540 156.920 37.720 157.060 ;
        RECT 26.540 156.720 26.680 156.920 ;
        RECT 21.940 156.580 26.680 156.720 ;
        RECT 26.925 156.720 27.215 156.765 ;
        RECT 27.370 156.720 27.690 156.780 ;
        RECT 26.925 156.580 27.690 156.720 ;
        RECT 26.925 156.535 27.215 156.580 ;
        RECT 21.020 156.380 21.160 156.535 ;
        RECT 27.370 156.520 27.690 156.580 ;
        RECT 32.905 156.720 33.195 156.765 ;
        RECT 36.570 156.720 36.890 156.780 ;
        RECT 32.905 156.580 36.890 156.720 ;
        RECT 37.580 156.720 37.720 156.920 ;
        RECT 37.965 156.920 40.110 157.060 ;
        RECT 37.965 156.875 38.255 156.920 ;
        RECT 39.790 156.860 40.110 156.920 ;
        RECT 49.080 156.920 53.360 157.060 ;
        RECT 54.140 156.920 55.750 157.060 ;
        RECT 49.080 156.780 49.220 156.920 ;
        RECT 38.885 156.720 39.175 156.765 ;
        RECT 43.010 156.720 43.330 156.780 ;
        RECT 37.580 156.580 43.330 156.720 ;
        RECT 32.905 156.535 33.195 156.580 ;
        RECT 36.570 156.520 36.890 156.580 ;
        RECT 38.885 156.535 39.175 156.580 ;
        RECT 43.010 156.520 43.330 156.580 ;
        RECT 48.545 156.720 48.835 156.765 ;
        RECT 48.990 156.720 49.310 156.780 ;
        RECT 48.545 156.580 49.310 156.720 ;
        RECT 48.545 156.535 48.835 156.580 ;
        RECT 48.990 156.520 49.310 156.580 ;
        RECT 49.925 156.720 50.215 156.765 ;
        RECT 50.830 156.720 51.150 156.780 ;
        RECT 49.925 156.580 51.150 156.720 ;
        RECT 49.925 156.535 50.215 156.580 ;
        RECT 50.830 156.520 51.150 156.580 ;
        RECT 52.210 156.520 52.530 156.780 ;
        RECT 53.220 156.720 53.360 156.920 ;
        RECT 55.430 156.860 55.750 156.920 ;
        RECT 57.360 156.920 59.415 157.060 ;
        RECT 57.360 156.720 57.500 156.920 ;
        RECT 59.125 156.875 59.415 156.920 ;
        RECT 53.220 156.580 57.500 156.720 ;
        RECT 57.745 156.720 58.035 156.765 ;
        RECT 58.190 156.720 58.510 156.780 ;
        RECT 57.745 156.580 58.510 156.720 ;
        RECT 57.745 156.535 58.035 156.580 ;
        RECT 58.190 156.520 58.510 156.580 ;
        RECT 22.325 156.380 22.615 156.425 ;
        RECT 26.450 156.380 26.770 156.440 ;
        RECT 21.020 156.240 26.770 156.380 ;
        RECT 43.100 156.380 43.240 156.520 ;
        RECT 59.200 156.380 59.340 156.875 ;
        RECT 59.660 156.720 59.800 157.260 ;
        RECT 64.185 157.260 70.930 157.400 ;
        RECT 64.185 157.215 64.475 157.260 ;
        RECT 70.610 157.200 70.930 157.260 ;
        RECT 71.160 157.260 80.960 157.400 ;
        RECT 63.710 157.060 64.030 157.120 ;
        RECT 65.565 157.060 65.855 157.105 ;
        RECT 63.710 156.920 65.855 157.060 ;
        RECT 63.710 156.860 64.030 156.920 ;
        RECT 65.565 156.875 65.855 156.920 ;
        RECT 66.010 157.060 66.330 157.120 ;
        RECT 71.160 157.060 71.300 157.260 ;
        RECT 80.820 157.105 80.960 157.260 ;
        RECT 66.010 156.920 71.300 157.060 ;
        RECT 80.745 157.060 81.035 157.105 ;
        RECT 80.745 156.920 86.940 157.060 ;
        RECT 66.010 156.860 66.330 156.920 ;
        RECT 80.745 156.875 81.035 156.920 ;
        RECT 86.800 156.780 86.940 156.920 ;
        RECT 60.045 156.720 60.335 156.765 ;
        RECT 61.870 156.720 62.190 156.780 ;
        RECT 59.660 156.580 62.190 156.720 ;
        RECT 60.045 156.535 60.335 156.580 ;
        RECT 61.870 156.520 62.190 156.580 ;
        RECT 62.330 156.720 62.650 156.780 ;
        RECT 62.805 156.720 63.095 156.765 ;
        RECT 62.330 156.580 63.095 156.720 ;
        RECT 62.330 156.520 62.650 156.580 ;
        RECT 62.805 156.535 63.095 156.580 ;
        RECT 63.250 156.520 63.570 156.780 ;
        RECT 65.090 156.520 65.410 156.780 ;
        RECT 66.485 156.535 66.775 156.765 ;
        RECT 70.150 156.720 70.470 156.780 ;
        RECT 73.370 156.720 73.690 156.780 ;
        RECT 70.150 156.580 73.690 156.720 ;
        RECT 64.185 156.380 64.475 156.425 ;
        RECT 64.630 156.380 64.950 156.440 ;
        RECT 66.560 156.380 66.700 156.535 ;
        RECT 70.150 156.520 70.470 156.580 ;
        RECT 73.370 156.520 73.690 156.580 ;
        RECT 74.305 156.720 74.595 156.765 ;
        RECT 76.590 156.720 76.910 156.780 ;
        RECT 74.305 156.580 76.910 156.720 ;
        RECT 74.305 156.535 74.595 156.580 ;
        RECT 71.085 156.380 71.375 156.425 ;
        RECT 74.380 156.380 74.520 156.535 ;
        RECT 76.590 156.520 76.910 156.580 ;
        RECT 79.365 156.720 79.655 156.765 ;
        RECT 81.190 156.720 81.510 156.780 ;
        RECT 79.365 156.580 81.510 156.720 ;
        RECT 79.365 156.535 79.655 156.580 ;
        RECT 81.190 156.520 81.510 156.580 ;
        RECT 83.505 156.535 83.795 156.765 ;
        RECT 43.100 156.240 54.280 156.380 ;
        RECT 59.200 156.240 64.950 156.380 ;
        RECT 22.325 156.195 22.615 156.240 ;
        RECT 26.450 156.180 26.770 156.240 ;
        RECT 24.625 156.040 24.915 156.085 ;
        RECT 31.050 156.040 31.370 156.100 ;
        RECT 24.625 155.900 31.370 156.040 ;
        RECT 24.625 155.855 24.915 155.900 ;
        RECT 31.050 155.840 31.370 155.900 ;
        RECT 47.610 155.840 47.930 156.100 ;
        RECT 54.140 156.040 54.280 156.240 ;
        RECT 64.185 156.195 64.475 156.240 ;
        RECT 64.630 156.180 64.950 156.240 ;
        RECT 65.180 156.240 71.375 156.380 ;
        RECT 65.180 156.100 65.320 156.240 ;
        RECT 71.085 156.195 71.375 156.240 ;
        RECT 72.540 156.240 74.520 156.380 ;
        RECT 81.665 156.380 81.955 156.425 ;
        RECT 82.110 156.380 82.430 156.440 ;
        RECT 81.665 156.240 82.430 156.380 ;
        RECT 58.205 156.040 58.495 156.085 ;
        RECT 54.140 155.900 58.495 156.040 ;
        RECT 58.205 155.855 58.495 155.900 ;
        RECT 58.650 155.840 58.970 156.100 ;
        RECT 59.110 155.840 59.430 156.100 ;
        RECT 65.090 155.840 65.410 156.100 ;
        RECT 70.610 156.040 70.930 156.100 ;
        RECT 72.085 156.040 72.375 156.085 ;
        RECT 72.540 156.040 72.680 156.240 ;
        RECT 81.665 156.195 81.955 156.240 ;
        RECT 82.110 156.180 82.430 156.240 ;
        RECT 70.610 155.900 72.680 156.040 ;
        RECT 81.190 156.040 81.510 156.100 ;
        RECT 83.580 156.040 83.720 156.535 ;
        RECT 86.250 156.520 86.570 156.780 ;
        RECT 86.710 156.720 87.030 156.780 ;
        RECT 87.185 156.720 87.475 156.765 ;
        RECT 86.710 156.580 87.475 156.720 ;
        RECT 86.710 156.520 87.030 156.580 ;
        RECT 87.185 156.535 87.475 156.580 ;
        RECT 81.190 155.900 83.720 156.040 ;
        RECT 84.425 156.040 84.715 156.085 ;
        RECT 84.870 156.040 85.190 156.100 ;
        RECT 84.425 155.900 85.190 156.040 ;
        RECT 70.610 155.840 70.930 155.900 ;
        RECT 72.085 155.855 72.375 155.900 ;
        RECT 81.190 155.840 81.510 155.900 ;
        RECT 84.425 155.855 84.715 155.900 ;
        RECT 84.870 155.840 85.190 155.900 ;
        RECT 86.725 156.040 87.015 156.085 ;
        RECT 87.630 156.040 87.950 156.100 ;
        RECT 86.725 155.900 87.950 156.040 ;
        RECT 86.725 155.855 87.015 155.900 ;
        RECT 87.630 155.840 87.950 155.900 ;
        RECT 18.100 155.220 89.400 155.700 ;
        RECT 25.530 155.020 25.850 155.080 ;
        RECT 26.465 155.020 26.755 155.065 ;
        RECT 25.530 154.880 26.755 155.020 ;
        RECT 25.530 154.820 25.850 154.880 ;
        RECT 26.465 154.835 26.755 154.880 ;
        RECT 28.305 155.020 28.595 155.065 ;
        RECT 42.550 155.020 42.870 155.080 ;
        RECT 28.305 154.880 42.870 155.020 ;
        RECT 28.305 154.835 28.595 154.880 ;
        RECT 42.550 154.820 42.870 154.880 ;
        RECT 44.390 154.820 44.710 155.080 ;
        RECT 60.030 155.020 60.350 155.080 ;
        RECT 46.320 154.880 60.350 155.020 ;
        RECT 29.210 154.480 29.530 154.740 ;
        RECT 29.670 154.680 29.990 154.740 ;
        RECT 39.345 154.680 39.635 154.725 ;
        RECT 46.320 154.680 46.460 154.880 ;
        RECT 60.030 154.820 60.350 154.880 ;
        RECT 71.070 155.020 71.390 155.080 ;
        RECT 71.070 154.880 72.220 155.020 ;
        RECT 71.070 154.820 71.390 154.880 ;
        RECT 47.610 154.680 47.930 154.740 ;
        RECT 29.670 154.540 38.640 154.680 ;
        RECT 29.670 154.480 29.990 154.540 ;
        RECT 29.760 154.200 32.200 154.340 ;
        RECT 19.550 153.800 19.870 154.060 ;
        RECT 20.945 154.000 21.235 154.045 ;
        RECT 25.085 154.000 25.375 154.045 ;
        RECT 20.945 153.860 25.375 154.000 ;
        RECT 20.945 153.815 21.235 153.860 ;
        RECT 25.085 153.815 25.375 153.860 ;
        RECT 25.160 153.660 25.300 153.815 ;
        RECT 26.910 153.800 27.230 154.060 ;
        RECT 27.370 154.045 27.690 154.060 ;
        RECT 27.370 154.000 27.800 154.045 ;
        RECT 29.760 154.000 29.900 154.200 ;
        RECT 32.060 154.060 32.200 154.200 ;
        RECT 36.110 154.140 36.430 154.400 ;
        RECT 37.030 154.140 37.350 154.400 ;
        RECT 38.500 154.385 38.640 154.540 ;
        RECT 39.345 154.540 46.460 154.680 ;
        RECT 46.780 154.540 47.930 154.680 ;
        RECT 39.345 154.495 39.635 154.540 ;
        RECT 38.425 154.340 38.715 154.385 ;
        RECT 39.790 154.340 40.110 154.400 ;
        RECT 38.425 154.200 40.110 154.340 ;
        RECT 38.425 154.155 38.715 154.200 ;
        RECT 39.790 154.140 40.110 154.200 ;
        RECT 45.325 154.155 45.615 154.385 ;
        RECT 45.785 154.340 46.075 154.385 ;
        RECT 46.230 154.340 46.550 154.400 ;
        RECT 46.780 154.385 46.920 154.540 ;
        RECT 47.610 154.480 47.930 154.540 ;
        RECT 48.070 154.680 48.390 154.740 ;
        RECT 52.670 154.680 52.990 154.740 ;
        RECT 64.645 154.680 64.935 154.725 ;
        RECT 48.070 154.540 52.440 154.680 ;
        RECT 48.070 154.480 48.390 154.540 ;
        RECT 45.785 154.200 46.550 154.340 ;
        RECT 45.785 154.155 46.075 154.200 ;
        RECT 27.370 153.860 29.900 154.000 ;
        RECT 27.370 153.815 27.800 153.860 ;
        RECT 27.370 153.800 27.690 153.815 ;
        RECT 31.510 153.800 31.830 154.060 ;
        RECT 31.970 153.800 32.290 154.060 ;
        RECT 45.400 154.000 45.540 154.155 ;
        RECT 46.230 154.140 46.550 154.200 ;
        RECT 46.705 154.155 46.995 154.385 ;
        RECT 47.150 154.140 47.470 154.400 ;
        RECT 48.545 154.340 48.835 154.385 ;
        RECT 48.990 154.340 49.310 154.400 ;
        RECT 48.545 154.200 49.310 154.340 ;
        RECT 48.545 154.155 48.835 154.200 ;
        RECT 47.625 154.000 47.915 154.045 ;
        RECT 45.400 153.860 47.915 154.000 ;
        RECT 47.625 153.815 47.915 153.860 ;
        RECT 26.450 153.660 26.770 153.720 ;
        RECT 29.210 153.660 29.530 153.720 ;
        RECT 25.160 153.520 29.530 153.660 ;
        RECT 31.600 153.660 31.740 153.800 ;
        RECT 32.905 153.660 33.195 153.705 ;
        RECT 48.620 153.660 48.760 154.155 ;
        RECT 48.990 154.140 49.310 154.200 ;
        RECT 49.450 154.140 49.770 154.400 ;
        RECT 49.910 154.140 50.230 154.400 ;
        RECT 52.300 154.385 52.440 154.540 ;
        RECT 52.670 154.540 64.935 154.680 ;
        RECT 52.670 154.480 52.990 154.540 ;
        RECT 64.645 154.495 64.935 154.540 ;
        RECT 52.225 154.155 52.515 154.385 ;
        RECT 53.145 154.340 53.435 154.385 ;
        RECT 54.050 154.340 54.370 154.400 ;
        RECT 53.145 154.200 54.370 154.340 ;
        RECT 53.145 154.155 53.435 154.200 ;
        RECT 52.300 154.000 52.440 154.155 ;
        RECT 54.050 154.140 54.370 154.200 ;
        RECT 65.105 154.155 65.395 154.385 ;
        RECT 69.690 154.340 70.010 154.400 ;
        RECT 70.165 154.340 70.455 154.385 ;
        RECT 69.690 154.200 70.455 154.340 ;
        RECT 53.590 154.000 53.910 154.060 ;
        RECT 52.300 153.860 53.910 154.000 ;
        RECT 65.180 154.000 65.320 154.155 ;
        RECT 69.690 154.140 70.010 154.200 ;
        RECT 70.165 154.155 70.455 154.200 ;
        RECT 70.625 154.340 70.915 154.385 ;
        RECT 71.070 154.340 71.390 154.400 ;
        RECT 70.625 154.200 71.390 154.340 ;
        RECT 70.625 154.155 70.915 154.200 ;
        RECT 70.700 154.000 70.840 154.155 ;
        RECT 71.070 154.140 71.390 154.200 ;
        RECT 71.545 154.155 71.835 154.385 ;
        RECT 72.080 154.340 72.220 154.880 ;
        RECT 72.450 154.820 72.770 155.080 ;
        RECT 83.965 155.020 84.255 155.065 ;
        RECT 84.410 155.020 84.730 155.080 ;
        RECT 83.965 154.880 84.730 155.020 ;
        RECT 83.965 154.835 84.255 154.880 ;
        RECT 84.410 154.820 84.730 154.880 ;
        RECT 84.885 154.835 85.175 155.065 ;
        RECT 81.190 154.680 81.510 154.740 ;
        RECT 84.960 154.680 85.100 154.835 ;
        RECT 87.170 154.820 87.490 155.080 ;
        RECT 86.710 154.680 87.030 154.740 ;
        RECT 89.010 154.680 89.330 154.740 ;
        RECT 74.380 154.540 85.100 154.680 ;
        RECT 85.880 154.540 89.330 154.680 ;
        RECT 73.845 154.340 74.135 154.385 ;
        RECT 72.080 154.200 74.135 154.340 ;
        RECT 73.845 154.155 74.135 154.200 ;
        RECT 71.620 154.000 71.760 154.155 ;
        RECT 71.990 154.000 72.310 154.060 ;
        RECT 65.180 153.860 70.840 154.000 ;
        RECT 71.160 153.860 72.310 154.000 ;
        RECT 53.590 153.800 53.910 153.860 ;
        RECT 54.970 153.660 55.290 153.720 ;
        RECT 31.600 153.520 32.200 153.660 ;
        RECT 26.450 153.460 26.770 153.520 ;
        RECT 29.210 153.460 29.530 153.520 ;
        RECT 32.060 153.320 32.200 153.520 ;
        RECT 32.905 153.520 48.760 153.660 ;
        RECT 49.080 153.520 55.290 153.660 ;
        RECT 32.905 153.475 33.195 153.520 ;
        RECT 43.930 153.320 44.250 153.380 ;
        RECT 49.080 153.320 49.220 153.520 ;
        RECT 54.970 153.460 55.290 153.520 ;
        RECT 55.430 153.660 55.750 153.720 ;
        RECT 60.030 153.660 60.350 153.720 ;
        RECT 68.310 153.660 68.630 153.720 ;
        RECT 71.160 153.660 71.300 153.860 ;
        RECT 71.990 153.800 72.310 153.860 ;
        RECT 55.430 153.520 71.300 153.660 ;
        RECT 71.530 153.660 71.850 153.720 ;
        RECT 72.925 153.660 73.215 153.705 ;
        RECT 71.530 153.520 73.215 153.660 ;
        RECT 55.430 153.460 55.750 153.520 ;
        RECT 60.030 153.460 60.350 153.520 ;
        RECT 68.310 153.460 68.630 153.520 ;
        RECT 71.530 153.460 71.850 153.520 ;
        RECT 72.925 153.475 73.215 153.520 ;
        RECT 32.060 153.180 49.220 153.320 ;
        RECT 43.930 153.120 44.250 153.180 ;
        RECT 53.130 153.120 53.450 153.380 ;
        RECT 53.590 153.320 53.910 153.380 ;
        RECT 55.520 153.320 55.660 153.460 ;
        RECT 53.590 153.180 55.660 153.320 ;
        RECT 60.950 153.320 61.270 153.380 ;
        RECT 74.380 153.320 74.520 154.540 ;
        RECT 81.190 154.480 81.510 154.540 ;
        RECT 82.570 154.140 82.890 154.400 ;
        RECT 83.045 154.340 83.335 154.385 ;
        RECT 83.950 154.340 84.270 154.400 ;
        RECT 85.880 154.385 86.020 154.540 ;
        RECT 86.710 154.480 87.030 154.540 ;
        RECT 89.010 154.480 89.330 154.540 ;
        RECT 83.045 154.200 84.270 154.340 ;
        RECT 83.045 154.155 83.335 154.200 ;
        RECT 83.950 154.140 84.270 154.200 ;
        RECT 85.805 154.155 86.095 154.385 ;
        RECT 86.265 154.155 86.555 154.385 ;
        RECT 74.765 153.815 75.055 154.045 ;
        RECT 83.490 154.000 83.810 154.060 ;
        RECT 86.340 154.000 86.480 154.155 ;
        RECT 83.490 153.860 86.480 154.000 ;
        RECT 74.840 153.660 74.980 153.815 ;
        RECT 83.490 153.800 83.810 153.860 ;
        RECT 87.630 153.660 87.950 153.720 ;
        RECT 74.840 153.520 87.950 153.660 ;
        RECT 87.630 153.460 87.950 153.520 ;
        RECT 60.950 153.180 74.520 153.320 ;
        RECT 53.590 153.120 53.910 153.180 ;
        RECT 60.950 153.120 61.270 153.180 ;
        RECT 81.650 153.120 81.970 153.380 ;
        RECT 18.100 152.500 89.400 152.980 ;
        RECT 24.625 152.300 24.915 152.345 ;
        RECT 25.070 152.300 25.390 152.360 ;
        RECT 24.625 152.160 25.390 152.300 ;
        RECT 24.625 152.115 24.915 152.160 ;
        RECT 25.070 152.100 25.390 152.160 ;
        RECT 25.530 152.300 25.850 152.360 ;
        RECT 29.225 152.300 29.515 152.345 ;
        RECT 32.430 152.300 32.750 152.360 ;
        RECT 33.365 152.300 33.655 152.345 ;
        RECT 25.530 152.160 29.515 152.300 ;
        RECT 25.530 152.100 25.850 152.160 ;
        RECT 29.225 152.115 29.515 152.160 ;
        RECT 29.760 152.160 33.655 152.300 ;
        RECT 24.165 151.960 24.455 152.005 ;
        RECT 26.450 151.960 26.770 152.020 ;
        RECT 24.165 151.820 26.770 151.960 ;
        RECT 24.165 151.775 24.455 151.820 ;
        RECT 24.240 151.620 24.380 151.775 ;
        RECT 26.450 151.760 26.770 151.820 ;
        RECT 26.910 151.960 27.230 152.020 ;
        RECT 27.385 151.960 27.675 152.005 ;
        RECT 29.760 151.960 29.900 152.160 ;
        RECT 32.430 152.100 32.750 152.160 ;
        RECT 33.365 152.115 33.655 152.160 ;
        RECT 37.030 152.300 37.350 152.360 ;
        RECT 45.325 152.300 45.615 152.345 ;
        RECT 47.150 152.300 47.470 152.360 ;
        RECT 37.030 152.160 44.620 152.300 ;
        RECT 37.030 152.100 37.350 152.160 ;
        RECT 26.910 151.820 29.900 151.960 ;
        RECT 34.285 151.960 34.575 152.005 ;
        RECT 36.110 151.960 36.430 152.020 ;
        RECT 34.285 151.820 37.260 151.960 ;
        RECT 26.910 151.760 27.230 151.820 ;
        RECT 27.385 151.775 27.675 151.820 ;
        RECT 34.285 151.775 34.575 151.820 ;
        RECT 36.110 151.760 36.430 151.820 ;
        RECT 21.020 151.480 24.380 151.620 ;
        RECT 31.600 151.480 36.800 151.620 ;
        RECT 21.020 151.325 21.160 151.480 ;
        RECT 20.945 151.095 21.235 151.325 ;
        RECT 21.865 151.095 22.155 151.325 ;
        RECT 25.530 151.280 25.850 151.340 ;
        RECT 31.600 151.325 31.740 151.480 ;
        RECT 31.525 151.280 31.815 151.325 ;
        RECT 25.530 151.140 31.815 151.280 ;
        RECT 21.390 150.940 21.710 151.000 ;
        RECT 21.940 150.940 22.080 151.095 ;
        RECT 25.530 151.080 25.850 151.140 ;
        RECT 31.525 151.095 31.815 151.140 ;
        RECT 35.650 151.080 35.970 151.340 ;
        RECT 36.110 151.280 36.430 151.340 ;
        RECT 36.660 151.325 36.800 151.480 ;
        RECT 36.585 151.280 36.875 151.325 ;
        RECT 36.110 151.140 36.875 151.280 ;
        RECT 37.120 151.280 37.260 151.820 ;
        RECT 37.505 151.620 37.795 151.665 ;
        RECT 37.505 151.480 42.780 151.620 ;
        RECT 37.505 151.435 37.795 151.480 ;
        RECT 42.640 151.340 42.780 151.480 ;
        RECT 37.965 151.280 38.255 151.325 ;
        RECT 41.645 151.280 41.935 151.325 ;
        RECT 37.120 151.140 41.935 151.280 ;
        RECT 36.110 151.080 36.430 151.140 ;
        RECT 36.585 151.095 36.875 151.140 ;
        RECT 37.965 151.095 38.255 151.140 ;
        RECT 41.645 151.095 41.935 151.140 ;
        RECT 22.325 150.940 22.615 150.985 ;
        RECT 27.370 150.940 27.690 151.000 ;
        RECT 21.390 150.800 27.690 150.940 ;
        RECT 21.390 150.740 21.710 150.800 ;
        RECT 22.325 150.755 22.615 150.800 ;
        RECT 27.370 150.740 27.690 150.800 ;
        RECT 29.210 150.740 29.530 151.000 ;
        RECT 31.970 150.940 32.290 151.000 ;
        RECT 33.365 150.940 33.655 150.985 ;
        RECT 31.970 150.800 33.655 150.940 ;
        RECT 36.660 150.940 36.800 151.095 ;
        RECT 42.550 151.080 42.870 151.340 ;
        RECT 43.930 151.080 44.250 151.340 ;
        RECT 44.480 151.325 44.620 152.160 ;
        RECT 45.325 152.160 47.470 152.300 ;
        RECT 45.325 152.115 45.615 152.160 ;
        RECT 47.150 152.100 47.470 152.160 ;
        RECT 48.530 152.300 48.850 152.360 ;
        RECT 50.385 152.300 50.675 152.345 ;
        RECT 48.530 152.160 50.675 152.300 ;
        RECT 48.530 152.100 48.850 152.160 ;
        RECT 50.385 152.115 50.675 152.160 ;
        RECT 54.985 152.300 55.275 152.345 ;
        RECT 55.430 152.300 55.750 152.360 ;
        RECT 54.985 152.160 55.750 152.300 ;
        RECT 54.985 152.115 55.275 152.160 ;
        RECT 55.430 152.100 55.750 152.160 ;
        RECT 57.270 152.100 57.590 152.360 ;
        RECT 58.650 152.300 58.970 152.360 ;
        RECT 59.585 152.300 59.875 152.345 ;
        RECT 58.650 152.160 59.875 152.300 ;
        RECT 58.650 152.100 58.970 152.160 ;
        RECT 59.585 152.115 59.875 152.160 ;
        RECT 63.265 152.300 63.555 152.345 ;
        RECT 66.010 152.300 66.330 152.360 ;
        RECT 63.265 152.160 66.330 152.300 ;
        RECT 63.265 152.115 63.555 152.160 ;
        RECT 66.010 152.100 66.330 152.160 ;
        RECT 70.150 152.100 70.470 152.360 ;
        RECT 85.790 152.100 86.110 152.360 ;
        RECT 47.625 151.960 47.915 152.005 ;
        RECT 51.290 151.960 51.610 152.020 ;
        RECT 54.510 151.960 54.830 152.020 ;
        RECT 47.625 151.820 54.830 151.960 ;
        RECT 47.625 151.775 47.915 151.820 ;
        RECT 51.290 151.760 51.610 151.820 ;
        RECT 54.510 151.760 54.830 151.820 ;
        RECT 55.890 151.960 56.210 152.020 ;
        RECT 55.890 151.820 61.640 151.960 ;
        RECT 55.890 151.760 56.210 151.820 ;
        RECT 52.210 151.620 52.530 151.680 ;
        RECT 45.860 151.480 52.530 151.620 ;
        RECT 44.405 151.095 44.695 151.325 ;
        RECT 45.310 151.280 45.630 151.340 ;
        RECT 45.860 151.325 46.000 151.480 ;
        RECT 52.210 151.420 52.530 151.480 ;
        RECT 53.680 151.480 60.720 151.620 ;
        RECT 46.690 151.325 47.010 151.340 ;
        RECT 45.785 151.280 46.075 151.325 ;
        RECT 45.310 151.140 46.075 151.280 ;
        RECT 45.310 151.080 45.630 151.140 ;
        RECT 45.785 151.095 46.075 151.140 ;
        RECT 46.555 151.095 47.010 151.325 ;
        RECT 51.305 151.280 51.595 151.325 ;
        RECT 51.305 151.140 52.900 151.280 ;
        RECT 51.305 151.095 51.595 151.140 ;
        RECT 46.690 151.080 47.010 151.095 ;
        RECT 36.660 150.800 40.480 150.940 ;
        RECT 31.970 150.740 32.290 150.800 ;
        RECT 33.365 150.755 33.655 150.800 ;
        RECT 20.025 150.600 20.315 150.645 ;
        RECT 29.670 150.600 29.990 150.660 ;
        RECT 20.025 150.460 29.990 150.600 ;
        RECT 20.025 150.415 20.315 150.460 ;
        RECT 29.670 150.400 29.990 150.460 ;
        RECT 30.145 150.600 30.435 150.645 ;
        RECT 35.190 150.600 35.510 150.660 ;
        RECT 37.030 150.600 37.350 150.660 ;
        RECT 30.145 150.460 37.350 150.600 ;
        RECT 30.145 150.415 30.435 150.460 ;
        RECT 35.190 150.400 35.510 150.460 ;
        RECT 37.030 150.400 37.350 150.460 ;
        RECT 39.345 150.600 39.635 150.645 ;
        RECT 39.790 150.600 40.110 150.660 ;
        RECT 40.340 150.645 40.480 150.800 ;
        RECT 40.710 150.740 41.030 151.000 ;
        RECT 46.780 150.940 46.920 151.080 ;
        RECT 51.750 150.940 52.070 151.000 ;
        RECT 46.780 150.800 52.070 150.940 ;
        RECT 51.750 150.740 52.070 150.800 ;
        RECT 52.210 150.740 52.530 151.000 ;
        RECT 52.760 150.940 52.900 151.140 ;
        RECT 53.130 151.080 53.450 151.340 ;
        RECT 53.680 151.325 53.820 151.480 ;
        RECT 53.605 151.095 53.895 151.325 ;
        RECT 54.065 151.290 54.355 151.325 ;
        RECT 54.065 151.280 54.740 151.290 ;
        RECT 54.970 151.280 55.290 151.340 ;
        RECT 54.065 151.150 55.290 151.280 ;
        RECT 54.065 151.095 54.355 151.150 ;
        RECT 54.600 151.140 55.290 151.150 ;
        RECT 54.970 151.080 55.290 151.140 ;
        RECT 58.190 151.080 58.510 151.340 ;
        RECT 58.665 151.280 58.955 151.325 ;
        RECT 59.110 151.280 59.430 151.340 ;
        RECT 58.665 151.140 59.430 151.280 ;
        RECT 58.665 151.095 58.955 151.140 ;
        RECT 57.270 150.940 57.590 151.000 ;
        RECT 58.740 150.940 58.880 151.095 ;
        RECT 59.110 151.080 59.430 151.140 ;
        RECT 60.030 151.080 60.350 151.340 ;
        RECT 52.760 150.800 54.050 150.940 ;
        RECT 39.345 150.460 40.110 150.600 ;
        RECT 39.345 150.415 39.635 150.460 ;
        RECT 39.790 150.400 40.110 150.460 ;
        RECT 40.265 150.415 40.555 150.645 ;
        RECT 42.090 150.400 42.410 150.660 ;
        RECT 53.910 150.600 54.050 150.800 ;
        RECT 57.270 150.800 58.880 150.940 ;
        RECT 60.580 150.940 60.720 151.480 ;
        RECT 60.950 151.080 61.270 151.340 ;
        RECT 61.500 151.325 61.640 151.820 ;
        RECT 64.185 151.775 64.475 152.005 ;
        RECT 65.550 151.960 65.870 152.020 ;
        RECT 72.005 151.960 72.295 152.005 ;
        RECT 75.670 151.960 75.990 152.020 ;
        RECT 65.550 151.820 75.990 151.960 ;
        RECT 64.260 151.620 64.400 151.775 ;
        RECT 65.550 151.760 65.870 151.820 ;
        RECT 72.005 151.775 72.295 151.820 ;
        RECT 75.670 151.760 75.990 151.820 ;
        RECT 87.630 151.760 87.950 152.020 ;
        RECT 64.260 151.480 71.300 151.620 ;
        RECT 61.425 151.095 61.715 151.325 ;
        RECT 63.250 151.080 63.570 151.340 ;
        RECT 65.180 151.325 65.320 151.480 ;
        RECT 71.160 151.340 71.300 151.480 ;
        RECT 65.105 151.095 65.395 151.325 ;
        RECT 66.075 151.280 66.365 151.325 ;
        RECT 66.075 151.140 66.700 151.280 ;
        RECT 66.075 151.095 66.365 151.140 ;
        RECT 64.630 150.940 64.950 151.000 ;
        RECT 60.580 150.800 64.950 150.940 ;
        RECT 66.560 150.940 66.700 151.140 ;
        RECT 67.850 151.080 68.170 151.340 ;
        RECT 69.230 151.080 69.550 151.340 ;
        RECT 69.690 151.280 70.010 151.340 ;
        RECT 70.625 151.280 70.915 151.325 ;
        RECT 69.690 151.140 70.915 151.280 ;
        RECT 69.690 151.080 70.010 151.140 ;
        RECT 70.625 151.095 70.915 151.140 ;
        RECT 71.070 151.080 71.390 151.340 ;
        RECT 71.990 151.080 72.310 151.340 ;
        RECT 84.870 151.080 85.190 151.340 ;
        RECT 66.930 150.940 67.250 151.000 ;
        RECT 69.780 150.940 69.920 151.080 ;
        RECT 66.560 150.800 69.920 150.940 ;
        RECT 81.650 150.940 81.970 151.000 ;
        RECT 86.725 150.940 87.015 150.985 ;
        RECT 81.650 150.800 87.015 150.940 ;
        RECT 57.270 150.740 57.590 150.800 ;
        RECT 64.630 150.740 64.950 150.800 ;
        RECT 66.930 150.740 67.250 150.800 ;
        RECT 81.650 150.740 81.970 150.800 ;
        RECT 86.725 150.755 87.015 150.800 ;
        RECT 55.890 150.600 56.210 150.660 ;
        RECT 65.105 150.600 65.395 150.645 ;
        RECT 53.910 150.460 65.395 150.600 ;
        RECT 55.890 150.400 56.210 150.460 ;
        RECT 65.105 150.415 65.395 150.460 ;
        RECT 68.310 150.400 68.630 150.660 ;
        RECT 18.100 149.780 89.400 150.260 ;
        RECT 36.110 149.380 36.430 149.640 ;
        RECT 37.965 149.580 38.255 149.625 ;
        RECT 49.910 149.580 50.230 149.640 ;
        RECT 65.550 149.580 65.870 149.640 ;
        RECT 36.660 149.440 50.230 149.580 ;
        RECT 35.190 149.040 35.510 149.300 ;
        RECT 35.650 149.240 35.970 149.300 ;
        RECT 36.660 149.240 36.800 149.440 ;
        RECT 37.965 149.395 38.255 149.440 ;
        RECT 49.910 149.380 50.230 149.440 ;
        RECT 53.680 149.440 65.870 149.580 ;
        RECT 35.650 149.100 36.800 149.240 ;
        RECT 35.650 149.040 35.970 149.100 ;
        RECT 20.945 148.715 21.235 148.945 ;
        RECT 21.020 148.560 21.160 148.715 ;
        RECT 21.390 148.700 21.710 148.960 ;
        RECT 36.660 148.945 36.800 149.100 ;
        RECT 51.750 149.040 52.070 149.300 ;
        RECT 21.865 148.900 22.155 148.945 ;
        RECT 23.705 148.900 23.995 148.945 ;
        RECT 21.865 148.760 23.995 148.900 ;
        RECT 21.865 148.715 22.155 148.760 ;
        RECT 23.705 148.715 23.995 148.760 ;
        RECT 36.585 148.715 36.875 148.945 ;
        RECT 37.045 148.715 37.335 148.945 ;
        RECT 51.305 148.715 51.595 148.945 ;
        RECT 25.070 148.560 25.390 148.620 ;
        RECT 37.120 148.560 37.260 148.715 ;
        RECT 21.020 148.420 23.000 148.560 ;
        RECT 20.010 148.020 20.330 148.280 ;
        RECT 22.860 148.265 23.000 148.420 ;
        RECT 25.070 148.420 37.260 148.560 ;
        RECT 25.070 148.360 25.390 148.420 ;
        RECT 22.785 148.035 23.075 148.265 ;
        RECT 50.370 148.020 50.690 148.280 ;
        RECT 35.205 147.880 35.495 147.925 ;
        RECT 35.650 147.880 35.970 147.940 ;
        RECT 35.205 147.740 35.970 147.880 ;
        RECT 51.380 147.880 51.520 148.715 ;
        RECT 52.210 148.700 52.530 148.960 ;
        RECT 53.680 148.945 53.820 149.440 ;
        RECT 65.550 149.380 65.870 149.440 ;
        RECT 66.100 149.440 69.460 149.580 ;
        RECT 56.810 149.240 57.130 149.300 ;
        RECT 57.745 149.240 58.035 149.285 ;
        RECT 60.030 149.240 60.350 149.300 ;
        RECT 66.100 149.240 66.240 149.440 ;
        RECT 69.320 149.300 69.460 149.440 ;
        RECT 68.310 149.240 68.630 149.300 ;
        RECT 54.140 149.100 56.580 149.240 ;
        RECT 54.140 148.960 54.280 149.100 ;
        RECT 53.145 148.715 53.435 148.945 ;
        RECT 53.605 148.715 53.895 148.945 ;
        RECT 53.220 148.560 53.360 148.715 ;
        RECT 54.050 148.700 54.370 148.960 ;
        RECT 54.970 148.700 55.290 148.960 ;
        RECT 55.890 148.700 56.210 148.960 ;
        RECT 56.440 148.945 56.580 149.100 ;
        RECT 56.810 149.100 58.035 149.240 ;
        RECT 56.810 149.040 57.130 149.100 ;
        RECT 57.745 149.055 58.035 149.100 ;
        RECT 59.200 149.100 60.350 149.240 ;
        RECT 56.365 148.715 56.655 148.945 ;
        RECT 57.270 148.700 57.590 148.960 ;
        RECT 58.190 148.900 58.510 148.960 ;
        RECT 59.200 148.945 59.340 149.100 ;
        RECT 60.030 149.040 60.350 149.100 ;
        RECT 60.580 149.100 66.240 149.240 ;
        RECT 67.480 149.100 68.630 149.240 ;
        RECT 58.665 148.900 58.955 148.945 ;
        RECT 58.190 148.760 58.955 148.900 ;
        RECT 58.190 148.700 58.510 148.760 ;
        RECT 58.665 148.715 58.955 148.760 ;
        RECT 59.125 148.715 59.415 148.945 ;
        RECT 59.570 148.900 59.890 148.960 ;
        RECT 60.580 148.945 60.720 149.100 ;
        RECT 60.505 148.900 60.795 148.945 ;
        RECT 59.570 148.760 60.795 148.900 ;
        RECT 56.825 148.560 57.115 148.605 ;
        RECT 53.220 148.420 57.115 148.560 ;
        RECT 58.740 148.560 58.880 148.715 ;
        RECT 59.570 148.700 59.890 148.760 ;
        RECT 60.505 148.715 60.795 148.760 ;
        RECT 60.965 148.715 61.255 148.945 ;
        RECT 61.870 148.900 62.190 148.960 ;
        RECT 67.480 148.900 67.620 149.100 ;
        RECT 68.310 149.040 68.630 149.100 ;
        RECT 69.230 149.040 69.550 149.300 ;
        RECT 61.870 148.760 67.620 148.900 ;
        RECT 60.030 148.560 60.350 148.620 ;
        RECT 61.040 148.560 61.180 148.715 ;
        RECT 61.870 148.700 62.190 148.760 ;
        RECT 67.850 148.700 68.170 148.960 ;
        RECT 87.630 148.700 87.950 148.960 ;
        RECT 67.940 148.560 68.080 148.700 ;
        RECT 58.740 148.420 68.080 148.560 ;
        RECT 56.825 148.375 57.115 148.420 ;
        RECT 60.030 148.360 60.350 148.420 ;
        RECT 61.425 148.220 61.715 148.265 ;
        RECT 58.280 148.080 61.715 148.220 ;
        RECT 54.970 147.880 55.290 147.940 ;
        RECT 58.280 147.880 58.420 148.080 ;
        RECT 61.425 148.035 61.715 148.080 ;
        RECT 64.630 148.220 64.950 148.280 ;
        RECT 69.245 148.220 69.535 148.265 ;
        RECT 64.630 148.080 69.535 148.220 ;
        RECT 64.630 148.020 64.950 148.080 ;
        RECT 69.245 148.035 69.535 148.080 ;
        RECT 82.110 148.220 82.430 148.280 ;
        RECT 86.725 148.220 87.015 148.265 ;
        RECT 82.110 148.080 87.015 148.220 ;
        RECT 82.110 148.020 82.430 148.080 ;
        RECT 86.725 148.035 87.015 148.080 ;
        RECT 51.380 147.740 58.420 147.880 ;
        RECT 58.650 147.880 58.970 147.940 ;
        RECT 60.045 147.880 60.335 147.925 ;
        RECT 66.930 147.880 67.250 147.940 ;
        RECT 58.650 147.740 67.250 147.880 ;
        RECT 35.205 147.695 35.495 147.740 ;
        RECT 35.650 147.680 35.970 147.740 ;
        RECT 54.970 147.680 55.290 147.740 ;
        RECT 58.650 147.680 58.970 147.740 ;
        RECT 60.045 147.695 60.335 147.740 ;
        RECT 66.930 147.680 67.250 147.740 ;
        RECT 18.100 147.060 89.400 147.540 ;
        RECT 35.650 146.660 35.970 146.920 ;
        RECT 38.885 146.860 39.175 146.905 ;
        RECT 39.330 146.860 39.650 146.920 ;
        RECT 38.885 146.720 39.650 146.860 ;
        RECT 38.885 146.675 39.175 146.720 ;
        RECT 39.330 146.660 39.650 146.720 ;
        RECT 41.170 146.860 41.490 146.920 ;
        RECT 47.165 146.860 47.455 146.905 ;
        RECT 57.270 146.860 57.590 146.920 ;
        RECT 41.170 146.720 57.590 146.860 ;
        RECT 41.170 146.660 41.490 146.720 ;
        RECT 47.165 146.675 47.455 146.720 ;
        RECT 57.270 146.660 57.590 146.720 ;
        RECT 60.045 146.860 60.335 146.905 ;
        RECT 60.950 146.860 61.270 146.920 ;
        RECT 60.045 146.720 61.270 146.860 ;
        RECT 60.045 146.675 60.335 146.720 ;
        RECT 60.950 146.660 61.270 146.720 ;
        RECT 61.425 146.860 61.715 146.905 ;
        RECT 61.870 146.860 62.190 146.920 ;
        RECT 61.425 146.720 62.190 146.860 ;
        RECT 61.425 146.675 61.715 146.720 ;
        RECT 61.870 146.660 62.190 146.720 ;
        RECT 62.805 146.860 63.095 146.905 ;
        RECT 63.250 146.860 63.570 146.920 ;
        RECT 62.805 146.720 63.570 146.860 ;
        RECT 62.805 146.675 63.095 146.720 ;
        RECT 34.285 146.180 34.575 146.225 ;
        RECT 37.965 146.180 38.255 146.225 ;
        RECT 38.870 146.180 39.190 146.240 ;
        RECT 34.285 146.040 36.800 146.180 ;
        RECT 34.285 145.995 34.575 146.040 ;
        RECT 33.810 145.640 34.130 145.900 ;
        RECT 36.660 145.885 36.800 146.040 ;
        RECT 37.965 146.040 39.190 146.180 ;
        RECT 37.965 145.995 38.255 146.040 ;
        RECT 38.870 145.980 39.190 146.040 ;
        RECT 57.730 146.180 58.050 146.240 ;
        RECT 58.205 146.180 58.495 146.225 ;
        RECT 62.880 146.180 63.020 146.675 ;
        RECT 63.250 146.660 63.570 146.720 ;
        RECT 86.710 146.660 87.030 146.920 ;
        RECT 66.930 146.320 67.250 146.580 ;
        RECT 57.730 146.040 58.495 146.180 ;
        RECT 57.730 145.980 58.050 146.040 ;
        RECT 58.205 145.995 58.495 146.040 ;
        RECT 60.580 146.040 64.860 146.180 ;
        RECT 34.745 145.655 35.035 145.885 ;
        RECT 35.205 145.655 35.495 145.885 ;
        RECT 36.585 145.655 36.875 145.885 ;
        RECT 37.045 145.840 37.335 145.885 ;
        RECT 39.790 145.840 40.110 145.900 ;
        RECT 37.045 145.700 40.110 145.840 ;
        RECT 37.045 145.655 37.335 145.700 ;
        RECT 34.820 145.160 34.960 145.655 ;
        RECT 35.280 145.500 35.420 145.655 ;
        RECT 39.790 145.640 40.110 145.700 ;
        RECT 40.250 145.640 40.570 145.900 ;
        RECT 40.710 145.640 41.030 145.900 ;
        RECT 41.185 145.655 41.475 145.885 ;
        RECT 36.110 145.500 36.430 145.560 ;
        RECT 41.260 145.500 41.400 145.655 ;
        RECT 42.090 145.640 42.410 145.900 ;
        RECT 45.310 145.640 45.630 145.900 ;
        RECT 46.690 145.840 47.010 145.900 ;
        RECT 47.625 145.840 47.915 145.885 ;
        RECT 46.690 145.700 47.915 145.840 ;
        RECT 46.690 145.640 47.010 145.700 ;
        RECT 47.625 145.655 47.915 145.700 ;
        RECT 55.430 145.840 55.750 145.900 ;
        RECT 60.580 145.885 60.720 146.040 ;
        RECT 58.665 145.840 58.955 145.885 ;
        RECT 55.430 145.700 58.955 145.840 ;
        RECT 55.430 145.640 55.750 145.700 ;
        RECT 58.665 145.655 58.955 145.700 ;
        RECT 60.505 145.655 60.795 145.885 ;
        RECT 61.410 145.840 61.730 145.900 ;
        RECT 64.720 145.885 64.860 146.040 ;
        RECT 61.885 145.840 62.175 145.885 ;
        RECT 61.410 145.700 62.175 145.840 ;
        RECT 61.410 145.640 61.730 145.700 ;
        RECT 61.885 145.655 62.175 145.700 ;
        RECT 64.185 145.655 64.475 145.885 ;
        RECT 64.645 145.840 64.935 145.885 ;
        RECT 65.090 145.840 65.410 145.900 ;
        RECT 64.645 145.700 65.410 145.840 ;
        RECT 64.645 145.655 64.935 145.700 ;
        RECT 35.280 145.360 41.400 145.500 ;
        RECT 60.950 145.500 61.270 145.560 ;
        RECT 64.260 145.500 64.400 145.655 ;
        RECT 65.090 145.640 65.410 145.700 ;
        RECT 66.010 145.640 66.330 145.900 ;
        RECT 60.950 145.360 64.400 145.500 ;
        RECT 36.110 145.300 36.430 145.360 ;
        RECT 60.950 145.300 61.270 145.360 ;
        RECT 87.170 145.300 87.490 145.560 ;
        RECT 40.250 145.160 40.570 145.220 ;
        RECT 34.820 145.020 40.570 145.160 ;
        RECT 40.250 144.960 40.570 145.020 ;
        RECT 18.100 144.340 89.400 144.820 ;
        RECT 36.110 143.940 36.430 144.200 ;
        RECT 45.310 144.140 45.630 144.200 ;
        RECT 42.180 144.000 45.630 144.140 ;
        RECT 33.810 143.800 34.130 143.860 ;
        RECT 37.965 143.800 38.255 143.845 ;
        RECT 40.710 143.800 41.030 143.860 ;
        RECT 42.180 143.845 42.320 144.000 ;
        RECT 45.310 143.940 45.630 144.000 ;
        RECT 33.810 143.660 41.030 143.800 ;
        RECT 33.810 143.600 34.130 143.660 ;
        RECT 37.965 143.615 38.255 143.660 ;
        RECT 40.710 143.600 41.030 143.660 ;
        RECT 42.105 143.615 42.395 143.845 ;
        RECT 44.405 143.800 44.695 143.845 ;
        RECT 46.690 143.800 47.010 143.860 ;
        RECT 44.405 143.660 47.010 143.800 ;
        RECT 44.405 143.615 44.695 143.660 ;
        RECT 28.750 143.460 29.070 143.520 ;
        RECT 37.505 143.460 37.795 143.505 ;
        RECT 28.750 143.320 37.795 143.460 ;
        RECT 28.750 143.260 29.070 143.320 ;
        RECT 37.505 143.275 37.795 143.320 ;
        RECT 38.885 143.460 39.175 143.505 ;
        RECT 41.185 143.460 41.475 143.505 ;
        RECT 44.480 143.460 44.620 143.615 ;
        RECT 46.690 143.600 47.010 143.660 ;
        RECT 60.030 143.800 60.350 143.860 ;
        RECT 62.805 143.800 63.095 143.845 ;
        RECT 60.030 143.660 63.095 143.800 ;
        RECT 60.030 143.600 60.350 143.660 ;
        RECT 62.805 143.615 63.095 143.660 ;
        RECT 38.885 143.320 44.620 143.460 ;
        RECT 44.850 143.460 45.170 143.520 ;
        RECT 45.325 143.460 45.615 143.505 ;
        RECT 44.850 143.320 45.615 143.460 ;
        RECT 38.885 143.275 39.175 143.320 ;
        RECT 41.185 143.275 41.475 143.320 ;
        RECT 35.650 143.120 35.970 143.180 ;
        RECT 36.125 143.120 36.415 143.165 ;
        RECT 35.650 142.980 36.415 143.120 ;
        RECT 37.580 143.120 37.720 143.275 ;
        RECT 44.850 143.260 45.170 143.320 ;
        RECT 45.325 143.275 45.615 143.320 ;
        RECT 46.245 143.460 46.535 143.505 ;
        RECT 49.450 143.460 49.770 143.520 ;
        RECT 46.245 143.320 49.770 143.460 ;
        RECT 46.245 143.275 46.535 143.320 ;
        RECT 49.450 143.260 49.770 143.320 ;
        RECT 63.725 143.275 64.015 143.505 ;
        RECT 39.805 143.120 40.095 143.165 ;
        RECT 60.950 143.120 61.270 143.180 ;
        RECT 63.800 143.120 63.940 143.275 ;
        RECT 65.090 143.260 65.410 143.520 ;
        RECT 66.010 143.260 66.330 143.520 ;
        RECT 37.580 142.980 63.940 143.120 ;
        RECT 35.650 142.920 35.970 142.980 ;
        RECT 36.125 142.935 36.415 142.980 ;
        RECT 39.805 142.935 40.095 142.980 ;
        RECT 36.200 142.780 36.340 142.935 ;
        RECT 60.950 142.920 61.270 142.980 ;
        RECT 87.630 142.920 87.950 143.180 ;
        RECT 43.025 142.780 43.315 142.825 ;
        RECT 57.730 142.780 58.050 142.840 ;
        RECT 36.200 142.640 43.315 142.780 ;
        RECT 43.025 142.595 43.315 142.640 ;
        RECT 46.780 142.640 58.050 142.780 ;
        RECT 37.045 142.440 37.335 142.485 ;
        RECT 42.550 142.440 42.870 142.500 ;
        RECT 46.780 142.440 46.920 142.640 ;
        RECT 57.730 142.580 58.050 142.640 ;
        RECT 37.045 142.300 46.920 142.440 ;
        RECT 47.165 142.440 47.455 142.485 ;
        RECT 48.530 142.440 48.850 142.500 ;
        RECT 47.165 142.300 48.850 142.440 ;
        RECT 37.045 142.255 37.335 142.300 ;
        RECT 42.550 142.240 42.870 142.300 ;
        RECT 47.165 142.255 47.455 142.300 ;
        RECT 48.530 142.240 48.850 142.300 ;
        RECT 18.100 141.620 89.400 142.100 ;
        RECT 35.665 141.420 35.955 141.465 ;
        RECT 36.570 141.420 36.890 141.480 ;
        RECT 35.665 141.280 36.890 141.420 ;
        RECT 35.665 141.235 35.955 141.280 ;
        RECT 36.570 141.220 36.890 141.280 ;
        RECT 40.250 141.420 40.570 141.480 ;
        RECT 41.185 141.420 41.475 141.465 ;
        RECT 40.250 141.280 41.475 141.420 ;
        RECT 40.250 141.220 40.570 141.280 ;
        RECT 41.185 141.235 41.475 141.280 ;
        RECT 43.025 141.420 43.315 141.465 ;
        RECT 44.850 141.420 45.170 141.480 ;
        RECT 43.025 141.280 45.170 141.420 ;
        RECT 43.025 141.235 43.315 141.280 ;
        RECT 44.850 141.220 45.170 141.280 ;
        RECT 45.310 141.420 45.630 141.480 ;
        RECT 46.245 141.420 46.535 141.465 ;
        RECT 45.310 141.280 46.535 141.420 ;
        RECT 45.310 141.220 45.630 141.280 ;
        RECT 46.245 141.235 46.535 141.280 ;
        RECT 39.805 141.080 40.095 141.125 ;
        RECT 43.930 141.080 44.250 141.140 ;
        RECT 39.805 140.940 44.250 141.080 ;
        RECT 39.805 140.895 40.095 140.940 ;
        RECT 43.930 140.880 44.250 140.940 ;
        RECT 42.550 140.740 42.870 140.800 ;
        RECT 40.800 140.600 42.870 140.740 ;
        RECT 25.530 140.400 25.850 140.460 ;
        RECT 26.005 140.400 26.295 140.445 ;
        RECT 25.530 140.260 26.295 140.400 ;
        RECT 25.530 140.200 25.850 140.260 ;
        RECT 26.005 140.215 26.295 140.260 ;
        RECT 35.190 140.400 35.510 140.460 ;
        RECT 36.585 140.400 36.875 140.445 ;
        RECT 35.190 140.260 36.875 140.400 ;
        RECT 35.190 140.200 35.510 140.260 ;
        RECT 36.585 140.215 36.875 140.260 ;
        RECT 38.870 140.200 39.190 140.460 ;
        RECT 40.800 140.445 40.940 140.600 ;
        RECT 42.550 140.540 42.870 140.600 ;
        RECT 40.725 140.215 41.015 140.445 ;
        RECT 41.645 140.215 41.935 140.445 ;
        RECT 41.720 140.060 41.860 140.215 ;
        RECT 42.090 140.200 42.410 140.460 ;
        RECT 45.310 140.400 45.630 140.460 ;
        RECT 42.640 140.260 45.630 140.400 ;
        RECT 42.640 140.060 42.780 140.260 ;
        RECT 45.310 140.200 45.630 140.260 ;
        RECT 48.530 140.200 48.850 140.460 ;
        RECT 41.720 139.920 42.780 140.060 ;
        RECT 44.850 140.060 45.170 140.120 ;
        RECT 45.785 140.060 46.075 140.105 ;
        RECT 44.850 139.920 46.075 140.060 ;
        RECT 44.850 139.860 45.170 139.920 ;
        RECT 45.785 139.875 46.075 139.920 ;
        RECT 48.070 139.720 48.390 139.780 ;
        RECT 49.465 139.720 49.755 139.765 ;
        RECT 48.070 139.580 49.755 139.720 ;
        RECT 48.070 139.520 48.390 139.580 ;
        RECT 49.465 139.535 49.755 139.580 ;
        RECT 18.100 138.900 89.400 139.380 ;
      LAYER met2 ;
        RECT 12.670 217.330 12.950 221.330 ;
        RECT 15.890 217.330 16.170 221.330 ;
        RECT 19.110 217.330 19.390 221.330 ;
        RECT 22.330 217.330 22.610 221.330 ;
        RECT 25.550 217.330 25.830 221.330 ;
        RECT 28.770 217.330 29.050 221.330 ;
        RECT 31.990 217.330 32.270 221.330 ;
        RECT 35.210 217.330 35.490 221.330 ;
        RECT 38.430 217.330 38.710 221.330 ;
        RECT 38.960 217.610 40.480 217.750 ;
        RECT 12.740 214.465 12.880 217.330 ;
        RECT 12.670 214.095 12.950 214.465 ;
        RECT 15.960 181.145 16.100 217.330 ;
        RECT 16.820 211.230 17.080 211.550 ;
        RECT 16.880 191.910 17.020 211.230 ;
        RECT 17.730 210.015 18.010 210.385 ;
        RECT 17.800 206.790 17.940 210.015 ;
        RECT 19.180 208.230 19.320 217.330 ;
        RECT 21.880 213.950 22.140 214.270 ;
        RECT 19.580 211.910 19.840 212.230 ;
        RECT 18.720 208.090 19.320 208.230 ;
        RECT 17.740 206.470 18.000 206.790 ;
        RECT 17.280 205.110 17.540 205.430 ;
        RECT 17.340 198.030 17.480 205.110 ;
        RECT 18.200 204.770 18.460 205.090 ;
        RECT 17.740 200.690 18.000 201.010 ;
        RECT 17.800 200.185 17.940 200.690 ;
        RECT 17.730 199.815 18.010 200.185 ;
        RECT 17.340 197.890 17.940 198.030 ;
        RECT 17.270 193.015 17.550 193.385 ;
        RECT 17.340 192.850 17.480 193.015 ;
        RECT 17.280 192.530 17.540 192.850 ;
        RECT 16.880 191.770 17.480 191.910 ;
        RECT 16.820 191.170 17.080 191.490 ;
        RECT 16.880 190.665 17.020 191.170 ;
        RECT 16.810 190.295 17.090 190.665 ;
        RECT 16.810 187.575 17.090 187.945 ;
        RECT 16.820 187.430 17.080 187.575 ;
        RECT 15.890 180.775 16.170 181.145 ;
        RECT 17.340 175.850 17.480 191.770 ;
        RECT 17.800 176.530 17.940 197.890 ;
        RECT 18.260 181.630 18.400 204.770 ;
        RECT 18.720 204.070 18.860 208.090 ;
        RECT 19.110 206.615 19.390 206.985 ;
        RECT 18.660 203.750 18.920 204.070 ;
        RECT 18.650 203.215 18.930 203.585 ;
        RECT 18.720 182.310 18.860 203.215 ;
        RECT 18.660 181.990 18.920 182.310 ;
        RECT 18.200 181.310 18.460 181.630 ;
        RECT 19.180 180.950 19.320 206.615 ;
        RECT 19.640 190.130 19.780 211.910 ;
        RECT 20.950 210.695 21.230 211.065 ;
        RECT 21.020 208.830 21.160 210.695 ;
        RECT 21.940 209.510 22.080 213.950 ;
        RECT 22.400 211.550 22.540 217.330 ;
        RECT 22.790 216.815 23.070 217.185 ;
        RECT 22.340 211.230 22.600 211.550 ;
        RECT 21.880 209.190 22.140 209.510 ;
        RECT 20.960 208.510 21.220 208.830 ;
        RECT 21.880 206.130 22.140 206.450 ;
        RECT 21.420 205.625 21.680 205.770 ;
        RECT 21.410 205.255 21.690 205.625 ;
        RECT 21.420 204.770 21.680 205.090 ;
        RECT 21.480 203.390 21.620 204.770 ;
        RECT 21.940 204.070 22.080 206.130 ;
        RECT 21.880 203.750 22.140 204.070 ;
        RECT 20.500 203.070 20.760 203.390 ;
        RECT 21.420 203.070 21.680 203.390 ;
        RECT 20.040 196.785 20.300 196.930 ;
        RECT 20.030 196.415 20.310 196.785 ;
        RECT 20.040 191.850 20.300 192.170 ;
        RECT 19.580 189.810 19.840 190.130 ;
        RECT 19.580 183.690 19.840 184.010 ;
        RECT 19.640 183.185 19.780 183.690 ;
        RECT 19.570 182.815 19.850 183.185 ;
        RECT 19.120 180.630 19.380 180.950 ;
        RECT 17.740 176.210 18.000 176.530 ;
        RECT 19.570 176.015 19.850 176.385 ;
        RECT 19.580 175.870 19.840 176.015 ;
        RECT 17.280 175.530 17.540 175.850 ;
        RECT 20.100 173.470 20.240 191.850 ;
        RECT 20.560 180.610 20.700 203.070 ;
        RECT 21.880 200.010 22.140 200.330 ;
        RECT 20.960 197.630 21.220 197.950 ;
        RECT 21.020 193.190 21.160 197.630 ;
        RECT 21.940 194.890 22.080 200.010 ;
        RECT 22.340 199.330 22.600 199.650 ;
        RECT 22.400 195.230 22.540 199.330 ;
        RECT 22.860 198.630 23.000 216.815 ;
        RECT 24.640 212.930 24.900 213.250 ;
        RECT 24.180 210.210 24.440 210.530 ;
        RECT 23.250 209.335 23.530 209.705 ;
        RECT 23.320 198.630 23.460 209.335 ;
        RECT 24.240 203.390 24.380 210.210 ;
        RECT 23.720 203.070 23.980 203.390 ;
        RECT 24.180 203.070 24.440 203.390 ;
        RECT 23.780 201.545 23.920 203.070 ;
        RECT 23.710 201.175 23.990 201.545 ;
        RECT 24.700 201.350 24.840 212.930 ;
        RECT 25.100 212.250 25.360 212.570 ;
        RECT 25.160 209.510 25.300 212.250 ;
        RECT 25.620 211.745 25.760 217.330 ;
        RECT 26.480 212.590 26.740 212.910 ;
        RECT 25.550 211.375 25.830 211.745 ;
        RECT 25.100 209.190 25.360 209.510 ;
        RECT 26.540 209.170 26.680 212.590 ;
        RECT 26.480 208.850 26.740 209.170 ;
        RECT 26.020 208.510 26.280 208.830 ;
        RECT 26.080 208.345 26.220 208.510 ;
        RECT 26.010 207.975 26.290 208.345 ;
        RECT 25.560 206.130 25.820 206.450 ;
        RECT 25.620 205.090 25.760 206.130 ;
        RECT 26.540 205.770 26.680 208.850 ;
        RECT 27.400 208.510 27.660 208.830 ;
        RECT 26.940 206.470 27.200 206.790 ;
        RECT 26.480 205.450 26.740 205.770 ;
        RECT 25.560 204.770 25.820 205.090 ;
        RECT 26.010 204.575 26.290 204.945 ;
        RECT 25.550 203.895 25.830 204.265 ;
        RECT 26.080 204.070 26.220 204.575 ;
        RECT 24.640 201.030 24.900 201.350 ;
        RECT 25.620 200.330 25.760 203.895 ;
        RECT 26.020 203.750 26.280 204.070 ;
        RECT 26.480 203.070 26.740 203.390 ;
        RECT 26.020 202.050 26.280 202.370 ;
        RECT 23.720 200.010 23.980 200.330 ;
        RECT 25.100 200.185 25.360 200.330 ;
        RECT 22.800 198.310 23.060 198.630 ;
        RECT 23.260 198.310 23.520 198.630 ;
        RECT 22.340 194.910 22.600 195.230 ;
        RECT 21.880 194.570 22.140 194.890 ;
        RECT 21.420 194.230 21.680 194.550 ;
        RECT 20.960 192.870 21.220 193.190 ;
        RECT 20.960 192.190 21.220 192.510 ;
        RECT 21.020 189.450 21.160 192.190 ;
        RECT 21.480 191.490 21.620 194.230 ;
        RECT 21.420 191.170 21.680 191.490 ;
        RECT 20.960 189.130 21.220 189.450 ;
        RECT 20.960 188.450 21.220 188.770 ;
        RECT 21.020 187.070 21.160 188.450 ;
        RECT 20.960 186.750 21.220 187.070 ;
        RECT 20.960 181.650 21.220 181.970 ;
        RECT 20.500 180.290 20.760 180.610 ;
        RECT 21.020 179.670 21.160 181.650 ;
        RECT 21.480 181.200 21.620 191.170 ;
        RECT 21.940 185.030 22.080 194.570 ;
        RECT 22.400 189.870 22.540 194.910 ;
        RECT 22.800 194.230 23.060 194.550 ;
        RECT 22.860 191.490 23.000 194.230 ;
        RECT 23.260 192.870 23.520 193.190 ;
        RECT 22.800 191.170 23.060 191.490 ;
        RECT 22.400 189.730 23.000 189.870 ;
        RECT 22.340 189.130 22.600 189.450 ;
        RECT 21.880 184.710 22.140 185.030 ;
        RECT 21.880 181.200 22.140 181.290 ;
        RECT 21.480 181.060 22.140 181.200 ;
        RECT 21.880 180.970 22.140 181.060 ;
        RECT 20.560 179.530 21.160 179.670 ;
        RECT 20.560 175.170 20.700 179.530 ;
        RECT 22.400 178.570 22.540 189.130 ;
        RECT 22.860 187.945 23.000 189.730 ;
        RECT 23.320 189.450 23.460 192.870 ;
        RECT 23.780 190.470 23.920 200.010 ;
        RECT 25.090 199.815 25.370 200.185 ;
        RECT 25.560 200.010 25.820 200.330 ;
        RECT 25.560 199.330 25.820 199.650 ;
        RECT 24.640 197.970 24.900 198.290 ;
        RECT 24.180 197.290 24.440 197.610 ;
        RECT 23.720 190.150 23.980 190.470 ;
        RECT 23.260 189.130 23.520 189.450 ;
        RECT 22.790 187.575 23.070 187.945 ;
        RECT 24.240 187.750 24.380 197.290 ;
        RECT 24.700 194.800 24.840 197.970 ;
        RECT 25.620 197.950 25.760 199.330 ;
        RECT 25.100 197.630 25.360 197.950 ;
        RECT 25.560 197.630 25.820 197.950 ;
        RECT 25.160 195.910 25.300 197.630 ;
        RECT 25.100 195.590 25.360 195.910 ;
        RECT 25.620 195.570 25.760 197.630 ;
        RECT 25.560 195.250 25.820 195.570 ;
        RECT 25.100 194.800 25.360 194.890 ;
        RECT 24.700 194.660 25.360 194.800 ;
        RECT 25.100 194.570 25.360 194.660 ;
        RECT 24.630 193.695 24.910 194.065 ;
        RECT 24.700 192.510 24.840 193.695 ;
        RECT 24.640 192.190 24.900 192.510 ;
        RECT 25.160 192.080 25.300 194.570 ;
        RECT 25.550 193.015 25.830 193.385 ;
        RECT 25.560 192.870 25.820 193.015 ;
        RECT 25.560 192.080 25.820 192.170 ;
        RECT 25.160 191.940 25.820 192.080 ;
        RECT 25.160 189.790 25.300 191.940 ;
        RECT 25.560 191.850 25.820 191.940 ;
        RECT 26.080 191.910 26.220 202.050 ;
        RECT 26.540 201.545 26.680 203.070 ;
        RECT 26.470 201.175 26.750 201.545 ;
        RECT 26.480 199.670 26.740 199.990 ;
        RECT 26.540 199.505 26.680 199.670 ;
        RECT 27.000 199.650 27.140 206.470 ;
        RECT 27.460 205.430 27.600 208.510 ;
        RECT 28.320 207.490 28.580 207.810 ;
        RECT 28.380 206.305 28.520 207.490 ;
        RECT 28.310 205.935 28.590 206.305 ;
        RECT 28.320 205.450 28.580 205.770 ;
        RECT 27.400 205.110 27.660 205.430 ;
        RECT 27.860 205.110 28.120 205.430 ;
        RECT 27.460 203.050 27.600 205.110 ;
        RECT 27.920 204.070 28.060 205.110 ;
        RECT 27.860 203.750 28.120 204.070 ;
        RECT 27.850 203.215 28.130 203.585 ;
        RECT 28.380 203.390 28.520 205.450 ;
        RECT 27.860 203.070 28.120 203.215 ;
        RECT 28.320 203.070 28.580 203.390 ;
        RECT 27.400 202.730 27.660 203.050 ;
        RECT 28.380 202.790 28.520 203.070 ;
        RECT 27.920 202.650 28.520 202.790 ;
        RECT 27.390 201.855 27.670 202.225 ;
        RECT 27.460 199.650 27.600 201.855 ;
        RECT 26.470 199.135 26.750 199.505 ;
        RECT 26.940 199.330 27.200 199.650 ;
        RECT 27.400 199.330 27.660 199.650 ;
        RECT 27.920 198.825 28.060 202.650 ;
        RECT 28.320 202.050 28.580 202.370 ;
        RECT 27.850 198.455 28.130 198.825 ;
        RECT 27.400 198.200 27.660 198.290 ;
        RECT 27.400 198.060 28.060 198.200 ;
        RECT 27.400 197.970 27.660 198.060 ;
        RECT 26.480 197.630 26.740 197.950 ;
        RECT 26.540 195.230 26.680 197.630 ;
        RECT 27.400 197.290 27.660 197.610 ;
        RECT 26.930 195.735 27.210 196.105 ;
        RECT 26.480 194.910 26.740 195.230 ;
        RECT 27.000 194.210 27.140 195.735 ;
        RECT 27.460 194.890 27.600 197.290 ;
        RECT 27.920 196.105 28.060 198.060 ;
        RECT 28.380 197.610 28.520 202.050 ;
        RECT 28.320 197.290 28.580 197.610 ;
        RECT 27.850 195.735 28.130 196.105 ;
        RECT 27.400 194.800 27.660 194.890 ;
        RECT 27.400 194.660 28.060 194.800 ;
        RECT 27.400 194.570 27.660 194.660 ;
        RECT 26.940 193.890 27.200 194.210 ;
        RECT 27.400 193.890 27.660 194.210 ;
        RECT 27.460 192.510 27.600 193.890 ;
        RECT 27.920 193.190 28.060 194.660 ;
        RECT 28.320 194.570 28.580 194.890 ;
        RECT 28.840 194.745 28.980 217.330 ;
        RECT 31.530 212.055 31.810 212.425 ;
        RECT 32.060 212.230 32.200 217.330 ;
        RECT 32.460 212.590 32.720 212.910 ;
        RECT 30.150 211.375 30.430 211.745 ;
        RECT 29.700 210.890 29.960 211.210 ;
        RECT 29.240 209.190 29.500 209.510 ;
        RECT 29.300 206.790 29.440 209.190 ;
        RECT 29.760 208.830 29.900 210.890 ;
        RECT 29.700 208.510 29.960 208.830 ;
        RECT 30.220 207.810 30.360 211.375 ;
        RECT 31.080 210.550 31.340 210.870 ;
        RECT 30.610 208.655 30.890 209.025 ;
        RECT 30.620 208.510 30.880 208.655 ;
        RECT 31.140 208.490 31.280 210.550 ;
        RECT 31.080 208.170 31.340 208.490 ;
        RECT 31.600 208.150 31.740 212.055 ;
        RECT 32.000 211.910 32.260 212.230 ;
        RECT 32.000 208.170 32.260 208.490 ;
        RECT 31.540 207.830 31.800 208.150 ;
        RECT 30.160 207.490 30.420 207.810 ;
        RECT 30.620 207.490 30.880 207.810 ;
        RECT 29.240 206.470 29.500 206.790 ;
        RECT 29.700 206.130 29.960 206.450 ;
        RECT 29.230 205.255 29.510 205.625 ;
        RECT 29.300 195.910 29.440 205.255 ;
        RECT 29.760 202.370 29.900 206.130 ;
        RECT 30.680 206.110 30.820 207.490 ;
        RECT 31.540 206.470 31.800 206.790 ;
        RECT 30.620 205.790 30.880 206.110 ;
        RECT 30.160 205.450 30.420 205.770 ;
        RECT 30.220 204.945 30.360 205.450 ;
        RECT 30.150 204.575 30.430 204.945 ;
        RECT 31.080 204.770 31.340 205.090 ;
        RECT 30.620 203.585 30.880 203.730 ;
        RECT 30.610 203.215 30.890 203.585 ;
        RECT 31.140 203.390 31.280 204.770 ;
        RECT 31.080 203.070 31.340 203.390 ;
        RECT 30.160 202.390 30.420 202.710 ;
        RECT 29.700 202.050 29.960 202.370 ;
        RECT 29.700 200.350 29.960 200.670 ;
        RECT 29.240 195.590 29.500 195.910 ;
        RECT 27.860 192.870 28.120 193.190 ;
        RECT 27.400 192.190 27.660 192.510 ;
        RECT 26.080 191.770 27.140 191.910 ;
        RECT 26.480 191.170 26.740 191.490 ;
        RECT 26.020 190.040 26.280 190.130 ;
        RECT 25.620 189.900 26.280 190.040 ;
        RECT 25.100 189.470 25.360 189.790 ;
        RECT 25.090 188.935 25.370 189.305 ;
        RECT 24.640 188.450 24.900 188.770 ;
        RECT 24.180 187.430 24.440 187.750 ;
        RECT 23.720 187.320 23.980 187.410 ;
        RECT 22.860 187.180 23.980 187.320 ;
        RECT 22.860 184.010 23.000 187.180 ;
        RECT 23.720 187.090 23.980 187.180 ;
        RECT 24.240 187.070 24.380 187.430 ;
        RECT 24.700 187.070 24.840 188.450 ;
        RECT 24.180 186.750 24.440 187.070 ;
        RECT 24.640 186.750 24.900 187.070 ;
        RECT 24.240 184.690 24.380 186.750 ;
        RECT 24.180 184.370 24.440 184.690 ;
        RECT 22.800 183.920 23.060 184.010 ;
        RECT 22.800 183.780 23.460 183.920 ;
        RECT 22.800 183.690 23.060 183.780 ;
        RECT 22.790 181.455 23.070 181.825 ;
        RECT 22.800 181.310 23.060 181.455 ;
        RECT 23.320 179.590 23.460 183.780 ;
        RECT 24.240 183.670 24.380 184.370 ;
        RECT 24.700 184.010 24.840 186.750 ;
        RECT 25.160 186.730 25.300 188.935 ;
        RECT 25.100 186.410 25.360 186.730 ;
        RECT 25.620 186.390 25.760 189.900 ;
        RECT 26.020 189.810 26.280 189.900 ;
        RECT 26.540 189.110 26.680 191.170 ;
        RECT 26.480 189.020 26.740 189.110 ;
        RECT 26.080 188.880 26.740 189.020 ;
        RECT 26.080 187.750 26.220 188.880 ;
        RECT 26.480 188.790 26.740 188.880 ;
        RECT 26.020 187.430 26.280 187.750 ;
        RECT 26.470 187.575 26.750 187.945 ;
        RECT 25.560 186.070 25.820 186.390 ;
        RECT 25.620 184.350 25.760 186.070 ;
        RECT 25.560 184.030 25.820 184.350 ;
        RECT 24.640 183.690 24.900 184.010 ;
        RECT 24.180 183.350 24.440 183.670 ;
        RECT 24.700 182.310 24.840 183.690 ;
        RECT 26.080 183.330 26.220 187.430 ;
        RECT 26.540 186.730 26.680 187.575 ;
        RECT 26.480 186.410 26.740 186.730 ;
        RECT 26.020 183.010 26.280 183.330 ;
        RECT 24.640 181.990 24.900 182.310 ;
        RECT 26.010 182.135 26.290 182.505 ;
        RECT 23.260 179.270 23.520 179.590 ;
        RECT 22.340 178.250 22.600 178.570 ;
        RECT 21.880 177.570 22.140 177.890 ;
        RECT 22.340 177.570 22.600 177.890 ;
        RECT 21.940 176.190 22.080 177.570 ;
        RECT 21.880 175.870 22.140 176.190 ;
        RECT 20.500 174.850 20.760 175.170 ;
        RECT 20.040 173.150 20.300 173.470 ;
        RECT 20.560 170.265 20.700 174.850 ;
        RECT 21.420 172.810 21.680 173.130 ;
        RECT 20.490 169.895 20.770 170.265 ;
        RECT 21.480 168.710 21.620 172.810 ;
        RECT 21.420 168.390 21.680 168.710 ;
        RECT 21.420 166.690 21.680 167.010 ;
        RECT 20.030 159.015 20.310 159.385 ;
        RECT 20.040 158.870 20.300 159.015 ;
        RECT 21.480 157.830 21.620 166.690 ;
        RECT 22.400 165.990 22.540 177.570 ;
        RECT 22.800 173.150 23.060 173.470 ;
        RECT 22.860 171.430 23.000 173.150 ;
        RECT 22.800 171.110 23.060 171.430 ;
        RECT 23.320 170.830 23.460 179.270 ;
        RECT 24.700 178.230 24.840 181.990 ;
        RECT 26.080 181.630 26.220 182.135 ;
        RECT 25.100 181.310 25.360 181.630 ;
        RECT 26.020 181.310 26.280 181.630 ;
        RECT 25.160 180.610 25.300 181.310 ;
        RECT 25.100 180.290 25.360 180.610 ;
        RECT 26.080 178.570 26.220 181.310 ;
        RECT 26.540 181.030 26.680 186.410 ;
        RECT 27.000 181.630 27.140 191.770 ;
        RECT 28.380 191.490 28.520 194.570 ;
        RECT 28.770 194.375 29.050 194.745 ;
        RECT 29.240 194.230 29.500 194.550 ;
        RECT 28.780 192.190 29.040 192.510 ;
        RECT 28.840 191.830 28.980 192.190 ;
        RECT 28.780 191.510 29.040 191.830 ;
        RECT 28.320 191.170 28.580 191.490 ;
        RECT 28.840 189.985 28.980 191.510 ;
        RECT 29.300 190.470 29.440 194.230 ;
        RECT 29.240 190.150 29.500 190.470 ;
        RECT 28.770 189.615 29.050 189.985 ;
        RECT 28.780 189.360 29.040 189.450 ;
        RECT 29.300 189.360 29.440 190.150 ;
        RECT 29.760 189.700 29.900 200.350 ;
        RECT 30.220 190.665 30.360 202.390 ;
        RECT 30.620 202.050 30.880 202.370 ;
        RECT 31.080 202.050 31.340 202.370 ;
        RECT 30.680 195.910 30.820 202.050 ;
        RECT 30.620 195.590 30.880 195.910 ;
        RECT 30.610 195.055 30.890 195.425 ;
        RECT 30.680 194.890 30.820 195.055 ;
        RECT 30.620 194.570 30.880 194.890 ;
        RECT 30.620 193.890 30.880 194.210 ;
        RECT 30.680 192.850 30.820 193.890 ;
        RECT 30.620 192.530 30.880 192.850 ;
        RECT 30.150 190.295 30.430 190.665 ;
        RECT 29.760 189.560 30.820 189.700 ;
        RECT 28.780 189.220 29.440 189.360 ;
        RECT 28.780 189.130 29.040 189.220 ;
        RECT 28.320 188.450 28.580 188.770 ;
        RECT 28.380 187.070 28.520 188.450 ;
        RECT 28.320 186.750 28.580 187.070 ;
        RECT 27.860 185.730 28.120 186.050 ;
        RECT 27.920 184.690 28.060 185.730 ;
        RECT 27.400 184.545 27.660 184.690 ;
        RECT 27.390 184.175 27.670 184.545 ;
        RECT 27.860 184.370 28.120 184.690 ;
        RECT 28.380 184.350 28.520 186.750 ;
        RECT 28.320 184.030 28.580 184.350 ;
        RECT 27.850 183.495 28.130 183.865 ;
        RECT 27.920 182.310 28.060 183.495 ;
        RECT 28.320 183.010 28.580 183.330 ;
        RECT 27.860 181.990 28.120 182.310 ;
        RECT 26.940 181.310 27.200 181.630 ;
        RECT 27.860 181.310 28.120 181.630 ;
        RECT 27.920 181.145 28.060 181.310 ;
        RECT 26.540 180.890 27.140 181.030 ;
        RECT 26.480 180.290 26.740 180.610 ;
        RECT 26.540 179.250 26.680 180.290 ;
        RECT 27.000 179.590 27.140 180.890 ;
        RECT 27.850 180.775 28.130 181.145 ;
        RECT 27.850 180.095 28.130 180.465 ;
        RECT 26.940 179.270 27.200 179.590 ;
        RECT 26.480 178.930 26.740 179.250 ;
        RECT 27.400 178.930 27.660 179.250 ;
        RECT 26.940 178.590 27.200 178.910 ;
        RECT 26.020 178.250 26.280 178.570 ;
        RECT 24.640 177.910 24.900 178.230 ;
        RECT 26.080 176.630 26.220 178.250 ;
        RECT 25.620 176.490 26.220 176.630 ;
        RECT 24.640 175.870 24.900 176.190 ;
        RECT 25.100 175.870 25.360 176.190 ;
        RECT 23.720 175.190 23.980 175.510 ;
        RECT 23.780 171.430 23.920 175.190 ;
        RECT 24.700 175.170 24.840 175.870 ;
        RECT 24.640 174.850 24.900 175.170 ;
        RECT 24.700 173.470 24.840 174.850 ;
        RECT 24.640 173.150 24.900 173.470 ;
        RECT 23.720 171.110 23.980 171.430 ;
        RECT 22.860 170.690 23.460 170.830 ;
        RECT 22.340 165.670 22.600 165.990 ;
        RECT 22.400 162.250 22.540 165.670 ;
        RECT 22.340 161.930 22.600 162.250 ;
        RECT 22.860 160.550 23.000 170.690 ;
        RECT 23.780 168.030 23.920 171.110 ;
        RECT 24.180 170.090 24.440 170.410 ;
        RECT 24.640 170.090 24.900 170.410 ;
        RECT 23.720 167.710 23.980 168.030 ;
        RECT 23.260 167.370 23.520 167.690 ;
        RECT 23.320 164.970 23.460 167.370 ;
        RECT 24.240 167.010 24.380 170.090 ;
        RECT 24.700 168.030 24.840 170.090 ;
        RECT 24.640 167.710 24.900 168.030 ;
        RECT 24.180 166.690 24.440 167.010 ;
        RECT 23.720 164.990 23.980 165.310 ;
        RECT 23.260 164.650 23.520 164.970 ;
        RECT 23.320 162.590 23.460 164.650 ;
        RECT 23.260 162.270 23.520 162.590 ;
        RECT 23.780 161.570 23.920 164.990 ;
        RECT 23.720 161.250 23.980 161.570 ;
        RECT 22.800 160.230 23.060 160.550 ;
        RECT 21.880 159.550 22.140 159.870 ;
        RECT 21.420 157.510 21.680 157.830 ;
        RECT 21.940 155.985 22.080 159.550 ;
        RECT 22.340 158.530 22.600 158.850 ;
        RECT 22.400 157.490 22.540 158.530 ;
        RECT 23.780 157.830 23.920 161.250 ;
        RECT 24.640 160.230 24.900 160.550 ;
        RECT 23.720 157.510 23.980 157.830 ;
        RECT 22.340 157.170 22.600 157.490 ;
        RECT 24.700 157.150 24.840 160.230 ;
        RECT 24.640 156.830 24.900 157.150 ;
        RECT 21.870 155.615 22.150 155.985 ;
        RECT 19.580 153.770 19.840 154.090 ;
        RECT 19.640 153.265 19.780 153.770 ;
        RECT 19.570 152.895 19.850 153.265 ;
        RECT 25.160 152.390 25.300 175.870 ;
        RECT 25.620 155.110 25.760 176.490 ;
        RECT 27.000 176.190 27.140 178.590 ;
        RECT 26.940 175.870 27.200 176.190 ;
        RECT 27.460 165.505 27.600 178.930 ;
        RECT 27.920 173.550 28.060 180.095 ;
        RECT 28.380 179.250 28.520 183.010 ;
        RECT 28.320 178.930 28.580 179.250 ;
        RECT 28.310 178.055 28.590 178.425 ;
        RECT 28.380 175.510 28.520 178.055 ;
        RECT 28.320 175.190 28.580 175.510 ;
        RECT 27.920 173.410 28.520 173.550 ;
        RECT 27.860 172.810 28.120 173.130 ;
        RECT 27.920 171.090 28.060 172.810 ;
        RECT 27.860 170.770 28.120 171.090 ;
        RECT 27.390 165.135 27.670 165.505 ;
        RECT 27.920 165.310 28.060 170.770 ;
        RECT 28.380 166.070 28.520 173.410 ;
        RECT 28.840 173.130 28.980 189.130 ;
        RECT 30.160 188.790 30.420 189.110 ;
        RECT 29.240 188.450 29.500 188.770 ;
        RECT 29.300 185.030 29.440 188.450 ;
        RECT 30.220 187.660 30.360 188.790 ;
        RECT 29.760 187.520 30.360 187.660 ;
        RECT 29.240 184.710 29.500 185.030 ;
        RECT 29.760 183.330 29.900 187.520 ;
        RECT 30.680 187.070 30.820 189.560 ;
        RECT 30.160 186.750 30.420 187.070 ;
        RECT 30.620 186.750 30.880 187.070 ;
        RECT 30.220 184.545 30.360 186.750 ;
        RECT 30.150 184.175 30.430 184.545 ;
        RECT 29.230 182.815 29.510 183.185 ;
        RECT 29.700 183.010 29.960 183.330 ;
        RECT 29.300 181.630 29.440 182.815 ;
        RECT 29.240 181.310 29.500 181.630 ;
        RECT 29.240 180.290 29.500 180.610 ;
        RECT 29.300 179.590 29.440 180.290 ;
        RECT 29.240 179.270 29.500 179.590 ;
        RECT 29.300 177.890 29.440 179.270 ;
        RECT 29.240 177.570 29.500 177.890 ;
        RECT 28.780 173.040 29.040 173.130 ;
        RECT 28.780 172.900 29.440 173.040 ;
        RECT 28.780 172.810 29.040 172.900 ;
        RECT 28.780 172.130 29.040 172.450 ;
        RECT 28.840 170.750 28.980 172.130 ;
        RECT 29.300 170.750 29.440 172.900 ;
        RECT 29.760 171.510 29.900 183.010 ;
        RECT 30.150 182.135 30.430 182.505 ;
        RECT 30.680 182.310 30.820 186.750 ;
        RECT 31.140 184.690 31.280 202.050 ;
        RECT 31.600 201.010 31.740 206.470 ;
        RECT 32.060 203.050 32.200 208.170 ;
        RECT 32.000 202.730 32.260 203.050 ;
        RECT 31.990 201.175 32.270 201.545 ;
        RECT 31.540 200.690 31.800 201.010 ;
        RECT 32.060 200.670 32.200 201.175 ;
        RECT 32.000 200.350 32.260 200.670 ;
        RECT 31.540 199.670 31.800 199.990 ;
        RECT 31.600 198.290 31.740 199.670 ;
        RECT 32.060 198.630 32.200 200.350 ;
        RECT 32.520 200.330 32.660 212.590 ;
        RECT 35.280 211.550 35.420 217.330 ;
        RECT 38.500 217.070 38.640 217.330 ;
        RECT 38.960 217.070 39.100 217.610 ;
        RECT 38.500 216.930 39.100 217.070 ;
        RECT 36.600 211.910 36.860 212.230 ;
        RECT 35.220 211.230 35.480 211.550 ;
        RECT 35.210 209.335 35.490 209.705 ;
        RECT 35.280 208.490 35.420 209.335 ;
        RECT 36.660 208.830 36.800 211.910 ;
        RECT 39.810 210.695 40.090 211.065 ;
        RECT 36.950 209.675 38.490 210.045 ;
        RECT 38.890 209.420 39.170 209.705 ;
        RECT 37.580 209.335 39.170 209.420 ;
        RECT 37.580 209.280 39.100 209.335 ;
        RECT 37.060 208.850 37.320 209.170 ;
        RECT 36.600 208.510 36.860 208.830 ;
        RECT 33.840 208.345 34.100 208.490 ;
        RECT 32.920 207.830 33.180 208.150 ;
        RECT 33.830 207.975 34.110 208.345 ;
        RECT 35.220 208.170 35.480 208.490 ;
        RECT 35.680 207.830 35.940 208.150 ;
        RECT 32.980 206.700 33.120 207.830 ;
        RECT 33.650 206.955 35.190 207.325 ;
        RECT 32.980 206.560 34.960 206.700 ;
        RECT 34.300 205.790 34.560 206.110 ;
        RECT 33.840 205.450 34.100 205.770 ;
        RECT 32.920 204.770 33.180 205.090 ;
        RECT 32.980 200.865 33.120 204.770 ;
        RECT 33.380 203.070 33.640 203.390 ;
        RECT 33.440 202.710 33.580 203.070 ;
        RECT 33.900 202.905 34.040 205.450 ;
        RECT 34.360 203.730 34.500 205.790 ;
        RECT 34.820 203.730 34.960 206.560 ;
        RECT 35.220 206.470 35.480 206.790 ;
        RECT 35.280 205.090 35.420 206.470 ;
        RECT 35.220 204.770 35.480 205.090 ;
        RECT 34.300 203.410 34.560 203.730 ;
        RECT 34.760 203.410 35.020 203.730 ;
        RECT 33.380 202.390 33.640 202.710 ;
        RECT 33.830 202.535 34.110 202.905 ;
        RECT 33.650 201.515 35.190 201.885 ;
        RECT 32.910 200.495 33.190 200.865 ;
        RECT 33.380 200.690 33.640 201.010 ;
        RECT 32.460 200.010 32.720 200.330 ;
        RECT 32.460 199.560 32.720 199.650 ;
        RECT 33.440 199.560 33.580 200.690 ;
        RECT 33.830 200.495 34.110 200.865 ;
        RECT 33.900 200.330 34.040 200.495 ;
        RECT 33.840 200.010 34.100 200.330 ;
        RECT 34.300 200.010 34.560 200.330 ;
        RECT 35.740 200.185 35.880 207.830 ;
        RECT 37.120 206.870 37.260 208.850 ;
        RECT 37.580 208.345 37.720 209.280 ;
        RECT 39.880 208.830 40.020 210.695 ;
        RECT 37.980 208.510 38.240 208.830 ;
        RECT 38.440 208.510 38.700 208.830 ;
        RECT 39.820 208.510 40.080 208.830 ;
        RECT 37.510 207.975 37.790 208.345 ;
        RECT 38.040 207.665 38.180 208.510 ;
        RECT 38.500 208.345 38.640 208.510 ;
        RECT 38.430 207.975 38.710 208.345 ;
        RECT 38.900 208.170 39.160 208.490 ;
        RECT 37.970 207.295 38.250 207.665 ;
        RECT 37.120 206.730 38.180 206.870 ;
        RECT 36.200 205.880 37.260 206.020 ;
        RECT 37.510 205.935 37.790 206.305 ;
        RECT 36.200 204.265 36.340 205.880 ;
        RECT 36.600 205.110 36.860 205.430 ;
        RECT 36.130 203.895 36.410 204.265 ;
        RECT 36.140 202.730 36.400 203.050 ;
        RECT 36.200 201.545 36.340 202.730 ;
        RECT 36.660 202.225 36.800 205.110 ;
        RECT 37.120 205.000 37.260 205.880 ;
        RECT 37.580 205.770 37.720 205.935 ;
        RECT 38.040 205.770 38.180 206.730 ;
        RECT 38.960 206.110 39.100 208.170 ;
        RECT 39.360 207.490 39.620 207.810 ;
        RECT 38.900 205.790 39.160 206.110 ;
        RECT 37.520 205.450 37.780 205.770 ;
        RECT 37.980 205.450 38.240 205.770 ;
        RECT 37.120 204.860 39.100 205.000 ;
        RECT 39.420 204.945 39.560 207.490 ;
        RECT 39.880 205.770 40.020 208.510 ;
        RECT 39.820 205.450 40.080 205.770 ;
        RECT 36.950 204.235 38.490 204.605 ;
        RECT 38.960 204.265 39.100 204.860 ;
        RECT 39.350 204.575 39.630 204.945 ;
        RECT 38.890 203.895 39.170 204.265 ;
        RECT 37.060 203.070 37.320 203.390 ;
        RECT 37.120 202.370 37.260 203.070 ;
        RECT 37.520 202.730 37.780 203.050 ;
        RECT 36.590 201.855 36.870 202.225 ;
        RECT 37.060 202.050 37.320 202.370 ;
        RECT 36.130 201.175 36.410 201.545 ;
        RECT 37.580 201.350 37.720 202.730 ;
        RECT 38.900 202.390 39.160 202.710 ;
        RECT 39.360 202.390 39.620 202.710 ;
        RECT 37.520 201.030 37.780 201.350 ;
        RECT 37.980 201.030 38.240 201.350 ;
        RECT 38.430 201.175 38.710 201.545 ;
        RECT 38.040 200.580 38.180 201.030 ;
        RECT 36.200 200.440 38.180 200.580 ;
        RECT 32.460 199.420 33.580 199.560 ;
        RECT 32.460 199.330 32.720 199.420 ;
        RECT 33.840 199.330 34.100 199.650 ;
        RECT 33.900 198.710 34.040 199.330 ;
        RECT 34.360 198.825 34.500 200.010 ;
        RECT 35.670 199.815 35.950 200.185 ;
        RECT 36.200 199.505 36.340 200.440 ;
        RECT 38.500 199.990 38.640 201.175 ;
        RECT 38.960 199.990 39.100 202.390 ;
        RECT 38.440 199.670 38.700 199.990 ;
        RECT 38.900 199.670 39.160 199.990 ;
        RECT 36.130 199.135 36.410 199.505 ;
        RECT 32.000 198.310 32.260 198.630 ;
        RECT 33.440 198.570 34.040 198.710 ;
        RECT 33.440 198.540 33.580 198.570 ;
        RECT 32.980 198.400 33.580 198.540 ;
        RECT 34.290 198.455 34.570 198.825 ;
        RECT 36.950 198.795 38.490 199.165 ;
        RECT 31.540 198.145 31.800 198.290 ;
        RECT 31.530 197.775 31.810 198.145 ;
        RECT 31.540 197.290 31.800 197.610 ;
        RECT 31.600 195.570 31.740 197.290 ;
        RECT 32.980 197.180 33.120 198.400 ;
        RECT 35.680 198.310 35.940 198.630 ;
        RECT 38.890 198.455 39.170 198.825 ;
        RECT 39.420 198.630 39.560 202.390 ;
        RECT 39.820 201.030 40.080 201.350 ;
        RECT 39.880 199.505 40.020 201.030 ;
        RECT 39.810 199.135 40.090 199.505 ;
        RECT 33.370 197.775 33.650 198.145 ;
        RECT 33.380 197.630 33.640 197.775 ;
        RECT 34.300 197.630 34.560 197.950 ;
        RECT 32.425 197.040 33.120 197.180 ;
        RECT 32.000 196.610 32.260 196.930 ;
        RECT 31.540 195.250 31.800 195.570 ;
        RECT 31.530 194.375 31.810 194.745 ;
        RECT 31.600 192.510 31.740 194.375 ;
        RECT 32.060 192.510 32.200 196.610 ;
        RECT 32.425 195.990 32.565 197.040 ;
        RECT 34.360 196.840 34.500 197.630 ;
        RECT 35.740 196.840 35.880 198.310 ;
        RECT 38.440 198.200 38.700 198.290 ;
        RECT 38.040 198.060 38.700 198.200 ;
        RECT 37.060 197.630 37.320 197.950 ;
        RECT 34.360 196.700 35.880 196.840 ;
        RECT 33.650 196.075 35.190 196.445 ;
        RECT 32.425 195.850 32.660 195.990 ;
        RECT 31.540 192.190 31.800 192.510 ;
        RECT 32.000 192.190 32.260 192.510 ;
        RECT 31.530 191.655 31.810 192.025 ;
        RECT 32.000 191.740 32.260 191.830 ;
        RECT 32.520 191.740 32.660 195.850 ;
        RECT 33.380 195.480 33.640 195.570 ;
        RECT 33.380 195.340 34.500 195.480 ;
        RECT 33.380 195.250 33.640 195.340 ;
        RECT 33.380 194.570 33.640 194.890 ;
        RECT 33.440 194.210 33.580 194.570 ;
        RECT 33.380 193.890 33.640 194.210 ;
        RECT 33.840 193.890 34.100 194.210 ;
        RECT 33.440 192.705 33.580 193.890 ;
        RECT 33.900 193.385 34.040 193.890 ;
        RECT 33.830 193.015 34.110 193.385 ;
        RECT 33.840 192.760 34.100 192.850 ;
        RECT 34.360 192.760 34.500 195.340 ;
        RECT 35.220 194.800 35.480 194.890 ;
        RECT 35.740 194.800 35.880 196.700 ;
        RECT 36.130 195.735 36.410 196.105 ;
        RECT 36.200 195.570 36.340 195.735 ;
        RECT 36.140 195.250 36.400 195.570 ;
        RECT 36.600 194.800 36.860 194.890 ;
        RECT 35.220 194.660 35.880 194.800 ;
        RECT 36.200 194.660 36.860 194.800 ;
        RECT 35.220 194.570 35.480 194.660 ;
        RECT 33.370 192.335 33.650 192.705 ;
        RECT 33.840 192.620 34.500 192.760 ;
        RECT 33.840 192.530 34.100 192.620 ;
        RECT 35.280 192.025 35.420 194.570 ;
        RECT 36.200 192.510 36.340 194.660 ;
        RECT 36.600 194.570 36.860 194.660 ;
        RECT 37.120 194.120 37.260 197.630 ;
        RECT 38.040 194.210 38.180 198.060 ;
        RECT 38.440 197.970 38.700 198.060 ;
        RECT 38.960 197.950 39.100 198.455 ;
        RECT 39.360 198.310 39.620 198.630 ;
        RECT 38.900 197.630 39.160 197.950 ;
        RECT 38.440 196.610 38.700 196.930 ;
        RECT 36.660 193.980 37.260 194.120 ;
        RECT 35.680 192.190 35.940 192.510 ;
        RECT 36.140 192.190 36.400 192.510 ;
        RECT 31.600 189.790 31.740 191.655 ;
        RECT 32.000 191.600 32.660 191.740 ;
        RECT 35.210 191.655 35.490 192.025 ;
        RECT 32.000 191.510 32.260 191.600 ;
        RECT 31.540 189.470 31.800 189.790 ;
        RECT 32.060 187.945 32.200 191.510 ;
        RECT 32.910 190.975 33.190 191.345 ;
        RECT 32.450 190.295 32.730 190.665 ;
        RECT 31.990 187.575 32.270 187.945 ;
        RECT 32.520 187.320 32.660 190.295 ;
        RECT 31.600 187.180 32.660 187.320 ;
        RECT 31.080 184.370 31.340 184.690 ;
        RECT 30.160 181.990 30.420 182.135 ;
        RECT 30.620 181.990 30.880 182.310 ;
        RECT 30.680 178.910 30.820 181.990 ;
        RECT 31.600 181.970 31.740 187.180 ;
        RECT 31.990 186.215 32.270 186.585 ;
        RECT 32.460 186.410 32.720 186.730 ;
        RECT 32.060 186.050 32.200 186.215 ;
        RECT 32.000 185.730 32.260 186.050 ;
        RECT 31.990 184.855 32.270 185.225 ;
        RECT 32.000 184.710 32.260 184.855 ;
        RECT 32.000 183.920 32.260 184.010 ;
        RECT 32.520 183.920 32.660 186.410 ;
        RECT 32.000 183.780 32.660 183.920 ;
        RECT 32.000 183.690 32.260 183.780 ;
        RECT 32.460 183.010 32.720 183.330 ;
        RECT 32.520 182.505 32.660 183.010 ;
        RECT 32.450 182.135 32.730 182.505 ;
        RECT 31.540 181.650 31.800 181.970 ;
        RECT 32.980 181.630 33.120 190.975 ;
        RECT 33.650 190.635 35.190 191.005 ;
        RECT 33.380 189.470 33.640 189.790 ;
        RECT 34.760 189.470 35.020 189.790 ;
        RECT 33.440 187.070 33.580 189.470 ;
        RECT 33.830 188.935 34.110 189.305 ;
        RECT 33.380 186.750 33.640 187.070 ;
        RECT 33.900 186.050 34.040 188.935 ;
        RECT 34.300 188.625 34.560 188.770 ;
        RECT 34.290 188.255 34.570 188.625 ;
        RECT 34.820 187.070 34.960 189.470 ;
        RECT 35.740 188.770 35.880 192.190 ;
        RECT 36.140 191.510 36.400 191.830 ;
        RECT 36.200 189.790 36.340 191.510 ;
        RECT 36.140 189.470 36.400 189.790 ;
        RECT 35.220 188.450 35.480 188.770 ;
        RECT 35.680 188.450 35.940 188.770 ;
        RECT 35.280 187.945 35.420 188.450 ;
        RECT 35.210 187.575 35.490 187.945 ;
        RECT 34.760 186.750 35.020 187.070 ;
        RECT 33.840 185.730 34.100 186.050 ;
        RECT 35.740 185.960 35.880 188.450 ;
        RECT 36.130 187.575 36.410 187.945 ;
        RECT 36.660 187.660 36.800 193.980 ;
        RECT 37.980 193.890 38.240 194.210 ;
        RECT 38.500 194.120 38.640 196.610 ;
        RECT 38.960 195.570 39.100 197.630 ;
        RECT 39.420 196.105 39.560 198.310 ;
        RECT 39.820 196.950 40.080 197.270 ;
        RECT 39.350 195.735 39.630 196.105 ;
        RECT 38.900 195.250 39.160 195.570 ;
        RECT 39.880 194.890 40.020 196.950 ;
        RECT 38.900 194.630 39.160 194.890 ;
        RECT 39.820 194.745 40.080 194.890 ;
        RECT 38.900 194.570 39.560 194.630 ;
        RECT 38.960 194.490 39.560 194.570 ;
        RECT 38.500 193.980 39.100 194.120 ;
        RECT 36.950 193.355 38.490 193.725 ;
        RECT 37.060 192.870 37.320 193.190 ;
        RECT 37.120 191.830 37.260 192.870 ;
        RECT 37.520 192.190 37.780 192.510 ;
        RECT 37.060 191.510 37.320 191.830 ;
        RECT 37.580 191.345 37.720 192.190 ;
        RECT 37.980 191.850 38.240 192.170 ;
        RECT 37.510 190.975 37.790 191.345 ;
        RECT 37.510 190.295 37.790 190.665 ;
        RECT 37.580 190.130 37.720 190.295 ;
        RECT 37.050 189.615 37.330 189.985 ;
        RECT 37.520 189.810 37.780 190.130 ;
        RECT 37.120 189.450 37.260 189.615 ;
        RECT 37.060 189.130 37.320 189.450 ;
        RECT 38.040 189.305 38.180 191.850 ;
        RECT 38.440 191.170 38.700 191.490 ;
        RECT 38.500 189.360 38.640 191.170 ;
        RECT 38.960 190.130 39.100 193.980 ;
        RECT 39.420 192.170 39.560 194.490 ;
        RECT 39.810 194.375 40.090 194.745 ;
        RECT 39.820 193.890 40.080 194.210 ;
        RECT 39.880 192.850 40.020 193.890 ;
        RECT 39.820 192.530 40.080 192.850 ;
        RECT 39.360 192.025 39.620 192.170 ;
        RECT 39.350 191.655 39.630 192.025 ;
        RECT 38.900 189.810 39.160 190.130 ;
        RECT 39.360 189.810 39.620 190.130 ;
        RECT 37.970 188.935 38.250 189.305 ;
        RECT 38.500 189.220 39.100 189.360 ;
        RECT 36.950 187.915 38.490 188.285 ;
        RECT 36.200 186.470 36.340 187.575 ;
        RECT 36.660 187.520 37.260 187.660 ;
        RECT 36.200 186.330 36.800 186.470 ;
        RECT 35.740 185.820 36.340 185.960 ;
        RECT 33.650 185.195 35.190 185.565 ;
        RECT 33.380 184.710 33.640 185.030 ;
        RECT 35.220 184.710 35.480 185.030 ;
        RECT 33.440 184.545 33.580 184.710 ;
        RECT 33.370 184.175 33.650 184.545 ;
        RECT 34.290 184.175 34.570 184.545 ;
        RECT 34.360 184.010 34.500 184.175 ;
        RECT 33.830 183.495 34.110 183.865 ;
        RECT 34.300 183.690 34.560 184.010 ;
        RECT 33.900 181.970 34.040 183.495 ;
        RECT 35.280 182.310 35.420 184.710 ;
        RECT 35.680 183.350 35.940 183.670 ;
        RECT 35.740 183.185 35.880 183.350 ;
        RECT 35.670 182.815 35.950 183.185 ;
        RECT 35.220 181.990 35.480 182.310 ;
        RECT 33.840 181.650 34.100 181.970 ;
        RECT 32.920 181.310 33.180 181.630 ;
        RECT 31.990 180.860 32.270 181.145 ;
        RECT 32.460 180.860 32.720 180.950 ;
        RECT 31.990 180.775 32.720 180.860 ;
        RECT 32.910 180.775 33.190 181.145 ;
        RECT 32.060 180.720 32.720 180.775 ;
        RECT 30.620 178.590 30.880 178.910 ;
        RECT 31.540 172.810 31.800 173.130 ;
        RECT 30.620 172.130 30.880 172.450 ;
        RECT 29.760 171.370 30.360 171.510 ;
        RECT 30.680 171.430 30.820 172.130 ;
        RECT 31.600 171.430 31.740 172.810 ;
        RECT 28.780 170.430 29.040 170.750 ;
        RECT 29.240 170.660 29.500 170.750 ;
        RECT 29.240 170.520 29.900 170.660 ;
        RECT 29.240 170.430 29.500 170.520 ;
        RECT 29.760 167.690 29.900 170.520 ;
        RECT 29.240 167.370 29.500 167.690 ;
        RECT 29.700 167.370 29.960 167.690 ;
        RECT 28.380 165.930 28.980 166.070 ;
        RECT 29.300 165.990 29.440 167.370 ;
        RECT 27.860 164.990 28.120 165.310 ;
        RECT 28.320 164.990 28.580 165.310 ;
        RECT 27.920 163.270 28.060 164.990 ;
        RECT 27.860 162.950 28.120 163.270 ;
        RECT 28.380 161.570 28.520 164.990 ;
        RECT 28.320 161.250 28.580 161.570 ;
        RECT 26.480 157.510 26.740 157.830 ;
        RECT 26.540 156.470 26.680 157.510 ;
        RECT 27.400 157.170 27.660 157.490 ;
        RECT 27.460 156.810 27.600 157.170 ;
        RECT 27.400 156.490 27.660 156.810 ;
        RECT 26.480 156.150 26.740 156.470 ;
        RECT 25.560 154.790 25.820 155.110 ;
        RECT 25.620 152.390 25.760 154.790 ;
        RECT 26.540 153.750 26.680 156.150 ;
        RECT 27.460 154.090 27.600 156.490 ;
        RECT 26.940 153.770 27.200 154.090 ;
        RECT 27.400 153.770 27.660 154.090 ;
        RECT 26.480 153.430 26.740 153.750 ;
        RECT 25.100 152.070 25.360 152.390 ;
        RECT 25.560 152.070 25.820 152.390 ;
        RECT 21.420 150.710 21.680 151.030 ;
        RECT 21.480 148.990 21.620 150.710 ;
        RECT 21.420 148.670 21.680 148.990 ;
        RECT 25.160 148.650 25.300 152.070 ;
        RECT 25.620 151.370 25.760 152.070 ;
        RECT 26.540 152.050 26.680 153.430 ;
        RECT 27.000 152.050 27.140 153.770 ;
        RECT 26.480 151.730 26.740 152.050 ;
        RECT 26.940 151.730 27.200 152.050 ;
        RECT 25.560 151.050 25.820 151.370 ;
        RECT 27.460 151.030 27.600 153.770 ;
        RECT 27.400 150.710 27.660 151.030 ;
        RECT 20.030 148.135 20.310 148.505 ;
        RECT 25.100 148.330 25.360 148.650 ;
        RECT 20.040 147.990 20.300 148.135 ;
        RECT 28.840 143.550 28.980 165.930 ;
        RECT 29.240 165.670 29.500 165.990 ;
        RECT 30.220 164.290 30.360 171.370 ;
        RECT 30.620 171.110 30.880 171.430 ;
        RECT 31.540 171.110 31.800 171.430 ;
        RECT 31.540 170.430 31.800 170.750 ;
        RECT 31.600 168.370 31.740 170.430 ;
        RECT 31.080 168.225 31.340 168.370 ;
        RECT 31.070 167.855 31.350 168.225 ;
        RECT 31.540 168.050 31.800 168.370 ;
        RECT 31.600 167.690 31.740 168.050 ;
        RECT 31.540 167.370 31.800 167.690 ;
        RECT 30.160 163.970 30.420 164.290 ;
        RECT 32.060 162.500 32.200 180.720 ;
        RECT 32.460 180.630 32.720 180.720 ;
        RECT 32.980 179.590 33.120 180.775 ;
        RECT 33.650 179.755 35.190 180.125 ;
        RECT 32.920 179.270 33.180 179.590 ;
        RECT 33.380 178.250 33.640 178.570 ;
        RECT 33.840 178.250 34.100 178.570 ;
        RECT 34.300 178.250 34.560 178.570 ;
        RECT 33.440 176.870 33.580 178.250 ;
        RECT 33.380 176.550 33.640 176.870 ;
        RECT 33.900 175.850 34.040 178.250 ;
        RECT 34.360 176.190 34.500 178.250 ;
        RECT 35.220 177.910 35.480 178.230 ;
        RECT 34.300 175.870 34.560 176.190 ;
        RECT 33.840 175.530 34.100 175.850 ;
        RECT 35.280 175.760 35.420 177.910 ;
        RECT 35.740 176.530 35.880 182.815 ;
        RECT 36.200 182.310 36.340 185.820 ;
        RECT 36.660 183.330 36.800 186.330 ;
        RECT 37.120 183.330 37.260 187.520 ;
        RECT 37.980 187.430 38.240 187.750 ;
        RECT 37.520 186.750 37.780 187.070 ;
        RECT 37.580 185.030 37.720 186.750 ;
        RECT 38.040 185.030 38.180 187.430 ;
        RECT 37.520 184.710 37.780 185.030 ;
        RECT 37.980 184.710 38.240 185.030 ;
        RECT 37.970 184.175 38.250 184.545 ;
        RECT 38.040 184.010 38.180 184.175 ;
        RECT 37.980 183.690 38.240 184.010 ;
        RECT 36.600 183.010 36.860 183.330 ;
        RECT 37.060 183.010 37.320 183.330 ;
        RECT 36.140 181.990 36.400 182.310 ;
        RECT 36.140 180.970 36.400 181.290 ;
        RECT 35.680 176.210 35.940 176.530 ;
        RECT 36.200 175.850 36.340 180.970 ;
        RECT 36.660 179.250 36.800 183.010 ;
        RECT 36.950 182.475 38.490 182.845 ;
        RECT 37.060 181.990 37.320 182.310 ;
        RECT 38.960 182.220 39.100 189.220 ;
        RECT 39.420 186.390 39.560 189.810 ;
        RECT 39.880 189.450 40.020 192.530 ;
        RECT 39.820 189.130 40.080 189.450 ;
        RECT 39.810 186.895 40.090 187.265 ;
        RECT 39.360 186.070 39.620 186.390 ;
        RECT 39.420 184.350 39.560 186.070 ;
        RECT 39.360 184.030 39.620 184.350 ;
        RECT 39.880 183.750 40.020 186.895 ;
        RECT 40.340 185.030 40.480 217.610 ;
        RECT 41.650 217.330 41.930 221.330 ;
        RECT 44.870 217.330 45.150 221.330 ;
        RECT 48.090 217.330 48.370 221.330 ;
        RECT 51.310 217.330 51.590 221.330 ;
        RECT 54.530 217.330 54.810 221.330 ;
        RECT 57.750 217.330 58.030 221.330 ;
        RECT 60.970 217.330 61.250 221.330 ;
        RECT 64.190 217.330 64.470 221.330 ;
        RECT 67.410 217.330 67.690 221.330 ;
        RECT 70.630 217.330 70.910 221.330 ;
        RECT 71.160 217.610 72.680 217.750 ;
        RECT 41.720 214.270 41.860 217.330 ;
        RECT 41.660 213.950 41.920 214.270 ;
        RECT 42.120 211.230 42.380 211.550 ;
        RECT 41.660 210.210 41.920 210.530 ;
        RECT 41.720 208.830 41.860 210.210 ;
        RECT 41.660 208.510 41.920 208.830 ;
        RECT 41.200 208.170 41.460 208.490 ;
        RECT 40.740 207.490 41.000 207.810 ;
        RECT 40.800 198.630 40.940 207.490 ;
        RECT 41.260 202.370 41.400 208.170 ;
        RECT 41.660 205.110 41.920 205.430 ;
        RECT 41.200 202.050 41.460 202.370 ;
        RECT 41.720 201.430 41.860 205.110 ;
        RECT 41.260 201.290 41.860 201.430 ;
        RECT 41.260 198.630 41.400 201.290 ;
        RECT 41.660 199.330 41.920 199.650 ;
        RECT 40.740 198.310 41.000 198.630 ;
        RECT 41.200 198.310 41.460 198.630 ;
        RECT 41.720 197.950 41.860 199.330 ;
        RECT 41.200 197.630 41.460 197.950 ;
        RECT 41.660 197.630 41.920 197.950 ;
        RECT 40.740 197.290 41.000 197.610 ;
        RECT 40.800 196.105 40.940 197.290 ;
        RECT 40.730 195.735 41.010 196.105 ;
        RECT 40.740 194.230 41.000 194.550 ;
        RECT 40.280 184.710 40.540 185.030 ;
        RECT 38.040 182.080 39.100 182.220 ;
        RECT 39.420 183.610 40.020 183.750 ;
        RECT 36.600 178.930 36.860 179.250 ;
        RECT 37.120 178.480 37.260 181.990 ;
        RECT 37.510 179.415 37.790 179.785 ;
        RECT 37.580 178.570 37.720 179.415 ;
        RECT 38.040 178.570 38.180 182.080 ;
        RECT 38.890 179.415 39.170 179.785 ;
        RECT 38.960 178.570 39.100 179.415 ;
        RECT 36.660 178.340 37.260 178.480 ;
        RECT 35.280 175.620 35.880 175.760 ;
        RECT 33.650 174.315 35.190 174.685 ;
        RECT 34.300 173.490 34.560 173.810 ;
        RECT 32.450 170.750 32.730 170.945 ;
        RECT 34.360 170.750 34.500 173.490 ;
        RECT 32.365 170.575 32.730 170.750 ;
        RECT 32.365 170.520 32.660 170.575 ;
        RECT 32.365 170.430 32.625 170.520 ;
        RECT 34.300 170.430 34.560 170.750 ;
        RECT 34.360 169.730 34.500 170.430 ;
        RECT 34.300 169.410 34.560 169.730 ;
        RECT 33.650 168.875 35.190 169.245 ;
        RECT 35.740 168.710 35.880 175.620 ;
        RECT 36.140 175.530 36.400 175.850 ;
        RECT 36.200 173.130 36.340 175.530 ;
        RECT 36.140 172.810 36.400 173.130 ;
        RECT 33.380 168.390 33.640 168.710 ;
        RECT 35.680 168.390 35.940 168.710 ;
        RECT 33.440 167.690 33.580 168.390 ;
        RECT 33.380 167.370 33.640 167.690 ;
        RECT 35.680 167.370 35.940 167.690 ;
        RECT 32.920 167.030 33.180 167.350 ;
        RECT 32.450 165.135 32.730 165.505 ;
        RECT 31.140 162.360 32.200 162.500 ;
        RECT 30.620 161.930 30.880 162.250 ;
        RECT 30.680 160.210 30.820 161.930 ;
        RECT 30.620 159.890 30.880 160.210 ;
        RECT 29.240 157.510 29.500 157.830 ;
        RECT 29.300 154.770 29.440 157.510 ;
        RECT 31.140 156.130 31.280 162.360 ;
        RECT 32.000 161.590 32.260 161.910 ;
        RECT 32.060 159.870 32.200 161.590 ;
        RECT 31.540 159.550 31.800 159.870 ;
        RECT 32.000 159.550 32.260 159.870 ;
        RECT 31.080 155.810 31.340 156.130 ;
        RECT 29.240 154.450 29.500 154.770 ;
        RECT 29.700 154.450 29.960 154.770 ;
        RECT 29.240 153.430 29.500 153.750 ;
        RECT 29.300 151.030 29.440 153.430 ;
        RECT 29.240 150.710 29.500 151.030 ;
        RECT 29.760 150.690 29.900 154.450 ;
        RECT 31.600 154.090 31.740 159.550 ;
        RECT 32.060 157.830 32.200 159.550 ;
        RECT 32.000 157.510 32.260 157.830 ;
        RECT 31.540 153.770 31.800 154.090 ;
        RECT 32.000 153.770 32.260 154.090 ;
        RECT 32.060 151.030 32.200 153.770 ;
        RECT 32.520 152.390 32.660 165.135 ;
        RECT 32.980 164.970 33.120 167.030 ;
        RECT 33.440 165.990 33.580 167.370 ;
        RECT 33.380 165.670 33.640 165.990 ;
        RECT 32.920 164.650 33.180 164.970 ;
        RECT 33.650 163.435 35.190 163.805 ;
        RECT 35.740 163.270 35.880 167.370 ;
        RECT 35.680 162.950 35.940 163.270 ;
        RECT 34.760 161.930 35.020 162.250 ;
        RECT 35.680 162.160 35.940 162.250 ;
        RECT 36.200 162.160 36.340 172.810 ;
        RECT 35.680 162.020 36.340 162.160 ;
        RECT 35.680 161.930 35.940 162.020 ;
        RECT 34.820 160.550 34.960 161.930 ;
        RECT 34.760 160.230 35.020 160.550 ;
        RECT 33.650 157.995 35.190 158.365 ;
        RECT 33.650 152.555 35.190 152.925 ;
        RECT 32.460 152.070 32.720 152.390 ;
        RECT 35.740 152.300 35.880 161.930 ;
        RECT 36.140 161.250 36.400 161.570 ;
        RECT 36.200 159.870 36.340 161.250 ;
        RECT 36.140 159.550 36.400 159.870 ;
        RECT 36.660 157.490 36.800 178.340 ;
        RECT 37.520 178.250 37.780 178.570 ;
        RECT 37.980 178.250 38.240 178.570 ;
        RECT 38.900 178.250 39.160 178.570 ;
        RECT 38.900 177.570 39.160 177.890 ;
        RECT 36.950 177.035 38.490 177.405 ;
        RECT 38.960 177.065 39.100 177.570 ;
        RECT 38.890 176.695 39.170 177.065 ;
        RECT 38.960 175.170 39.100 176.695 ;
        RECT 38.900 174.850 39.160 175.170 ;
        RECT 39.420 173.810 39.560 183.610 ;
        RECT 39.820 183.010 40.080 183.330 ;
        RECT 39.880 177.890 40.020 183.010 ;
        RECT 40.800 181.630 40.940 194.230 ;
        RECT 41.260 194.210 41.400 197.630 ;
        RECT 41.650 197.095 41.930 197.465 ;
        RECT 41.720 195.230 41.860 197.095 ;
        RECT 41.660 194.910 41.920 195.230 ;
        RECT 41.200 193.890 41.460 194.210 ;
        RECT 42.180 192.420 42.320 211.230 ;
        RECT 42.580 208.510 42.840 208.830 ;
        RECT 42.640 206.450 42.780 208.510 ;
        RECT 43.950 207.975 44.230 208.345 ;
        RECT 43.030 207.295 43.310 207.665 ;
        RECT 42.580 206.130 42.840 206.450 ;
        RECT 42.580 202.905 42.840 203.050 ;
        RECT 42.570 202.535 42.850 202.905 ;
        RECT 42.570 201.430 42.850 201.545 ;
        RECT 43.100 201.430 43.240 207.295 ;
        RECT 43.500 205.450 43.760 205.770 ;
        RECT 42.570 201.290 43.240 201.430 ;
        RECT 42.570 201.175 42.850 201.290 ;
        RECT 42.640 197.610 42.780 201.175 ;
        RECT 42.580 197.290 42.840 197.610 ;
        RECT 43.040 197.465 43.300 197.610 ;
        RECT 43.030 197.095 43.310 197.465 ;
        RECT 42.580 196.610 42.840 196.930 ;
        RECT 43.560 196.840 43.700 205.450 ;
        RECT 44.020 197.950 44.160 207.975 ;
        RECT 44.420 204.770 44.680 205.090 ;
        RECT 44.480 197.950 44.620 204.770 ;
        RECT 43.960 197.630 44.220 197.950 ;
        RECT 44.420 197.630 44.680 197.950 ;
        RECT 43.100 196.700 43.700 196.840 ;
        RECT 41.260 192.280 42.320 192.420 ;
        RECT 41.260 185.225 41.400 192.280 ;
        RECT 41.660 191.740 41.920 191.830 ;
        RECT 41.660 191.600 42.320 191.740 ;
        RECT 41.660 191.510 41.920 191.600 ;
        RECT 41.660 190.150 41.920 190.470 ;
        RECT 41.720 186.050 41.860 190.150 ;
        RECT 42.180 187.660 42.320 191.600 ;
        RECT 42.640 190.470 42.780 196.610 ;
        RECT 43.100 194.065 43.240 196.700 ;
        RECT 43.500 194.570 43.760 194.890 ;
        RECT 44.020 194.745 44.160 197.630 ;
        RECT 44.410 197.095 44.690 197.465 ;
        RECT 44.480 195.910 44.620 197.095 ;
        RECT 44.420 195.590 44.680 195.910 ;
        RECT 44.420 194.910 44.680 195.230 ;
        RECT 43.030 193.695 43.310 194.065 ;
        RECT 43.040 192.190 43.300 192.510 ;
        RECT 42.580 190.150 42.840 190.470 ;
        RECT 43.100 187.945 43.240 192.190 ;
        RECT 43.560 190.470 43.700 194.570 ;
        RECT 43.950 194.375 44.230 194.745 ;
        RECT 44.480 194.210 44.620 194.910 ;
        RECT 43.960 193.890 44.220 194.210 ;
        RECT 44.420 193.890 44.680 194.210 ;
        RECT 44.020 191.490 44.160 193.890 ;
        RECT 44.420 191.850 44.680 192.170 ;
        RECT 43.960 191.170 44.220 191.490 ;
        RECT 43.500 190.150 43.760 190.470 ;
        RECT 43.500 189.130 43.760 189.450 ;
        RECT 42.180 187.520 42.780 187.660 ;
        RECT 43.030 187.575 43.310 187.945 ;
        RECT 43.560 187.750 43.700 189.130 ;
        RECT 43.950 188.255 44.230 188.625 ;
        RECT 44.020 187.750 44.160 188.255 ;
        RECT 42.120 186.750 42.380 187.070 ;
        RECT 42.180 186.585 42.320 186.750 ;
        RECT 42.110 186.215 42.390 186.585 ;
        RECT 41.660 185.730 41.920 186.050 ;
        RECT 41.190 184.855 41.470 185.225 ;
        RECT 41.200 183.690 41.460 184.010 ;
        RECT 41.660 183.690 41.920 184.010 ;
        RECT 41.260 182.310 41.400 183.690 ;
        RECT 41.200 181.990 41.460 182.310 ;
        RECT 40.740 181.310 41.000 181.630 ;
        RECT 40.800 178.990 40.940 181.310 ;
        RECT 41.190 179.415 41.470 179.785 ;
        RECT 40.340 178.850 40.940 178.990 ;
        RECT 40.340 178.570 40.480 178.850 ;
        RECT 40.280 178.250 40.540 178.570 ;
        RECT 40.740 178.250 41.000 178.570 ;
        RECT 39.820 177.800 40.080 177.890 ;
        RECT 39.820 177.660 40.480 177.800 ;
        RECT 39.820 177.570 40.080 177.660 ;
        RECT 40.340 176.870 40.480 177.660 ;
        RECT 40.280 176.550 40.540 176.870 ;
        RECT 39.820 175.870 40.080 176.190 ;
        RECT 39.360 173.490 39.620 173.810 ;
        RECT 38.900 172.130 39.160 172.450 ;
        RECT 36.950 171.595 38.490 171.965 ;
        RECT 38.960 171.430 39.100 172.130 ;
        RECT 38.900 171.110 39.160 171.430 ;
        RECT 37.060 170.430 37.320 170.750 ;
        RECT 37.120 168.710 37.260 170.430 ;
        RECT 37.520 169.410 37.780 169.730 ;
        RECT 37.060 168.390 37.320 168.710 ;
        RECT 37.580 167.545 37.720 169.410 ;
        RECT 37.980 168.390 38.240 168.710 ;
        RECT 37.510 167.175 37.790 167.545 ;
        RECT 38.040 167.010 38.180 168.390 ;
        RECT 38.960 168.030 39.100 171.110 ;
        RECT 39.350 170.575 39.630 170.945 ;
        RECT 39.420 170.410 39.560 170.575 ;
        RECT 39.360 170.090 39.620 170.410 ;
        RECT 38.900 167.710 39.160 168.030 ;
        RECT 38.890 167.175 39.170 167.545 ;
        RECT 37.980 166.690 38.240 167.010 ;
        RECT 36.950 166.155 38.490 166.525 ;
        RECT 38.960 165.650 39.100 167.175 ;
        RECT 38.900 165.330 39.160 165.650 ;
        RECT 38.960 163.180 39.100 165.330 ;
        RECT 38.500 163.040 39.100 163.180 ;
        RECT 38.500 161.910 38.640 163.040 ;
        RECT 38.900 162.500 39.160 162.590 ;
        RECT 39.420 162.500 39.560 170.090 ;
        RECT 39.880 169.730 40.020 175.870 ;
        RECT 40.340 170.410 40.480 176.550 ;
        RECT 40.800 176.385 40.940 178.250 ;
        RECT 40.730 176.015 41.010 176.385 ;
        RECT 40.740 174.850 41.000 175.170 ;
        RECT 40.280 170.090 40.540 170.410 ;
        RECT 39.820 169.410 40.080 169.730 ;
        RECT 39.820 167.710 40.080 168.030 ;
        RECT 39.880 165.990 40.020 167.710 ;
        RECT 39.820 165.670 40.080 165.990 ;
        RECT 38.900 162.360 39.560 162.500 ;
        RECT 38.900 162.270 39.160 162.360 ;
        RECT 38.440 161.590 38.700 161.910 ;
        RECT 38.900 161.250 39.160 161.570 ;
        RECT 36.950 160.715 38.490 161.085 ;
        RECT 38.960 160.550 39.100 161.250 ;
        RECT 38.900 160.230 39.160 160.550 ;
        RECT 38.440 159.550 38.700 159.870 ;
        RECT 38.500 157.490 38.640 159.550 ;
        RECT 38.900 159.210 39.160 159.530 ;
        RECT 36.600 157.170 36.860 157.490 ;
        RECT 38.440 157.170 38.700 157.490 ;
        RECT 36.600 156.490 36.860 156.810 ;
        RECT 36.140 154.110 36.400 154.430 ;
        RECT 34.820 152.160 35.880 152.300 ;
        RECT 32.000 150.710 32.260 151.030 ;
        RECT 29.700 150.370 29.960 150.690 ;
        RECT 34.820 148.560 34.960 152.160 ;
        RECT 36.200 152.050 36.340 154.110 ;
        RECT 36.140 151.730 36.400 152.050 ;
        RECT 35.680 151.050 35.940 151.370 ;
        RECT 36.140 151.050 36.400 151.370 ;
        RECT 35.220 150.370 35.480 150.690 ;
        RECT 35.280 149.330 35.420 150.370 ;
        RECT 35.740 149.330 35.880 151.050 ;
        RECT 36.200 149.670 36.340 151.050 ;
        RECT 36.140 149.350 36.400 149.670 ;
        RECT 35.220 149.010 35.480 149.330 ;
        RECT 35.680 149.010 35.940 149.330 ;
        RECT 34.820 148.420 36.340 148.560 ;
        RECT 35.680 147.650 35.940 147.970 ;
        RECT 33.650 147.115 35.190 147.485 ;
        RECT 35.740 146.950 35.880 147.650 ;
        RECT 35.680 146.630 35.940 146.950 ;
        RECT 36.200 146.350 36.340 148.420 ;
        RECT 35.740 146.210 36.340 146.350 ;
        RECT 33.840 145.610 34.100 145.930 ;
        RECT 33.900 143.890 34.040 145.610 ;
        RECT 33.840 143.570 34.100 143.890 ;
        RECT 28.780 143.230 29.040 143.550 ;
        RECT 35.740 143.210 35.880 146.210 ;
        RECT 36.140 145.270 36.400 145.590 ;
        RECT 36.200 144.230 36.340 145.270 ;
        RECT 36.140 143.910 36.400 144.230 ;
        RECT 35.680 142.890 35.940 143.210 ;
        RECT 33.650 141.675 35.190 142.045 ;
        RECT 36.660 141.510 36.800 156.490 ;
        RECT 36.950 155.275 38.490 155.645 ;
        RECT 37.060 154.110 37.320 154.430 ;
        RECT 37.120 152.390 37.260 154.110 ;
        RECT 37.060 152.070 37.320 152.390 ;
        RECT 37.120 150.690 37.260 152.070 ;
        RECT 37.060 150.370 37.320 150.690 ;
        RECT 36.950 149.835 38.490 150.205 ;
        RECT 38.960 146.270 39.100 159.210 ;
        RECT 39.420 146.950 39.560 162.360 ;
        RECT 39.880 160.630 40.020 165.670 ;
        RECT 40.340 162.250 40.480 170.090 ;
        RECT 40.800 168.370 40.940 174.850 ;
        RECT 41.260 172.360 41.400 179.415 ;
        RECT 41.720 174.150 41.860 183.690 ;
        RECT 42.640 181.145 42.780 187.520 ;
        RECT 43.100 184.010 43.240 187.575 ;
        RECT 43.500 187.430 43.760 187.750 ;
        RECT 43.960 187.430 44.220 187.750 ;
        RECT 43.500 186.410 43.760 186.730 ;
        RECT 43.560 185.030 43.700 186.410 ;
        RECT 43.960 186.070 44.220 186.390 ;
        RECT 43.500 184.710 43.760 185.030 ;
        RECT 43.040 183.690 43.300 184.010 ;
        RECT 44.020 183.920 44.160 186.070 ;
        RECT 44.480 184.690 44.620 191.850 ;
        RECT 44.940 190.130 45.080 217.330 ;
        RECT 46.250 206.615 46.530 206.985 ;
        RECT 45.340 200.350 45.600 200.670 ;
        RECT 45.400 197.950 45.540 200.350 ;
        RECT 45.800 199.330 46.060 199.650 ;
        RECT 45.340 197.630 45.600 197.950 ;
        RECT 45.340 194.570 45.600 194.890 ;
        RECT 45.400 193.190 45.540 194.570 ;
        RECT 45.340 192.870 45.600 193.190 ;
        RECT 45.340 192.190 45.600 192.510 ;
        RECT 44.880 189.810 45.140 190.130 ;
        RECT 45.400 187.660 45.540 192.190 ;
        RECT 44.940 187.520 45.540 187.660 ;
        RECT 44.420 184.370 44.680 184.690 ;
        RECT 43.490 183.495 43.770 183.865 ;
        RECT 44.020 183.780 44.620 183.920 ;
        RECT 42.570 180.775 42.850 181.145 ;
        RECT 42.110 178.735 42.390 179.105 ;
        RECT 42.180 178.570 42.320 178.735 ;
        RECT 42.120 178.250 42.380 178.570 ;
        RECT 43.040 178.425 43.300 178.570 ;
        RECT 41.660 173.830 41.920 174.150 ;
        RECT 42.180 173.130 42.320 178.250 ;
        RECT 42.580 177.910 42.840 178.230 ;
        RECT 43.030 178.055 43.310 178.425 ;
        RECT 42.640 176.530 42.780 177.910 ;
        RECT 42.580 176.210 42.840 176.530 ;
        RECT 42.120 172.810 42.380 173.130 ;
        RECT 41.260 172.220 42.320 172.360 ;
        RECT 41.200 170.430 41.460 170.750 ;
        RECT 40.740 168.050 41.000 168.370 ;
        RECT 40.280 161.930 40.540 162.250 ;
        RECT 39.880 160.490 40.480 160.630 ;
        RECT 39.820 159.890 40.080 160.210 ;
        RECT 39.880 157.830 40.020 159.890 ;
        RECT 40.340 159.530 40.480 160.490 ;
        RECT 40.280 159.210 40.540 159.530 ;
        RECT 40.800 159.190 40.940 168.050 ;
        RECT 40.740 158.870 41.000 159.190 ;
        RECT 39.820 157.510 40.080 157.830 ;
        RECT 39.820 156.830 40.080 157.150 ;
        RECT 39.880 154.430 40.020 156.830 ;
        RECT 39.820 154.110 40.080 154.430 ;
        RECT 40.730 150.855 41.010 151.225 ;
        RECT 40.740 150.710 41.000 150.855 ;
        RECT 39.820 150.370 40.080 150.690 ;
        RECT 39.360 146.630 39.620 146.950 ;
        RECT 38.900 145.950 39.160 146.270 ;
        RECT 39.880 145.930 40.020 150.370 ;
        RECT 41.260 146.950 41.400 170.430 ;
        RECT 42.180 167.600 42.320 172.220 ;
        RECT 43.100 168.710 43.240 178.055 ;
        RECT 43.560 173.470 43.700 183.495 ;
        RECT 43.960 183.185 44.220 183.330 ;
        RECT 43.950 182.815 44.230 183.185 ;
        RECT 43.960 181.310 44.220 181.630 ;
        RECT 44.020 180.950 44.160 181.310 ;
        RECT 44.480 181.145 44.620 183.780 ;
        RECT 44.940 182.505 45.080 187.520 ;
        RECT 45.340 186.980 45.600 187.070 ;
        RECT 45.860 186.980 46.000 199.330 ;
        RECT 46.320 194.745 46.460 206.615 ;
        RECT 47.180 205.450 47.440 205.770 ;
        RECT 47.240 203.730 47.380 205.450 ;
        RECT 47.640 205.110 47.900 205.430 ;
        RECT 47.180 203.410 47.440 203.730 ;
        RECT 46.710 201.855 46.990 202.225 ;
        RECT 46.780 201.010 46.920 201.855 ;
        RECT 46.720 200.690 46.980 201.010 ;
        RECT 46.720 199.670 46.980 199.990 ;
        RECT 47.180 199.670 47.440 199.990 ;
        RECT 46.250 194.375 46.530 194.745 ;
        RECT 46.780 194.210 46.920 199.670 ;
        RECT 47.240 198.145 47.380 199.670 ;
        RECT 47.170 197.775 47.450 198.145 ;
        RECT 47.180 195.250 47.440 195.570 ;
        RECT 46.260 193.890 46.520 194.210 ;
        RECT 46.720 193.890 46.980 194.210 ;
        RECT 46.320 187.750 46.460 193.890 ;
        RECT 46.780 192.850 46.920 193.890 ;
        RECT 47.240 193.385 47.380 195.250 ;
        RECT 47.700 194.890 47.840 205.110 ;
        RECT 47.640 194.570 47.900 194.890 ;
        RECT 47.170 193.015 47.450 193.385 ;
        RECT 46.720 192.530 46.980 192.850 ;
        RECT 47.640 192.530 47.900 192.850 ;
        RECT 47.180 192.190 47.440 192.510 ;
        RECT 47.240 190.430 47.380 192.190 ;
        RECT 47.700 191.830 47.840 192.530 ;
        RECT 47.640 191.510 47.900 191.830 ;
        RECT 46.780 190.290 47.380 190.430 ;
        RECT 47.630 190.295 47.910 190.665 ;
        RECT 46.780 189.110 46.920 190.290 ;
        RECT 47.180 189.810 47.440 190.130 ;
        RECT 46.720 188.790 46.980 189.110 ;
        RECT 46.260 187.430 46.520 187.750 ;
        RECT 45.340 186.840 46.000 186.980 ;
        RECT 45.340 186.750 45.600 186.840 ;
        RECT 45.340 185.730 45.600 186.050 ;
        RECT 44.870 182.135 45.150 182.505 ;
        RECT 45.400 181.970 45.540 185.730 ;
        RECT 45.790 184.855 46.070 185.225 ;
        RECT 45.340 181.650 45.600 181.970 ;
        RECT 43.960 180.630 44.220 180.950 ;
        RECT 44.410 180.775 44.690 181.145 ;
        RECT 45.860 180.950 46.000 184.855 ;
        RECT 46.320 184.690 46.460 187.430 ;
        RECT 46.780 187.265 46.920 188.790 ;
        RECT 46.710 186.895 46.990 187.265 ;
        RECT 46.720 186.410 46.980 186.730 ;
        RECT 46.260 184.370 46.520 184.690 ;
        RECT 46.780 182.220 46.920 186.410 ;
        RECT 47.240 182.310 47.380 189.810 ;
        RECT 47.700 184.545 47.840 190.295 ;
        RECT 47.630 184.175 47.910 184.545 ;
        RECT 47.640 183.700 47.900 184.020 ;
        RECT 46.320 182.080 46.920 182.220 ;
        RECT 45.800 180.630 46.060 180.950 ;
        RECT 44.420 180.290 44.680 180.610 ;
        RECT 44.880 180.290 45.140 180.610 ;
        RECT 43.960 178.930 44.220 179.250 ;
        RECT 44.020 178.570 44.160 178.930 ;
        RECT 43.960 178.250 44.220 178.570 ;
        RECT 43.500 173.150 43.760 173.470 ;
        RECT 44.480 172.450 44.620 180.290 ;
        RECT 44.940 179.590 45.080 180.290 ;
        RECT 44.880 179.270 45.140 179.590 ;
        RECT 45.340 178.590 45.600 178.910 ;
        RECT 44.880 178.250 45.140 178.570 ;
        RECT 44.940 175.850 45.080 178.250 ;
        RECT 45.400 177.890 45.540 178.590 ;
        RECT 45.340 177.570 45.600 177.890 ;
        RECT 46.320 176.950 46.460 182.080 ;
        RECT 47.180 181.990 47.440 182.310 ;
        RECT 46.720 181.310 46.980 181.630 ;
        RECT 46.780 178.310 46.920 181.310 ;
        RECT 46.780 178.170 47.380 178.310 ;
        RECT 46.720 177.570 46.980 177.890 ;
        RECT 45.860 176.810 46.460 176.950 ;
        RECT 45.860 176.630 46.000 176.810 ;
        RECT 45.860 176.490 46.460 176.630 ;
        RECT 45.800 176.100 46.060 176.190 ;
        RECT 45.400 175.960 46.060 176.100 ;
        RECT 44.880 175.530 45.140 175.850 ;
        RECT 44.420 172.130 44.680 172.450 ;
        RECT 44.480 171.430 44.620 172.130 ;
        RECT 44.420 171.110 44.680 171.430 ;
        RECT 43.500 170.430 43.760 170.750 ;
        RECT 43.040 168.390 43.300 168.710 ;
        RECT 42.580 168.225 42.840 168.370 ;
        RECT 42.570 167.855 42.850 168.225 ;
        RECT 43.040 167.600 43.300 167.690 ;
        RECT 42.180 167.460 43.300 167.600 ;
        RECT 43.040 167.370 43.300 167.460 ;
        RECT 42.580 162.270 42.840 162.590 ;
        RECT 42.640 161.480 42.780 162.270 ;
        RECT 43.100 161.990 43.240 167.370 ;
        RECT 43.560 163.270 43.700 170.430 ;
        RECT 44.480 168.110 44.620 171.110 ;
        RECT 44.020 168.030 44.620 168.110 ;
        RECT 43.960 167.970 44.620 168.030 ;
        RECT 43.960 167.710 44.220 167.970 ;
        RECT 44.020 165.310 44.160 167.710 ;
        RECT 44.420 167.370 44.680 167.690 ;
        RECT 43.960 164.990 44.220 165.310 ;
        RECT 43.500 162.950 43.760 163.270 ;
        RECT 43.100 161.850 44.160 161.990 ;
        RECT 42.640 161.340 43.240 161.480 ;
        RECT 43.100 159.870 43.240 161.340 ;
        RECT 42.580 159.550 42.840 159.870 ;
        RECT 43.040 159.550 43.300 159.870 ;
        RECT 42.640 155.110 42.780 159.550 ;
        RECT 43.100 156.810 43.240 159.550 ;
        RECT 43.490 159.015 43.770 159.385 ;
        RECT 43.500 158.870 43.760 159.015 ;
        RECT 43.040 156.490 43.300 156.810 ;
        RECT 42.580 154.790 42.840 155.110 ;
        RECT 42.640 151.370 42.780 154.790 ;
        RECT 44.020 153.410 44.160 161.850 ;
        RECT 44.480 155.110 44.620 167.370 ;
        RECT 44.420 154.790 44.680 155.110 ;
        RECT 43.960 153.090 44.220 153.410 ;
        RECT 44.020 151.370 44.160 153.090 ;
        RECT 42.580 151.050 42.840 151.370 ;
        RECT 43.960 151.050 44.220 151.370 ;
        RECT 42.120 150.370 42.380 150.690 ;
        RECT 41.200 146.630 41.460 146.950 ;
        RECT 42.180 145.930 42.320 150.370 ;
        RECT 39.820 145.610 40.080 145.930 ;
        RECT 40.280 145.610 40.540 145.930 ;
        RECT 40.740 145.610 41.000 145.930 ;
        RECT 42.120 145.610 42.380 145.930 ;
        RECT 40.340 145.250 40.480 145.610 ;
        RECT 40.280 144.930 40.540 145.250 ;
        RECT 36.950 144.395 38.490 144.765 ;
        RECT 40.340 141.510 40.480 144.930 ;
        RECT 40.800 143.890 40.940 145.610 ;
        RECT 40.740 143.570 41.000 143.890 ;
        RECT 42.580 142.210 42.840 142.530 ;
        RECT 36.600 141.190 36.860 141.510 ;
        RECT 40.280 141.190 40.540 141.510 ;
        RECT 42.640 140.830 42.780 142.210 ;
        RECT 44.020 141.170 44.160 151.050 ;
        RECT 44.940 143.550 45.080 175.530 ;
        RECT 45.400 167.010 45.540 175.960 ;
        RECT 45.800 175.870 46.060 175.960 ;
        RECT 45.800 175.190 46.060 175.510 ;
        RECT 45.340 166.690 45.600 167.010 ;
        RECT 45.400 163.270 45.540 166.690 ;
        RECT 45.340 162.950 45.600 163.270 ;
        RECT 45.860 162.670 46.000 175.190 ;
        RECT 46.320 171.430 46.460 176.490 ;
        RECT 46.780 175.170 46.920 177.570 ;
        RECT 47.240 176.870 47.380 178.170 ;
        RECT 47.180 176.550 47.440 176.870 ;
        RECT 47.170 176.015 47.450 176.385 ;
        RECT 47.180 175.870 47.440 176.015 ;
        RECT 46.720 174.850 46.980 175.170 ;
        RECT 47.240 174.230 47.380 175.870 ;
        RECT 46.780 174.090 47.380 174.230 ;
        RECT 46.260 171.110 46.520 171.430 ;
        RECT 46.780 170.945 46.920 174.090 ;
        RECT 47.170 171.255 47.450 171.625 ;
        RECT 46.710 170.575 46.990 170.945 ;
        RECT 47.240 170.750 47.380 171.255 ;
        RECT 47.180 170.430 47.440 170.750 ;
        RECT 46.720 170.090 46.980 170.410 ;
        RECT 46.780 169.730 46.920 170.090 ;
        RECT 46.260 169.410 46.520 169.730 ;
        RECT 46.720 169.410 46.980 169.730 ;
        RECT 47.240 169.585 47.380 170.430 ;
        RECT 46.320 167.690 46.460 169.410 ;
        RECT 47.170 169.215 47.450 169.585 ;
        RECT 46.720 168.390 46.980 168.710 ;
        RECT 46.260 167.370 46.520 167.690 ;
        RECT 45.400 162.530 46.000 162.670 ;
        RECT 45.400 151.370 45.540 162.530 ;
        RECT 45.800 161.930 46.060 162.250 ;
        RECT 45.860 160.550 46.000 161.930 ;
        RECT 45.800 160.230 46.060 160.550 ;
        RECT 46.260 160.230 46.520 160.550 ;
        RECT 45.800 159.210 46.060 159.530 ;
        RECT 45.860 157.830 46.000 159.210 ;
        RECT 45.800 157.510 46.060 157.830 ;
        RECT 46.320 154.430 46.460 160.230 ;
        RECT 46.260 154.110 46.520 154.430 ;
        RECT 46.780 151.370 46.920 168.390 ;
        RECT 47.170 167.175 47.450 167.545 ;
        RECT 47.180 167.030 47.440 167.175 ;
        RECT 47.700 165.990 47.840 183.700 ;
        RECT 48.160 182.310 48.300 217.330 ;
        RECT 51.380 212.425 51.520 217.330 ;
        RECT 54.600 212.570 54.740 217.330 ;
        RECT 51.310 212.055 51.590 212.425 ;
        RECT 54.540 212.250 54.800 212.570 ;
        RECT 56.370 210.695 56.650 211.065 ;
        RECT 55.000 208.510 55.260 208.830 ;
        RECT 49.940 207.830 50.200 208.150 ;
        RECT 49.480 206.130 49.740 206.450 ;
        RECT 49.020 205.450 49.280 205.770 ;
        RECT 48.560 204.770 48.820 205.090 ;
        RECT 48.100 181.990 48.360 182.310 ;
        RECT 48.620 181.630 48.760 204.770 ;
        RECT 49.080 198.630 49.220 205.450 ;
        RECT 49.020 198.310 49.280 198.630 ;
        RECT 49.010 196.415 49.290 196.785 ;
        RECT 49.080 189.450 49.220 196.415 ;
        RECT 49.540 195.230 49.680 206.130 ;
        RECT 50.000 205.770 50.140 207.830 ;
        RECT 54.540 206.130 54.800 206.450 ;
        RECT 49.940 205.450 50.200 205.770 ;
        RECT 52.700 205.450 52.960 205.770 ;
        RECT 53.160 205.450 53.420 205.770 ;
        RECT 54.080 205.450 54.340 205.770 ;
        RECT 50.400 205.340 50.660 205.430 ;
        RECT 50.400 205.200 51.060 205.340 ;
        RECT 50.400 205.110 50.660 205.200 ;
        RECT 50.400 202.050 50.660 202.370 ;
        RECT 49.940 197.630 50.200 197.950 ;
        RECT 50.000 195.910 50.140 197.630 ;
        RECT 49.940 195.590 50.200 195.910 ;
        RECT 50.460 195.570 50.600 202.050 ;
        RECT 50.400 195.250 50.660 195.570 ;
        RECT 49.480 194.910 49.740 195.230 ;
        RECT 50.390 194.375 50.670 194.745 ;
        RECT 49.940 193.890 50.200 194.210 ;
        RECT 49.470 192.335 49.750 192.705 ;
        RECT 50.000 192.510 50.140 193.890 ;
        RECT 50.460 193.190 50.600 194.375 ;
        RECT 50.400 192.870 50.660 193.190 ;
        RECT 50.460 192.510 50.600 192.870 ;
        RECT 49.020 189.130 49.280 189.450 ;
        RECT 49.010 187.575 49.290 187.945 ;
        RECT 49.020 187.430 49.280 187.575 ;
        RECT 49.540 187.265 49.680 192.335 ;
        RECT 49.940 192.190 50.200 192.510 ;
        RECT 50.400 192.190 50.660 192.510 ;
        RECT 50.400 191.170 50.660 191.490 ;
        RECT 50.460 190.470 50.600 191.170 ;
        RECT 50.400 190.150 50.660 190.470 ;
        RECT 50.460 189.190 50.600 190.150 ;
        RECT 50.920 190.130 51.060 205.200 ;
        RECT 51.320 205.110 51.580 205.430 ;
        RECT 51.380 203.390 51.520 205.110 ;
        RECT 51.320 203.070 51.580 203.390 ;
        RECT 51.780 203.070 52.040 203.390 ;
        RECT 51.380 201.010 51.520 203.070 ;
        RECT 51.320 200.690 51.580 201.010 ;
        RECT 51.840 198.825 51.980 203.070 ;
        RECT 52.230 200.495 52.510 200.865 ;
        RECT 51.770 198.455 52.050 198.825 ;
        RECT 51.780 194.230 52.040 194.550 ;
        RECT 51.840 192.850 51.980 194.230 ;
        RECT 51.780 192.530 52.040 192.850 ;
        RECT 50.860 189.810 51.120 190.130 ;
        RECT 51.320 189.810 51.580 190.130 ;
        RECT 52.300 189.870 52.440 200.495 ;
        RECT 52.760 190.470 52.900 205.450 ;
        RECT 53.220 198.290 53.360 205.450 ;
        RECT 53.620 203.410 53.880 203.730 ;
        RECT 53.680 203.050 53.820 203.410 ;
        RECT 53.620 202.730 53.880 203.050 ;
        RECT 53.620 199.670 53.880 199.990 ;
        RECT 53.160 197.970 53.420 198.290 ;
        RECT 53.150 195.735 53.430 196.105 ;
        RECT 53.220 190.495 53.360 195.735 ;
        RECT 52.700 190.150 52.960 190.470 ;
        RECT 53.150 190.125 53.430 190.495 ;
        RECT 50.000 189.050 50.600 189.190 ;
        RECT 50.860 189.130 51.120 189.450 ;
        RECT 49.470 186.895 49.750 187.265 ;
        RECT 50.000 187.070 50.140 189.050 ;
        RECT 50.400 188.450 50.660 188.770 ;
        RECT 49.480 186.750 49.740 186.895 ;
        RECT 49.940 186.750 50.200 187.070 ;
        RECT 49.540 183.865 49.680 186.750 ;
        RECT 49.940 186.070 50.200 186.390 ;
        RECT 50.000 184.690 50.140 186.070 ;
        RECT 50.460 185.030 50.600 188.450 ;
        RECT 50.400 184.710 50.660 185.030 ;
        RECT 49.940 184.370 50.200 184.690 ;
        RECT 49.470 183.495 49.750 183.865 ;
        RECT 50.000 183.670 50.140 184.370 ;
        RECT 50.400 183.690 50.660 184.010 ;
        RECT 49.940 183.350 50.200 183.670 ;
        RECT 49.470 182.815 49.750 183.185 ;
        RECT 50.460 183.070 50.600 183.690 ;
        RECT 50.000 182.930 50.600 183.070 ;
        RECT 49.540 181.630 49.680 182.815 ;
        RECT 48.560 181.310 48.820 181.630 ;
        RECT 49.480 181.310 49.740 181.630 ;
        RECT 49.470 180.775 49.750 181.145 ;
        RECT 48.100 178.590 48.360 178.910 ;
        RECT 48.550 178.735 48.830 179.105 ;
        RECT 47.640 165.670 47.900 165.990 ;
        RECT 47.640 162.950 47.900 163.270 ;
        RECT 47.700 160.210 47.840 162.950 ;
        RECT 47.640 159.890 47.900 160.210 ;
        RECT 48.160 160.065 48.300 178.590 ;
        RECT 48.620 178.230 48.760 178.735 ;
        RECT 49.540 178.230 49.680 180.775 ;
        RECT 50.000 180.465 50.140 182.930 ;
        RECT 49.930 180.095 50.210 180.465 ;
        RECT 50.400 180.290 50.660 180.610 ;
        RECT 49.930 179.415 50.210 179.785 ;
        RECT 49.940 179.270 50.200 179.415 ;
        RECT 49.940 178.250 50.200 178.570 ;
        RECT 48.560 177.910 48.820 178.230 ;
        RECT 49.480 177.910 49.740 178.230 ;
        RECT 49.010 177.375 49.290 177.745 ;
        RECT 48.550 176.695 48.830 177.065 ;
        RECT 48.560 176.550 48.820 176.695 ;
        RECT 49.080 176.310 49.220 177.375 ;
        RECT 49.020 175.990 49.280 176.310 ;
        RECT 49.480 175.190 49.740 175.510 ;
        RECT 49.540 173.665 49.680 175.190 ;
        RECT 49.470 173.295 49.750 173.665 ;
        RECT 48.550 171.935 48.830 172.305 ;
        RECT 48.620 166.750 48.760 171.935 ;
        RECT 49.020 170.430 49.280 170.750 ;
        RECT 49.080 168.710 49.220 170.430 ;
        RECT 49.020 168.390 49.280 168.710 ;
        RECT 48.620 166.610 49.220 166.750 ;
        RECT 48.560 165.670 48.820 165.990 ;
        RECT 47.180 159.550 47.440 159.870 ;
        RECT 47.240 158.025 47.380 159.550 ;
        RECT 47.700 158.850 47.840 159.890 ;
        RECT 48.090 159.695 48.370 160.065 ;
        RECT 48.100 159.550 48.360 159.695 ;
        RECT 48.090 159.015 48.370 159.385 ;
        RECT 48.100 158.870 48.360 159.015 ;
        RECT 47.640 158.530 47.900 158.850 ;
        RECT 47.170 157.655 47.450 158.025 ;
        RECT 48.100 157.170 48.360 157.490 ;
        RECT 47.640 155.810 47.900 156.130 ;
        RECT 47.700 154.770 47.840 155.810 ;
        RECT 48.160 154.770 48.300 157.170 ;
        RECT 47.640 154.450 47.900 154.770 ;
        RECT 48.100 154.450 48.360 154.770 ;
        RECT 47.180 154.110 47.440 154.430 ;
        RECT 47.240 152.390 47.380 154.110 ;
        RECT 48.620 152.390 48.760 165.670 ;
        RECT 49.080 162.590 49.220 166.610 ;
        RECT 49.020 162.270 49.280 162.590 ;
        RECT 50.000 161.570 50.140 178.250 ;
        RECT 50.460 176.190 50.600 180.290 ;
        RECT 50.920 177.065 51.060 189.130 ;
        RECT 51.380 188.770 51.520 189.810 ;
        RECT 51.840 189.730 52.440 189.870 ;
        RECT 51.320 188.450 51.580 188.770 ;
        RECT 51.380 187.750 51.520 188.450 ;
        RECT 51.840 187.945 51.980 189.730 ;
        RECT 53.160 189.130 53.420 189.450 ;
        RECT 52.700 188.790 52.960 189.110 ;
        RECT 52.760 188.625 52.900 188.790 ;
        RECT 52.690 188.255 52.970 188.625 ;
        RECT 51.320 187.430 51.580 187.750 ;
        RECT 51.770 187.575 52.050 187.945 ;
        RECT 52.760 187.410 52.900 188.255 ;
        RECT 52.700 187.090 52.960 187.410 ;
        RECT 52.240 186.410 52.500 186.730 ;
        RECT 52.700 186.410 52.960 186.730 ;
        RECT 53.220 186.585 53.360 189.130 ;
        RECT 51.780 184.030 52.040 184.350 ;
        RECT 51.320 178.590 51.580 178.910 ;
        RECT 50.850 176.695 51.130 177.065 ;
        RECT 50.400 175.870 50.660 176.190 ;
        RECT 50.390 175.335 50.670 175.705 ;
        RECT 50.400 175.190 50.660 175.335 ;
        RECT 50.860 175.190 51.120 175.510 ;
        RECT 50.920 175.025 51.060 175.190 ;
        RECT 51.380 175.170 51.520 178.590 ;
        RECT 51.840 178.570 51.980 184.030 ;
        RECT 51.780 178.250 52.040 178.570 ;
        RECT 50.850 174.655 51.130 175.025 ;
        RECT 51.320 174.850 51.580 175.170 ;
        RECT 52.300 173.720 52.440 186.410 ;
        RECT 52.760 184.690 52.900 186.410 ;
        RECT 53.150 186.215 53.430 186.585 ;
        RECT 53.680 186.390 53.820 199.670 ;
        RECT 54.140 193.190 54.280 205.450 ;
        RECT 54.600 200.330 54.740 206.130 ;
        RECT 54.540 200.010 54.800 200.330 ;
        RECT 54.600 196.930 54.740 200.010 ;
        RECT 54.540 196.610 54.800 196.930 ;
        RECT 54.540 195.590 54.800 195.910 ;
        RECT 54.080 192.870 54.340 193.190 ;
        RECT 54.070 190.975 54.350 191.345 ;
        RECT 54.140 190.470 54.280 190.975 ;
        RECT 54.080 190.150 54.340 190.470 ;
        RECT 54.070 189.615 54.350 189.985 ;
        RECT 53.620 186.070 53.880 186.390 ;
        RECT 53.160 185.730 53.420 186.050 ;
        RECT 52.700 184.370 52.960 184.690 ;
        RECT 53.220 184.010 53.360 185.730 ;
        RECT 52.700 183.690 52.960 184.010 ;
        RECT 53.160 183.690 53.420 184.010 ;
        RECT 52.760 181.290 52.900 183.690 ;
        RECT 53.150 182.815 53.430 183.185 ;
        RECT 53.620 183.010 53.880 183.330 ;
        RECT 53.220 181.630 53.360 182.815 ;
        RECT 53.680 181.630 53.820 183.010 ;
        RECT 54.140 182.310 54.280 189.615 ;
        RECT 54.600 189.110 54.740 195.590 ;
        RECT 54.540 188.790 54.800 189.110 ;
        RECT 54.600 184.350 54.740 188.790 ;
        RECT 55.060 185.030 55.200 208.510 ;
        RECT 55.920 207.490 56.180 207.810 ;
        RECT 55.460 204.945 55.720 205.090 ;
        RECT 55.450 204.575 55.730 204.945 ;
        RECT 55.460 200.010 55.720 200.330 ;
        RECT 55.520 198.630 55.660 200.010 ;
        RECT 55.460 198.310 55.720 198.630 ;
        RECT 55.980 197.950 56.120 207.490 ;
        RECT 55.920 197.630 56.180 197.950 ;
        RECT 55.460 194.570 55.720 194.890 ;
        RECT 55.520 193.385 55.660 194.570 ;
        RECT 55.450 193.015 55.730 193.385 ;
        RECT 55.460 190.150 55.720 190.470 ;
        RECT 56.440 190.430 56.580 210.695 ;
        RECT 57.820 210.385 57.960 217.330 ;
        RECT 59.140 211.910 59.400 212.230 ;
        RECT 57.750 210.015 58.030 210.385 ;
        RECT 56.840 208.850 57.100 209.170 ;
        RECT 56.900 202.370 57.040 208.850 ;
        RECT 57.760 208.170 58.020 208.490 ;
        RECT 58.220 208.170 58.480 208.490 ;
        RECT 58.680 208.170 58.940 208.490 ;
        RECT 57.290 203.895 57.570 204.265 ;
        RECT 57.820 204.070 57.960 208.170 ;
        RECT 58.280 207.665 58.420 208.170 ;
        RECT 58.210 207.295 58.490 207.665 ;
        RECT 58.740 206.450 58.880 208.170 ;
        RECT 58.680 206.130 58.940 206.450 ;
        RECT 56.840 202.050 57.100 202.370 ;
        RECT 56.900 198.630 57.040 202.050 ;
        RECT 56.840 198.310 57.100 198.630 ;
        RECT 56.840 196.950 57.100 197.270 ;
        RECT 56.900 191.490 57.040 196.950 ;
        RECT 56.840 191.170 57.100 191.490 ;
        RECT 56.900 190.470 57.040 191.170 ;
        RECT 55.980 190.290 56.580 190.430 ;
        RECT 55.520 187.410 55.660 190.150 ;
        RECT 55.460 187.090 55.720 187.410 ;
        RECT 55.450 186.215 55.730 186.585 ;
        RECT 55.000 184.710 55.260 185.030 ;
        RECT 54.540 184.030 54.800 184.350 ;
        RECT 54.990 183.495 55.270 183.865 ;
        RECT 54.080 181.990 54.340 182.310 ;
        RECT 53.160 181.310 53.420 181.630 ;
        RECT 53.620 181.310 53.880 181.630 ;
        RECT 54.080 181.310 54.340 181.630 ;
        RECT 54.540 181.310 54.800 181.630 ;
        RECT 52.700 180.970 52.960 181.290 ;
        RECT 52.700 180.465 52.960 180.610 ;
        RECT 52.690 180.095 52.970 180.465 ;
        RECT 52.700 178.250 52.960 178.570 ;
        RECT 52.760 174.230 52.900 178.250 ;
        RECT 53.150 178.055 53.430 178.425 ;
        RECT 53.160 177.910 53.420 178.055 ;
        RECT 54.140 177.065 54.280 181.310 ;
        RECT 54.600 179.590 54.740 181.310 ;
        RECT 55.060 181.145 55.200 183.495 ;
        RECT 54.990 180.775 55.270 181.145 ;
        RECT 54.540 179.270 54.800 179.590 ;
        RECT 55.060 178.230 55.200 180.775 ;
        RECT 55.000 177.910 55.260 178.230 ;
        RECT 53.150 176.695 53.430 177.065 ;
        RECT 54.070 176.695 54.350 177.065 ;
        RECT 53.160 176.550 53.420 176.695 ;
        RECT 53.160 175.870 53.420 176.190 ;
        RECT 53.620 175.870 53.880 176.190 ;
        RECT 54.070 176.015 54.350 176.385 ;
        RECT 54.080 175.870 54.340 176.015 ;
        RECT 53.220 175.705 53.360 175.870 ;
        RECT 53.150 175.335 53.430 175.705 ;
        RECT 52.760 174.090 53.360 174.230 ;
        RECT 53.220 173.810 53.360 174.090 ;
        RECT 52.300 173.580 52.900 173.720 ;
        RECT 51.310 171.935 51.590 172.305 ;
        RECT 51.780 172.130 52.040 172.450 ;
        RECT 52.760 172.360 52.900 173.580 ;
        RECT 53.160 173.490 53.420 173.810 ;
        RECT 53.160 172.810 53.420 173.130 ;
        RECT 53.680 172.985 53.820 175.870 ;
        RECT 55.520 175.590 55.660 186.215 ;
        RECT 55.980 183.330 56.120 190.290 ;
        RECT 56.840 190.150 57.100 190.470 ;
        RECT 57.360 189.870 57.500 203.895 ;
        RECT 57.760 203.750 58.020 204.070 ;
        RECT 57.820 198.825 57.960 203.750 ;
        RECT 58.680 203.410 58.940 203.730 ;
        RECT 58.740 201.010 58.880 203.410 ;
        RECT 59.200 202.905 59.340 211.910 ;
        RECT 61.040 211.630 61.180 217.330 ;
        RECT 64.260 214.465 64.400 217.330 ;
        RECT 64.190 214.095 64.470 214.465 ;
        RECT 67.480 213.785 67.620 217.330 ;
        RECT 70.700 217.070 70.840 217.330 ;
        RECT 71.160 217.070 71.300 217.610 ;
        RECT 70.700 216.930 71.300 217.070 ;
        RECT 67.410 213.415 67.690 213.785 ;
        RECT 68.790 213.415 69.070 213.785 ;
        RECT 59.600 211.230 59.860 211.550 ;
        RECT 60.580 211.490 61.180 211.630 ;
        RECT 59.130 202.535 59.410 202.905 ;
        RECT 58.680 200.690 58.940 201.010 ;
        RECT 59.140 200.690 59.400 201.010 ;
        RECT 58.220 200.010 58.480 200.330 ;
        RECT 58.680 200.010 58.940 200.330 ;
        RECT 57.750 198.455 58.030 198.825 ;
        RECT 58.280 198.290 58.420 200.010 ;
        RECT 58.220 197.970 58.480 198.290 ;
        RECT 58.740 197.465 58.880 200.010 ;
        RECT 58.670 197.095 58.950 197.465 ;
        RECT 58.680 196.610 58.940 196.930 ;
        RECT 58.220 191.850 58.480 192.170 ;
        RECT 57.760 191.170 58.020 191.490 ;
        RECT 57.820 190.470 57.960 191.170 ;
        RECT 57.760 190.150 58.020 190.470 ;
        RECT 57.360 189.730 57.960 189.870 ;
        RECT 56.380 189.130 56.640 189.450 ;
        RECT 56.440 185.905 56.580 189.130 ;
        RECT 57.300 186.750 57.560 187.070 ;
        RECT 56.840 186.410 57.100 186.730 ;
        RECT 56.370 185.535 56.650 185.905 ;
        RECT 56.900 185.030 57.040 186.410 ;
        RECT 56.840 184.710 57.100 185.030 ;
        RECT 56.370 183.495 56.650 183.865 ;
        RECT 55.920 183.010 56.180 183.330 ;
        RECT 55.920 181.310 56.180 181.630 ;
        RECT 55.980 181.145 56.120 181.310 ;
        RECT 55.910 180.775 56.190 181.145 ;
        RECT 55.920 180.290 56.180 180.610 ;
        RECT 55.980 179.785 56.120 180.290 ;
        RECT 55.910 179.415 56.190 179.785 ;
        RECT 55.910 178.735 56.190 179.105 ;
        RECT 55.980 176.190 56.120 178.735 ;
        RECT 56.440 176.190 56.580 183.495 ;
        RECT 56.840 181.650 57.100 181.970 ;
        RECT 56.900 178.570 57.040 181.650 ;
        RECT 56.840 178.250 57.100 178.570 ;
        RECT 57.360 176.950 57.500 186.750 ;
        RECT 56.900 176.810 57.500 176.950 ;
        RECT 55.920 175.870 56.180 176.190 ;
        RECT 56.380 175.870 56.640 176.190 ;
        RECT 55.060 175.510 55.660 175.590 ;
        RECT 55.000 175.450 55.660 175.510 ;
        RECT 55.980 175.590 56.120 175.870 ;
        RECT 55.980 175.450 56.580 175.590 ;
        RECT 55.000 175.190 55.260 175.450 ;
        RECT 55.920 174.850 56.180 175.170 ;
        RECT 55.460 173.830 55.720 174.150 ;
        RECT 55.000 173.490 55.260 173.810 ;
        RECT 52.300 172.220 52.900 172.360 ;
        RECT 50.850 171.255 51.130 171.625 ;
        RECT 50.920 168.370 51.060 171.255 ;
        RECT 50.860 168.050 51.120 168.370 ;
        RECT 50.400 167.370 50.660 167.690 ;
        RECT 49.940 161.250 50.200 161.570 ;
        RECT 49.940 160.065 50.200 160.210 ;
        RECT 49.930 159.695 50.210 160.065 ;
        RECT 49.940 159.210 50.200 159.530 ;
        RECT 49.480 158.530 49.740 158.850 ;
        RECT 49.020 156.490 49.280 156.810 ;
        RECT 49.080 154.430 49.220 156.490 ;
        RECT 49.540 154.430 49.680 158.530 ;
        RECT 50.000 158.025 50.140 159.210 ;
        RECT 49.930 157.655 50.210 158.025 ;
        RECT 50.000 154.430 50.140 157.655 ;
        RECT 49.020 154.110 49.280 154.430 ;
        RECT 49.480 154.110 49.740 154.430 ;
        RECT 49.940 154.110 50.200 154.430 ;
        RECT 47.180 152.070 47.440 152.390 ;
        RECT 48.560 152.070 48.820 152.390 ;
        RECT 45.340 151.050 45.600 151.370 ;
        RECT 46.720 151.050 46.980 151.370 ;
        RECT 45.400 145.930 45.540 151.050 ;
        RECT 46.780 145.930 46.920 151.050 ;
        RECT 45.340 145.610 45.600 145.930 ;
        RECT 46.720 145.610 46.980 145.930 ;
        RECT 45.400 144.230 45.540 145.610 ;
        RECT 45.340 143.910 45.600 144.230 ;
        RECT 44.880 143.230 45.140 143.550 ;
        RECT 44.940 141.510 45.080 143.230 ;
        RECT 45.400 141.510 45.540 143.910 ;
        RECT 46.780 143.890 46.920 145.610 ;
        RECT 46.720 143.570 46.980 143.890 ;
        RECT 49.540 143.550 49.680 154.110 ;
        RECT 50.000 149.670 50.140 154.110 ;
        RECT 49.940 149.350 50.200 149.670 ;
        RECT 50.460 148.310 50.600 167.370 ;
        RECT 50.860 163.970 51.120 164.290 ;
        RECT 50.920 158.850 51.060 163.970 ;
        RECT 50.860 158.530 51.120 158.850 ;
        RECT 50.920 156.810 51.060 158.530 ;
        RECT 50.860 156.490 51.120 156.810 ;
        RECT 51.380 152.050 51.520 171.935 ;
        RECT 51.840 171.625 51.980 172.130 ;
        RECT 51.770 171.255 52.050 171.625 ;
        RECT 51.770 170.575 52.050 170.945 ;
        RECT 51.840 165.390 51.980 170.575 ;
        RECT 52.300 170.070 52.440 172.220 ;
        RECT 52.700 170.770 52.960 171.090 ;
        RECT 52.240 169.750 52.500 170.070 ;
        RECT 52.760 165.990 52.900 170.770 ;
        RECT 53.220 168.370 53.360 172.810 ;
        RECT 53.610 172.615 53.890 172.985 ;
        RECT 54.540 172.470 54.800 172.790 ;
        RECT 53.620 172.130 53.880 172.450 ;
        RECT 54.080 172.130 54.340 172.450 ;
        RECT 53.680 171.625 53.820 172.130 ;
        RECT 53.610 171.255 53.890 171.625 ;
        RECT 54.140 171.090 54.280 172.130 ;
        RECT 54.600 171.090 54.740 172.470 ;
        RECT 54.080 170.770 54.340 171.090 ;
        RECT 54.540 170.770 54.800 171.090 ;
        RECT 53.620 170.430 53.880 170.750 ;
        RECT 53.160 168.050 53.420 168.370 ;
        RECT 53.680 167.350 53.820 170.430 ;
        RECT 53.620 167.030 53.880 167.350 ;
        RECT 53.160 166.690 53.420 167.010 ;
        RECT 52.700 165.670 52.960 165.990 ;
        RECT 51.840 165.250 52.900 165.390 ;
        RECT 51.780 161.930 52.040 162.250 ;
        RECT 51.840 160.550 51.980 161.930 ;
        RECT 52.240 161.250 52.500 161.570 ;
        RECT 51.780 160.230 52.040 160.550 ;
        RECT 52.300 156.810 52.440 161.250 ;
        RECT 52.240 156.490 52.500 156.810 ;
        RECT 52.760 154.770 52.900 165.250 ;
        RECT 53.220 160.210 53.360 166.690 ;
        RECT 54.600 165.650 54.740 170.770 ;
        RECT 55.060 169.585 55.200 173.490 ;
        RECT 55.520 173.470 55.660 173.830 ;
        RECT 55.460 173.150 55.720 173.470 ;
        RECT 55.980 173.130 56.120 174.850 ;
        RECT 55.920 172.810 56.180 173.130 ;
        RECT 56.440 172.790 56.580 175.450 ;
        RECT 56.380 172.470 56.640 172.790 ;
        RECT 55.460 172.130 55.720 172.450 ;
        RECT 54.990 169.215 55.270 169.585 ;
        RECT 55.000 166.690 55.260 167.010 ;
        RECT 54.540 165.390 54.800 165.650 ;
        RECT 53.680 165.330 54.800 165.390 ;
        RECT 53.680 165.250 54.740 165.330 ;
        RECT 55.060 165.310 55.200 166.690 ;
        RECT 55.520 165.990 55.660 172.130 ;
        RECT 56.370 171.935 56.650 172.305 ;
        RECT 55.920 170.430 56.180 170.750 ;
        RECT 55.460 165.670 55.720 165.990 ;
        RECT 55.980 165.310 56.120 170.430 ;
        RECT 53.680 164.970 53.820 165.250 ;
        RECT 55.000 164.990 55.260 165.310 ;
        RECT 55.920 164.990 56.180 165.310 ;
        RECT 53.620 164.650 53.880 164.970 ;
        RECT 55.980 163.270 56.120 164.990 ;
        RECT 55.920 162.950 56.180 163.270 ;
        RECT 54.080 161.930 54.340 162.250 ;
        RECT 53.620 161.250 53.880 161.570 ;
        RECT 53.680 160.210 53.820 161.250 ;
        RECT 53.160 159.890 53.420 160.210 ;
        RECT 53.620 159.890 53.880 160.210 ;
        RECT 53.220 159.190 53.360 159.890 ;
        RECT 53.160 158.870 53.420 159.190 ;
        RECT 54.140 158.850 54.280 161.930 ;
        RECT 55.000 161.590 55.260 161.910 ;
        RECT 55.060 160.550 55.200 161.590 ;
        RECT 56.440 160.550 56.580 171.935 ;
        RECT 56.900 171.430 57.040 176.810 ;
        RECT 57.290 172.615 57.570 172.985 ;
        RECT 56.840 171.110 57.100 171.430 ;
        RECT 57.360 166.070 57.500 172.615 ;
        RECT 57.820 171.430 57.960 189.730 ;
        RECT 58.280 186.730 58.420 191.850 ;
        RECT 58.220 186.410 58.480 186.730 ;
        RECT 58.210 182.135 58.490 182.505 ;
        RECT 58.280 179.590 58.420 182.135 ;
        RECT 58.220 179.270 58.480 179.590 ;
        RECT 58.740 178.990 58.880 196.610 ;
        RECT 59.200 189.450 59.340 200.690 ;
        RECT 59.660 200.185 59.800 211.230 ;
        RECT 60.580 206.110 60.720 211.490 ;
        RECT 61.440 210.890 61.700 211.210 ;
        RECT 60.980 208.510 61.240 208.830 ;
        RECT 60.520 205.790 60.780 206.110 ;
        RECT 61.040 205.430 61.180 208.510 ;
        RECT 61.500 205.770 61.640 210.890 ;
        RECT 62.820 209.190 63.080 209.510 ;
        RECT 67.420 209.190 67.680 209.510 ;
        RECT 61.440 205.450 61.700 205.770 ;
        RECT 60.980 205.110 61.240 205.430 ;
        RECT 61.500 203.980 61.640 205.450 ;
        RECT 60.120 203.840 61.640 203.980 ;
        RECT 60.120 200.330 60.260 203.840 ;
        RECT 60.980 203.070 61.240 203.390 ;
        RECT 60.520 202.730 60.780 203.050 ;
        RECT 59.590 199.815 59.870 200.185 ;
        RECT 60.060 200.010 60.320 200.330 ;
        RECT 60.120 195.910 60.260 200.010 ;
        RECT 60.580 199.990 60.720 202.730 ;
        RECT 60.520 199.670 60.780 199.990 ;
        RECT 60.520 197.290 60.780 197.610 ;
        RECT 60.580 196.785 60.720 197.290 ;
        RECT 60.510 196.415 60.790 196.785 ;
        RECT 60.060 195.590 60.320 195.910 ;
        RECT 60.060 192.530 60.320 192.850 ;
        RECT 59.600 192.190 59.860 192.510 ;
        RECT 59.140 189.130 59.400 189.450 ;
        RECT 59.140 187.090 59.400 187.410 ;
        RECT 59.200 183.330 59.340 187.090 ;
        RECT 59.660 184.690 59.800 192.190 ;
        RECT 60.120 187.410 60.260 192.530 ;
        RECT 61.040 191.490 61.180 203.070 ;
        RECT 61.440 202.730 61.700 203.050 ;
        RECT 61.500 199.650 61.640 202.730 ;
        RECT 61.900 202.390 62.160 202.710 ;
        RECT 61.440 199.330 61.700 199.650 ;
        RECT 60.980 191.170 61.240 191.490 ;
        RECT 60.970 190.295 61.250 190.665 ;
        RECT 61.040 190.130 61.180 190.295 ;
        RECT 60.980 189.810 61.240 190.130 ;
        RECT 60.060 187.090 60.320 187.410 ;
        RECT 60.060 186.410 60.320 186.730 ;
        RECT 59.600 184.370 59.860 184.690 ;
        RECT 59.140 183.010 59.400 183.330 ;
        RECT 60.120 182.310 60.260 186.410 ;
        RECT 61.040 184.010 61.180 189.810 ;
        RECT 61.500 189.450 61.640 199.330 ;
        RECT 61.960 197.950 62.100 202.390 ;
        RECT 62.360 199.330 62.620 199.650 ;
        RECT 61.900 197.630 62.160 197.950 ;
        RECT 62.420 197.610 62.560 199.330 ;
        RECT 62.880 197.950 63.020 209.190 ;
        RECT 66.040 208.850 66.300 209.170 ;
        RECT 63.740 205.110 64.000 205.430 ;
        RECT 63.280 200.010 63.540 200.330 ;
        RECT 62.820 197.630 63.080 197.950 ;
        RECT 62.360 197.290 62.620 197.610 ;
        RECT 62.820 196.950 63.080 197.270 ;
        RECT 62.880 195.230 63.020 196.950 ;
        RECT 62.820 194.910 63.080 195.230 ;
        RECT 61.900 194.570 62.160 194.890 ;
        RECT 61.960 191.490 62.100 194.570 ;
        RECT 61.900 191.170 62.160 191.490 ;
        RECT 63.340 191.345 63.480 200.010 ;
        RECT 63.800 199.650 63.940 205.110 ;
        RECT 65.120 203.070 65.380 203.390 ;
        RECT 64.200 202.730 64.460 203.050 ;
        RECT 63.740 199.330 64.000 199.650 ;
        RECT 63.800 197.950 63.940 199.330 ;
        RECT 63.740 197.630 64.000 197.950 ;
        RECT 63.740 196.950 64.000 197.270 ;
        RECT 63.270 190.975 63.550 191.345 ;
        RECT 61.890 190.295 62.170 190.665 ;
        RECT 61.960 189.450 62.100 190.295 ;
        RECT 63.800 189.870 63.940 196.950 ;
        RECT 64.260 196.670 64.400 202.730 ;
        RECT 64.260 196.530 64.860 196.670 ;
        RECT 64.200 193.890 64.460 194.210 ;
        RECT 63.340 189.730 63.940 189.870 ;
        RECT 61.440 189.130 61.700 189.450 ;
        RECT 61.900 189.130 62.160 189.450 ;
        RECT 61.500 186.050 61.640 189.130 ;
        RECT 61.440 185.730 61.700 186.050 ;
        RECT 61.430 184.855 61.710 185.225 ;
        RECT 60.980 183.690 61.240 184.010 ;
        RECT 61.500 182.310 61.640 184.855 ;
        RECT 60.060 181.990 60.320 182.310 ;
        RECT 60.980 181.990 61.240 182.310 ;
        RECT 61.440 181.990 61.700 182.310 ;
        RECT 59.600 180.970 59.860 181.290 ;
        RECT 59.660 179.250 59.800 180.970 ;
        RECT 61.040 180.610 61.180 181.990 ;
        RECT 61.430 181.455 61.710 181.825 ;
        RECT 61.440 181.310 61.700 181.455 ;
        RECT 61.960 181.290 62.100 189.130 ;
        RECT 63.340 187.265 63.480 189.730 ;
        RECT 64.260 189.450 64.400 193.890 ;
        RECT 63.740 189.130 64.000 189.450 ;
        RECT 64.200 189.130 64.460 189.450 ;
        RECT 63.270 186.895 63.550 187.265 ;
        RECT 62.350 185.535 62.630 185.905 ;
        RECT 62.820 185.730 63.080 186.050 ;
        RECT 62.420 182.310 62.560 185.535 ;
        RECT 62.360 181.990 62.620 182.310 ;
        RECT 61.900 180.970 62.160 181.290 ;
        RECT 60.980 180.290 61.240 180.610 ;
        RECT 61.900 180.290 62.160 180.610 ;
        RECT 58.280 178.850 58.880 178.990 ;
        RECT 59.600 178.930 59.860 179.250 ;
        RECT 60.520 178.930 60.780 179.250 ;
        RECT 61.040 179.105 61.180 180.290 ;
        RECT 61.430 179.415 61.710 179.785 ;
        RECT 58.280 175.170 58.420 178.850 ;
        RECT 58.670 178.055 58.950 178.425 ;
        RECT 59.600 178.250 59.860 178.570 ;
        RECT 58.680 177.910 58.940 178.055 ;
        RECT 58.740 177.065 58.880 177.910 ;
        RECT 58.670 176.695 58.950 177.065 ;
        RECT 59.660 176.440 59.800 178.250 ;
        RECT 60.580 177.065 60.720 178.930 ;
        RECT 60.970 178.735 61.250 179.105 ;
        RECT 61.500 178.570 61.640 179.415 ;
        RECT 61.960 178.570 62.100 180.290 ;
        RECT 61.440 178.480 61.700 178.570 ;
        RECT 61.040 178.340 61.700 178.480 ;
        RECT 60.510 176.695 60.790 177.065 ;
        RECT 60.060 176.440 60.320 176.530 ;
        RECT 58.670 176.015 58.950 176.385 ;
        RECT 59.660 176.300 60.320 176.440 ;
        RECT 60.060 176.210 60.320 176.300 ;
        RECT 58.220 174.850 58.480 175.170 ;
        RECT 58.220 173.490 58.480 173.810 ;
        RECT 58.280 172.985 58.420 173.490 ;
        RECT 58.210 172.615 58.490 172.985 ;
        RECT 58.220 172.130 58.480 172.450 ;
        RECT 58.280 171.430 58.420 172.130 ;
        RECT 57.760 171.110 58.020 171.430 ;
        RECT 58.220 171.110 58.480 171.430 ;
        RECT 58.740 170.750 58.880 176.015 ;
        RECT 59.140 175.530 59.400 175.850 ;
        RECT 59.200 175.170 59.340 175.530 ;
        RECT 59.590 175.335 59.870 175.705 ;
        RECT 59.140 174.850 59.400 175.170 ;
        RECT 58.680 170.430 58.940 170.750 ;
        RECT 59.200 170.150 59.340 174.850 ;
        RECT 59.660 172.450 59.800 175.335 ;
        RECT 60.120 173.130 60.260 176.210 ;
        RECT 60.510 176.015 60.790 176.385 ;
        RECT 61.040 176.190 61.180 178.340 ;
        RECT 61.440 178.250 61.700 178.340 ;
        RECT 61.900 178.250 62.160 178.570 ;
        RECT 60.060 172.810 60.320 173.130 ;
        RECT 59.600 172.130 59.860 172.450 ;
        RECT 60.060 172.305 60.320 172.450 ;
        RECT 60.050 171.935 60.330 172.305 ;
        RECT 60.060 170.660 60.320 170.750 ;
        RECT 60.580 170.660 60.720 176.015 ;
        RECT 60.980 175.870 61.240 176.190 ;
        RECT 61.440 176.100 61.700 176.190 ;
        RECT 61.960 176.100 62.100 178.250 ;
        RECT 62.360 177.910 62.620 178.230 ;
        RECT 62.420 176.190 62.560 177.910 ;
        RECT 61.440 175.960 62.100 176.100 ;
        RECT 61.440 175.870 61.700 175.960 ;
        RECT 62.360 175.870 62.620 176.190 ;
        RECT 61.440 174.850 61.700 175.170 ;
        RECT 60.980 172.130 61.240 172.450 ;
        RECT 61.040 170.750 61.180 172.130 ;
        RECT 60.060 170.520 60.720 170.660 ;
        RECT 60.060 170.430 60.320 170.520 ;
        RECT 60.980 170.430 61.240 170.750 ;
        RECT 59.200 170.010 60.720 170.150 ;
        RECT 58.220 168.390 58.480 168.710 ;
        RECT 57.360 165.930 57.960 166.070 ;
        RECT 57.300 164.990 57.560 165.310 ;
        RECT 56.840 164.650 57.100 164.970 ;
        RECT 55.000 160.230 55.260 160.550 ;
        RECT 56.380 160.230 56.640 160.550 ;
        RECT 56.440 159.870 56.580 160.230 ;
        RECT 56.380 159.550 56.640 159.870 ;
        RECT 55.460 158.870 55.720 159.190 ;
        RECT 54.080 158.530 54.340 158.850 ;
        RECT 53.620 157.400 53.880 157.490 ;
        RECT 53.620 157.260 55.200 157.400 ;
        RECT 53.620 157.170 53.880 157.260 ;
        RECT 52.700 154.450 52.960 154.770 ;
        RECT 54.080 154.110 54.340 154.430 ;
        RECT 53.620 153.770 53.880 154.090 ;
        RECT 53.680 153.410 53.820 153.770 ;
        RECT 53.160 153.090 53.420 153.410 ;
        RECT 53.620 153.090 53.880 153.410 ;
        RECT 51.320 151.730 51.580 152.050 ;
        RECT 52.240 151.390 52.500 151.710 ;
        RECT 52.300 151.030 52.440 151.390 ;
        RECT 53.220 151.370 53.360 153.090 ;
        RECT 53.160 151.050 53.420 151.370 ;
        RECT 51.780 150.710 52.040 151.030 ;
        RECT 52.240 150.710 52.500 151.030 ;
        RECT 51.840 149.330 51.980 150.710 ;
        RECT 51.780 149.010 52.040 149.330 ;
        RECT 52.300 148.990 52.440 150.710 ;
        RECT 54.140 148.990 54.280 154.110 ;
        RECT 55.060 153.750 55.200 157.260 ;
        RECT 55.520 157.150 55.660 158.870 ;
        RECT 55.460 156.830 55.720 157.150 ;
        RECT 55.000 153.430 55.260 153.750 ;
        RECT 55.460 153.430 55.720 153.750 ;
        RECT 54.540 151.730 54.800 152.050 ;
        RECT 55.060 151.790 55.200 153.430 ;
        RECT 55.520 152.390 55.660 153.430 ;
        RECT 55.460 152.070 55.720 152.390 ;
        RECT 55.920 151.790 56.180 152.050 ;
        RECT 55.060 151.730 56.180 151.790 ;
        RECT 54.600 151.280 54.740 151.730 ;
        RECT 55.060 151.650 56.120 151.730 ;
        RECT 55.000 151.280 55.260 151.370 ;
        RECT 54.600 151.140 55.260 151.280 ;
        RECT 55.000 151.050 55.260 151.140 ;
        RECT 52.240 148.670 52.500 148.990 ;
        RECT 54.080 148.670 54.340 148.990 ;
        RECT 55.000 148.670 55.260 148.990 ;
        RECT 50.400 147.990 50.660 148.310 ;
        RECT 55.060 147.970 55.200 148.670 ;
        RECT 55.000 147.650 55.260 147.970 ;
        RECT 55.520 145.930 55.660 151.650 ;
        RECT 55.920 150.370 56.180 150.690 ;
        RECT 55.980 148.990 56.120 150.370 ;
        RECT 56.900 149.330 57.040 164.650 ;
        RECT 57.360 152.390 57.500 164.990 ;
        RECT 57.300 152.070 57.560 152.390 ;
        RECT 57.300 150.710 57.560 151.030 ;
        RECT 56.840 149.010 57.100 149.330 ;
        RECT 57.360 148.990 57.500 150.710 ;
        RECT 55.920 148.670 56.180 148.990 ;
        RECT 57.300 148.670 57.560 148.990 ;
        RECT 57.360 146.950 57.500 148.670 ;
        RECT 57.300 146.630 57.560 146.950 ;
        RECT 57.820 146.270 57.960 165.930 ;
        RECT 58.280 165.310 58.420 168.390 ;
        RECT 58.680 167.370 58.940 167.690 ;
        RECT 60.060 167.370 60.320 167.690 ;
        RECT 58.220 164.990 58.480 165.310 ;
        RECT 58.740 162.590 58.880 167.370 ;
        RECT 59.140 164.990 59.400 165.310 ;
        RECT 58.680 162.270 58.940 162.590 ;
        RECT 58.220 159.210 58.480 159.530 ;
        RECT 58.280 156.810 58.420 159.210 ;
        RECT 58.680 158.870 58.940 159.190 ;
        RECT 58.220 156.490 58.480 156.810 ;
        RECT 58.740 156.130 58.880 158.870 ;
        RECT 59.200 156.130 59.340 164.990 ;
        RECT 60.120 162.250 60.260 167.370 ;
        RECT 60.580 165.310 60.720 170.010 ;
        RECT 61.040 165.650 61.180 170.430 ;
        RECT 61.500 170.410 61.640 174.850 ;
        RECT 61.890 173.975 62.170 174.345 ;
        RECT 61.960 172.450 62.100 173.975 ;
        RECT 62.360 172.810 62.620 173.130 ;
        RECT 61.900 172.130 62.160 172.450 ;
        RECT 62.420 170.945 62.560 172.810 ;
        RECT 62.350 170.575 62.630 170.945 ;
        RECT 61.440 170.090 61.700 170.410 ;
        RECT 60.980 165.330 61.240 165.650 ;
        RECT 60.520 164.990 60.780 165.310 ;
        RECT 60.580 163.270 60.720 164.990 ;
        RECT 60.520 162.950 60.780 163.270 ;
        RECT 60.060 161.930 60.320 162.250 ;
        RECT 58.680 155.810 58.940 156.130 ;
        RECT 59.140 155.810 59.400 156.130 ;
        RECT 60.120 155.110 60.260 161.930 ;
        RECT 60.520 159.890 60.780 160.210 ;
        RECT 60.580 158.850 60.720 159.890 ;
        RECT 60.520 158.530 60.780 158.850 ;
        RECT 60.060 154.790 60.320 155.110 ;
        RECT 60.060 153.430 60.320 153.750 ;
        RECT 58.680 152.070 58.940 152.390 ;
        RECT 58.220 151.050 58.480 151.370 ;
        RECT 58.280 148.990 58.420 151.050 ;
        RECT 58.220 148.670 58.480 148.990 ;
        RECT 58.740 147.970 58.880 152.070 ;
        RECT 60.120 151.370 60.260 153.430 ;
        RECT 60.980 153.090 61.240 153.410 ;
        RECT 61.040 151.370 61.180 153.090 ;
        RECT 59.140 151.280 59.400 151.370 ;
        RECT 59.140 151.140 59.800 151.280 ;
        RECT 59.140 151.050 59.400 151.140 ;
        RECT 59.660 148.990 59.800 151.140 ;
        RECT 60.060 151.050 60.320 151.370 ;
        RECT 60.980 151.050 61.240 151.370 ;
        RECT 60.120 149.330 60.260 151.050 ;
        RECT 60.060 149.010 60.320 149.330 ;
        RECT 59.600 148.670 59.860 148.990 ;
        RECT 60.060 148.330 60.320 148.650 ;
        RECT 58.680 147.650 58.940 147.970 ;
        RECT 57.760 145.950 58.020 146.270 ;
        RECT 55.460 145.610 55.720 145.930 ;
        RECT 49.480 143.230 49.740 143.550 ;
        RECT 57.820 142.870 57.960 145.950 ;
        RECT 60.120 143.890 60.260 148.330 ;
        RECT 61.040 146.950 61.180 151.050 ;
        RECT 60.980 146.630 61.240 146.950 ;
        RECT 61.040 145.590 61.180 146.630 ;
        RECT 61.500 145.930 61.640 170.090 ;
        RECT 61.900 169.980 62.160 170.070 ;
        RECT 62.420 169.980 62.560 170.575 ;
        RECT 61.900 169.840 62.560 169.980 ;
        RECT 61.900 169.750 62.160 169.840 ;
        RECT 62.880 168.905 63.020 185.730 ;
        RECT 63.800 182.310 63.940 189.130 ;
        RECT 64.720 186.050 64.860 196.530 ;
        RECT 65.180 187.750 65.320 203.070 ;
        RECT 65.580 202.730 65.840 203.050 ;
        RECT 65.640 190.665 65.780 202.730 ;
        RECT 66.100 201.545 66.240 208.850 ;
        RECT 67.480 206.790 67.620 209.190 ;
        RECT 68.340 207.490 68.600 207.810 ;
        RECT 67.420 206.470 67.680 206.790 ;
        RECT 67.880 205.625 68.140 205.770 ;
        RECT 67.870 205.255 68.150 205.625 ;
        RECT 67.420 203.410 67.680 203.730 ;
        RECT 66.960 202.730 67.220 203.050 ;
        RECT 66.500 202.050 66.760 202.370 ;
        RECT 66.030 201.175 66.310 201.545 ;
        RECT 66.560 194.210 66.700 202.050 ;
        RECT 67.020 197.465 67.160 202.730 ;
        RECT 66.950 197.095 67.230 197.465 ;
        RECT 67.480 196.670 67.620 203.410 ;
        RECT 67.880 203.070 68.140 203.390 ;
        RECT 67.020 196.530 67.620 196.670 ;
        RECT 66.500 193.890 66.760 194.210 ;
        RECT 65.570 190.295 65.850 190.665 ;
        RECT 65.120 187.430 65.380 187.750 ;
        RECT 65.580 186.410 65.840 186.730 ;
        RECT 64.660 185.730 64.920 186.050 ;
        RECT 65.640 185.030 65.780 186.410 ;
        RECT 65.580 184.710 65.840 185.030 ;
        RECT 64.200 183.010 64.460 183.330 ;
        RECT 63.740 181.990 64.000 182.310 ;
        RECT 63.740 181.540 64.000 181.630 ;
        RECT 64.260 181.540 64.400 183.010 ;
        RECT 63.740 181.400 64.400 181.540 ;
        RECT 64.650 181.455 64.930 181.825 ;
        RECT 65.640 181.630 65.780 184.710 ;
        RECT 66.040 184.030 66.300 184.350 ;
        RECT 63.740 181.310 64.000 181.400 ;
        RECT 64.260 179.590 64.400 181.400 ;
        RECT 64.660 181.310 64.920 181.455 ;
        RECT 65.580 181.310 65.840 181.630 ;
        RECT 64.660 180.630 64.920 180.950 ;
        RECT 65.120 180.630 65.380 180.950 ;
        RECT 64.200 179.270 64.460 179.590 ;
        RECT 63.740 178.590 64.000 178.910 ;
        RECT 63.280 178.250 63.540 178.570 ;
        RECT 63.340 176.870 63.480 178.250 ;
        RECT 63.280 176.550 63.540 176.870 ;
        RECT 63.280 175.870 63.540 176.190 ;
        RECT 63.340 174.150 63.480 175.870 ;
        RECT 63.800 175.170 63.940 178.590 ;
        RECT 63.740 174.850 64.000 175.170 ;
        RECT 63.280 173.830 63.540 174.150 ;
        RECT 63.340 173.470 63.480 173.830 ;
        RECT 63.280 173.150 63.540 173.470 ;
        RECT 63.740 173.150 64.000 173.470 ;
        RECT 63.270 172.615 63.550 172.985 ;
        RECT 63.280 172.470 63.540 172.615 ;
        RECT 62.810 168.535 63.090 168.905 ;
        RECT 63.340 168.030 63.480 172.470 ;
        RECT 63.800 170.750 63.940 173.150 ;
        RECT 64.260 173.130 64.400 179.270 ;
        RECT 64.720 176.530 64.860 180.630 ;
        RECT 64.660 176.210 64.920 176.530 ;
        RECT 64.660 175.530 64.920 175.850 ;
        RECT 64.720 175.170 64.860 175.530 ;
        RECT 64.660 174.850 64.920 175.170 ;
        RECT 64.660 173.830 64.920 174.150 ;
        RECT 64.720 173.665 64.860 173.830 ;
        RECT 64.650 173.295 64.930 173.665 ;
        RECT 64.200 172.810 64.460 173.130 ;
        RECT 64.660 172.810 64.920 173.130 ;
        RECT 63.740 170.430 64.000 170.750 ;
        RECT 64.720 170.070 64.860 172.810 ;
        RECT 65.180 170.945 65.320 180.630 ;
        RECT 65.640 178.570 65.780 181.310 ;
        RECT 66.100 179.590 66.240 184.030 ;
        RECT 67.020 180.610 67.160 196.530 ;
        RECT 67.420 193.890 67.680 194.210 ;
        RECT 67.480 192.590 67.620 193.890 ;
        RECT 67.940 193.190 68.080 203.070 ;
        RECT 68.400 194.550 68.540 207.490 ;
        RECT 68.860 196.785 69.000 213.415 ;
        RECT 71.560 210.550 71.820 210.870 ;
        RECT 71.620 209.170 71.760 210.550 ;
        RECT 72.010 209.335 72.290 209.705 ;
        RECT 71.560 208.850 71.820 209.170 ;
        RECT 69.260 208.510 69.520 208.830 ;
        RECT 69.720 208.510 69.980 208.830 ;
        RECT 70.640 208.510 70.900 208.830 ;
        RECT 69.320 204.945 69.460 208.510 ;
        RECT 69.250 204.575 69.530 204.945 ;
        RECT 69.260 203.750 69.520 204.070 ;
        RECT 69.320 203.050 69.460 203.750 ;
        RECT 69.260 202.730 69.520 203.050 ;
        RECT 69.320 198.630 69.460 202.730 ;
        RECT 69.260 198.310 69.520 198.630 ;
        RECT 69.780 197.950 69.920 208.510 ;
        RECT 70.180 205.790 70.440 206.110 ;
        RECT 70.240 204.070 70.380 205.790 ;
        RECT 70.180 203.750 70.440 204.070 ;
        RECT 70.700 203.050 70.840 208.510 ;
        RECT 72.080 205.625 72.220 209.335 ;
        RECT 71.100 205.110 71.360 205.430 ;
        RECT 72.010 205.255 72.290 205.625 ;
        RECT 71.160 203.050 71.300 205.110 ;
        RECT 71.560 204.770 71.820 205.090 ;
        RECT 71.620 204.070 71.760 204.770 ;
        RECT 71.560 203.750 71.820 204.070 ;
        RECT 72.010 203.215 72.290 203.585 ;
        RECT 70.640 202.730 70.900 203.050 ;
        RECT 71.100 202.730 71.360 203.050 ;
        RECT 71.560 202.730 71.820 203.050 ;
        RECT 71.620 199.505 71.760 202.730 ;
        RECT 71.550 199.135 71.830 199.505 ;
        RECT 70.180 198.310 70.440 198.630 ;
        RECT 69.720 197.630 69.980 197.950 ;
        RECT 68.790 196.415 69.070 196.785 ;
        RECT 69.250 195.055 69.530 195.425 ;
        RECT 68.340 194.230 68.600 194.550 ;
        RECT 68.800 193.890 69.060 194.210 ;
        RECT 67.880 192.870 68.140 193.190 ;
        RECT 67.480 192.450 68.080 192.590 ;
        RECT 67.940 192.170 68.080 192.450 ;
        RECT 67.880 191.850 68.140 192.170 ;
        RECT 67.420 184.710 67.680 185.030 ;
        RECT 67.480 183.240 67.620 184.710 ;
        RECT 67.940 184.010 68.080 191.850 ;
        RECT 68.340 189.470 68.600 189.790 ;
        RECT 67.880 183.690 68.140 184.010 ;
        RECT 67.480 183.100 68.080 183.240 ;
        RECT 66.960 180.290 67.220 180.610 ;
        RECT 66.040 179.270 66.300 179.590 ;
        RECT 66.960 178.590 67.220 178.910 ;
        RECT 65.580 178.250 65.840 178.570 ;
        RECT 66.030 178.055 66.310 178.425 ;
        RECT 66.100 177.630 66.240 178.055 ;
        RECT 65.640 177.490 66.240 177.630 ;
        RECT 65.640 175.850 65.780 177.490 ;
        RECT 67.020 175.850 67.160 178.590 ;
        RECT 67.940 176.950 68.080 183.100 ;
        RECT 68.400 182.310 68.540 189.470 ;
        RECT 68.340 181.990 68.600 182.310 ;
        RECT 67.480 176.810 68.080 176.950 ;
        RECT 67.480 176.190 67.620 176.810 ;
        RECT 68.330 176.695 68.610 177.065 ;
        RECT 67.420 175.870 67.680 176.190 ;
        RECT 67.870 176.015 68.150 176.385 ;
        RECT 65.580 175.530 65.840 175.850 ;
        RECT 66.960 175.530 67.220 175.850 ;
        RECT 67.020 175.170 67.160 175.530 ;
        RECT 65.580 174.850 65.840 175.170 ;
        RECT 66.960 174.850 67.220 175.170 ;
        RECT 65.110 170.575 65.390 170.945 ;
        RECT 64.660 169.750 64.920 170.070 ;
        RECT 65.640 169.585 65.780 174.850 ;
        RECT 66.500 172.985 66.760 173.130 ;
        RECT 66.490 172.615 66.770 172.985 ;
        RECT 66.960 172.810 67.220 173.130 ;
        RECT 67.020 172.450 67.160 172.810 ;
        RECT 66.960 172.130 67.220 172.450 ;
        RECT 66.950 171.255 67.230 171.625 ;
        RECT 67.020 170.070 67.160 171.255 ;
        RECT 67.480 170.150 67.620 175.870 ;
        RECT 67.940 173.130 68.080 176.015 ;
        RECT 67.880 172.810 68.140 173.130 ;
        RECT 67.870 171.935 68.150 172.305 ;
        RECT 67.940 170.750 68.080 171.935 ;
        RECT 68.400 171.430 68.540 176.695 ;
        RECT 68.340 171.110 68.600 171.430 ;
        RECT 68.860 171.090 69.000 193.890 ;
        RECT 69.320 181.825 69.460 195.055 ;
        RECT 70.240 192.170 70.380 198.310 ;
        RECT 72.080 198.290 72.220 203.215 ;
        RECT 72.020 197.970 72.280 198.290 ;
        RECT 70.640 197.630 70.900 197.950 ;
        RECT 70.700 195.230 70.840 197.630 ;
        RECT 70.640 194.910 70.900 195.230 ;
        RECT 72.020 194.910 72.280 195.230 ;
        RECT 71.560 194.570 71.820 194.890 ;
        RECT 71.100 192.190 71.360 192.510 ;
        RECT 70.180 191.850 70.440 192.170 ;
        RECT 70.170 190.295 70.450 190.665 ;
        RECT 69.720 188.450 69.980 188.770 ;
        RECT 69.250 181.455 69.530 181.825 ;
        RECT 69.260 180.630 69.520 180.950 ;
        RECT 69.320 178.570 69.460 180.630 ;
        RECT 69.780 178.570 69.920 188.450 ;
        RECT 69.260 178.250 69.520 178.570 ;
        RECT 69.720 178.250 69.980 178.570 ;
        RECT 69.260 177.570 69.520 177.890 ;
        RECT 69.320 176.530 69.460 177.570 ;
        RECT 69.260 176.210 69.520 176.530 ;
        RECT 68.800 170.770 69.060 171.090 ;
        RECT 67.880 170.430 68.140 170.750 ;
        RECT 69.320 170.320 69.460 176.210 ;
        RECT 69.710 176.015 69.990 176.385 ;
        RECT 69.780 173.470 69.920 176.015 ;
        RECT 70.240 174.150 70.380 190.295 ;
        RECT 71.160 188.770 71.300 192.190 ;
        RECT 71.620 190.470 71.760 194.570 ;
        RECT 71.560 190.150 71.820 190.470 ;
        RECT 71.620 189.450 71.760 190.150 ;
        RECT 71.560 189.130 71.820 189.450 ;
        RECT 71.100 188.450 71.360 188.770 ;
        RECT 70.640 183.010 70.900 183.330 ;
        RECT 70.700 177.890 70.840 183.010 ;
        RECT 71.160 178.570 71.300 188.450 ;
        RECT 71.560 187.430 71.820 187.750 ;
        RECT 71.620 179.590 71.760 187.430 ;
        RECT 71.560 179.270 71.820 179.590 ;
        RECT 71.550 178.735 71.830 179.105 ;
        RECT 71.100 178.250 71.360 178.570 ;
        RECT 70.640 177.570 70.900 177.890 ;
        RECT 70.180 173.830 70.440 174.150 ;
        RECT 69.720 173.150 69.980 173.470 ;
        RECT 70.700 172.870 70.840 177.570 ;
        RECT 71.100 176.780 71.360 176.870 ;
        RECT 71.620 176.780 71.760 178.735 ;
        RECT 71.100 176.640 71.760 176.780 ;
        RECT 71.100 176.550 71.360 176.640 ;
        RECT 71.100 175.870 71.360 176.190 ;
        RECT 71.160 175.170 71.300 175.870 ;
        RECT 71.560 175.190 71.820 175.510 ;
        RECT 71.100 174.850 71.360 175.170 ;
        RECT 69.780 172.730 70.840 172.870 ;
        RECT 69.780 170.750 69.920 172.730 ;
        RECT 70.180 172.305 70.440 172.450 ;
        RECT 70.170 171.935 70.450 172.305 ;
        RECT 69.720 170.430 69.980 170.750 ;
        RECT 68.400 170.180 69.460 170.320 ;
        RECT 66.040 169.750 66.300 170.070 ;
        RECT 66.960 169.750 67.220 170.070 ;
        RECT 67.480 170.010 68.080 170.150 ;
        RECT 65.570 169.215 65.850 169.585 ;
        RECT 65.120 168.390 65.380 168.710 ;
        RECT 61.900 167.710 62.160 168.030 ;
        RECT 63.280 167.710 63.540 168.030 ;
        RECT 61.960 156.810 62.100 167.710 ;
        RECT 65.180 167.690 65.320 168.390 ;
        RECT 65.120 167.370 65.380 167.690 ;
        RECT 65.580 167.370 65.840 167.690 ;
        RECT 66.100 167.600 66.240 169.750 ;
        RECT 66.960 168.225 67.220 168.370 ;
        RECT 66.950 167.855 67.230 168.225 ;
        RECT 67.420 167.600 67.680 167.690 ;
        RECT 66.100 167.460 67.680 167.600 ;
        RECT 65.640 164.630 65.780 167.370 ;
        RECT 65.580 164.310 65.840 164.630 ;
        RECT 66.100 162.590 66.240 167.460 ;
        RECT 67.420 167.370 67.680 167.460 ;
        RECT 66.960 166.690 67.220 167.010 ;
        RECT 67.020 165.650 67.160 166.690 ;
        RECT 66.960 165.330 67.220 165.650 ;
        RECT 67.940 165.390 68.080 170.010 ;
        RECT 68.400 165.990 68.540 170.180 ;
        RECT 69.250 169.215 69.530 169.585 ;
        RECT 68.800 167.370 69.060 167.690 ;
        RECT 68.340 165.670 68.600 165.990 ;
        RECT 66.040 162.270 66.300 162.590 ;
        RECT 63.280 161.250 63.540 161.570 ;
        RECT 63.740 161.250 64.000 161.570 ;
        RECT 63.340 160.550 63.480 161.250 ;
        RECT 63.280 160.230 63.540 160.550 ;
        RECT 63.340 159.870 63.480 160.230 ;
        RECT 63.280 159.550 63.540 159.870 ;
        RECT 62.360 159.210 62.620 159.530 ;
        RECT 62.420 156.810 62.560 159.210 ;
        RECT 63.340 156.810 63.480 159.550 ;
        RECT 63.800 157.150 63.940 161.250 ;
        RECT 64.660 159.890 64.920 160.210 ;
        RECT 63.740 156.830 64.000 157.150 ;
        RECT 61.900 156.490 62.160 156.810 ;
        RECT 62.360 156.490 62.620 156.810 ;
        RECT 63.280 156.490 63.540 156.810 ;
        RECT 63.340 151.370 63.480 156.490 ;
        RECT 64.720 156.470 64.860 159.890 ;
        RECT 65.120 159.210 65.380 159.530 ;
        RECT 65.180 156.810 65.320 159.210 ;
        RECT 67.020 157.830 67.160 165.330 ;
        RECT 67.940 165.250 68.540 165.390 ;
        RECT 67.880 164.650 68.140 164.970 ;
        RECT 67.940 160.550 68.080 164.650 ;
        RECT 67.880 160.230 68.140 160.550 ;
        RECT 65.580 157.510 65.840 157.830 ;
        RECT 66.960 157.510 67.220 157.830 ;
        RECT 65.120 156.490 65.380 156.810 ;
        RECT 64.660 156.150 64.920 156.470 ;
        RECT 65.120 155.810 65.380 156.130 ;
        RECT 63.280 151.050 63.540 151.370 ;
        RECT 61.900 148.670 62.160 148.990 ;
        RECT 61.960 146.950 62.100 148.670 ;
        RECT 63.340 146.950 63.480 151.050 ;
        RECT 64.660 150.940 64.920 151.030 ;
        RECT 65.180 150.940 65.320 155.810 ;
        RECT 65.640 152.050 65.780 157.510 ;
        RECT 66.040 156.830 66.300 157.150 ;
        RECT 66.100 152.390 66.240 156.830 ;
        RECT 68.400 153.750 68.540 165.250 ;
        RECT 68.860 158.850 69.000 167.370 ;
        RECT 68.800 158.530 69.060 158.850 ;
        RECT 68.340 153.430 68.600 153.750 ;
        RECT 66.040 152.070 66.300 152.390 ;
        RECT 65.580 151.730 65.840 152.050 ;
        RECT 64.660 150.800 65.320 150.940 ;
        RECT 64.660 150.710 64.920 150.800 ;
        RECT 64.720 148.310 64.860 150.710 ;
        RECT 65.640 149.670 65.780 151.730 ;
        RECT 65.580 149.350 65.840 149.670 ;
        RECT 64.660 147.990 64.920 148.310 ;
        RECT 61.900 146.630 62.160 146.950 ;
        RECT 63.280 146.630 63.540 146.950 ;
        RECT 66.100 145.930 66.240 152.070 ;
        RECT 69.320 151.370 69.460 169.215 ;
        RECT 69.720 167.420 69.980 167.740 ;
        RECT 69.780 164.630 69.920 167.420 ;
        RECT 70.240 165.650 70.380 171.935 ;
        RECT 70.640 170.430 70.900 170.750 ;
        RECT 70.700 168.030 70.840 170.430 ;
        RECT 70.640 167.710 70.900 168.030 ;
        RECT 71.160 167.350 71.300 174.850 ;
        RECT 71.620 173.130 71.760 175.190 ;
        RECT 72.080 173.810 72.220 194.910 ;
        RECT 72.020 173.490 72.280 173.810 ;
        RECT 71.560 172.810 71.820 173.130 ;
        RECT 72.020 170.945 72.280 171.090 ;
        RECT 72.010 170.575 72.290 170.945 ;
        RECT 72.020 167.600 72.280 167.690 ;
        RECT 71.620 167.460 72.280 167.600 ;
        RECT 71.100 167.030 71.360 167.350 ;
        RECT 70.180 165.330 70.440 165.650 ;
        RECT 71.090 165.135 71.370 165.505 ;
        RECT 69.720 164.310 69.980 164.630 ;
        RECT 70.640 159.550 70.900 159.870 ;
        RECT 70.700 157.490 70.840 159.550 ;
        RECT 70.640 157.170 70.900 157.490 ;
        RECT 70.180 156.490 70.440 156.810 ;
        RECT 69.720 154.110 69.980 154.430 ;
        RECT 69.780 151.370 69.920 154.110 ;
        RECT 70.240 152.390 70.380 156.490 ;
        RECT 70.700 156.130 70.840 157.170 ;
        RECT 70.640 155.810 70.900 156.130 ;
        RECT 71.160 155.110 71.300 165.135 ;
        RECT 71.620 158.850 71.760 167.460 ;
        RECT 72.020 167.370 72.280 167.460 ;
        RECT 72.020 165.220 72.280 165.310 ;
        RECT 72.540 165.220 72.680 217.610 ;
        RECT 73.850 217.330 74.130 221.330 ;
        RECT 77.070 217.330 77.350 221.330 ;
        RECT 78.520 217.610 80.040 217.750 ;
        RECT 73.920 211.745 74.060 217.330 ;
        RECT 77.140 216.505 77.280 217.330 ;
        RECT 77.070 216.135 77.350 216.505 ;
        RECT 73.850 211.375 74.130 211.745 ;
        RECT 73.400 208.850 73.660 209.170 ;
        RECT 72.940 206.470 73.200 206.790 ;
        RECT 73.000 202.225 73.140 206.470 ;
        RECT 72.930 201.855 73.210 202.225 ;
        RECT 72.940 200.350 73.200 200.670 ;
        RECT 73.000 194.890 73.140 200.350 ;
        RECT 72.940 194.570 73.200 194.890 ;
        RECT 73.460 191.490 73.600 208.850 ;
        RECT 75.240 208.510 75.500 208.830 ;
        RECT 75.300 208.150 75.440 208.510 ;
        RECT 75.240 207.830 75.500 208.150 ;
        RECT 73.860 203.070 74.120 203.390 ;
        RECT 74.310 203.215 74.590 203.585 ;
        RECT 74.320 203.070 74.580 203.215 ;
        RECT 73.920 202.370 74.060 203.070 ;
        RECT 73.860 202.050 74.120 202.370 ;
        RECT 74.780 191.850 75.040 192.170 ;
        RECT 73.400 191.170 73.660 191.490 ;
        RECT 74.320 191.170 74.580 191.490 ;
        RECT 73.460 186.730 73.600 191.170 ;
        RECT 74.380 187.070 74.520 191.170 ;
        RECT 74.320 186.750 74.580 187.070 ;
        RECT 73.400 186.410 73.660 186.730 ;
        RECT 74.840 186.470 74.980 191.850 ;
        RECT 75.300 187.410 75.440 207.830 ;
        RECT 77.540 206.130 77.800 206.450 ;
        RECT 77.600 205.770 77.740 206.130 ;
        RECT 75.700 205.450 75.960 205.770 ;
        RECT 77.540 205.450 77.800 205.770 ;
        RECT 75.760 201.545 75.900 205.450 ;
        RECT 76.620 202.050 76.880 202.370 ;
        RECT 75.690 201.175 75.970 201.545 ;
        RECT 76.160 201.030 76.420 201.350 ;
        RECT 75.690 193.015 75.970 193.385 ;
        RECT 75.240 187.090 75.500 187.410 ;
        RECT 72.940 184.710 73.200 185.030 ;
        RECT 73.000 179.250 73.140 184.710 ;
        RECT 72.940 178.930 73.200 179.250 ;
        RECT 72.940 177.910 73.200 178.230 ;
        RECT 72.020 165.080 72.680 165.220 ;
        RECT 72.020 164.990 72.280 165.080 ;
        RECT 72.010 164.455 72.290 164.825 ;
        RECT 72.020 164.310 72.280 164.455 ;
        RECT 72.540 163.270 72.680 165.080 ;
        RECT 73.000 164.630 73.140 177.910 ;
        RECT 73.460 175.510 73.600 186.410 ;
        RECT 74.840 186.330 75.440 186.470 ;
        RECT 74.780 185.730 75.040 186.050 ;
        RECT 74.840 184.010 74.980 185.730 ;
        RECT 75.300 184.690 75.440 186.330 ;
        RECT 75.240 184.370 75.500 184.690 ;
        RECT 74.780 183.690 75.040 184.010 ;
        RECT 73.860 181.990 74.120 182.310 ;
        RECT 73.920 178.570 74.060 181.990 ;
        RECT 74.780 181.650 75.040 181.970 ;
        RECT 73.860 178.250 74.120 178.570 ;
        RECT 74.320 178.250 74.580 178.570 ;
        RECT 73.400 175.190 73.660 175.510 ;
        RECT 74.380 174.910 74.520 178.250 ;
        RECT 74.840 175.850 74.980 181.650 ;
        RECT 75.240 175.870 75.500 176.190 ;
        RECT 74.780 175.530 75.040 175.850 ;
        RECT 73.460 174.770 74.520 174.910 ;
        RECT 73.460 174.150 73.600 174.770 ;
        RECT 74.840 174.150 74.980 175.530 ;
        RECT 73.400 173.830 73.660 174.150 ;
        RECT 74.320 173.830 74.580 174.150 ;
        RECT 74.780 173.830 75.040 174.150 ;
        RECT 73.400 170.430 73.660 170.750 ;
        RECT 73.860 170.430 74.120 170.750 ;
        RECT 73.460 168.370 73.600 170.430 ;
        RECT 73.400 168.050 73.660 168.370 ;
        RECT 73.920 167.690 74.060 170.430 ;
        RECT 73.860 167.370 74.120 167.690 ;
        RECT 73.400 165.560 73.660 165.650 ;
        RECT 73.920 165.560 74.060 167.370 ;
        RECT 73.400 165.420 74.060 165.560 ;
        RECT 73.400 165.330 73.660 165.420 ;
        RECT 72.940 164.310 73.200 164.630 ;
        RECT 72.480 162.950 72.740 163.270 ;
        RECT 72.940 162.950 73.200 163.270 ;
        RECT 72.020 161.590 72.280 161.910 ;
        RECT 72.080 160.210 72.220 161.590 ;
        RECT 72.020 159.890 72.280 160.210 ;
        RECT 72.480 159.550 72.740 159.870 ;
        RECT 72.020 158.870 72.280 159.190 ;
        RECT 71.560 158.530 71.820 158.850 ;
        RECT 71.100 154.790 71.360 155.110 ;
        RECT 71.100 154.110 71.360 154.430 ;
        RECT 70.180 152.070 70.440 152.390 ;
        RECT 71.160 151.370 71.300 154.110 ;
        RECT 71.620 153.750 71.760 158.530 ;
        RECT 72.080 157.830 72.220 158.870 ;
        RECT 72.540 158.760 72.680 159.550 ;
        RECT 73.000 158.850 73.140 162.950 ;
        RECT 73.400 159.890 73.660 160.210 ;
        RECT 72.940 158.760 73.200 158.850 ;
        RECT 72.540 158.620 73.200 158.760 ;
        RECT 72.020 157.510 72.280 157.830 ;
        RECT 72.540 155.110 72.680 158.620 ;
        RECT 72.940 158.530 73.200 158.620 ;
        RECT 73.460 156.810 73.600 159.890 ;
        RECT 73.920 157.830 74.060 165.420 ;
        RECT 74.380 165.310 74.520 173.830 ;
        RECT 74.780 173.150 75.040 173.470 ;
        RECT 74.840 167.690 74.980 173.150 ;
        RECT 74.780 167.370 75.040 167.690 ;
        RECT 74.320 164.990 74.580 165.310 ;
        RECT 74.840 164.630 74.980 167.370 ;
        RECT 75.300 165.505 75.440 175.870 ;
        RECT 75.760 170.070 75.900 193.015 ;
        RECT 76.220 187.070 76.360 201.030 ;
        RECT 76.680 192.510 76.820 202.050 ;
        RECT 76.620 192.190 76.880 192.510 ;
        RECT 77.540 192.190 77.800 192.510 ;
        RECT 76.610 190.975 76.890 191.345 ;
        RECT 76.160 186.750 76.420 187.070 ;
        RECT 76.680 183.865 76.820 190.975 ;
        RECT 77.600 189.790 77.740 192.190 ;
        RECT 77.540 189.470 77.800 189.790 ;
        RECT 77.540 188.790 77.800 189.110 ;
        RECT 77.080 187.430 77.340 187.750 ;
        RECT 77.140 185.225 77.280 187.430 ;
        RECT 77.070 184.855 77.350 185.225 ;
        RECT 77.600 184.350 77.740 188.790 ;
        RECT 78.000 186.750 78.260 187.070 ;
        RECT 77.540 184.030 77.800 184.350 ;
        RECT 76.610 183.495 76.890 183.865 ;
        RECT 76.160 183.010 76.420 183.330 ;
        RECT 76.220 181.630 76.360 183.010 ;
        RECT 76.160 181.310 76.420 181.630 ;
        RECT 77.080 181.310 77.340 181.630 ;
        RECT 77.140 176.190 77.280 181.310 ;
        RECT 77.600 179.250 77.740 184.030 ;
        RECT 77.540 178.930 77.800 179.250 ;
        RECT 78.060 178.570 78.200 186.750 ;
        RECT 78.000 178.250 78.260 178.570 ;
        RECT 78.520 177.630 78.660 217.610 ;
        RECT 79.900 217.070 80.040 217.610 ;
        RECT 80.290 217.330 80.570 221.330 ;
        RECT 83.510 217.330 83.790 221.330 ;
        RECT 86.730 217.330 87.010 221.330 ;
        RECT 89.950 217.330 90.230 221.330 ;
        RECT 93.170 217.330 93.450 221.330 ;
        RECT 80.360 217.070 80.500 217.330 ;
        RECT 79.900 216.930 80.500 217.070 ;
        RECT 79.830 214.095 80.110 214.465 ;
        RECT 79.370 207.295 79.650 207.665 ;
        RECT 79.440 206.110 79.580 207.295 ;
        RECT 79.380 205.790 79.640 206.110 ;
        RECT 79.900 201.010 80.040 214.095 ;
        RECT 80.300 212.930 80.560 213.250 ;
        RECT 80.360 202.280 80.500 212.930 ;
        RECT 81.680 212.590 81.940 212.910 ;
        RECT 81.740 209.510 81.880 212.590 ;
        RECT 83.580 212.425 83.720 217.330 ;
        RECT 83.510 212.055 83.790 212.425 ;
        RECT 82.600 211.230 82.860 211.550 ;
        RECT 81.680 209.190 81.940 209.510 ;
        RECT 81.220 208.510 81.480 208.830 ;
        RECT 82.130 208.655 82.410 209.025 ;
        RECT 80.760 208.170 81.020 208.490 ;
        RECT 80.820 203.050 80.960 208.170 ;
        RECT 81.280 205.625 81.420 208.510 ;
        RECT 82.200 208.150 82.340 208.655 ;
        RECT 82.140 207.830 82.400 208.150 ;
        RECT 82.200 205.770 82.340 207.830 ;
        RECT 81.210 205.255 81.490 205.625 ;
        RECT 82.140 205.450 82.400 205.770 ;
        RECT 81.680 204.770 81.940 205.090 ;
        RECT 80.760 202.730 81.020 203.050 ;
        RECT 80.360 202.140 81.420 202.280 ;
        RECT 79.840 200.690 80.100 201.010 ;
        RECT 81.280 199.390 81.420 202.140 ;
        RECT 81.740 200.330 81.880 204.770 ;
        RECT 82.660 200.330 82.800 211.230 ;
        RECT 83.060 208.345 83.320 208.490 ;
        RECT 83.050 207.975 83.330 208.345 ;
        RECT 86.270 207.975 86.550 208.345 ;
        RECT 84.440 207.490 84.700 207.810 ;
        RECT 85.360 207.490 85.620 207.810 ;
        RECT 83.980 203.070 84.240 203.390 ;
        RECT 84.500 203.300 84.640 207.490 ;
        RECT 85.420 206.110 85.560 207.490 ;
        RECT 85.360 205.790 85.620 206.110 ;
        RECT 84.900 205.450 85.160 205.770 ;
        RECT 84.960 204.945 85.100 205.450 ;
        RECT 85.820 205.110 86.080 205.430 ;
        RECT 84.890 204.575 85.170 204.945 ;
        RECT 85.880 204.150 86.020 205.110 ;
        RECT 86.340 205.090 86.480 207.975 ;
        RECT 86.280 204.770 86.540 205.090 ;
        RECT 85.880 204.070 86.480 204.150 ;
        RECT 85.880 204.010 86.540 204.070 ;
        RECT 86.280 203.750 86.540 204.010 ;
        RECT 85.820 203.300 86.080 203.390 ;
        RECT 84.500 203.160 86.080 203.300 ;
        RECT 85.820 203.070 86.080 203.160 ;
        RECT 81.680 200.010 81.940 200.330 ;
        RECT 82.600 200.010 82.860 200.330 ;
        RECT 83.520 200.010 83.780 200.330 ;
        RECT 80.360 199.250 81.420 199.390 ;
        RECT 78.920 197.290 79.180 197.610 ;
        RECT 78.980 195.230 79.120 197.290 ;
        RECT 80.360 196.930 80.500 199.250 ;
        RECT 80.750 198.455 81.030 198.825 ;
        RECT 80.760 198.310 81.020 198.455 ;
        RECT 80.820 197.950 80.960 198.310 ;
        RECT 81.280 197.950 81.420 199.250 ;
        RECT 80.760 197.630 81.020 197.950 ;
        RECT 81.220 197.630 81.480 197.950 ;
        RECT 81.670 197.775 81.950 198.145 ;
        RECT 81.220 196.950 81.480 197.270 ;
        RECT 80.300 196.610 80.560 196.930 ;
        RECT 80.760 195.590 81.020 195.910 ;
        RECT 78.920 194.910 79.180 195.230 ;
        RECT 79.840 191.510 80.100 191.830 ;
        RECT 79.900 190.430 80.040 191.510 ;
        RECT 79.440 190.290 80.040 190.430 ;
        RECT 78.920 189.810 79.180 190.130 ;
        RECT 78.060 177.490 78.660 177.630 ;
        RECT 77.080 175.870 77.340 176.190 ;
        RECT 76.160 175.530 76.420 175.850 ;
        RECT 78.060 175.705 78.200 177.490 ;
        RECT 78.460 176.550 78.720 176.870 ;
        RECT 76.220 175.170 76.360 175.530 ;
        RECT 77.990 175.335 78.270 175.705 ;
        RECT 76.160 174.850 76.420 175.170 ;
        RECT 77.540 173.830 77.800 174.150 ;
        RECT 76.160 172.810 76.420 173.130 ;
        RECT 76.620 172.810 76.880 173.130 ;
        RECT 76.220 170.070 76.360 172.810 ;
        RECT 76.680 171.510 76.820 172.810 ;
        RECT 76.680 171.370 77.280 171.510 ;
        RECT 76.620 170.430 76.880 170.750 ;
        RECT 75.700 169.750 75.960 170.070 ;
        RECT 76.160 169.750 76.420 170.070 ;
        RECT 76.680 169.730 76.820 170.430 ;
        RECT 77.140 170.265 77.280 171.370 ;
        RECT 77.070 169.895 77.350 170.265 ;
        RECT 77.600 169.730 77.740 173.830 ;
        RECT 78.520 173.665 78.660 176.550 ;
        RECT 78.980 175.025 79.120 189.810 ;
        RECT 79.440 183.750 79.580 190.290 ;
        RECT 79.840 184.430 80.100 184.690 ;
        RECT 79.840 184.370 80.500 184.430 ;
        RECT 79.900 184.290 80.500 184.370 ;
        RECT 80.360 184.010 80.500 184.290 ;
        RECT 79.840 183.750 80.100 184.010 ;
        RECT 79.440 183.690 80.100 183.750 ;
        RECT 80.300 183.690 80.560 184.010 ;
        RECT 79.440 183.610 80.040 183.690 ;
        RECT 79.440 175.850 79.580 183.610 ;
        RECT 80.300 183.010 80.560 183.330 ;
        RECT 80.360 180.610 80.500 183.010 ;
        RECT 80.300 180.290 80.560 180.610 ;
        RECT 79.380 175.530 79.640 175.850 ;
        RECT 78.910 174.655 79.190 175.025 ;
        RECT 78.450 173.295 78.730 173.665 ;
        RECT 78.920 173.490 79.180 173.810 ;
        RECT 79.380 173.490 79.640 173.810 ;
        RECT 78.000 172.810 78.260 173.130 ;
        RECT 78.060 171.090 78.200 172.810 ;
        RECT 78.000 170.770 78.260 171.090 ;
        RECT 78.460 170.430 78.720 170.750 ;
        RECT 78.000 169.750 78.260 170.070 ;
        RECT 76.680 169.590 77.740 169.730 ;
        RECT 76.610 168.535 76.890 168.905 ;
        RECT 77.600 168.790 77.740 169.590 ;
        RECT 78.060 169.585 78.200 169.750 ;
        RECT 77.990 169.215 78.270 169.585 ;
        RECT 77.600 168.650 78.200 168.790 ;
        RECT 76.680 167.690 76.820 168.535 ;
        RECT 77.540 168.050 77.800 168.370 ;
        RECT 76.620 167.370 76.880 167.690 ;
        RECT 75.700 166.690 75.960 167.010 ;
        RECT 75.230 165.135 75.510 165.505 ;
        RECT 75.240 164.990 75.500 165.135 ;
        RECT 74.780 164.310 75.040 164.630 ;
        RECT 74.840 163.270 74.980 164.310 ;
        RECT 75.240 163.970 75.500 164.290 ;
        RECT 74.780 162.950 75.040 163.270 ;
        RECT 74.780 161.930 75.040 162.250 ;
        RECT 74.840 159.190 74.980 161.930 ;
        RECT 75.300 160.550 75.440 163.970 ;
        RECT 75.760 162.930 75.900 166.690 ;
        RECT 76.160 164.990 76.420 165.310 ;
        RECT 76.620 164.990 76.880 165.310 ;
        RECT 76.220 163.270 76.360 164.990 ;
        RECT 76.160 162.950 76.420 163.270 ;
        RECT 75.700 162.610 75.960 162.930 ;
        RECT 76.150 162.415 76.430 162.785 ;
        RECT 76.680 162.590 76.820 164.990 ;
        RECT 77.600 164.290 77.740 168.050 ;
        RECT 78.060 167.350 78.200 168.650 ;
        RECT 78.520 168.370 78.660 170.430 ;
        RECT 78.460 168.050 78.720 168.370 ;
        RECT 78.000 167.030 78.260 167.350 ;
        RECT 78.060 165.650 78.200 167.030 ;
        RECT 78.000 165.330 78.260 165.650 ;
        RECT 78.460 164.990 78.720 165.310 ;
        RECT 78.520 164.630 78.660 164.990 ;
        RECT 78.460 164.310 78.720 164.630 ;
        RECT 77.540 163.970 77.800 164.290 ;
        RECT 77.540 162.950 77.800 163.270 ;
        RECT 76.220 162.250 76.360 162.415 ;
        RECT 76.620 162.270 76.880 162.590 ;
        RECT 76.160 161.930 76.420 162.250 ;
        RECT 77.070 161.735 77.350 162.105 ;
        RECT 77.140 161.570 77.280 161.735 ;
        RECT 77.080 161.250 77.340 161.570 ;
        RECT 77.600 160.550 77.740 162.950 ;
        RECT 78.980 162.250 79.120 173.490 ;
        RECT 79.440 170.945 79.580 173.490 ;
        RECT 79.370 170.575 79.650 170.945 ;
        RECT 79.370 167.855 79.650 168.225 ;
        RECT 79.440 164.630 79.580 167.855 ;
        RECT 80.360 167.350 80.500 180.290 ;
        RECT 80.820 179.250 80.960 195.590 ;
        RECT 81.280 190.665 81.420 196.950 ;
        RECT 81.740 191.830 81.880 197.775 ;
        RECT 82.600 194.745 82.860 194.890 ;
        RECT 82.140 194.230 82.400 194.550 ;
        RECT 82.590 194.375 82.870 194.745 ;
        RECT 83.060 194.570 83.320 194.890 ;
        RECT 82.200 191.830 82.340 194.230 ;
        RECT 82.600 193.890 82.860 194.210 ;
        RECT 83.120 194.065 83.260 194.570 ;
        RECT 81.680 191.510 81.940 191.830 ;
        RECT 82.140 191.510 82.400 191.830 ;
        RECT 81.210 190.295 81.490 190.665 ;
        RECT 81.220 189.470 81.480 189.790 ;
        RECT 81.280 183.330 81.420 189.470 ;
        RECT 81.220 183.010 81.480 183.330 ;
        RECT 81.220 180.630 81.480 180.950 ;
        RECT 80.760 178.930 81.020 179.250 ;
        RECT 81.280 178.570 81.420 180.630 ;
        RECT 81.220 178.250 81.480 178.570 ;
        RECT 81.220 176.550 81.480 176.870 ;
        RECT 81.280 175.760 81.420 176.550 ;
        RECT 81.740 176.530 81.880 191.510 ;
        RECT 82.660 189.450 82.800 193.890 ;
        RECT 83.050 193.695 83.330 194.065 ;
        RECT 83.580 192.025 83.720 200.010 ;
        RECT 83.510 191.655 83.790 192.025 ;
        RECT 83.520 190.150 83.780 190.470 ;
        RECT 83.060 189.470 83.320 189.790 ;
        RECT 82.600 189.130 82.860 189.450 ;
        RECT 82.140 188.790 82.400 189.110 ;
        RECT 81.680 176.210 81.940 176.530 ;
        RECT 81.280 175.620 81.880 175.760 ;
        RECT 80.300 167.030 80.560 167.350 ;
        RECT 80.300 164.650 80.560 164.970 ;
        RECT 80.760 164.650 81.020 164.970 ;
        RECT 79.380 164.310 79.640 164.630 ;
        RECT 80.360 162.590 80.500 164.650 ;
        RECT 80.300 162.270 80.560 162.590 ;
        RECT 78.920 161.930 79.180 162.250 ;
        RECT 75.240 160.230 75.500 160.550 ;
        RECT 77.540 160.230 77.800 160.550 ;
        RECT 75.700 159.890 75.960 160.210 ;
        RECT 76.620 159.890 76.880 160.210 ;
        RECT 74.780 158.870 75.040 159.190 ;
        RECT 73.860 157.510 74.120 157.830 ;
        RECT 73.400 156.490 73.660 156.810 ;
        RECT 72.480 154.790 72.740 155.110 ;
        RECT 72.020 153.770 72.280 154.090 ;
        RECT 71.560 153.430 71.820 153.750 ;
        RECT 72.080 151.370 72.220 153.770 ;
        RECT 75.760 152.050 75.900 159.890 ;
        RECT 76.680 156.810 76.820 159.890 ;
        RECT 78.980 157.830 79.120 161.930 ;
        RECT 80.820 161.910 80.960 164.650 ;
        RECT 81.740 164.290 81.880 175.620 ;
        RECT 82.200 174.150 82.340 188.790 ;
        RECT 83.120 188.625 83.260 189.470 ;
        RECT 83.050 188.255 83.330 188.625 ;
        RECT 82.590 186.215 82.870 186.585 ;
        RECT 82.140 173.830 82.400 174.150 ;
        RECT 82.130 173.295 82.410 173.665 ;
        RECT 82.200 165.560 82.340 173.295 ;
        RECT 82.660 171.430 82.800 186.215 ;
        RECT 83.060 183.690 83.320 184.010 ;
        RECT 83.120 175.170 83.260 183.690 ;
        RECT 83.060 174.850 83.320 175.170 ;
        RECT 83.050 173.975 83.330 174.345 ;
        RECT 82.600 171.110 82.860 171.430 ;
        RECT 82.200 165.420 82.800 165.560 ;
        RECT 82.140 164.650 82.400 164.970 ;
        RECT 81.680 163.970 81.940 164.290 ;
        RECT 80.760 161.590 81.020 161.910 ;
        RECT 80.290 159.015 80.570 159.385 ;
        RECT 80.360 157.830 80.500 159.015 ;
        RECT 78.920 157.510 79.180 157.830 ;
        RECT 80.300 157.510 80.560 157.830 ;
        RECT 76.620 156.490 76.880 156.810 ;
        RECT 80.820 155.870 80.960 161.590 ;
        RECT 81.220 161.250 81.480 161.570 ;
        RECT 81.280 156.810 81.420 161.250 ;
        RECT 81.220 156.490 81.480 156.810 ;
        RECT 82.200 156.470 82.340 164.650 ;
        RECT 82.660 162.250 82.800 165.420 ;
        RECT 83.120 164.970 83.260 173.975 ;
        RECT 83.580 171.430 83.720 190.150 ;
        RECT 84.040 189.870 84.180 203.070 ;
        RECT 86.800 202.790 86.940 217.330 ;
        RECT 87.650 210.015 87.930 210.385 ;
        RECT 87.720 208.830 87.860 210.015 ;
        RECT 87.660 208.510 87.920 208.830 ;
        RECT 87.200 208.170 87.460 208.490 ;
        RECT 86.340 202.650 86.940 202.790 ;
        RECT 84.440 199.670 84.700 199.990 ;
        RECT 84.500 199.505 84.640 199.670 ;
        RECT 84.430 199.135 84.710 199.505 ;
        RECT 84.440 198.310 84.700 198.630 ;
        RECT 84.500 197.950 84.640 198.310 ;
        RECT 84.440 197.630 84.700 197.950 ;
        RECT 85.820 197.630 86.080 197.950 ;
        RECT 84.900 195.250 85.160 195.570 ;
        RECT 84.440 191.510 84.700 191.830 ;
        RECT 84.500 190.470 84.640 191.510 ;
        RECT 84.440 190.150 84.700 190.470 ;
        RECT 84.040 189.730 84.640 189.870 ;
        RECT 84.500 186.050 84.640 189.730 ;
        RECT 84.440 185.730 84.700 186.050 ;
        RECT 83.980 183.010 84.240 183.330 ;
        RECT 84.040 179.250 84.180 183.010 ;
        RECT 84.500 181.970 84.640 185.730 ;
        RECT 84.440 181.650 84.700 181.970 ;
        RECT 83.980 178.930 84.240 179.250 ;
        RECT 84.440 178.250 84.700 178.570 ;
        RECT 84.500 176.870 84.640 178.250 ;
        RECT 84.440 176.550 84.700 176.870 ;
        RECT 83.980 175.190 84.240 175.510 ;
        RECT 84.040 174.150 84.180 175.190 ;
        RECT 84.440 174.850 84.700 175.170 ;
        RECT 83.980 173.830 84.240 174.150 ;
        RECT 83.520 171.110 83.780 171.430 ;
        RECT 83.060 164.650 83.320 164.970 ;
        RECT 83.060 163.970 83.320 164.290 ;
        RECT 82.600 161.930 82.860 162.250 ;
        RECT 83.120 159.270 83.260 163.970 ;
        RECT 83.580 160.210 83.720 171.110 ;
        RECT 84.040 167.600 84.180 173.830 ;
        RECT 84.500 173.470 84.640 174.850 ;
        RECT 84.440 173.150 84.700 173.470 ;
        RECT 84.960 168.030 85.100 195.250 ;
        RECT 85.360 194.570 85.620 194.890 ;
        RECT 85.420 190.470 85.560 194.570 ;
        RECT 85.360 190.150 85.620 190.470 ;
        RECT 85.360 188.790 85.620 189.110 ;
        RECT 85.420 187.750 85.560 188.790 ;
        RECT 85.360 187.430 85.620 187.750 ;
        RECT 85.360 186.750 85.620 187.070 ;
        RECT 85.420 185.030 85.560 186.750 ;
        RECT 85.360 184.710 85.620 185.030 ;
        RECT 85.360 183.350 85.620 183.670 ;
        RECT 85.420 179.250 85.560 183.350 ;
        RECT 85.880 181.710 86.020 197.630 ;
        RECT 86.340 187.410 86.480 202.650 ;
        RECT 87.260 195.910 87.400 208.170 ;
        RECT 87.650 205.935 87.930 206.305 ;
        RECT 87.720 205.770 87.860 205.935 ;
        RECT 87.660 205.450 87.920 205.770 ;
        RECT 89.500 198.310 89.760 198.630 ;
        RECT 88.120 197.630 88.380 197.950 ;
        RECT 87.200 195.590 87.460 195.910 ;
        RECT 86.740 194.570 87.000 194.890 ;
        RECT 86.800 193.190 86.940 194.570 ;
        RECT 87.200 193.890 87.460 194.210 ;
        RECT 86.740 192.870 87.000 193.190 ;
        RECT 87.260 192.850 87.400 193.890 ;
        RECT 87.200 192.530 87.460 192.850 ;
        RECT 87.660 192.190 87.920 192.510 ;
        RECT 87.200 189.130 87.460 189.450 ;
        RECT 86.740 188.450 87.000 188.770 ;
        RECT 86.280 187.090 86.540 187.410 ;
        RECT 85.880 181.570 86.480 181.710 ;
        RECT 86.340 181.290 86.480 181.570 ;
        RECT 86.280 180.970 86.540 181.290 ;
        RECT 85.360 178.930 85.620 179.250 ;
        RECT 85.820 173.830 86.080 174.150 ;
        RECT 85.880 173.470 86.020 173.830 ;
        RECT 85.820 173.150 86.080 173.470 ;
        RECT 85.360 172.810 85.620 173.130 ;
        RECT 85.420 171.625 85.560 172.810 ;
        RECT 85.350 171.255 85.630 171.625 ;
        RECT 84.900 167.710 85.160 168.030 ;
        RECT 84.440 167.600 84.700 167.690 ;
        RECT 84.040 167.460 84.700 167.600 ;
        RECT 84.440 167.370 84.700 167.460 ;
        RECT 83.970 165.815 84.250 166.185 ;
        RECT 83.980 165.670 84.240 165.815 ;
        RECT 84.440 164.650 84.700 164.970 ;
        RECT 84.500 164.290 84.640 164.650 ;
        RECT 83.980 163.970 84.240 164.290 ;
        RECT 84.440 163.970 84.700 164.290 ;
        RECT 83.520 159.890 83.780 160.210 ;
        RECT 83.120 159.130 83.720 159.270 ;
        RECT 82.140 156.150 82.400 156.470 ;
        RECT 81.220 155.870 81.480 156.130 ;
        RECT 80.820 155.810 81.480 155.870 ;
        RECT 80.820 155.730 81.420 155.810 ;
        RECT 81.280 154.770 81.420 155.730 ;
        RECT 81.220 154.450 81.480 154.770 ;
        RECT 81.680 153.090 81.940 153.410 ;
        RECT 75.700 151.730 75.960 152.050 ;
        RECT 67.880 151.050 68.140 151.370 ;
        RECT 69.260 151.050 69.520 151.370 ;
        RECT 69.720 151.050 69.980 151.370 ;
        RECT 71.100 151.050 71.360 151.370 ;
        RECT 72.020 151.050 72.280 151.370 ;
        RECT 81.740 151.225 81.880 153.090 ;
        RECT 66.960 150.710 67.220 151.030 ;
        RECT 67.020 147.970 67.160 150.710 ;
        RECT 67.940 148.990 68.080 151.050 ;
        RECT 68.340 150.370 68.600 150.690 ;
        RECT 68.400 149.330 68.540 150.370 ;
        RECT 69.320 149.330 69.460 151.050 ;
        RECT 81.670 150.855 81.950 151.225 ;
        RECT 81.680 150.710 81.940 150.855 ;
        RECT 68.340 149.010 68.600 149.330 ;
        RECT 69.260 149.010 69.520 149.330 ;
        RECT 67.880 148.670 68.140 148.990 ;
        RECT 82.200 148.310 82.340 156.150 ;
        RECT 82.600 154.110 82.860 154.430 ;
        RECT 82.660 152.585 82.800 154.110 ;
        RECT 83.580 154.090 83.720 159.130 ;
        RECT 84.040 154.430 84.180 163.970 ;
        RECT 84.430 162.415 84.710 162.785 ;
        RECT 84.500 155.110 84.640 162.415 ;
        RECT 84.960 162.250 85.100 167.710 ;
        RECT 85.420 164.630 85.560 171.255 ;
        RECT 86.340 165.990 86.480 180.970 ;
        RECT 86.800 172.450 86.940 188.450 ;
        RECT 87.260 184.545 87.400 189.130 ;
        RECT 87.190 184.175 87.470 184.545 ;
        RECT 87.200 183.690 87.460 184.010 ;
        RECT 87.260 182.310 87.400 183.690 ;
        RECT 87.200 181.990 87.460 182.310 ;
        RECT 87.720 179.785 87.860 192.190 ;
        RECT 88.180 183.185 88.320 197.630 ;
        RECT 89.030 191.655 89.310 192.025 ;
        RECT 88.580 183.350 88.840 183.670 ;
        RECT 88.110 182.815 88.390 183.185 ;
        RECT 87.650 179.415 87.930 179.785 ;
        RECT 87.200 177.570 87.460 177.890 ;
        RECT 87.260 176.385 87.400 177.570 ;
        RECT 87.190 176.015 87.470 176.385 ;
        RECT 87.190 172.615 87.470 172.985 ;
        RECT 88.640 172.790 88.780 183.350 ;
        RECT 89.100 174.150 89.240 191.655 ;
        RECT 89.560 183.670 89.700 198.310 ;
        RECT 89.500 183.350 89.760 183.670 ;
        RECT 90.020 178.425 90.160 217.330 ;
        RECT 93.240 211.745 93.380 217.330 ;
        RECT 93.170 211.375 93.450 211.745 ;
        RECT 89.950 178.055 90.230 178.425 ;
        RECT 89.040 173.830 89.300 174.150 ;
        RECT 87.260 172.450 87.400 172.615 ;
        RECT 88.580 172.470 88.840 172.790 ;
        RECT 86.740 172.130 87.000 172.450 ;
        RECT 87.200 172.130 87.460 172.450 ;
        RECT 86.280 165.670 86.540 165.990 ;
        RECT 85.360 164.310 85.620 164.630 ;
        RECT 84.900 161.930 85.160 162.250 ;
        RECT 85.360 161.930 85.620 162.250 ;
        RECT 85.420 160.550 85.560 161.930 ;
        RECT 85.360 160.230 85.620 160.550 ;
        RECT 86.340 156.810 86.480 165.670 ;
        RECT 87.660 165.330 87.920 165.650 ;
        RECT 86.740 164.200 87.000 164.290 ;
        RECT 86.740 164.060 87.400 164.200 ;
        RECT 86.740 163.970 87.000 164.060 ;
        RECT 86.740 161.930 87.000 162.250 ;
        RECT 86.800 156.810 86.940 161.930 ;
        RECT 86.280 156.490 86.540 156.810 ;
        RECT 86.740 156.490 87.000 156.810 ;
        RECT 84.900 155.810 85.160 156.130 ;
        RECT 84.440 154.790 84.700 155.110 ;
        RECT 83.980 154.110 84.240 154.430 ;
        RECT 83.520 153.770 83.780 154.090 ;
        RECT 82.590 152.215 82.870 152.585 ;
        RECT 84.960 151.370 85.100 155.810 ;
        RECT 85.810 155.615 86.090 155.985 ;
        RECT 85.880 152.390 86.020 155.615 ;
        RECT 87.260 155.110 87.400 164.060 ;
        RECT 87.720 156.130 87.860 165.330 ;
        RECT 87.660 155.810 87.920 156.130 ;
        RECT 87.200 154.790 87.460 155.110 ;
        RECT 86.740 154.450 87.000 154.770 ;
        RECT 85.820 152.070 86.080 152.390 ;
        RECT 84.900 151.050 85.160 151.370 ;
        RECT 82.140 147.990 82.400 148.310 ;
        RECT 66.960 147.650 67.220 147.970 ;
        RECT 67.020 146.610 67.160 147.650 ;
        RECT 86.800 146.950 86.940 154.450 ;
        RECT 87.720 153.750 87.860 155.810 ;
        RECT 89.100 154.770 89.240 173.830 ;
        RECT 89.040 154.450 89.300 154.770 ;
        RECT 87.660 153.430 87.920 153.750 ;
        RECT 87.720 152.050 87.860 153.430 ;
        RECT 87.660 151.730 87.920 152.050 ;
        RECT 87.650 148.815 87.930 149.185 ;
        RECT 87.660 148.670 87.920 148.815 ;
        RECT 86.740 146.630 87.000 146.950 ;
        RECT 66.960 146.290 67.220 146.610 ;
        RECT 61.440 145.610 61.700 145.930 ;
        RECT 65.120 145.610 65.380 145.930 ;
        RECT 66.040 145.610 66.300 145.930 ;
        RECT 60.980 145.270 61.240 145.590 ;
        RECT 60.060 143.570 60.320 143.890 ;
        RECT 61.040 143.210 61.180 145.270 ;
        RECT 65.180 143.550 65.320 145.610 ;
        RECT 66.100 143.550 66.240 145.610 ;
        RECT 87.190 145.415 87.470 145.785 ;
        RECT 87.200 145.270 87.460 145.415 ;
        RECT 65.120 143.230 65.380 143.550 ;
        RECT 66.040 143.230 66.300 143.550 ;
        RECT 60.980 142.890 61.240 143.210 ;
        RECT 87.660 142.890 87.920 143.210 ;
        RECT 57.760 142.550 58.020 142.870 ;
        RECT 48.560 142.210 48.820 142.530 ;
        RECT 87.720 142.385 87.860 142.890 ;
        RECT 44.880 141.190 45.140 141.510 ;
        RECT 45.340 141.190 45.600 141.510 ;
        RECT 43.960 140.850 44.220 141.170 ;
        RECT 42.580 140.510 42.840 140.830 ;
        RECT 45.400 140.490 45.540 141.190 ;
        RECT 48.620 140.490 48.760 142.210 ;
        RECT 87.650 142.015 87.930 142.385 ;
        RECT 25.560 140.170 25.820 140.490 ;
        RECT 35.220 140.170 35.480 140.490 ;
        RECT 38.900 140.170 39.160 140.490 ;
        RECT 42.120 140.400 42.380 140.490 ;
        RECT 41.720 140.260 42.380 140.400 ;
        RECT 25.620 132.260 25.760 140.170 ;
        RECT 35.280 132.260 35.420 140.170 ;
        RECT 36.950 138.955 38.490 139.325 ;
        RECT 38.960 134.790 39.100 140.170 ;
        RECT 38.500 134.650 39.100 134.790 ;
        RECT 38.500 132.260 38.640 134.650 ;
        RECT 41.720 132.260 41.860 140.260 ;
        RECT 42.120 140.170 42.380 140.260 ;
        RECT 45.340 140.170 45.600 140.490 ;
        RECT 48.560 140.170 48.820 140.490 ;
        RECT 44.880 139.830 45.140 140.150 ;
        RECT 44.940 132.260 45.080 139.830 ;
        RECT 48.100 139.490 48.360 139.810 ;
        RECT 48.160 132.260 48.300 139.490 ;
        RECT 25.550 128.260 25.830 132.260 ;
        RECT 35.210 128.260 35.490 132.260 ;
        RECT 38.430 128.260 38.710 132.260 ;
        RECT 41.650 128.260 41.930 132.260 ;
        RECT 44.870 128.260 45.150 132.260 ;
        RECT 48.090 128.260 48.370 132.260 ;
      LAYER met3 ;
        RECT 31.250 220.550 31.630 220.560 ;
        RECT 90.930 220.550 94.930 220.700 ;
        RECT 31.250 220.250 94.930 220.550 ;
        RECT 31.250 220.240 31.630 220.250 ;
        RECT 90.930 220.100 94.930 220.250 ;
        RECT 22.765 217.150 23.095 217.165 ;
        RECT 90.930 217.150 94.930 217.300 ;
        RECT 22.765 216.850 94.930 217.150 ;
        RECT 22.765 216.835 23.095 216.850 ;
        RECT 90.930 216.700 94.930 216.850 ;
        RECT 18.370 216.470 18.750 216.480 ;
        RECT 77.045 216.470 77.375 216.485 ;
        RECT 18.370 216.170 77.375 216.470 ;
        RECT 18.370 216.160 18.750 216.170 ;
        RECT 77.045 216.155 77.375 216.170 ;
        RECT 12.645 214.430 12.975 214.445 ;
        RECT 26.650 214.430 27.030 214.440 ;
        RECT 12.645 214.130 27.030 214.430 ;
        RECT 12.645 214.115 12.975 214.130 ;
        RECT 26.650 214.120 27.030 214.130 ;
        RECT 64.165 214.430 64.495 214.445 ;
        RECT 79.805 214.430 80.135 214.445 ;
        RECT 64.165 214.130 80.135 214.430 ;
        RECT 64.165 214.115 64.495 214.130 ;
        RECT 79.805 214.115 80.135 214.130 ;
        RECT 42.290 213.750 42.670 213.760 ;
        RECT 67.385 213.750 67.715 213.765 ;
        RECT 42.290 213.450 67.715 213.750 ;
        RECT 42.290 213.440 42.670 213.450 ;
        RECT 67.385 213.435 67.715 213.450 ;
        RECT 68.765 213.750 69.095 213.765 ;
        RECT 90.930 213.750 94.930 213.900 ;
        RECT 68.765 213.450 94.930 213.750 ;
        RECT 68.765 213.435 69.095 213.450 ;
        RECT 90.930 213.300 94.930 213.450 ;
        RECT 31.505 212.390 31.835 212.405 ;
        RECT 51.285 212.390 51.615 212.405 ;
        RECT 31.505 212.090 51.615 212.390 ;
        RECT 31.505 212.075 31.835 212.090 ;
        RECT 51.285 212.075 51.615 212.090 ;
        RECT 58.850 212.390 59.230 212.400 ;
        RECT 83.485 212.390 83.815 212.405 ;
        RECT 58.850 212.090 83.815 212.390 ;
        RECT 58.850 212.080 59.230 212.090 ;
        RECT 83.485 212.075 83.815 212.090 ;
        RECT 22.970 211.710 23.350 211.720 ;
        RECT 25.525 211.710 25.855 211.725 ;
        RECT 22.970 211.410 25.855 211.710 ;
        RECT 22.970 211.400 23.350 211.410 ;
        RECT 25.525 211.395 25.855 211.410 ;
        RECT 30.125 211.710 30.455 211.725 ;
        RECT 45.050 211.710 45.430 211.720 ;
        RECT 30.125 211.410 45.430 211.710 ;
        RECT 30.125 211.395 30.455 211.410 ;
        RECT 45.050 211.400 45.430 211.410 ;
        RECT 56.090 211.710 56.470 211.720 ;
        RECT 73.825 211.710 74.155 211.725 ;
        RECT 93.145 211.710 93.475 211.725 ;
        RECT 56.090 211.410 74.155 211.710 ;
        RECT 56.090 211.400 56.470 211.410 ;
        RECT 73.825 211.395 74.155 211.410 ;
        RECT 74.530 211.410 93.475 211.710 ;
        RECT 20.925 211.030 21.255 211.045 ;
        RECT 39.785 211.030 40.115 211.045 ;
        RECT 20.925 210.730 40.115 211.030 ;
        RECT 20.925 210.715 21.255 210.730 ;
        RECT 39.785 210.715 40.115 210.730 ;
        RECT 56.345 211.030 56.675 211.045 ;
        RECT 74.530 211.030 74.830 211.410 ;
        RECT 93.145 211.395 93.475 211.410 ;
        RECT 56.345 210.730 74.830 211.030 ;
        RECT 56.345 210.715 56.675 210.730 ;
        RECT 12.580 210.350 16.580 210.500 ;
        RECT 17.705 210.350 18.035 210.365 ;
        RECT 12.580 210.050 18.035 210.350 ;
        RECT 12.580 209.900 16.580 210.050 ;
        RECT 17.705 210.035 18.035 210.050 ;
        RECT 57.725 210.350 58.055 210.365 ;
        RECT 87.625 210.350 87.955 210.365 ;
        RECT 90.930 210.350 94.930 210.500 ;
        RECT 57.725 210.050 87.955 210.350 ;
        RECT 57.725 210.035 58.055 210.050 ;
        RECT 87.625 210.035 87.955 210.050 ;
        RECT 88.330 210.050 94.930 210.350 ;
        RECT 36.930 209.695 38.510 210.025 ;
        RECT 23.225 209.670 23.555 209.685 ;
        RECT 35.185 209.670 35.515 209.685 ;
        RECT 23.225 209.370 35.515 209.670 ;
        RECT 23.225 209.355 23.555 209.370 ;
        RECT 35.185 209.355 35.515 209.370 ;
        RECT 38.865 209.670 39.195 209.685 ;
        RECT 71.985 209.670 72.315 209.685 ;
        RECT 38.865 209.370 72.315 209.670 ;
        RECT 38.865 209.355 39.195 209.370 ;
        RECT 71.985 209.355 72.315 209.370 ;
        RECT 79.090 209.670 79.470 209.680 ;
        RECT 88.330 209.670 88.630 210.050 ;
        RECT 90.930 209.900 94.930 210.050 ;
        RECT 79.090 209.370 88.630 209.670 ;
        RECT 79.090 209.360 79.470 209.370 ;
        RECT 30.585 208.990 30.915 209.005 ;
        RECT 82.105 208.990 82.435 209.005 ;
        RECT 30.585 208.690 82.435 208.990 ;
        RECT 30.585 208.675 30.915 208.690 ;
        RECT 82.105 208.675 82.435 208.690 ;
        RECT 24.810 208.310 25.190 208.320 ;
        RECT 25.985 208.310 26.315 208.325 ;
        RECT 33.805 208.310 34.135 208.325 ;
        RECT 37.485 208.310 37.815 208.325 ;
        RECT 24.810 208.010 26.315 208.310 ;
        RECT 24.810 208.000 25.190 208.010 ;
        RECT 25.985 207.995 26.315 208.010 ;
        RECT 27.610 208.010 37.815 208.310 ;
        RECT 12.580 206.950 16.580 207.100 ;
        RECT 19.085 206.950 19.415 206.965 ;
        RECT 12.580 206.650 19.415 206.950 ;
        RECT 12.580 206.500 16.580 206.650 ;
        RECT 19.085 206.635 19.415 206.650 ;
        RECT 21.385 205.590 21.715 205.605 ;
        RECT 27.610 205.600 27.910 208.010 ;
        RECT 33.805 207.995 34.135 208.010 ;
        RECT 37.485 207.995 37.815 208.010 ;
        RECT 38.405 208.310 38.735 208.325 ;
        RECT 43.925 208.310 44.255 208.325 ;
        RECT 83.025 208.310 83.355 208.325 ;
        RECT 38.405 208.010 83.355 208.310 ;
        RECT 38.405 207.995 38.735 208.010 ;
        RECT 43.925 207.995 44.255 208.010 ;
        RECT 83.025 207.995 83.355 208.010 ;
        RECT 85.530 208.310 85.910 208.320 ;
        RECT 86.245 208.310 86.575 208.325 ;
        RECT 85.530 208.010 86.575 208.310 ;
        RECT 85.530 208.000 85.910 208.010 ;
        RECT 86.245 207.995 86.575 208.010 ;
        RECT 37.945 207.630 38.275 207.645 ;
        RECT 43.005 207.630 43.335 207.645 ;
        RECT 37.945 207.330 43.335 207.630 ;
        RECT 37.945 207.315 38.275 207.330 ;
        RECT 43.005 207.315 43.335 207.330 ;
        RECT 57.010 207.630 57.390 207.640 ;
        RECT 58.185 207.630 58.515 207.645 ;
        RECT 79.345 207.630 79.675 207.645 ;
        RECT 57.010 207.330 79.675 207.630 ;
        RECT 57.010 207.320 57.390 207.330 ;
        RECT 58.185 207.315 58.515 207.330 ;
        RECT 79.345 207.315 79.675 207.330 ;
        RECT 33.630 206.975 35.210 207.305 ;
        RECT 46.225 206.950 46.555 206.965 ;
        RECT 77.250 206.950 77.630 206.960 ;
        RECT 90.930 206.950 94.930 207.100 ;
        RECT 35.890 206.650 61.030 206.950 ;
        RECT 28.285 206.270 28.615 206.285 ;
        RECT 35.890 206.270 36.190 206.650 ;
        RECT 46.225 206.635 46.555 206.650 ;
        RECT 28.285 205.970 36.190 206.270 ;
        RECT 37.485 206.270 37.815 206.285 ;
        RECT 46.890 206.270 47.270 206.280 ;
        RECT 37.485 205.970 47.270 206.270 ;
        RECT 60.730 206.270 61.030 206.650 ;
        RECT 77.250 206.650 94.930 206.950 ;
        RECT 77.250 206.640 77.630 206.650 ;
        RECT 90.930 206.500 94.930 206.650 ;
        RECT 87.625 206.270 87.955 206.285 ;
        RECT 60.730 205.970 87.955 206.270 ;
        RECT 28.285 205.955 28.615 205.970 ;
        RECT 37.485 205.955 37.815 205.970 ;
        RECT 46.890 205.960 47.270 205.970 ;
        RECT 87.625 205.955 87.955 205.970 ;
        RECT 27.570 205.590 27.950 205.600 ;
        RECT 21.385 205.290 27.950 205.590 ;
        RECT 21.385 205.275 21.715 205.290 ;
        RECT 27.570 205.280 27.950 205.290 ;
        RECT 29.205 205.590 29.535 205.605 ;
        RECT 67.845 205.590 68.175 205.605 ;
        RECT 29.205 205.290 68.175 205.590 ;
        RECT 29.205 205.275 29.535 205.290 ;
        RECT 67.845 205.275 68.175 205.290 ;
        RECT 71.985 205.590 72.315 205.605 ;
        RECT 81.185 205.590 81.515 205.605 ;
        RECT 71.985 205.290 81.515 205.590 ;
        RECT 71.985 205.275 72.315 205.290 ;
        RECT 81.185 205.275 81.515 205.290 ;
        RECT 25.985 204.910 26.315 204.925 ;
        RECT 29.220 204.910 29.520 205.275 ;
        RECT 25.985 204.610 29.520 204.910 ;
        RECT 30.125 204.910 30.455 204.925 ;
        RECT 39.325 204.920 39.655 204.925 ;
        RECT 35.850 204.910 36.230 204.920 ;
        RECT 30.125 204.610 36.230 204.910 ;
        RECT 25.985 204.595 26.315 204.610 ;
        RECT 30.125 204.595 30.455 204.610 ;
        RECT 35.850 204.600 36.230 204.610 ;
        RECT 39.325 204.910 39.910 204.920 ;
        RECT 54.250 204.910 54.630 204.920 ;
        RECT 55.425 204.910 55.755 204.925 ;
        RECT 39.325 204.610 40.110 204.910 ;
        RECT 54.250 204.610 55.755 204.910 ;
        RECT 39.325 204.600 39.910 204.610 ;
        RECT 54.250 204.600 54.630 204.610 ;
        RECT 39.325 204.595 39.655 204.600 ;
        RECT 55.425 204.595 55.755 204.610 ;
        RECT 69.225 204.910 69.555 204.925 ;
        RECT 69.890 204.910 70.270 204.920 ;
        RECT 69.225 204.610 70.270 204.910 ;
        RECT 69.225 204.595 69.555 204.610 ;
        RECT 69.890 204.600 70.270 204.610 ;
        RECT 71.730 204.910 72.110 204.920 ;
        RECT 84.865 204.910 85.195 204.925 ;
        RECT 71.730 204.610 85.195 204.910 ;
        RECT 71.730 204.600 72.110 204.610 ;
        RECT 84.865 204.595 85.195 204.610 ;
        RECT 36.930 204.255 38.510 204.585 ;
        RECT 25.525 204.230 25.855 204.245 ;
        RECT 36.105 204.230 36.435 204.245 ;
        RECT 25.525 203.930 36.435 204.230 ;
        RECT 25.525 203.915 25.855 203.930 ;
        RECT 36.105 203.915 36.435 203.930 ;
        RECT 38.865 204.230 39.195 204.245 ;
        RECT 57.265 204.230 57.595 204.245 ;
        RECT 38.865 203.930 73.910 204.230 ;
        RECT 38.865 203.915 39.195 203.930 ;
        RECT 57.265 203.915 57.595 203.930 ;
        RECT 12.580 203.550 16.580 203.700 ;
        RECT 18.625 203.550 18.955 203.565 ;
        RECT 12.580 203.250 18.955 203.550 ;
        RECT 12.580 203.100 16.580 203.250 ;
        RECT 18.625 203.235 18.955 203.250 ;
        RECT 27.825 203.550 28.155 203.565 ;
        RECT 30.585 203.550 30.915 203.565 ;
        RECT 68.970 203.550 69.350 203.560 ;
        RECT 71.985 203.550 72.315 203.565 ;
        RECT 27.825 203.250 30.915 203.550 ;
        RECT 27.825 203.235 28.155 203.250 ;
        RECT 30.585 203.235 30.915 203.250 ;
        RECT 32.210 203.250 72.315 203.550 ;
        RECT 73.610 203.550 73.910 203.930 ;
        RECT 74.285 203.550 74.615 203.565 ;
        RECT 73.610 203.250 74.615 203.550 ;
        RECT 27.365 202.190 27.695 202.205 ;
        RECT 32.210 202.190 32.510 203.250 ;
        RECT 68.970 203.240 69.350 203.250 ;
        RECT 71.985 203.235 72.315 203.250 ;
        RECT 74.285 203.235 74.615 203.250 ;
        RECT 78.170 203.550 78.550 203.560 ;
        RECT 90.930 203.550 94.930 203.700 ;
        RECT 78.170 203.250 94.930 203.550 ;
        RECT 78.170 203.240 78.550 203.250 ;
        RECT 90.930 203.100 94.930 203.250 ;
        RECT 33.805 202.870 34.135 202.885 ;
        RECT 41.370 202.870 41.750 202.880 ;
        RECT 33.805 202.570 41.750 202.870 ;
        RECT 33.805 202.555 34.135 202.570 ;
        RECT 41.370 202.560 41.750 202.570 ;
        RECT 42.545 202.870 42.875 202.885 ;
        RECT 57.010 202.870 57.390 202.880 ;
        RECT 42.545 202.570 57.390 202.870 ;
        RECT 42.545 202.555 42.875 202.570 ;
        RECT 57.010 202.560 57.390 202.570 ;
        RECT 59.105 202.870 59.435 202.885 ;
        RECT 59.770 202.870 60.150 202.880 ;
        RECT 59.105 202.570 60.150 202.870 ;
        RECT 59.105 202.555 59.435 202.570 ;
        RECT 59.770 202.560 60.150 202.570 ;
        RECT 27.365 201.890 32.510 202.190 ;
        RECT 36.565 202.190 36.895 202.205 ;
        RECT 44.130 202.190 44.510 202.200 ;
        RECT 36.565 201.890 44.510 202.190 ;
        RECT 27.365 201.875 27.695 201.890 ;
        RECT 36.565 201.875 36.895 201.890 ;
        RECT 44.130 201.880 44.510 201.890 ;
        RECT 46.685 202.190 47.015 202.205 ;
        RECT 52.410 202.190 52.790 202.200 ;
        RECT 72.905 202.190 73.235 202.205 ;
        RECT 46.685 201.890 73.235 202.190 ;
        RECT 46.685 201.875 47.015 201.890 ;
        RECT 52.410 201.880 52.790 201.890 ;
        RECT 72.905 201.875 73.235 201.890 ;
        RECT 33.630 201.535 35.210 201.865 ;
        RECT 23.685 201.510 24.015 201.525 ;
        RECT 24.810 201.510 25.190 201.520 ;
        RECT 23.685 201.210 25.190 201.510 ;
        RECT 23.685 201.195 24.015 201.210 ;
        RECT 24.810 201.200 25.190 201.210 ;
        RECT 26.445 201.510 26.775 201.525 ;
        RECT 31.965 201.510 32.295 201.525 ;
        RECT 26.445 201.210 32.295 201.510 ;
        RECT 26.445 201.195 26.775 201.210 ;
        RECT 31.965 201.195 32.295 201.210 ;
        RECT 36.105 201.510 36.435 201.525 ;
        RECT 38.405 201.510 38.735 201.525 ;
        RECT 40.450 201.510 40.830 201.520 ;
        RECT 36.105 201.210 40.830 201.510 ;
        RECT 36.105 201.195 36.435 201.210 ;
        RECT 38.405 201.195 38.735 201.210 ;
        RECT 40.450 201.200 40.830 201.210 ;
        RECT 42.545 201.510 42.875 201.525 ;
        RECT 65.290 201.510 65.670 201.520 ;
        RECT 66.005 201.510 66.335 201.525 ;
        RECT 42.545 201.210 66.335 201.510 ;
        RECT 42.545 201.195 42.875 201.210 ;
        RECT 65.290 201.200 65.670 201.210 ;
        RECT 66.005 201.195 66.335 201.210 ;
        RECT 73.570 201.510 73.950 201.520 ;
        RECT 75.665 201.510 75.995 201.525 ;
        RECT 73.570 201.210 75.995 201.510 ;
        RECT 73.570 201.200 73.950 201.210 ;
        RECT 75.665 201.195 75.995 201.210 ;
        RECT 28.490 200.830 28.870 200.840 ;
        RECT 32.885 200.830 33.215 200.845 ;
        RECT 28.490 200.530 33.215 200.830 ;
        RECT 28.490 200.520 28.870 200.530 ;
        RECT 32.885 200.515 33.215 200.530 ;
        RECT 33.805 200.830 34.135 200.845 ;
        RECT 52.205 200.830 52.535 200.845 ;
        RECT 33.805 200.530 52.535 200.830 ;
        RECT 33.805 200.515 34.135 200.530 ;
        RECT 52.205 200.515 52.535 200.530 ;
        RECT 12.580 200.150 16.580 200.300 ;
        RECT 17.705 200.150 18.035 200.165 ;
        RECT 12.580 199.850 18.035 200.150 ;
        RECT 12.580 199.700 16.580 199.850 ;
        RECT 17.705 199.835 18.035 199.850 ;
        RECT 25.065 200.150 25.395 200.165 ;
        RECT 35.645 200.150 35.975 200.165 ;
        RECT 45.970 200.150 46.350 200.160 ;
        RECT 25.065 199.850 31.820 200.150 ;
        RECT 25.065 199.835 25.395 199.850 ;
        RECT 26.445 199.470 26.775 199.485 ;
        RECT 30.330 199.470 30.710 199.480 ;
        RECT 26.445 199.170 30.710 199.470 ;
        RECT 31.520 199.470 31.820 199.850 ;
        RECT 35.645 199.850 46.350 200.150 ;
        RECT 35.645 199.835 35.975 199.850 ;
        RECT 45.970 199.840 46.350 199.850 ;
        RECT 55.170 200.150 55.550 200.160 ;
        RECT 59.565 200.150 59.895 200.165 ;
        RECT 55.170 199.850 59.895 200.150 ;
        RECT 55.170 199.840 55.550 199.850 ;
        RECT 59.565 199.835 59.895 199.850 ;
        RECT 75.410 200.150 75.790 200.160 ;
        RECT 90.930 200.150 94.930 200.300 ;
        RECT 75.410 199.850 94.930 200.150 ;
        RECT 75.410 199.840 75.790 199.850 ;
        RECT 90.930 199.700 94.930 199.850 ;
        RECT 36.105 199.470 36.435 199.485 ;
        RECT 31.520 199.170 36.435 199.470 ;
        RECT 26.445 199.155 26.775 199.170 ;
        RECT 30.330 199.160 30.710 199.170 ;
        RECT 36.105 199.155 36.435 199.170 ;
        RECT 39.785 199.470 40.115 199.485 ;
        RECT 60.690 199.470 61.070 199.480 ;
        RECT 71.525 199.470 71.855 199.485 ;
        RECT 39.785 199.170 71.855 199.470 ;
        RECT 39.785 199.155 40.115 199.170 ;
        RECT 60.690 199.160 61.070 199.170 ;
        RECT 71.525 199.155 71.855 199.170 ;
        RECT 82.770 199.470 83.150 199.480 ;
        RECT 84.405 199.470 84.735 199.485 ;
        RECT 82.770 199.170 84.735 199.470 ;
        RECT 82.770 199.160 83.150 199.170 ;
        RECT 84.405 199.155 84.735 199.170 ;
        RECT 36.930 198.815 38.510 199.145 ;
        RECT 24.810 198.790 25.190 198.800 ;
        RECT 27.825 198.790 28.155 198.805 ;
        RECT 24.810 198.490 28.155 198.790 ;
        RECT 24.810 198.480 25.190 198.490 ;
        RECT 27.825 198.475 28.155 198.490 ;
        RECT 32.170 198.790 32.550 198.800 ;
        RECT 34.265 198.790 34.595 198.805 ;
        RECT 32.170 198.490 34.595 198.790 ;
        RECT 32.170 198.480 32.550 198.490 ;
        RECT 34.265 198.475 34.595 198.490 ;
        RECT 38.865 198.790 39.195 198.805 ;
        RECT 51.745 198.790 52.075 198.805 ;
        RECT 38.865 198.490 52.075 198.790 ;
        RECT 38.865 198.475 39.195 198.490 ;
        RECT 51.745 198.475 52.075 198.490 ;
        RECT 57.725 198.790 58.055 198.805 ;
        RECT 80.725 198.790 81.055 198.805 ;
        RECT 57.725 198.490 81.055 198.790 ;
        RECT 57.725 198.475 58.055 198.490 ;
        RECT 80.725 198.475 81.055 198.490 ;
        RECT 31.505 198.110 31.835 198.125 ;
        RECT 33.345 198.110 33.675 198.125 ;
        RECT 38.880 198.110 39.180 198.475 ;
        RECT 31.505 197.810 39.180 198.110 ;
        RECT 47.145 198.110 47.475 198.125 ;
        RECT 81.645 198.110 81.975 198.125 ;
        RECT 47.145 197.810 81.975 198.110 ;
        RECT 31.505 197.795 31.835 197.810 ;
        RECT 33.345 197.795 33.675 197.810 ;
        RECT 47.145 197.795 47.475 197.810 ;
        RECT 81.645 197.795 81.975 197.810 ;
        RECT 40.450 197.430 40.830 197.440 ;
        RECT 41.625 197.430 41.955 197.445 ;
        RECT 32.210 197.130 36.190 197.430 ;
        RECT 12.580 196.750 16.580 196.900 ;
        RECT 20.005 196.750 20.335 196.765 ;
        RECT 12.580 196.450 20.335 196.750 ;
        RECT 12.580 196.300 16.580 196.450 ;
        RECT 20.005 196.435 20.335 196.450 ;
        RECT 26.905 196.070 27.235 196.085 ;
        RECT 27.825 196.070 28.155 196.085 ;
        RECT 32.210 196.070 32.510 197.130 ;
        RECT 35.890 196.750 36.190 197.130 ;
        RECT 40.450 197.130 41.955 197.430 ;
        RECT 40.450 197.120 40.830 197.130 ;
        RECT 41.625 197.115 41.955 197.130 ;
        RECT 43.005 197.440 43.335 197.445 ;
        RECT 43.005 197.430 43.590 197.440 ;
        RECT 44.385 197.430 44.715 197.445 ;
        RECT 58.645 197.430 58.975 197.445 ;
        RECT 43.005 197.130 43.790 197.430 ;
        RECT 44.385 197.130 58.975 197.430 ;
        RECT 43.005 197.120 43.590 197.130 ;
        RECT 43.005 197.115 43.335 197.120 ;
        RECT 44.385 197.115 44.715 197.130 ;
        RECT 58.645 197.115 58.975 197.130 ;
        RECT 66.925 197.440 67.255 197.445 ;
        RECT 66.925 197.430 67.510 197.440 ;
        RECT 66.925 197.130 67.710 197.430 ;
        RECT 66.925 197.120 67.510 197.130 ;
        RECT 66.925 197.115 67.255 197.120 ;
        RECT 48.985 196.750 49.315 196.765 ;
        RECT 60.485 196.750 60.815 196.765 ;
        RECT 35.890 196.450 43.550 196.750 ;
        RECT 33.630 196.095 35.210 196.425 ;
        RECT 26.905 195.770 32.510 196.070 ;
        RECT 36.105 196.070 36.435 196.085 ;
        RECT 39.325 196.070 39.655 196.085 ;
        RECT 40.705 196.080 41.035 196.085 ;
        RECT 40.450 196.070 41.035 196.080 ;
        RECT 36.105 195.770 39.655 196.070 ;
        RECT 40.250 195.770 41.035 196.070 ;
        RECT 26.905 195.755 27.235 195.770 ;
        RECT 27.825 195.755 28.155 195.770 ;
        RECT 36.105 195.755 36.435 195.770 ;
        RECT 39.325 195.755 39.655 195.770 ;
        RECT 40.450 195.760 41.035 195.770 ;
        RECT 40.705 195.755 41.035 195.760 ;
        RECT 30.585 195.390 30.915 195.405 ;
        RECT 42.290 195.390 42.670 195.400 ;
        RECT 30.585 195.090 42.670 195.390 ;
        RECT 43.250 195.390 43.550 196.450 ;
        RECT 48.985 196.450 60.815 196.750 ;
        RECT 48.985 196.435 49.315 196.450 ;
        RECT 60.485 196.435 60.815 196.450 ;
        RECT 66.210 196.750 66.590 196.760 ;
        RECT 68.765 196.750 69.095 196.765 ;
        RECT 90.930 196.750 94.930 196.900 ;
        RECT 66.210 196.450 69.095 196.750 ;
        RECT 66.210 196.440 66.590 196.450 ;
        RECT 68.765 196.435 69.095 196.450 ;
        RECT 74.530 196.450 94.930 196.750 ;
        RECT 53.125 196.070 53.455 196.085 ;
        RECT 74.530 196.070 74.830 196.450 ;
        RECT 90.930 196.300 94.930 196.450 ;
        RECT 53.125 195.770 74.830 196.070 ;
        RECT 53.125 195.755 53.455 195.770 ;
        RECT 69.225 195.390 69.555 195.405 ;
        RECT 43.250 195.090 69.555 195.390 ;
        RECT 30.585 195.075 30.915 195.090 ;
        RECT 42.290 195.080 42.670 195.090 ;
        RECT 69.225 195.075 69.555 195.090 ;
        RECT 25.730 194.710 26.110 194.720 ;
        RECT 28.745 194.710 29.075 194.725 ;
        RECT 31.505 194.720 31.835 194.725 ;
        RECT 31.250 194.710 31.835 194.720 ;
        RECT 39.785 194.710 40.115 194.725 ;
        RECT 25.730 194.410 29.075 194.710 ;
        RECT 31.050 194.410 31.835 194.710 ;
        RECT 25.730 194.400 26.110 194.410 ;
        RECT 28.745 194.395 29.075 194.410 ;
        RECT 31.250 194.400 31.835 194.410 ;
        RECT 31.505 194.395 31.835 194.400 ;
        RECT 36.120 194.410 40.115 194.710 ;
        RECT 24.605 194.030 24.935 194.045 ;
        RECT 36.120 194.030 36.420 194.410 ;
        RECT 39.785 194.395 40.115 194.410 ;
        RECT 42.290 194.710 42.670 194.720 ;
        RECT 43.925 194.710 44.255 194.725 ;
        RECT 42.290 194.410 44.255 194.710 ;
        RECT 42.290 194.400 42.670 194.410 ;
        RECT 43.925 194.395 44.255 194.410 ;
        RECT 46.225 194.710 46.555 194.725 ;
        RECT 50.365 194.710 50.695 194.725 ;
        RECT 46.225 194.410 50.695 194.710 ;
        RECT 46.225 194.395 46.555 194.410 ;
        RECT 50.365 194.395 50.695 194.410 ;
        RECT 59.770 194.710 60.150 194.720 ;
        RECT 82.565 194.710 82.895 194.725 ;
        RECT 59.770 194.410 82.895 194.710 ;
        RECT 59.770 194.400 60.150 194.410 ;
        RECT 82.565 194.395 82.895 194.410 ;
        RECT 24.605 193.730 36.420 194.030 ;
        RECT 43.005 194.030 43.335 194.045 ;
        RECT 47.810 194.030 48.190 194.040 ;
        RECT 83.025 194.030 83.355 194.045 ;
        RECT 43.005 193.730 83.355 194.030 ;
        RECT 24.605 193.715 24.935 193.730 ;
        RECT 43.005 193.715 43.335 193.730 ;
        RECT 47.810 193.720 48.190 193.730 ;
        RECT 83.025 193.715 83.355 193.730 ;
        RECT 12.580 193.350 16.580 193.500 ;
        RECT 36.930 193.375 38.510 193.705 ;
        RECT 17.245 193.350 17.575 193.365 ;
        RECT 12.580 193.050 17.575 193.350 ;
        RECT 12.580 192.900 16.580 193.050 ;
        RECT 17.245 193.035 17.575 193.050 ;
        RECT 25.525 193.350 25.855 193.365 ;
        RECT 33.805 193.350 34.135 193.365 ;
        RECT 25.525 193.050 34.135 193.350 ;
        RECT 25.525 193.035 25.855 193.050 ;
        RECT 33.805 193.035 34.135 193.050 ;
        RECT 47.145 193.350 47.475 193.365 ;
        RECT 55.425 193.350 55.755 193.365 ;
        RECT 47.145 193.050 55.755 193.350 ;
        RECT 47.145 193.035 47.475 193.050 ;
        RECT 55.425 193.035 55.755 193.050 ;
        RECT 75.665 193.350 75.995 193.365 ;
        RECT 90.930 193.350 94.930 193.500 ;
        RECT 75.665 193.050 94.930 193.350 ;
        RECT 75.665 193.035 75.995 193.050 ;
        RECT 90.930 192.900 94.930 193.050 ;
        RECT 33.345 192.670 33.675 192.685 ;
        RECT 49.445 192.670 49.775 192.685 ;
        RECT 33.345 192.370 49.775 192.670 ;
        RECT 33.345 192.355 33.675 192.370 ;
        RECT 49.445 192.355 49.775 192.370 ;
        RECT 31.505 191.990 31.835 192.005 ;
        RECT 35.185 191.990 35.515 192.005 ;
        RECT 31.505 191.690 35.515 191.990 ;
        RECT 31.505 191.675 31.835 191.690 ;
        RECT 35.185 191.675 35.515 191.690 ;
        RECT 39.325 191.990 39.655 192.005 ;
        RECT 83.485 191.990 83.815 192.005 ;
        RECT 89.005 191.990 89.335 192.005 ;
        RECT 39.325 191.690 89.335 191.990 ;
        RECT 39.325 191.675 39.655 191.690 ;
        RECT 83.485 191.675 83.815 191.690 ;
        RECT 89.005 191.675 89.335 191.690 ;
        RECT 28.490 191.310 28.870 191.320 ;
        RECT 32.885 191.310 33.215 191.325 ;
        RECT 37.485 191.310 37.815 191.325 ;
        RECT 28.490 191.010 33.215 191.310 ;
        RECT 28.490 191.000 28.870 191.010 ;
        RECT 32.885 190.995 33.215 191.010 ;
        RECT 35.660 191.010 37.815 191.310 ;
        RECT 33.630 190.655 35.210 190.985 ;
        RECT 16.785 190.630 17.115 190.645 ;
        RECT 16.570 190.315 17.115 190.630 ;
        RECT 30.125 190.630 30.455 190.645 ;
        RECT 32.425 190.630 32.755 190.645 ;
        RECT 30.125 190.330 32.755 190.630 ;
        RECT 30.125 190.315 30.455 190.330 ;
        RECT 32.425 190.315 32.755 190.330 ;
        RECT 16.570 190.100 16.870 190.315 ;
        RECT 12.580 189.650 16.870 190.100 ;
        RECT 28.745 189.960 29.075 189.965 ;
        RECT 28.490 189.950 29.075 189.960 ;
        RECT 28.290 189.650 29.075 189.950 ;
        RECT 12.580 189.500 16.580 189.650 ;
        RECT 28.490 189.640 29.075 189.650 ;
        RECT 29.410 189.950 29.790 189.960 ;
        RECT 35.660 189.950 35.960 191.010 ;
        RECT 37.485 190.995 37.815 191.010 ;
        RECT 40.450 191.310 40.830 191.320 ;
        RECT 54.045 191.310 54.375 191.325 ;
        RECT 63.245 191.310 63.575 191.325 ;
        RECT 40.450 191.010 54.375 191.310 ;
        RECT 40.450 191.000 40.830 191.010 ;
        RECT 54.045 190.995 54.375 191.010 ;
        RECT 60.960 191.010 63.575 191.310 ;
        RECT 60.960 190.645 61.260 191.010 ;
        RECT 63.245 190.995 63.575 191.010 ;
        RECT 76.585 191.310 76.915 191.325 ;
        RECT 79.090 191.310 79.470 191.320 ;
        RECT 76.585 191.010 79.470 191.310 ;
        RECT 76.585 190.995 76.915 191.010 ;
        RECT 79.090 191.000 79.470 191.010 ;
        RECT 37.485 190.630 37.815 190.645 ;
        RECT 47.605 190.630 47.935 190.645 ;
        RECT 37.485 190.330 47.935 190.630 ;
        RECT 53.125 190.460 53.455 190.475 ;
        RECT 37.485 190.315 37.815 190.330 ;
        RECT 47.605 190.315 47.935 190.330 ;
        RECT 52.450 190.160 53.455 190.460 ;
        RECT 60.945 190.315 61.275 190.645 ;
        RECT 61.865 190.630 62.195 190.645 ;
        RECT 65.545 190.630 65.875 190.645 ;
        RECT 61.865 190.330 65.875 190.630 ;
        RECT 61.865 190.315 62.195 190.330 ;
        RECT 65.545 190.315 65.875 190.330 ;
        RECT 70.145 190.630 70.475 190.645 ;
        RECT 81.185 190.630 81.515 190.645 ;
        RECT 70.145 190.330 81.515 190.630 ;
        RECT 70.145 190.315 70.475 190.330 ;
        RECT 81.185 190.315 81.515 190.330 ;
        RECT 29.410 189.650 35.960 189.950 ;
        RECT 37.025 189.950 37.355 189.965 ;
        RECT 52.450 189.950 52.750 190.160 ;
        RECT 53.125 190.145 53.455 190.160 ;
        RECT 37.025 189.650 52.750 189.950 ;
        RECT 54.045 189.950 54.375 189.965 ;
        RECT 90.930 189.950 94.930 190.100 ;
        RECT 54.045 189.650 94.930 189.950 ;
        RECT 29.410 189.640 29.790 189.650 ;
        RECT 28.745 189.635 29.075 189.640 ;
        RECT 37.025 189.635 37.355 189.650 ;
        RECT 54.045 189.635 54.375 189.650 ;
        RECT 90.930 189.500 94.930 189.650 ;
        RECT 25.065 189.270 25.395 189.285 ;
        RECT 33.805 189.270 34.135 189.285 ;
        RECT 25.065 188.970 34.135 189.270 ;
        RECT 25.065 188.955 25.395 188.970 ;
        RECT 33.805 188.955 34.135 188.970 ;
        RECT 37.945 189.270 38.275 189.285 ;
        RECT 55.170 189.270 55.550 189.280 ;
        RECT 75.410 189.270 75.790 189.280 ;
        RECT 37.945 188.970 55.550 189.270 ;
        RECT 37.945 188.955 38.275 188.970 ;
        RECT 55.170 188.960 55.550 188.970 ;
        RECT 63.490 188.970 75.790 189.270 ;
        RECT 31.250 188.590 31.630 188.600 ;
        RECT 34.265 188.590 34.595 188.605 ;
        RECT 43.925 188.600 44.255 188.605 ;
        RECT 43.925 188.590 44.510 188.600 ;
        RECT 52.665 188.590 52.995 188.605 ;
        RECT 31.250 188.290 34.595 188.590 ;
        RECT 43.700 188.290 44.510 188.590 ;
        RECT 31.250 188.280 31.630 188.290 ;
        RECT 34.265 188.275 34.595 188.290 ;
        RECT 43.925 188.280 44.510 188.290 ;
        RECT 45.320 188.290 52.995 188.590 ;
        RECT 43.925 188.275 44.255 188.280 ;
        RECT 36.930 187.935 38.510 188.265 ;
        RECT 16.785 187.920 17.115 187.925 ;
        RECT 16.530 187.910 17.115 187.920 ;
        RECT 16.330 187.610 17.115 187.910 ;
        RECT 16.530 187.600 17.115 187.610 ;
        RECT 16.785 187.595 17.115 187.600 ;
        RECT 22.765 187.910 23.095 187.925 ;
        RECT 26.445 187.910 26.775 187.925 ;
        RECT 22.765 187.610 26.775 187.910 ;
        RECT 22.765 187.595 23.095 187.610 ;
        RECT 26.445 187.595 26.775 187.610 ;
        RECT 31.965 187.595 32.295 187.925 ;
        RECT 35.185 187.910 35.515 187.925 ;
        RECT 36.105 187.910 36.435 187.925 ;
        RECT 35.185 187.610 36.435 187.910 ;
        RECT 35.185 187.595 35.515 187.610 ;
        RECT 36.105 187.595 36.435 187.610 ;
        RECT 43.005 187.910 43.335 187.925 ;
        RECT 45.320 187.910 45.620 188.290 ;
        RECT 52.665 188.275 52.995 188.290 ;
        RECT 57.930 188.590 58.310 188.600 ;
        RECT 63.490 188.590 63.790 188.970 ;
        RECT 75.410 188.960 75.790 188.970 ;
        RECT 83.025 188.590 83.355 188.605 ;
        RECT 57.930 188.290 63.790 188.590 ;
        RECT 74.530 188.290 83.355 188.590 ;
        RECT 57.930 188.280 58.310 188.290 ;
        RECT 43.005 187.610 45.620 187.910 ;
        RECT 46.890 187.910 47.270 187.920 ;
        RECT 48.985 187.910 49.315 187.925 ;
        RECT 46.890 187.610 49.315 187.910 ;
        RECT 43.005 187.595 43.335 187.610 ;
        RECT 46.890 187.600 47.270 187.610 ;
        RECT 48.985 187.595 49.315 187.610 ;
        RECT 51.745 187.910 52.075 187.925 ;
        RECT 53.330 187.910 53.710 187.920 ;
        RECT 74.530 187.910 74.830 188.290 ;
        RECT 83.025 188.275 83.355 188.290 ;
        RECT 51.745 187.610 74.830 187.910 ;
        RECT 51.745 187.595 52.075 187.610 ;
        RECT 53.330 187.600 53.710 187.610 ;
        RECT 31.980 187.230 32.280 187.595 ;
        RECT 39.785 187.230 40.115 187.245 ;
        RECT 31.980 186.930 40.115 187.230 ;
        RECT 39.785 186.915 40.115 186.930 ;
        RECT 46.685 187.230 47.015 187.245 ;
        RECT 49.445 187.230 49.775 187.245 ;
        RECT 63.245 187.230 63.575 187.245 ;
        RECT 46.685 186.930 49.070 187.230 ;
        RECT 46.685 186.915 47.015 186.930 ;
        RECT 12.580 186.560 16.580 186.700 ;
        RECT 12.580 186.240 16.910 186.560 ;
        RECT 31.965 186.550 32.295 186.565 ;
        RECT 42.085 186.550 42.415 186.565 ;
        RECT 31.965 186.250 42.415 186.550 ;
        RECT 12.580 186.100 16.580 186.240 ;
        RECT 31.965 186.235 32.295 186.250 ;
        RECT 42.085 186.235 42.415 186.250 ;
        RECT 48.770 185.880 49.070 186.930 ;
        RECT 49.445 186.930 63.575 187.230 ;
        RECT 49.445 186.915 49.775 186.930 ;
        RECT 63.245 186.915 63.575 186.930 ;
        RECT 51.490 186.550 51.870 186.560 ;
        RECT 53.125 186.550 53.455 186.565 ;
        RECT 51.490 186.250 53.455 186.550 ;
        RECT 51.490 186.240 51.870 186.250 ;
        RECT 53.125 186.235 53.455 186.250 ;
        RECT 55.425 186.550 55.755 186.565 ;
        RECT 57.010 186.550 57.390 186.560 ;
        RECT 55.425 186.250 57.390 186.550 ;
        RECT 55.425 186.235 55.755 186.250 ;
        RECT 57.010 186.240 57.390 186.250 ;
        RECT 82.565 186.550 82.895 186.565 ;
        RECT 90.930 186.550 94.930 186.700 ;
        RECT 82.565 186.250 94.930 186.550 ;
        RECT 82.565 186.235 82.895 186.250 ;
        RECT 90.930 186.100 94.930 186.250 ;
        RECT 48.730 185.870 49.110 185.880 ;
        RECT 56.345 185.870 56.675 185.885 ;
        RECT 62.325 185.870 62.655 185.885 ;
        RECT 48.730 185.570 62.655 185.870 ;
        RECT 48.730 185.560 49.110 185.570 ;
        RECT 56.345 185.555 56.675 185.570 ;
        RECT 62.325 185.555 62.655 185.570 ;
        RECT 33.630 185.215 35.210 185.545 ;
        RECT 25.730 185.190 26.110 185.200 ;
        RECT 31.965 185.190 32.295 185.205 ;
        RECT 41.165 185.190 41.495 185.205 ;
        RECT 25.730 184.890 32.295 185.190 ;
        RECT 25.730 184.880 26.110 184.890 ;
        RECT 31.965 184.875 32.295 184.890 ;
        RECT 37.960 184.890 41.495 185.190 ;
        RECT 37.960 184.525 38.260 184.890 ;
        RECT 41.165 184.875 41.495 184.890 ;
        RECT 42.290 185.190 42.670 185.200 ;
        RECT 45.765 185.190 46.095 185.205 ;
        RECT 42.290 184.890 46.095 185.190 ;
        RECT 42.290 184.880 42.670 184.890 ;
        RECT 45.765 184.875 46.095 184.890 ;
        RECT 61.405 185.190 61.735 185.205 ;
        RECT 77.045 185.190 77.375 185.205 ;
        RECT 61.405 184.890 77.375 185.190 ;
        RECT 61.405 184.875 61.735 184.890 ;
        RECT 77.045 184.875 77.375 184.890 ;
        RECT 27.365 184.510 27.695 184.525 ;
        RECT 30.125 184.510 30.455 184.525 ;
        RECT 33.345 184.510 33.675 184.525 ;
        RECT 27.365 184.210 29.750 184.510 ;
        RECT 27.365 184.195 27.695 184.210 ;
        RECT 26.650 183.830 27.030 183.840 ;
        RECT 27.825 183.830 28.155 183.845 ;
        RECT 26.650 183.530 28.155 183.830 ;
        RECT 29.450 183.830 29.750 184.210 ;
        RECT 30.125 184.210 33.675 184.510 ;
        RECT 30.125 184.195 30.455 184.210 ;
        RECT 33.345 184.195 33.675 184.210 ;
        RECT 34.265 184.510 34.595 184.525 ;
        RECT 35.850 184.510 36.230 184.520 ;
        RECT 34.265 184.210 36.230 184.510 ;
        RECT 34.265 184.195 34.595 184.210 ;
        RECT 35.850 184.200 36.230 184.210 ;
        RECT 37.945 184.195 38.275 184.525 ;
        RECT 47.605 184.510 47.935 184.525 ;
        RECT 87.165 184.510 87.495 184.525 ;
        RECT 47.605 184.210 87.495 184.510 ;
        RECT 47.605 184.195 47.935 184.210 ;
        RECT 87.165 184.195 87.495 184.210 ;
        RECT 33.805 183.830 34.135 183.845 ;
        RECT 29.450 183.530 34.135 183.830 ;
        RECT 26.650 183.520 27.030 183.530 ;
        RECT 27.825 183.515 28.155 183.530 ;
        RECT 33.805 183.515 34.135 183.530 ;
        RECT 43.465 183.830 43.795 183.845 ;
        RECT 49.445 183.830 49.775 183.845 ;
        RECT 54.965 183.830 55.295 183.845 ;
        RECT 56.345 183.840 56.675 183.845 ;
        RECT 56.090 183.830 56.675 183.840 ;
        RECT 76.585 183.830 76.915 183.845 ;
        RECT 43.465 183.530 55.295 183.830 ;
        RECT 55.890 183.530 56.675 183.830 ;
        RECT 43.465 183.515 43.795 183.530 ;
        RECT 49.445 183.515 49.775 183.530 ;
        RECT 54.965 183.515 55.295 183.530 ;
        RECT 56.090 183.520 56.675 183.530 ;
        RECT 56.345 183.515 56.675 183.520 ;
        RECT 63.490 183.530 76.915 183.830 ;
        RECT 12.580 183.150 16.580 183.300 ;
        RECT 19.545 183.150 19.875 183.165 ;
        RECT 12.580 182.850 19.875 183.150 ;
        RECT 12.580 182.700 16.580 182.850 ;
        RECT 19.545 182.835 19.875 182.850 ;
        RECT 22.970 183.150 23.350 183.160 ;
        RECT 29.205 183.150 29.535 183.165 ;
        RECT 22.970 182.850 29.535 183.150 ;
        RECT 22.970 182.840 23.350 182.850 ;
        RECT 29.205 182.835 29.535 182.850 ;
        RECT 31.250 183.150 31.630 183.160 ;
        RECT 35.645 183.150 35.975 183.165 ;
        RECT 31.250 182.850 35.975 183.150 ;
        RECT 31.250 182.840 31.630 182.850 ;
        RECT 35.645 182.835 35.975 182.850 ;
        RECT 43.925 183.150 44.255 183.165 ;
        RECT 45.050 183.150 45.430 183.160 ;
        RECT 43.925 182.850 45.430 183.150 ;
        RECT 43.925 182.835 44.255 182.850 ;
        RECT 45.050 182.840 45.430 182.850 ;
        RECT 45.970 183.150 46.350 183.160 ;
        RECT 49.445 183.150 49.775 183.165 ;
        RECT 45.970 182.850 49.775 183.150 ;
        RECT 45.970 182.840 46.350 182.850 ;
        RECT 49.445 182.835 49.775 182.850 ;
        RECT 53.125 183.150 53.455 183.165 ;
        RECT 63.490 183.150 63.790 183.530 ;
        RECT 76.585 183.515 76.915 183.530 ;
        RECT 53.125 182.850 63.790 183.150 ;
        RECT 88.085 183.150 88.415 183.165 ;
        RECT 90.930 183.150 94.930 183.300 ;
        RECT 88.085 182.850 94.930 183.150 ;
        RECT 53.125 182.835 53.455 182.850 ;
        RECT 88.085 182.835 88.415 182.850 ;
        RECT 36.930 182.495 38.510 182.825 ;
        RECT 90.930 182.700 94.930 182.850 ;
        RECT 24.810 182.470 25.190 182.480 ;
        RECT 25.985 182.470 26.315 182.485 ;
        RECT 24.810 182.170 26.315 182.470 ;
        RECT 24.810 182.160 25.190 182.170 ;
        RECT 25.985 182.155 26.315 182.170 ;
        RECT 27.570 182.470 27.950 182.480 ;
        RECT 30.125 182.470 30.455 182.485 ;
        RECT 27.570 182.170 30.455 182.470 ;
        RECT 27.570 182.160 27.950 182.170 ;
        RECT 30.125 182.155 30.455 182.170 ;
        RECT 32.425 182.470 32.755 182.485 ;
        RECT 35.850 182.470 36.230 182.480 ;
        RECT 32.425 182.170 36.230 182.470 ;
        RECT 32.425 182.155 32.755 182.170 ;
        RECT 35.850 182.160 36.230 182.170 ;
        RECT 44.845 182.470 45.175 182.485 ;
        RECT 58.185 182.470 58.515 182.485 ;
        RECT 44.845 182.170 58.515 182.470 ;
        RECT 44.845 182.155 45.175 182.170 ;
        RECT 58.185 182.155 58.515 182.170 ;
        RECT 67.130 182.470 67.510 182.480 ;
        RECT 75.410 182.470 75.790 182.480 ;
        RECT 67.130 182.170 75.790 182.470 ;
        RECT 67.130 182.160 67.510 182.170 ;
        RECT 75.410 182.160 75.790 182.170 ;
        RECT 22.765 181.790 23.095 181.805 ;
        RECT 54.250 181.790 54.630 181.800 ;
        RECT 22.765 181.490 54.630 181.790 ;
        RECT 22.765 181.475 23.095 181.490 ;
        RECT 54.250 181.480 54.630 181.490 ;
        RECT 61.405 181.790 61.735 181.805 ;
        RECT 63.450 181.790 63.830 181.800 ;
        RECT 64.625 181.790 64.955 181.805 ;
        RECT 61.405 181.490 64.955 181.790 ;
        RECT 61.405 181.475 61.735 181.490 ;
        RECT 63.450 181.480 63.830 181.490 ;
        RECT 64.625 181.475 64.955 181.490 ;
        RECT 69.225 181.790 69.555 181.805 ;
        RECT 71.730 181.790 72.110 181.800 ;
        RECT 69.225 181.490 72.110 181.790 ;
        RECT 69.225 181.475 69.555 181.490 ;
        RECT 71.730 181.480 72.110 181.490 ;
        RECT 15.865 181.110 16.195 181.125 ;
        RECT 27.825 181.110 28.155 181.125 ;
        RECT 15.865 180.810 28.155 181.110 ;
        RECT 15.865 180.795 16.195 180.810 ;
        RECT 27.825 180.795 28.155 180.810 ;
        RECT 28.490 181.110 28.870 181.120 ;
        RECT 31.965 181.110 32.295 181.125 ;
        RECT 28.490 180.810 32.295 181.110 ;
        RECT 28.490 180.800 28.870 180.810 ;
        RECT 31.965 180.795 32.295 180.810 ;
        RECT 32.885 181.110 33.215 181.125 ;
        RECT 42.545 181.110 42.875 181.125 ;
        RECT 32.885 180.810 42.875 181.110 ;
        RECT 32.885 180.795 33.215 180.810 ;
        RECT 42.545 180.795 42.875 180.810 ;
        RECT 44.385 181.110 44.715 181.125 ;
        RECT 49.445 181.110 49.775 181.125 ;
        RECT 44.385 180.810 49.775 181.110 ;
        RECT 44.385 180.795 44.715 180.810 ;
        RECT 49.445 180.795 49.775 180.810 ;
        RECT 54.965 181.110 55.295 181.125 ;
        RECT 55.885 181.110 56.215 181.125 ;
        RECT 54.965 180.810 56.215 181.110 ;
        RECT 54.965 180.795 55.295 180.810 ;
        RECT 55.885 180.795 56.215 180.810 ;
        RECT 27.825 180.430 28.155 180.445 ;
        RECT 29.410 180.430 29.790 180.440 ;
        RECT 27.825 180.130 29.790 180.430 ;
        RECT 27.825 180.115 28.155 180.130 ;
        RECT 29.410 180.120 29.790 180.130 ;
        RECT 35.850 180.430 36.230 180.440 ;
        RECT 49.905 180.430 50.235 180.445 ;
        RECT 52.665 180.440 52.995 180.445 ;
        RECT 35.850 180.130 50.235 180.430 ;
        RECT 35.850 180.120 36.230 180.130 ;
        RECT 49.905 180.115 50.235 180.130 ;
        RECT 52.410 180.430 52.995 180.440 ;
        RECT 52.410 180.130 53.220 180.430 ;
        RECT 52.410 180.120 52.995 180.130 ;
        RECT 52.665 180.115 52.995 180.120 ;
        RECT 33.630 179.775 35.210 180.105 ;
        RECT 37.485 179.750 37.815 179.765 ;
        RECT 38.865 179.750 39.195 179.765 ;
        RECT 41.165 179.750 41.495 179.765 ;
        RECT 49.905 179.750 50.235 179.765 ;
        RECT 37.485 179.450 50.235 179.750 ;
        RECT 37.485 179.435 37.815 179.450 ;
        RECT 38.865 179.435 39.195 179.450 ;
        RECT 41.165 179.435 41.495 179.450 ;
        RECT 49.905 179.435 50.235 179.450 ;
        RECT 55.885 179.750 56.215 179.765 ;
        RECT 61.405 179.750 61.735 179.765 ;
        RECT 55.885 179.450 61.735 179.750 ;
        RECT 55.885 179.435 56.215 179.450 ;
        RECT 61.405 179.435 61.735 179.450 ;
        RECT 87.625 179.750 87.955 179.765 ;
        RECT 90.930 179.750 94.930 179.900 ;
        RECT 87.625 179.450 94.930 179.750 ;
        RECT 87.625 179.435 87.955 179.450 ;
        RECT 90.930 179.300 94.930 179.450 ;
        RECT 40.450 179.070 40.830 179.080 ;
        RECT 42.085 179.070 42.415 179.085 ;
        RECT 48.525 179.070 48.855 179.085 ;
        RECT 40.450 178.770 48.855 179.070 ;
        RECT 40.450 178.760 40.830 178.770 ;
        RECT 42.085 178.755 42.415 178.770 ;
        RECT 48.525 178.755 48.855 178.770 ;
        RECT 55.885 179.070 56.215 179.085 ;
        RECT 59.770 179.070 60.150 179.080 ;
        RECT 55.885 178.770 60.150 179.070 ;
        RECT 55.885 178.755 56.215 178.770 ;
        RECT 59.770 178.760 60.150 178.770 ;
        RECT 60.945 179.070 61.275 179.085 ;
        RECT 71.525 179.070 71.855 179.085 ;
        RECT 60.945 178.770 71.855 179.070 ;
        RECT 60.945 178.755 61.275 178.770 ;
        RECT 71.525 178.755 71.855 178.770 ;
        RECT 28.285 178.390 28.615 178.405 ;
        RECT 41.370 178.390 41.750 178.400 ;
        RECT 28.285 178.090 41.750 178.390 ;
        RECT 28.285 178.075 28.615 178.090 ;
        RECT 41.370 178.080 41.750 178.090 ;
        RECT 43.005 178.390 43.335 178.405 ;
        RECT 53.125 178.390 53.455 178.405 ;
        RECT 43.005 178.090 53.455 178.390 ;
        RECT 43.005 178.075 43.335 178.090 ;
        RECT 53.125 178.075 53.455 178.090 ;
        RECT 58.645 178.390 58.975 178.405 ;
        RECT 66.005 178.390 66.335 178.405 ;
        RECT 58.645 178.090 66.335 178.390 ;
        RECT 58.645 178.075 58.975 178.090 ;
        RECT 66.005 178.075 66.335 178.090 ;
        RECT 67.130 178.390 67.510 178.400 ;
        RECT 89.925 178.390 90.255 178.405 ;
        RECT 67.130 178.090 90.255 178.390 ;
        RECT 67.130 178.080 67.510 178.090 ;
        RECT 89.925 178.075 90.255 178.090 ;
        RECT 48.985 177.710 49.315 177.725 ;
        RECT 55.170 177.710 55.550 177.720 ;
        RECT 57.010 177.710 57.390 177.720 ;
        RECT 70.810 177.710 71.190 177.720 ;
        RECT 48.985 177.410 71.190 177.710 ;
        RECT 48.985 177.395 49.315 177.410 ;
        RECT 55.170 177.400 55.550 177.410 ;
        RECT 57.010 177.400 57.390 177.410 ;
        RECT 70.810 177.400 71.190 177.410 ;
        RECT 36.930 177.055 38.510 177.385 ;
        RECT 38.865 177.030 39.195 177.045 ;
        RECT 48.525 177.030 48.855 177.045 ;
        RECT 50.825 177.040 51.155 177.045 ;
        RECT 50.570 177.030 51.155 177.040 ;
        RECT 53.125 177.040 53.455 177.045 ;
        RECT 53.125 177.030 53.710 177.040 ;
        RECT 38.865 176.730 48.855 177.030 ;
        RECT 50.370 176.730 51.155 177.030 ;
        RECT 52.900 176.730 53.710 177.030 ;
        RECT 38.865 176.715 39.195 176.730 ;
        RECT 48.525 176.715 48.855 176.730 ;
        RECT 50.570 176.720 51.155 176.730 ;
        RECT 50.825 176.715 51.155 176.720 ;
        RECT 53.125 176.720 53.710 176.730 ;
        RECT 54.045 177.030 54.375 177.045 ;
        RECT 56.090 177.030 56.470 177.040 ;
        RECT 58.645 177.030 58.975 177.045 ;
        RECT 54.045 176.730 58.975 177.030 ;
        RECT 53.125 176.715 53.455 176.720 ;
        RECT 54.045 176.715 54.375 176.730 ;
        RECT 56.090 176.720 56.470 176.730 ;
        RECT 58.645 176.715 58.975 176.730 ;
        RECT 60.485 176.715 60.815 177.045 ;
        RECT 68.305 177.030 68.635 177.045 ;
        RECT 78.170 177.030 78.550 177.040 ;
        RECT 68.305 176.730 78.550 177.030 ;
        RECT 68.305 176.715 68.635 176.730 ;
        RECT 78.170 176.720 78.550 176.730 ;
        RECT 12.580 176.350 16.580 176.500 ;
        RECT 60.500 176.365 60.800 176.715 ;
        RECT 19.545 176.350 19.875 176.365 ;
        RECT 12.580 176.050 19.875 176.350 ;
        RECT 12.580 175.900 16.580 176.050 ;
        RECT 19.545 176.035 19.875 176.050 ;
        RECT 40.705 176.350 41.035 176.365 ;
        RECT 47.145 176.350 47.475 176.365 ;
        RECT 40.705 176.050 47.475 176.350 ;
        RECT 40.705 176.035 41.035 176.050 ;
        RECT 47.145 176.035 47.475 176.050 ;
        RECT 47.810 176.350 48.190 176.360 ;
        RECT 54.045 176.350 54.375 176.365 ;
        RECT 47.810 176.050 54.375 176.350 ;
        RECT 47.810 176.040 48.190 176.050 ;
        RECT 54.045 176.035 54.375 176.050 ;
        RECT 58.645 176.360 58.975 176.365 ;
        RECT 58.645 176.350 59.230 176.360 ;
        RECT 58.645 176.050 59.430 176.350 ;
        RECT 58.645 176.040 59.230 176.050 ;
        RECT 58.645 176.035 58.975 176.040 ;
        RECT 60.485 176.035 60.815 176.365 ;
        RECT 67.845 176.350 68.175 176.365 ;
        RECT 69.685 176.360 70.015 176.365 ;
        RECT 68.970 176.350 69.350 176.360 ;
        RECT 67.845 176.050 69.350 176.350 ;
        RECT 67.845 176.035 68.175 176.050 ;
        RECT 68.970 176.040 69.350 176.050 ;
        RECT 69.685 176.350 70.270 176.360 ;
        RECT 87.165 176.350 87.495 176.365 ;
        RECT 90.930 176.350 94.930 176.500 ;
        RECT 69.685 176.050 70.470 176.350 ;
        RECT 87.165 176.050 94.930 176.350 ;
        RECT 69.685 176.040 70.270 176.050 ;
        RECT 69.685 176.035 70.015 176.040 ;
        RECT 87.165 176.035 87.495 176.050 ;
        RECT 90.930 175.900 94.930 176.050 ;
        RECT 32.170 175.670 32.550 175.680 ;
        RECT 43.210 175.670 43.590 175.680 ;
        RECT 50.365 175.670 50.695 175.685 ;
        RECT 32.170 175.370 42.860 175.670 ;
        RECT 32.170 175.360 32.550 175.370 ;
        RECT 42.560 174.990 42.860 175.370 ;
        RECT 43.210 175.370 50.695 175.670 ;
        RECT 43.210 175.360 43.590 175.370 ;
        RECT 50.365 175.355 50.695 175.370 ;
        RECT 53.125 175.670 53.455 175.685 ;
        RECT 57.930 175.670 58.310 175.680 ;
        RECT 53.125 175.370 58.310 175.670 ;
        RECT 53.125 175.355 53.455 175.370 ;
        RECT 57.930 175.360 58.310 175.370 ;
        RECT 59.565 175.670 59.895 175.685 ;
        RECT 77.965 175.670 78.295 175.685 ;
        RECT 59.565 175.370 78.295 175.670 ;
        RECT 59.565 175.355 59.895 175.370 ;
        RECT 77.965 175.355 78.295 175.370 ;
        RECT 50.825 174.990 51.155 175.005 ;
        RECT 78.885 174.990 79.215 175.005 ;
        RECT 42.560 174.690 51.155 174.990 ;
        RECT 50.825 174.675 51.155 174.690 ;
        RECT 65.330 174.690 79.215 174.990 ;
        RECT 33.630 174.335 35.210 174.665 ;
        RECT 39.530 174.310 39.910 174.320 ;
        RECT 61.865 174.310 62.195 174.325 ;
        RECT 39.530 174.010 62.195 174.310 ;
        RECT 39.530 174.000 39.910 174.010 ;
        RECT 61.865 173.995 62.195 174.010 ;
        RECT 30.330 173.630 30.710 173.640 ;
        RECT 49.445 173.630 49.775 173.645 ;
        RECT 64.625 173.630 64.955 173.645 ;
        RECT 30.330 173.330 64.955 173.630 ;
        RECT 30.330 173.320 30.710 173.330 ;
        RECT 49.445 173.315 49.775 173.330 ;
        RECT 64.625 173.315 64.955 173.330 ;
        RECT 18.370 172.950 18.750 172.960 ;
        RECT 53.585 172.950 53.915 172.965 ;
        RECT 57.265 172.960 57.595 172.965 ;
        RECT 18.370 172.650 53.915 172.950 ;
        RECT 18.370 172.640 18.750 172.650 ;
        RECT 53.585 172.635 53.915 172.650 ;
        RECT 57.010 172.950 57.595 172.960 ;
        RECT 58.185 172.950 58.515 172.965 ;
        RECT 63.245 172.960 63.575 172.965 ;
        RECT 60.690 172.950 61.070 172.960 ;
        RECT 57.010 172.650 57.820 172.950 ;
        RECT 58.185 172.650 61.070 172.950 ;
        RECT 57.010 172.640 57.595 172.650 ;
        RECT 57.265 172.635 57.595 172.640 ;
        RECT 58.185 172.635 58.515 172.650 ;
        RECT 60.690 172.640 61.070 172.650 ;
        RECT 63.245 172.950 63.830 172.960 ;
        RECT 63.245 172.650 64.030 172.950 ;
        RECT 63.245 172.640 63.830 172.650 ;
        RECT 63.245 172.635 63.575 172.640 ;
        RECT 48.525 172.280 48.855 172.285 ;
        RECT 51.285 172.280 51.615 172.285 ;
        RECT 56.345 172.280 56.675 172.285 ;
        RECT 48.525 172.270 49.110 172.280 ;
        RECT 51.285 172.270 51.870 172.280 ;
        RECT 56.090 172.270 56.675 172.280 ;
        RECT 48.300 171.970 49.110 172.270 ;
        RECT 51.060 171.970 51.870 172.270 ;
        RECT 55.890 171.970 56.675 172.270 ;
        RECT 48.525 171.960 49.110 171.970 ;
        RECT 51.285 171.960 51.870 171.970 ;
        RECT 56.090 171.960 56.675 171.970 ;
        RECT 48.525 171.955 48.855 171.960 ;
        RECT 51.285 171.955 51.615 171.960 ;
        RECT 56.345 171.955 56.675 171.960 ;
        RECT 60.025 172.270 60.355 172.285 ;
        RECT 65.330 172.270 65.630 174.690 ;
        RECT 78.885 174.675 79.215 174.690 ;
        RECT 83.025 174.310 83.355 174.325 ;
        RECT 74.530 174.010 83.355 174.310 ;
        RECT 66.465 172.950 66.795 172.965 ;
        RECT 67.130 172.950 67.510 172.960 ;
        RECT 74.530 172.950 74.830 174.010 ;
        RECT 83.025 173.995 83.355 174.010 ;
        RECT 78.425 173.630 78.755 173.645 ;
        RECT 82.105 173.630 82.435 173.645 ;
        RECT 82.770 173.630 83.150 173.640 ;
        RECT 78.425 173.330 83.150 173.630 ;
        RECT 78.425 173.315 78.755 173.330 ;
        RECT 82.105 173.315 82.435 173.330 ;
        RECT 82.770 173.320 83.150 173.330 ;
        RECT 66.465 172.650 67.510 172.950 ;
        RECT 66.465 172.635 66.795 172.650 ;
        RECT 67.130 172.640 67.510 172.650 ;
        RECT 69.010 172.650 74.830 172.950 ;
        RECT 87.165 172.950 87.495 172.965 ;
        RECT 90.930 172.950 94.930 173.100 ;
        RECT 87.165 172.650 94.930 172.950 ;
        RECT 60.025 171.970 65.630 172.270 ;
        RECT 66.210 172.270 66.590 172.280 ;
        RECT 67.845 172.270 68.175 172.285 ;
        RECT 66.210 171.970 68.175 172.270 ;
        RECT 60.025 171.955 60.355 171.970 ;
        RECT 66.210 171.960 66.590 171.970 ;
        RECT 67.845 171.955 68.175 171.970 ;
        RECT 36.930 171.615 38.510 171.945 ;
        RECT 45.050 171.590 45.430 171.600 ;
        RECT 47.145 171.590 47.475 171.605 ;
        RECT 50.825 171.600 51.155 171.605 ;
        RECT 45.050 171.290 47.475 171.590 ;
        RECT 45.050 171.280 45.430 171.290 ;
        RECT 47.145 171.275 47.475 171.290 ;
        RECT 50.570 171.590 51.155 171.600 ;
        RECT 51.745 171.590 52.075 171.605 ;
        RECT 53.585 171.590 53.915 171.605 ;
        RECT 50.570 171.290 51.380 171.590 ;
        RECT 51.745 171.290 53.915 171.590 ;
        RECT 50.570 171.280 51.155 171.290 ;
        RECT 50.825 171.275 51.155 171.280 ;
        RECT 51.745 171.275 52.075 171.290 ;
        RECT 53.585 171.275 53.915 171.290 ;
        RECT 65.290 171.590 65.670 171.600 ;
        RECT 66.925 171.590 67.255 171.605 ;
        RECT 65.290 171.290 67.255 171.590 ;
        RECT 65.290 171.280 65.670 171.290 ;
        RECT 66.925 171.275 67.255 171.290 ;
        RECT 32.425 170.910 32.755 170.925 ;
        RECT 39.325 170.910 39.655 170.925 ;
        RECT 32.425 170.610 39.655 170.910 ;
        RECT 32.425 170.595 32.755 170.610 ;
        RECT 39.325 170.595 39.655 170.610 ;
        RECT 46.685 170.910 47.015 170.925 ;
        RECT 51.745 170.910 52.075 170.925 ;
        RECT 46.685 170.610 52.075 170.910 ;
        RECT 46.685 170.595 47.015 170.610 ;
        RECT 51.745 170.595 52.075 170.610 ;
        RECT 62.325 170.910 62.655 170.925 ;
        RECT 65.085 170.910 65.415 170.925 ;
        RECT 69.010 170.910 69.310 172.650 ;
        RECT 87.165 172.635 87.495 172.650 ;
        RECT 90.930 172.500 94.930 172.650 ;
        RECT 70.145 172.270 70.475 172.285 ;
        RECT 71.730 172.270 72.110 172.280 ;
        RECT 70.145 171.970 72.110 172.270 ;
        RECT 70.145 171.955 70.475 171.970 ;
        RECT 71.730 171.960 72.110 171.970 ;
        RECT 70.810 171.590 71.190 171.600 ;
        RECT 85.325 171.590 85.655 171.605 ;
        RECT 70.810 171.290 85.655 171.590 ;
        RECT 70.810 171.280 71.190 171.290 ;
        RECT 85.325 171.275 85.655 171.290 ;
        RECT 62.325 170.610 69.310 170.910 ;
        RECT 71.985 170.910 72.315 170.925 ;
        RECT 79.345 170.910 79.675 170.925 ;
        RECT 71.985 170.610 79.675 170.910 ;
        RECT 62.325 170.595 62.655 170.610 ;
        RECT 65.085 170.595 65.415 170.610 ;
        RECT 71.985 170.595 72.315 170.610 ;
        RECT 79.345 170.595 79.675 170.610 ;
        RECT 20.465 170.230 20.795 170.245 ;
        RECT 77.045 170.230 77.375 170.245 ;
        RECT 20.465 169.930 77.375 170.230 ;
        RECT 20.465 169.915 20.795 169.930 ;
        RECT 77.045 169.915 77.375 169.930 ;
        RECT 47.145 169.550 47.475 169.565 ;
        RECT 54.965 169.550 55.295 169.565 ;
        RECT 47.145 169.250 55.295 169.550 ;
        RECT 47.145 169.235 47.475 169.250 ;
        RECT 54.965 169.235 55.295 169.250 ;
        RECT 65.545 169.550 65.875 169.565 ;
        RECT 69.225 169.550 69.555 169.565 ;
        RECT 65.545 169.250 69.555 169.550 ;
        RECT 65.545 169.235 65.875 169.250 ;
        RECT 69.225 169.235 69.555 169.250 ;
        RECT 77.965 169.550 78.295 169.565 ;
        RECT 90.930 169.550 94.930 169.700 ;
        RECT 77.965 169.250 94.930 169.550 ;
        RECT 77.965 169.235 78.295 169.250 ;
        RECT 33.630 168.895 35.210 169.225 ;
        RECT 90.930 169.100 94.930 169.250 ;
        RECT 62.785 168.870 63.115 168.885 ;
        RECT 76.585 168.870 76.915 168.885 ;
        RECT 62.785 168.570 76.915 168.870 ;
        RECT 62.785 168.555 63.115 168.570 ;
        RECT 76.585 168.555 76.915 168.570 ;
        RECT 31.045 168.190 31.375 168.205 ;
        RECT 42.545 168.190 42.875 168.205 ;
        RECT 31.045 167.890 42.875 168.190 ;
        RECT 31.045 167.875 31.375 167.890 ;
        RECT 42.545 167.875 42.875 167.890 ;
        RECT 66.925 168.190 67.255 168.205 ;
        RECT 79.345 168.190 79.675 168.205 ;
        RECT 66.925 167.890 79.675 168.190 ;
        RECT 66.925 167.875 67.255 167.890 ;
        RECT 79.345 167.875 79.675 167.890 ;
        RECT 37.485 167.510 37.815 167.525 ;
        RECT 38.865 167.510 39.195 167.525 ;
        RECT 47.145 167.510 47.475 167.525 ;
        RECT 37.485 167.210 47.475 167.510 ;
        RECT 37.485 167.195 37.815 167.210 ;
        RECT 38.865 167.195 39.195 167.210 ;
        RECT 47.145 167.195 47.475 167.210 ;
        RECT 36.930 166.175 38.510 166.505 ;
        RECT 83.945 166.150 84.275 166.165 ;
        RECT 90.930 166.150 94.930 166.300 ;
        RECT 83.945 165.850 94.930 166.150 ;
        RECT 83.945 165.835 84.275 165.850 ;
        RECT 90.930 165.700 94.930 165.850 ;
        RECT 27.365 165.470 27.695 165.485 ;
        RECT 32.425 165.470 32.755 165.485 ;
        RECT 71.065 165.470 71.395 165.485 ;
        RECT 75.205 165.470 75.535 165.485 ;
        RECT 27.365 165.170 75.535 165.470 ;
        RECT 27.365 165.155 27.695 165.170 ;
        RECT 32.425 165.155 32.755 165.170 ;
        RECT 71.065 165.155 71.395 165.170 ;
        RECT 75.205 165.155 75.535 165.170 ;
        RECT 71.985 164.790 72.315 164.805 ;
        RECT 73.570 164.790 73.950 164.800 ;
        RECT 71.985 164.490 73.950 164.790 ;
        RECT 71.985 164.475 72.315 164.490 ;
        RECT 73.570 164.480 73.950 164.490 ;
        RECT 33.630 163.455 35.210 163.785 ;
        RECT 75.410 162.750 75.790 162.760 ;
        RECT 76.125 162.750 76.455 162.765 ;
        RECT 75.410 162.450 76.455 162.750 ;
        RECT 75.410 162.440 75.790 162.450 ;
        RECT 76.125 162.435 76.455 162.450 ;
        RECT 84.405 162.750 84.735 162.765 ;
        RECT 90.930 162.750 94.930 162.900 ;
        RECT 84.405 162.450 94.930 162.750 ;
        RECT 84.405 162.435 84.735 162.450 ;
        RECT 90.930 162.300 94.930 162.450 ;
        RECT 77.045 162.080 77.375 162.085 ;
        RECT 77.045 162.070 77.630 162.080 ;
        RECT 76.820 161.770 77.630 162.070 ;
        RECT 77.045 161.760 77.630 161.770 ;
        RECT 77.045 161.755 77.375 161.760 ;
        RECT 36.930 160.735 38.510 161.065 ;
        RECT 48.065 160.030 48.395 160.045 ;
        RECT 49.905 160.030 50.235 160.045 ;
        RECT 48.065 159.730 50.235 160.030 ;
        RECT 48.065 159.715 48.395 159.730 ;
        RECT 49.905 159.715 50.235 159.730 ;
        RECT 12.580 159.350 16.580 159.500 ;
        RECT 20.005 159.350 20.335 159.365 ;
        RECT 12.580 159.050 20.335 159.350 ;
        RECT 12.580 158.900 16.580 159.050 ;
        RECT 20.005 159.035 20.335 159.050 ;
        RECT 43.465 159.350 43.795 159.365 ;
        RECT 48.065 159.350 48.395 159.365 ;
        RECT 43.465 159.050 48.395 159.350 ;
        RECT 43.465 159.035 43.795 159.050 ;
        RECT 48.065 159.035 48.395 159.050 ;
        RECT 80.265 159.350 80.595 159.365 ;
        RECT 90.930 159.350 94.930 159.500 ;
        RECT 80.265 159.050 94.930 159.350 ;
        RECT 80.265 159.035 80.595 159.050 ;
        RECT 90.930 158.900 94.930 159.050 ;
        RECT 33.630 158.015 35.210 158.345 ;
        RECT 47.145 157.990 47.475 158.005 ;
        RECT 49.905 157.990 50.235 158.005 ;
        RECT 47.145 157.690 50.235 157.990 ;
        RECT 47.145 157.675 47.475 157.690 ;
        RECT 49.905 157.675 50.235 157.690 ;
        RECT 12.580 155.950 16.580 156.100 ;
        RECT 21.845 155.950 22.175 155.965 ;
        RECT 12.580 155.650 22.175 155.950 ;
        RECT 12.580 155.500 16.580 155.650 ;
        RECT 21.845 155.635 22.175 155.650 ;
        RECT 85.785 155.950 86.115 155.965 ;
        RECT 90.930 155.950 94.930 156.100 ;
        RECT 85.785 155.650 94.930 155.950 ;
        RECT 85.785 155.635 86.115 155.650 ;
        RECT 36.930 155.295 38.510 155.625 ;
        RECT 90.930 155.500 94.930 155.650 ;
        RECT 19.545 153.230 19.875 153.245 ;
        RECT 16.570 152.930 19.875 153.230 ;
        RECT 16.570 152.700 16.870 152.930 ;
        RECT 19.545 152.915 19.875 152.930 ;
        RECT 12.580 152.250 16.870 152.700 ;
        RECT 33.630 152.575 35.210 152.905 ;
        RECT 82.565 152.550 82.895 152.565 ;
        RECT 90.930 152.550 94.930 152.700 ;
        RECT 82.565 152.250 94.930 152.550 ;
        RECT 12.580 152.100 16.580 152.250 ;
        RECT 82.565 152.235 82.895 152.250 ;
        RECT 90.930 152.100 94.930 152.250 ;
        RECT 40.705 151.190 41.035 151.205 ;
        RECT 81.645 151.190 81.975 151.205 ;
        RECT 40.705 150.890 81.975 151.190 ;
        RECT 40.705 150.875 41.035 150.890 ;
        RECT 81.645 150.875 81.975 150.890 ;
        RECT 36.930 149.855 38.510 150.185 ;
        RECT 12.580 149.150 16.580 149.300 ;
        RECT 87.625 149.150 87.955 149.165 ;
        RECT 90.930 149.150 94.930 149.300 ;
        RECT 12.580 148.700 16.870 149.150 ;
        RECT 87.625 148.850 94.930 149.150 ;
        RECT 87.625 148.835 87.955 148.850 ;
        RECT 90.930 148.700 94.930 148.850 ;
        RECT 16.570 148.470 16.870 148.700 ;
        RECT 20.005 148.470 20.335 148.485 ;
        RECT 16.570 148.170 20.335 148.470 ;
        RECT 20.005 148.155 20.335 148.170 ;
        RECT 33.630 147.135 35.210 147.465 ;
        RECT 87.165 145.750 87.495 145.765 ;
        RECT 90.930 145.750 94.930 145.900 ;
        RECT 87.165 145.450 94.930 145.750 ;
        RECT 87.165 145.435 87.495 145.450 ;
        RECT 90.930 145.300 94.930 145.450 ;
        RECT 36.930 144.415 38.510 144.745 ;
        RECT 87.625 142.350 87.955 142.365 ;
        RECT 90.930 142.350 94.930 142.500 ;
        RECT 87.625 142.050 94.930 142.350 ;
        RECT 87.625 142.035 87.955 142.050 ;
        RECT 33.630 141.695 35.210 142.025 ;
        RECT 90.930 141.900 94.930 142.050 ;
        RECT 36.930 138.975 38.510 139.305 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 31.275 220.235 31.605 220.565 ;
        RECT 18.395 216.155 18.725 216.485 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 16.555 187.595 16.885 187.925 ;
        RECT 16.570 186.565 16.870 187.595 ;
        RECT 16.555 186.235 16.885 186.565 ;
        RECT 18.410 172.965 18.710 216.155 ;
        RECT 26.675 214.115 27.005 214.445 ;
        RECT 22.995 211.395 23.325 211.725 ;
        RECT 23.010 183.165 23.310 211.395 ;
        RECT 24.410 207.570 25.590 208.750 ;
        RECT 24.410 200.770 25.590 201.950 ;
        RECT 24.835 198.475 25.165 198.805 ;
        RECT 22.995 182.835 23.325 183.165 ;
        RECT 24.850 182.485 25.150 198.475 ;
        RECT 25.755 194.395 26.085 194.725 ;
        RECT 25.770 185.205 26.070 194.395 ;
        RECT 25.755 184.875 26.085 185.205 ;
        RECT 26.690 183.845 26.990 214.115 ;
        RECT 27.595 205.275 27.925 205.605 ;
        RECT 26.675 183.515 27.005 183.845 ;
        RECT 27.610 182.485 27.910 205.275 ;
        RECT 28.515 200.515 28.845 200.845 ;
        RECT 28.530 191.325 28.830 200.515 ;
        RECT 30.355 199.155 30.685 199.485 ;
        RECT 30.370 191.750 30.670 199.155 ;
        RECT 31.290 194.725 31.590 220.235 ;
        RECT 42.315 213.435 42.645 213.765 ;
        RECT 32.195 198.475 32.525 198.805 ;
        RECT 31.275 194.395 31.605 194.725 ;
        RECT 28.515 190.995 28.845 191.325 ;
        RECT 29.930 190.570 31.110 191.750 ;
        RECT 28.515 189.635 28.845 189.965 ;
        RECT 29.435 189.635 29.765 189.965 ;
        RECT 24.835 182.155 25.165 182.485 ;
        RECT 27.595 182.155 27.925 182.485 ;
        RECT 28.530 181.125 28.830 189.635 ;
        RECT 28.515 180.795 28.845 181.125 ;
        RECT 29.450 180.445 29.750 189.635 ;
        RECT 29.435 180.115 29.765 180.445 ;
        RECT 30.370 173.645 30.670 190.570 ;
        RECT 31.275 188.275 31.605 188.605 ;
        RECT 31.290 183.165 31.590 188.275 ;
        RECT 31.275 182.835 31.605 183.165 ;
        RECT 32.210 175.685 32.510 198.475 ;
        RECT 32.195 175.355 32.525 175.685 ;
        RECT 30.355 173.315 30.685 173.645 ;
        RECT 18.395 172.635 18.725 172.965 ;
        RECT 33.620 138.900 35.220 210.100 ;
        RECT 35.875 204.595 36.205 204.925 ;
        RECT 35.890 184.525 36.190 204.595 ;
        RECT 35.875 184.195 36.205 184.525 ;
        RECT 35.875 182.155 36.205 182.485 ;
        RECT 35.890 180.445 36.190 182.155 ;
        RECT 35.875 180.115 36.205 180.445 ;
        RECT 36.920 138.900 38.520 210.100 ;
        RECT 39.555 204.595 39.885 204.925 ;
        RECT 39.570 174.325 39.870 204.595 ;
        RECT 41.395 202.555 41.725 202.885 ;
        RECT 40.475 201.195 40.805 201.525 ;
        RECT 40.490 197.445 40.790 201.195 ;
        RECT 40.475 197.115 40.805 197.445 ;
        RECT 40.475 195.755 40.805 196.085 ;
        RECT 40.490 191.325 40.790 195.755 ;
        RECT 40.475 190.995 40.805 191.325 ;
        RECT 40.490 179.085 40.790 190.995 ;
        RECT 40.475 178.755 40.805 179.085 ;
        RECT 41.410 178.405 41.710 202.555 ;
        RECT 42.330 195.405 42.630 213.435 ;
        RECT 58.875 212.075 59.205 212.405 ;
        RECT 45.075 211.395 45.405 211.725 ;
        RECT 56.115 211.395 56.445 211.725 ;
        RECT 44.155 201.875 44.485 202.205 ;
        RECT 43.235 197.115 43.565 197.445 ;
        RECT 42.315 195.075 42.645 195.405 ;
        RECT 42.315 194.395 42.645 194.725 ;
        RECT 42.330 185.205 42.630 194.395 ;
        RECT 42.315 184.875 42.645 185.205 ;
        RECT 41.395 178.075 41.725 178.405 ;
        RECT 43.250 175.685 43.550 197.115 ;
        RECT 44.170 188.605 44.470 201.875 ;
        RECT 44.155 188.275 44.485 188.605 ;
        RECT 45.090 183.165 45.390 211.395 ;
        RECT 46.915 205.955 47.245 206.285 ;
        RECT 45.995 199.835 46.325 200.165 ;
        RECT 46.010 183.165 46.310 199.835 ;
        RECT 46.930 187.925 47.230 205.955 ;
        RECT 54.275 204.595 54.605 204.925 ;
        RECT 52.435 201.875 52.765 202.205 ;
        RECT 47.835 193.715 48.165 194.045 ;
        RECT 46.915 187.595 47.245 187.925 ;
        RECT 45.075 182.835 45.405 183.165 ;
        RECT 45.995 182.835 46.325 183.165 ;
        RECT 43.235 175.355 43.565 175.685 ;
        RECT 39.555 173.995 39.885 174.325 ;
        RECT 45.090 171.605 45.390 182.835 ;
        RECT 47.850 176.365 48.150 193.715 ;
        RECT 51.515 186.235 51.845 186.565 ;
        RECT 48.755 185.555 49.085 185.885 ;
        RECT 47.835 176.035 48.165 176.365 ;
        RECT 48.770 172.285 49.070 185.555 ;
        RECT 50.595 176.715 50.925 177.045 ;
        RECT 48.755 171.955 49.085 172.285 ;
        RECT 50.610 171.605 50.910 176.715 ;
        RECT 51.530 172.285 51.830 186.235 ;
        RECT 52.450 180.445 52.750 201.875 ;
        RECT 53.355 187.595 53.685 187.925 ;
        RECT 52.435 180.115 52.765 180.445 ;
        RECT 53.370 177.045 53.670 187.595 ;
        RECT 54.290 181.805 54.590 204.595 ;
        RECT 55.195 199.835 55.525 200.165 ;
        RECT 55.210 189.285 55.510 199.835 ;
        RECT 55.195 188.955 55.525 189.285 ;
        RECT 54.275 181.475 54.605 181.805 ;
        RECT 55.210 177.725 55.510 188.955 ;
        RECT 56.130 183.845 56.430 211.395 ;
        RECT 57.035 207.315 57.365 207.645 ;
        RECT 57.050 202.885 57.350 207.315 ;
        RECT 57.035 202.555 57.365 202.885 ;
        RECT 57.050 186.565 57.350 202.555 ;
        RECT 57.955 188.275 58.285 188.605 ;
        RECT 57.035 186.235 57.365 186.565 ;
        RECT 56.115 183.515 56.445 183.845 ;
        RECT 55.195 177.395 55.525 177.725 ;
        RECT 57.035 177.395 57.365 177.725 ;
        RECT 53.355 176.715 53.685 177.045 ;
        RECT 56.115 176.715 56.445 177.045 ;
        RECT 56.130 172.285 56.430 176.715 ;
        RECT 57.050 172.965 57.350 177.395 ;
        RECT 57.970 175.685 58.270 188.275 ;
        RECT 58.890 176.365 59.190 212.075 ;
        RECT 79.115 209.355 79.445 209.685 ;
        RECT 77.275 206.635 77.605 206.965 ;
        RECT 69.915 204.595 70.245 204.925 ;
        RECT 71.755 204.595 72.085 204.925 ;
        RECT 68.995 203.235 69.325 203.565 ;
        RECT 59.795 202.555 60.125 202.885 ;
        RECT 59.810 194.725 60.110 202.555 ;
        RECT 65.315 201.195 65.645 201.525 ;
        RECT 60.715 199.155 61.045 199.485 ;
        RECT 59.795 194.395 60.125 194.725 ;
        RECT 59.810 179.085 60.110 194.395 ;
        RECT 59.795 178.755 60.125 179.085 ;
        RECT 58.875 176.035 59.205 176.365 ;
        RECT 57.955 175.355 58.285 175.685 ;
        RECT 60.730 172.965 61.030 199.155 ;
        RECT 63.475 181.475 63.805 181.805 ;
        RECT 63.490 172.965 63.790 181.475 ;
        RECT 57.035 172.635 57.365 172.965 ;
        RECT 60.715 172.635 61.045 172.965 ;
        RECT 63.475 172.635 63.805 172.965 ;
        RECT 51.515 171.955 51.845 172.285 ;
        RECT 56.115 171.955 56.445 172.285 ;
        RECT 65.330 171.605 65.630 201.195 ;
        RECT 67.155 197.115 67.485 197.445 ;
        RECT 66.235 196.435 66.565 196.765 ;
        RECT 66.250 172.285 66.550 196.435 ;
        RECT 67.170 182.485 67.470 197.115 ;
        RECT 67.155 182.155 67.485 182.485 ;
        RECT 67.155 178.075 67.485 178.405 ;
        RECT 67.170 172.965 67.470 178.075 ;
        RECT 69.010 176.365 69.310 203.235 ;
        RECT 69.930 176.365 70.230 204.595 ;
        RECT 71.770 191.750 72.070 204.595 ;
        RECT 73.170 200.770 74.350 201.950 ;
        RECT 71.330 190.570 72.510 191.750 ;
        RECT 71.755 181.475 72.085 181.805 ;
        RECT 70.835 177.395 71.165 177.725 ;
        RECT 68.995 176.035 69.325 176.365 ;
        RECT 69.915 176.035 70.245 176.365 ;
        RECT 67.155 172.635 67.485 172.965 ;
        RECT 66.235 171.955 66.565 172.285 ;
        RECT 70.850 171.605 71.150 177.395 ;
        RECT 71.770 172.285 72.070 181.475 ;
        RECT 71.755 171.955 72.085 172.285 ;
        RECT 45.075 171.275 45.405 171.605 ;
        RECT 50.595 171.275 50.925 171.605 ;
        RECT 65.315 171.275 65.645 171.605 ;
        RECT 70.835 171.275 71.165 171.605 ;
        RECT 73.610 164.805 73.910 200.770 ;
        RECT 75.435 199.835 75.765 200.165 ;
        RECT 75.450 189.285 75.750 199.835 ;
        RECT 75.435 188.955 75.765 189.285 ;
        RECT 75.435 182.155 75.765 182.485 ;
        RECT 73.595 164.475 73.925 164.805 ;
        RECT 75.450 162.765 75.750 182.155 ;
        RECT 75.435 162.435 75.765 162.765 ;
        RECT 77.290 162.085 77.590 206.635 ;
        RECT 78.195 203.235 78.525 203.565 ;
        RECT 78.210 177.045 78.510 203.235 ;
        RECT 79.130 191.325 79.430 209.355 ;
        RECT 85.130 207.570 86.310 208.750 ;
        RECT 82.795 199.155 83.125 199.485 ;
        RECT 79.115 190.995 79.445 191.325 ;
        RECT 78.195 176.715 78.525 177.045 ;
        RECT 82.810 173.645 83.110 199.155 ;
        RECT 82.795 173.315 83.125 173.645 ;
        RECT 77.275 161.755 77.605 162.085 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
      LAYER met5 ;
        RECT 24.200 207.360 86.520 208.960 ;
        RECT 24.200 200.560 74.560 202.160 ;
        RECT 29.720 190.360 72.720 191.960 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

