VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 16.075 211.425 16.245 211.615 ;
        RECT 18.375 211.425 18.545 211.615 ;
        RECT 18.835 211.425 19.005 211.615 ;
        RECT 22.055 211.425 22.225 211.615 ;
        RECT 23.895 211.425 24.065 211.615 ;
        RECT 24.355 211.445 24.525 211.615 ;
        RECT 24.360 211.425 24.525 211.445 ;
        RECT 28.490 211.425 28.660 211.615 ;
        RECT 31.250 211.425 31.420 211.615 ;
        RECT 31.715 211.445 31.885 211.615 ;
        RECT 31.745 211.425 31.885 211.445 ;
        RECT 34.475 211.425 34.645 211.615 ;
        RECT 37.670 211.425 37.840 211.615 ;
        RECT 42.305 211.470 42.465 211.580 ;
        RECT 51.955 211.425 52.125 211.615 ;
        RECT 52.420 211.425 52.590 211.615 ;
        RECT 57.930 211.425 58.100 211.615 ;
        RECT 67.135 211.425 67.305 211.615 ;
        RECT 69.435 211.425 69.605 211.615 ;
        RECT 69.895 211.425 70.065 211.615 ;
        RECT 79.095 211.425 79.265 211.615 ;
        RECT 80.935 211.445 81.105 211.615 ;
        RECT 80.935 211.425 81.135 211.445 ;
        RECT 85.525 211.425 85.695 211.615 ;
        RECT 86.915 211.425 87.085 211.615 ;
        RECT 15.935 210.615 17.305 211.425 ;
        RECT 17.325 210.515 18.675 211.425 ;
        RECT 18.695 210.745 20.525 211.425 ;
        RECT 19.180 210.515 20.525 210.745 ;
        RECT 20.535 210.745 22.365 211.425 ;
        RECT 22.375 210.745 24.205 211.425 ;
        RECT 24.360 210.745 26.195 211.425 ;
        RECT 20.535 210.515 21.880 210.745 ;
        RECT 22.375 210.515 23.720 210.745 ;
        RECT 25.265 210.515 26.195 210.745 ;
        RECT 26.615 210.515 28.805 211.425 ;
        RECT 28.825 210.555 29.255 211.340 ;
        RECT 29.375 210.515 31.565 211.425 ;
        RECT 31.745 210.605 34.315 211.425 ;
        RECT 34.335 210.745 37.545 211.425 ;
        RECT 32.725 210.515 34.315 210.605 ;
        RECT 36.410 210.515 37.545 210.745 ;
        RECT 37.610 210.515 41.685 211.425 ;
        RECT 41.705 210.555 42.135 211.340 ;
        RECT 43.160 210.745 52.265 211.425 ;
        RECT 52.275 210.745 54.550 211.425 ;
        RECT 53.180 210.515 54.550 210.745 ;
        RECT 54.585 210.555 55.015 211.340 ;
        RECT 55.325 210.515 58.245 211.425 ;
        RECT 58.340 210.745 67.445 211.425 ;
        RECT 67.465 210.555 67.895 211.340 ;
        RECT 67.915 210.515 69.730 211.425 ;
        RECT 69.755 210.745 78.860 211.425 ;
        RECT 78.965 210.515 80.315 211.425 ;
        RECT 80.345 210.555 80.775 211.340 ;
        RECT 80.935 210.745 84.465 211.425 ;
        RECT 81.640 210.515 84.465 210.745 ;
        RECT 84.475 210.645 85.845 211.425 ;
        RECT 85.855 210.615 87.225 211.425 ;
      LAYER nwell ;
        RECT 15.740 207.395 87.420 210.225 ;
      LAYER pwell ;
        RECT 18.435 207.015 19.385 207.105 ;
        RECT 15.935 206.195 17.305 207.005 ;
        RECT 18.435 206.195 20.365 207.015 ;
        RECT 20.535 206.875 21.880 207.105 ;
        RECT 23.515 207.015 24.465 207.105 ;
        RECT 20.535 206.195 22.365 206.875 ;
        RECT 22.535 206.195 24.465 207.015 ;
        RECT 26.960 206.905 28.345 207.105 ;
        RECT 24.675 206.225 28.345 206.905 ;
        RECT 28.825 206.280 29.255 207.065 ;
        RECT 16.075 205.985 16.245 206.195 ;
        RECT 20.215 206.175 20.365 206.195 ;
        RECT 17.465 206.040 17.625 206.150 ;
        RECT 18.835 205.985 19.005 206.175 ;
        RECT 19.290 205.985 19.460 206.175 ;
        RECT 20.215 206.005 20.385 206.175 ;
        RECT 20.670 205.985 20.840 206.175 ;
        RECT 22.055 206.005 22.225 206.195 ;
        RECT 22.535 206.175 22.685 206.195 ;
        RECT 22.515 206.005 22.685 206.175 ;
        RECT 23.890 205.985 24.060 206.175 ;
        RECT 24.815 206.005 24.985 206.225 ;
        RECT 26.975 206.195 28.345 206.225 ;
        RECT 29.735 206.195 33.405 207.105 ;
        RECT 33.415 206.875 35.005 207.105 ;
        RECT 33.415 206.195 37.085 206.875 ;
        RECT 37.180 206.195 46.285 206.875 ;
        RECT 46.295 206.195 50.395 207.105 ;
        RECT 50.435 206.195 54.105 207.105 ;
        RECT 54.585 206.280 55.015 207.065 ;
        RECT 58.455 206.875 62.385 207.105 ;
        RECT 72.440 206.875 75.265 207.105 ;
        RECT 76.120 206.875 78.945 207.105 ;
        RECT 55.035 206.195 57.775 206.875 ;
        RECT 57.970 206.195 62.385 206.875 ;
        RECT 62.395 206.195 71.500 206.875 ;
        RECT 71.735 206.195 75.265 206.875 ;
        RECT 75.415 206.195 78.945 206.875 ;
        RECT 78.965 206.195 80.315 207.105 ;
        RECT 80.345 206.280 80.775 207.065 ;
        RECT 81.640 206.875 84.465 207.105 ;
        RECT 80.935 206.195 84.465 206.875 ;
        RECT 84.475 206.195 85.845 206.975 ;
        RECT 85.855 206.195 87.225 207.005 ;
        RECT 15.935 205.175 17.305 205.985 ;
        RECT 17.315 205.305 19.145 205.985 ;
        RECT 17.315 205.075 18.660 205.305 ;
        RECT 19.175 205.075 20.525 205.985 ;
        RECT 20.555 205.075 21.905 205.985 ;
        RECT 22.370 205.755 24.060 205.985 ;
        RECT 24.215 205.955 25.610 205.985 ;
        RECT 26.655 205.955 26.825 206.175 ;
        RECT 27.115 206.005 27.285 206.175 ;
        RECT 28.490 206.035 28.610 206.145 ;
        RECT 29.410 206.035 29.530 206.145 ;
        RECT 29.880 206.005 30.050 206.195 ;
        RECT 27.145 205.985 27.285 206.005 ;
        RECT 32.175 205.985 32.345 206.175 ;
        RECT 36.770 206.005 36.940 206.195 ;
        RECT 41.375 205.985 41.545 206.175 ;
        RECT 42.305 206.030 42.465 206.140 ;
        RECT 43.215 205.985 43.385 206.175 ;
        RECT 45.975 206.005 46.145 206.195 ;
        RECT 46.440 206.005 46.610 206.195 ;
        RECT 53.790 206.005 53.960 206.195 ;
        RECT 54.250 206.035 54.370 206.145 ;
        RECT 55.175 206.005 55.345 206.195 ;
        RECT 57.970 206.175 58.080 206.195 ;
        RECT 62.535 206.175 62.705 206.195 ;
        RECT 71.735 206.175 71.935 206.195 ;
        RECT 75.415 206.175 75.615 206.195 ;
        RECT 57.910 206.005 58.080 206.175 ;
        RECT 61.155 205.985 61.325 206.175 ;
        RECT 62.530 206.005 62.705 206.175 ;
        RECT 62.530 205.985 62.700 206.005 ;
        RECT 63.000 205.985 63.170 206.175 ;
        RECT 66.685 206.030 66.845 206.140 ;
        RECT 71.275 206.005 71.445 206.175 ;
        RECT 71.245 205.985 71.445 206.005 ;
        RECT 71.735 205.985 71.905 206.175 ;
        RECT 75.415 206.005 75.585 206.175 ;
        RECT 80.015 206.005 80.185 206.195 ;
        RECT 80.935 206.175 81.135 206.195 ;
        RECT 80.935 206.005 81.105 206.175 ;
        RECT 81.855 205.985 82.025 206.175 ;
        RECT 85.070 205.985 85.240 206.175 ;
        RECT 85.535 206.145 85.705 206.195 ;
        RECT 85.530 206.035 85.705 206.145 ;
        RECT 85.535 206.005 85.705 206.035 ;
        RECT 86.915 205.985 87.085 206.195 ;
        RECT 22.370 205.075 24.205 205.755 ;
        RECT 24.215 205.275 26.950 205.955 ;
        RECT 24.215 205.075 25.625 205.275 ;
        RECT 27.145 205.165 29.715 205.985 ;
        RECT 29.745 205.305 32.485 205.985 ;
        RECT 32.580 205.305 41.685 205.985 ;
        RECT 28.125 205.075 29.715 205.165 ;
        RECT 41.705 205.115 42.135 205.900 ;
        RECT 43.075 205.305 52.180 205.985 ;
        RECT 52.360 205.305 61.465 205.985 ;
        RECT 61.495 205.075 62.845 205.985 ;
        RECT 62.855 205.075 66.455 205.985 ;
        RECT 67.465 205.115 67.895 205.900 ;
        RECT 67.915 205.305 71.445 205.985 ;
        RECT 67.915 205.075 70.740 205.305 ;
        RECT 71.605 205.075 72.955 205.985 ;
        RECT 73.060 205.305 82.165 205.985 ;
        RECT 82.175 205.075 85.385 205.985 ;
        RECT 85.855 205.175 87.225 205.985 ;
      LAYER nwell ;
        RECT 15.740 201.955 87.420 204.785 ;
      LAYER pwell ;
        RECT 15.935 200.755 17.305 201.565 ;
        RECT 18.720 201.435 20.065 201.665 ;
        RECT 18.235 200.755 20.065 201.435 ;
        RECT 20.075 201.435 21.420 201.665 ;
        RECT 20.075 200.755 21.905 201.435 ;
        RECT 22.855 200.755 24.205 201.665 ;
        RECT 25.355 201.575 26.305 201.665 ;
        RECT 24.375 200.755 26.305 201.575 ;
        RECT 26.515 200.755 28.805 201.665 ;
        RECT 28.825 200.840 29.255 201.625 ;
        RECT 29.275 200.755 30.645 201.535 ;
        RECT 30.665 200.755 33.395 201.665 ;
        RECT 33.415 200.755 36.155 201.435 ;
        RECT 36.260 200.755 45.365 201.435 ;
        RECT 45.460 200.755 54.565 201.435 ;
        RECT 54.585 200.840 55.015 201.625 ;
        RECT 55.035 200.755 59.165 201.665 ;
        RECT 59.195 200.755 60.545 201.665 ;
        RECT 60.555 200.755 69.660 201.435 ;
        RECT 69.755 200.755 78.860 201.435 ;
        RECT 78.955 200.755 80.325 201.535 ;
        RECT 80.345 200.840 80.775 201.625 ;
        RECT 80.805 200.985 84.005 201.665 ;
        RECT 84.500 201.435 85.845 201.665 ;
        RECT 80.805 200.755 83.860 200.985 ;
        RECT 84.015 200.755 85.845 201.435 ;
        RECT 85.855 200.755 87.225 201.565 ;
        RECT 16.075 200.545 16.245 200.755 ;
        RECT 17.465 200.600 17.625 200.710 ;
        RECT 18.375 200.565 18.545 200.755 ;
        RECT 18.835 200.545 19.005 200.735 ;
        RECT 19.290 200.595 19.410 200.705 ;
        RECT 20.215 200.585 20.385 200.735 ;
        RECT 15.935 199.735 17.305 200.545 ;
        RECT 17.315 199.865 19.145 200.545 ;
        RECT 17.315 199.635 18.660 199.865 ;
        RECT 19.615 199.635 20.505 200.585 ;
        RECT 20.685 200.545 20.855 200.735 ;
        RECT 21.595 200.565 21.765 200.755 ;
        RECT 22.060 200.545 22.230 200.735 ;
        RECT 22.970 200.565 23.140 200.755 ;
        RECT 24.375 200.735 24.525 200.755 ;
        RECT 24.355 200.565 24.525 200.735 ;
        RECT 25.735 200.545 25.905 200.735 ;
        RECT 28.490 200.565 28.660 200.755 ;
        RECT 30.335 200.565 30.505 200.755 ;
        RECT 30.335 200.545 30.500 200.565 ;
        RECT 30.795 200.545 30.965 200.735 ;
        RECT 33.095 200.565 33.265 200.755 ;
        RECT 33.555 200.565 33.725 200.755 ;
        RECT 36.775 200.545 36.945 200.735 ;
        RECT 38.160 200.545 38.330 200.735 ;
        RECT 38.620 200.545 38.790 200.735 ;
        RECT 20.535 199.765 21.905 200.545 ;
        RECT 21.915 199.635 25.585 200.545 ;
        RECT 25.595 199.635 28.345 200.545 ;
        RECT 28.665 199.865 30.500 200.545 ;
        RECT 28.665 199.635 29.595 199.865 ;
        RECT 30.655 199.635 33.865 200.545 ;
        RECT 33.875 199.635 37.085 200.545 ;
        RECT 37.095 199.635 38.445 200.545 ;
        RECT 38.475 199.635 41.395 200.545 ;
        RECT 41.705 199.675 42.135 200.460 ;
        RECT 42.300 200.315 42.470 200.735 ;
        RECT 45.055 200.565 45.225 200.755 ;
        RECT 46.900 200.545 47.070 200.735 ;
        RECT 50.575 200.545 50.745 200.735 ;
        RECT 54.255 200.565 54.425 200.755 ;
        RECT 58.850 200.565 59.020 200.755 ;
        RECT 60.230 200.565 60.400 200.755 ;
        RECT 60.695 200.565 60.865 200.755 ;
        RECT 63.450 200.545 63.620 200.735 ;
        RECT 63.920 200.565 64.090 200.735 ;
        RECT 67.130 200.595 67.250 200.705 ;
        RECT 63.945 200.545 64.090 200.565 ;
        RECT 68.055 200.545 68.225 200.735 ;
        RECT 69.895 200.565 70.065 200.755 ;
        RECT 77.260 200.545 77.430 200.735 ;
        RECT 79.095 200.565 79.265 200.755 ;
        RECT 80.940 200.545 81.110 200.735 ;
        RECT 83.690 200.565 83.860 200.755 ;
        RECT 84.155 200.565 84.325 200.755 ;
        RECT 85.525 200.545 85.695 200.735 ;
        RECT 86.915 200.545 87.085 200.755 ;
        RECT 43.580 200.315 46.740 200.545 ;
        RECT 42.195 199.865 46.740 200.315 ;
        RECT 42.195 199.635 43.570 199.865 ;
        RECT 45.360 199.635 46.740 199.865 ;
        RECT 46.755 199.635 50.410 200.545 ;
        RECT 50.435 199.865 59.540 200.545 ;
        RECT 59.635 199.635 63.765 200.545 ;
        RECT 63.945 199.635 66.985 200.545 ;
        RECT 67.465 199.675 67.895 200.460 ;
        RECT 67.915 199.865 77.020 200.545 ;
        RECT 77.115 199.635 80.660 200.545 ;
        RECT 80.795 199.635 84.340 200.545 ;
        RECT 84.475 199.765 85.845 200.545 ;
        RECT 85.855 199.735 87.225 200.545 ;
      LAYER nwell ;
        RECT 15.740 196.515 87.420 199.345 ;
      LAYER pwell ;
        RECT 17.785 196.135 19.375 196.225 ;
        RECT 15.935 195.315 17.305 196.125 ;
        RECT 17.785 195.315 20.355 196.135 ;
        RECT 21.585 195.995 22.515 196.225 ;
        RECT 16.075 195.105 16.245 195.315 ;
        RECT 20.215 195.295 20.355 195.315 ;
        RECT 20.680 195.315 22.515 195.995 ;
        RECT 22.835 195.315 26.505 196.225 ;
        RECT 27.435 195.315 28.805 196.095 ;
        RECT 28.825 195.400 29.255 196.185 ;
        RECT 29.275 195.315 30.625 196.225 ;
        RECT 30.655 195.315 32.485 196.225 ;
        RECT 32.645 195.315 36.300 196.225 ;
        RECT 37.095 195.315 40.305 196.225 ;
        RECT 40.400 195.315 49.505 195.995 ;
        RECT 49.515 195.315 53.645 196.225 ;
        RECT 54.585 195.400 55.015 196.185 ;
        RECT 55.120 195.315 64.225 195.995 ;
        RECT 64.235 195.315 67.445 196.225 ;
        RECT 67.455 195.315 71.125 196.225 ;
        RECT 71.220 195.315 80.325 195.995 ;
        RECT 80.345 195.400 80.775 196.185 ;
        RECT 81.640 195.995 84.465 196.225 ;
        RECT 80.935 195.315 84.465 195.995 ;
        RECT 84.485 195.315 85.835 196.225 ;
        RECT 85.855 195.315 87.225 196.125 ;
        RECT 20.680 195.295 20.845 195.315 ;
        RECT 17.450 195.155 17.570 195.265 ;
        RECT 18.835 195.105 19.005 195.295 ;
        RECT 19.305 195.105 19.475 195.295 ;
        RECT 20.215 195.125 20.385 195.295 ;
        RECT 20.675 195.125 20.845 195.295 ;
        RECT 21.595 195.105 21.765 195.295 ;
        RECT 22.975 195.105 23.145 195.295 ;
        RECT 23.430 195.155 23.550 195.265 ;
        RECT 23.895 195.105 24.065 195.295 ;
        RECT 26.190 195.125 26.360 195.315 ;
        RECT 26.665 195.160 26.825 195.270 ;
        RECT 28.495 195.125 28.665 195.315 ;
        RECT 28.950 195.155 29.070 195.265 ;
        RECT 28.495 195.105 28.660 195.125 ;
        RECT 29.425 195.105 29.595 195.295 ;
        RECT 30.340 195.125 30.510 195.315 ;
        RECT 30.800 195.125 30.970 195.315 ;
        RECT 32.645 195.295 32.805 195.315 ;
        RECT 32.175 195.105 32.345 195.295 ;
        RECT 32.635 195.125 32.805 195.295 ;
        RECT 35.395 195.125 35.565 195.295 ;
        RECT 35.395 195.105 35.545 195.125 ;
        RECT 35.855 195.105 36.025 195.295 ;
        RECT 36.770 195.155 36.890 195.265 ;
        RECT 37.235 195.125 37.405 195.315 ;
        RECT 41.370 195.105 41.540 195.295 ;
        RECT 45.055 195.105 45.225 195.295 ;
        RECT 45.515 195.105 45.685 195.295 ;
        RECT 49.195 195.125 49.365 195.315 ;
        RECT 49.660 195.125 49.830 195.315 ;
        RECT 53.805 195.160 53.965 195.270 ;
        RECT 57.475 195.105 57.645 195.295 ;
        RECT 57.930 195.155 58.050 195.265 ;
        RECT 63.915 195.125 64.085 195.315 ;
        RECT 67.130 195.295 67.300 195.315 ;
        RECT 67.130 195.125 67.305 195.295 ;
        RECT 67.600 195.125 67.770 195.315 ;
        RECT 67.135 195.105 67.305 195.125 ;
        RECT 68.055 195.105 68.225 195.295 ;
        RECT 71.270 195.155 71.390 195.265 ;
        RECT 71.740 195.105 71.910 195.295 ;
        RECT 75.885 195.150 76.045 195.260 ;
        RECT 80.015 195.125 80.185 195.315 ;
        RECT 80.935 195.295 81.135 195.315 ;
        RECT 80.935 195.125 81.105 195.295 ;
        RECT 84.615 195.125 84.785 195.315 ;
        RECT 85.535 195.105 85.705 195.295 ;
        RECT 86.915 195.105 87.085 195.315 ;
        RECT 15.935 194.295 17.305 195.105 ;
        RECT 17.315 194.425 19.145 195.105 ;
        RECT 17.315 194.195 18.660 194.425 ;
        RECT 19.155 194.325 20.525 195.105 ;
        RECT 20.535 194.325 21.905 195.105 ;
        RECT 21.925 194.195 23.275 195.105 ;
        RECT 23.765 194.195 26.495 195.105 ;
        RECT 26.825 194.425 28.660 195.105 ;
        RECT 26.825 194.195 27.755 194.425 ;
        RECT 29.275 194.325 30.645 195.105 ;
        RECT 30.655 194.195 32.470 195.105 ;
        RECT 33.615 194.285 35.545 195.105 ;
        RECT 35.715 194.425 38.465 195.105 ;
        RECT 33.615 194.195 34.565 194.285 ;
        RECT 37.535 194.195 38.465 194.425 ;
        RECT 38.475 194.195 41.685 195.105 ;
        RECT 41.705 194.235 42.135 195.020 ;
        RECT 42.155 194.195 45.365 195.105 ;
        RECT 45.375 194.195 48.585 195.105 ;
        RECT 48.680 194.425 57.785 195.105 ;
        RECT 58.340 194.425 67.445 195.105 ;
        RECT 67.915 195.075 69.755 195.105 ;
        RECT 67.465 194.235 67.895 195.020 ;
        RECT 67.915 194.425 71.080 195.075 ;
        RECT 68.400 194.395 71.080 194.425 ;
        RECT 68.400 194.195 69.755 194.395 ;
        RECT 71.595 194.195 75.725 195.105 ;
        RECT 76.740 194.425 85.845 195.105 ;
        RECT 85.855 194.295 87.225 195.105 ;
      LAYER nwell ;
        RECT 15.740 191.075 87.420 193.905 ;
      LAYER pwell ;
        RECT 15.935 189.875 17.305 190.685 ;
        RECT 18.235 189.875 19.605 190.655 ;
        RECT 19.615 189.875 20.985 190.655 ;
        RECT 20.995 189.875 22.365 190.655 ;
        RECT 24.805 190.555 25.735 190.785 ;
        RECT 23.900 189.875 25.735 190.555 ;
        RECT 26.055 190.555 27.400 190.785 ;
        RECT 26.055 189.875 27.885 190.555 ;
        RECT 28.825 189.960 29.255 190.745 ;
        RECT 30.195 190.555 31.125 190.785 ;
        RECT 30.195 189.875 34.095 190.555 ;
        RECT 34.795 189.875 36.165 190.655 ;
        RECT 36.175 189.875 37.990 190.785 ;
        RECT 38.100 189.875 47.205 190.555 ;
        RECT 47.215 189.875 50.870 190.785 ;
        RECT 50.895 189.875 54.565 190.785 ;
        RECT 54.585 189.960 55.015 190.745 ;
        RECT 55.045 189.875 57.785 190.555 ;
        RECT 57.795 189.875 61.870 190.785 ;
        RECT 61.935 189.875 71.040 190.555 ;
        RECT 71.220 189.875 80.325 190.555 ;
        RECT 80.345 189.960 80.775 190.745 ;
        RECT 80.795 189.875 83.835 190.785 ;
        RECT 84.015 189.875 85.845 190.785 ;
        RECT 85.855 189.875 87.225 190.685 ;
        RECT 16.075 189.665 16.245 189.875 ;
        RECT 19.295 189.855 19.465 189.875 ;
        RECT 17.465 189.720 17.625 189.830 ;
        RECT 18.835 189.665 19.005 189.855 ;
        RECT 19.290 189.685 19.465 189.855 ;
        RECT 20.675 189.685 20.845 189.875 ;
        RECT 22.055 189.685 22.225 189.875 ;
        RECT 23.900 189.855 24.065 189.875 ;
        RECT 22.515 189.685 22.685 189.855 ;
        RECT 19.290 189.665 19.460 189.685 ;
        RECT 23.435 189.665 23.605 189.855 ;
        RECT 23.895 189.685 24.065 189.855 ;
        RECT 24.820 189.665 24.990 189.855 ;
        RECT 27.575 189.685 27.745 189.875 ;
        RECT 28.045 189.720 28.205 189.830 ;
        RECT 28.500 189.665 28.670 189.855 ;
        RECT 29.425 189.720 29.585 189.830 ;
        RECT 29.875 189.665 30.045 189.855 ;
        RECT 30.610 189.685 30.780 189.875 ;
        RECT 31.530 189.665 31.700 189.855 ;
        RECT 34.470 189.715 34.590 189.825 ;
        RECT 34.935 189.685 35.105 189.875 ;
        RECT 35.670 189.665 35.840 189.855 ;
        RECT 37.695 189.685 37.865 189.875 ;
        RECT 39.530 189.715 39.650 189.825 ;
        RECT 39.995 189.665 40.165 189.855 ;
        RECT 42.300 189.665 42.470 189.855 ;
        RECT 46.895 189.685 47.065 189.875 ;
        RECT 47.360 189.685 47.530 189.875 ;
        RECT 47.820 189.665 47.990 189.855 ;
        RECT 48.250 189.665 48.420 189.855 ;
        RECT 54.250 189.685 54.420 189.875 ;
        RECT 55.180 189.665 55.350 189.855 ;
        RECT 57.475 189.685 57.645 189.875 ;
        RECT 57.935 189.665 58.105 189.855 ;
        RECT 61.640 189.685 61.810 189.875 ;
        RECT 62.075 189.685 62.245 189.875 ;
        RECT 67.135 189.665 67.305 189.855 ;
        RECT 68.045 189.665 68.215 189.855 ;
        RECT 74.495 189.685 74.665 189.855 ;
        RECT 80.015 189.685 80.185 189.875 ;
        RECT 83.690 189.855 83.835 189.875 ;
        RECT 85.530 189.855 85.700 189.875 ;
        RECT 83.690 189.685 83.865 189.855 ;
        RECT 85.530 189.685 85.705 189.855 ;
        RECT 74.495 189.665 74.635 189.685 ;
        RECT 83.695 189.665 83.865 189.685 ;
        RECT 85.535 189.665 85.705 189.685 ;
        RECT 86.915 189.665 87.085 189.875 ;
        RECT 15.935 188.855 17.305 189.665 ;
        RECT 17.315 188.985 19.145 189.665 ;
        RECT 17.315 188.755 18.660 188.985 ;
        RECT 19.175 188.755 20.525 189.665 ;
        RECT 20.665 188.755 23.665 189.665 ;
        RECT 24.675 188.985 28.345 189.665 ;
        RECT 24.675 188.755 25.600 188.985 ;
        RECT 28.355 188.755 29.705 189.665 ;
        RECT 29.745 188.755 31.095 189.665 ;
        RECT 31.115 188.985 35.015 189.665 ;
        RECT 35.255 188.985 39.155 189.665 ;
        RECT 39.855 188.985 41.685 189.665 ;
        RECT 31.115 188.755 32.045 188.985 ;
        RECT 35.255 188.755 36.185 188.985 ;
        RECT 40.340 188.755 41.685 188.985 ;
        RECT 41.705 188.795 42.135 189.580 ;
        RECT 42.155 188.755 46.455 189.665 ;
        RECT 46.755 188.755 48.105 189.665 ;
        RECT 48.190 188.755 52.265 189.665 ;
        RECT 52.275 188.755 55.475 189.665 ;
        RECT 55.505 188.985 58.245 189.665 ;
        RECT 58.340 188.985 67.445 189.665 ;
        RECT 67.465 188.795 67.895 189.580 ;
        RECT 67.915 188.985 72.045 189.665 ;
        RECT 67.915 188.755 69.285 188.985 ;
        RECT 72.065 188.845 74.635 189.665 ;
        RECT 74.900 188.985 84.005 189.665 ;
        RECT 84.015 188.985 85.845 189.665 ;
        RECT 85.855 188.855 87.225 189.665 ;
        RECT 72.065 188.755 73.655 188.845 ;
      LAYER nwell ;
        RECT 15.740 185.635 87.420 188.465 ;
      LAYER pwell ;
        RECT 15.935 184.435 17.305 185.245 ;
        RECT 17.315 184.435 18.685 185.215 ;
        RECT 19.175 184.435 20.525 185.345 ;
        RECT 20.665 184.435 23.665 185.345 ;
        RECT 24.215 185.115 25.140 185.345 ;
        RECT 24.215 184.435 27.885 185.115 ;
        RECT 28.825 184.520 29.255 185.305 ;
        RECT 29.275 184.435 30.645 185.215 ;
        RECT 30.655 185.115 31.585 185.345 ;
        RECT 30.655 184.435 34.555 185.115 ;
        RECT 34.795 184.435 36.165 185.215 ;
        RECT 36.635 184.435 38.005 185.215 ;
        RECT 38.945 184.435 41.675 185.345 ;
        RECT 42.155 184.435 46.230 185.345 ;
        RECT 47.215 184.435 50.425 185.345 ;
        RECT 50.435 184.435 52.250 185.345 ;
        RECT 52.375 184.435 54.565 185.345 ;
        RECT 54.585 184.520 55.015 185.305 ;
        RECT 55.120 184.435 64.225 185.115 ;
        RECT 64.245 184.435 66.985 185.115 ;
        RECT 66.995 184.435 76.100 185.115 ;
        RECT 76.195 184.435 79.850 185.345 ;
        RECT 80.345 184.520 80.775 185.305 ;
        RECT 80.795 184.665 83.995 185.345 ;
        RECT 80.940 184.435 83.995 184.665 ;
        RECT 84.015 184.435 85.365 185.345 ;
        RECT 85.855 184.435 87.225 185.245 ;
        RECT 16.075 184.225 16.245 184.435 ;
        RECT 17.465 184.245 17.635 184.435 ;
        RECT 19.290 184.415 19.460 184.435 ;
        RECT 18.830 184.275 18.950 184.385 ;
        RECT 19.290 184.245 19.465 184.415 ;
        RECT 19.295 184.225 19.465 184.245 ;
        RECT 20.665 184.225 20.835 184.415 ;
        RECT 21.135 184.225 21.305 184.415 ;
        RECT 22.980 184.225 23.150 184.415 ;
        RECT 23.435 184.245 23.605 184.435 ;
        RECT 23.890 184.275 24.010 184.385 ;
        RECT 24.360 184.245 24.530 184.435 ;
        RECT 25.265 184.225 25.435 184.415 ;
        RECT 25.745 184.225 25.915 184.415 ;
        RECT 27.125 184.225 27.295 184.415 ;
        RECT 28.045 184.280 28.205 184.390 ;
        RECT 28.495 184.225 28.665 184.415 ;
        RECT 30.325 184.245 30.495 184.435 ;
        RECT 30.785 184.225 30.955 184.415 ;
        RECT 31.070 184.245 31.240 184.435 ;
        RECT 31.265 184.270 31.425 184.380 ;
        RECT 32.170 184.225 32.340 184.415 ;
        RECT 33.555 184.225 33.725 184.415 ;
        RECT 34.935 184.245 35.105 184.435 ;
        RECT 36.310 184.275 36.430 184.385 ;
        RECT 37.685 184.245 37.855 184.435 ;
        RECT 38.165 184.280 38.325 184.390 ;
        RECT 39.075 184.225 39.245 184.415 ;
        RECT 41.375 184.245 41.545 184.435 ;
        RECT 46.000 184.415 46.170 184.435 ;
        RECT 47.355 184.415 47.525 184.435 ;
        RECT 41.830 184.275 41.950 184.385 ;
        RECT 44.595 184.225 44.765 184.415 ;
        RECT 45.965 184.245 46.170 184.415 ;
        RECT 46.445 184.280 46.605 184.390 ;
        RECT 47.345 184.245 47.525 184.415 ;
        RECT 45.965 184.225 46.135 184.245 ;
        RECT 47.345 184.225 47.515 184.245 ;
        RECT 47.825 184.225 47.995 184.415 ;
        RECT 50.105 184.225 50.275 184.415 ;
        RECT 51.485 184.225 51.655 184.415 ;
        RECT 51.955 184.225 52.125 184.435 ;
        RECT 54.250 184.245 54.420 184.435 ;
        RECT 58.855 184.245 59.025 184.415 ;
        RECT 58.855 184.225 59.015 184.245 ;
        RECT 62.075 184.225 62.245 184.415 ;
        RECT 62.545 184.270 62.705 184.380 ;
        RECT 63.915 184.245 64.085 184.435 ;
        RECT 66.675 184.245 66.845 184.435 ;
        RECT 67.135 184.385 67.305 184.435 ;
        RECT 67.130 184.275 67.305 184.385 ;
        RECT 67.135 184.245 67.305 184.275 ;
        RECT 66.645 184.225 66.845 184.245 ;
        RECT 74.030 184.225 74.200 184.415 ;
        RECT 74.500 184.225 74.670 184.415 ;
        RECT 76.340 184.245 76.510 184.435 ;
        RECT 80.010 184.275 80.130 184.385 ;
        RECT 80.940 184.245 81.110 184.435 ;
        RECT 84.160 184.245 84.330 184.435 ;
        RECT 85.535 184.385 85.705 184.415 ;
        RECT 85.530 184.275 85.705 184.385 ;
        RECT 85.535 184.225 85.705 184.275 ;
        RECT 86.915 184.225 87.085 184.435 ;
        RECT 15.935 183.415 17.305 184.225 ;
        RECT 18.235 183.445 19.605 184.225 ;
        RECT 19.615 183.445 20.985 184.225 ;
        RECT 20.995 183.545 22.825 184.225 ;
        RECT 22.835 183.315 24.185 184.225 ;
        RECT 24.215 183.445 25.585 184.225 ;
        RECT 25.595 183.445 26.965 184.225 ;
        RECT 26.975 183.445 28.345 184.225 ;
        RECT 28.365 183.315 29.715 184.225 ;
        RECT 29.735 183.445 31.105 184.225 ;
        RECT 32.055 183.315 33.405 184.225 ;
        RECT 33.415 183.415 38.925 184.225 ;
        RECT 38.935 183.415 41.685 184.225 ;
        RECT 41.705 183.355 42.135 184.140 ;
        RECT 42.185 183.315 44.905 184.225 ;
        RECT 44.915 183.445 46.285 184.225 ;
        RECT 46.295 183.445 47.665 184.225 ;
        RECT 47.675 183.445 49.045 184.225 ;
        RECT 49.055 183.445 50.425 184.225 ;
        RECT 50.435 183.445 51.805 184.225 ;
        RECT 51.815 183.315 55.025 184.225 ;
        RECT 55.360 183.315 59.015 184.225 ;
        RECT 59.175 183.315 62.385 184.225 ;
        RECT 63.315 183.545 66.845 184.225 ;
        RECT 63.315 183.315 66.140 183.545 ;
        RECT 67.465 183.355 67.895 184.140 ;
        RECT 68.275 183.315 74.345 184.225 ;
        RECT 74.500 183.995 76.190 184.225 ;
        RECT 74.355 183.315 76.190 183.995 ;
        RECT 76.740 183.545 85.845 184.225 ;
        RECT 85.855 183.415 87.225 184.225 ;
      LAYER nwell ;
        RECT 15.740 180.195 87.420 183.025 ;
      LAYER pwell ;
        RECT 15.935 178.995 17.305 179.805 ;
        RECT 19.285 179.675 20.215 179.905 ;
        RECT 18.380 178.995 20.215 179.675 ;
        RECT 20.535 179.675 21.900 179.905 ;
        RECT 25.575 179.675 26.505 179.905 ;
        RECT 20.535 178.995 23.745 179.675 ;
        RECT 23.755 178.995 26.505 179.675 ;
        RECT 26.975 178.995 28.790 179.905 ;
        RECT 28.825 179.080 29.255 179.865 ;
        RECT 30.195 178.995 33.115 179.905 ;
        RECT 33.415 178.995 35.245 179.905 ;
        RECT 35.270 178.995 38.925 179.905 ;
        RECT 38.935 178.995 42.605 179.905 ;
        RECT 42.615 179.675 43.535 179.905 ;
        RECT 42.615 178.995 46.200 179.675 ;
        RECT 46.755 178.995 48.585 179.905 ;
        RECT 48.595 179.675 49.525 179.905 ;
        RECT 53.175 179.675 54.105 179.905 ;
        RECT 48.595 178.995 51.345 179.675 ;
        RECT 51.355 178.995 54.105 179.675 ;
        RECT 54.585 179.080 55.015 179.865 ;
        RECT 55.035 178.995 58.245 179.905 ;
        RECT 59.175 178.995 61.925 179.905 ;
        RECT 62.420 179.675 63.765 179.905 ;
        RECT 61.935 178.995 63.765 179.675 ;
        RECT 63.775 178.995 67.250 179.905 ;
        RECT 67.465 178.995 68.815 179.905 ;
        RECT 68.835 178.995 77.940 179.675 ;
        RECT 78.035 178.995 80.245 179.905 ;
        RECT 80.345 179.080 80.775 179.865 ;
        RECT 80.795 178.995 84.005 179.905 ;
        RECT 84.500 179.675 85.845 179.905 ;
        RECT 84.015 178.995 85.845 179.675 ;
        RECT 85.855 178.995 87.225 179.805 ;
        RECT 16.075 178.785 16.245 178.995 ;
        RECT 18.380 178.975 18.545 178.995 ;
        RECT 23.430 178.975 23.600 178.995 ;
        RECT 17.465 178.785 17.635 178.975 ;
        RECT 18.375 178.805 18.545 178.975 ;
        RECT 18.845 178.830 19.005 178.940 ;
        RECT 19.760 178.785 19.930 178.975 ;
        RECT 23.430 178.805 23.605 178.975 ;
        RECT 23.895 178.805 24.065 178.995 ;
        RECT 23.435 178.785 23.605 178.805 ;
        RECT 24.815 178.785 24.985 178.975 ;
        RECT 25.275 178.785 25.445 178.975 ;
        RECT 26.655 178.945 26.825 178.975 ;
        RECT 26.650 178.835 26.825 178.945 ;
        RECT 26.655 178.785 26.825 178.835 ;
        RECT 28.495 178.805 28.665 178.995 ;
        RECT 29.425 178.840 29.585 178.950 ;
        RECT 30.340 178.805 30.510 178.995 ;
        RECT 31.250 178.785 31.420 178.975 ;
        RECT 32.635 178.785 32.805 178.975 ;
        RECT 33.560 178.805 33.730 178.995 ;
        RECT 38.155 178.785 38.325 178.975 ;
        RECT 38.610 178.805 38.780 178.995 ;
        RECT 39.080 178.805 39.250 178.995 ;
        RECT 42.295 178.785 42.465 178.975 ;
        RECT 42.760 178.805 42.930 178.995 ;
        RECT 45.515 178.785 45.685 178.975 ;
        RECT 46.430 178.835 46.550 178.945 ;
        RECT 47.350 178.835 47.470 178.945 ;
        RECT 48.270 178.805 48.440 178.995 ;
        RECT 48.740 178.785 48.910 178.975 ;
        RECT 50.115 178.785 50.285 178.975 ;
        RECT 51.035 178.805 51.205 178.995 ;
        RECT 51.495 178.975 51.665 178.995 ;
        RECT 51.485 178.805 51.665 178.975 ;
        RECT 51.485 178.785 51.655 178.805 ;
        RECT 52.880 178.785 53.050 178.975 ;
        RECT 54.245 178.785 54.415 178.975 ;
        RECT 55.175 178.805 55.345 178.995 ;
        RECT 57.935 178.805 58.105 178.975 ;
        RECT 58.405 178.840 58.565 178.950 ;
        RECT 57.905 178.785 58.105 178.805 ;
        RECT 59.320 178.785 59.490 178.995 ;
        RECT 59.780 178.785 59.950 178.975 ;
        RECT 62.075 178.805 62.245 178.995 ;
        RECT 62.530 178.835 62.650 178.945 ;
        RECT 63.000 178.785 63.170 178.975 ;
        RECT 63.920 178.805 64.090 178.995 ;
        RECT 66.685 178.830 66.845 178.940 ;
        RECT 67.595 178.805 67.765 178.995 ;
        RECT 68.975 178.805 69.145 178.995 ;
        RECT 70.815 178.785 70.985 178.975 ;
        RECT 71.270 178.835 71.390 178.945 ;
        RECT 71.740 178.785 71.910 178.975 ;
        RECT 74.965 178.830 75.125 178.940 ;
        RECT 75.875 178.785 76.045 178.975 ;
        RECT 78.180 178.805 78.350 178.995 ;
        RECT 80.940 178.805 81.110 178.995 ;
        RECT 84.155 178.805 84.325 178.995 ;
        RECT 85.085 178.830 85.245 178.940 ;
        RECT 86.915 178.785 87.085 178.995 ;
        RECT 15.935 177.975 17.305 178.785 ;
        RECT 17.315 178.005 18.685 178.785 ;
        RECT 19.760 178.555 21.450 178.785 ;
        RECT 19.615 177.875 21.450 178.555 ;
        RECT 21.915 178.105 23.745 178.785 ;
        RECT 21.915 177.875 23.260 178.105 ;
        RECT 23.755 178.005 25.125 178.785 ;
        RECT 25.135 178.005 26.505 178.785 ;
        RECT 26.515 177.975 30.185 178.785 ;
        RECT 31.135 177.875 32.485 178.785 ;
        RECT 32.495 177.975 38.005 178.785 ;
        RECT 38.015 177.975 41.685 178.785 ;
        RECT 41.705 177.915 42.135 178.700 ;
        RECT 42.155 178.105 45.365 178.785 ;
        RECT 44.230 177.875 45.365 178.105 ;
        RECT 45.390 177.875 47.205 178.785 ;
        RECT 47.675 177.875 49.025 178.785 ;
        RECT 49.055 178.005 50.425 178.785 ;
        RECT 50.435 178.005 51.805 178.785 ;
        RECT 51.815 177.875 53.165 178.785 ;
        RECT 53.195 178.005 54.565 178.785 ;
        RECT 54.575 178.105 58.105 178.785 ;
        RECT 54.575 177.875 57.400 178.105 ;
        RECT 58.255 177.875 59.605 178.785 ;
        RECT 59.635 177.875 62.385 178.785 ;
        RECT 62.855 178.105 66.440 178.785 ;
        RECT 62.855 177.875 63.775 178.105 ;
        RECT 67.465 177.915 67.895 178.700 ;
        RECT 67.915 177.875 71.125 178.785 ;
        RECT 71.740 178.555 74.795 178.785 ;
        RECT 71.595 177.875 74.795 178.555 ;
        RECT 75.735 178.105 84.840 178.785 ;
        RECT 85.855 177.975 87.225 178.785 ;
      LAYER nwell ;
        RECT 15.740 174.755 87.420 177.585 ;
      LAYER pwell ;
        RECT 15.935 173.555 17.305 174.365 ;
        RECT 18.235 173.555 21.445 174.465 ;
        RECT 21.455 173.555 26.965 174.365 ;
        RECT 26.975 173.555 28.805 174.365 ;
        RECT 28.825 173.640 29.255 174.425 ;
        RECT 29.285 173.555 32.015 174.465 ;
        RECT 32.035 173.555 35.705 174.365 ;
        RECT 36.175 173.555 37.525 174.465 ;
        RECT 37.555 173.555 43.065 174.365 ;
        RECT 43.075 173.555 48.585 174.365 ;
        RECT 49.530 173.555 51.345 174.465 ;
        RECT 52.290 173.555 54.105 174.465 ;
        RECT 54.585 173.640 55.015 174.425 ;
        RECT 55.495 173.555 56.865 174.335 ;
        RECT 56.885 173.555 58.235 174.465 ;
        RECT 58.275 173.555 59.625 174.465 ;
        RECT 59.635 173.555 62.845 174.465 ;
        RECT 63.315 173.555 64.685 174.335 ;
        RECT 64.715 173.555 66.065 174.465 ;
        RECT 66.085 173.555 67.435 174.465 ;
        RECT 67.555 173.555 69.745 174.465 ;
        RECT 70.020 173.555 72.955 174.465 ;
        RECT 72.985 173.555 75.920 174.465 ;
        RECT 76.665 173.785 79.865 174.465 ;
        RECT 76.665 173.555 79.720 173.785 ;
        RECT 80.345 173.640 80.775 174.425 ;
        RECT 80.805 173.785 84.005 174.465 ;
        RECT 84.500 174.235 85.845 174.465 ;
        RECT 80.805 173.555 83.860 173.785 ;
        RECT 84.015 173.555 85.845 174.235 ;
        RECT 85.855 173.555 87.225 174.365 ;
        RECT 16.075 173.345 16.245 173.555 ;
        RECT 17.455 173.345 17.625 173.535 ;
        RECT 18.375 173.365 18.545 173.555 ;
        RECT 19.290 173.395 19.410 173.505 ;
        RECT 20.030 173.345 20.200 173.535 ;
        RECT 21.595 173.365 21.765 173.555 ;
        RECT 23.895 173.345 24.065 173.535 ;
        RECT 27.115 173.365 27.285 173.555 ;
        RECT 28.035 173.345 28.205 173.535 ;
        RECT 30.335 173.365 30.505 173.535 ;
        RECT 31.715 173.365 31.885 173.555 ;
        RECT 32.175 173.365 32.345 173.555 ;
        RECT 30.335 173.345 30.500 173.365 ;
        RECT 33.555 173.345 33.725 173.535 ;
        RECT 34.025 173.390 34.185 173.500 ;
        RECT 35.210 173.345 35.380 173.535 ;
        RECT 35.850 173.395 35.970 173.505 ;
        RECT 37.240 173.365 37.410 173.555 ;
        RECT 37.695 173.365 37.865 173.555 ;
        RECT 39.075 173.345 39.245 173.535 ;
        RECT 43.215 173.365 43.385 173.555 ;
        RECT 43.675 173.345 43.845 173.535 ;
        RECT 44.130 173.395 44.250 173.505 ;
        RECT 44.595 173.345 44.765 173.535 ;
        RECT 47.355 173.345 47.525 173.535 ;
        RECT 48.745 173.400 48.905 173.510 ;
        RECT 49.655 173.365 49.825 173.555 ;
        RECT 50.115 173.345 50.285 173.535 ;
        RECT 51.505 173.400 51.665 173.510 ;
        RECT 51.965 173.390 52.125 173.500 ;
        RECT 52.415 173.365 52.585 173.555 ;
        RECT 52.875 173.345 53.045 173.535 ;
        RECT 54.250 173.395 54.370 173.505 ;
        RECT 54.725 173.390 54.885 173.500 ;
        RECT 55.170 173.395 55.290 173.505 ;
        RECT 56.545 173.345 56.715 173.555 ;
        RECT 57.015 173.365 57.185 173.555 ;
        RECT 58.390 173.365 58.560 173.555 ;
        RECT 60.235 173.365 60.405 173.535 ;
        RECT 60.205 173.345 60.405 173.365 ;
        RECT 60.695 173.345 60.865 173.535 ;
        RECT 62.535 173.365 62.705 173.555 ;
        RECT 62.995 173.505 63.165 173.535 ;
        RECT 62.990 173.395 63.165 173.505 ;
        RECT 62.995 173.345 63.165 173.395 ;
        RECT 63.465 173.345 63.635 173.535 ;
        RECT 64.365 173.365 64.535 173.555 ;
        RECT 65.750 173.535 65.920 173.555 ;
        RECT 65.745 173.365 65.920 173.535 ;
        RECT 65.745 173.345 65.915 173.365 ;
        RECT 66.215 173.345 66.385 173.555 ;
        RECT 68.050 173.395 68.170 173.505 ;
        RECT 68.525 173.345 68.695 173.535 ;
        RECT 69.430 173.365 69.600 173.555 ;
        RECT 70.020 173.535 70.065 173.555 ;
        RECT 75.875 173.535 75.920 173.555 ;
        RECT 69.895 173.365 70.065 173.535 ;
        RECT 70.815 173.345 70.985 173.535 ;
        RECT 74.495 173.345 74.665 173.535 ;
        RECT 74.955 173.345 75.125 173.535 ;
        RECT 75.875 173.365 76.045 173.535 ;
        RECT 76.330 173.395 76.450 173.505 ;
        RECT 76.795 173.345 76.965 173.535 ;
        RECT 79.550 173.365 79.720 173.555 ;
        RECT 80.010 173.395 80.130 173.505 ;
        RECT 83.690 173.365 83.860 173.555 ;
        RECT 84.155 173.365 84.325 173.555 ;
        RECT 86.915 173.345 87.085 173.555 ;
        RECT 15.935 172.535 17.305 173.345 ;
        RECT 17.315 172.535 19.145 173.345 ;
        RECT 19.615 172.665 23.515 173.345 ;
        RECT 19.615 172.435 20.545 172.665 ;
        RECT 23.755 172.535 26.505 173.345 ;
        RECT 26.515 172.435 28.330 173.345 ;
        RECT 28.665 172.665 30.500 173.345 ;
        RECT 28.665 172.435 29.595 172.665 ;
        RECT 30.655 172.435 33.865 173.345 ;
        RECT 34.795 172.665 38.695 173.345 ;
        RECT 34.795 172.435 35.725 172.665 ;
        RECT 38.935 172.535 41.685 173.345 ;
        RECT 41.705 172.475 42.135 173.260 ;
        RECT 42.155 172.435 43.970 173.345 ;
        RECT 44.465 172.435 47.195 173.345 ;
        RECT 47.215 172.535 49.965 173.345 ;
        RECT 49.990 172.435 51.805 173.345 ;
        RECT 52.750 172.435 54.565 173.345 ;
        RECT 55.495 172.565 56.865 173.345 ;
        RECT 56.875 172.665 60.405 173.345 ;
        RECT 56.875 172.435 59.700 172.665 ;
        RECT 60.555 172.565 61.925 173.345 ;
        RECT 61.935 172.565 63.305 173.345 ;
        RECT 63.315 172.565 64.685 173.345 ;
        RECT 64.695 172.565 66.065 173.345 ;
        RECT 66.075 172.565 67.445 173.345 ;
        RECT 67.465 172.475 67.895 173.260 ;
        RECT 68.375 172.565 69.745 173.345 ;
        RECT 69.765 172.435 71.115 173.345 ;
        RECT 71.275 172.435 74.725 173.345 ;
        RECT 74.815 172.665 76.645 173.345 ;
        RECT 76.655 172.665 85.760 173.345 ;
        RECT 75.300 172.435 76.645 172.665 ;
        RECT 85.855 172.535 87.225 173.345 ;
      LAYER nwell ;
        RECT 15.740 169.315 87.420 172.145 ;
      LAYER pwell ;
        RECT 15.935 168.115 17.305 168.925 ;
        RECT 17.315 168.115 19.145 168.925 ;
        RECT 19.155 168.795 20.085 169.025 ;
        RECT 19.155 168.115 23.055 168.795 ;
        RECT 23.295 168.115 26.045 168.925 ;
        RECT 26.055 168.115 27.870 169.025 ;
        RECT 28.825 168.200 29.255 168.985 ;
        RECT 29.585 168.795 30.515 169.025 ;
        RECT 29.585 168.115 31.420 168.795 ;
        RECT 31.575 168.115 33.390 169.025 ;
        RECT 34.335 168.795 35.265 169.025 ;
        RECT 34.335 168.115 38.235 168.795 ;
        RECT 38.485 168.115 39.835 169.025 ;
        RECT 39.855 168.115 41.205 169.025 ;
        RECT 42.155 168.115 43.970 169.025 ;
        RECT 44.005 168.115 45.355 169.025 ;
        RECT 45.375 168.115 46.745 168.925 ;
        RECT 46.755 168.115 48.105 169.025 ;
        RECT 48.135 168.115 53.645 168.925 ;
        RECT 54.585 168.200 55.015 168.985 ;
        RECT 55.035 168.825 55.980 169.025 ;
        RECT 57.315 168.825 58.245 169.025 ;
        RECT 55.035 168.345 58.245 168.825 ;
        RECT 55.035 168.145 58.105 168.345 ;
        RECT 55.035 168.115 55.980 168.145 ;
        RECT 16.075 167.905 16.245 168.115 ;
        RECT 17.455 167.905 17.625 168.115 ;
        RECT 19.570 167.925 19.740 168.115 ;
        RECT 23.435 167.925 23.605 168.115 ;
        RECT 23.620 167.905 23.790 168.095 ;
        RECT 27.115 167.905 27.285 168.095 ;
        RECT 27.575 167.905 27.745 168.115 ;
        RECT 31.255 168.095 31.420 168.115 ;
        RECT 28.045 167.960 28.205 168.070 ;
        RECT 31.255 167.925 31.425 168.095 ;
        RECT 33.095 167.905 33.265 168.115 ;
        RECT 33.565 167.960 33.725 168.070 ;
        RECT 34.750 167.925 34.920 168.115 ;
        RECT 38.615 167.905 38.785 168.115 ;
        RECT 40.920 167.925 41.090 168.115 ;
        RECT 41.385 168.065 41.545 168.070 ;
        RECT 41.370 167.960 41.545 168.065 ;
        RECT 41.370 167.955 41.490 167.960 ;
        RECT 42.295 167.905 42.465 168.095 ;
        RECT 43.675 167.925 43.845 168.115 ;
        RECT 44.135 167.925 44.305 168.115 ;
        RECT 45.515 168.095 45.685 168.115 ;
        RECT 45.050 167.955 45.170 168.065 ;
        RECT 45.515 167.925 45.690 168.095 ;
        RECT 47.820 167.925 47.990 168.115 ;
        RECT 48.275 167.925 48.445 168.115 ;
        RECT 45.520 167.905 45.690 167.925 ;
        RECT 49.195 167.905 49.365 168.095 ;
        RECT 51.040 167.905 51.210 168.095 ;
        RECT 53.805 167.960 53.965 168.070 ;
        RECT 57.470 167.905 57.640 168.095 ;
        RECT 57.935 167.925 58.105 168.145 ;
        RECT 58.255 168.115 60.085 168.925 ;
        RECT 60.555 168.115 63.765 169.025 ;
        RECT 63.790 168.115 67.445 169.025 ;
        RECT 67.455 168.115 69.270 169.025 ;
        RECT 70.345 168.115 73.345 169.025 ;
        RECT 75.260 168.795 76.630 169.025 ;
        RECT 74.355 168.115 76.630 168.795 ;
        RECT 76.665 168.115 79.405 168.795 ;
        RECT 80.345 168.200 80.775 168.985 ;
        RECT 80.875 168.115 83.085 169.025 ;
        RECT 83.095 168.115 85.835 168.795 ;
        RECT 85.855 168.115 87.225 168.925 ;
        RECT 58.395 167.925 58.565 168.115 ;
        RECT 60.230 167.955 60.350 168.065 ;
        RECT 60.685 167.925 60.855 168.115 ;
        RECT 57.940 167.905 58.105 167.925 ;
        RECT 61.160 167.905 61.330 168.095 ;
        RECT 61.615 167.905 61.785 168.095 ;
        RECT 64.375 167.905 64.545 168.095 ;
        RECT 66.225 167.905 66.395 168.095 ;
        RECT 67.130 167.925 67.300 168.115 ;
        RECT 68.065 167.950 68.225 168.060 ;
        RECT 68.975 167.905 69.145 168.115 ;
        RECT 69.445 167.960 69.605 168.070 ;
        RECT 70.355 167.905 70.525 168.095 ;
        RECT 71.735 167.905 71.905 168.095 ;
        RECT 73.115 167.925 73.285 168.115 ;
        RECT 73.585 167.960 73.745 168.070 ;
        RECT 74.500 167.925 74.670 168.115 ;
        RECT 15.935 167.095 17.305 167.905 ;
        RECT 17.315 167.095 20.065 167.905 ;
        RECT 20.305 167.225 24.205 167.905 ;
        RECT 23.275 166.995 24.205 167.225 ;
        RECT 24.215 166.995 27.425 167.905 ;
        RECT 27.435 167.095 32.945 167.905 ;
        RECT 32.955 167.095 38.465 167.905 ;
        RECT 38.475 167.095 41.225 167.905 ;
        RECT 41.705 167.035 42.135 167.820 ;
        RECT 42.155 167.095 44.905 167.905 ;
        RECT 45.375 167.225 49.045 167.905 ;
        RECT 45.375 166.995 46.300 167.225 ;
        RECT 49.055 167.095 50.885 167.905 ;
        RECT 50.895 166.995 53.815 167.905 ;
        RECT 54.310 166.995 57.785 167.905 ;
        RECT 57.940 167.225 59.775 167.905 ;
        RECT 58.845 166.995 59.775 167.225 ;
        RECT 60.095 166.995 61.445 167.905 ;
        RECT 61.475 167.095 64.225 167.905 ;
        RECT 64.250 166.995 66.065 167.905 ;
        RECT 66.075 167.125 67.445 167.905 ;
        RECT 67.465 167.035 67.895 167.820 ;
        RECT 68.835 167.125 70.205 167.905 ;
        RECT 70.215 167.125 71.585 167.905 ;
        RECT 71.675 166.995 75.125 167.905 ;
        RECT 75.410 167.875 75.580 168.095 ;
        RECT 77.725 167.950 77.885 168.060 ;
        RECT 78.635 167.905 78.805 168.095 ;
        RECT 79.095 167.925 79.265 168.115 ;
        RECT 79.565 167.960 79.725 168.070 ;
        RECT 82.770 167.925 82.940 168.115 ;
        RECT 83.235 167.925 83.405 168.115 ;
        RECT 76.610 167.875 77.565 167.905 ;
        RECT 75.285 167.195 77.565 167.875 ;
        RECT 78.495 167.225 81.245 167.905 ;
        RECT 76.610 166.995 77.565 167.195 ;
        RECT 80.315 166.995 81.245 167.225 ;
        RECT 81.255 167.875 82.650 167.905 ;
        RECT 83.695 167.875 83.865 168.095 ;
        RECT 84.155 167.905 84.325 168.095 ;
        RECT 86.915 167.905 87.085 168.115 ;
        RECT 81.255 167.195 83.990 167.875 ;
        RECT 84.015 167.225 85.845 167.905 ;
        RECT 81.255 166.995 82.665 167.195 ;
        RECT 84.500 166.995 85.845 167.225 ;
        RECT 85.855 167.095 87.225 167.905 ;
      LAYER nwell ;
        RECT 15.740 163.875 87.420 166.705 ;
      LAYER pwell ;
        RECT 15.935 162.675 17.305 163.485 ;
        RECT 17.315 162.675 20.065 163.485 ;
        RECT 23.275 163.355 24.205 163.585 ;
        RECT 20.305 162.675 24.205 163.355 ;
        RECT 24.215 162.675 26.965 163.485 ;
        RECT 27.435 162.675 28.785 163.585 ;
        RECT 28.825 162.760 29.255 163.545 ;
        RECT 29.275 162.675 32.485 163.585 ;
        RECT 32.955 163.355 33.885 163.585 ;
        RECT 32.955 162.675 36.855 163.355 ;
        RECT 37.095 162.675 38.445 163.585 ;
        RECT 38.475 162.675 41.225 163.485 ;
        RECT 41.235 162.675 44.445 163.585 ;
        RECT 44.455 162.675 49.965 163.485 ;
        RECT 49.975 162.675 53.645 163.485 ;
        RECT 54.585 162.760 55.015 163.545 ;
        RECT 55.035 163.385 55.980 163.585 ;
        RECT 57.315 163.385 58.245 163.585 ;
        RECT 55.035 162.905 58.245 163.385 ;
        RECT 55.035 162.705 58.105 162.905 ;
        RECT 55.035 162.675 55.980 162.705 ;
        RECT 16.075 162.465 16.245 162.675 ;
        RECT 17.455 162.485 17.625 162.675 ;
        RECT 18.835 162.465 19.005 162.655 ;
        RECT 19.295 162.465 19.465 162.655 ;
        RECT 22.055 162.465 22.225 162.655 ;
        RECT 22.515 162.465 22.685 162.655 ;
        RECT 23.620 162.485 23.790 162.675 ;
        RECT 24.355 162.485 24.525 162.675 ;
        RECT 27.110 162.515 27.230 162.625 ;
        RECT 28.030 162.515 28.150 162.625 ;
        RECT 28.500 162.485 28.670 162.675 ;
        RECT 29.415 162.465 29.585 162.655 ;
        RECT 29.875 162.485 30.045 162.655 ;
        RECT 32.175 162.485 32.345 162.675 ;
        RECT 32.630 162.515 32.750 162.625 ;
        RECT 29.905 162.465 30.045 162.485 ;
        RECT 32.910 162.465 33.080 162.655 ;
        RECT 33.370 162.485 33.540 162.675 ;
        RECT 36.775 162.465 36.945 162.655 ;
        RECT 38.160 162.485 38.330 162.675 ;
        RECT 38.615 162.485 38.785 162.675 ;
        RECT 40.925 162.510 41.085 162.620 ;
        RECT 41.365 162.485 41.535 162.675 ;
        RECT 44.595 162.485 44.765 162.675 ;
        RECT 45.975 162.485 46.145 162.655 ;
        RECT 38.620 162.465 38.785 162.485 ;
        RECT 45.975 162.465 46.135 162.485 ;
        RECT 49.650 162.465 49.820 162.655 ;
        RECT 50.115 162.465 50.285 162.675 ;
        RECT 53.335 162.465 53.505 162.655 ;
        RECT 53.805 162.520 53.965 162.630 ;
        RECT 57.935 162.485 58.105 162.705 ;
        RECT 58.255 162.675 63.765 163.485 ;
        RECT 63.775 162.675 67.445 163.485 ;
        RECT 67.455 162.675 68.825 163.485 ;
        RECT 58.395 162.485 58.565 162.675 ;
        RECT 58.860 162.465 59.030 162.655 ;
        RECT 63.915 162.485 64.085 162.675 ;
        RECT 65.755 162.465 65.925 162.655 ;
        RECT 66.215 162.465 66.385 162.655 ;
        RECT 67.595 162.485 67.765 162.675 ;
        RECT 68.055 162.465 68.225 162.655 ;
        RECT 68.835 162.635 69.725 163.585 ;
        RECT 71.125 163.355 72.045 163.585 ;
        RECT 69.755 162.675 72.045 163.355 ;
        RECT 72.075 162.675 73.425 163.585 ;
        RECT 73.895 162.675 75.265 163.455 ;
        RECT 76.610 163.385 77.565 163.585 ;
        RECT 75.285 162.705 77.565 163.385 ;
        RECT 69.435 162.485 69.605 162.635 ;
        RECT 69.895 162.485 70.065 162.675 ;
        RECT 71.275 162.465 71.445 162.655 ;
        RECT 73.110 162.485 73.280 162.675 ;
        RECT 73.575 162.625 73.745 162.655 ;
        RECT 73.570 162.515 73.745 162.625 ;
        RECT 73.575 162.465 73.745 162.515 ;
        RECT 74.045 162.485 74.215 162.675 ;
        RECT 75.410 162.485 75.580 162.705 ;
        RECT 76.610 162.675 77.565 162.705 ;
        RECT 78.115 162.675 80.325 163.585 ;
        RECT 80.345 162.760 80.775 163.545 ;
        RECT 80.805 162.675 82.155 163.585 ;
        RECT 82.255 162.675 85.840 163.585 ;
        RECT 85.855 162.675 87.225 163.485 ;
        RECT 75.885 162.510 76.045 162.620 ;
        RECT 76.795 162.465 76.965 162.655 ;
        RECT 77.710 162.515 77.830 162.625 ;
        RECT 80.010 162.485 80.180 162.675 ;
        RECT 80.935 162.485 81.105 162.675 ;
        RECT 85.530 162.485 85.700 162.675 ;
        RECT 86.915 162.465 87.085 162.675 ;
        RECT 15.935 161.655 17.305 162.465 ;
        RECT 17.315 161.785 19.145 162.465 ;
        RECT 19.155 161.785 20.985 162.465 ;
        RECT 17.315 161.555 18.660 161.785 ;
        RECT 20.995 161.685 22.365 162.465 ;
        RECT 22.375 161.655 27.885 162.465 ;
        RECT 28.365 161.555 29.715 162.465 ;
        RECT 29.905 161.645 32.475 162.465 ;
        RECT 30.885 161.555 32.475 161.645 ;
        RECT 32.495 161.785 36.395 162.465 ;
        RECT 32.495 161.555 33.425 161.785 ;
        RECT 36.635 161.655 38.465 162.465 ;
        RECT 38.620 161.785 40.455 162.465 ;
        RECT 39.525 161.555 40.455 161.785 ;
        RECT 41.705 161.595 42.135 162.380 ;
        RECT 42.480 161.555 46.135 162.465 ;
        RECT 46.295 161.555 49.965 162.465 ;
        RECT 49.975 161.555 53.185 162.465 ;
        RECT 53.195 161.655 58.705 162.465 ;
        RECT 58.715 161.555 63.105 162.465 ;
        RECT 63.325 161.555 66.055 162.465 ;
        RECT 66.075 161.655 67.445 162.465 ;
        RECT 67.465 161.595 67.895 162.380 ;
        RECT 67.915 161.555 71.125 162.465 ;
        RECT 71.135 161.785 73.425 162.465 ;
        RECT 73.435 161.785 75.725 162.465 ;
        RECT 76.655 161.785 85.760 162.465 ;
        RECT 72.505 161.555 73.425 161.785 ;
        RECT 74.805 161.555 75.725 161.785 ;
        RECT 85.855 161.655 87.225 162.465 ;
      LAYER nwell ;
        RECT 15.740 158.435 87.420 161.265 ;
      LAYER pwell ;
        RECT 15.935 157.235 17.305 158.045 ;
        RECT 18.235 157.235 20.065 158.145 ;
        RECT 21.920 157.915 23.285 158.145 ;
        RECT 20.075 157.235 23.285 157.915 ;
        RECT 23.295 157.235 25.125 158.145 ;
        RECT 25.135 157.235 28.805 158.045 ;
        RECT 28.825 157.320 29.255 158.105 ;
        RECT 29.275 157.915 30.620 158.145 ;
        RECT 36.855 158.055 37.805 158.145 ;
        RECT 29.275 157.235 31.105 157.915 ;
        RECT 31.115 157.235 34.785 158.045 ;
        RECT 35.875 157.235 37.805 158.055 ;
        RECT 38.015 157.235 43.525 158.045 ;
        RECT 43.535 157.235 45.365 158.045 ;
        RECT 45.375 157.235 48.125 158.145 ;
        RECT 48.135 157.235 49.965 158.045 ;
        RECT 51.820 157.915 53.185 158.145 ;
        RECT 49.975 157.235 53.185 157.915 ;
        RECT 53.195 157.235 54.565 158.045 ;
        RECT 54.585 157.320 55.015 158.105 ;
        RECT 55.465 157.235 58.245 158.145 ;
        RECT 58.255 157.235 60.085 158.045 ;
        RECT 60.555 157.235 62.370 158.145 ;
        RECT 64.660 157.945 65.605 158.145 ;
        RECT 62.855 157.265 65.605 157.945 ;
        RECT 16.075 157.025 16.245 157.235 ;
        RECT 17.430 157.190 17.600 157.215 ;
        RECT 17.430 157.080 17.625 157.190 ;
        RECT 17.430 157.045 17.600 157.080 ;
        RECT 18.380 157.045 18.550 157.235 ;
        RECT 20.220 157.045 20.390 157.235 ;
        RECT 22.065 157.070 22.225 157.180 ;
        RECT 17.490 157.025 17.600 157.045 ;
        RECT 22.975 157.025 23.145 157.215 ;
        RECT 24.810 157.045 24.980 157.235 ;
        RECT 25.275 157.045 25.445 157.235 ;
        RECT 26.655 157.025 26.825 157.215 ;
        RECT 30.795 157.045 30.965 157.235 ;
        RECT 31.255 157.025 31.425 157.235 ;
        RECT 35.875 157.215 36.025 157.235 ;
        RECT 34.945 157.080 35.105 157.190 ;
        RECT 35.855 157.045 36.025 157.215 ;
        RECT 37.235 157.025 37.405 157.215 ;
        RECT 37.695 157.025 37.865 157.215 ;
        RECT 38.155 157.045 38.325 157.235 ;
        RECT 41.370 157.075 41.490 157.185 ;
        RECT 42.285 157.025 42.455 157.215 ;
        RECT 43.675 157.045 43.845 157.235 ;
        RECT 45.515 157.025 45.685 157.235 ;
        RECT 48.275 157.025 48.445 157.235 ;
        RECT 50.120 157.045 50.290 157.235 ;
        RECT 51.030 157.025 51.200 157.215 ;
        RECT 51.495 157.025 51.665 157.215 ;
        RECT 53.335 157.045 53.505 157.235 ;
        RECT 57.015 157.025 57.185 157.215 ;
        RECT 57.935 157.045 58.105 157.235 ;
        RECT 58.395 157.045 58.565 157.235 ;
        RECT 60.230 157.075 60.350 157.185 ;
        RECT 60.695 157.025 60.865 157.215 ;
        RECT 62.075 157.045 62.245 157.235 ;
        RECT 63.000 157.215 63.170 157.265 ;
        RECT 64.660 157.235 65.605 157.265 ;
        RECT 65.615 157.235 68.365 158.045 ;
        RECT 70.205 157.915 71.125 158.145 ;
        RECT 68.835 157.235 71.125 157.915 ;
        RECT 71.155 157.235 72.505 158.145 ;
        RECT 72.515 157.235 76.185 158.045 ;
        RECT 77.115 157.235 78.485 158.015 ;
        RECT 78.495 157.235 80.325 157.915 ;
        RECT 80.345 157.320 80.775 158.105 ;
        RECT 81.740 157.915 83.080 158.145 ;
        RECT 81.255 157.235 85.845 157.915 ;
        RECT 85.855 157.235 87.225 158.045 ;
        RECT 62.530 157.075 62.650 157.185 ;
        RECT 62.995 157.045 63.170 157.215 ;
        RECT 62.995 157.025 63.165 157.045 ;
        RECT 63.455 157.025 63.625 157.215 ;
        RECT 65.755 157.045 65.925 157.235 ;
        RECT 67.130 157.075 67.250 157.185 ;
        RECT 68.510 157.075 68.630 157.185 ;
        RECT 68.975 157.045 69.145 157.235 ;
        RECT 70.355 157.025 70.525 157.215 ;
        RECT 72.190 157.045 72.360 157.235 ;
        RECT 72.655 157.045 72.825 157.235 ;
        RECT 72.655 157.025 72.805 157.045 ;
        RECT 73.115 157.025 73.285 157.215 ;
        RECT 76.345 157.080 76.505 157.190 ;
        RECT 77.265 157.045 77.435 157.235 ;
        RECT 78.645 157.070 78.805 157.180 ;
        RECT 80.015 157.045 80.185 157.235 ;
        RECT 80.465 157.025 80.635 157.215 ;
        RECT 80.945 157.185 81.115 157.215 ;
        RECT 80.930 157.075 81.115 157.185 ;
        RECT 80.945 157.025 81.115 157.075 ;
        RECT 81.400 157.045 81.570 157.235 ;
        RECT 83.695 157.025 83.865 157.215 ;
        RECT 84.155 157.025 84.325 157.215 ;
        RECT 86.915 157.025 87.085 157.235 ;
        RECT 15.935 156.215 17.305 157.025 ;
        RECT 17.490 156.345 21.905 157.025 ;
        RECT 22.835 156.345 26.505 157.025 ;
        RECT 26.515 156.795 28.085 157.025 ;
        RECT 30.175 156.985 31.095 157.025 ;
        RECT 30.175 156.795 31.105 156.985 ;
        RECT 26.515 156.435 31.105 156.795 ;
        RECT 26.515 156.345 31.095 156.435 ;
        RECT 17.975 156.115 21.905 156.345 ;
        RECT 25.575 156.115 26.505 156.345 ;
        RECT 28.095 156.115 31.095 156.345 ;
        RECT 31.115 156.215 33.865 157.025 ;
        RECT 34.015 156.115 37.465 157.025 ;
        RECT 37.555 156.215 41.225 157.025 ;
        RECT 41.705 156.155 42.135 156.940 ;
        RECT 42.155 156.115 45.365 157.025 ;
        RECT 45.385 156.115 48.115 157.025 ;
        RECT 48.135 156.215 49.965 157.025 ;
        RECT 49.995 156.115 51.345 157.025 ;
        RECT 51.355 156.215 56.865 157.025 ;
        RECT 56.875 156.215 60.545 157.025 ;
        RECT 60.555 156.215 61.925 157.025 ;
        RECT 61.945 156.115 63.295 157.025 ;
        RECT 63.315 156.215 66.985 157.025 ;
        RECT 67.465 156.155 67.895 156.940 ;
        RECT 67.925 156.115 70.655 157.025 ;
        RECT 70.875 156.205 72.805 157.025 ;
        RECT 72.975 156.215 78.485 157.025 ;
        RECT 79.415 156.245 80.785 157.025 ;
        RECT 80.795 156.245 82.165 157.025 ;
        RECT 82.175 156.345 84.005 157.025 ;
        RECT 84.015 156.345 85.845 157.025 ;
        RECT 70.875 156.115 71.825 156.205 ;
        RECT 82.175 156.115 83.520 156.345 ;
        RECT 84.500 156.115 85.845 156.345 ;
        RECT 85.855 156.215 87.225 157.025 ;
      LAYER nwell ;
        RECT 15.740 152.995 87.420 155.825 ;
      LAYER pwell ;
        RECT 17.325 152.615 18.915 152.705 ;
        RECT 15.935 151.795 17.305 152.605 ;
        RECT 17.325 151.795 19.895 152.615 ;
        RECT 21.895 152.475 22.825 152.705 ;
        RECT 20.075 151.795 22.825 152.475 ;
        RECT 22.835 151.795 24.665 152.605 ;
        RECT 25.135 152.505 26.065 152.705 ;
        RECT 27.395 152.505 28.345 152.705 ;
        RECT 25.135 152.025 28.345 152.505 ;
        RECT 25.280 151.825 28.345 152.025 ;
        RECT 28.825 151.880 29.255 152.665 ;
        RECT 29.275 152.505 30.205 152.705 ;
        RECT 31.535 152.505 32.485 152.705 ;
        RECT 29.275 152.025 32.485 152.505 ;
        RECT 16.075 151.585 16.245 151.795 ;
        RECT 19.755 151.775 19.895 151.795 ;
        RECT 18.835 151.585 19.005 151.775 ;
        RECT 19.295 151.585 19.465 151.775 ;
        RECT 19.755 151.605 19.925 151.775 ;
        RECT 20.215 151.605 20.385 151.795 ;
        RECT 21.595 151.585 21.765 151.775 ;
        RECT 22.055 151.585 22.225 151.775 ;
        RECT 22.975 151.605 23.145 151.795 ;
        RECT 24.810 151.635 24.930 151.745 ;
        RECT 25.280 151.605 25.450 151.825 ;
        RECT 27.410 151.795 28.345 151.825 ;
        RECT 29.420 151.825 32.485 152.025 ;
        RECT 27.575 151.585 27.745 151.775 ;
        RECT 28.490 151.635 28.610 151.745 ;
        RECT 29.420 151.605 29.590 151.825 ;
        RECT 31.550 151.795 32.485 151.825 ;
        RECT 33.425 151.795 37.545 152.705 ;
        RECT 37.555 151.795 39.385 152.475 ;
        RECT 39.415 151.795 40.765 152.705 ;
        RECT 42.375 152.615 43.325 152.705 ;
        RECT 41.395 151.795 43.325 152.615 ;
        RECT 43.535 152.025 45.370 152.705 ;
        RECT 43.680 151.795 45.370 152.025 ;
        RECT 45.835 151.795 47.665 152.605 ;
        RECT 48.135 151.795 51.805 152.705 ;
        RECT 52.300 152.475 53.645 152.705 ;
        RECT 51.815 151.795 53.645 152.475 ;
        RECT 54.585 151.880 55.015 152.665 ;
        RECT 55.035 151.795 58.245 152.705 ;
        RECT 58.295 152.475 59.670 152.705 ;
        RECT 61.460 152.475 62.840 152.705 ;
        RECT 58.295 152.025 62.840 152.475 ;
        RECT 32.645 151.640 32.805 151.750 ;
        RECT 33.095 151.585 33.265 151.775 ;
        RECT 34.935 151.585 35.105 151.775 ;
        RECT 35.395 151.605 35.565 151.795 ;
        RECT 36.775 151.585 36.945 151.775 ;
        RECT 37.235 151.605 37.405 151.795 ;
        RECT 39.075 151.605 39.245 151.795 ;
        RECT 40.450 151.775 40.620 151.795 ;
        RECT 41.395 151.775 41.545 151.795 ;
        RECT 40.450 151.605 40.625 151.775 ;
        RECT 40.910 151.635 41.030 151.745 ;
        RECT 41.375 151.605 41.545 151.775 ;
        RECT 40.455 151.585 40.625 151.605 ;
        RECT 42.295 151.585 42.465 151.775 ;
        RECT 43.680 151.605 43.850 151.795 ;
        RECT 45.975 151.605 46.145 151.795 ;
        RECT 47.810 151.635 47.930 151.745 ;
        RECT 48.275 151.585 48.445 151.795 ;
        RECT 51.955 151.605 52.125 151.795 ;
        RECT 53.795 151.605 53.965 151.775 ;
        RECT 53.795 151.585 53.960 151.605 ;
        RECT 54.260 151.585 54.430 151.775 ;
        RECT 55.175 151.605 55.345 151.795 ;
        RECT 55.635 151.585 55.805 151.775 ;
        RECT 58.400 151.605 58.570 152.025 ;
        RECT 59.680 151.795 62.840 152.025 ;
        RECT 62.855 151.795 64.205 152.705 ;
        RECT 64.235 151.795 65.605 152.605 ;
        RECT 65.625 151.795 68.355 152.705 ;
        RECT 68.375 151.795 70.190 152.705 ;
        RECT 70.215 151.795 75.725 152.605 ;
        RECT 75.735 151.795 79.405 152.605 ;
        RECT 80.345 151.880 80.775 152.665 ;
        RECT 80.795 151.795 82.625 152.605 ;
        RECT 82.635 151.795 84.005 152.575 ;
        RECT 84.015 151.795 85.845 152.475 ;
        RECT 85.855 151.795 87.225 152.605 ;
        RECT 58.850 151.585 59.020 151.775 ;
        RECT 60.235 151.585 60.405 151.775 ;
        RECT 63.920 151.605 64.090 151.795 ;
        RECT 64.375 151.605 64.545 151.795 ;
        RECT 67.135 151.585 67.305 151.775 ;
        RECT 68.055 151.585 68.225 151.795 ;
        RECT 69.895 151.605 70.065 151.795 ;
        RECT 70.355 151.605 70.525 151.795 ;
        RECT 73.575 151.585 73.745 151.775 ;
        RECT 75.875 151.605 76.045 151.795 ;
        RECT 79.095 151.585 79.265 151.775 ;
        RECT 79.565 151.640 79.725 151.750 ;
        RECT 80.935 151.605 81.105 151.795 ;
        RECT 82.785 151.605 82.955 151.795 ;
        RECT 84.155 151.605 84.325 151.795 ;
        RECT 85.535 151.585 85.705 151.775 ;
        RECT 86.915 151.585 87.085 151.795 ;
        RECT 15.935 150.775 17.305 151.585 ;
        RECT 17.315 150.905 19.145 151.585 ;
        RECT 17.315 150.675 18.660 150.905 ;
        RECT 19.165 150.675 20.515 151.585 ;
        RECT 20.535 150.805 21.905 151.585 ;
        RECT 21.915 150.775 27.425 151.585 ;
        RECT 27.435 150.775 32.945 151.585 ;
        RECT 32.970 150.675 34.785 151.585 ;
        RECT 34.795 150.905 36.625 151.585 ;
        RECT 35.280 150.675 36.625 150.905 ;
        RECT 36.635 150.775 40.305 151.585 ;
        RECT 40.315 150.775 41.685 151.585 ;
        RECT 41.705 150.715 42.135 151.500 ;
        RECT 42.155 150.775 47.665 151.585 ;
        RECT 48.135 150.675 51.805 151.585 ;
        RECT 52.125 150.905 53.960 151.585 ;
        RECT 52.125 150.675 53.055 150.905 ;
        RECT 54.115 150.675 55.465 151.585 ;
        RECT 55.495 150.675 58.705 151.585 ;
        RECT 58.735 150.675 60.085 151.585 ;
        RECT 60.095 150.775 65.605 151.585 ;
        RECT 65.615 150.675 67.430 151.585 ;
        RECT 67.465 150.715 67.895 151.500 ;
        RECT 67.915 150.775 73.425 151.585 ;
        RECT 73.435 150.775 78.945 151.585 ;
        RECT 78.955 150.775 84.465 151.585 ;
        RECT 84.475 150.805 85.845 151.585 ;
        RECT 85.855 150.775 87.225 151.585 ;
      LAYER nwell ;
        RECT 15.740 147.555 87.420 150.385 ;
      LAYER pwell ;
        RECT 15.935 146.355 17.305 147.165 ;
        RECT 17.315 146.355 22.825 147.165 ;
        RECT 22.835 146.355 28.345 147.165 ;
        RECT 28.825 146.440 29.255 147.225 ;
        RECT 29.275 146.355 31.105 147.165 ;
        RECT 31.595 146.355 32.945 147.265 ;
        RECT 32.955 146.355 36.615 147.265 ;
        RECT 36.805 146.355 40.305 147.265 ;
        RECT 40.315 146.355 43.065 147.165 ;
        RECT 43.085 146.585 46.285 147.265 ;
        RECT 43.085 146.355 46.140 146.585 ;
        RECT 46.295 146.355 51.805 147.165 ;
        RECT 51.815 146.355 54.565 147.165 ;
        RECT 54.585 146.440 55.015 147.225 ;
        RECT 55.530 147.035 56.905 147.265 ;
        RECT 58.675 147.035 59.625 147.265 ;
        RECT 60.120 147.035 61.465 147.265 ;
        RECT 61.960 147.035 65.570 147.265 ;
        RECT 55.530 146.585 59.625 147.035 ;
        RECT 16.075 146.145 16.245 146.355 ;
        RECT 17.455 146.145 17.625 146.355 ;
        RECT 22.975 146.145 23.145 146.355 ;
        RECT 28.495 146.305 28.665 146.335 ;
        RECT 28.490 146.195 28.665 146.305 ;
        RECT 28.495 146.145 28.665 146.195 ;
        RECT 29.415 146.165 29.585 146.355 ;
        RECT 31.250 146.195 31.370 146.305 ;
        RECT 31.710 146.165 31.880 146.355 ;
        RECT 35.390 146.145 35.560 146.335 ;
        RECT 36.330 146.165 36.500 146.355 ;
        RECT 36.805 146.335 36.940 146.355 ;
        RECT 36.770 146.165 36.940 146.335 ;
        RECT 37.695 146.165 37.865 146.335 ;
        RECT 38.165 146.190 38.325 146.300 ;
        RECT 37.695 146.145 37.845 146.165 ;
        RECT 39.080 146.145 39.250 146.335 ;
        RECT 40.455 146.165 40.625 146.355 ;
        RECT 41.370 146.195 41.490 146.305 ;
        RECT 43.675 146.145 43.845 146.335 ;
        RECT 44.135 146.145 44.305 146.335 ;
        RECT 45.515 146.145 45.685 146.335 ;
        RECT 45.970 146.165 46.140 146.355 ;
        RECT 46.435 146.165 46.605 146.355 ;
        RECT 51.035 146.145 51.205 146.335 ;
        RECT 51.955 146.165 52.125 146.355 ;
        RECT 55.170 146.195 55.290 146.305 ;
        RECT 55.635 146.165 55.805 146.585 ;
        RECT 56.915 146.355 59.625 146.585 ;
        RECT 59.635 146.355 61.465 147.035 ;
        RECT 61.475 146.355 65.570 147.035 ;
        RECT 65.615 146.355 71.125 147.165 ;
        RECT 71.135 146.355 76.645 147.165 ;
        RECT 76.655 146.355 80.325 147.165 ;
        RECT 80.345 146.440 80.775 147.225 ;
        RECT 80.795 146.355 83.545 147.165 ;
        RECT 84.015 146.355 85.845 147.035 ;
        RECT 85.855 146.355 87.225 147.165 ;
        RECT 56.555 146.145 56.725 146.335 ;
        RECT 59.775 146.165 59.945 146.355 ;
        RECT 60.230 146.195 60.350 146.305 ;
        RECT 61.620 146.165 61.790 146.355 ;
        RECT 64.370 146.145 64.540 146.335 ;
        RECT 64.835 146.145 65.005 146.335 ;
        RECT 65.755 146.165 65.925 146.355 ;
        RECT 68.055 146.145 68.225 146.335 ;
        RECT 71.275 146.165 71.445 146.355 ;
        RECT 73.575 146.145 73.745 146.335 ;
        RECT 76.795 146.165 76.965 146.355 ;
        RECT 79.095 146.145 79.265 146.335 ;
        RECT 80.935 146.165 81.105 146.355 ;
        RECT 83.690 146.195 83.810 146.305 ;
        RECT 85.535 146.165 85.705 146.355 ;
        RECT 86.915 146.145 87.085 146.355 ;
        RECT 15.935 145.335 17.305 146.145 ;
        RECT 17.315 145.335 22.825 146.145 ;
        RECT 22.835 145.335 28.345 146.145 ;
        RECT 28.355 145.335 33.865 146.145 ;
        RECT 33.875 145.235 35.705 146.145 ;
        RECT 35.915 145.325 37.845 146.145 ;
        RECT 38.935 145.465 41.210 146.145 ;
        RECT 35.915 145.235 36.865 145.325 ;
        RECT 39.840 145.235 41.210 145.465 ;
        RECT 41.705 145.275 42.135 146.060 ;
        RECT 42.155 145.465 43.985 146.145 ;
        RECT 43.995 145.365 45.365 146.145 ;
        RECT 45.375 145.335 50.885 146.145 ;
        RECT 50.895 145.335 56.405 146.145 ;
        RECT 56.415 145.335 60.085 146.145 ;
        RECT 60.590 145.465 64.685 146.145 ;
        RECT 60.590 145.235 64.200 145.465 ;
        RECT 64.695 145.335 67.445 146.145 ;
        RECT 67.465 145.275 67.895 146.060 ;
        RECT 67.915 145.335 73.425 146.145 ;
        RECT 73.435 145.335 78.945 146.145 ;
        RECT 78.955 145.335 84.465 146.145 ;
        RECT 85.855 145.335 87.225 146.145 ;
      LAYER nwell ;
        RECT 15.740 142.115 87.420 144.945 ;
      LAYER pwell ;
        RECT 15.935 140.915 17.305 141.725 ;
        RECT 17.315 140.915 22.825 141.725 ;
        RECT 25.135 140.915 28.805 141.725 ;
        RECT 28.825 141.000 29.255 141.785 ;
        RECT 29.275 140.915 32.945 141.725 ;
        RECT 33.415 140.915 34.785 141.695 ;
        RECT 34.795 140.915 36.625 141.725 ;
        RECT 37.120 141.595 38.465 141.825 ;
        RECT 36.635 140.915 38.465 141.595 ;
        RECT 38.475 140.915 39.825 141.825 ;
        RECT 39.855 140.915 41.225 141.695 ;
        RECT 41.705 141.000 42.135 141.785 ;
        RECT 43.075 140.915 44.905 141.595 ;
        RECT 44.915 140.915 46.285 141.725 ;
        RECT 46.780 141.595 48.125 141.825 ;
        RECT 46.295 140.915 48.125 141.595 ;
        RECT 48.135 140.915 53.645 141.725 ;
        RECT 54.585 141.000 55.015 141.785 ;
        RECT 55.035 140.915 60.545 141.725 ;
        RECT 60.555 140.915 66.065 141.725 ;
        RECT 66.075 140.915 67.445 141.725 ;
        RECT 67.465 141.000 67.895 141.785 ;
        RECT 67.915 140.915 73.425 141.725 ;
        RECT 73.435 140.915 78.945 141.725 ;
        RECT 78.955 140.915 80.325 141.725 ;
        RECT 80.345 141.000 80.775 141.785 ;
        RECT 80.795 140.915 84.465 141.725 ;
        RECT 84.475 140.915 85.845 141.725 ;
        RECT 85.855 140.915 87.225 141.725 ;
        RECT 16.075 140.725 16.245 140.915 ;
        RECT 17.455 140.725 17.625 140.915 ;
        RECT 22.985 140.760 23.145 140.870 ;
        RECT 24.815 140.725 24.985 140.895 ;
        RECT 25.275 140.725 25.445 140.915 ;
        RECT 29.415 140.725 29.585 140.915 ;
        RECT 33.090 140.755 33.210 140.865 ;
        RECT 34.475 140.725 34.645 140.915 ;
        RECT 34.935 140.725 35.105 140.915 ;
        RECT 36.775 140.725 36.945 140.915 ;
        RECT 39.540 140.725 39.710 140.915 ;
        RECT 40.005 140.725 40.175 140.915 ;
        RECT 41.370 140.755 41.490 140.865 ;
        RECT 42.305 140.760 42.465 140.870 ;
        RECT 43.215 140.725 43.385 140.915 ;
        RECT 45.055 140.725 45.225 140.915 ;
        RECT 46.435 140.725 46.605 140.915 ;
        RECT 48.275 140.725 48.445 140.915 ;
        RECT 53.805 140.760 53.965 140.870 ;
        RECT 55.175 140.725 55.345 140.915 ;
        RECT 60.695 140.725 60.865 140.915 ;
        RECT 66.215 140.725 66.385 140.915 ;
        RECT 68.055 140.725 68.225 140.915 ;
        RECT 73.575 140.725 73.745 140.915 ;
        RECT 79.095 140.725 79.265 140.915 ;
        RECT 80.935 140.725 81.105 140.915 ;
        RECT 84.615 140.725 84.785 140.915 ;
        RECT 86.915 140.725 87.085 140.915 ;
      LAYER li1 ;
        RECT 15.930 211.445 87.230 211.615 ;
        RECT 16.015 210.695 17.225 211.445 ;
        RECT 16.015 210.155 16.535 210.695 ;
        RECT 17.455 210.625 17.665 211.445 ;
        RECT 17.835 210.645 18.165 211.275 ;
        RECT 16.705 209.985 17.225 210.525 ;
        RECT 17.835 210.045 18.085 210.645 ;
        RECT 18.335 210.625 18.565 211.445 ;
        RECT 18.865 210.895 19.035 211.275 ;
        RECT 19.250 211.065 19.580 211.445 ;
        RECT 18.865 210.725 19.580 210.895 ;
        RECT 18.255 210.205 18.585 210.455 ;
        RECT 18.775 210.175 19.130 210.545 ;
        RECT 19.410 210.535 19.580 210.725 ;
        RECT 19.750 210.700 20.005 211.275 ;
        RECT 19.410 210.205 19.665 210.535 ;
        RECT 16.015 208.895 17.225 209.985 ;
        RECT 17.455 208.895 17.665 210.035 ;
        RECT 17.835 209.065 18.165 210.045 ;
        RECT 18.335 208.895 18.565 210.035 ;
        RECT 19.410 209.995 19.580 210.205 ;
        RECT 18.865 209.825 19.580 209.995 ;
        RECT 19.835 209.970 20.005 210.700 ;
        RECT 20.180 210.605 20.440 211.445 ;
        RECT 20.620 210.605 20.880 211.445 ;
        RECT 21.055 210.700 21.310 211.275 ;
        RECT 21.480 211.065 21.810 211.445 ;
        RECT 22.025 210.895 22.195 211.275 ;
        RECT 21.480 210.725 22.195 210.895 ;
        RECT 18.865 209.065 19.035 209.825 ;
        RECT 19.250 208.895 19.580 209.655 ;
        RECT 19.750 209.065 20.005 209.970 ;
        RECT 20.180 208.895 20.440 210.045 ;
        RECT 20.620 208.895 20.880 210.045 ;
        RECT 21.055 209.970 21.225 210.700 ;
        RECT 21.480 210.535 21.650 210.725 ;
        RECT 22.460 210.605 22.720 211.445 ;
        RECT 22.895 210.700 23.150 211.275 ;
        RECT 23.320 211.065 23.650 211.445 ;
        RECT 23.865 210.895 24.035 211.275 ;
        RECT 24.460 210.935 24.700 211.445 ;
        RECT 24.880 210.935 25.160 211.265 ;
        RECT 25.390 210.935 25.605 211.445 ;
        RECT 23.320 210.725 24.035 210.895 ;
        RECT 21.395 210.205 21.650 210.535 ;
        RECT 21.480 209.995 21.650 210.205 ;
        RECT 21.930 210.175 22.285 210.545 ;
        RECT 21.055 209.065 21.310 209.970 ;
        RECT 21.480 209.825 22.195 209.995 ;
        RECT 21.480 208.895 21.810 209.655 ;
        RECT 22.025 209.065 22.195 209.825 ;
        RECT 22.460 208.895 22.720 210.045 ;
        RECT 22.895 209.970 23.065 210.700 ;
        RECT 23.320 210.535 23.490 210.725 ;
        RECT 23.235 210.205 23.490 210.535 ;
        RECT 23.320 209.995 23.490 210.205 ;
        RECT 23.770 210.175 24.125 210.545 ;
        RECT 24.355 210.205 24.710 210.765 ;
        RECT 24.880 210.035 25.050 210.935 ;
        RECT 25.220 210.205 25.485 210.765 ;
        RECT 25.775 210.705 26.390 211.275 ;
        RECT 26.705 211.065 27.875 211.275 ;
        RECT 26.705 211.045 27.035 211.065 ;
        RECT 25.735 210.035 25.905 210.535 ;
        RECT 22.895 209.065 23.150 209.970 ;
        RECT 23.320 209.825 24.035 209.995 ;
        RECT 23.320 208.895 23.650 209.655 ;
        RECT 23.865 209.065 24.035 209.825 ;
        RECT 24.480 209.865 25.905 210.035 ;
        RECT 24.480 209.690 24.870 209.865 ;
        RECT 25.355 208.895 25.685 209.695 ;
        RECT 26.075 209.685 26.390 210.705 ;
        RECT 26.595 210.625 27.455 210.875 ;
        RECT 27.625 210.815 27.875 211.065 ;
        RECT 28.045 210.985 28.215 211.445 ;
        RECT 28.385 210.815 28.725 211.275 ;
        RECT 27.625 210.645 28.725 210.815 ;
        RECT 28.895 210.720 29.185 211.445 ;
        RECT 29.465 211.065 30.635 211.275 ;
        RECT 29.465 211.045 29.795 211.065 ;
        RECT 29.355 210.625 30.215 210.875 ;
        RECT 30.385 210.815 30.635 211.065 ;
        RECT 30.805 210.985 30.975 211.445 ;
        RECT 31.145 210.815 31.485 211.275 ;
        RECT 30.385 210.645 31.485 210.815 ;
        RECT 31.855 210.815 32.185 211.175 ;
        RECT 32.815 210.985 33.065 211.445 ;
        RECT 33.235 210.985 33.785 211.275 ;
        RECT 31.855 210.625 33.245 210.815 ;
        RECT 26.595 210.035 26.875 210.625 ;
        RECT 27.045 210.205 27.795 210.455 ;
        RECT 27.965 210.205 28.725 210.455 ;
        RECT 26.595 209.865 28.295 210.035 ;
        RECT 25.855 209.065 26.390 209.685 ;
        RECT 26.700 208.895 26.955 209.695 ;
        RECT 27.125 209.065 27.455 209.865 ;
        RECT 27.625 208.895 27.795 209.695 ;
        RECT 27.965 209.065 28.295 209.865 ;
        RECT 28.465 208.895 28.725 210.035 ;
        RECT 28.895 208.895 29.185 210.060 ;
        RECT 29.355 210.035 29.635 210.625 ;
        RECT 33.075 210.535 33.245 210.625 ;
        RECT 29.805 210.205 30.555 210.455 ;
        RECT 30.725 210.205 31.485 210.455 ;
        RECT 31.655 210.205 32.345 210.455 ;
        RECT 32.575 210.205 32.905 210.455 ;
        RECT 33.075 210.205 33.365 210.535 ;
        RECT 29.355 209.865 31.055 210.035 ;
        RECT 29.460 208.895 29.715 209.695 ;
        RECT 29.885 209.065 30.215 209.865 ;
        RECT 30.385 208.895 30.555 209.695 ;
        RECT 30.725 209.065 31.055 209.865 ;
        RECT 31.225 208.895 31.485 210.035 ;
        RECT 31.655 209.765 31.970 210.205 ;
        RECT 33.075 209.955 33.245 210.205 ;
        RECT 32.305 209.785 33.245 209.955 ;
        RECT 31.855 208.895 32.135 209.565 ;
        RECT 32.305 209.235 32.605 209.785 ;
        RECT 33.535 209.615 33.785 210.985 ;
        RECT 33.955 210.645 34.245 211.445 ;
        RECT 34.500 210.945 34.995 211.275 ;
        RECT 32.815 208.895 33.145 209.615 ;
        RECT 33.335 209.065 33.785 209.615 ;
        RECT 33.955 208.895 34.245 210.035 ;
        RECT 34.415 209.455 34.655 210.765 ;
        RECT 34.825 210.035 34.995 210.945 ;
        RECT 35.215 210.205 35.565 211.170 ;
        RECT 35.745 210.205 36.045 211.175 ;
        RECT 36.225 210.205 36.505 211.175 ;
        RECT 36.685 210.645 36.955 211.445 ;
        RECT 37.125 210.725 37.465 211.235 ;
        RECT 37.720 210.895 38.050 211.275 ;
        RECT 38.220 211.065 39.405 211.235 ;
        RECT 39.665 210.975 39.835 211.445 ;
        RECT 37.720 210.725 38.265 210.895 ;
        RECT 36.700 210.205 37.030 210.455 ;
        RECT 36.700 210.035 37.015 210.205 ;
        RECT 34.825 209.865 37.015 210.035 ;
        RECT 34.420 208.895 34.755 209.275 ;
        RECT 34.925 209.065 35.175 209.865 ;
        RECT 35.395 208.895 35.725 209.615 ;
        RECT 35.910 209.065 36.160 209.865 ;
        RECT 36.625 208.895 36.955 209.695 ;
        RECT 37.205 209.325 37.465 210.725 ;
        RECT 37.635 210.205 37.895 210.555 ;
        RECT 38.095 210.085 38.265 210.725 ;
        RECT 38.635 210.795 39.020 210.885 ;
        RECT 40.005 210.795 40.335 211.260 ;
        RECT 38.635 210.625 40.335 210.795 ;
        RECT 40.505 210.625 40.675 211.445 ;
        RECT 40.845 210.795 41.175 211.265 ;
        RECT 41.345 210.965 41.515 211.445 ;
        RECT 40.845 210.625 41.605 210.795 ;
        RECT 41.775 210.720 42.065 211.445 ;
        RECT 43.245 210.965 43.545 211.445 ;
        RECT 43.715 210.795 43.975 211.250 ;
        RECT 44.145 210.965 44.405 211.445 ;
        RECT 44.585 210.795 44.845 211.250 ;
        RECT 45.015 210.965 45.265 211.445 ;
        RECT 45.445 210.795 45.705 211.250 ;
        RECT 45.875 210.965 46.125 211.445 ;
        RECT 46.305 210.795 46.565 211.250 ;
        RECT 46.735 210.965 46.980 211.445 ;
        RECT 47.150 210.795 47.425 211.250 ;
        RECT 47.595 210.965 47.840 211.445 ;
        RECT 48.010 210.795 48.270 211.250 ;
        RECT 48.440 210.965 48.700 211.445 ;
        RECT 48.870 210.795 49.130 211.250 ;
        RECT 49.300 210.965 49.560 211.445 ;
        RECT 49.730 210.795 49.990 211.250 ;
        RECT 50.160 210.885 50.420 211.445 ;
        RECT 43.245 210.765 49.990 210.795 ;
        RECT 38.435 210.255 38.780 210.455 ;
        RECT 38.950 210.255 39.340 210.455 ;
        RECT 38.095 210.035 38.880 210.085 ;
        RECT 37.125 209.065 37.465 209.325 ;
        RECT 37.800 209.860 38.880 210.035 ;
        RECT 37.800 209.065 38.130 209.860 ;
        RECT 38.300 208.895 38.540 209.680 ;
        RECT 38.710 209.655 38.880 209.860 ;
        RECT 39.050 209.825 39.340 210.255 ;
        RECT 39.530 210.245 40.015 210.455 ;
        RECT 40.185 210.245 40.625 210.455 ;
        RECT 40.795 210.245 41.125 210.455 ;
        RECT 39.530 209.825 39.835 210.245 ;
        RECT 40.795 210.075 40.965 210.245 ;
        RECT 40.005 209.905 40.965 210.075 ;
        RECT 40.005 209.655 40.175 209.905 ;
        RECT 38.710 209.485 40.175 209.655 ;
        RECT 39.100 209.065 39.855 209.485 ;
        RECT 40.345 208.895 40.675 209.735 ;
        RECT 41.295 209.655 41.605 210.625 ;
        RECT 43.215 210.625 49.990 210.765 ;
        RECT 43.215 210.595 44.410 210.625 ;
        RECT 40.845 209.485 41.605 209.655 ;
        RECT 40.845 209.065 41.095 209.485 ;
        RECT 41.265 208.895 41.605 209.315 ;
        RECT 41.775 208.895 42.065 210.060 ;
        RECT 43.245 210.035 44.410 210.595 ;
        RECT 50.590 210.455 50.840 211.265 ;
        RECT 51.020 210.920 51.280 211.445 ;
        RECT 51.450 210.455 51.700 211.265 ;
        RECT 51.880 210.935 52.185 211.445 ;
        RECT 52.375 210.935 52.615 211.445 ;
        RECT 52.785 210.935 53.075 211.275 ;
        RECT 53.305 210.935 53.620 211.445 ;
        RECT 44.580 210.205 51.700 210.455 ;
        RECT 51.870 210.205 52.185 210.765 ;
        RECT 52.420 210.425 52.615 210.765 ;
        RECT 52.415 210.255 52.615 210.425 ;
        RECT 52.420 210.205 52.615 210.255 ;
        RECT 43.245 209.810 49.990 210.035 ;
        RECT 43.245 208.895 43.515 209.640 ;
        RECT 43.685 209.070 43.975 209.810 ;
        RECT 44.585 209.795 49.990 209.810 ;
        RECT 44.145 208.900 44.400 209.625 ;
        RECT 44.585 209.070 44.845 209.795 ;
        RECT 45.015 208.900 45.260 209.625 ;
        RECT 45.445 209.070 45.705 209.795 ;
        RECT 45.875 208.900 46.120 209.625 ;
        RECT 46.305 209.070 46.565 209.795 ;
        RECT 46.735 208.900 46.980 209.625 ;
        RECT 47.150 209.070 47.410 209.795 ;
        RECT 47.580 208.900 47.840 209.625 ;
        RECT 48.010 209.070 48.270 209.795 ;
        RECT 48.440 208.900 48.700 209.625 ;
        RECT 48.870 209.070 49.130 209.795 ;
        RECT 49.300 208.900 49.560 209.625 ;
        RECT 49.730 209.070 49.990 209.795 ;
        RECT 50.160 208.900 50.420 209.695 ;
        RECT 50.590 209.070 50.840 210.205 ;
        RECT 44.145 208.895 50.420 208.900 ;
        RECT 51.020 208.895 51.280 209.705 ;
        RECT 51.455 209.065 51.700 210.205 ;
        RECT 52.785 210.035 52.965 210.935 ;
        RECT 53.790 210.875 53.960 211.145 ;
        RECT 54.130 211.045 54.460 211.445 ;
        RECT 53.135 210.205 53.545 210.765 ;
        RECT 53.790 210.705 54.485 210.875 ;
        RECT 54.655 210.720 54.945 211.445 ;
        RECT 55.445 211.045 55.775 211.445 ;
        RECT 55.945 210.875 56.275 211.215 ;
        RECT 57.325 211.045 57.655 211.445 ;
        RECT 53.715 210.035 53.885 210.535 ;
        RECT 52.425 209.865 53.885 210.035 ;
        RECT 51.880 208.895 52.175 209.705 ;
        RECT 52.425 209.690 52.785 209.865 ;
        RECT 54.055 209.695 54.485 210.705 ;
        RECT 55.290 210.705 57.655 210.875 ;
        RECT 57.825 210.720 58.155 211.230 ;
        RECT 58.425 210.965 58.725 211.445 ;
        RECT 58.895 210.795 59.155 211.250 ;
        RECT 59.325 210.965 59.585 211.445 ;
        RECT 59.765 210.795 60.025 211.250 ;
        RECT 60.195 210.965 60.445 211.445 ;
        RECT 60.625 210.795 60.885 211.250 ;
        RECT 61.055 210.965 61.305 211.445 ;
        RECT 61.485 210.795 61.745 211.250 ;
        RECT 61.915 210.965 62.160 211.445 ;
        RECT 62.330 210.795 62.605 211.250 ;
        RECT 62.775 210.965 63.020 211.445 ;
        RECT 63.190 210.795 63.450 211.250 ;
        RECT 63.620 210.965 63.880 211.445 ;
        RECT 64.050 210.795 64.310 211.250 ;
        RECT 64.480 210.965 64.740 211.445 ;
        RECT 64.910 210.795 65.170 211.250 ;
        RECT 65.340 210.885 65.600 211.445 ;
        RECT 53.370 208.895 53.540 209.695 ;
        RECT 53.710 209.525 54.485 209.695 ;
        RECT 53.710 209.065 54.040 209.525 ;
        RECT 54.210 208.895 54.380 209.355 ;
        RECT 54.655 208.895 54.945 210.060 ;
        RECT 55.290 209.705 55.460 210.705 ;
        RECT 57.485 210.535 57.655 210.705 ;
        RECT 55.630 209.875 55.875 210.535 ;
        RECT 56.090 209.875 56.355 210.535 ;
        RECT 56.550 209.875 56.835 210.535 ;
        RECT 57.010 210.205 57.315 210.535 ;
        RECT 57.485 210.205 57.795 210.535 ;
        RECT 57.010 209.875 57.225 210.205 ;
        RECT 57.965 210.085 58.155 210.720 ;
        RECT 55.290 209.535 55.745 209.705 ;
        RECT 55.415 209.105 55.745 209.535 ;
        RECT 55.925 209.535 57.215 209.705 ;
        RECT 55.925 209.115 56.175 209.535 ;
        RECT 56.405 208.895 56.735 209.365 ;
        RECT 56.965 209.115 57.215 209.535 ;
        RECT 57.405 208.895 57.655 210.035 ;
        RECT 57.935 209.955 58.155 210.085 ;
        RECT 57.825 209.105 58.155 209.955 ;
        RECT 58.425 210.625 65.170 210.795 ;
        RECT 58.425 210.035 59.590 210.625 ;
        RECT 65.770 210.455 66.020 211.265 ;
        RECT 66.200 210.920 66.460 211.445 ;
        RECT 66.630 210.455 66.880 211.265 ;
        RECT 67.060 210.935 67.365 211.445 ;
        RECT 59.760 210.205 66.880 210.455 ;
        RECT 67.050 210.205 67.365 210.765 ;
        RECT 67.535 210.720 67.825 211.445 ;
        RECT 68.005 210.715 68.305 211.445 ;
        RECT 68.485 210.535 68.715 211.155 ;
        RECT 68.915 210.885 69.140 211.265 ;
        RECT 69.310 211.055 69.640 211.445 ;
        RECT 69.835 210.935 70.140 211.445 ;
        RECT 68.915 210.705 69.245 210.885 ;
        RECT 68.010 210.205 68.305 210.535 ;
        RECT 68.485 210.205 68.900 210.535 ;
        RECT 58.425 209.810 65.170 210.035 ;
        RECT 58.425 208.895 58.695 209.640 ;
        RECT 58.865 209.070 59.155 209.810 ;
        RECT 59.765 209.795 65.170 209.810 ;
        RECT 59.325 208.900 59.580 209.625 ;
        RECT 59.765 209.070 60.025 209.795 ;
        RECT 60.195 208.900 60.440 209.625 ;
        RECT 60.625 209.070 60.885 209.795 ;
        RECT 61.055 208.900 61.300 209.625 ;
        RECT 61.485 209.070 61.745 209.795 ;
        RECT 61.915 208.900 62.160 209.625 ;
        RECT 62.330 209.070 62.590 209.795 ;
        RECT 62.760 208.900 63.020 209.625 ;
        RECT 63.190 209.070 63.450 209.795 ;
        RECT 63.620 208.900 63.880 209.625 ;
        RECT 64.050 209.070 64.310 209.795 ;
        RECT 64.480 208.900 64.740 209.625 ;
        RECT 64.910 209.070 65.170 209.795 ;
        RECT 65.340 208.900 65.600 209.695 ;
        RECT 65.770 209.070 66.020 210.205 ;
        RECT 59.325 208.895 65.600 208.900 ;
        RECT 66.200 208.895 66.460 209.705 ;
        RECT 66.635 209.065 66.880 210.205 ;
        RECT 67.060 208.895 67.355 209.705 ;
        RECT 67.535 208.895 67.825 210.060 ;
        RECT 69.070 210.035 69.245 210.705 ;
        RECT 69.415 210.205 69.655 210.855 ;
        RECT 69.835 210.205 70.150 210.765 ;
        RECT 70.320 210.455 70.570 211.265 ;
        RECT 70.740 210.920 71.000 211.445 ;
        RECT 71.180 210.455 71.430 211.265 ;
        RECT 71.600 210.885 71.860 211.445 ;
        RECT 72.030 210.795 72.290 211.250 ;
        RECT 72.460 210.965 72.720 211.445 ;
        RECT 72.890 210.795 73.150 211.250 ;
        RECT 73.320 210.965 73.580 211.445 ;
        RECT 73.750 210.795 74.010 211.250 ;
        RECT 74.180 210.965 74.425 211.445 ;
        RECT 74.595 210.795 74.870 211.250 ;
        RECT 75.040 210.965 75.285 211.445 ;
        RECT 75.455 210.795 75.715 211.250 ;
        RECT 75.895 210.965 76.145 211.445 ;
        RECT 76.315 210.795 76.575 211.250 ;
        RECT 76.755 210.965 77.005 211.445 ;
        RECT 77.175 210.795 77.435 211.250 ;
        RECT 77.615 210.965 77.875 211.445 ;
        RECT 78.045 210.795 78.305 211.250 ;
        RECT 78.475 210.965 78.775 211.445 ;
        RECT 72.030 210.625 78.775 210.795 ;
        RECT 79.075 210.625 79.305 211.445 ;
        RECT 79.475 210.645 79.805 211.275 ;
        RECT 70.320 210.205 77.440 210.455 ;
        RECT 68.005 209.675 68.900 210.005 ;
        RECT 69.070 209.845 69.655 210.035 ;
        RECT 68.005 209.505 69.210 209.675 ;
        RECT 68.005 209.075 68.335 209.505 ;
        RECT 68.515 208.895 68.710 209.335 ;
        RECT 68.880 209.075 69.210 209.505 ;
        RECT 69.380 209.075 69.655 209.845 ;
        RECT 69.845 208.895 70.140 209.705 ;
        RECT 70.320 209.065 70.565 210.205 ;
        RECT 70.740 208.895 71.000 209.705 ;
        RECT 71.180 209.070 71.430 210.205 ;
        RECT 77.610 210.085 78.775 210.625 ;
        RECT 79.055 210.205 79.385 210.455 ;
        RECT 77.610 210.035 78.805 210.085 ;
        RECT 79.555 210.045 79.805 210.645 ;
        RECT 79.975 210.625 80.185 211.445 ;
        RECT 80.415 210.720 80.705 211.445 ;
        RECT 72.030 209.915 78.805 210.035 ;
        RECT 72.030 209.810 78.775 209.915 ;
        RECT 72.030 209.795 77.435 209.810 ;
        RECT 71.600 208.900 71.860 209.695 ;
        RECT 72.030 209.070 72.290 209.795 ;
        RECT 72.460 208.900 72.720 209.625 ;
        RECT 72.890 209.070 73.150 209.795 ;
        RECT 73.320 208.900 73.580 209.625 ;
        RECT 73.750 209.070 74.010 209.795 ;
        RECT 74.180 208.900 74.440 209.625 ;
        RECT 74.610 209.070 74.870 209.795 ;
        RECT 75.040 208.900 75.285 209.625 ;
        RECT 75.455 209.070 75.715 209.795 ;
        RECT 75.900 208.900 76.145 209.625 ;
        RECT 76.315 209.070 76.575 209.795 ;
        RECT 76.760 208.900 77.005 209.625 ;
        RECT 77.175 209.070 77.435 209.795 ;
        RECT 77.620 208.900 77.875 209.625 ;
        RECT 78.045 209.070 78.335 209.810 ;
        RECT 71.600 208.895 77.875 208.900 ;
        RECT 78.505 208.895 78.775 209.640 ;
        RECT 79.075 208.895 79.305 210.035 ;
        RECT 79.475 209.065 79.805 210.045 ;
        RECT 79.975 208.895 80.185 210.035 ;
        RECT 80.415 208.895 80.705 210.060 ;
        RECT 80.895 209.865 81.125 211.205 ;
        RECT 81.305 210.365 81.535 211.265 ;
        RECT 81.735 210.665 81.980 211.445 ;
        RECT 82.150 210.905 82.580 211.265 ;
        RECT 83.160 211.075 83.890 211.445 ;
        RECT 82.150 210.715 83.890 210.905 ;
        RECT 82.150 210.485 82.370 210.715 ;
        RECT 81.305 209.685 81.645 210.365 ;
        RECT 80.895 209.485 81.645 209.685 ;
        RECT 81.825 210.185 82.370 210.485 ;
        RECT 80.895 209.095 81.135 209.485 ;
        RECT 81.305 208.895 81.655 209.305 ;
        RECT 81.825 209.075 82.155 210.185 ;
        RECT 82.540 209.915 82.965 210.535 ;
        RECT 83.160 209.915 83.420 210.535 ;
        RECT 83.630 210.205 83.890 210.715 ;
        RECT 82.325 209.545 83.350 209.745 ;
        RECT 82.325 209.075 82.505 209.545 ;
        RECT 82.675 208.895 83.005 209.375 ;
        RECT 83.180 209.075 83.350 209.545 ;
        RECT 83.615 208.895 83.900 210.035 ;
        RECT 84.090 209.075 84.370 211.265 ;
        RECT 84.555 210.770 84.815 211.275 ;
        RECT 84.995 211.065 85.325 211.445 ;
        RECT 85.505 210.895 85.675 211.275 ;
        RECT 84.555 209.970 84.735 210.770 ;
        RECT 85.010 210.725 85.675 210.895 ;
        RECT 85.010 210.470 85.180 210.725 ;
        RECT 85.935 210.695 87.145 211.445 ;
        RECT 84.905 210.140 85.180 210.470 ;
        RECT 85.405 210.175 85.745 210.545 ;
        RECT 85.010 209.995 85.180 210.140 ;
        RECT 84.555 209.065 84.825 209.970 ;
        RECT 85.010 209.825 85.685 209.995 ;
        RECT 84.995 208.895 85.325 209.655 ;
        RECT 85.505 209.065 85.685 209.825 ;
        RECT 85.935 209.985 86.455 210.525 ;
        RECT 86.625 210.155 87.145 210.695 ;
        RECT 85.935 208.895 87.145 209.985 ;
        RECT 15.930 208.725 87.230 208.895 ;
        RECT 16.015 207.635 17.225 208.725 ;
        RECT 16.015 206.925 16.535 207.465 ;
        RECT 16.705 207.095 17.225 207.635 ;
        RECT 18.315 208.005 18.775 208.555 ;
        RECT 18.965 208.005 19.295 208.725 ;
        RECT 16.015 206.175 17.225 206.925 ;
        RECT 18.315 206.635 18.565 208.005 ;
        RECT 19.495 207.835 19.795 208.385 ;
        RECT 19.965 208.055 20.245 208.725 ;
        RECT 18.855 207.665 19.795 207.835 ;
        RECT 18.855 207.415 19.025 207.665 ;
        RECT 20.165 207.415 20.430 207.775 ;
        RECT 20.620 207.575 20.880 208.725 ;
        RECT 21.055 207.650 21.310 208.555 ;
        RECT 21.480 207.965 21.810 208.725 ;
        RECT 22.025 207.795 22.195 208.555 ;
        RECT 22.655 208.055 22.935 208.725 ;
        RECT 18.735 207.085 19.025 207.415 ;
        RECT 19.195 207.165 19.535 207.415 ;
        RECT 19.755 207.165 20.430 207.415 ;
        RECT 18.855 206.995 19.025 207.085 ;
        RECT 18.855 206.805 20.245 206.995 ;
        RECT 18.315 206.345 18.875 206.635 ;
        RECT 19.045 206.175 19.295 206.635 ;
        RECT 19.915 206.445 20.245 206.805 ;
        RECT 20.620 206.175 20.880 207.015 ;
        RECT 21.055 206.920 21.225 207.650 ;
        RECT 21.480 207.625 22.195 207.795 ;
        RECT 23.105 207.835 23.405 208.385 ;
        RECT 23.605 208.005 23.935 208.725 ;
        RECT 24.125 208.005 24.585 208.555 ;
        RECT 21.480 207.415 21.650 207.625 ;
        RECT 21.395 207.085 21.650 207.415 ;
        RECT 21.055 206.345 21.310 206.920 ;
        RECT 21.480 206.895 21.650 207.085 ;
        RECT 21.930 207.075 22.285 207.445 ;
        RECT 22.470 207.415 22.735 207.775 ;
        RECT 23.105 207.665 24.045 207.835 ;
        RECT 23.875 207.415 24.045 207.665 ;
        RECT 22.470 207.165 23.145 207.415 ;
        RECT 23.365 207.165 23.705 207.415 ;
        RECT 23.875 207.085 24.165 207.415 ;
        RECT 23.875 206.995 24.045 207.085 ;
        RECT 21.480 206.725 22.195 206.895 ;
        RECT 21.480 206.175 21.810 206.555 ;
        RECT 22.025 206.345 22.195 206.725 ;
        RECT 22.655 206.805 24.045 206.995 ;
        RECT 22.655 206.445 22.985 206.805 ;
        RECT 24.335 206.635 24.585 208.005 ;
        RECT 24.755 207.665 25.070 208.725 ;
        RECT 25.700 208.220 26.315 208.725 ;
        RECT 24.815 206.835 25.080 207.415 ;
        RECT 25.250 207.335 25.525 207.995 ;
        RECT 25.720 207.685 25.955 208.050 ;
        RECT 26.125 208.045 26.315 208.220 ;
        RECT 26.485 208.215 26.960 208.555 ;
        RECT 26.125 207.855 26.455 208.045 ;
        RECT 26.680 207.685 26.870 207.980 ;
        RECT 27.130 207.880 27.345 208.725 ;
        RECT 27.545 207.885 27.830 208.555 ;
        RECT 25.720 207.515 27.490 207.685 ;
        RECT 25.250 207.105 26.085 207.335 ;
        RECT 23.605 206.175 23.855 206.635 ;
        RECT 24.025 206.345 24.585 206.635 ;
        RECT 24.755 206.175 25.025 206.665 ;
        RECT 25.250 206.395 25.525 207.105 ;
        RECT 26.255 206.660 26.510 207.515 ;
        RECT 25.725 206.395 26.510 206.660 ;
        RECT 26.680 206.855 27.090 207.335 ;
        RECT 27.260 207.085 27.490 207.515 ;
        RECT 27.660 207.535 27.830 207.885 ;
        RECT 28.000 207.715 28.265 208.725 ;
        RECT 28.895 207.560 29.185 208.725 ;
        RECT 29.820 207.580 30.115 208.725 ;
        RECT 27.660 207.015 28.265 207.535 ;
        RECT 26.680 206.395 26.890 206.855 ;
        RECT 27.660 206.805 27.830 207.015 ;
        RECT 27.080 206.175 27.410 206.670 ;
        RECT 27.585 206.345 27.830 206.805 ;
        RECT 28.000 206.175 28.265 206.835 ;
        RECT 28.895 206.175 29.185 206.900 ;
        RECT 29.820 206.175 30.115 206.995 ;
        RECT 30.285 206.725 30.515 208.425 ;
        RECT 30.730 207.920 30.985 208.725 ;
        RECT 31.185 208.110 31.515 208.555 ;
        RECT 31.685 208.280 31.960 208.725 ;
        RECT 32.195 208.110 32.525 208.555 ;
        RECT 31.185 207.930 32.525 208.110 ;
        RECT 32.985 207.750 33.315 208.415 ;
        RECT 33.515 207.925 33.845 208.725 ;
        RECT 30.730 207.580 33.315 207.750 ;
        RECT 34.020 207.585 34.355 208.555 ;
        RECT 34.525 207.925 34.855 208.725 ;
        RECT 35.255 207.755 35.505 208.555 ;
        RECT 35.690 208.005 36.020 208.725 ;
        RECT 36.240 207.755 36.490 208.555 ;
        RECT 36.665 208.345 36.995 208.725 ;
        RECT 34.535 207.585 36.590 207.755 ;
        RECT 30.730 206.965 31.040 207.580 ;
        RECT 34.020 207.365 34.195 207.585 ;
        RECT 34.535 207.405 34.760 207.585 ;
        RECT 31.210 207.135 31.540 207.365 ;
        RECT 31.710 207.135 32.180 207.365 ;
        RECT 32.350 207.195 32.805 207.365 ;
        RECT 32.350 207.135 32.800 207.195 ;
        RECT 32.990 207.135 33.325 207.365 ;
        RECT 34.015 207.195 34.195 207.365 ;
        RECT 30.730 206.785 33.315 206.965 ;
        RECT 30.285 206.345 30.505 206.725 ;
        RECT 30.675 206.175 31.525 206.535 ;
        RECT 32.005 206.365 32.335 206.785 ;
        RECT 32.540 206.175 32.815 206.615 ;
        RECT 32.985 206.365 33.315 206.785 ;
        RECT 33.505 206.175 33.835 206.900 ;
        RECT 34.020 206.895 34.195 207.195 ;
        RECT 34.365 207.165 34.760 207.405 ;
        RECT 34.020 206.430 34.355 206.895 ;
        RECT 34.025 206.385 34.355 206.430 ;
        RECT 34.525 206.175 34.760 206.980 ;
        RECT 34.930 206.505 35.190 207.415 ;
        RECT 35.500 207.395 35.670 207.415 ;
        RECT 35.370 206.505 35.670 207.395 ;
        RECT 35.845 206.510 36.200 207.415 ;
        RECT 36.420 206.675 36.590 207.585 ;
        RECT 36.760 206.845 36.965 208.165 ;
        RECT 37.265 207.980 37.535 208.725 ;
        RECT 38.165 208.720 44.440 208.725 ;
        RECT 37.705 207.810 37.995 208.550 ;
        RECT 38.165 207.995 38.420 208.720 ;
        RECT 38.605 207.825 38.865 208.550 ;
        RECT 39.035 207.995 39.280 208.720 ;
        RECT 39.465 207.825 39.725 208.550 ;
        RECT 39.895 207.995 40.140 208.720 ;
        RECT 40.325 207.825 40.585 208.550 ;
        RECT 40.755 207.995 41.000 208.720 ;
        RECT 41.170 207.825 41.430 208.550 ;
        RECT 41.600 207.995 41.860 208.720 ;
        RECT 42.030 207.825 42.290 208.550 ;
        RECT 42.460 207.995 42.720 208.720 ;
        RECT 42.890 207.825 43.150 208.550 ;
        RECT 43.320 207.995 43.580 208.720 ;
        RECT 43.750 207.825 44.010 208.550 ;
        RECT 44.180 207.925 44.440 208.720 ;
        RECT 38.605 207.810 44.010 207.825 ;
        RECT 37.265 207.585 44.010 207.810 ;
        RECT 37.265 206.995 38.430 207.585 ;
        RECT 44.610 207.415 44.860 208.550 ;
        RECT 45.040 207.915 45.300 208.725 ;
        RECT 45.475 207.415 45.720 208.555 ;
        RECT 45.900 207.915 46.195 208.725 ;
        RECT 46.465 207.715 46.635 208.555 ;
        RECT 46.805 208.385 47.975 208.555 ;
        RECT 46.805 207.885 47.135 208.385 ;
        RECT 47.645 208.345 47.975 208.385 ;
        RECT 48.165 208.305 48.520 208.725 ;
        RECT 47.305 208.125 47.535 208.215 ;
        RECT 48.690 208.125 48.940 208.555 ;
        RECT 47.305 207.885 48.940 208.125 ;
        RECT 49.110 207.965 49.440 208.725 ;
        RECT 49.610 207.885 49.865 208.555 ;
        RECT 46.465 207.545 49.525 207.715 ;
        RECT 38.600 207.165 45.720 207.415 ;
        RECT 37.265 206.825 44.010 206.995 ;
        RECT 36.420 206.345 36.915 206.675 ;
        RECT 37.265 206.175 37.565 206.655 ;
        RECT 37.735 206.370 37.995 206.825 ;
        RECT 38.165 206.175 38.425 206.655 ;
        RECT 38.605 206.370 38.865 206.825 ;
        RECT 39.035 206.175 39.285 206.655 ;
        RECT 39.465 206.370 39.725 206.825 ;
        RECT 39.895 206.175 40.145 206.655 ;
        RECT 40.325 206.370 40.585 206.825 ;
        RECT 40.755 206.175 41.000 206.655 ;
        RECT 41.170 206.370 41.445 206.825 ;
        RECT 41.615 206.175 41.860 206.655 ;
        RECT 42.030 206.370 42.290 206.825 ;
        RECT 42.460 206.175 42.720 206.655 ;
        RECT 42.890 206.370 43.150 206.825 ;
        RECT 43.320 206.175 43.580 206.655 ;
        RECT 43.750 206.370 44.010 206.825 ;
        RECT 44.180 206.175 44.440 206.735 ;
        RECT 44.610 206.355 44.860 207.165 ;
        RECT 45.040 206.175 45.300 206.700 ;
        RECT 45.470 206.355 45.720 207.165 ;
        RECT 45.890 206.855 46.205 207.415 ;
        RECT 46.375 207.165 46.730 207.375 ;
        RECT 46.900 207.165 47.345 207.365 ;
        RECT 47.515 207.165 47.990 207.365 ;
        RECT 46.465 206.825 47.530 206.995 ;
        RECT 45.900 206.175 46.205 206.685 ;
        RECT 46.465 206.345 46.635 206.825 ;
        RECT 46.805 206.175 47.135 206.655 ;
        RECT 47.360 206.595 47.530 206.825 ;
        RECT 47.710 206.765 47.990 207.165 ;
        RECT 48.260 207.165 48.590 207.365 ;
        RECT 48.760 207.165 49.125 207.365 ;
        RECT 48.260 206.765 48.545 207.165 ;
        RECT 49.355 206.995 49.525 207.545 ;
        RECT 48.725 206.825 49.525 206.995 ;
        RECT 48.725 206.595 48.895 206.825 ;
        RECT 49.695 206.755 49.865 207.885 ;
        RECT 50.035 207.535 50.205 208.725 ;
        RECT 50.525 207.750 50.855 208.415 ;
        RECT 51.315 208.110 51.645 208.555 ;
        RECT 51.880 208.280 52.155 208.725 ;
        RECT 52.325 208.110 52.655 208.555 ;
        RECT 51.315 207.930 52.655 208.110 ;
        RECT 52.855 207.920 53.110 208.725 ;
        RECT 50.525 207.580 53.110 207.750 ;
        RECT 50.515 207.135 50.850 207.365 ;
        RECT 51.035 207.195 51.490 207.365 ;
        RECT 51.040 207.135 51.490 207.195 ;
        RECT 51.660 207.135 52.130 207.365 ;
        RECT 52.300 207.135 52.630 207.365 ;
        RECT 49.680 206.685 49.865 206.755 ;
        RECT 49.655 206.675 49.865 206.685 ;
        RECT 47.360 206.345 48.895 206.595 ;
        RECT 49.065 206.175 49.395 206.655 ;
        RECT 49.610 206.345 49.865 206.675 ;
        RECT 50.035 206.175 50.205 207.070 ;
        RECT 52.800 206.965 53.110 207.580 ;
        RECT 50.525 206.785 53.110 206.965 ;
        RECT 50.525 206.365 50.855 206.785 ;
        RECT 51.025 206.175 51.300 206.615 ;
        RECT 51.505 206.365 51.835 206.785 ;
        RECT 53.325 206.725 53.555 208.425 ;
        RECT 53.725 207.580 54.020 208.725 ;
        RECT 54.655 207.560 54.945 208.725 ;
        RECT 55.115 207.755 55.425 208.555 ;
        RECT 55.595 207.925 55.905 208.725 ;
        RECT 56.075 208.095 56.335 208.555 ;
        RECT 56.505 208.265 56.760 208.725 ;
        RECT 56.935 208.095 57.195 208.555 ;
        RECT 56.075 207.925 57.195 208.095 ;
        RECT 55.115 207.585 56.145 207.755 ;
        RECT 52.315 206.175 53.165 206.535 ;
        RECT 53.335 206.345 53.555 206.725 ;
        RECT 53.725 206.175 54.020 206.995 ;
        RECT 54.655 206.175 54.945 206.900 ;
        RECT 55.115 206.675 55.285 207.585 ;
        RECT 55.455 206.845 55.805 207.415 ;
        RECT 55.975 207.335 56.145 207.585 ;
        RECT 56.935 207.675 57.195 207.925 ;
        RECT 57.365 207.855 57.650 208.725 ;
        RECT 57.875 208.130 58.310 208.555 ;
        RECT 58.480 208.300 58.865 208.725 ;
        RECT 57.875 207.960 58.865 208.130 ;
        RECT 56.935 207.505 57.690 207.675 ;
        RECT 55.975 207.165 57.115 207.335 ;
        RECT 57.285 206.995 57.690 207.505 ;
        RECT 57.875 207.085 58.360 207.790 ;
        RECT 58.530 207.415 58.865 207.960 ;
        RECT 59.035 207.765 59.460 208.555 ;
        RECT 59.630 208.130 59.905 208.555 ;
        RECT 60.075 208.300 60.460 208.725 ;
        RECT 59.630 207.935 60.460 208.130 ;
        RECT 59.035 207.585 59.940 207.765 ;
        RECT 58.530 207.085 58.940 207.415 ;
        RECT 59.110 207.085 59.940 207.585 ;
        RECT 60.110 207.415 60.460 207.935 ;
        RECT 60.630 207.765 60.875 208.555 ;
        RECT 61.065 208.130 61.320 208.555 ;
        RECT 61.490 208.300 61.875 208.725 ;
        RECT 61.065 207.935 61.875 208.130 ;
        RECT 60.630 207.585 61.355 207.765 ;
        RECT 60.110 207.085 60.535 207.415 ;
        RECT 60.705 207.085 61.355 207.585 ;
        RECT 61.525 207.415 61.875 207.935 ;
        RECT 62.045 207.585 62.305 208.555 ;
        RECT 62.485 207.915 62.780 208.725 ;
        RECT 61.525 207.085 61.950 207.415 ;
        RECT 56.040 206.825 57.690 206.995 ;
        RECT 58.530 206.915 58.865 207.085 ;
        RECT 59.110 206.915 59.460 207.085 ;
        RECT 60.110 206.915 60.460 207.085 ;
        RECT 60.705 206.915 60.875 207.085 ;
        RECT 61.525 206.915 61.875 207.085 ;
        RECT 62.120 206.915 62.305 207.585 ;
        RECT 62.960 207.415 63.205 208.555 ;
        RECT 63.380 207.915 63.640 208.725 ;
        RECT 64.240 208.720 70.515 208.725 ;
        RECT 63.820 207.415 64.070 208.550 ;
        RECT 64.240 207.925 64.500 208.720 ;
        RECT 64.670 207.825 64.930 208.550 ;
        RECT 65.100 207.995 65.360 208.720 ;
        RECT 65.530 207.825 65.790 208.550 ;
        RECT 65.960 207.995 66.220 208.720 ;
        RECT 66.390 207.825 66.650 208.550 ;
        RECT 66.820 207.995 67.080 208.720 ;
        RECT 67.250 207.825 67.510 208.550 ;
        RECT 67.680 207.995 67.925 208.720 ;
        RECT 68.095 207.825 68.355 208.550 ;
        RECT 68.540 207.995 68.785 208.720 ;
        RECT 68.955 207.825 69.215 208.550 ;
        RECT 69.400 207.995 69.645 208.720 ;
        RECT 69.815 207.825 70.075 208.550 ;
        RECT 70.260 207.995 70.515 208.720 ;
        RECT 64.670 207.810 70.075 207.825 ;
        RECT 70.685 207.810 70.975 208.550 ;
        RECT 71.145 207.980 71.415 208.725 ;
        RECT 71.695 208.135 71.935 208.525 ;
        RECT 72.105 208.315 72.455 208.725 ;
        RECT 71.695 207.935 72.445 208.135 ;
        RECT 64.670 207.585 71.415 207.810 ;
        RECT 55.115 206.345 55.415 206.675 ;
        RECT 55.585 206.175 55.860 206.655 ;
        RECT 56.040 206.435 56.335 206.825 ;
        RECT 56.505 206.175 56.760 206.655 ;
        RECT 56.935 206.435 57.195 206.825 ;
        RECT 57.875 206.745 58.865 206.915 ;
        RECT 57.365 206.175 57.645 206.655 ;
        RECT 57.875 206.345 58.310 206.745 ;
        RECT 58.480 206.175 58.865 206.575 ;
        RECT 59.035 206.345 59.460 206.915 ;
        RECT 59.650 206.745 60.460 206.915 ;
        RECT 59.650 206.345 59.905 206.745 ;
        RECT 60.075 206.175 60.460 206.575 ;
        RECT 60.630 206.345 60.875 206.915 ;
        RECT 61.065 206.745 61.875 206.915 ;
        RECT 61.065 206.345 61.320 206.745 ;
        RECT 61.490 206.175 61.875 206.575 ;
        RECT 62.045 206.345 62.305 206.915 ;
        RECT 62.475 206.855 62.790 207.415 ;
        RECT 62.960 207.165 70.080 207.415 ;
        RECT 62.475 206.175 62.780 206.685 ;
        RECT 62.960 206.355 63.210 207.165 ;
        RECT 63.380 206.175 63.640 206.700 ;
        RECT 63.820 206.355 64.070 207.165 ;
        RECT 70.250 206.995 71.415 207.585 ;
        RECT 64.670 206.825 71.415 206.995 ;
        RECT 64.240 206.175 64.500 206.735 ;
        RECT 64.670 206.370 64.930 206.825 ;
        RECT 65.100 206.175 65.360 206.655 ;
        RECT 65.530 206.370 65.790 206.825 ;
        RECT 65.960 206.175 66.220 206.655 ;
        RECT 66.390 206.370 66.650 206.825 ;
        RECT 66.820 206.175 67.065 206.655 ;
        RECT 67.235 206.370 67.510 206.825 ;
        RECT 67.680 206.175 67.925 206.655 ;
        RECT 68.095 206.370 68.355 206.825 ;
        RECT 68.535 206.175 68.785 206.655 ;
        RECT 68.955 206.370 69.215 206.825 ;
        RECT 69.395 206.175 69.645 206.655 ;
        RECT 69.815 206.370 70.075 206.825 ;
        RECT 70.255 206.175 70.515 206.655 ;
        RECT 70.685 206.370 70.945 206.825 ;
        RECT 71.115 206.175 71.415 206.655 ;
        RECT 71.695 206.415 71.925 207.755 ;
        RECT 72.105 207.255 72.445 207.935 ;
        RECT 72.625 207.435 72.955 208.545 ;
        RECT 73.125 208.075 73.305 208.545 ;
        RECT 73.475 208.245 73.805 208.725 ;
        RECT 73.980 208.075 74.150 208.545 ;
        RECT 73.125 207.875 74.150 208.075 ;
        RECT 72.105 206.355 72.335 207.255 ;
        RECT 72.625 207.135 73.170 207.435 ;
        RECT 72.535 206.175 72.780 206.955 ;
        RECT 72.950 206.905 73.170 207.135 ;
        RECT 73.340 207.085 73.765 207.705 ;
        RECT 73.960 207.085 74.220 207.705 ;
        RECT 74.415 207.585 74.700 208.725 ;
        RECT 74.430 206.905 74.690 207.415 ;
        RECT 72.950 206.715 74.690 206.905 ;
        RECT 72.950 206.355 73.380 206.715 ;
        RECT 73.960 206.175 74.690 206.545 ;
        RECT 74.890 206.355 75.170 208.545 ;
        RECT 75.375 208.135 75.615 208.525 ;
        RECT 75.785 208.315 76.135 208.725 ;
        RECT 75.375 207.935 76.125 208.135 ;
        RECT 75.375 206.415 75.605 207.755 ;
        RECT 75.785 207.255 76.125 207.935 ;
        RECT 76.305 207.435 76.635 208.545 ;
        RECT 76.805 208.075 76.985 208.545 ;
        RECT 77.155 208.245 77.485 208.725 ;
        RECT 77.660 208.075 77.830 208.545 ;
        RECT 76.805 207.875 77.830 208.075 ;
        RECT 75.785 206.355 76.015 207.255 ;
        RECT 76.305 207.135 76.850 207.435 ;
        RECT 76.215 206.175 76.460 206.955 ;
        RECT 76.630 206.905 76.850 207.135 ;
        RECT 77.020 207.085 77.445 207.705 ;
        RECT 77.640 207.085 77.900 207.705 ;
        RECT 78.095 207.585 78.380 208.725 ;
        RECT 78.110 206.905 78.370 207.415 ;
        RECT 76.630 206.715 78.370 206.905 ;
        RECT 76.630 206.355 77.060 206.715 ;
        RECT 77.640 206.175 78.370 206.545 ;
        RECT 78.570 206.355 78.850 208.545 ;
        RECT 79.095 207.585 79.305 208.725 ;
        RECT 79.475 207.575 79.805 208.555 ;
        RECT 79.975 207.585 80.205 208.725 ;
        RECT 79.095 206.175 79.305 206.995 ;
        RECT 79.475 206.975 79.725 207.575 ;
        RECT 80.415 207.560 80.705 208.725 ;
        RECT 80.895 208.135 81.135 208.525 ;
        RECT 81.305 208.315 81.655 208.725 ;
        RECT 80.895 207.935 81.645 208.135 ;
        RECT 79.895 207.165 80.225 207.415 ;
        RECT 79.475 206.345 79.805 206.975 ;
        RECT 79.975 206.175 80.205 206.995 ;
        RECT 80.415 206.175 80.705 206.900 ;
        RECT 80.895 206.415 81.125 207.755 ;
        RECT 81.305 207.255 81.645 207.935 ;
        RECT 81.825 207.435 82.155 208.545 ;
        RECT 82.325 208.075 82.505 208.545 ;
        RECT 82.675 208.245 83.005 208.725 ;
        RECT 83.180 208.075 83.350 208.545 ;
        RECT 82.325 207.875 83.350 208.075 ;
        RECT 81.305 206.355 81.535 207.255 ;
        RECT 81.825 207.135 82.370 207.435 ;
        RECT 81.735 206.175 81.980 206.955 ;
        RECT 82.150 206.905 82.370 207.135 ;
        RECT 82.540 207.085 82.965 207.705 ;
        RECT 83.160 207.085 83.420 207.705 ;
        RECT 83.615 207.585 83.900 208.725 ;
        RECT 83.630 206.905 83.890 207.415 ;
        RECT 82.150 206.715 83.890 206.905 ;
        RECT 82.150 206.355 82.580 206.715 ;
        RECT 83.160 206.175 83.890 206.545 ;
        RECT 84.090 206.355 84.370 208.545 ;
        RECT 84.555 207.650 84.825 208.555 ;
        RECT 84.995 207.965 85.325 208.725 ;
        RECT 85.505 207.795 85.675 208.555 ;
        RECT 84.555 206.850 84.725 207.650 ;
        RECT 85.010 207.625 85.675 207.795 ;
        RECT 85.935 207.635 87.145 208.725 ;
        RECT 85.010 207.480 85.180 207.625 ;
        RECT 84.895 207.150 85.180 207.480 ;
        RECT 85.010 206.895 85.180 207.150 ;
        RECT 85.415 207.075 85.745 207.445 ;
        RECT 85.935 207.095 86.455 207.635 ;
        RECT 86.625 206.925 87.145 207.465 ;
        RECT 84.555 206.345 84.815 206.850 ;
        RECT 85.010 206.725 85.675 206.895 ;
        RECT 84.995 206.175 85.325 206.555 ;
        RECT 85.505 206.345 85.675 206.725 ;
        RECT 85.935 206.175 87.145 206.925 ;
        RECT 15.930 206.005 87.230 206.175 ;
        RECT 16.015 205.255 17.225 206.005 ;
        RECT 16.015 204.715 16.535 205.255 ;
        RECT 17.400 205.165 17.660 206.005 ;
        RECT 17.835 205.260 18.090 205.835 ;
        RECT 18.260 205.625 18.590 206.005 ;
        RECT 18.805 205.455 18.975 205.835 ;
        RECT 18.260 205.285 18.975 205.455 ;
        RECT 16.705 204.545 17.225 205.085 ;
        RECT 16.015 203.455 17.225 204.545 ;
        RECT 17.400 203.455 17.660 204.605 ;
        RECT 17.835 204.530 18.005 205.260 ;
        RECT 18.260 205.095 18.430 205.285 ;
        RECT 19.235 205.205 19.545 206.005 ;
        RECT 19.750 205.205 20.445 205.835 ;
        RECT 20.615 205.205 20.925 206.005 ;
        RECT 21.130 205.205 21.825 205.835 ;
        RECT 22.040 205.545 22.790 205.835 ;
        RECT 23.300 205.545 23.630 206.005 ;
        RECT 18.175 204.765 18.430 205.095 ;
        RECT 18.260 204.555 18.430 204.765 ;
        RECT 18.710 204.735 19.065 205.105 ;
        RECT 19.245 204.765 19.580 205.035 ;
        RECT 19.750 204.605 19.920 205.205 ;
        RECT 21.130 205.155 21.305 205.205 ;
        RECT 20.090 204.765 20.425 205.015 ;
        RECT 20.625 204.765 20.960 205.035 ;
        RECT 21.130 204.605 21.300 205.155 ;
        RECT 21.470 204.765 21.805 205.015 ;
        RECT 17.835 203.625 18.090 204.530 ;
        RECT 18.260 204.385 18.975 204.555 ;
        RECT 18.260 203.455 18.590 204.215 ;
        RECT 18.805 203.625 18.975 204.385 ;
        RECT 19.235 203.455 19.515 204.595 ;
        RECT 19.685 203.625 20.015 204.605 ;
        RECT 20.185 203.455 20.445 204.595 ;
        RECT 20.615 203.455 20.895 204.595 ;
        RECT 21.065 203.625 21.395 204.605 ;
        RECT 21.565 203.455 21.825 204.595 ;
        RECT 22.040 204.255 22.410 205.545 ;
        RECT 23.850 205.355 24.120 205.565 ;
        RECT 22.785 205.185 24.120 205.355 ;
        RECT 24.295 205.345 24.570 206.005 ;
        RECT 24.740 205.375 24.990 205.835 ;
        RECT 25.165 205.510 25.495 206.005 ;
        RECT 22.785 205.015 22.955 205.185 ;
        RECT 24.740 205.165 24.910 205.375 ;
        RECT 25.675 205.340 25.905 205.785 ;
        RECT 22.580 204.765 22.955 205.015 ;
        RECT 23.125 204.775 23.600 205.015 ;
        RECT 23.770 204.775 24.120 205.015 ;
        RECT 22.785 204.595 22.955 204.765 ;
        RECT 24.295 204.645 24.910 205.165 ;
        RECT 25.080 204.665 25.310 205.095 ;
        RECT 25.495 204.845 25.905 205.340 ;
        RECT 26.075 205.520 26.865 205.785 ;
        RECT 26.075 204.665 26.330 205.520 ;
        RECT 27.255 205.375 27.585 205.735 ;
        RECT 28.215 205.545 28.465 206.005 ;
        RECT 28.635 205.545 29.185 205.835 ;
        RECT 26.500 204.845 26.885 205.325 ;
        RECT 27.255 205.185 28.645 205.375 ;
        RECT 28.475 205.095 28.645 205.185 ;
        RECT 27.055 204.765 27.745 205.015 ;
        RECT 27.975 204.765 28.305 205.015 ;
        RECT 28.475 204.765 28.765 205.095 ;
        RECT 22.785 204.425 24.120 204.595 ;
        RECT 23.840 204.265 24.120 204.425 ;
        RECT 22.040 204.085 23.210 204.255 ;
        RECT 22.495 203.455 22.710 203.915 ;
        RECT 22.880 203.625 23.210 204.085 ;
        RECT 23.380 203.455 23.630 204.255 ;
        RECT 24.295 203.455 24.555 204.465 ;
        RECT 24.725 204.295 24.895 204.645 ;
        RECT 25.080 204.495 26.870 204.665 ;
        RECT 24.725 203.625 25.000 204.295 ;
        RECT 25.200 203.455 25.415 204.300 ;
        RECT 25.640 204.200 25.890 204.495 ;
        RECT 26.115 204.135 26.445 204.325 ;
        RECT 25.600 203.625 26.075 203.965 ;
        RECT 26.255 203.960 26.445 204.135 ;
        RECT 26.615 204.130 26.870 204.495 ;
        RECT 27.055 204.325 27.370 204.765 ;
        RECT 28.475 204.515 28.645 204.765 ;
        RECT 27.705 204.345 28.645 204.515 ;
        RECT 26.255 203.455 26.885 203.960 ;
        RECT 27.255 203.455 27.535 204.125 ;
        RECT 27.705 203.795 28.005 204.345 ;
        RECT 28.935 204.175 29.185 205.545 ;
        RECT 29.355 205.205 29.645 206.005 ;
        RECT 29.875 205.525 30.155 206.005 ;
        RECT 30.325 205.355 30.585 205.745 ;
        RECT 30.760 205.525 31.015 206.005 ;
        RECT 31.185 205.355 31.480 205.745 ;
        RECT 31.660 205.525 31.935 206.005 ;
        RECT 32.105 205.505 32.405 205.835 ;
        RECT 32.665 205.525 32.965 206.005 ;
        RECT 29.830 205.185 31.480 205.355 ;
        RECT 29.830 204.675 30.235 205.185 ;
        RECT 30.405 204.845 31.545 205.015 ;
        RECT 28.215 203.455 28.545 204.175 ;
        RECT 28.735 203.625 29.185 204.175 ;
        RECT 29.355 203.455 29.645 204.595 ;
        RECT 29.830 204.505 30.585 204.675 ;
        RECT 29.870 203.455 30.155 204.325 ;
        RECT 30.325 204.255 30.585 204.505 ;
        RECT 31.375 204.595 31.545 204.845 ;
        RECT 31.715 204.765 32.065 205.335 ;
        RECT 32.235 204.595 32.405 205.505 ;
        RECT 33.135 205.355 33.395 205.810 ;
        RECT 33.565 205.525 33.825 206.005 ;
        RECT 34.005 205.355 34.265 205.810 ;
        RECT 34.435 205.525 34.685 206.005 ;
        RECT 34.865 205.355 35.125 205.810 ;
        RECT 35.295 205.525 35.545 206.005 ;
        RECT 35.725 205.355 35.985 205.810 ;
        RECT 36.155 205.525 36.400 206.005 ;
        RECT 36.570 205.355 36.845 205.810 ;
        RECT 37.015 205.525 37.260 206.005 ;
        RECT 37.430 205.355 37.690 205.810 ;
        RECT 37.860 205.525 38.120 206.005 ;
        RECT 38.290 205.355 38.550 205.810 ;
        RECT 38.720 205.525 38.980 206.005 ;
        RECT 39.150 205.355 39.410 205.810 ;
        RECT 39.580 205.445 39.840 206.005 ;
        RECT 31.375 204.425 32.405 204.595 ;
        RECT 30.325 204.085 31.445 204.255 ;
        RECT 30.325 203.625 30.585 204.085 ;
        RECT 30.760 203.455 31.015 203.915 ;
        RECT 31.185 203.625 31.445 204.085 ;
        RECT 31.615 203.455 31.925 204.255 ;
        RECT 32.095 203.625 32.405 204.425 ;
        RECT 32.665 205.185 39.410 205.355 ;
        RECT 32.665 204.595 33.830 205.185 ;
        RECT 40.010 205.015 40.260 205.825 ;
        RECT 40.440 205.480 40.700 206.005 ;
        RECT 40.870 205.015 41.120 205.825 ;
        RECT 41.300 205.495 41.605 206.005 ;
        RECT 34.000 204.765 41.120 205.015 ;
        RECT 41.290 204.765 41.605 205.325 ;
        RECT 41.775 205.280 42.065 206.005 ;
        RECT 43.155 205.495 43.460 206.005 ;
        RECT 43.155 204.765 43.470 205.325 ;
        RECT 43.640 205.015 43.890 205.825 ;
        RECT 44.060 205.480 44.320 206.005 ;
        RECT 44.500 205.015 44.750 205.825 ;
        RECT 44.920 205.445 45.180 206.005 ;
        RECT 45.350 205.355 45.610 205.810 ;
        RECT 45.780 205.525 46.040 206.005 ;
        RECT 46.210 205.355 46.470 205.810 ;
        RECT 46.640 205.525 46.900 206.005 ;
        RECT 47.070 205.355 47.330 205.810 ;
        RECT 47.500 205.525 47.745 206.005 ;
        RECT 47.915 205.355 48.190 205.810 ;
        RECT 48.360 205.525 48.605 206.005 ;
        RECT 48.775 205.355 49.035 205.810 ;
        RECT 49.215 205.525 49.465 206.005 ;
        RECT 49.635 205.355 49.895 205.810 ;
        RECT 50.075 205.525 50.325 206.005 ;
        RECT 50.495 205.355 50.755 205.810 ;
        RECT 50.935 205.525 51.195 206.005 ;
        RECT 51.365 205.355 51.625 205.810 ;
        RECT 51.795 205.525 52.095 206.005 ;
        RECT 52.445 205.525 52.745 206.005 ;
        RECT 52.915 205.355 53.175 205.810 ;
        RECT 53.345 205.525 53.605 206.005 ;
        RECT 53.785 205.355 54.045 205.810 ;
        RECT 54.215 205.525 54.465 206.005 ;
        RECT 54.645 205.355 54.905 205.810 ;
        RECT 55.075 205.525 55.325 206.005 ;
        RECT 55.505 205.355 55.765 205.810 ;
        RECT 55.935 205.525 56.180 206.005 ;
        RECT 56.350 205.355 56.625 205.810 ;
        RECT 56.795 205.525 57.040 206.005 ;
        RECT 57.210 205.355 57.470 205.810 ;
        RECT 57.640 205.525 57.900 206.005 ;
        RECT 58.070 205.355 58.330 205.810 ;
        RECT 58.500 205.525 58.760 206.005 ;
        RECT 58.930 205.355 59.190 205.810 ;
        RECT 59.360 205.445 59.620 206.005 ;
        RECT 45.350 205.185 52.095 205.355 ;
        RECT 43.640 204.765 50.760 205.015 ;
        RECT 32.665 204.370 39.410 204.595 ;
        RECT 32.665 203.455 32.935 204.200 ;
        RECT 33.105 203.630 33.395 204.370 ;
        RECT 34.005 204.355 39.410 204.370 ;
        RECT 33.565 203.460 33.820 204.185 ;
        RECT 34.005 203.630 34.265 204.355 ;
        RECT 34.435 203.460 34.680 204.185 ;
        RECT 34.865 203.630 35.125 204.355 ;
        RECT 35.295 203.460 35.540 204.185 ;
        RECT 35.725 203.630 35.985 204.355 ;
        RECT 36.155 203.460 36.400 204.185 ;
        RECT 36.570 203.630 36.830 204.355 ;
        RECT 37.000 203.460 37.260 204.185 ;
        RECT 37.430 203.630 37.690 204.355 ;
        RECT 37.860 203.460 38.120 204.185 ;
        RECT 38.290 203.630 38.550 204.355 ;
        RECT 38.720 203.460 38.980 204.185 ;
        RECT 39.150 203.630 39.410 204.355 ;
        RECT 39.580 203.460 39.840 204.255 ;
        RECT 40.010 203.630 40.260 204.765 ;
        RECT 33.565 203.455 39.840 203.460 ;
        RECT 40.440 203.455 40.700 204.265 ;
        RECT 40.875 203.625 41.120 204.765 ;
        RECT 41.300 203.455 41.595 204.265 ;
        RECT 41.775 203.455 42.065 204.620 ;
        RECT 43.165 203.455 43.460 204.265 ;
        RECT 43.640 203.625 43.885 204.765 ;
        RECT 44.060 203.455 44.320 204.265 ;
        RECT 44.500 203.630 44.750 204.765 ;
        RECT 50.930 204.595 52.095 205.185 ;
        RECT 45.350 204.370 52.095 204.595 ;
        RECT 52.445 205.185 59.190 205.355 ;
        RECT 52.445 204.595 53.610 205.185 ;
        RECT 59.790 205.015 60.040 205.825 ;
        RECT 60.220 205.480 60.480 206.005 ;
        RECT 60.650 205.015 60.900 205.825 ;
        RECT 61.080 205.495 61.385 206.005 ;
        RECT 53.780 204.765 60.900 205.015 ;
        RECT 61.070 204.765 61.385 205.325 ;
        RECT 61.565 205.195 61.835 206.005 ;
        RECT 62.005 205.195 62.335 205.835 ;
        RECT 62.505 205.195 62.745 206.005 ;
        RECT 62.940 205.625 64.955 205.795 ;
        RECT 65.145 205.625 65.475 206.005 ;
        RECT 62.940 205.305 63.195 205.625 ;
        RECT 61.555 204.765 61.905 205.015 ;
        RECT 52.445 204.370 59.190 204.595 ;
        RECT 45.350 204.355 50.755 204.370 ;
        RECT 44.920 203.460 45.180 204.255 ;
        RECT 45.350 203.630 45.610 204.355 ;
        RECT 45.780 203.460 46.040 204.185 ;
        RECT 46.210 203.630 46.470 204.355 ;
        RECT 46.640 203.460 46.900 204.185 ;
        RECT 47.070 203.630 47.330 204.355 ;
        RECT 47.500 203.460 47.760 204.185 ;
        RECT 47.930 203.630 48.190 204.355 ;
        RECT 48.360 203.460 48.605 204.185 ;
        RECT 48.775 203.630 49.035 204.355 ;
        RECT 49.220 203.460 49.465 204.185 ;
        RECT 49.635 203.630 49.895 204.355 ;
        RECT 50.080 203.460 50.325 204.185 ;
        RECT 50.495 203.630 50.755 204.355 ;
        RECT 50.940 203.460 51.195 204.185 ;
        RECT 51.365 203.630 51.655 204.370 ;
        RECT 44.920 203.455 51.195 203.460 ;
        RECT 51.825 203.455 52.095 204.200 ;
        RECT 52.445 203.455 52.715 204.200 ;
        RECT 52.885 203.630 53.175 204.370 ;
        RECT 53.785 204.355 59.190 204.370 ;
        RECT 53.345 203.460 53.600 204.185 ;
        RECT 53.785 203.630 54.045 204.355 ;
        RECT 54.215 203.460 54.460 204.185 ;
        RECT 54.645 203.630 54.905 204.355 ;
        RECT 55.075 203.460 55.320 204.185 ;
        RECT 55.505 203.630 55.765 204.355 ;
        RECT 55.935 203.460 56.180 204.185 ;
        RECT 56.350 203.630 56.610 204.355 ;
        RECT 56.780 203.460 57.040 204.185 ;
        RECT 57.210 203.630 57.470 204.355 ;
        RECT 57.640 203.460 57.900 204.185 ;
        RECT 58.070 203.630 58.330 204.355 ;
        RECT 58.500 203.460 58.760 204.185 ;
        RECT 58.930 203.630 59.190 204.355 ;
        RECT 59.360 203.460 59.620 204.255 ;
        RECT 59.790 203.630 60.040 204.765 ;
        RECT 53.345 203.455 59.620 203.460 ;
        RECT 60.220 203.455 60.480 204.265 ;
        RECT 60.655 203.625 60.900 204.765 ;
        RECT 62.075 204.595 62.245 205.195 ;
        RECT 62.415 204.765 62.765 205.015 ;
        RECT 62.940 204.765 63.180 205.095 ;
        RECT 63.365 204.645 63.695 205.455 ;
        RECT 64.205 205.185 65.895 205.455 ;
        RECT 66.065 205.205 66.445 206.005 ;
        RECT 67.535 205.280 67.825 206.005 ;
        RECT 63.920 204.815 65.010 205.015 ;
        RECT 65.320 204.815 66.445 205.015 ;
        RECT 61.080 203.455 61.375 204.265 ;
        RECT 61.565 203.455 61.895 204.595 ;
        RECT 62.075 204.425 62.755 204.595 ;
        RECT 62.425 203.640 62.755 204.425 ;
        RECT 62.940 203.455 63.195 204.595 ;
        RECT 63.365 204.425 65.895 204.645 ;
        RECT 63.365 203.625 63.695 204.425 ;
        RECT 63.865 203.455 64.035 204.255 ;
        RECT 64.205 203.625 64.535 204.425 ;
        RECT 64.705 203.455 65.395 204.255 ;
        RECT 65.565 203.625 65.895 204.425 ;
        RECT 66.065 203.455 66.445 204.645 ;
        RECT 67.535 203.455 67.825 204.620 ;
        RECT 68.010 203.635 68.290 205.825 ;
        RECT 68.490 205.635 69.220 206.005 ;
        RECT 69.800 205.465 70.230 205.825 ;
        RECT 68.490 205.275 70.230 205.465 ;
        RECT 68.490 204.765 68.750 205.275 ;
        RECT 68.480 203.455 68.765 204.595 ;
        RECT 68.960 204.475 69.220 205.095 ;
        RECT 69.415 204.475 69.840 205.095 ;
        RECT 70.010 205.045 70.230 205.275 ;
        RECT 70.400 205.225 70.645 206.005 ;
        RECT 70.010 204.745 70.555 205.045 ;
        RECT 70.845 204.925 71.075 205.825 ;
        RECT 69.030 204.105 70.055 204.305 ;
        RECT 69.030 203.635 69.200 204.105 ;
        RECT 69.375 203.455 69.705 203.935 ;
        RECT 69.875 203.635 70.055 204.105 ;
        RECT 70.225 203.635 70.555 204.745 ;
        RECT 70.735 204.245 71.075 204.925 ;
        RECT 71.255 204.425 71.485 205.765 ;
        RECT 71.715 205.185 71.945 206.005 ;
        RECT 72.115 205.205 72.445 205.835 ;
        RECT 71.695 204.765 72.025 205.015 ;
        RECT 72.195 204.605 72.445 205.205 ;
        RECT 72.615 205.185 72.825 206.005 ;
        RECT 73.145 205.525 73.445 206.005 ;
        RECT 73.615 205.355 73.875 205.810 ;
        RECT 74.045 205.525 74.305 206.005 ;
        RECT 74.485 205.355 74.745 205.810 ;
        RECT 74.915 205.525 75.165 206.005 ;
        RECT 75.345 205.355 75.605 205.810 ;
        RECT 75.775 205.525 76.025 206.005 ;
        RECT 76.205 205.355 76.465 205.810 ;
        RECT 76.635 205.525 76.880 206.005 ;
        RECT 77.050 205.355 77.325 205.810 ;
        RECT 77.495 205.525 77.740 206.005 ;
        RECT 77.910 205.355 78.170 205.810 ;
        RECT 78.340 205.525 78.600 206.005 ;
        RECT 78.770 205.355 79.030 205.810 ;
        RECT 79.200 205.525 79.460 206.005 ;
        RECT 79.630 205.355 79.890 205.810 ;
        RECT 80.060 205.445 80.320 206.005 ;
        RECT 73.145 205.185 79.890 205.355 ;
        RECT 70.735 204.045 71.485 204.245 ;
        RECT 70.725 203.455 71.075 203.865 ;
        RECT 71.245 203.655 71.485 204.045 ;
        RECT 71.715 203.455 71.945 204.595 ;
        RECT 72.115 203.625 72.445 204.605 ;
        RECT 73.145 204.595 74.310 205.185 ;
        RECT 80.490 205.015 80.740 205.825 ;
        RECT 80.920 205.480 81.180 206.005 ;
        RECT 81.350 205.015 81.600 205.825 ;
        RECT 81.780 205.495 82.085 206.005 ;
        RECT 82.255 205.525 82.515 206.005 ;
        RECT 82.685 205.755 82.930 205.835 ;
        RECT 82.685 205.585 83.015 205.755 ;
        RECT 74.480 204.765 81.600 205.015 ;
        RECT 81.770 204.765 82.085 205.325 ;
        RECT 82.300 204.765 82.495 205.335 ;
        RECT 72.615 203.455 72.825 204.595 ;
        RECT 73.145 204.370 79.890 204.595 ;
        RECT 73.145 203.455 73.415 204.200 ;
        RECT 73.585 203.630 73.875 204.370 ;
        RECT 74.485 204.355 79.890 204.370 ;
        RECT 74.045 203.460 74.300 204.185 ;
        RECT 74.485 203.630 74.745 204.355 ;
        RECT 74.915 203.460 75.160 204.185 ;
        RECT 75.345 203.630 75.605 204.355 ;
        RECT 75.775 203.460 76.020 204.185 ;
        RECT 76.205 203.630 76.465 204.355 ;
        RECT 76.635 203.460 76.880 204.185 ;
        RECT 77.050 203.630 77.310 204.355 ;
        RECT 77.480 203.460 77.740 204.185 ;
        RECT 77.910 203.630 78.170 204.355 ;
        RECT 78.340 203.460 78.600 204.185 ;
        RECT 78.770 203.630 79.030 204.355 ;
        RECT 79.200 203.460 79.460 204.185 ;
        RECT 79.630 203.630 79.890 204.355 ;
        RECT 80.060 203.460 80.320 204.255 ;
        RECT 80.490 203.630 80.740 204.765 ;
        RECT 74.045 203.455 80.320 203.460 ;
        RECT 80.920 203.455 81.180 204.265 ;
        RECT 81.355 203.625 81.600 204.765 ;
        RECT 82.685 204.595 82.855 205.585 ;
        RECT 83.215 205.390 83.425 205.675 ;
        RECT 83.690 205.665 83.860 205.690 ;
        RECT 83.690 205.495 83.865 205.665 ;
        RECT 84.105 205.625 84.435 206.005 ;
        RECT 84.625 205.665 84.795 205.835 ;
        RECT 84.205 205.545 84.375 205.625 ;
        RECT 84.615 205.495 84.795 205.665 ;
        RECT 85.045 205.545 85.300 206.005 ;
        RECT 83.690 205.395 83.860 205.495 ;
        RECT 83.035 205.220 83.425 205.390 ;
        RECT 83.595 205.225 83.860 205.395 ;
        RECT 84.625 205.375 84.795 205.495 ;
        RECT 83.035 205.155 83.315 205.220 ;
        RECT 83.035 204.765 83.205 205.155 ;
        RECT 83.595 205.015 83.765 205.225 ;
        RECT 84.120 205.095 84.325 205.330 ;
        RECT 84.625 205.205 85.300 205.375 ;
        RECT 85.935 205.255 87.145 206.005 ;
        RECT 83.435 204.845 83.765 205.015 ;
        RECT 83.595 204.830 83.765 204.845 ;
        RECT 83.995 204.765 84.325 205.095 ;
        RECT 84.505 204.845 84.835 205.015 ;
        RECT 84.665 204.595 84.835 204.845 ;
        RECT 82.345 204.425 84.835 204.595 ;
        RECT 81.780 203.455 82.075 204.265 ;
        RECT 82.345 203.625 82.515 204.425 ;
        RECT 85.045 204.255 85.300 205.205 ;
        RECT 82.745 204.085 84.035 204.255 ;
        RECT 82.805 203.665 83.055 204.085 ;
        RECT 83.245 203.455 83.575 203.915 ;
        RECT 83.785 203.665 84.035 204.085 ;
        RECT 84.205 203.455 84.455 204.255 ;
        RECT 84.625 204.085 85.300 204.255 ;
        RECT 85.935 204.545 86.455 205.085 ;
        RECT 86.625 204.715 87.145 205.255 ;
        RECT 84.625 203.625 84.795 204.085 ;
        RECT 85.005 203.455 85.255 203.915 ;
        RECT 85.935 203.455 87.145 204.545 ;
        RECT 15.930 203.285 87.230 203.455 ;
        RECT 16.015 202.195 17.225 203.285 ;
        RECT 16.015 201.485 16.535 202.025 ;
        RECT 16.705 201.655 17.225 202.195 ;
        RECT 18.405 202.355 18.575 203.115 ;
        RECT 18.790 202.525 19.120 203.285 ;
        RECT 18.405 202.185 19.120 202.355 ;
        RECT 19.290 202.210 19.545 203.115 ;
        RECT 18.315 201.635 18.670 202.005 ;
        RECT 18.950 201.975 19.120 202.185 ;
        RECT 18.950 201.645 19.205 201.975 ;
        RECT 16.015 200.735 17.225 201.485 ;
        RECT 18.950 201.455 19.120 201.645 ;
        RECT 19.375 201.480 19.545 202.210 ;
        RECT 19.720 202.135 19.980 203.285 ;
        RECT 20.160 202.135 20.420 203.285 ;
        RECT 20.595 202.210 20.850 203.115 ;
        RECT 21.020 202.525 21.350 203.285 ;
        RECT 21.565 202.355 21.735 203.115 ;
        RECT 18.405 201.285 19.120 201.455 ;
        RECT 18.405 200.905 18.575 201.285 ;
        RECT 18.790 200.735 19.120 201.115 ;
        RECT 19.290 200.905 19.545 201.480 ;
        RECT 19.720 200.735 19.980 201.575 ;
        RECT 20.160 200.735 20.420 201.575 ;
        RECT 20.595 201.480 20.765 202.210 ;
        RECT 21.020 202.185 21.735 202.355 ;
        RECT 21.020 201.975 21.190 202.185 ;
        RECT 22.915 202.145 23.195 203.285 ;
        RECT 23.365 202.135 23.695 203.115 ;
        RECT 23.865 202.145 24.125 203.285 ;
        RECT 24.495 202.615 24.775 203.285 ;
        RECT 24.945 202.395 25.245 202.945 ;
        RECT 25.445 202.565 25.775 203.285 ;
        RECT 25.965 202.565 26.425 203.115 ;
        RECT 20.935 201.645 21.190 201.975 ;
        RECT 20.595 200.905 20.850 201.480 ;
        RECT 21.020 201.455 21.190 201.645 ;
        RECT 21.470 201.635 21.825 202.005 ;
        RECT 22.925 201.705 23.260 201.975 ;
        RECT 23.430 201.535 23.600 202.135 ;
        RECT 24.310 201.975 24.575 202.335 ;
        RECT 24.945 202.225 25.885 202.395 ;
        RECT 25.715 201.975 25.885 202.225 ;
        RECT 23.770 201.725 24.105 201.975 ;
        RECT 24.310 201.725 24.985 201.975 ;
        RECT 25.205 201.725 25.545 201.975 ;
        RECT 25.715 201.645 26.005 201.975 ;
        RECT 25.715 201.555 25.885 201.645 ;
        RECT 21.020 201.285 21.735 201.455 ;
        RECT 21.020 200.735 21.350 201.115 ;
        RECT 21.565 200.905 21.735 201.285 ;
        RECT 22.915 200.735 23.225 201.535 ;
        RECT 23.430 200.905 24.125 201.535 ;
        RECT 24.495 201.365 25.885 201.555 ;
        RECT 24.495 201.005 24.825 201.365 ;
        RECT 26.175 201.195 26.425 202.565 ;
        RECT 26.615 202.485 26.895 203.285 ;
        RECT 27.095 202.315 27.425 203.115 ;
        RECT 27.625 202.485 27.795 203.285 ;
        RECT 27.965 202.315 28.295 203.115 ;
        RECT 26.595 201.645 26.835 202.315 ;
        RECT 27.015 202.145 28.295 202.315 ;
        RECT 28.465 202.145 28.725 203.285 ;
        RECT 27.015 201.475 27.185 202.145 ;
        RECT 28.895 202.120 29.185 203.285 ;
        RECT 29.355 202.210 29.625 203.115 ;
        RECT 29.795 202.525 30.125 203.285 ;
        RECT 30.305 202.355 30.475 203.115 ;
        RECT 27.355 201.645 27.665 201.975 ;
        RECT 27.835 201.645 28.215 201.975 ;
        RECT 28.415 201.645 28.700 201.975 ;
        RECT 27.460 201.475 27.665 201.645 ;
        RECT 25.445 200.735 25.695 201.195 ;
        RECT 25.865 200.905 26.425 201.195 ;
        RECT 26.595 200.905 27.290 201.475 ;
        RECT 27.460 200.950 27.810 201.475 ;
        RECT 28.000 200.950 28.215 201.645 ;
        RECT 28.385 200.735 28.720 201.475 ;
        RECT 28.895 200.735 29.185 201.460 ;
        RECT 29.355 201.410 29.525 202.210 ;
        RECT 29.810 202.185 30.475 202.355 ;
        RECT 30.755 202.395 31.015 203.105 ;
        RECT 31.185 202.575 31.515 203.285 ;
        RECT 31.685 202.395 31.915 203.105 ;
        RECT 29.810 202.040 29.980 202.185 ;
        RECT 30.755 202.155 31.915 202.395 ;
        RECT 32.095 202.375 32.365 203.105 ;
        RECT 32.545 202.555 32.885 203.285 ;
        RECT 32.095 202.155 32.865 202.375 ;
        RECT 29.695 201.710 29.980 202.040 ;
        RECT 29.810 201.455 29.980 201.710 ;
        RECT 30.215 201.635 30.545 202.005 ;
        RECT 30.745 201.645 31.045 201.975 ;
        RECT 31.225 201.665 31.750 201.975 ;
        RECT 31.930 201.665 32.395 201.975 ;
        RECT 29.355 200.905 29.615 201.410 ;
        RECT 29.810 201.285 30.475 201.455 ;
        RECT 29.795 200.735 30.125 201.115 ;
        RECT 30.305 200.905 30.475 201.285 ;
        RECT 30.755 200.735 31.045 201.465 ;
        RECT 31.225 201.025 31.455 201.665 ;
        RECT 32.575 201.485 32.865 202.155 ;
        RECT 31.635 201.285 32.865 201.485 ;
        RECT 31.635 200.915 31.945 201.285 ;
        RECT 32.125 200.735 32.795 201.105 ;
        RECT 33.055 200.915 33.315 203.105 ;
        RECT 33.495 202.315 33.805 203.115 ;
        RECT 33.975 202.485 34.285 203.285 ;
        RECT 34.455 202.655 34.715 203.115 ;
        RECT 34.885 202.825 35.140 203.285 ;
        RECT 35.315 202.655 35.575 203.115 ;
        RECT 34.455 202.485 35.575 202.655 ;
        RECT 33.495 202.145 34.525 202.315 ;
        RECT 33.495 201.235 33.665 202.145 ;
        RECT 33.835 201.405 34.185 201.975 ;
        RECT 34.355 201.895 34.525 202.145 ;
        RECT 35.315 202.235 35.575 202.485 ;
        RECT 35.745 202.415 36.030 203.285 ;
        RECT 36.345 202.540 36.615 203.285 ;
        RECT 37.245 203.280 43.520 203.285 ;
        RECT 36.785 202.370 37.075 203.110 ;
        RECT 37.245 202.555 37.500 203.280 ;
        RECT 37.685 202.385 37.945 203.110 ;
        RECT 38.115 202.555 38.360 203.280 ;
        RECT 38.545 202.385 38.805 203.110 ;
        RECT 38.975 202.555 39.220 203.280 ;
        RECT 39.405 202.385 39.665 203.110 ;
        RECT 39.835 202.555 40.080 203.280 ;
        RECT 40.250 202.385 40.510 203.110 ;
        RECT 40.680 202.555 40.940 203.280 ;
        RECT 41.110 202.385 41.370 203.110 ;
        RECT 41.540 202.555 41.800 203.280 ;
        RECT 41.970 202.385 42.230 203.110 ;
        RECT 42.400 202.555 42.660 203.280 ;
        RECT 42.830 202.385 43.090 203.110 ;
        RECT 43.260 202.485 43.520 203.280 ;
        RECT 37.685 202.370 43.090 202.385 ;
        RECT 35.315 202.065 36.070 202.235 ;
        RECT 34.355 201.725 35.495 201.895 ;
        RECT 35.665 201.555 36.070 202.065 ;
        RECT 34.420 201.385 36.070 201.555 ;
        RECT 36.345 202.145 43.090 202.370 ;
        RECT 36.345 201.555 37.510 202.145 ;
        RECT 43.690 201.975 43.940 203.110 ;
        RECT 44.120 202.475 44.380 203.285 ;
        RECT 44.555 201.975 44.800 203.115 ;
        RECT 44.980 202.475 45.275 203.285 ;
        RECT 45.545 202.540 45.815 203.285 ;
        RECT 46.445 203.280 52.720 203.285 ;
        RECT 45.985 202.370 46.275 203.110 ;
        RECT 46.445 202.555 46.700 203.280 ;
        RECT 46.885 202.385 47.145 203.110 ;
        RECT 47.315 202.555 47.560 203.280 ;
        RECT 47.745 202.385 48.005 203.110 ;
        RECT 48.175 202.555 48.420 203.280 ;
        RECT 48.605 202.385 48.865 203.110 ;
        RECT 49.035 202.555 49.280 203.280 ;
        RECT 49.450 202.385 49.710 203.110 ;
        RECT 49.880 202.555 50.140 203.280 ;
        RECT 50.310 202.385 50.570 203.110 ;
        RECT 50.740 202.555 51.000 203.280 ;
        RECT 51.170 202.385 51.430 203.110 ;
        RECT 51.600 202.555 51.860 203.280 ;
        RECT 52.030 202.385 52.290 203.110 ;
        RECT 52.460 202.485 52.720 203.280 ;
        RECT 46.885 202.370 52.290 202.385 ;
        RECT 45.545 202.145 52.290 202.370 ;
        RECT 37.680 201.725 44.800 201.975 ;
        RECT 36.345 201.385 43.090 201.555 ;
        RECT 33.495 200.905 33.795 201.235 ;
        RECT 33.965 200.735 34.240 201.215 ;
        RECT 34.420 200.995 34.715 201.385 ;
        RECT 34.885 200.735 35.140 201.215 ;
        RECT 35.315 200.995 35.575 201.385 ;
        RECT 35.745 200.735 36.025 201.215 ;
        RECT 36.345 200.735 36.645 201.215 ;
        RECT 36.815 200.930 37.075 201.385 ;
        RECT 37.245 200.735 37.505 201.215 ;
        RECT 37.685 200.930 37.945 201.385 ;
        RECT 38.115 200.735 38.365 201.215 ;
        RECT 38.545 200.930 38.805 201.385 ;
        RECT 38.975 200.735 39.225 201.215 ;
        RECT 39.405 200.930 39.665 201.385 ;
        RECT 39.835 200.735 40.080 201.215 ;
        RECT 40.250 200.930 40.525 201.385 ;
        RECT 40.695 200.735 40.940 201.215 ;
        RECT 41.110 200.930 41.370 201.385 ;
        RECT 41.540 200.735 41.800 201.215 ;
        RECT 41.970 200.930 42.230 201.385 ;
        RECT 42.400 200.735 42.660 201.215 ;
        RECT 42.830 200.930 43.090 201.385 ;
        RECT 43.260 200.735 43.520 201.295 ;
        RECT 43.690 200.915 43.940 201.725 ;
        RECT 44.120 200.735 44.380 201.260 ;
        RECT 44.550 200.915 44.800 201.725 ;
        RECT 44.970 201.415 45.285 201.975 ;
        RECT 45.545 201.555 46.710 202.145 ;
        RECT 52.890 201.975 53.140 203.110 ;
        RECT 53.320 202.475 53.580 203.285 ;
        RECT 53.755 201.975 54.000 203.115 ;
        RECT 54.180 202.475 54.475 203.285 ;
        RECT 54.655 202.120 54.945 203.285 ;
        RECT 55.115 202.315 55.405 203.115 ;
        RECT 55.575 202.485 55.810 203.285 ;
        RECT 55.995 202.945 57.530 203.115 ;
        RECT 55.995 202.315 56.325 202.945 ;
        RECT 55.115 202.145 56.325 202.315 ;
        RECT 46.880 201.725 54.000 201.975 ;
        RECT 45.545 201.385 52.290 201.555 ;
        RECT 44.980 200.735 45.285 201.245 ;
        RECT 45.545 200.735 45.845 201.215 ;
        RECT 46.015 200.930 46.275 201.385 ;
        RECT 46.445 200.735 46.705 201.215 ;
        RECT 46.885 200.930 47.145 201.385 ;
        RECT 47.315 200.735 47.565 201.215 ;
        RECT 47.745 200.930 48.005 201.385 ;
        RECT 48.175 200.735 48.425 201.215 ;
        RECT 48.605 200.930 48.865 201.385 ;
        RECT 49.035 200.735 49.280 201.215 ;
        RECT 49.450 200.930 49.725 201.385 ;
        RECT 49.895 200.735 50.140 201.215 ;
        RECT 50.310 200.930 50.570 201.385 ;
        RECT 50.740 200.735 51.000 201.215 ;
        RECT 51.170 200.930 51.430 201.385 ;
        RECT 51.600 200.735 51.860 201.215 ;
        RECT 52.030 200.930 52.290 201.385 ;
        RECT 52.460 200.735 52.720 201.295 ;
        RECT 52.890 200.915 53.140 201.725 ;
        RECT 53.320 200.735 53.580 201.260 ;
        RECT 53.750 200.915 54.000 201.725 ;
        RECT 54.170 201.415 54.485 201.975 ;
        RECT 55.115 201.645 55.360 201.975 ;
        RECT 55.530 201.475 55.700 202.145 ;
        RECT 56.495 201.975 56.730 202.720 ;
        RECT 55.870 201.645 56.270 201.975 ;
        RECT 56.440 201.645 56.730 201.975 ;
        RECT 56.920 201.975 57.190 202.720 ;
        RECT 57.360 202.315 57.530 202.945 ;
        RECT 57.700 202.485 58.095 203.285 ;
        RECT 57.360 202.145 58.095 202.315 ;
        RECT 56.920 201.645 57.250 201.975 ;
        RECT 57.420 201.645 57.755 201.975 ;
        RECT 57.925 201.645 58.095 202.145 ;
        RECT 58.265 201.965 58.620 203.115 ;
        RECT 58.790 202.135 59.085 203.285 ;
        RECT 59.265 202.145 59.595 203.285 ;
        RECT 60.125 202.315 60.455 203.100 ;
        RECT 60.645 202.475 60.940 203.285 ;
        RECT 59.775 202.145 60.455 202.315 ;
        RECT 58.265 201.705 59.085 201.965 ;
        RECT 59.255 201.725 59.605 201.975 ;
        RECT 58.265 201.645 58.620 201.705 ;
        RECT 54.180 200.735 54.485 201.245 ;
        RECT 54.655 200.735 54.945 201.460 ;
        RECT 55.115 200.905 55.700 201.475 ;
        RECT 55.950 201.305 57.335 201.475 ;
        RECT 55.950 200.960 56.280 201.305 ;
        RECT 56.495 200.735 56.870 201.135 ;
        RECT 57.050 200.960 57.335 201.305 ;
        RECT 57.505 200.735 58.175 201.475 ;
        RECT 58.345 200.905 58.620 201.645 ;
        RECT 59.775 201.545 59.945 202.145 ;
        RECT 61.120 201.975 61.365 203.115 ;
        RECT 61.540 202.475 61.800 203.285 ;
        RECT 62.400 203.280 68.675 203.285 ;
        RECT 61.980 201.975 62.230 203.110 ;
        RECT 62.400 202.485 62.660 203.280 ;
        RECT 62.830 202.385 63.090 203.110 ;
        RECT 63.260 202.555 63.520 203.280 ;
        RECT 63.690 202.385 63.950 203.110 ;
        RECT 64.120 202.555 64.380 203.280 ;
        RECT 64.550 202.385 64.810 203.110 ;
        RECT 64.980 202.555 65.240 203.280 ;
        RECT 65.410 202.385 65.670 203.110 ;
        RECT 65.840 202.555 66.085 203.280 ;
        RECT 66.255 202.385 66.515 203.110 ;
        RECT 66.700 202.555 66.945 203.280 ;
        RECT 67.115 202.385 67.375 203.110 ;
        RECT 67.560 202.555 67.805 203.280 ;
        RECT 67.975 202.385 68.235 203.110 ;
        RECT 68.420 202.555 68.675 203.280 ;
        RECT 62.830 202.370 68.235 202.385 ;
        RECT 68.845 202.370 69.135 203.110 ;
        RECT 69.305 202.540 69.575 203.285 ;
        RECT 69.845 202.475 70.140 203.285 ;
        RECT 62.830 202.145 69.575 202.370 ;
        RECT 60.115 201.725 60.465 201.975 ;
        RECT 58.790 200.735 59.085 201.535 ;
        RECT 59.265 200.735 59.535 201.545 ;
        RECT 59.705 200.905 60.035 201.545 ;
        RECT 60.205 200.735 60.445 201.545 ;
        RECT 60.635 201.415 60.950 201.975 ;
        RECT 61.120 201.725 68.240 201.975 ;
        RECT 60.635 200.735 60.940 201.245 ;
        RECT 61.120 200.915 61.370 201.725 ;
        RECT 61.540 200.735 61.800 201.260 ;
        RECT 61.980 200.915 62.230 201.725 ;
        RECT 68.410 201.555 69.575 202.145 ;
        RECT 70.320 201.975 70.565 203.115 ;
        RECT 70.740 202.475 71.000 203.285 ;
        RECT 71.600 203.280 77.875 203.285 ;
        RECT 71.180 201.975 71.430 203.110 ;
        RECT 71.600 202.485 71.860 203.280 ;
        RECT 72.030 202.385 72.290 203.110 ;
        RECT 72.460 202.555 72.720 203.280 ;
        RECT 72.890 202.385 73.150 203.110 ;
        RECT 73.320 202.555 73.580 203.280 ;
        RECT 73.750 202.385 74.010 203.110 ;
        RECT 74.180 202.555 74.440 203.280 ;
        RECT 74.610 202.385 74.870 203.110 ;
        RECT 75.040 202.555 75.285 203.280 ;
        RECT 75.455 202.385 75.715 203.110 ;
        RECT 75.900 202.555 76.145 203.280 ;
        RECT 76.315 202.385 76.575 203.110 ;
        RECT 76.760 202.555 77.005 203.280 ;
        RECT 77.175 202.385 77.435 203.110 ;
        RECT 77.620 202.555 77.875 203.280 ;
        RECT 72.030 202.370 77.435 202.385 ;
        RECT 78.045 202.370 78.335 203.110 ;
        RECT 78.505 202.540 78.775 203.285 ;
        RECT 72.030 202.145 78.775 202.370 ;
        RECT 79.125 202.355 79.295 203.115 ;
        RECT 79.475 202.525 79.805 203.285 ;
        RECT 79.125 202.185 79.790 202.355 ;
        RECT 79.975 202.210 80.245 203.115 ;
        RECT 62.830 201.385 69.575 201.555 ;
        RECT 69.835 201.415 70.150 201.975 ;
        RECT 70.320 201.725 77.440 201.975 ;
        RECT 62.400 200.735 62.660 201.295 ;
        RECT 62.830 200.930 63.090 201.385 ;
        RECT 63.260 200.735 63.520 201.215 ;
        RECT 63.690 200.930 63.950 201.385 ;
        RECT 64.120 200.735 64.380 201.215 ;
        RECT 64.550 200.930 64.810 201.385 ;
        RECT 64.980 200.735 65.225 201.215 ;
        RECT 65.395 200.930 65.670 201.385 ;
        RECT 65.840 200.735 66.085 201.215 ;
        RECT 66.255 200.930 66.515 201.385 ;
        RECT 66.695 200.735 66.945 201.215 ;
        RECT 67.115 200.930 67.375 201.385 ;
        RECT 67.555 200.735 67.805 201.215 ;
        RECT 67.975 200.930 68.235 201.385 ;
        RECT 68.415 200.735 68.675 201.215 ;
        RECT 68.845 200.930 69.105 201.385 ;
        RECT 69.275 200.735 69.575 201.215 ;
        RECT 69.835 200.735 70.140 201.245 ;
        RECT 70.320 200.915 70.570 201.725 ;
        RECT 70.740 200.735 71.000 201.260 ;
        RECT 71.180 200.915 71.430 201.725 ;
        RECT 77.610 201.555 78.775 202.145 ;
        RECT 79.620 202.040 79.790 202.185 ;
        RECT 79.055 201.635 79.385 202.005 ;
        RECT 79.620 201.710 79.905 202.040 ;
        RECT 72.030 201.385 78.775 201.555 ;
        RECT 79.620 201.455 79.790 201.710 ;
        RECT 71.600 200.735 71.860 201.295 ;
        RECT 72.030 200.930 72.290 201.385 ;
        RECT 72.460 200.735 72.720 201.215 ;
        RECT 72.890 200.930 73.150 201.385 ;
        RECT 73.320 200.735 73.580 201.215 ;
        RECT 73.750 200.930 74.010 201.385 ;
        RECT 74.180 200.735 74.425 201.215 ;
        RECT 74.595 200.930 74.870 201.385 ;
        RECT 75.040 200.735 75.285 201.215 ;
        RECT 75.455 200.930 75.715 201.385 ;
        RECT 75.895 200.735 76.145 201.215 ;
        RECT 76.315 200.930 76.575 201.385 ;
        RECT 76.755 200.735 77.005 201.215 ;
        RECT 77.175 200.930 77.435 201.385 ;
        RECT 77.615 200.735 77.875 201.215 ;
        RECT 78.045 200.930 78.305 201.385 ;
        RECT 79.125 201.285 79.790 201.455 ;
        RECT 80.075 201.410 80.245 202.210 ;
        RECT 80.415 202.120 80.705 203.285 ;
        RECT 80.875 202.145 81.205 203.285 ;
        RECT 81.375 202.655 81.730 203.115 ;
        RECT 81.900 202.825 82.475 203.285 ;
        RECT 82.645 202.655 82.975 203.115 ;
        RECT 81.375 202.485 82.975 202.655 ;
        RECT 83.175 202.485 83.430 203.285 ;
        RECT 81.375 202.145 81.650 202.485 ;
        RECT 81.830 201.925 82.020 202.305 ;
        RECT 80.875 201.725 82.020 201.925 ;
        RECT 82.200 201.585 82.480 202.485 ;
        RECT 83.600 202.315 83.900 202.510 ;
        RECT 82.650 202.145 83.900 202.315 ;
        RECT 84.185 202.355 84.355 203.115 ;
        RECT 84.570 202.525 84.900 203.285 ;
        RECT 84.185 202.185 84.900 202.355 ;
        RECT 85.070 202.210 85.325 203.115 ;
        RECT 82.650 201.725 82.980 202.145 ;
        RECT 83.210 201.645 83.555 201.975 ;
        RECT 82.200 201.555 82.485 201.585 ;
        RECT 78.475 200.735 78.775 201.215 ;
        RECT 79.125 200.905 79.295 201.285 ;
        RECT 79.475 200.735 79.805 201.115 ;
        RECT 79.985 200.905 80.245 201.410 ;
        RECT 80.415 200.735 80.705 201.460 ;
        RECT 80.875 201.345 81.985 201.555 ;
        RECT 80.875 200.905 81.225 201.345 ;
        RECT 81.395 200.735 81.565 201.175 ;
        RECT 81.735 201.115 81.985 201.345 ;
        RECT 82.155 201.285 82.485 201.555 ;
        RECT 82.655 201.115 82.930 201.555 ;
        RECT 83.730 201.490 83.900 202.145 ;
        RECT 84.095 201.635 84.450 202.005 ;
        RECT 84.730 201.975 84.900 202.185 ;
        RECT 84.730 201.645 84.985 201.975 ;
        RECT 81.735 200.905 82.930 201.115 ;
        RECT 83.165 200.735 83.495 201.475 ;
        RECT 83.665 201.160 83.900 201.490 ;
        RECT 84.730 201.455 84.900 201.645 ;
        RECT 85.155 201.480 85.325 202.210 ;
        RECT 85.500 202.135 85.760 203.285 ;
        RECT 85.935 202.195 87.145 203.285 ;
        RECT 85.935 201.655 86.455 202.195 ;
        RECT 84.185 201.285 84.900 201.455 ;
        RECT 84.185 200.905 84.355 201.285 ;
        RECT 84.570 200.735 84.900 201.115 ;
        RECT 85.070 200.905 85.325 201.480 ;
        RECT 85.500 200.735 85.760 201.575 ;
        RECT 86.625 201.485 87.145 202.025 ;
        RECT 85.935 200.735 87.145 201.485 ;
        RECT 15.930 200.565 87.230 200.735 ;
        RECT 16.015 199.815 17.225 200.565 ;
        RECT 16.015 199.275 16.535 199.815 ;
        RECT 17.400 199.725 17.660 200.565 ;
        RECT 17.835 199.820 18.090 200.395 ;
        RECT 18.260 200.185 18.590 200.565 ;
        RECT 18.805 200.015 18.975 200.395 ;
        RECT 18.260 199.845 18.975 200.015 ;
        RECT 16.705 199.105 17.225 199.645 ;
        RECT 16.015 198.015 17.225 199.105 ;
        RECT 17.400 198.015 17.660 199.165 ;
        RECT 17.835 199.090 18.005 199.820 ;
        RECT 18.260 199.655 18.430 199.845 ;
        RECT 18.175 199.325 18.430 199.655 ;
        RECT 18.260 199.115 18.430 199.325 ;
        RECT 18.710 199.295 19.065 199.665 ;
        RECT 17.835 198.185 18.090 199.090 ;
        RECT 18.260 198.945 18.975 199.115 ;
        RECT 18.260 198.015 18.590 198.775 ;
        RECT 18.805 198.185 18.975 198.945 ;
        RECT 19.695 198.185 20.445 200.395 ;
        RECT 20.705 200.015 20.875 200.395 ;
        RECT 21.055 200.185 21.385 200.565 ;
        RECT 20.705 199.845 21.370 200.015 ;
        RECT 21.565 199.890 21.825 200.395 ;
        RECT 20.635 199.295 20.975 199.665 ;
        RECT 21.200 199.590 21.370 199.845 ;
        RECT 21.200 199.260 21.475 199.590 ;
        RECT 21.200 199.115 21.370 199.260 ;
        RECT 20.695 198.945 21.370 199.115 ;
        RECT 21.645 199.090 21.825 199.890 ;
        RECT 20.695 198.185 20.875 198.945 ;
        RECT 21.055 198.015 21.385 198.775 ;
        RECT 21.555 198.185 21.825 199.090 ;
        RECT 22.000 200.090 22.335 200.350 ;
        RECT 22.505 200.165 22.835 200.565 ;
        RECT 23.005 200.165 24.620 200.335 ;
        RECT 22.000 198.735 22.255 200.090 ;
        RECT 23.005 199.995 23.175 200.165 ;
        RECT 22.615 199.825 23.175 199.995 ;
        RECT 22.615 199.655 22.785 199.825 ;
        RECT 22.480 199.325 22.785 199.655 ;
        RECT 22.980 199.545 23.230 199.655 ;
        RECT 23.440 199.545 23.710 199.985 ;
        RECT 23.900 199.885 24.190 199.985 ;
        RECT 23.895 199.715 24.190 199.885 ;
        RECT 22.975 199.375 23.230 199.545 ;
        RECT 23.435 199.375 23.710 199.545 ;
        RECT 22.980 199.325 23.230 199.375 ;
        RECT 23.440 199.325 23.710 199.375 ;
        RECT 23.900 199.325 24.190 199.715 ;
        RECT 24.360 199.325 24.780 199.990 ;
        RECT 25.165 199.845 25.495 200.565 ;
        RECT 25.090 199.325 25.440 199.655 ;
        RECT 22.615 199.155 22.785 199.325 ;
        RECT 25.235 199.205 25.440 199.325 ;
        RECT 25.675 199.620 26.015 200.395 ;
        RECT 26.185 200.105 26.355 200.565 ;
        RECT 26.595 200.130 26.955 200.395 ;
        RECT 26.595 200.125 26.950 200.130 ;
        RECT 26.595 200.115 26.945 200.125 ;
        RECT 26.595 200.110 26.940 200.115 ;
        RECT 26.595 200.100 26.935 200.110 ;
        RECT 27.585 200.105 27.755 200.565 ;
        RECT 26.595 200.095 26.930 200.100 ;
        RECT 26.595 200.085 26.920 200.095 ;
        RECT 26.595 200.075 26.910 200.085 ;
        RECT 26.595 199.935 26.895 200.075 ;
        RECT 26.185 199.745 26.895 199.935 ;
        RECT 27.085 199.935 27.415 200.015 ;
        RECT 27.925 199.935 28.265 200.395 ;
        RECT 27.085 199.745 28.265 199.935 ;
        RECT 28.470 199.825 29.085 200.395 ;
        RECT 29.255 200.055 29.470 200.565 ;
        RECT 29.700 200.055 29.980 200.385 ;
        RECT 30.160 200.055 30.400 200.565 ;
        RECT 22.615 198.985 24.985 199.155 ;
        RECT 25.235 199.035 25.445 199.205 ;
        RECT 22.000 198.225 22.335 198.735 ;
        RECT 22.585 198.015 22.915 198.815 ;
        RECT 23.160 198.605 24.585 198.775 ;
        RECT 23.160 198.185 23.445 198.605 ;
        RECT 23.700 198.015 24.030 198.435 ;
        RECT 24.255 198.355 24.585 198.605 ;
        RECT 24.815 198.525 24.985 198.985 ;
        RECT 25.245 198.355 25.415 198.855 ;
        RECT 24.255 198.185 25.415 198.355 ;
        RECT 25.675 198.185 25.955 199.620 ;
        RECT 26.185 199.175 26.470 199.745 ;
        RECT 26.655 199.345 27.125 199.575 ;
        RECT 27.295 199.555 27.625 199.575 ;
        RECT 27.295 199.375 27.745 199.555 ;
        RECT 27.935 199.375 28.265 199.575 ;
        RECT 26.185 198.960 27.335 199.175 ;
        RECT 26.125 198.015 26.835 198.790 ;
        RECT 27.005 198.185 27.335 198.960 ;
        RECT 27.530 198.260 27.745 199.375 ;
        RECT 28.035 199.035 28.265 199.375 ;
        RECT 28.470 198.805 28.785 199.825 ;
        RECT 28.955 199.155 29.125 199.655 ;
        RECT 29.375 199.325 29.640 199.885 ;
        RECT 29.810 199.155 29.980 200.055 ;
        RECT 30.150 199.325 30.505 199.885 ;
        RECT 30.740 199.800 31.195 200.565 ;
        RECT 31.470 200.185 32.770 200.395 ;
        RECT 33.025 200.205 33.355 200.565 ;
        RECT 32.600 200.035 32.770 200.185 ;
        RECT 33.525 200.065 33.785 200.395 ;
        RECT 31.670 199.575 31.890 199.975 ;
        RECT 30.735 199.375 31.225 199.575 ;
        RECT 31.415 199.365 31.890 199.575 ;
        RECT 32.135 199.575 32.345 199.975 ;
        RECT 32.600 199.910 33.355 200.035 ;
        RECT 32.600 199.865 33.445 199.910 ;
        RECT 33.175 199.745 33.445 199.865 ;
        RECT 32.135 199.365 32.465 199.575 ;
        RECT 32.635 199.305 33.045 199.610 ;
        RECT 28.955 198.985 30.380 199.155 ;
        RECT 27.925 198.015 28.255 198.735 ;
        RECT 28.470 198.185 29.005 198.805 ;
        RECT 29.175 198.015 29.505 198.815 ;
        RECT 29.990 198.810 30.380 198.985 ;
        RECT 30.740 199.135 31.915 199.195 ;
        RECT 33.275 199.170 33.445 199.745 ;
        RECT 33.245 199.135 33.445 199.170 ;
        RECT 30.740 199.025 33.445 199.135 ;
        RECT 30.740 198.405 30.995 199.025 ;
        RECT 31.585 198.965 33.385 199.025 ;
        RECT 31.585 198.935 31.915 198.965 ;
        RECT 33.615 198.865 33.785 200.065 ;
        RECT 31.245 198.765 31.430 198.855 ;
        RECT 32.020 198.765 32.855 198.775 ;
        RECT 31.245 198.565 32.855 198.765 ;
        RECT 31.245 198.525 31.475 198.565 ;
        RECT 30.740 198.185 31.075 198.405 ;
        RECT 32.080 198.015 32.435 198.395 ;
        RECT 32.605 198.185 32.855 198.565 ;
        RECT 33.105 198.015 33.355 198.795 ;
        RECT 33.525 198.185 33.785 198.865 ;
        RECT 33.955 200.065 34.215 200.395 ;
        RECT 34.385 200.205 34.715 200.565 ;
        RECT 34.970 200.185 36.270 200.395 ;
        RECT 33.955 198.865 34.125 200.065 ;
        RECT 34.970 200.035 35.140 200.185 ;
        RECT 34.385 199.910 35.140 200.035 ;
        RECT 34.295 199.865 35.140 199.910 ;
        RECT 34.295 199.745 34.565 199.865 ;
        RECT 34.295 199.170 34.465 199.745 ;
        RECT 34.695 199.305 35.105 199.610 ;
        RECT 35.395 199.575 35.605 199.975 ;
        RECT 35.275 199.365 35.605 199.575 ;
        RECT 35.850 199.575 36.070 199.975 ;
        RECT 36.545 199.800 37.000 200.565 ;
        RECT 37.175 199.765 37.870 200.395 ;
        RECT 38.075 199.765 38.385 200.565 ;
        RECT 38.565 199.840 38.895 200.350 ;
        RECT 39.065 200.165 39.395 200.565 ;
        RECT 40.445 199.995 40.775 200.335 ;
        RECT 40.945 200.165 41.275 200.565 ;
        RECT 35.850 199.365 36.325 199.575 ;
        RECT 36.515 199.375 37.005 199.575 ;
        RECT 37.195 199.325 37.530 199.575 ;
        RECT 34.295 199.135 34.495 199.170 ;
        RECT 35.825 199.135 37.000 199.195 ;
        RECT 37.700 199.165 37.870 199.765 ;
        RECT 38.040 199.325 38.375 199.595 ;
        RECT 34.295 199.025 37.000 199.135 ;
        RECT 34.355 198.965 36.155 199.025 ;
        RECT 35.825 198.935 36.155 198.965 ;
        RECT 33.955 198.185 34.215 198.865 ;
        RECT 34.385 198.015 34.635 198.795 ;
        RECT 34.885 198.765 35.720 198.775 ;
        RECT 36.310 198.765 36.495 198.855 ;
        RECT 34.885 198.565 36.495 198.765 ;
        RECT 34.885 198.185 35.135 198.565 ;
        RECT 36.265 198.525 36.495 198.565 ;
        RECT 36.745 198.405 37.000 199.025 ;
        RECT 35.305 198.015 35.660 198.395 ;
        RECT 36.665 198.185 37.000 198.405 ;
        RECT 37.175 198.015 37.435 199.155 ;
        RECT 37.605 198.185 37.935 199.165 ;
        RECT 38.105 198.015 38.385 199.155 ;
        RECT 38.565 199.075 38.755 199.840 ;
        RECT 39.065 199.825 41.430 199.995 ;
        RECT 41.775 199.840 42.065 200.565 ;
        RECT 39.065 199.655 39.235 199.825 ;
        RECT 38.925 199.325 39.235 199.655 ;
        RECT 39.405 199.325 39.710 199.655 ;
        RECT 38.565 198.225 38.895 199.075 ;
        RECT 39.065 198.015 39.315 199.155 ;
        RECT 39.495 198.995 39.710 199.325 ;
        RECT 39.885 198.995 40.170 199.655 ;
        RECT 40.365 198.995 40.630 199.655 ;
        RECT 40.845 198.995 41.090 199.655 ;
        RECT 41.260 198.825 41.430 199.825 ;
        RECT 42.235 199.825 42.555 200.200 ;
        RECT 42.810 199.825 42.980 200.565 ;
        RECT 43.230 199.995 43.400 200.200 ;
        RECT 43.645 200.165 44.000 200.565 ;
        RECT 44.175 199.995 44.345 200.345 ;
        RECT 44.545 200.165 44.875 200.565 ;
        RECT 45.045 199.995 45.215 200.345 ;
        RECT 45.385 200.165 45.765 200.565 ;
        RECT 43.230 199.825 43.750 199.995 ;
        RECT 44.175 199.825 45.785 199.995 ;
        RECT 45.955 199.890 46.230 200.235 ;
        RECT 39.505 198.655 40.795 198.825 ;
        RECT 39.505 198.235 39.755 198.655 ;
        RECT 39.985 198.015 40.315 198.485 ;
        RECT 40.545 198.235 40.795 198.655 ;
        RECT 40.975 198.655 41.430 198.825 ;
        RECT 40.975 198.225 41.305 198.655 ;
        RECT 41.775 198.015 42.065 199.180 ;
        RECT 42.235 198.785 42.410 199.825 ;
        RECT 42.580 198.955 42.930 199.655 ;
        RECT 43.100 199.325 43.390 199.655 ;
        RECT 43.560 199.575 43.750 199.825 ;
        RECT 45.615 199.655 45.785 199.825 ;
        RECT 43.560 199.405 44.005 199.575 ;
        RECT 43.560 199.125 43.750 199.405 ;
        RECT 44.400 199.235 44.570 199.655 ;
        RECT 44.790 199.325 45.445 199.655 ;
        RECT 45.615 199.325 45.890 199.655 ;
        RECT 43.145 198.955 43.750 199.125 ;
        RECT 43.920 199.065 44.570 199.235 ;
        RECT 45.615 199.155 45.785 199.325 ;
        RECT 46.060 199.155 46.230 199.890 ;
        RECT 46.400 199.625 46.570 200.565 ;
        RECT 46.845 200.225 47.180 200.395 ;
        RECT 46.845 199.825 47.460 200.225 ;
        RECT 48.140 200.185 48.475 200.565 ;
        RECT 49.065 200.125 49.300 200.565 ;
        RECT 49.470 200.035 49.800 200.395 ;
        RECT 49.970 200.205 50.300 200.565 ;
        RECT 50.515 200.055 50.820 200.565 ;
        RECT 47.630 199.825 48.900 200.015 ;
        RECT 49.470 199.865 50.290 200.035 ;
        RECT 46.835 199.325 47.110 199.655 ;
        RECT 43.920 198.785 44.090 199.065 ;
        RECT 45.125 198.985 45.785 199.155 ;
        RECT 45.125 198.865 45.295 198.985 ;
        RECT 42.235 198.615 44.090 198.785 ;
        RECT 44.260 198.695 45.295 198.865 ;
        RECT 42.235 198.195 42.495 198.615 ;
        RECT 44.260 198.445 44.430 198.695 ;
        RECT 42.665 198.015 42.995 198.445 ;
        RECT 43.685 198.275 44.430 198.445 ;
        RECT 44.655 198.195 45.295 198.525 ;
        RECT 45.465 198.015 45.745 198.815 ;
        RECT 45.955 198.185 46.230 199.155 ;
        RECT 46.400 198.015 46.570 199.210 ;
        RECT 47.280 199.140 47.460 199.825 ;
        RECT 47.630 199.325 47.990 199.655 ;
        RECT 48.280 199.545 48.570 199.655 ;
        RECT 48.275 199.375 48.570 199.545 ;
        RECT 48.280 199.325 48.570 199.375 ;
        RECT 48.740 199.325 49.075 199.655 ;
        RECT 49.245 199.325 49.925 199.655 ;
        RECT 49.245 199.140 49.415 199.325 ;
        RECT 46.840 198.885 49.415 199.140 ;
        RECT 46.840 198.185 47.105 198.885 ;
        RECT 47.275 198.015 47.605 198.715 ;
        RECT 47.775 198.185 48.445 198.885 ;
        RECT 50.095 198.745 50.290 199.865 ;
        RECT 50.515 199.325 50.830 199.885 ;
        RECT 51.000 199.575 51.250 200.385 ;
        RECT 51.420 200.040 51.680 200.565 ;
        RECT 51.860 199.575 52.110 200.385 ;
        RECT 52.280 200.005 52.540 200.565 ;
        RECT 52.710 199.915 52.970 200.370 ;
        RECT 53.140 200.085 53.400 200.565 ;
        RECT 53.570 199.915 53.830 200.370 ;
        RECT 54.000 200.085 54.260 200.565 ;
        RECT 54.430 199.915 54.690 200.370 ;
        RECT 54.860 200.085 55.105 200.565 ;
        RECT 55.275 199.915 55.550 200.370 ;
        RECT 55.720 200.085 55.965 200.565 ;
        RECT 56.135 199.915 56.395 200.370 ;
        RECT 56.575 200.085 56.825 200.565 ;
        RECT 56.995 199.915 57.255 200.370 ;
        RECT 57.435 200.085 57.685 200.565 ;
        RECT 57.855 199.915 58.115 200.370 ;
        RECT 58.295 200.085 58.555 200.565 ;
        RECT 58.725 199.915 58.985 200.370 ;
        RECT 59.155 200.085 59.455 200.565 ;
        RECT 59.715 200.225 61.075 200.395 ;
        RECT 52.710 199.745 59.455 199.915 ;
        RECT 59.715 199.745 60.075 200.225 ;
        RECT 60.245 199.825 60.575 200.055 ;
        RECT 60.745 199.995 61.075 200.225 ;
        RECT 61.245 200.165 61.575 200.565 ;
        RECT 61.745 199.995 62.075 200.395 ;
        RECT 60.745 199.825 62.075 199.995 ;
        RECT 62.345 199.825 62.675 200.565 ;
        RECT 51.000 199.325 58.120 199.575 ;
        RECT 48.950 198.015 49.380 198.715 ;
        RECT 49.560 198.575 50.290 198.745 ;
        RECT 49.560 198.185 49.750 198.575 ;
        RECT 49.920 198.015 50.250 198.395 ;
        RECT 50.525 198.015 50.820 198.825 ;
        RECT 51.000 198.185 51.245 199.325 ;
        RECT 51.420 198.015 51.680 198.825 ;
        RECT 51.860 198.190 52.110 199.325 ;
        RECT 58.290 199.155 59.455 199.745 ;
        RECT 59.715 199.405 60.075 199.575 ;
        RECT 59.715 199.325 60.045 199.405 ;
        RECT 52.710 198.930 59.455 199.155 ;
        RECT 52.710 198.915 58.115 198.930 ;
        RECT 52.280 198.020 52.540 198.815 ;
        RECT 52.710 198.190 52.970 198.915 ;
        RECT 53.140 198.020 53.400 198.745 ;
        RECT 53.570 198.190 53.830 198.915 ;
        RECT 54.000 198.020 54.260 198.745 ;
        RECT 54.430 198.190 54.690 198.915 ;
        RECT 54.860 198.020 55.120 198.745 ;
        RECT 55.290 198.190 55.550 198.915 ;
        RECT 55.720 198.020 55.965 198.745 ;
        RECT 56.135 198.190 56.395 198.915 ;
        RECT 56.580 198.020 56.825 198.745 ;
        RECT 56.995 198.190 57.255 198.915 ;
        RECT 57.440 198.020 57.685 198.745 ;
        RECT 57.855 198.190 58.115 198.915 ;
        RECT 58.300 198.020 58.555 198.745 ;
        RECT 58.725 198.190 59.015 198.930 ;
        RECT 52.280 198.015 58.555 198.020 ;
        RECT 59.185 198.015 59.455 198.760 ;
        RECT 59.715 198.015 60.075 199.155 ;
        RECT 60.245 198.865 60.445 199.825 ;
        RECT 60.615 199.545 60.860 199.655 ;
        RECT 60.615 199.375 60.865 199.545 ;
        RECT 60.615 199.035 60.860 199.375 ;
        RECT 61.135 199.035 61.355 199.655 ;
        RECT 61.610 199.035 61.785 199.655 ;
        RECT 62.055 199.035 62.275 199.655 ;
        RECT 62.445 198.865 62.755 199.655 ;
        RECT 60.245 198.695 62.755 198.865 ;
        RECT 60.745 198.185 61.075 198.695 ;
        RECT 62.245 198.015 62.755 198.525 ;
        RECT 62.925 198.185 63.255 200.395 ;
        RECT 63.425 199.765 63.685 200.565 ;
        RECT 64.035 200.185 64.365 200.565 ;
        RECT 64.535 200.015 64.725 200.395 ;
        RECT 64.895 200.205 65.225 200.565 ;
        RECT 64.325 199.825 64.725 200.015 ;
        RECT 65.445 199.995 65.635 200.395 ;
        RECT 64.895 199.825 65.635 199.995 ;
        RECT 63.425 198.015 63.685 199.155 ;
        RECT 63.865 198.015 64.155 198.985 ;
        RECT 64.325 198.185 64.555 199.825 ;
        RECT 64.895 199.655 65.065 199.825 ;
        RECT 64.725 198.960 65.065 199.655 ;
        RECT 65.235 199.240 65.560 199.655 ;
        RECT 66.010 199.325 66.390 200.285 ;
        RECT 66.575 200.085 66.905 200.565 ;
        RECT 66.580 199.325 66.895 199.900 ;
        RECT 67.535 199.840 67.825 200.565 ;
        RECT 67.995 200.055 68.300 200.565 ;
        RECT 67.995 199.325 68.310 199.885 ;
        RECT 68.480 199.575 68.730 200.385 ;
        RECT 68.900 200.040 69.160 200.565 ;
        RECT 69.340 199.575 69.590 200.385 ;
        RECT 69.760 200.005 70.020 200.565 ;
        RECT 70.190 199.915 70.450 200.370 ;
        RECT 70.620 200.085 70.880 200.565 ;
        RECT 71.050 199.915 71.310 200.370 ;
        RECT 71.480 200.085 71.740 200.565 ;
        RECT 71.910 199.915 72.170 200.370 ;
        RECT 72.340 200.085 72.585 200.565 ;
        RECT 72.755 199.915 73.030 200.370 ;
        RECT 73.200 200.085 73.445 200.565 ;
        RECT 73.615 199.915 73.875 200.370 ;
        RECT 74.055 200.085 74.305 200.565 ;
        RECT 74.475 199.915 74.735 200.370 ;
        RECT 74.915 200.085 75.165 200.565 ;
        RECT 75.335 199.915 75.595 200.370 ;
        RECT 75.775 200.085 76.035 200.565 ;
        RECT 76.205 199.915 76.465 200.370 ;
        RECT 76.635 200.085 76.935 200.565 ;
        RECT 70.190 199.745 76.935 199.915 ;
        RECT 77.195 199.745 77.490 200.565 ;
        RECT 77.660 199.825 78.100 200.385 ;
        RECT 78.270 199.825 78.720 200.565 ;
        RECT 78.890 199.995 79.060 200.395 ;
        RECT 79.230 200.165 79.650 200.565 ;
        RECT 79.820 199.995 80.050 200.395 ;
        RECT 78.890 199.825 80.050 199.995 ;
        RECT 80.220 199.825 80.705 200.395 ;
        RECT 68.480 199.325 75.600 199.575 ;
        RECT 64.725 198.730 65.560 198.960 ;
        RECT 64.725 198.015 65.055 198.430 ;
        RECT 65.245 198.185 65.560 198.730 ;
        RECT 65.730 198.715 66.845 198.980 ;
        RECT 65.730 198.185 65.955 198.715 ;
        RECT 66.125 198.015 66.455 198.525 ;
        RECT 66.625 198.185 66.845 198.715 ;
        RECT 67.535 198.015 67.825 199.180 ;
        RECT 68.005 198.015 68.300 198.825 ;
        RECT 68.480 198.185 68.725 199.325 ;
        RECT 68.900 198.015 69.160 198.825 ;
        RECT 69.340 198.190 69.590 199.325 ;
        RECT 75.770 199.155 76.935 199.745 ;
        RECT 77.660 199.575 77.970 199.825 ;
        RECT 77.195 199.355 77.970 199.575 ;
        RECT 70.190 198.930 76.935 199.155 ;
        RECT 70.190 198.915 75.595 198.930 ;
        RECT 69.760 198.020 70.020 198.815 ;
        RECT 70.190 198.190 70.450 198.915 ;
        RECT 70.620 198.020 70.880 198.745 ;
        RECT 71.050 198.190 71.310 198.915 ;
        RECT 71.480 198.020 71.740 198.745 ;
        RECT 71.910 198.190 72.170 198.915 ;
        RECT 72.340 198.020 72.600 198.745 ;
        RECT 72.770 198.190 73.030 198.915 ;
        RECT 73.200 198.020 73.445 198.745 ;
        RECT 73.615 198.190 73.875 198.915 ;
        RECT 74.060 198.020 74.305 198.745 ;
        RECT 74.475 198.190 74.735 198.915 ;
        RECT 74.920 198.020 75.165 198.745 ;
        RECT 75.335 198.190 75.595 198.915 ;
        RECT 75.780 198.020 76.035 198.745 ;
        RECT 76.205 198.190 76.495 198.930 ;
        RECT 69.760 198.015 76.035 198.020 ;
        RECT 76.665 198.015 76.935 198.760 ;
        RECT 77.195 198.015 77.490 199.185 ;
        RECT 77.660 198.815 77.970 199.355 ;
        RECT 78.140 199.205 78.310 199.655 ;
        RECT 78.480 199.375 78.870 199.655 ;
        RECT 79.055 199.325 79.300 199.655 ;
        RECT 78.140 199.035 78.930 199.205 ;
        RECT 77.660 198.185 78.100 198.815 ;
        RECT 78.275 198.015 78.590 198.865 ;
        RECT 78.760 198.355 78.930 199.035 ;
        RECT 79.100 198.525 79.300 199.325 ;
        RECT 79.500 198.525 79.750 199.655 ;
        RECT 79.965 199.325 80.365 199.655 ;
        RECT 80.535 199.155 80.705 199.825 ;
        RECT 80.875 199.745 81.170 200.565 ;
        RECT 81.340 199.825 81.780 200.385 ;
        RECT 81.950 199.825 82.400 200.565 ;
        RECT 82.570 199.995 82.740 200.395 ;
        RECT 82.910 200.165 83.330 200.565 ;
        RECT 83.500 199.995 83.730 200.395 ;
        RECT 82.570 199.825 83.730 199.995 ;
        RECT 83.900 199.825 84.385 200.395 ;
        RECT 81.340 199.575 81.650 199.825 ;
        RECT 80.875 199.355 81.650 199.575 ;
        RECT 79.940 198.985 80.705 199.155 ;
        RECT 79.940 198.355 80.190 198.985 ;
        RECT 78.760 198.185 80.190 198.355 ;
        RECT 80.365 198.015 80.700 198.815 ;
        RECT 80.875 198.015 81.170 199.185 ;
        RECT 81.340 198.815 81.650 199.355 ;
        RECT 81.820 199.205 81.990 199.655 ;
        RECT 82.160 199.375 82.550 199.655 ;
        RECT 82.735 199.325 82.980 199.655 ;
        RECT 81.820 199.035 82.610 199.205 ;
        RECT 81.340 198.185 81.780 198.815 ;
        RECT 81.955 198.015 82.270 198.865 ;
        RECT 82.440 198.355 82.610 199.035 ;
        RECT 82.780 198.525 82.980 199.325 ;
        RECT 83.180 198.525 83.430 199.655 ;
        RECT 83.645 199.325 84.045 199.655 ;
        RECT 84.215 199.155 84.385 199.825 ;
        RECT 83.620 198.985 84.385 199.155 ;
        RECT 84.555 199.890 84.815 200.395 ;
        RECT 84.995 200.185 85.325 200.565 ;
        RECT 85.505 200.015 85.675 200.395 ;
        RECT 84.555 199.090 84.735 199.890 ;
        RECT 85.010 199.845 85.675 200.015 ;
        RECT 85.010 199.590 85.180 199.845 ;
        RECT 85.935 199.815 87.145 200.565 ;
        RECT 84.905 199.260 85.180 199.590 ;
        RECT 85.405 199.295 85.745 199.665 ;
        RECT 85.010 199.115 85.180 199.260 ;
        RECT 83.620 198.355 83.870 198.985 ;
        RECT 82.440 198.185 83.870 198.355 ;
        RECT 84.045 198.015 84.380 198.815 ;
        RECT 84.555 198.185 84.825 199.090 ;
        RECT 85.010 198.945 85.685 199.115 ;
        RECT 84.995 198.015 85.325 198.775 ;
        RECT 85.505 198.185 85.685 198.945 ;
        RECT 85.935 199.105 86.455 199.645 ;
        RECT 86.625 199.275 87.145 199.815 ;
        RECT 85.935 198.015 87.145 199.105 ;
        RECT 15.930 197.845 87.230 198.015 ;
        RECT 16.015 196.755 17.225 197.845 ;
        RECT 16.015 196.045 16.535 196.585 ;
        RECT 16.705 196.215 17.225 196.755 ;
        RECT 17.855 196.705 18.145 197.845 ;
        RECT 18.315 197.125 18.765 197.675 ;
        RECT 18.955 197.125 19.285 197.845 ;
        RECT 16.015 195.295 17.225 196.045 ;
        RECT 17.855 195.295 18.145 196.095 ;
        RECT 18.315 195.755 18.565 197.125 ;
        RECT 19.495 196.955 19.795 197.505 ;
        RECT 19.965 197.175 20.245 197.845 ;
        RECT 18.855 196.785 19.795 196.955 ;
        RECT 18.855 196.535 19.025 196.785 ;
        RECT 20.130 196.535 20.445 196.975 ;
        RECT 20.800 196.875 21.190 197.050 ;
        RECT 21.675 197.045 22.005 197.845 ;
        RECT 22.175 197.055 22.710 197.675 ;
        RECT 20.800 196.705 22.225 196.875 ;
        RECT 18.735 196.205 19.025 196.535 ;
        RECT 19.195 196.285 19.525 196.535 ;
        RECT 19.755 196.285 20.445 196.535 ;
        RECT 18.855 196.115 19.025 196.205 ;
        RECT 18.855 195.925 20.245 196.115 ;
        RECT 20.675 195.975 21.030 196.535 ;
        RECT 18.315 195.465 18.865 195.755 ;
        RECT 19.035 195.295 19.285 195.755 ;
        RECT 19.915 195.565 20.245 195.925 ;
        RECT 21.200 195.805 21.370 196.705 ;
        RECT 21.540 195.975 21.805 196.535 ;
        RECT 22.055 196.205 22.225 196.705 ;
        RECT 22.395 196.035 22.710 197.055 ;
        RECT 23.005 197.505 24.165 197.675 ;
        RECT 23.005 197.005 23.175 197.505 ;
        RECT 23.435 196.875 23.605 197.335 ;
        RECT 23.835 197.255 24.165 197.505 ;
        RECT 24.390 197.425 24.720 197.845 ;
        RECT 24.975 197.255 25.260 197.675 ;
        RECT 23.835 197.085 25.260 197.255 ;
        RECT 25.505 197.045 25.835 197.845 ;
        RECT 26.085 197.125 26.420 197.635 ;
        RECT 22.980 196.535 23.185 196.825 ;
        RECT 23.435 196.705 25.805 196.875 ;
        RECT 25.635 196.535 25.805 196.705 ;
        RECT 22.980 196.485 23.330 196.535 ;
        RECT 22.975 196.315 23.330 196.485 ;
        RECT 22.980 196.205 23.330 196.315 ;
        RECT 20.780 195.295 21.020 195.805 ;
        RECT 21.200 195.475 21.480 195.805 ;
        RECT 21.710 195.295 21.925 195.805 ;
        RECT 22.095 195.465 22.710 196.035 ;
        RECT 22.925 195.295 23.255 196.015 ;
        RECT 23.640 195.870 24.060 196.535 ;
        RECT 24.230 195.875 24.520 196.535 ;
        RECT 24.710 196.485 24.980 196.535 ;
        RECT 25.190 196.485 25.440 196.535 ;
        RECT 24.710 196.315 24.985 196.485 ;
        RECT 25.190 196.315 25.445 196.485 ;
        RECT 24.710 195.875 24.980 196.315 ;
        RECT 25.190 196.205 25.440 196.315 ;
        RECT 25.635 196.205 25.940 196.535 ;
        RECT 25.635 196.035 25.805 196.205 ;
        RECT 25.245 195.865 25.805 196.035 ;
        RECT 25.245 195.695 25.415 195.865 ;
        RECT 26.165 195.770 26.420 197.125 ;
        RECT 23.800 195.525 25.415 195.695 ;
        RECT 25.585 195.295 25.915 195.695 ;
        RECT 26.085 195.510 26.420 195.770 ;
        RECT 27.515 196.770 27.785 197.675 ;
        RECT 27.955 197.085 28.285 197.845 ;
        RECT 28.465 196.915 28.635 197.675 ;
        RECT 27.515 195.970 27.685 196.770 ;
        RECT 27.970 196.745 28.635 196.915 ;
        RECT 27.970 196.600 28.140 196.745 ;
        RECT 28.895 196.680 29.185 197.845 ;
        RECT 29.355 196.705 29.615 197.845 ;
        RECT 29.785 196.695 30.115 197.675 ;
        RECT 30.285 196.705 30.565 197.845 ;
        RECT 30.740 196.705 31.060 197.845 ;
        RECT 27.855 196.270 28.140 196.600 ;
        RECT 27.970 196.015 28.140 196.270 ;
        RECT 28.375 196.195 28.705 196.565 ;
        RECT 29.375 196.285 29.710 196.535 ;
        RECT 29.880 196.095 30.050 196.695 ;
        RECT 31.240 196.535 31.435 197.585 ;
        RECT 31.615 196.995 31.945 197.675 ;
        RECT 32.145 197.045 32.400 197.845 ;
        RECT 31.615 196.715 31.965 196.995 ;
        RECT 30.220 196.265 30.555 196.535 ;
        RECT 30.800 196.485 31.060 196.535 ;
        RECT 30.795 196.315 31.060 196.485 ;
        RECT 30.800 196.205 31.060 196.315 ;
        RECT 31.240 196.205 31.625 196.535 ;
        RECT 31.795 196.335 31.965 196.715 ;
        RECT 32.155 196.505 32.400 196.865 ;
        RECT 32.730 196.835 33.030 197.675 ;
        RECT 33.225 197.005 33.475 197.845 ;
        RECT 34.065 197.255 34.870 197.675 ;
        RECT 33.645 197.085 35.210 197.255 ;
        RECT 33.645 196.835 33.815 197.085 ;
        RECT 32.730 196.665 33.815 196.835 ;
        RECT 31.795 196.165 32.315 196.335 ;
        RECT 32.575 196.205 32.905 196.495 ;
        RECT 27.515 195.465 27.775 195.970 ;
        RECT 27.970 195.845 28.635 196.015 ;
        RECT 27.955 195.295 28.285 195.675 ;
        RECT 28.465 195.465 28.635 195.845 ;
        RECT 28.895 195.295 29.185 196.020 ;
        RECT 29.355 195.465 30.050 196.095 ;
        RECT 30.255 195.295 30.565 196.095 ;
        RECT 30.740 195.825 31.955 195.995 ;
        RECT 30.740 195.475 31.030 195.825 ;
        RECT 31.225 195.295 31.555 195.655 ;
        RECT 31.725 195.520 31.955 195.825 ;
        RECT 32.145 195.600 32.315 196.165 ;
        RECT 33.075 196.035 33.245 196.665 ;
        RECT 33.985 196.535 34.305 196.915 ;
        RECT 33.415 196.285 33.745 196.495 ;
        RECT 33.925 196.285 34.305 196.535 ;
        RECT 34.495 196.495 34.870 196.915 ;
        RECT 35.040 196.835 35.210 197.085 ;
        RECT 35.380 197.005 35.710 197.845 ;
        RECT 35.880 197.085 36.545 197.675 ;
        RECT 35.040 196.665 35.960 196.835 ;
        RECT 35.790 196.495 35.960 196.665 ;
        RECT 34.495 196.485 34.980 196.495 ;
        RECT 34.475 196.315 34.980 196.485 ;
        RECT 34.495 196.285 34.980 196.315 ;
        RECT 35.170 196.285 35.620 196.495 ;
        RECT 35.790 196.285 36.125 196.495 ;
        RECT 36.295 196.115 36.545 197.085 ;
        RECT 37.180 197.455 37.515 197.675 ;
        RECT 38.520 197.465 38.875 197.845 ;
        RECT 37.180 196.835 37.435 197.455 ;
        RECT 37.685 197.295 37.915 197.335 ;
        RECT 39.045 197.295 39.295 197.675 ;
        RECT 37.685 197.095 39.295 197.295 ;
        RECT 37.685 197.005 37.870 197.095 ;
        RECT 38.460 197.085 39.295 197.095 ;
        RECT 39.545 197.065 39.795 197.845 ;
        RECT 39.965 196.995 40.225 197.675 ;
        RECT 40.485 197.100 40.755 197.845 ;
        RECT 41.385 197.840 47.660 197.845 ;
        RECT 38.025 196.895 38.355 196.925 ;
        RECT 38.025 196.835 39.825 196.895 ;
        RECT 37.180 196.725 39.885 196.835 ;
        RECT 37.180 196.665 38.355 196.725 ;
        RECT 39.685 196.690 39.885 196.725 ;
        RECT 37.175 196.285 37.665 196.485 ;
        RECT 37.855 196.285 38.330 196.495 ;
        RECT 32.735 195.855 33.245 196.035 ;
        RECT 33.650 195.945 35.350 196.115 ;
        RECT 33.650 195.855 34.035 195.945 ;
        RECT 32.735 195.465 33.065 195.855 ;
        RECT 33.235 195.515 34.420 195.685 ;
        RECT 34.680 195.295 34.850 195.765 ;
        RECT 35.020 195.480 35.350 195.945 ;
        RECT 35.520 195.295 35.690 196.115 ;
        RECT 35.860 195.475 36.545 196.115 ;
        RECT 37.180 195.295 37.635 196.060 ;
        RECT 38.110 195.885 38.330 196.285 ;
        RECT 38.575 196.285 38.905 196.495 ;
        RECT 38.575 195.885 38.785 196.285 ;
        RECT 39.075 196.250 39.485 196.555 ;
        RECT 39.715 196.115 39.885 196.690 ;
        RECT 39.615 195.995 39.885 196.115 ;
        RECT 39.040 195.950 39.885 195.995 ;
        RECT 39.040 195.825 39.795 195.950 ;
        RECT 39.040 195.675 39.210 195.825 ;
        RECT 40.055 195.795 40.225 196.995 ;
        RECT 40.925 196.930 41.215 197.670 ;
        RECT 41.385 197.115 41.640 197.840 ;
        RECT 41.825 196.945 42.085 197.670 ;
        RECT 42.255 197.115 42.500 197.840 ;
        RECT 42.685 196.945 42.945 197.670 ;
        RECT 43.115 197.115 43.360 197.840 ;
        RECT 43.545 196.945 43.805 197.670 ;
        RECT 43.975 197.115 44.220 197.840 ;
        RECT 44.390 196.945 44.650 197.670 ;
        RECT 44.820 197.115 45.080 197.840 ;
        RECT 45.250 196.945 45.510 197.670 ;
        RECT 45.680 197.115 45.940 197.840 ;
        RECT 46.110 196.945 46.370 197.670 ;
        RECT 46.540 197.115 46.800 197.840 ;
        RECT 46.970 196.945 47.230 197.670 ;
        RECT 47.400 197.045 47.660 197.840 ;
        RECT 41.825 196.930 47.230 196.945 ;
        RECT 40.485 196.705 47.230 196.930 ;
        RECT 40.485 196.115 41.650 196.705 ;
        RECT 47.830 196.535 48.080 197.670 ;
        RECT 48.260 197.035 48.520 197.845 ;
        RECT 48.695 196.535 48.940 197.675 ;
        RECT 49.120 197.035 49.415 197.845 ;
        RECT 49.595 196.705 49.855 197.845 ;
        RECT 41.820 196.285 48.940 196.535 ;
        RECT 40.485 195.945 47.230 196.115 ;
        RECT 37.910 195.465 39.210 195.675 ;
        RECT 39.465 195.295 39.795 195.655 ;
        RECT 39.965 195.465 40.225 195.795 ;
        RECT 40.485 195.295 40.785 195.775 ;
        RECT 40.955 195.490 41.215 195.945 ;
        RECT 41.385 195.295 41.645 195.775 ;
        RECT 41.825 195.490 42.085 195.945 ;
        RECT 42.255 195.295 42.505 195.775 ;
        RECT 42.685 195.490 42.945 195.945 ;
        RECT 43.115 195.295 43.365 195.775 ;
        RECT 43.545 195.490 43.805 195.945 ;
        RECT 43.975 195.295 44.220 195.775 ;
        RECT 44.390 195.490 44.665 195.945 ;
        RECT 44.835 195.295 45.080 195.775 ;
        RECT 45.250 195.490 45.510 195.945 ;
        RECT 45.680 195.295 45.940 195.775 ;
        RECT 46.110 195.490 46.370 195.945 ;
        RECT 46.540 195.295 46.800 195.775 ;
        RECT 46.970 195.490 47.230 195.945 ;
        RECT 47.400 195.295 47.660 195.855 ;
        RECT 47.830 195.475 48.080 196.285 ;
        RECT 48.260 195.295 48.520 195.820 ;
        RECT 48.690 195.475 48.940 196.285 ;
        RECT 49.110 195.975 49.425 196.535 ;
        RECT 49.120 195.295 49.425 195.805 ;
        RECT 49.595 195.295 49.855 196.095 ;
        RECT 50.025 195.465 50.355 197.675 ;
        RECT 50.525 197.335 51.035 197.845 ;
        RECT 52.205 197.165 52.535 197.675 ;
        RECT 50.525 196.995 53.035 197.165 ;
        RECT 50.525 196.205 50.835 196.995 ;
        RECT 51.005 196.205 51.225 196.825 ;
        RECT 51.495 196.205 51.670 196.825 ;
        RECT 51.925 196.205 52.145 196.825 ;
        RECT 52.415 196.655 52.665 196.825 ;
        RECT 52.420 196.205 52.665 196.655 ;
        RECT 52.835 196.035 53.035 196.995 ;
        RECT 53.205 196.705 53.565 197.845 ;
        RECT 54.655 196.680 54.945 197.845 ;
        RECT 55.205 197.100 55.475 197.845 ;
        RECT 56.105 197.840 62.380 197.845 ;
        RECT 55.645 196.930 55.935 197.670 ;
        RECT 56.105 197.115 56.360 197.840 ;
        RECT 56.545 196.945 56.805 197.670 ;
        RECT 56.975 197.115 57.220 197.840 ;
        RECT 57.405 196.945 57.665 197.670 ;
        RECT 57.835 197.115 58.080 197.840 ;
        RECT 58.265 196.945 58.525 197.670 ;
        RECT 58.695 197.115 58.940 197.840 ;
        RECT 59.110 196.945 59.370 197.670 ;
        RECT 59.540 197.115 59.800 197.840 ;
        RECT 59.970 196.945 60.230 197.670 ;
        RECT 60.400 197.115 60.660 197.840 ;
        RECT 60.830 196.945 61.090 197.670 ;
        RECT 61.260 197.115 61.520 197.840 ;
        RECT 61.690 196.945 61.950 197.670 ;
        RECT 62.120 197.045 62.380 197.840 ;
        RECT 56.545 196.930 61.950 196.945 ;
        RECT 55.205 196.705 61.950 196.930 ;
        RECT 53.235 196.455 53.565 196.535 ;
        RECT 53.205 196.285 53.565 196.455 ;
        RECT 55.205 196.145 56.370 196.705 ;
        RECT 62.550 196.535 62.800 197.670 ;
        RECT 62.980 197.035 63.240 197.845 ;
        RECT 63.415 196.535 63.660 197.675 ;
        RECT 63.840 197.035 64.135 197.845 ;
        RECT 64.405 196.875 64.575 197.675 ;
        RECT 64.865 197.215 65.115 197.635 ;
        RECT 65.305 197.385 65.635 197.845 ;
        RECT 65.845 197.215 66.095 197.635 ;
        RECT 64.805 197.045 66.095 197.215 ;
        RECT 66.265 197.045 66.515 197.845 ;
        RECT 66.685 197.215 66.855 197.675 ;
        RECT 67.065 197.385 67.315 197.845 ;
        RECT 66.685 197.045 67.360 197.215 ;
        RECT 64.405 196.705 66.895 196.875 ;
        RECT 56.540 196.285 63.660 196.535 ;
        RECT 55.175 196.115 56.370 196.145 ;
        RECT 50.605 195.295 50.935 196.035 ;
        RECT 51.205 195.865 52.535 196.035 ;
        RECT 51.205 195.465 51.535 195.865 ;
        RECT 51.705 195.295 52.035 195.695 ;
        RECT 52.205 195.635 52.535 195.865 ;
        RECT 52.705 195.805 53.035 196.035 ;
        RECT 53.205 195.635 53.565 196.115 ;
        RECT 52.205 195.465 53.565 195.635 ;
        RECT 54.655 195.295 54.945 196.020 ;
        RECT 55.175 195.975 61.950 196.115 ;
        RECT 55.205 195.945 61.950 195.975 ;
        RECT 55.205 195.295 55.505 195.775 ;
        RECT 55.675 195.490 55.935 195.945 ;
        RECT 56.105 195.295 56.365 195.775 ;
        RECT 56.545 195.490 56.805 195.945 ;
        RECT 56.975 195.295 57.225 195.775 ;
        RECT 57.405 195.490 57.665 195.945 ;
        RECT 57.835 195.295 58.085 195.775 ;
        RECT 58.265 195.490 58.525 195.945 ;
        RECT 58.695 195.295 58.940 195.775 ;
        RECT 59.110 195.490 59.385 195.945 ;
        RECT 59.555 195.295 59.800 195.775 ;
        RECT 59.970 195.490 60.230 195.945 ;
        RECT 60.400 195.295 60.660 195.775 ;
        RECT 60.830 195.490 61.090 195.945 ;
        RECT 61.260 195.295 61.520 195.775 ;
        RECT 61.690 195.490 61.950 195.945 ;
        RECT 62.120 195.295 62.380 195.855 ;
        RECT 62.550 195.475 62.800 196.285 ;
        RECT 62.980 195.295 63.240 195.820 ;
        RECT 63.410 195.475 63.660 196.285 ;
        RECT 63.830 195.975 64.145 196.535 ;
        RECT 64.360 195.965 64.555 196.535 ;
        RECT 63.840 195.295 64.145 195.805 ;
        RECT 64.315 195.295 64.575 195.775 ;
        RECT 64.745 195.715 64.915 196.705 ;
        RECT 65.095 196.080 65.265 196.535 ;
        RECT 65.655 196.455 65.825 196.470 ;
        RECT 65.495 196.285 65.825 196.455 ;
        RECT 65.095 195.910 65.485 196.080 ;
        RECT 64.745 195.545 65.075 195.715 ;
        RECT 65.275 195.625 65.485 195.910 ;
        RECT 65.655 196.075 65.825 196.285 ;
        RECT 66.055 196.205 66.385 196.535 ;
        RECT 66.725 196.455 66.895 196.705 ;
        RECT 66.565 196.285 66.895 196.455 ;
        RECT 65.655 195.905 65.920 196.075 ;
        RECT 66.180 195.970 66.385 196.205 ;
        RECT 67.105 196.095 67.360 197.045 ;
        RECT 67.540 196.700 67.835 197.845 ;
        RECT 65.750 195.805 65.920 195.905 ;
        RECT 66.685 195.925 67.360 196.095 ;
        RECT 65.750 195.635 65.925 195.805 ;
        RECT 66.265 195.675 66.435 195.755 ;
        RECT 65.750 195.610 65.920 195.635 ;
        RECT 64.745 195.465 64.990 195.545 ;
        RECT 66.165 195.295 66.495 195.675 ;
        RECT 66.685 195.465 66.855 195.925 ;
        RECT 67.105 195.295 67.360 195.755 ;
        RECT 67.540 195.295 67.835 196.115 ;
        RECT 68.005 195.845 68.235 197.545 ;
        RECT 68.450 197.040 68.705 197.845 ;
        RECT 68.905 197.230 69.235 197.675 ;
        RECT 69.405 197.400 69.680 197.845 ;
        RECT 69.915 197.230 70.245 197.675 ;
        RECT 68.905 197.050 70.245 197.230 ;
        RECT 70.705 196.870 71.035 197.535 ;
        RECT 71.305 197.100 71.575 197.845 ;
        RECT 72.205 197.840 78.480 197.845 ;
        RECT 71.745 196.930 72.035 197.670 ;
        RECT 72.205 197.115 72.460 197.840 ;
        RECT 72.645 196.945 72.905 197.670 ;
        RECT 73.075 197.115 73.320 197.840 ;
        RECT 73.505 196.945 73.765 197.670 ;
        RECT 73.935 197.115 74.180 197.840 ;
        RECT 74.365 196.945 74.625 197.670 ;
        RECT 74.795 197.115 75.040 197.840 ;
        RECT 75.210 196.945 75.470 197.670 ;
        RECT 75.640 197.115 75.900 197.840 ;
        RECT 76.070 196.945 76.330 197.670 ;
        RECT 76.500 197.115 76.760 197.840 ;
        RECT 76.930 196.945 77.190 197.670 ;
        RECT 77.360 197.115 77.620 197.840 ;
        RECT 77.790 196.945 78.050 197.670 ;
        RECT 78.220 197.045 78.480 197.840 ;
        RECT 72.645 196.930 78.050 196.945 ;
        RECT 68.450 196.700 71.035 196.870 ;
        RECT 71.305 196.705 78.050 196.930 ;
        RECT 68.450 196.085 68.760 196.700 ;
        RECT 68.930 196.255 69.260 196.485 ;
        RECT 69.430 196.255 69.900 196.485 ;
        RECT 70.070 196.315 70.525 196.485 ;
        RECT 70.070 196.255 70.520 196.315 ;
        RECT 70.710 196.255 71.045 196.485 ;
        RECT 71.305 196.115 72.470 196.705 ;
        RECT 78.650 196.535 78.900 197.670 ;
        RECT 79.080 197.035 79.340 197.845 ;
        RECT 79.515 196.535 79.760 197.675 ;
        RECT 79.940 197.035 80.235 197.845 ;
        RECT 80.415 196.680 80.705 197.845 ;
        RECT 80.895 197.255 81.135 197.645 ;
        RECT 81.305 197.435 81.655 197.845 ;
        RECT 80.895 197.055 81.645 197.255 ;
        RECT 72.640 196.285 79.760 196.535 ;
        RECT 68.450 195.905 71.035 196.085 ;
        RECT 71.305 195.945 78.050 196.115 ;
        RECT 68.005 195.465 68.225 195.845 ;
        RECT 68.395 195.295 69.245 195.655 ;
        RECT 69.725 195.485 70.055 195.905 ;
        RECT 70.260 195.295 70.535 195.735 ;
        RECT 70.705 195.485 71.035 195.905 ;
        RECT 71.305 195.295 71.605 195.775 ;
        RECT 71.775 195.490 72.035 195.945 ;
        RECT 72.205 195.295 72.465 195.775 ;
        RECT 72.645 195.490 72.905 195.945 ;
        RECT 73.075 195.295 73.325 195.775 ;
        RECT 73.505 195.490 73.765 195.945 ;
        RECT 73.935 195.295 74.185 195.775 ;
        RECT 74.365 195.490 74.625 195.945 ;
        RECT 74.795 195.295 75.040 195.775 ;
        RECT 75.210 195.490 75.485 195.945 ;
        RECT 75.655 195.295 75.900 195.775 ;
        RECT 76.070 195.490 76.330 195.945 ;
        RECT 76.500 195.295 76.760 195.775 ;
        RECT 76.930 195.490 77.190 195.945 ;
        RECT 77.360 195.295 77.620 195.775 ;
        RECT 77.790 195.490 78.050 195.945 ;
        RECT 78.220 195.295 78.480 195.855 ;
        RECT 78.650 195.475 78.900 196.285 ;
        RECT 79.080 195.295 79.340 195.820 ;
        RECT 79.510 195.475 79.760 196.285 ;
        RECT 79.930 195.975 80.245 196.535 ;
        RECT 79.940 195.295 80.245 195.805 ;
        RECT 80.415 195.295 80.705 196.020 ;
        RECT 80.895 195.535 81.125 196.875 ;
        RECT 81.305 196.375 81.645 197.055 ;
        RECT 81.825 196.555 82.155 197.665 ;
        RECT 82.325 197.195 82.505 197.665 ;
        RECT 82.675 197.365 83.005 197.845 ;
        RECT 83.180 197.195 83.350 197.665 ;
        RECT 82.325 196.995 83.350 197.195 ;
        RECT 81.305 195.475 81.535 196.375 ;
        RECT 81.825 196.255 82.370 196.555 ;
        RECT 81.735 195.295 81.980 196.075 ;
        RECT 82.150 196.025 82.370 196.255 ;
        RECT 82.540 196.205 82.965 196.825 ;
        RECT 83.160 196.205 83.420 196.825 ;
        RECT 83.615 196.705 83.900 197.845 ;
        RECT 83.630 196.025 83.890 196.535 ;
        RECT 82.150 195.835 83.890 196.025 ;
        RECT 82.150 195.475 82.580 195.835 ;
        RECT 83.160 195.295 83.890 195.665 ;
        RECT 84.090 195.475 84.370 197.665 ;
        RECT 84.595 196.705 84.825 197.845 ;
        RECT 84.995 196.695 85.325 197.675 ;
        RECT 85.495 196.705 85.705 197.845 ;
        RECT 85.935 196.755 87.145 197.845 ;
        RECT 84.575 196.285 84.905 196.535 ;
        RECT 84.595 195.295 84.825 196.115 ;
        RECT 85.075 196.095 85.325 196.695 ;
        RECT 85.935 196.215 86.455 196.755 ;
        RECT 84.995 195.465 85.325 196.095 ;
        RECT 85.495 195.295 85.705 196.115 ;
        RECT 86.625 196.045 87.145 196.585 ;
        RECT 85.935 195.295 87.145 196.045 ;
        RECT 15.930 195.125 87.230 195.295 ;
        RECT 16.015 194.375 17.225 195.125 ;
        RECT 16.015 193.835 16.535 194.375 ;
        RECT 17.400 194.285 17.660 195.125 ;
        RECT 17.835 194.380 18.090 194.955 ;
        RECT 18.260 194.745 18.590 195.125 ;
        RECT 18.805 194.575 18.975 194.955 ;
        RECT 18.260 194.405 18.975 194.575 ;
        RECT 19.325 194.575 19.495 194.955 ;
        RECT 19.675 194.745 20.005 195.125 ;
        RECT 19.325 194.405 19.990 194.575 ;
        RECT 20.185 194.450 20.445 194.955 ;
        RECT 16.705 193.665 17.225 194.205 ;
        RECT 16.015 192.575 17.225 193.665 ;
        RECT 17.400 192.575 17.660 193.725 ;
        RECT 17.835 193.650 18.005 194.380 ;
        RECT 18.260 194.215 18.430 194.405 ;
        RECT 18.175 193.885 18.430 194.215 ;
        RECT 18.260 193.675 18.430 193.885 ;
        RECT 18.710 193.855 19.065 194.225 ;
        RECT 19.255 193.855 19.595 194.225 ;
        RECT 19.820 194.150 19.990 194.405 ;
        RECT 19.820 193.820 20.095 194.150 ;
        RECT 19.820 193.675 19.990 193.820 ;
        RECT 17.835 192.745 18.090 193.650 ;
        RECT 18.260 193.505 18.975 193.675 ;
        RECT 18.260 192.575 18.590 193.335 ;
        RECT 18.805 192.745 18.975 193.505 ;
        RECT 19.315 193.505 19.990 193.675 ;
        RECT 20.265 193.650 20.445 194.450 ;
        RECT 19.315 192.745 19.495 193.505 ;
        RECT 19.675 192.575 20.005 193.335 ;
        RECT 20.175 192.745 20.445 193.650 ;
        RECT 20.615 194.450 20.875 194.955 ;
        RECT 21.055 194.745 21.385 195.125 ;
        RECT 21.565 194.575 21.735 194.955 ;
        RECT 20.615 193.650 20.785 194.450 ;
        RECT 21.070 194.405 21.735 194.575 ;
        RECT 21.070 194.150 21.240 194.405 ;
        RECT 22.055 194.305 22.265 195.125 ;
        RECT 22.435 194.325 22.765 194.955 ;
        RECT 20.955 193.820 21.240 194.150 ;
        RECT 21.475 193.855 21.805 194.225 ;
        RECT 21.070 193.675 21.240 193.820 ;
        RECT 22.435 193.725 22.685 194.325 ;
        RECT 22.935 194.305 23.165 195.125 ;
        RECT 22.855 193.885 23.185 194.135 ;
        RECT 20.615 192.745 20.885 193.650 ;
        RECT 21.070 193.505 21.735 193.675 ;
        RECT 21.055 192.575 21.385 193.335 ;
        RECT 21.565 192.745 21.735 193.505 ;
        RECT 22.055 192.575 22.265 193.715 ;
        RECT 22.435 192.745 22.765 193.725 ;
        RECT 22.935 192.575 23.165 193.715 ;
        RECT 23.845 192.755 24.105 194.945 ;
        RECT 24.365 194.755 25.035 195.125 ;
        RECT 25.215 194.575 25.525 194.945 ;
        RECT 24.295 194.375 25.525 194.575 ;
        RECT 24.295 193.705 24.585 194.375 ;
        RECT 25.705 194.195 25.935 194.835 ;
        RECT 26.115 194.395 26.405 195.125 ;
        RECT 26.630 194.385 27.245 194.955 ;
        RECT 27.415 194.615 27.630 195.125 ;
        RECT 27.860 194.615 28.140 194.945 ;
        RECT 28.320 194.615 28.560 195.125 ;
        RECT 24.765 193.885 25.230 194.195 ;
        RECT 25.410 193.885 25.935 194.195 ;
        RECT 26.115 193.885 26.415 194.215 ;
        RECT 24.295 193.485 25.065 193.705 ;
        RECT 24.275 192.575 24.615 193.305 ;
        RECT 24.795 192.755 25.065 193.485 ;
        RECT 25.245 193.465 26.405 193.705 ;
        RECT 25.245 192.755 25.475 193.465 ;
        RECT 25.645 192.575 25.975 193.285 ;
        RECT 26.145 192.755 26.405 193.465 ;
        RECT 26.630 193.365 26.945 194.385 ;
        RECT 27.115 193.715 27.285 194.215 ;
        RECT 27.535 193.885 27.800 194.445 ;
        RECT 27.970 193.715 28.140 194.615 ;
        RECT 29.445 194.575 29.615 194.955 ;
        RECT 29.795 194.745 30.125 195.125 ;
        RECT 28.310 193.885 28.665 194.445 ;
        RECT 29.445 194.405 30.110 194.575 ;
        RECT 30.305 194.450 30.565 194.955 ;
        RECT 29.375 193.855 29.715 194.225 ;
        RECT 29.940 194.150 30.110 194.405 ;
        RECT 29.940 193.820 30.215 194.150 ;
        RECT 27.115 193.545 28.540 193.715 ;
        RECT 29.940 193.675 30.110 193.820 ;
        RECT 26.630 192.745 27.165 193.365 ;
        RECT 27.335 192.575 27.665 193.375 ;
        RECT 28.150 193.370 28.540 193.545 ;
        RECT 29.435 193.505 30.110 193.675 ;
        RECT 30.385 193.650 30.565 194.450 ;
        RECT 30.745 194.395 31.045 195.125 ;
        RECT 31.225 194.215 31.455 194.835 ;
        RECT 31.655 194.565 31.880 194.945 ;
        RECT 32.050 194.735 32.380 195.125 ;
        RECT 33.495 194.665 34.055 194.955 ;
        RECT 34.225 194.665 34.475 195.125 ;
        RECT 31.655 194.385 31.985 194.565 ;
        RECT 30.750 193.885 31.045 194.215 ;
        RECT 31.225 193.885 31.640 194.215 ;
        RECT 31.810 193.715 31.985 194.385 ;
        RECT 32.155 193.885 32.395 194.535 ;
        RECT 29.435 192.745 29.615 193.505 ;
        RECT 29.795 192.575 30.125 193.335 ;
        RECT 30.295 192.745 30.565 193.650 ;
        RECT 30.745 193.355 31.640 193.685 ;
        RECT 31.810 193.525 32.395 193.715 ;
        RECT 30.745 193.185 31.950 193.355 ;
        RECT 30.745 192.755 31.075 193.185 ;
        RECT 31.255 192.575 31.450 193.015 ;
        RECT 31.620 192.755 31.950 193.185 ;
        RECT 32.120 192.755 32.395 193.525 ;
        RECT 33.495 193.295 33.745 194.665 ;
        RECT 35.095 194.495 35.425 194.855 ;
        RECT 35.800 194.620 36.135 195.125 ;
        RECT 36.305 194.555 36.545 194.930 ;
        RECT 36.825 194.795 36.995 194.940 ;
        RECT 36.825 194.600 37.200 194.795 ;
        RECT 37.560 194.630 37.955 195.125 ;
        RECT 34.035 194.305 35.425 194.495 ;
        RECT 34.035 194.215 34.205 194.305 ;
        RECT 33.915 193.885 34.205 194.215 ;
        RECT 34.375 193.885 34.715 194.135 ;
        RECT 34.935 193.885 35.610 194.135 ;
        RECT 34.035 193.635 34.205 193.885 ;
        RECT 34.035 193.465 34.975 193.635 ;
        RECT 35.345 193.525 35.610 193.885 ;
        RECT 35.855 193.595 36.155 194.445 ;
        RECT 36.325 194.405 36.545 194.555 ;
        RECT 36.325 194.075 36.860 194.405 ;
        RECT 37.030 194.265 37.200 194.600 ;
        RECT 38.125 194.435 38.365 194.955 ;
        RECT 39.015 194.745 39.345 195.125 ;
        RECT 33.495 192.745 33.955 193.295 ;
        RECT 34.145 192.575 34.475 193.295 ;
        RECT 34.675 192.915 34.975 193.465 ;
        RECT 36.325 193.425 36.560 194.075 ;
        RECT 37.030 193.905 38.015 194.265 ;
        RECT 35.145 192.575 35.425 193.245 ;
        RECT 35.885 193.195 36.560 193.425 ;
        RECT 36.730 193.885 38.015 193.905 ;
        RECT 36.730 193.735 37.590 193.885 ;
        RECT 35.885 192.765 36.055 193.195 ;
        RECT 36.225 192.575 36.555 193.025 ;
        RECT 36.730 192.790 37.015 193.735 ;
        RECT 38.190 193.630 38.365 194.435 ;
        RECT 38.570 194.575 38.845 194.715 ;
        RECT 39.515 194.575 39.725 194.745 ;
        RECT 38.570 194.385 39.725 194.575 ;
        RECT 39.895 194.575 40.225 194.955 ;
        RECT 40.415 194.745 40.745 195.125 ;
        RECT 39.895 194.370 40.745 194.575 ;
        RECT 38.565 193.760 38.825 194.215 ;
        RECT 39.080 193.810 39.665 194.185 ;
        RECT 37.190 193.255 37.885 193.565 ;
        RECT 37.195 192.575 37.880 193.045 ;
        RECT 38.060 192.845 38.365 193.630 ;
        RECT 38.570 192.575 38.895 193.560 ;
        RECT 39.080 193.425 39.285 193.810 ;
        RECT 39.835 193.595 40.245 194.200 ;
        RECT 40.415 193.880 40.745 194.370 ;
        RECT 40.415 193.425 40.585 193.880 ;
        RECT 39.075 193.255 39.285 193.425 ;
        RECT 39.080 193.225 39.285 193.255 ;
        RECT 39.465 193.205 40.585 193.425 ;
        RECT 39.465 192.745 39.725 193.205 ;
        RECT 39.895 192.575 40.745 193.025 ;
        RECT 40.915 192.745 41.160 194.955 ;
        RECT 41.345 194.325 41.585 195.125 ;
        RECT 41.775 194.400 42.065 195.125 ;
        RECT 42.235 194.625 42.495 194.955 ;
        RECT 42.665 194.765 42.995 195.125 ;
        RECT 43.250 194.745 44.550 194.955 ;
        RECT 41.345 192.575 41.600 193.575 ;
        RECT 41.775 192.575 42.065 193.740 ;
        RECT 42.235 193.425 42.405 194.625 ;
        RECT 43.250 194.595 43.420 194.745 ;
        RECT 42.665 194.470 43.420 194.595 ;
        RECT 42.575 194.425 43.420 194.470 ;
        RECT 42.575 194.305 42.845 194.425 ;
        RECT 42.575 193.730 42.745 194.305 ;
        RECT 42.975 193.865 43.385 194.170 ;
        RECT 43.675 194.135 43.885 194.535 ;
        RECT 43.555 193.925 43.885 194.135 ;
        RECT 44.130 194.135 44.350 194.535 ;
        RECT 44.825 194.360 45.280 195.125 ;
        RECT 44.130 193.925 44.605 194.135 ;
        RECT 44.795 193.935 45.285 194.135 ;
        RECT 42.575 193.695 42.775 193.730 ;
        RECT 44.105 193.695 45.280 193.755 ;
        RECT 42.575 193.585 45.280 193.695 ;
        RECT 42.635 193.525 44.435 193.585 ;
        RECT 44.105 193.495 44.435 193.525 ;
        RECT 42.235 192.745 42.495 193.425 ;
        RECT 42.665 192.575 42.915 193.355 ;
        RECT 43.165 193.325 44.000 193.335 ;
        RECT 44.590 193.325 44.775 193.415 ;
        RECT 43.165 193.125 44.775 193.325 ;
        RECT 43.165 192.745 43.415 193.125 ;
        RECT 44.545 193.085 44.775 193.125 ;
        RECT 45.025 192.965 45.280 193.585 ;
        RECT 43.585 192.575 43.940 192.955 ;
        RECT 44.945 192.745 45.280 192.965 ;
        RECT 45.455 192.745 45.735 194.845 ;
        RECT 45.965 194.665 46.135 195.125 ;
        RECT 46.405 194.735 47.655 194.915 ;
        RECT 46.790 194.495 47.155 194.565 ;
        RECT 45.905 194.315 47.155 194.495 ;
        RECT 47.325 194.515 47.655 194.735 ;
        RECT 47.825 194.685 47.995 195.125 ;
        RECT 48.165 194.515 48.505 194.930 ;
        RECT 48.765 194.645 49.065 195.125 ;
        RECT 47.325 194.345 48.505 194.515 ;
        RECT 49.235 194.475 49.495 194.930 ;
        RECT 49.665 194.645 49.925 195.125 ;
        RECT 50.105 194.475 50.365 194.930 ;
        RECT 50.535 194.645 50.785 195.125 ;
        RECT 50.965 194.475 51.225 194.930 ;
        RECT 51.395 194.645 51.645 195.125 ;
        RECT 51.825 194.475 52.085 194.930 ;
        RECT 52.255 194.645 52.500 195.125 ;
        RECT 52.670 194.475 52.945 194.930 ;
        RECT 53.115 194.645 53.360 195.125 ;
        RECT 53.530 194.475 53.790 194.930 ;
        RECT 53.960 194.645 54.220 195.125 ;
        RECT 54.390 194.475 54.650 194.930 ;
        RECT 54.820 194.645 55.080 195.125 ;
        RECT 55.250 194.475 55.510 194.930 ;
        RECT 55.680 194.565 55.940 195.125 ;
        RECT 45.905 193.715 46.180 194.315 ;
        RECT 48.765 194.305 55.510 194.475 ;
        RECT 46.350 193.885 46.705 194.135 ;
        RECT 46.900 194.105 47.365 194.135 ;
        RECT 46.895 193.935 47.365 194.105 ;
        RECT 46.900 193.885 47.365 193.935 ;
        RECT 47.535 193.885 47.865 194.135 ;
        RECT 48.040 193.935 48.505 194.135 ;
        RECT 47.685 193.765 47.865 193.885 ;
        RECT 45.905 193.505 47.515 193.715 ;
        RECT 47.685 193.595 48.015 193.765 ;
        RECT 47.105 193.405 47.515 193.505 ;
        RECT 45.925 192.575 46.710 193.335 ;
        RECT 47.105 192.745 47.490 193.405 ;
        RECT 47.815 192.805 48.015 193.595 ;
        RECT 48.185 192.575 48.505 193.755 ;
        RECT 48.765 193.715 49.930 194.305 ;
        RECT 56.110 194.135 56.360 194.945 ;
        RECT 56.540 194.600 56.800 195.125 ;
        RECT 56.970 194.135 57.220 194.945 ;
        RECT 57.400 194.615 57.705 195.125 ;
        RECT 58.425 194.645 58.725 195.125 ;
        RECT 58.895 194.475 59.155 194.930 ;
        RECT 59.325 194.645 59.585 195.125 ;
        RECT 59.765 194.475 60.025 194.930 ;
        RECT 60.195 194.645 60.445 195.125 ;
        RECT 60.625 194.475 60.885 194.930 ;
        RECT 61.055 194.645 61.305 195.125 ;
        RECT 61.485 194.475 61.745 194.930 ;
        RECT 61.915 194.645 62.160 195.125 ;
        RECT 62.330 194.475 62.605 194.930 ;
        RECT 62.775 194.645 63.020 195.125 ;
        RECT 63.190 194.475 63.450 194.930 ;
        RECT 63.620 194.645 63.880 195.125 ;
        RECT 64.050 194.475 64.310 194.930 ;
        RECT 64.480 194.645 64.740 195.125 ;
        RECT 64.910 194.475 65.170 194.930 ;
        RECT 65.340 194.565 65.600 195.125 ;
        RECT 50.100 193.885 57.220 194.135 ;
        RECT 57.390 193.885 57.705 194.445 ;
        RECT 58.425 194.305 65.170 194.475 ;
        RECT 48.765 193.490 55.510 193.715 ;
        RECT 48.765 192.575 49.035 193.320 ;
        RECT 49.205 192.750 49.495 193.490 ;
        RECT 50.105 193.475 55.510 193.490 ;
        RECT 49.665 192.580 49.920 193.305 ;
        RECT 50.105 192.750 50.365 193.475 ;
        RECT 50.535 192.580 50.780 193.305 ;
        RECT 50.965 192.750 51.225 193.475 ;
        RECT 51.395 192.580 51.640 193.305 ;
        RECT 51.825 192.750 52.085 193.475 ;
        RECT 52.255 192.580 52.500 193.305 ;
        RECT 52.670 192.750 52.930 193.475 ;
        RECT 53.100 192.580 53.360 193.305 ;
        RECT 53.530 192.750 53.790 193.475 ;
        RECT 53.960 192.580 54.220 193.305 ;
        RECT 54.390 192.750 54.650 193.475 ;
        RECT 54.820 192.580 55.080 193.305 ;
        RECT 55.250 192.750 55.510 193.475 ;
        RECT 55.680 192.580 55.940 193.375 ;
        RECT 56.110 192.750 56.360 193.885 ;
        RECT 49.665 192.575 55.940 192.580 ;
        RECT 56.540 192.575 56.800 193.385 ;
        RECT 56.975 192.745 57.220 193.885 ;
        RECT 58.425 193.715 59.590 194.305 ;
        RECT 65.770 194.135 66.020 194.945 ;
        RECT 66.200 194.600 66.460 195.125 ;
        RECT 66.630 194.135 66.880 194.945 ;
        RECT 67.060 194.615 67.365 195.125 ;
        RECT 59.760 193.885 66.880 194.135 ;
        RECT 67.050 193.885 67.365 194.445 ;
        RECT 67.535 194.400 67.825 195.125 ;
        RECT 67.995 194.475 68.255 194.920 ;
        RECT 68.505 194.645 68.675 195.125 ;
        RECT 68.845 194.615 69.195 194.945 ;
        RECT 69.430 194.645 69.600 195.125 ;
        RECT 67.995 194.305 68.675 194.475 ;
        RECT 58.425 193.490 65.170 193.715 ;
        RECT 57.400 192.575 57.695 193.385 ;
        RECT 58.425 192.575 58.695 193.320 ;
        RECT 58.865 192.750 59.155 193.490 ;
        RECT 59.765 193.475 65.170 193.490 ;
        RECT 59.325 192.580 59.580 193.305 ;
        RECT 59.765 192.750 60.025 193.475 ;
        RECT 60.195 192.580 60.440 193.305 ;
        RECT 60.625 192.750 60.885 193.475 ;
        RECT 61.055 192.580 61.300 193.305 ;
        RECT 61.485 192.750 61.745 193.475 ;
        RECT 61.915 192.580 62.160 193.305 ;
        RECT 62.330 192.750 62.590 193.475 ;
        RECT 62.760 192.580 63.020 193.305 ;
        RECT 63.190 192.750 63.450 193.475 ;
        RECT 63.620 192.580 63.880 193.305 ;
        RECT 64.050 192.750 64.310 193.475 ;
        RECT 64.480 192.580 64.740 193.305 ;
        RECT 64.910 192.750 65.170 193.475 ;
        RECT 65.340 192.580 65.600 193.375 ;
        RECT 65.770 192.750 66.020 193.885 ;
        RECT 59.325 192.575 65.600 192.580 ;
        RECT 66.200 192.575 66.460 193.385 ;
        RECT 66.635 192.745 66.880 193.885 ;
        RECT 67.060 192.575 67.355 193.385 ;
        RECT 67.535 192.575 67.825 193.740 ;
        RECT 67.995 193.570 68.335 194.135 ;
        RECT 68.505 193.400 68.675 194.305 ;
        RECT 68.845 193.715 69.015 194.615 ;
        RECT 69.900 194.555 70.070 194.905 ;
        RECT 70.240 194.725 70.570 195.125 ;
        RECT 70.740 194.605 70.995 194.905 ;
        RECT 70.740 194.555 71.045 194.605 ;
        RECT 69.900 194.475 71.045 194.555 ;
        RECT 69.335 194.445 71.045 194.475 ;
        RECT 69.185 194.385 71.045 194.445 ;
        RECT 69.185 194.305 70.070 194.385 ;
        RECT 69.185 194.275 69.505 194.305 ;
        RECT 69.185 193.885 69.355 194.275 ;
        RECT 68.845 193.510 69.240 193.715 ;
        RECT 69.605 193.595 70.140 194.135 ;
        RECT 70.400 193.885 70.700 194.215 ;
        RECT 70.400 193.425 70.570 193.885 ;
        RECT 70.875 193.715 71.045 194.385 ;
        RECT 71.675 194.325 71.935 195.125 ;
        RECT 67.995 193.340 68.675 193.400 ;
        RECT 69.460 193.340 70.570 193.425 ;
        RECT 67.995 193.255 70.570 193.340 ;
        RECT 70.740 193.285 71.045 193.715 ;
        RECT 67.995 193.170 69.630 193.255 ;
        RECT 67.995 192.990 68.255 193.170 ;
        RECT 68.460 192.575 68.820 193.000 ;
        RECT 69.335 192.575 69.665 193.000 ;
        RECT 69.845 192.845 71.045 193.085 ;
        RECT 71.675 192.575 71.935 193.715 ;
        RECT 72.105 192.745 72.435 194.955 ;
        RECT 72.685 194.385 73.015 195.125 ;
        RECT 73.285 194.555 73.615 194.955 ;
        RECT 73.785 194.725 74.115 195.125 ;
        RECT 74.285 194.785 75.645 194.955 ;
        RECT 74.285 194.555 74.615 194.785 ;
        RECT 73.285 194.385 74.615 194.555 ;
        RECT 74.785 194.385 75.115 194.615 ;
        RECT 72.605 193.425 72.915 194.215 ;
        RECT 73.085 193.595 73.305 194.215 ;
        RECT 73.575 193.595 73.750 194.215 ;
        RECT 74.005 193.595 74.225 194.215 ;
        RECT 74.500 194.105 74.745 194.215 ;
        RECT 74.495 193.935 74.745 194.105 ;
        RECT 74.500 193.595 74.745 193.935 ;
        RECT 74.915 193.425 75.115 194.385 ;
        RECT 75.285 194.305 75.645 194.785 ;
        RECT 76.825 194.645 77.125 195.125 ;
        RECT 77.295 194.475 77.555 194.930 ;
        RECT 77.725 194.645 77.985 195.125 ;
        RECT 78.165 194.475 78.425 194.930 ;
        RECT 78.595 194.645 78.845 195.125 ;
        RECT 79.025 194.475 79.285 194.930 ;
        RECT 79.455 194.645 79.705 195.125 ;
        RECT 79.885 194.475 80.145 194.930 ;
        RECT 80.315 194.645 80.560 195.125 ;
        RECT 80.730 194.475 81.005 194.930 ;
        RECT 81.175 194.645 81.420 195.125 ;
        RECT 81.590 194.475 81.850 194.930 ;
        RECT 82.020 194.645 82.280 195.125 ;
        RECT 82.450 194.475 82.710 194.930 ;
        RECT 82.880 194.645 83.140 195.125 ;
        RECT 83.310 194.475 83.570 194.930 ;
        RECT 83.740 194.565 84.000 195.125 ;
        RECT 76.825 194.305 83.570 194.475 ;
        RECT 75.285 193.965 75.645 194.135 ;
        RECT 75.315 193.885 75.645 193.965 ;
        RECT 76.825 193.715 77.990 194.305 ;
        RECT 84.170 194.135 84.420 194.945 ;
        RECT 84.600 194.600 84.860 195.125 ;
        RECT 85.030 194.135 85.280 194.945 ;
        RECT 85.460 194.615 85.765 195.125 ;
        RECT 78.160 193.885 85.280 194.135 ;
        RECT 85.450 193.885 85.765 194.445 ;
        RECT 85.935 194.375 87.145 195.125 ;
        RECT 72.605 193.255 75.115 193.425 ;
        RECT 72.605 192.575 73.115 193.085 ;
        RECT 74.285 192.745 74.615 193.255 ;
        RECT 75.285 192.575 75.645 193.715 ;
        RECT 76.825 193.490 83.570 193.715 ;
        RECT 76.825 192.575 77.095 193.320 ;
        RECT 77.265 192.750 77.555 193.490 ;
        RECT 78.165 193.475 83.570 193.490 ;
        RECT 77.725 192.580 77.980 193.305 ;
        RECT 78.165 192.750 78.425 193.475 ;
        RECT 78.595 192.580 78.840 193.305 ;
        RECT 79.025 192.750 79.285 193.475 ;
        RECT 79.455 192.580 79.700 193.305 ;
        RECT 79.885 192.750 80.145 193.475 ;
        RECT 80.315 192.580 80.560 193.305 ;
        RECT 80.730 192.750 80.990 193.475 ;
        RECT 81.160 192.580 81.420 193.305 ;
        RECT 81.590 192.750 81.850 193.475 ;
        RECT 82.020 192.580 82.280 193.305 ;
        RECT 82.450 192.750 82.710 193.475 ;
        RECT 82.880 192.580 83.140 193.305 ;
        RECT 83.310 192.750 83.570 193.475 ;
        RECT 83.740 192.580 84.000 193.375 ;
        RECT 84.170 192.750 84.420 193.885 ;
        RECT 77.725 192.575 84.000 192.580 ;
        RECT 84.600 192.575 84.860 193.385 ;
        RECT 85.035 192.745 85.280 193.885 ;
        RECT 85.935 193.665 86.455 194.205 ;
        RECT 86.625 193.835 87.145 194.375 ;
        RECT 85.460 192.575 85.755 193.385 ;
        RECT 85.935 192.575 87.145 193.665 ;
        RECT 15.930 192.405 87.230 192.575 ;
        RECT 16.015 191.315 17.225 192.405 ;
        RECT 16.015 190.605 16.535 191.145 ;
        RECT 16.705 190.775 17.225 191.315 ;
        RECT 18.315 191.330 18.585 192.235 ;
        RECT 18.755 191.645 19.085 192.405 ;
        RECT 19.265 191.475 19.435 192.235 ;
        RECT 16.015 189.855 17.225 190.605 ;
        RECT 18.315 190.530 18.485 191.330 ;
        RECT 18.770 191.305 19.435 191.475 ;
        RECT 19.695 191.330 19.965 192.235 ;
        RECT 20.135 191.645 20.465 192.405 ;
        RECT 20.645 191.475 20.815 192.235 ;
        RECT 18.770 191.160 18.940 191.305 ;
        RECT 18.655 190.830 18.940 191.160 ;
        RECT 18.770 190.575 18.940 190.830 ;
        RECT 19.175 190.755 19.505 191.125 ;
        RECT 18.315 190.025 18.575 190.530 ;
        RECT 18.770 190.405 19.435 190.575 ;
        RECT 18.755 189.855 19.085 190.235 ;
        RECT 19.265 190.025 19.435 190.405 ;
        RECT 19.695 190.530 19.865 191.330 ;
        RECT 20.150 191.305 20.815 191.475 ;
        RECT 21.075 191.330 21.345 192.235 ;
        RECT 21.515 191.645 21.845 192.405 ;
        RECT 22.025 191.475 22.195 192.235 ;
        RECT 22.645 191.680 22.975 192.405 ;
        RECT 20.150 191.160 20.320 191.305 ;
        RECT 20.035 190.830 20.320 191.160 ;
        RECT 20.150 190.575 20.320 190.830 ;
        RECT 20.555 190.755 20.885 191.125 ;
        RECT 19.695 190.025 19.955 190.530 ;
        RECT 20.150 190.405 20.815 190.575 ;
        RECT 20.135 189.855 20.465 190.235 ;
        RECT 20.645 190.025 20.815 190.405 ;
        RECT 21.075 190.530 21.245 191.330 ;
        RECT 21.530 191.305 22.195 191.475 ;
        RECT 21.530 191.160 21.700 191.305 ;
        RECT 21.415 190.830 21.700 191.160 ;
        RECT 21.530 190.575 21.700 190.830 ;
        RECT 21.935 190.755 22.265 191.125 ;
        RECT 21.075 190.025 21.335 190.530 ;
        RECT 21.530 190.405 22.195 190.575 ;
        RECT 21.515 189.855 21.845 190.235 ;
        RECT 22.025 190.025 22.195 190.405 ;
        RECT 22.455 190.025 22.975 191.510 ;
        RECT 23.145 190.685 23.665 192.235 ;
        RECT 24.020 191.435 24.410 191.610 ;
        RECT 24.895 191.605 25.225 192.405 ;
        RECT 25.395 191.615 25.930 192.235 ;
        RECT 24.020 191.265 25.445 191.435 ;
        RECT 23.895 190.535 24.250 191.095 ;
        RECT 23.145 189.855 23.485 190.515 ;
        RECT 24.420 190.365 24.590 191.265 ;
        RECT 24.760 190.535 25.025 191.095 ;
        RECT 25.275 190.765 25.445 191.265 ;
        RECT 25.615 190.595 25.930 191.615 ;
        RECT 26.140 191.255 26.400 192.405 ;
        RECT 26.575 191.330 26.830 192.235 ;
        RECT 27.000 191.645 27.330 192.405 ;
        RECT 27.545 191.475 27.715 192.235 ;
        RECT 24.000 189.855 24.240 190.365 ;
        RECT 24.420 190.035 24.700 190.365 ;
        RECT 24.930 189.855 25.145 190.365 ;
        RECT 25.315 190.025 25.930 190.595 ;
        RECT 26.140 189.855 26.400 190.695 ;
        RECT 26.575 190.600 26.745 191.330 ;
        RECT 27.000 191.305 27.715 191.475 ;
        RECT 27.000 191.095 27.170 191.305 ;
        RECT 28.895 191.240 29.185 192.405 ;
        RECT 30.280 191.265 30.615 192.235 ;
        RECT 30.785 191.265 30.955 192.405 ;
        RECT 31.125 192.065 33.155 192.235 ;
        RECT 26.915 190.765 27.170 191.095 ;
        RECT 26.575 190.025 26.830 190.600 ;
        RECT 27.000 190.575 27.170 190.765 ;
        RECT 27.450 190.755 27.805 191.125 ;
        RECT 30.280 190.595 30.450 191.265 ;
        RECT 31.125 191.095 31.295 192.065 ;
        RECT 30.620 190.765 30.875 191.095 ;
        RECT 31.100 190.765 31.295 191.095 ;
        RECT 31.465 191.725 32.590 191.895 ;
        RECT 30.705 190.595 30.875 190.765 ;
        RECT 31.465 190.595 31.635 191.725 ;
        RECT 27.000 190.405 27.715 190.575 ;
        RECT 27.000 189.855 27.330 190.235 ;
        RECT 27.545 190.025 27.715 190.405 ;
        RECT 28.895 189.855 29.185 190.580 ;
        RECT 30.280 190.025 30.535 190.595 ;
        RECT 30.705 190.425 31.635 190.595 ;
        RECT 31.805 191.385 32.815 191.555 ;
        RECT 31.805 190.585 31.975 191.385 ;
        RECT 31.460 190.390 31.635 190.425 ;
        RECT 30.705 189.855 31.035 190.255 ;
        RECT 31.460 190.025 31.990 190.390 ;
        RECT 32.180 190.365 32.455 191.185 ;
        RECT 32.175 190.195 32.455 190.365 ;
        RECT 32.180 190.025 32.455 190.195 ;
        RECT 32.625 190.025 32.815 191.385 ;
        RECT 32.985 191.400 33.155 192.065 ;
        RECT 33.325 191.645 33.495 192.405 ;
        RECT 33.730 191.645 34.245 192.055 ;
        RECT 32.985 191.210 33.735 191.400 ;
        RECT 33.905 190.835 34.245 191.645 ;
        RECT 34.965 191.475 35.135 192.235 ;
        RECT 35.315 191.645 35.645 192.405 ;
        RECT 34.965 191.305 35.630 191.475 ;
        RECT 35.815 191.330 36.085 192.235 ;
        RECT 35.460 191.160 35.630 191.305 ;
        RECT 33.015 190.665 34.245 190.835 ;
        RECT 34.895 190.755 35.225 191.125 ;
        RECT 35.460 190.830 35.745 191.160 ;
        RECT 32.995 189.855 33.505 190.390 ;
        RECT 33.725 190.060 33.970 190.665 ;
        RECT 35.460 190.575 35.630 190.830 ;
        RECT 34.965 190.405 35.630 190.575 ;
        RECT 35.915 190.530 36.085 191.330 ;
        RECT 36.265 191.795 36.595 192.225 ;
        RECT 36.775 191.965 36.970 192.405 ;
        RECT 37.140 191.795 37.470 192.225 ;
        RECT 36.265 191.625 37.470 191.795 ;
        RECT 36.265 191.295 37.160 191.625 ;
        RECT 37.640 191.455 37.915 192.225 ;
        RECT 38.185 191.660 38.455 192.405 ;
        RECT 39.085 192.400 45.360 192.405 ;
        RECT 38.625 191.490 38.915 192.230 ;
        RECT 39.085 191.675 39.340 192.400 ;
        RECT 39.525 191.505 39.785 192.230 ;
        RECT 39.955 191.675 40.200 192.400 ;
        RECT 40.385 191.505 40.645 192.230 ;
        RECT 40.815 191.675 41.060 192.400 ;
        RECT 41.245 191.505 41.505 192.230 ;
        RECT 41.675 191.675 41.920 192.400 ;
        RECT 42.090 191.505 42.350 192.230 ;
        RECT 42.520 191.675 42.780 192.400 ;
        RECT 42.950 191.505 43.210 192.230 ;
        RECT 43.380 191.675 43.640 192.400 ;
        RECT 43.810 191.505 44.070 192.230 ;
        RECT 44.240 191.675 44.500 192.400 ;
        RECT 44.670 191.505 44.930 192.230 ;
        RECT 45.100 191.605 45.360 192.400 ;
        RECT 39.525 191.490 44.930 191.505 ;
        RECT 37.330 191.265 37.915 191.455 ;
        RECT 38.185 191.265 44.930 191.490 ;
        RECT 36.270 190.765 36.565 191.095 ;
        RECT 36.745 190.765 37.160 191.095 ;
        RECT 34.965 190.025 35.135 190.405 ;
        RECT 35.315 189.855 35.645 190.235 ;
        RECT 35.825 190.025 36.085 190.530 ;
        RECT 36.265 189.855 36.565 190.585 ;
        RECT 36.745 190.145 36.975 190.765 ;
        RECT 37.330 190.595 37.505 191.265 ;
        RECT 37.175 190.415 37.505 190.595 ;
        RECT 37.675 190.445 37.915 191.095 ;
        RECT 38.185 190.675 39.350 191.265 ;
        RECT 45.530 191.095 45.780 192.230 ;
        RECT 45.960 191.595 46.220 192.405 ;
        RECT 46.395 191.095 46.640 192.235 ;
        RECT 46.820 191.595 47.115 192.405 ;
        RECT 47.300 191.535 47.565 192.235 ;
        RECT 47.735 191.705 48.065 192.405 ;
        RECT 48.235 191.535 48.905 192.235 ;
        RECT 49.410 191.705 49.840 192.405 ;
        RECT 50.020 191.845 50.210 192.235 ;
        RECT 50.380 192.025 50.710 192.405 ;
        RECT 51.065 192.065 52.225 192.235 ;
        RECT 50.020 191.675 50.750 191.845 ;
        RECT 47.300 191.280 49.875 191.535 ;
        RECT 39.520 190.845 46.640 191.095 ;
        RECT 38.185 190.505 44.930 190.675 ;
        RECT 37.175 190.035 37.400 190.415 ;
        RECT 37.570 189.855 37.900 190.245 ;
        RECT 38.185 189.855 38.485 190.335 ;
        RECT 38.655 190.050 38.915 190.505 ;
        RECT 39.085 189.855 39.345 190.335 ;
        RECT 39.525 190.050 39.785 190.505 ;
        RECT 39.955 189.855 40.205 190.335 ;
        RECT 40.385 190.050 40.645 190.505 ;
        RECT 40.815 189.855 41.065 190.335 ;
        RECT 41.245 190.050 41.505 190.505 ;
        RECT 41.675 189.855 41.920 190.335 ;
        RECT 42.090 190.050 42.365 190.505 ;
        RECT 42.535 189.855 42.780 190.335 ;
        RECT 42.950 190.050 43.210 190.505 ;
        RECT 43.380 189.855 43.640 190.335 ;
        RECT 43.810 190.050 44.070 190.505 ;
        RECT 44.240 189.855 44.500 190.335 ;
        RECT 44.670 190.050 44.930 190.505 ;
        RECT 45.100 189.855 45.360 190.415 ;
        RECT 45.530 190.035 45.780 190.845 ;
        RECT 45.960 189.855 46.220 190.380 ;
        RECT 46.390 190.035 46.640 190.845 ;
        RECT 46.810 190.535 47.125 191.095 ;
        RECT 47.295 190.765 47.570 191.095 ;
        RECT 47.740 190.595 47.920 191.280 ;
        RECT 49.705 191.095 49.875 191.280 ;
        RECT 48.090 190.765 48.450 191.095 ;
        RECT 48.740 191.045 49.030 191.095 ;
        RECT 48.735 190.875 49.030 191.045 ;
        RECT 48.740 190.765 49.030 190.875 ;
        RECT 49.200 190.765 49.535 191.095 ;
        RECT 49.705 190.765 50.385 191.095 ;
        RECT 46.820 189.855 47.125 190.365 ;
        RECT 47.305 190.195 47.920 190.595 ;
        RECT 48.090 190.405 49.360 190.595 ;
        RECT 50.555 190.555 50.750 191.675 ;
        RECT 51.065 191.565 51.235 192.065 ;
        RECT 51.495 191.435 51.665 191.895 ;
        RECT 51.895 191.815 52.225 192.065 ;
        RECT 52.450 191.985 52.780 192.405 ;
        RECT 53.035 191.815 53.320 192.235 ;
        RECT 51.895 191.645 53.320 191.815 ;
        RECT 53.565 191.605 53.895 192.405 ;
        RECT 54.145 191.685 54.480 192.195 ;
        RECT 51.040 191.095 51.245 191.385 ;
        RECT 51.495 191.265 53.865 191.435 ;
        RECT 53.695 191.095 53.865 191.265 ;
        RECT 51.040 191.045 51.390 191.095 ;
        RECT 51.035 190.875 51.390 191.045 ;
        RECT 51.040 190.765 51.390 190.875 ;
        RECT 49.930 190.385 50.750 190.555 ;
        RECT 47.305 190.025 47.640 190.195 ;
        RECT 48.600 189.855 48.935 190.235 ;
        RECT 49.525 189.855 49.760 190.295 ;
        RECT 49.930 190.025 50.260 190.385 ;
        RECT 50.430 189.855 50.760 190.215 ;
        RECT 50.985 189.855 51.315 190.575 ;
        RECT 51.700 190.430 52.120 191.095 ;
        RECT 52.290 190.705 52.580 191.095 ;
        RECT 52.770 191.045 53.040 191.095 ;
        RECT 53.250 191.045 53.500 191.095 ;
        RECT 52.770 190.875 53.045 191.045 ;
        RECT 53.250 190.875 53.505 191.045 ;
        RECT 52.290 190.535 52.585 190.705 ;
        RECT 52.290 190.435 52.580 190.535 ;
        RECT 52.770 190.435 53.040 190.875 ;
        RECT 53.250 190.765 53.500 190.875 ;
        RECT 53.695 190.765 54.000 191.095 ;
        RECT 53.695 190.595 53.865 190.765 ;
        RECT 53.305 190.425 53.865 190.595 ;
        RECT 53.305 190.255 53.475 190.425 ;
        RECT 54.225 190.330 54.480 191.685 ;
        RECT 54.655 191.240 54.945 192.405 ;
        RECT 55.170 191.535 55.455 192.405 ;
        RECT 55.625 191.775 55.885 192.235 ;
        RECT 56.060 191.945 56.315 192.405 ;
        RECT 56.485 191.775 56.745 192.235 ;
        RECT 55.625 191.605 56.745 191.775 ;
        RECT 56.915 191.605 57.225 192.405 ;
        RECT 55.625 191.355 55.885 191.605 ;
        RECT 57.395 191.435 57.705 192.235 ;
        RECT 57.875 191.985 58.215 192.405 ;
        RECT 58.385 191.815 58.635 192.235 ;
        RECT 55.130 191.185 55.885 191.355 ;
        RECT 56.675 191.265 57.705 191.435 ;
        RECT 55.130 190.675 55.535 191.185 ;
        RECT 56.675 191.015 56.845 191.265 ;
        RECT 55.705 190.845 56.845 191.015 ;
        RECT 51.860 190.085 53.475 190.255 ;
        RECT 53.645 189.855 53.975 190.255 ;
        RECT 54.145 190.070 54.480 190.330 ;
        RECT 54.655 189.855 54.945 190.580 ;
        RECT 55.130 190.505 56.780 190.675 ;
        RECT 57.015 190.525 57.365 191.095 ;
        RECT 55.175 189.855 55.455 190.335 ;
        RECT 55.625 190.115 55.885 190.505 ;
        RECT 56.060 189.855 56.315 190.335 ;
        RECT 56.485 190.115 56.780 190.505 ;
        RECT 57.535 190.355 57.705 191.265 ;
        RECT 57.875 191.645 58.635 191.815 ;
        RECT 57.875 190.675 58.185 191.645 ;
        RECT 58.805 191.565 59.135 192.405 ;
        RECT 59.625 191.815 60.380 192.235 ;
        RECT 59.305 191.645 60.770 191.815 ;
        RECT 59.305 191.395 59.475 191.645 ;
        RECT 58.515 191.225 59.475 191.395 ;
        RECT 58.515 191.055 58.685 191.225 ;
        RECT 59.645 191.055 59.950 191.475 ;
        RECT 58.355 190.845 58.685 191.055 ;
        RECT 58.855 190.845 59.295 191.055 ;
        RECT 59.465 190.845 59.950 191.055 ;
        RECT 60.140 191.045 60.430 191.475 ;
        RECT 60.600 191.440 60.770 191.645 ;
        RECT 60.940 191.620 61.180 192.405 ;
        RECT 61.350 191.440 61.680 192.235 ;
        RECT 62.025 191.595 62.320 192.405 ;
        RECT 60.600 191.265 61.680 191.440 ;
        RECT 60.600 191.215 61.385 191.265 ;
        RECT 60.140 190.845 60.530 191.045 ;
        RECT 60.700 190.845 61.045 191.045 ;
        RECT 57.875 190.505 58.635 190.675 ;
        RECT 56.960 189.855 57.235 190.335 ;
        RECT 57.405 190.025 57.705 190.355 ;
        RECT 57.965 189.855 58.135 190.335 ;
        RECT 58.305 190.035 58.635 190.505 ;
        RECT 58.805 189.855 58.975 190.675 ;
        RECT 59.145 190.505 60.845 190.675 ;
        RECT 59.145 190.040 59.475 190.505 ;
        RECT 60.460 190.415 60.845 190.505 ;
        RECT 61.215 190.575 61.385 191.215 ;
        RECT 62.500 191.095 62.745 192.235 ;
        RECT 62.920 191.595 63.180 192.405 ;
        RECT 63.780 192.400 70.055 192.405 ;
        RECT 63.360 191.095 63.610 192.230 ;
        RECT 63.780 191.605 64.040 192.400 ;
        RECT 64.210 191.505 64.470 192.230 ;
        RECT 64.640 191.675 64.900 192.400 ;
        RECT 65.070 191.505 65.330 192.230 ;
        RECT 65.500 191.675 65.760 192.400 ;
        RECT 65.930 191.505 66.190 192.230 ;
        RECT 66.360 191.675 66.620 192.400 ;
        RECT 66.790 191.505 67.050 192.230 ;
        RECT 67.220 191.675 67.465 192.400 ;
        RECT 67.635 191.505 67.895 192.230 ;
        RECT 68.080 191.675 68.325 192.400 ;
        RECT 68.495 191.505 68.755 192.230 ;
        RECT 68.940 191.675 69.185 192.400 ;
        RECT 69.355 191.505 69.615 192.230 ;
        RECT 69.800 191.675 70.055 192.400 ;
        RECT 64.210 191.490 69.615 191.505 ;
        RECT 70.225 191.490 70.515 192.230 ;
        RECT 70.685 191.660 70.955 192.405 ;
        RECT 71.305 191.660 71.575 192.405 ;
        RECT 72.205 192.400 78.480 192.405 ;
        RECT 71.745 191.490 72.035 192.230 ;
        RECT 72.205 191.675 72.460 192.400 ;
        RECT 72.645 191.505 72.905 192.230 ;
        RECT 73.075 191.675 73.320 192.400 ;
        RECT 73.505 191.505 73.765 192.230 ;
        RECT 73.935 191.675 74.180 192.400 ;
        RECT 74.365 191.505 74.625 192.230 ;
        RECT 74.795 191.675 75.040 192.400 ;
        RECT 75.210 191.505 75.470 192.230 ;
        RECT 75.640 191.675 75.900 192.400 ;
        RECT 76.070 191.505 76.330 192.230 ;
        RECT 76.500 191.675 76.760 192.400 ;
        RECT 76.930 191.505 77.190 192.230 ;
        RECT 77.360 191.675 77.620 192.400 ;
        RECT 77.790 191.505 78.050 192.230 ;
        RECT 78.220 191.605 78.480 192.400 ;
        RECT 72.645 191.490 78.050 191.505 ;
        RECT 64.210 191.265 70.955 191.490 ;
        RECT 61.585 190.745 61.845 191.095 ;
        RECT 61.215 190.405 61.760 190.575 ;
        RECT 62.015 190.535 62.330 191.095 ;
        RECT 62.500 190.845 69.620 191.095 ;
        RECT 69.790 191.045 70.955 191.265 ;
        RECT 71.305 191.265 78.050 191.490 ;
        RECT 69.790 190.875 70.985 191.045 ;
        RECT 59.645 189.855 59.815 190.325 ;
        RECT 60.075 190.065 61.260 190.235 ;
        RECT 61.430 190.025 61.760 190.405 ;
        RECT 62.015 189.855 62.320 190.365 ;
        RECT 62.500 190.035 62.750 190.845 ;
        RECT 62.920 189.855 63.180 190.380 ;
        RECT 63.360 190.035 63.610 190.845 ;
        RECT 69.790 190.675 70.955 190.875 ;
        RECT 64.210 190.505 70.955 190.675 ;
        RECT 71.305 190.675 72.470 191.265 ;
        RECT 78.650 191.095 78.900 192.230 ;
        RECT 79.080 191.595 79.340 192.405 ;
        RECT 79.515 191.095 79.760 192.235 ;
        RECT 79.940 191.595 80.235 192.405 ;
        RECT 80.415 191.240 80.705 192.405 ;
        RECT 80.935 191.705 81.155 192.235 ;
        RECT 81.325 191.895 81.655 192.405 ;
        RECT 81.825 191.705 82.050 192.235 ;
        RECT 80.935 191.440 82.050 191.705 ;
        RECT 82.220 191.690 82.535 192.235 ;
        RECT 82.725 191.990 83.055 192.405 ;
        RECT 82.220 191.460 83.055 191.690 ;
        RECT 72.640 190.845 79.760 191.095 ;
        RECT 71.305 190.505 78.050 190.675 ;
        RECT 63.780 189.855 64.040 190.415 ;
        RECT 64.210 190.050 64.470 190.505 ;
        RECT 64.640 189.855 64.900 190.335 ;
        RECT 65.070 190.050 65.330 190.505 ;
        RECT 65.500 189.855 65.760 190.335 ;
        RECT 65.930 190.050 66.190 190.505 ;
        RECT 66.360 189.855 66.605 190.335 ;
        RECT 66.775 190.050 67.050 190.505 ;
        RECT 67.220 189.855 67.465 190.335 ;
        RECT 67.635 190.050 67.895 190.505 ;
        RECT 68.075 189.855 68.325 190.335 ;
        RECT 68.495 190.050 68.755 190.505 ;
        RECT 68.935 189.855 69.185 190.335 ;
        RECT 69.355 190.050 69.615 190.505 ;
        RECT 69.795 189.855 70.055 190.335 ;
        RECT 70.225 190.050 70.485 190.505 ;
        RECT 70.655 189.855 70.955 190.335 ;
        RECT 71.305 189.855 71.605 190.335 ;
        RECT 71.775 190.050 72.035 190.505 ;
        RECT 72.205 189.855 72.465 190.335 ;
        RECT 72.645 190.050 72.905 190.505 ;
        RECT 73.075 189.855 73.325 190.335 ;
        RECT 73.505 190.050 73.765 190.505 ;
        RECT 73.935 189.855 74.185 190.335 ;
        RECT 74.365 190.050 74.625 190.505 ;
        RECT 74.795 189.855 75.040 190.335 ;
        RECT 75.210 190.050 75.485 190.505 ;
        RECT 75.655 189.855 75.900 190.335 ;
        RECT 76.070 190.050 76.330 190.505 ;
        RECT 76.500 189.855 76.760 190.335 ;
        RECT 76.930 190.050 77.190 190.505 ;
        RECT 77.360 189.855 77.620 190.335 ;
        RECT 77.790 190.050 78.050 190.505 ;
        RECT 78.220 189.855 78.480 190.415 ;
        RECT 78.650 190.035 78.900 190.845 ;
        RECT 79.080 189.855 79.340 190.380 ;
        RECT 79.510 190.035 79.760 190.845 ;
        RECT 79.930 190.535 80.245 191.095 ;
        RECT 79.940 189.855 80.245 190.365 ;
        RECT 80.415 189.855 80.705 190.580 ;
        RECT 80.885 190.520 81.200 191.095 ;
        RECT 80.875 189.855 81.205 190.335 ;
        RECT 81.390 190.135 81.770 191.095 ;
        RECT 82.220 190.765 82.545 191.180 ;
        RECT 82.715 190.765 83.055 191.460 ;
        RECT 82.715 190.595 82.885 190.765 ;
        RECT 83.225 190.595 83.455 192.235 ;
        RECT 83.625 191.435 83.915 192.405 ;
        RECT 84.100 191.605 84.355 192.405 ;
        RECT 84.555 191.555 84.885 192.235 ;
        RECT 84.100 191.065 84.345 191.425 ;
        RECT 84.535 191.275 84.885 191.555 ;
        RECT 84.535 190.895 84.705 191.275 ;
        RECT 85.065 191.095 85.260 192.145 ;
        RECT 85.440 191.265 85.760 192.405 ;
        RECT 85.935 191.315 87.145 192.405 ;
        RECT 82.145 190.425 82.885 190.595 ;
        RECT 82.145 190.025 82.335 190.425 ;
        RECT 83.055 190.405 83.455 190.595 ;
        RECT 84.185 190.725 84.705 190.895 ;
        RECT 84.875 190.765 85.260 191.095 ;
        RECT 85.440 191.045 85.700 191.095 ;
        RECT 85.440 190.875 85.705 191.045 ;
        RECT 85.440 190.765 85.700 190.875 ;
        RECT 85.935 190.775 86.455 191.315 ;
        RECT 82.555 189.855 82.885 190.215 ;
        RECT 83.055 190.025 83.245 190.405 ;
        RECT 83.415 189.855 83.745 190.235 ;
        RECT 84.185 190.160 84.355 190.725 ;
        RECT 86.625 190.605 87.145 191.145 ;
        RECT 84.545 190.385 85.760 190.555 ;
        RECT 84.545 190.080 84.775 190.385 ;
        RECT 84.945 189.855 85.275 190.215 ;
        RECT 85.470 190.035 85.760 190.385 ;
        RECT 85.935 189.855 87.145 190.605 ;
        RECT 15.930 189.685 87.230 189.855 ;
        RECT 16.015 188.935 17.225 189.685 ;
        RECT 16.015 188.395 16.535 188.935 ;
        RECT 17.400 188.845 17.660 189.685 ;
        RECT 17.835 188.940 18.090 189.515 ;
        RECT 18.260 189.305 18.590 189.685 ;
        RECT 18.805 189.135 18.975 189.515 ;
        RECT 18.260 188.965 18.975 189.135 ;
        RECT 16.705 188.225 17.225 188.765 ;
        RECT 16.015 187.135 17.225 188.225 ;
        RECT 17.400 187.135 17.660 188.285 ;
        RECT 17.835 188.210 18.005 188.940 ;
        RECT 18.260 188.775 18.430 188.965 ;
        RECT 19.235 188.885 19.545 189.685 ;
        RECT 19.750 188.885 20.445 189.515 ;
        RECT 20.615 188.945 21.105 189.515 ;
        RECT 21.275 189.115 21.505 189.515 ;
        RECT 21.675 189.285 22.095 189.685 ;
        RECT 22.265 189.115 22.435 189.515 ;
        RECT 21.275 188.945 22.435 189.115 ;
        RECT 22.605 188.945 23.055 189.685 ;
        RECT 23.225 188.945 23.665 189.505 ;
        RECT 19.750 188.835 19.925 188.885 ;
        RECT 18.175 188.445 18.430 188.775 ;
        RECT 18.260 188.235 18.430 188.445 ;
        RECT 18.710 188.415 19.065 188.785 ;
        RECT 19.245 188.445 19.580 188.715 ;
        RECT 19.750 188.285 19.920 188.835 ;
        RECT 20.090 188.445 20.425 188.695 ;
        RECT 17.835 187.305 18.090 188.210 ;
        RECT 18.260 188.065 18.975 188.235 ;
        RECT 18.260 187.135 18.590 187.895 ;
        RECT 18.805 187.305 18.975 188.065 ;
        RECT 19.235 187.135 19.515 188.275 ;
        RECT 19.685 187.305 20.015 188.285 ;
        RECT 20.615 188.275 20.785 188.945 ;
        RECT 20.955 188.445 21.360 188.775 ;
        RECT 20.185 187.135 20.445 188.275 ;
        RECT 20.615 188.105 21.385 188.275 ;
        RECT 20.625 187.135 20.955 187.935 ;
        RECT 21.135 187.475 21.385 188.105 ;
        RECT 21.575 187.645 21.825 188.775 ;
        RECT 22.025 188.445 22.270 188.775 ;
        RECT 22.455 188.495 22.845 188.775 ;
        RECT 22.025 187.645 22.225 188.445 ;
        RECT 23.015 188.325 23.185 188.775 ;
        RECT 22.395 188.155 23.185 188.325 ;
        RECT 22.395 187.475 22.565 188.155 ;
        RECT 21.135 187.305 22.565 187.475 ;
        RECT 22.735 187.135 23.050 187.985 ;
        RECT 23.355 187.935 23.665 188.945 ;
        RECT 23.225 187.305 23.665 187.935 ;
        RECT 24.755 188.945 25.095 189.515 ;
        RECT 25.290 189.020 25.460 189.685 ;
        RECT 25.740 189.345 25.960 189.390 ;
        RECT 25.735 189.175 25.960 189.345 ;
        RECT 26.130 189.205 26.575 189.375 ;
        RECT 25.740 189.035 25.960 189.175 ;
        RECT 24.755 187.975 24.930 188.945 ;
        RECT 25.740 188.865 26.235 189.035 ;
        RECT 25.100 188.325 25.270 188.775 ;
        RECT 25.440 188.495 25.890 188.695 ;
        RECT 26.060 188.670 26.235 188.865 ;
        RECT 26.405 188.415 26.575 189.205 ;
        RECT 26.745 189.080 26.995 189.450 ;
        RECT 26.825 188.695 26.995 189.080 ;
        RECT 27.165 189.045 27.415 189.450 ;
        RECT 27.585 189.215 27.755 189.685 ;
        RECT 27.925 189.045 28.265 189.450 ;
        RECT 27.165 188.865 28.265 189.045 ;
        RECT 28.455 188.875 28.695 189.685 ;
        RECT 28.865 188.875 29.195 189.515 ;
        RECT 29.365 188.875 29.635 189.685 ;
        RECT 26.825 188.525 27.020 188.695 ;
        RECT 25.100 188.155 25.495 188.325 ;
        RECT 26.405 188.275 26.680 188.415 ;
        RECT 24.755 187.305 25.015 187.975 ;
        RECT 25.325 187.885 25.495 188.155 ;
        RECT 25.665 188.055 26.680 188.275 ;
        RECT 26.850 188.275 27.020 188.525 ;
        RECT 27.190 188.445 27.750 188.695 ;
        RECT 26.850 187.885 27.405 188.275 ;
        RECT 25.325 187.715 27.405 187.885 ;
        RECT 25.185 187.135 25.515 187.535 ;
        RECT 26.385 187.135 26.785 187.535 ;
        RECT 27.075 187.480 27.405 187.715 ;
        RECT 27.575 187.345 27.750 188.445 ;
        RECT 27.920 188.125 28.265 188.695 ;
        RECT 28.435 188.445 28.785 188.695 ;
        RECT 28.955 188.275 29.125 188.875 ;
        RECT 29.855 188.865 30.085 189.685 ;
        RECT 30.255 188.885 30.585 189.515 ;
        RECT 29.295 188.445 29.645 188.695 ;
        RECT 29.835 188.445 30.165 188.695 ;
        RECT 30.335 188.285 30.585 188.885 ;
        RECT 30.755 188.865 30.965 189.685 ;
        RECT 31.200 188.945 31.455 189.515 ;
        RECT 31.625 189.285 31.955 189.685 ;
        RECT 32.380 189.150 32.910 189.515 ;
        RECT 32.380 189.115 32.555 189.150 ;
        RECT 31.625 188.945 32.555 189.115 ;
        RECT 33.100 189.005 33.375 189.515 ;
        RECT 28.445 188.105 29.125 188.275 ;
        RECT 27.920 187.135 28.265 187.955 ;
        RECT 28.445 187.320 28.775 188.105 ;
        RECT 29.305 187.135 29.635 188.275 ;
        RECT 29.855 187.135 30.085 188.275 ;
        RECT 30.255 187.305 30.585 188.285 ;
        RECT 31.200 188.275 31.370 188.945 ;
        RECT 31.625 188.775 31.795 188.945 ;
        RECT 31.540 188.445 31.795 188.775 ;
        RECT 32.020 188.445 32.215 188.775 ;
        RECT 30.755 187.135 30.965 188.275 ;
        RECT 31.200 187.305 31.535 188.275 ;
        RECT 31.705 187.135 31.875 188.275 ;
        RECT 32.045 187.475 32.215 188.445 ;
        RECT 32.385 187.815 32.555 188.945 ;
        RECT 32.725 188.155 32.895 188.955 ;
        RECT 33.095 188.835 33.375 189.005 ;
        RECT 33.100 188.355 33.375 188.835 ;
        RECT 33.545 188.155 33.735 189.515 ;
        RECT 33.915 189.150 34.425 189.685 ;
        RECT 34.645 188.875 34.890 189.480 ;
        RECT 35.340 188.945 35.595 189.515 ;
        RECT 35.765 189.285 36.095 189.685 ;
        RECT 36.520 189.150 37.050 189.515 ;
        RECT 36.520 189.115 36.695 189.150 ;
        RECT 35.765 188.945 36.695 189.115 ;
        RECT 33.935 188.705 35.165 188.875 ;
        RECT 32.725 187.985 33.735 188.155 ;
        RECT 33.905 188.140 34.655 188.330 ;
        RECT 32.385 187.645 33.510 187.815 ;
        RECT 33.905 187.475 34.075 188.140 ;
        RECT 34.825 187.895 35.165 188.705 ;
        RECT 32.045 187.305 34.075 187.475 ;
        RECT 34.245 187.135 34.415 187.895 ;
        RECT 34.650 187.485 35.165 187.895 ;
        RECT 35.340 188.275 35.510 188.945 ;
        RECT 35.765 188.775 35.935 188.945 ;
        RECT 35.680 188.445 35.935 188.775 ;
        RECT 36.160 188.445 36.355 188.775 ;
        RECT 35.340 187.305 35.675 188.275 ;
        RECT 35.845 187.135 36.015 188.275 ;
        RECT 36.185 187.475 36.355 188.445 ;
        RECT 36.525 187.815 36.695 188.945 ;
        RECT 36.865 188.155 37.035 188.955 ;
        RECT 37.240 188.665 37.515 189.515 ;
        RECT 37.235 188.495 37.515 188.665 ;
        RECT 37.240 188.355 37.515 188.495 ;
        RECT 37.685 188.155 37.875 189.515 ;
        RECT 38.055 189.150 38.565 189.685 ;
        RECT 38.785 188.875 39.030 189.480 ;
        RECT 40.025 189.135 40.195 189.515 ;
        RECT 40.410 189.305 40.740 189.685 ;
        RECT 40.025 188.965 40.740 189.135 ;
        RECT 38.075 188.705 39.305 188.875 ;
        RECT 36.865 187.985 37.875 188.155 ;
        RECT 38.045 188.140 38.795 188.330 ;
        RECT 36.525 187.645 37.650 187.815 ;
        RECT 38.045 187.475 38.215 188.140 ;
        RECT 38.965 187.895 39.305 188.705 ;
        RECT 39.935 188.415 40.290 188.785 ;
        RECT 40.570 188.775 40.740 188.965 ;
        RECT 40.910 188.940 41.165 189.515 ;
        RECT 40.570 188.445 40.825 188.775 ;
        RECT 40.570 188.235 40.740 188.445 ;
        RECT 36.185 187.305 38.215 187.475 ;
        RECT 38.385 187.135 38.555 187.895 ;
        RECT 38.790 187.485 39.305 187.895 ;
        RECT 40.025 188.065 40.740 188.235 ;
        RECT 40.995 188.210 41.165 188.940 ;
        RECT 41.340 188.845 41.600 189.685 ;
        RECT 41.775 188.960 42.065 189.685 ;
        RECT 42.285 188.885 42.495 189.685 ;
        RECT 40.025 187.305 40.195 188.065 ;
        RECT 40.410 187.135 40.740 187.895 ;
        RECT 40.910 187.305 41.165 188.210 ;
        RECT 41.340 187.135 41.600 188.285 ;
        RECT 41.775 187.135 42.065 188.300 ;
        RECT 42.285 187.135 42.495 188.275 ;
        RECT 42.665 187.305 43.005 189.515 ;
        RECT 43.185 189.225 43.435 189.685 ;
        RECT 43.625 189.055 43.955 189.515 ;
        RECT 44.155 189.345 44.540 189.515 ;
        RECT 44.135 189.175 44.540 189.345 ;
        RECT 43.180 188.885 43.955 189.055 ;
        RECT 43.180 187.985 43.455 188.885 ;
        RECT 43.655 188.155 43.985 188.695 ;
        RECT 44.155 188.155 44.540 189.175 ;
        RECT 45.015 189.145 45.345 189.515 ;
        RECT 45.535 189.315 45.865 189.685 ;
        RECT 46.035 189.145 46.365 189.515 ;
        RECT 45.015 188.945 46.365 189.145 ;
        RECT 46.835 188.885 47.530 189.515 ;
        RECT 47.735 188.885 48.045 189.685 ;
        RECT 48.300 189.135 48.630 189.515 ;
        RECT 48.800 189.305 49.985 189.475 ;
        RECT 50.245 189.215 50.415 189.685 ;
        RECT 48.300 188.965 48.845 189.135 ;
        RECT 44.830 188.155 45.250 188.695 ;
        RECT 45.450 188.445 45.810 188.775 ;
        RECT 45.980 188.455 46.665 188.765 ;
        RECT 43.180 187.745 45.345 187.985 ;
        RECT 43.185 187.135 43.805 187.575 ;
        RECT 44.010 187.305 44.290 187.745 ;
        RECT 44.475 187.135 44.805 187.515 ;
        RECT 45.015 187.305 45.345 187.745 ;
        RECT 45.520 187.645 45.810 188.445 ;
        RECT 45.515 187.475 45.810 187.645 ;
        RECT 45.520 187.400 45.810 187.475 ;
        RECT 46.035 187.135 46.290 188.275 ;
        RECT 46.460 187.415 46.665 188.455 ;
        RECT 46.855 188.445 47.190 188.695 ;
        RECT 47.360 188.285 47.530 188.885 ;
        RECT 47.700 188.445 48.035 188.715 ;
        RECT 48.215 188.445 48.475 188.795 ;
        RECT 48.675 188.325 48.845 188.965 ;
        RECT 49.215 189.035 49.600 189.125 ;
        RECT 50.585 189.035 50.915 189.500 ;
        RECT 49.215 188.865 50.915 189.035 ;
        RECT 51.085 188.865 51.255 189.685 ;
        RECT 51.425 189.035 51.755 189.505 ;
        RECT 51.925 189.205 52.095 189.685 ;
        RECT 52.365 189.345 53.555 189.515 ;
        RECT 52.365 189.175 52.675 189.345 ;
        RECT 51.425 188.865 52.185 189.035 ;
        RECT 49.015 188.495 49.360 188.695 ;
        RECT 49.530 188.495 49.920 188.695 ;
        RECT 46.835 187.135 47.095 188.275 ;
        RECT 47.265 187.305 47.595 188.285 ;
        RECT 48.675 188.275 49.460 188.325 ;
        RECT 47.765 187.135 48.045 188.275 ;
        RECT 48.380 188.100 49.460 188.275 ;
        RECT 48.380 187.305 48.710 188.100 ;
        RECT 48.880 187.135 49.120 187.920 ;
        RECT 49.290 187.895 49.460 188.100 ;
        RECT 49.630 188.065 49.920 188.495 ;
        RECT 50.110 188.485 50.595 188.695 ;
        RECT 50.765 188.485 51.205 188.695 ;
        RECT 51.375 188.485 51.705 188.695 ;
        RECT 50.110 188.065 50.415 188.485 ;
        RECT 51.375 188.315 51.545 188.485 ;
        RECT 50.585 188.145 51.545 188.315 ;
        RECT 50.585 187.895 50.755 188.145 ;
        RECT 49.290 187.725 50.755 187.895 ;
        RECT 49.680 187.305 50.435 187.725 ;
        RECT 50.925 187.135 51.255 187.975 ;
        RECT 51.875 187.895 52.185 188.865 ;
        RECT 52.360 188.370 52.675 189.005 ;
        RECT 51.425 187.725 52.185 187.895 ;
        RECT 51.425 187.305 51.675 187.725 ;
        RECT 51.845 187.135 52.185 187.555 ;
        RECT 52.365 187.135 52.675 188.200 ;
        RECT 52.845 187.985 53.055 189.175 ;
        RECT 53.225 189.055 53.555 189.345 ;
        RECT 53.795 189.225 53.965 189.685 ;
        RECT 54.195 189.055 54.525 189.515 ;
        RECT 54.705 189.225 54.875 189.685 ;
        RECT 55.055 189.055 55.385 189.515 ;
        RECT 55.635 189.205 55.915 189.685 ;
        RECT 53.225 188.885 55.385 189.055 ;
        RECT 56.085 189.035 56.345 189.425 ;
        RECT 56.520 189.205 56.775 189.685 ;
        RECT 56.945 189.035 57.240 189.425 ;
        RECT 57.420 189.205 57.695 189.685 ;
        RECT 57.865 189.185 58.165 189.515 ;
        RECT 58.425 189.205 58.725 189.685 ;
        RECT 55.590 188.865 57.240 189.035 ;
        RECT 53.395 188.325 53.890 188.695 ;
        RECT 54.070 188.495 54.870 188.695 ;
        RECT 55.040 188.325 55.370 188.715 ;
        RECT 53.335 188.155 55.370 188.325 ;
        RECT 55.590 188.355 55.995 188.865 ;
        RECT 56.165 188.525 57.305 188.695 ;
        RECT 55.590 188.185 56.345 188.355 ;
        RECT 52.845 187.805 54.495 187.985 ;
        RECT 52.845 187.305 53.080 187.805 ;
        RECT 54.195 187.645 54.495 187.805 ;
        RECT 53.250 187.135 53.580 187.595 ;
        RECT 53.775 187.475 53.965 187.635 ;
        RECT 54.665 187.475 54.885 187.985 ;
        RECT 53.775 187.305 54.885 187.475 ;
        RECT 55.055 187.135 55.385 187.985 ;
        RECT 55.630 187.135 55.915 188.005 ;
        RECT 56.085 187.935 56.345 188.185 ;
        RECT 57.135 188.275 57.305 188.525 ;
        RECT 57.475 188.445 57.825 189.015 ;
        RECT 57.995 188.275 58.165 189.185 ;
        RECT 58.895 189.035 59.155 189.490 ;
        RECT 59.325 189.205 59.585 189.685 ;
        RECT 59.765 189.035 60.025 189.490 ;
        RECT 60.195 189.205 60.445 189.685 ;
        RECT 60.625 189.035 60.885 189.490 ;
        RECT 61.055 189.205 61.305 189.685 ;
        RECT 61.485 189.035 61.745 189.490 ;
        RECT 61.915 189.205 62.160 189.685 ;
        RECT 62.330 189.035 62.605 189.490 ;
        RECT 62.775 189.205 63.020 189.685 ;
        RECT 63.190 189.035 63.450 189.490 ;
        RECT 63.620 189.205 63.880 189.685 ;
        RECT 64.050 189.035 64.310 189.490 ;
        RECT 64.480 189.205 64.740 189.685 ;
        RECT 64.910 189.035 65.170 189.490 ;
        RECT 65.340 189.125 65.600 189.685 ;
        RECT 57.135 188.105 58.165 188.275 ;
        RECT 56.085 187.765 57.205 187.935 ;
        RECT 56.085 187.305 56.345 187.765 ;
        RECT 56.520 187.135 56.775 187.595 ;
        RECT 56.945 187.305 57.205 187.765 ;
        RECT 57.375 187.135 57.685 187.935 ;
        RECT 57.855 187.305 58.165 188.105 ;
        RECT 58.425 188.865 65.170 189.035 ;
        RECT 58.425 188.275 59.590 188.865 ;
        RECT 65.770 188.695 66.020 189.505 ;
        RECT 66.200 189.160 66.460 189.685 ;
        RECT 66.630 188.695 66.880 189.505 ;
        RECT 67.060 189.175 67.365 189.685 ;
        RECT 59.760 188.445 66.880 188.695 ;
        RECT 67.050 188.445 67.365 189.005 ;
        RECT 67.535 188.960 67.825 189.685 ;
        RECT 68.020 188.860 68.275 189.685 ;
        RECT 68.445 188.945 68.780 189.515 ;
        RECT 68.975 189.020 69.145 189.685 ;
        RECT 69.425 189.035 69.645 189.390 ;
        RECT 69.815 189.205 70.275 189.375 ;
        RECT 69.425 189.000 69.930 189.035 ;
        RECT 58.425 188.050 65.170 188.275 ;
        RECT 58.425 187.135 58.695 187.880 ;
        RECT 58.865 187.310 59.155 188.050 ;
        RECT 59.765 188.035 65.170 188.050 ;
        RECT 59.325 187.140 59.580 187.865 ;
        RECT 59.765 187.310 60.025 188.035 ;
        RECT 60.195 187.140 60.440 187.865 ;
        RECT 60.625 187.310 60.885 188.035 ;
        RECT 61.055 187.140 61.300 187.865 ;
        RECT 61.485 187.310 61.745 188.035 ;
        RECT 61.915 187.140 62.160 187.865 ;
        RECT 62.330 187.310 62.590 188.035 ;
        RECT 62.760 187.140 63.020 187.865 ;
        RECT 63.190 187.310 63.450 188.035 ;
        RECT 63.620 187.140 63.880 187.865 ;
        RECT 64.050 187.310 64.310 188.035 ;
        RECT 64.480 187.140 64.740 187.865 ;
        RECT 64.910 187.310 65.170 188.035 ;
        RECT 65.340 187.140 65.600 187.935 ;
        RECT 65.770 187.310 66.020 188.445 ;
        RECT 59.325 187.135 65.600 187.140 ;
        RECT 66.200 187.135 66.460 187.945 ;
        RECT 66.635 187.305 66.880 188.445 ;
        RECT 67.060 187.135 67.355 187.945 ;
        RECT 67.535 187.135 67.825 188.300 ;
        RECT 68.020 187.135 68.275 188.360 ;
        RECT 68.445 187.985 68.615 188.945 ;
        RECT 69.425 188.865 69.935 189.000 ;
        RECT 68.785 188.325 68.955 188.775 ;
        RECT 69.125 188.495 69.595 188.695 ;
        RECT 69.765 188.670 69.935 188.865 ;
        RECT 70.105 188.415 70.275 189.205 ;
        RECT 70.445 189.080 70.690 189.450 ;
        RECT 70.520 188.695 70.690 189.080 ;
        RECT 70.865 189.045 71.095 189.450 ;
        RECT 71.285 189.215 71.455 189.685 ;
        RECT 71.625 189.045 71.955 189.450 ;
        RECT 70.865 188.865 71.955 189.045 ;
        RECT 72.135 188.885 72.425 189.685 ;
        RECT 72.595 189.225 73.145 189.515 ;
        RECT 73.315 189.225 73.565 189.685 ;
        RECT 70.520 188.525 70.710 188.695 ;
        RECT 68.785 188.155 69.180 188.325 ;
        RECT 70.105 188.275 70.370 188.415 ;
        RECT 68.445 187.975 68.685 187.985 ;
        RECT 68.445 187.305 68.700 187.975 ;
        RECT 69.010 187.885 69.180 188.155 ;
        RECT 69.350 188.055 70.370 188.275 ;
        RECT 70.540 188.275 70.710 188.525 ;
        RECT 70.880 188.445 71.435 188.695 ;
        RECT 70.540 187.885 71.095 188.275 ;
        RECT 69.010 187.715 71.095 187.885 ;
        RECT 68.870 187.135 69.200 187.535 ;
        RECT 70.070 187.135 70.475 187.535 ;
        RECT 70.745 187.345 71.095 187.715 ;
        RECT 71.265 187.645 71.435 188.445 ;
        RECT 71.610 188.125 71.955 188.695 ;
        RECT 71.265 187.475 71.445 187.645 ;
        RECT 71.265 187.345 71.435 187.475 ;
        RECT 71.640 187.135 71.955 187.955 ;
        RECT 72.135 187.135 72.425 188.275 ;
        RECT 72.595 187.855 72.845 189.225 ;
        RECT 74.195 189.055 74.525 189.415 ;
        RECT 74.985 189.205 75.285 189.685 ;
        RECT 73.135 188.865 74.525 189.055 ;
        RECT 75.455 189.035 75.715 189.490 ;
        RECT 75.885 189.205 76.145 189.685 ;
        RECT 76.325 189.035 76.585 189.490 ;
        RECT 76.755 189.205 77.005 189.685 ;
        RECT 77.185 189.035 77.445 189.490 ;
        RECT 77.615 189.205 77.865 189.685 ;
        RECT 78.045 189.035 78.305 189.490 ;
        RECT 78.475 189.205 78.720 189.685 ;
        RECT 78.890 189.035 79.165 189.490 ;
        RECT 79.335 189.205 79.580 189.685 ;
        RECT 79.750 189.035 80.010 189.490 ;
        RECT 80.180 189.205 80.440 189.685 ;
        RECT 80.610 189.035 80.870 189.490 ;
        RECT 81.040 189.205 81.300 189.685 ;
        RECT 81.470 189.035 81.730 189.490 ;
        RECT 81.900 189.125 82.160 189.685 ;
        RECT 74.985 188.865 81.730 189.035 ;
        RECT 73.135 188.775 73.305 188.865 ;
        RECT 73.015 188.445 73.305 188.775 ;
        RECT 73.475 188.445 73.805 188.695 ;
        RECT 74.035 188.445 74.725 188.695 ;
        RECT 73.135 188.195 73.305 188.445 ;
        RECT 73.135 188.025 74.075 188.195 ;
        RECT 72.595 187.305 73.045 187.855 ;
        RECT 73.235 187.135 73.565 187.855 ;
        RECT 73.775 187.475 74.075 188.025 ;
        RECT 74.410 188.005 74.725 188.445 ;
        RECT 74.985 188.275 76.150 188.865 ;
        RECT 82.330 188.695 82.580 189.505 ;
        RECT 82.760 189.160 83.020 189.685 ;
        RECT 83.190 188.695 83.440 189.505 ;
        RECT 83.620 189.175 83.925 189.685 ;
        RECT 84.100 189.285 84.435 189.685 ;
        RECT 84.605 189.115 84.810 189.515 ;
        RECT 85.020 189.205 85.295 189.685 ;
        RECT 85.505 189.185 85.765 189.515 ;
        RECT 76.320 188.445 83.440 188.695 ;
        RECT 83.610 188.445 83.925 189.005 ;
        RECT 84.125 188.945 84.810 189.115 ;
        RECT 74.985 188.050 81.730 188.275 ;
        RECT 74.245 187.135 74.525 187.805 ;
        RECT 74.985 187.135 75.255 187.880 ;
        RECT 75.425 187.310 75.715 188.050 ;
        RECT 76.325 188.035 81.730 188.050 ;
        RECT 75.885 187.140 76.140 187.865 ;
        RECT 76.325 187.310 76.585 188.035 ;
        RECT 76.755 187.140 77.000 187.865 ;
        RECT 77.185 187.310 77.445 188.035 ;
        RECT 77.615 187.140 77.860 187.865 ;
        RECT 78.045 187.310 78.305 188.035 ;
        RECT 78.475 187.140 78.720 187.865 ;
        RECT 78.890 187.310 79.150 188.035 ;
        RECT 79.320 187.140 79.580 187.865 ;
        RECT 79.750 187.310 80.010 188.035 ;
        RECT 80.180 187.140 80.440 187.865 ;
        RECT 80.610 187.310 80.870 188.035 ;
        RECT 81.040 187.140 81.300 187.865 ;
        RECT 81.470 187.310 81.730 188.035 ;
        RECT 81.900 187.140 82.160 187.935 ;
        RECT 82.330 187.310 82.580 188.445 ;
        RECT 75.885 187.135 82.160 187.140 ;
        RECT 82.760 187.135 83.020 187.945 ;
        RECT 83.195 187.305 83.440 188.445 ;
        RECT 83.620 187.135 83.915 187.945 ;
        RECT 84.125 187.915 84.465 188.945 ;
        RECT 84.635 188.275 84.885 188.775 ;
        RECT 85.065 188.445 85.425 189.025 ;
        RECT 85.595 188.275 85.765 189.185 ;
        RECT 85.935 188.935 87.145 189.685 ;
        RECT 84.635 188.105 85.765 188.275 ;
        RECT 84.125 187.740 84.790 187.915 ;
        RECT 84.100 187.135 84.435 187.560 ;
        RECT 84.605 187.335 84.790 187.740 ;
        RECT 84.995 187.135 85.325 187.915 ;
        RECT 85.495 187.335 85.765 188.105 ;
        RECT 85.935 188.225 86.455 188.765 ;
        RECT 86.625 188.395 87.145 188.935 ;
        RECT 85.935 187.135 87.145 188.225 ;
        RECT 15.930 186.965 87.230 187.135 ;
        RECT 16.015 185.875 17.225 186.965 ;
        RECT 16.015 185.165 16.535 185.705 ;
        RECT 16.705 185.335 17.225 185.875 ;
        RECT 17.475 186.035 17.655 186.795 ;
        RECT 17.835 186.205 18.165 186.965 ;
        RECT 17.475 185.865 18.150 186.035 ;
        RECT 18.335 185.890 18.605 186.795 ;
        RECT 17.980 185.720 18.150 185.865 ;
        RECT 17.415 185.315 17.755 185.685 ;
        RECT 17.980 185.390 18.255 185.720 ;
        RECT 16.015 184.415 17.225 185.165 ;
        RECT 17.980 185.135 18.150 185.390 ;
        RECT 17.485 184.965 18.150 185.135 ;
        RECT 18.425 185.090 18.605 185.890 ;
        RECT 19.235 185.825 19.515 186.965 ;
        RECT 19.685 185.815 20.015 186.795 ;
        RECT 20.185 185.825 20.445 186.965 ;
        RECT 20.625 186.165 20.955 186.965 ;
        RECT 21.135 186.625 22.565 186.795 ;
        RECT 21.135 185.995 21.385 186.625 ;
        RECT 20.615 185.825 21.385 185.995 ;
        RECT 19.750 185.775 19.925 185.815 ;
        RECT 19.245 185.385 19.580 185.655 ;
        RECT 19.750 185.215 19.920 185.775 ;
        RECT 20.090 185.405 20.425 185.655 ;
        RECT 17.485 184.585 17.655 184.965 ;
        RECT 17.835 184.415 18.165 184.795 ;
        RECT 18.345 184.585 18.605 185.090 ;
        RECT 19.235 184.415 19.545 185.215 ;
        RECT 19.750 184.585 20.445 185.215 ;
        RECT 20.615 185.155 20.785 185.825 ;
        RECT 20.955 185.325 21.360 185.655 ;
        RECT 21.575 185.325 21.825 186.455 ;
        RECT 22.025 185.655 22.225 186.455 ;
        RECT 22.395 185.945 22.565 186.625 ;
        RECT 22.735 186.115 23.050 186.965 ;
        RECT 23.225 186.165 23.665 186.795 ;
        RECT 22.395 185.775 23.185 185.945 ;
        RECT 22.025 185.325 22.270 185.655 ;
        RECT 22.455 185.325 22.845 185.605 ;
        RECT 23.015 185.325 23.185 185.775 ;
        RECT 23.355 185.155 23.665 186.165 ;
        RECT 20.615 184.585 21.105 185.155 ;
        RECT 21.275 184.985 22.435 185.155 ;
        RECT 21.275 184.585 21.505 184.985 ;
        RECT 21.675 184.415 22.095 184.815 ;
        RECT 22.265 184.585 22.435 184.985 ;
        RECT 22.605 184.415 23.055 185.155 ;
        RECT 23.225 184.595 23.665 185.155 ;
        RECT 24.295 186.125 24.555 186.795 ;
        RECT 24.725 186.565 25.055 186.965 ;
        RECT 25.925 186.565 26.325 186.965 ;
        RECT 26.615 186.385 26.945 186.620 ;
        RECT 24.865 186.215 26.945 186.385 ;
        RECT 24.295 186.115 24.525 186.125 ;
        RECT 24.295 185.155 24.470 186.115 ;
        RECT 24.865 185.945 25.035 186.215 ;
        RECT 24.640 185.775 25.035 185.945 ;
        RECT 25.205 185.825 26.220 186.045 ;
        RECT 24.640 185.325 24.810 185.775 ;
        RECT 25.945 185.685 26.220 185.825 ;
        RECT 26.390 185.825 26.945 186.215 ;
        RECT 24.980 185.405 25.430 185.605 ;
        RECT 25.600 185.235 25.775 185.430 ;
        RECT 24.295 184.585 24.635 185.155 ;
        RECT 24.830 184.415 25.000 185.080 ;
        RECT 25.280 185.065 25.775 185.235 ;
        RECT 25.280 184.925 25.500 185.065 ;
        RECT 25.275 184.755 25.500 184.925 ;
        RECT 25.945 184.895 26.115 185.685 ;
        RECT 26.390 185.575 26.560 185.825 ;
        RECT 27.115 185.655 27.290 186.755 ;
        RECT 27.460 186.145 27.805 186.965 ;
        RECT 26.365 185.405 26.560 185.575 ;
        RECT 26.730 185.405 27.290 185.655 ;
        RECT 27.460 185.405 27.805 185.975 ;
        RECT 28.895 185.800 29.185 186.965 ;
        RECT 29.355 185.890 29.625 186.795 ;
        RECT 29.795 186.205 30.125 186.965 ;
        RECT 30.305 186.035 30.485 186.795 ;
        RECT 26.365 185.020 26.535 185.405 ;
        RECT 25.280 184.710 25.500 184.755 ;
        RECT 25.670 184.725 26.115 184.895 ;
        RECT 26.285 184.650 26.535 185.020 ;
        RECT 26.705 185.055 27.805 185.235 ;
        RECT 26.705 184.650 26.955 185.055 ;
        RECT 27.125 184.415 27.295 184.885 ;
        RECT 27.465 184.650 27.805 185.055 ;
        RECT 28.895 184.415 29.185 185.140 ;
        RECT 29.355 185.090 29.535 185.890 ;
        RECT 29.810 185.865 30.485 186.035 ;
        RECT 29.810 185.720 29.980 185.865 ;
        RECT 29.705 185.390 29.980 185.720 ;
        RECT 30.740 185.825 31.075 186.795 ;
        RECT 31.245 185.825 31.415 186.965 ;
        RECT 31.585 186.625 33.615 186.795 ;
        RECT 29.810 185.135 29.980 185.390 ;
        RECT 30.205 185.315 30.545 185.685 ;
        RECT 30.740 185.155 30.910 185.825 ;
        RECT 31.585 185.655 31.755 186.625 ;
        RECT 31.080 185.325 31.335 185.655 ;
        RECT 31.560 185.325 31.755 185.655 ;
        RECT 31.925 186.285 33.050 186.455 ;
        RECT 31.165 185.155 31.335 185.325 ;
        RECT 31.925 185.155 32.095 186.285 ;
        RECT 29.355 184.585 29.615 185.090 ;
        RECT 29.810 184.965 30.475 185.135 ;
        RECT 29.795 184.415 30.125 184.795 ;
        RECT 30.305 184.585 30.475 184.965 ;
        RECT 30.740 184.585 30.995 185.155 ;
        RECT 31.165 184.985 32.095 185.155 ;
        RECT 32.265 185.945 33.275 186.115 ;
        RECT 32.265 185.145 32.435 185.945 ;
        RECT 32.640 185.265 32.915 185.745 ;
        RECT 32.635 185.095 32.915 185.265 ;
        RECT 31.920 184.950 32.095 184.985 ;
        RECT 31.165 184.415 31.495 184.815 ;
        RECT 31.920 184.585 32.450 184.950 ;
        RECT 32.640 184.585 32.915 185.095 ;
        RECT 33.085 184.585 33.275 185.945 ;
        RECT 33.445 185.960 33.615 186.625 ;
        RECT 33.785 186.205 33.955 186.965 ;
        RECT 34.190 186.205 34.705 186.615 ;
        RECT 33.445 185.770 34.195 185.960 ;
        RECT 34.365 185.395 34.705 186.205 ;
        RECT 34.965 186.035 35.135 186.795 ;
        RECT 35.315 186.205 35.645 186.965 ;
        RECT 34.965 185.865 35.630 186.035 ;
        RECT 35.815 185.890 36.085 186.795 ;
        RECT 35.460 185.720 35.630 185.865 ;
        RECT 33.475 185.225 34.705 185.395 ;
        RECT 34.895 185.315 35.225 185.685 ;
        RECT 35.460 185.390 35.745 185.720 ;
        RECT 33.455 184.415 33.965 184.950 ;
        RECT 34.185 184.620 34.430 185.225 ;
        RECT 35.460 185.135 35.630 185.390 ;
        RECT 34.965 184.965 35.630 185.135 ;
        RECT 35.915 185.090 36.085 185.890 ;
        RECT 34.965 184.585 35.135 184.965 ;
        RECT 35.315 184.415 35.645 184.795 ;
        RECT 35.825 184.585 36.085 185.090 ;
        RECT 36.715 185.890 36.985 186.795 ;
        RECT 37.155 186.205 37.485 186.965 ;
        RECT 37.665 186.035 37.845 186.795 ;
        RECT 36.715 185.090 36.895 185.890 ;
        RECT 37.170 185.865 37.845 186.035 ;
        RECT 39.035 186.075 39.295 186.785 ;
        RECT 39.465 186.255 39.795 186.965 ;
        RECT 39.965 186.075 40.195 186.785 ;
        RECT 37.170 185.720 37.340 185.865 ;
        RECT 39.035 185.835 40.195 186.075 ;
        RECT 40.375 186.055 40.645 186.785 ;
        RECT 40.825 186.235 41.165 186.965 ;
        RECT 40.375 185.835 41.145 186.055 ;
        RECT 37.065 185.390 37.340 185.720 ;
        RECT 37.170 185.135 37.340 185.390 ;
        RECT 37.565 185.315 37.905 185.685 ;
        RECT 39.025 185.325 39.325 185.655 ;
        RECT 39.505 185.345 40.030 185.655 ;
        RECT 40.210 185.345 40.675 185.655 ;
        RECT 36.715 184.585 36.975 185.090 ;
        RECT 37.170 184.965 37.835 185.135 ;
        RECT 37.155 184.415 37.485 184.795 ;
        RECT 37.665 184.585 37.835 184.965 ;
        RECT 39.035 184.415 39.325 185.145 ;
        RECT 39.505 184.705 39.735 185.345 ;
        RECT 40.855 185.165 41.145 185.835 ;
        RECT 39.915 184.965 41.145 185.165 ;
        RECT 39.915 184.595 40.225 184.965 ;
        RECT 40.405 184.415 41.075 184.785 ;
        RECT 41.335 184.595 41.595 186.785 ;
        RECT 42.235 186.545 42.575 186.965 ;
        RECT 42.745 186.375 42.995 186.795 ;
        RECT 42.235 186.205 42.995 186.375 ;
        RECT 42.235 185.235 42.545 186.205 ;
        RECT 43.165 186.125 43.495 186.965 ;
        RECT 43.985 186.375 44.740 186.795 ;
        RECT 43.665 186.205 45.130 186.375 ;
        RECT 43.665 185.955 43.835 186.205 ;
        RECT 42.875 185.785 43.835 185.955 ;
        RECT 42.875 185.615 43.045 185.785 ;
        RECT 44.005 185.615 44.310 186.035 ;
        RECT 42.715 185.405 43.045 185.615 ;
        RECT 43.215 185.405 43.655 185.615 ;
        RECT 43.825 185.405 44.310 185.615 ;
        RECT 44.500 185.605 44.790 186.035 ;
        RECT 44.960 186.000 45.130 186.205 ;
        RECT 45.300 186.180 45.540 186.965 ;
        RECT 45.710 186.000 46.040 186.795 ;
        RECT 44.960 185.825 46.040 186.000 ;
        RECT 44.960 185.775 45.745 185.825 ;
        RECT 44.500 185.405 44.890 185.605 ;
        RECT 45.060 185.405 45.405 185.605 ;
        RECT 42.235 185.065 42.995 185.235 ;
        RECT 42.325 184.415 42.495 184.895 ;
        RECT 42.665 184.595 42.995 185.065 ;
        RECT 43.165 184.415 43.335 185.235 ;
        RECT 43.505 185.065 45.205 185.235 ;
        RECT 43.505 184.600 43.835 185.065 ;
        RECT 44.820 184.975 45.205 185.065 ;
        RECT 45.575 185.135 45.745 185.775 ;
        RECT 45.945 185.305 46.205 185.655 ;
        RECT 45.575 184.965 46.120 185.135 ;
        RECT 44.005 184.415 44.175 184.885 ;
        RECT 44.435 184.625 45.620 184.795 ;
        RECT 45.790 184.585 46.120 184.965 ;
        RECT 47.295 184.695 47.575 186.795 ;
        RECT 47.765 186.205 48.550 186.965 ;
        RECT 48.945 186.135 49.330 186.795 ;
        RECT 48.945 186.035 49.355 186.135 ;
        RECT 47.745 185.825 49.355 186.035 ;
        RECT 49.655 185.945 49.855 186.735 ;
        RECT 47.745 185.225 48.020 185.825 ;
        RECT 49.525 185.775 49.855 185.945 ;
        RECT 50.025 185.785 50.345 186.965 ;
        RECT 50.525 186.355 50.855 186.785 ;
        RECT 51.035 186.525 51.230 186.965 ;
        RECT 51.400 186.355 51.730 186.785 ;
        RECT 50.525 186.185 51.730 186.355 ;
        RECT 50.525 185.855 51.420 186.185 ;
        RECT 51.900 186.015 52.175 186.785 ;
        RECT 52.460 186.165 52.715 186.965 ;
        RECT 51.590 185.825 52.175 186.015 ;
        RECT 52.885 185.995 53.215 186.795 ;
        RECT 53.385 186.165 53.555 186.965 ;
        RECT 53.725 185.995 54.055 186.795 ;
        RECT 52.355 185.825 54.055 185.995 ;
        RECT 54.225 185.825 54.485 186.965 ;
        RECT 49.525 185.655 49.705 185.775 ;
        RECT 48.190 185.405 48.545 185.655 ;
        RECT 48.740 185.605 49.205 185.655 ;
        RECT 48.735 185.435 49.205 185.605 ;
        RECT 48.740 185.405 49.205 185.435 ;
        RECT 49.375 185.405 49.705 185.655 ;
        RECT 49.880 185.405 50.345 185.605 ;
        RECT 50.530 185.325 50.825 185.655 ;
        RECT 51.005 185.325 51.420 185.655 ;
        RECT 47.745 185.045 48.995 185.225 ;
        RECT 48.630 184.975 48.995 185.045 ;
        RECT 49.165 185.025 50.345 185.195 ;
        RECT 47.805 184.415 47.975 184.875 ;
        RECT 49.165 184.805 49.495 185.025 ;
        RECT 48.245 184.625 49.495 184.805 ;
        RECT 49.665 184.415 49.835 184.855 ;
        RECT 50.005 184.610 50.345 185.025 ;
        RECT 50.525 184.415 50.825 185.145 ;
        RECT 51.005 184.705 51.235 185.325 ;
        RECT 51.590 185.155 51.765 185.825 ;
        RECT 51.435 184.975 51.765 185.155 ;
        RECT 51.935 185.005 52.175 185.655 ;
        RECT 52.355 185.235 52.635 185.825 ;
        RECT 54.655 185.800 54.945 186.965 ;
        RECT 55.205 186.220 55.475 186.965 ;
        RECT 56.105 186.960 62.380 186.965 ;
        RECT 55.645 186.050 55.935 186.790 ;
        RECT 56.105 186.235 56.360 186.960 ;
        RECT 56.545 186.065 56.805 186.790 ;
        RECT 56.975 186.235 57.220 186.960 ;
        RECT 57.405 186.065 57.665 186.790 ;
        RECT 57.835 186.235 58.080 186.960 ;
        RECT 58.265 186.065 58.525 186.790 ;
        RECT 58.695 186.235 58.940 186.960 ;
        RECT 59.110 186.065 59.370 186.790 ;
        RECT 59.540 186.235 59.800 186.960 ;
        RECT 59.970 186.065 60.230 186.790 ;
        RECT 60.400 186.235 60.660 186.960 ;
        RECT 60.830 186.065 61.090 186.790 ;
        RECT 61.260 186.235 61.520 186.960 ;
        RECT 61.690 186.065 61.950 186.790 ;
        RECT 62.120 186.165 62.380 186.960 ;
        RECT 56.545 186.050 61.950 186.065 ;
        RECT 55.205 185.825 61.950 186.050 ;
        RECT 52.805 185.405 53.555 185.655 ;
        RECT 53.725 185.405 54.485 185.655 ;
        RECT 55.205 185.235 56.370 185.825 ;
        RECT 62.550 185.655 62.800 186.790 ;
        RECT 62.980 186.155 63.240 186.965 ;
        RECT 63.415 185.655 63.660 186.795 ;
        RECT 63.840 186.155 64.135 186.965 ;
        RECT 64.370 186.095 64.655 186.965 ;
        RECT 64.825 186.335 65.085 186.795 ;
        RECT 65.260 186.505 65.515 186.965 ;
        RECT 65.685 186.335 65.945 186.795 ;
        RECT 64.825 186.165 65.945 186.335 ;
        RECT 66.115 186.165 66.425 186.965 ;
        RECT 64.825 185.915 65.085 186.165 ;
        RECT 66.595 185.995 66.905 186.795 ;
        RECT 67.085 186.155 67.380 186.965 ;
        RECT 64.330 185.745 65.085 185.915 ;
        RECT 65.875 185.825 66.905 185.995 ;
        RECT 56.540 185.405 63.660 185.655 ;
        RECT 52.355 184.985 53.215 185.235 ;
        RECT 53.385 185.045 54.485 185.215 ;
        RECT 51.435 184.595 51.660 184.975 ;
        RECT 51.830 184.415 52.160 184.805 ;
        RECT 52.465 184.795 52.795 184.815 ;
        RECT 53.385 184.795 53.635 185.045 ;
        RECT 52.465 184.585 53.635 184.795 ;
        RECT 53.805 184.415 53.975 184.875 ;
        RECT 54.145 184.585 54.485 185.045 ;
        RECT 54.655 184.415 54.945 185.140 ;
        RECT 55.205 185.065 61.950 185.235 ;
        RECT 55.205 184.415 55.505 184.895 ;
        RECT 55.675 184.610 55.935 185.065 ;
        RECT 56.105 184.415 56.365 184.895 ;
        RECT 56.545 184.610 56.805 185.065 ;
        RECT 56.975 184.415 57.225 184.895 ;
        RECT 57.405 184.610 57.665 185.065 ;
        RECT 57.835 184.415 58.085 184.895 ;
        RECT 58.265 184.610 58.525 185.065 ;
        RECT 58.695 184.415 58.940 184.895 ;
        RECT 59.110 184.610 59.385 185.065 ;
        RECT 59.555 184.415 59.800 184.895 ;
        RECT 59.970 184.610 60.230 185.065 ;
        RECT 60.400 184.415 60.660 184.895 ;
        RECT 60.830 184.610 61.090 185.065 ;
        RECT 61.260 184.415 61.520 184.895 ;
        RECT 61.690 184.610 61.950 185.065 ;
        RECT 62.120 184.415 62.380 184.975 ;
        RECT 62.550 184.595 62.800 185.405 ;
        RECT 62.980 184.415 63.240 184.940 ;
        RECT 63.410 184.595 63.660 185.405 ;
        RECT 63.830 185.095 64.145 185.655 ;
        RECT 64.330 185.235 64.735 185.745 ;
        RECT 65.875 185.575 66.045 185.825 ;
        RECT 64.905 185.405 66.045 185.575 ;
        RECT 64.330 185.065 65.980 185.235 ;
        RECT 66.215 185.085 66.565 185.655 ;
        RECT 63.840 184.415 64.145 184.925 ;
        RECT 64.375 184.415 64.655 184.895 ;
        RECT 64.825 184.675 65.085 185.065 ;
        RECT 65.260 184.415 65.515 184.895 ;
        RECT 65.685 184.675 65.980 185.065 ;
        RECT 66.735 184.915 66.905 185.825 ;
        RECT 67.560 185.655 67.805 186.795 ;
        RECT 67.980 186.155 68.240 186.965 ;
        RECT 68.840 186.960 75.115 186.965 ;
        RECT 68.420 185.655 68.670 186.790 ;
        RECT 68.840 186.165 69.100 186.960 ;
        RECT 69.270 186.065 69.530 186.790 ;
        RECT 69.700 186.235 69.960 186.960 ;
        RECT 70.130 186.065 70.390 186.790 ;
        RECT 70.560 186.235 70.820 186.960 ;
        RECT 70.990 186.065 71.250 186.790 ;
        RECT 71.420 186.235 71.680 186.960 ;
        RECT 71.850 186.065 72.110 186.790 ;
        RECT 72.280 186.235 72.525 186.960 ;
        RECT 72.695 186.065 72.955 186.790 ;
        RECT 73.140 186.235 73.385 186.960 ;
        RECT 73.555 186.065 73.815 186.790 ;
        RECT 74.000 186.235 74.245 186.960 ;
        RECT 74.415 186.065 74.675 186.790 ;
        RECT 74.860 186.235 75.115 186.960 ;
        RECT 69.270 186.050 74.675 186.065 ;
        RECT 75.285 186.050 75.575 186.790 ;
        RECT 75.745 186.220 76.015 186.965 ;
        RECT 76.280 186.095 76.545 186.795 ;
        RECT 76.715 186.265 77.045 186.965 ;
        RECT 77.215 186.095 77.885 186.795 ;
        RECT 78.390 186.265 78.820 186.965 ;
        RECT 79.000 186.405 79.190 186.795 ;
        RECT 79.360 186.585 79.690 186.965 ;
        RECT 79.000 186.235 79.730 186.405 ;
        RECT 69.270 185.825 76.015 186.050 ;
        RECT 76.280 185.840 78.855 186.095 ;
        RECT 67.075 185.095 67.390 185.655 ;
        RECT 67.560 185.405 74.680 185.655 ;
        RECT 66.160 184.415 66.435 184.895 ;
        RECT 66.605 184.585 66.905 184.915 ;
        RECT 67.075 184.415 67.380 184.925 ;
        RECT 67.560 184.595 67.810 185.405 ;
        RECT 67.980 184.415 68.240 184.940 ;
        RECT 68.420 184.595 68.670 185.405 ;
        RECT 74.850 185.235 76.015 185.825 ;
        RECT 76.275 185.325 76.550 185.655 ;
        RECT 69.270 185.065 76.015 185.235 ;
        RECT 76.720 185.155 76.900 185.840 ;
        RECT 78.685 185.655 78.855 185.840 ;
        RECT 77.070 185.325 77.430 185.655 ;
        RECT 77.720 185.605 78.010 185.655 ;
        RECT 77.715 185.435 78.010 185.605 ;
        RECT 77.720 185.325 78.010 185.435 ;
        RECT 78.180 185.325 78.515 185.655 ;
        RECT 78.685 185.325 79.365 185.655 ;
        RECT 68.840 184.415 69.100 184.975 ;
        RECT 69.270 184.610 69.530 185.065 ;
        RECT 69.700 184.415 69.960 184.895 ;
        RECT 70.130 184.610 70.390 185.065 ;
        RECT 70.560 184.415 70.820 184.895 ;
        RECT 70.990 184.610 71.250 185.065 ;
        RECT 71.420 184.415 71.665 184.895 ;
        RECT 71.835 184.610 72.110 185.065 ;
        RECT 72.280 184.415 72.525 184.895 ;
        RECT 72.695 184.610 72.955 185.065 ;
        RECT 73.135 184.415 73.385 184.895 ;
        RECT 73.555 184.610 73.815 185.065 ;
        RECT 73.995 184.415 74.245 184.895 ;
        RECT 74.415 184.610 74.675 185.065 ;
        RECT 74.855 184.415 75.115 184.895 ;
        RECT 75.285 184.610 75.545 185.065 ;
        RECT 75.715 184.415 76.015 184.895 ;
        RECT 76.285 184.755 76.900 185.155 ;
        RECT 77.070 184.965 78.340 185.155 ;
        RECT 79.535 185.115 79.730 186.235 ;
        RECT 80.415 185.800 80.705 186.965 ;
        RECT 80.900 185.995 81.200 186.190 ;
        RECT 81.370 186.165 81.625 186.965 ;
        RECT 81.825 186.335 82.155 186.795 ;
        RECT 82.325 186.505 82.900 186.965 ;
        RECT 83.070 186.335 83.425 186.795 ;
        RECT 81.825 186.165 83.425 186.335 ;
        RECT 80.900 185.825 82.150 185.995 ;
        RECT 80.900 185.170 81.070 185.825 ;
        RECT 81.245 185.325 81.590 185.655 ;
        RECT 81.820 185.405 82.150 185.825 ;
        RECT 82.320 185.235 82.600 186.165 ;
        RECT 82.780 185.605 82.970 185.985 ;
        RECT 83.150 185.825 83.425 186.165 ;
        RECT 83.595 185.825 83.925 186.965 ;
        RECT 84.105 185.995 84.435 186.780 ;
        RECT 84.105 185.825 84.785 185.995 ;
        RECT 84.965 185.825 85.295 186.965 ;
        RECT 85.935 185.875 87.145 186.965 ;
        RECT 82.780 185.405 83.925 185.605 ;
        RECT 84.095 185.405 84.445 185.655 ;
        RECT 78.910 184.945 79.730 185.115 ;
        RECT 76.285 184.585 76.620 184.755 ;
        RECT 77.580 184.415 77.915 184.795 ;
        RECT 78.505 184.415 78.740 184.855 ;
        RECT 78.910 184.585 79.240 184.945 ;
        RECT 79.410 184.415 79.740 184.775 ;
        RECT 80.415 184.415 80.705 185.140 ;
        RECT 80.900 184.840 81.135 185.170 ;
        RECT 81.305 184.415 81.635 185.155 ;
        RECT 81.870 184.795 82.145 185.235 ;
        RECT 82.320 185.135 82.645 185.235 ;
        RECT 82.315 184.965 82.645 185.135 ;
        RECT 82.815 185.025 83.925 185.235 ;
        RECT 84.615 185.225 84.785 185.825 ;
        RECT 84.955 185.405 85.305 185.655 ;
        RECT 85.935 185.335 86.455 185.875 ;
        RECT 82.815 184.795 83.065 185.025 ;
        RECT 81.870 184.585 83.065 184.795 ;
        RECT 83.235 184.415 83.405 184.855 ;
        RECT 83.575 184.585 83.925 185.025 ;
        RECT 84.115 184.415 84.355 185.225 ;
        RECT 84.525 184.585 84.855 185.225 ;
        RECT 85.025 184.415 85.295 185.225 ;
        RECT 86.625 185.165 87.145 185.705 ;
        RECT 85.935 184.415 87.145 185.165 ;
        RECT 15.930 184.245 87.230 184.415 ;
        RECT 16.015 183.495 17.225 184.245 ;
        RECT 18.315 183.570 18.575 184.075 ;
        RECT 18.755 183.865 19.085 184.245 ;
        RECT 19.265 183.695 19.435 184.075 ;
        RECT 16.015 182.955 16.535 183.495 ;
        RECT 16.705 182.785 17.225 183.325 ;
        RECT 16.015 181.695 17.225 182.785 ;
        RECT 18.315 182.770 18.485 183.570 ;
        RECT 18.770 183.525 19.435 183.695 ;
        RECT 19.695 183.570 19.955 184.075 ;
        RECT 20.135 183.865 20.465 184.245 ;
        RECT 20.645 183.695 20.815 184.075 ;
        RECT 18.770 183.270 18.940 183.525 ;
        RECT 18.655 182.940 18.940 183.270 ;
        RECT 19.175 182.975 19.505 183.345 ;
        RECT 18.770 182.795 18.940 182.940 ;
        RECT 18.315 181.865 18.585 182.770 ;
        RECT 18.770 182.625 19.435 182.795 ;
        RECT 18.755 181.695 19.085 182.455 ;
        RECT 19.265 181.865 19.435 182.625 ;
        RECT 19.695 182.770 19.875 183.570 ;
        RECT 20.150 183.525 20.815 183.695 ;
        RECT 21.075 183.745 21.335 184.075 ;
        RECT 21.545 183.765 21.820 184.245 ;
        RECT 20.150 183.270 20.320 183.525 ;
        RECT 20.045 182.940 20.320 183.270 ;
        RECT 20.545 182.975 20.885 183.345 ;
        RECT 20.150 182.795 20.320 182.940 ;
        RECT 21.075 182.835 21.245 183.745 ;
        RECT 22.030 183.675 22.235 184.075 ;
        RECT 22.405 183.845 22.740 184.245 ;
        RECT 21.415 183.005 21.775 183.585 ;
        RECT 22.030 183.505 22.715 183.675 ;
        RECT 21.955 182.835 22.205 183.335 ;
        RECT 19.695 181.865 19.965 182.770 ;
        RECT 20.150 182.625 20.825 182.795 ;
        RECT 20.135 181.695 20.465 182.455 ;
        RECT 20.645 181.865 20.825 182.625 ;
        RECT 21.075 182.665 22.205 182.835 ;
        RECT 21.075 181.895 21.345 182.665 ;
        RECT 22.375 182.475 22.715 183.505 ;
        RECT 22.935 183.435 23.175 184.245 ;
        RECT 23.345 183.435 23.675 184.075 ;
        RECT 23.845 183.435 24.115 184.245 ;
        RECT 24.295 183.570 24.555 184.075 ;
        RECT 24.735 183.865 25.065 184.245 ;
        RECT 25.245 183.695 25.415 184.075 ;
        RECT 22.915 183.005 23.265 183.255 ;
        RECT 23.435 182.835 23.605 183.435 ;
        RECT 23.775 183.005 24.125 183.255 ;
        RECT 21.515 181.695 21.845 182.475 ;
        RECT 22.050 182.300 22.715 182.475 ;
        RECT 22.925 182.665 23.605 182.835 ;
        RECT 22.050 181.895 22.235 182.300 ;
        RECT 22.405 181.695 22.740 182.120 ;
        RECT 22.925 181.880 23.255 182.665 ;
        RECT 23.785 181.695 24.115 182.835 ;
        RECT 24.295 182.770 24.475 183.570 ;
        RECT 24.750 183.525 25.415 183.695 ;
        RECT 25.765 183.695 25.935 184.075 ;
        RECT 26.115 183.865 26.445 184.245 ;
        RECT 25.765 183.525 26.430 183.695 ;
        RECT 26.625 183.570 26.885 184.075 ;
        RECT 24.750 183.270 24.920 183.525 ;
        RECT 24.645 182.940 24.920 183.270 ;
        RECT 25.145 182.975 25.485 183.345 ;
        RECT 25.695 182.975 26.035 183.345 ;
        RECT 26.260 183.270 26.430 183.525 ;
        RECT 24.750 182.795 24.920 182.940 ;
        RECT 26.260 182.940 26.535 183.270 ;
        RECT 26.260 182.795 26.430 182.940 ;
        RECT 24.295 181.865 24.565 182.770 ;
        RECT 24.750 182.625 25.425 182.795 ;
        RECT 24.735 181.695 25.065 182.455 ;
        RECT 25.245 181.865 25.425 182.625 ;
        RECT 25.755 182.625 26.430 182.795 ;
        RECT 26.705 182.770 26.885 183.570 ;
        RECT 27.145 183.695 27.315 184.075 ;
        RECT 27.495 183.865 27.825 184.245 ;
        RECT 27.145 183.525 27.810 183.695 ;
        RECT 28.005 183.570 28.265 184.075 ;
        RECT 27.075 182.975 27.415 183.345 ;
        RECT 27.640 183.270 27.810 183.525 ;
        RECT 27.640 182.940 27.915 183.270 ;
        RECT 27.640 182.795 27.810 182.940 ;
        RECT 25.755 181.865 25.935 182.625 ;
        RECT 26.115 181.695 26.445 182.455 ;
        RECT 26.615 181.865 26.885 182.770 ;
        RECT 27.135 182.625 27.810 182.795 ;
        RECT 28.085 182.770 28.265 183.570 ;
        RECT 28.475 183.425 28.705 184.245 ;
        RECT 28.875 183.445 29.205 184.075 ;
        RECT 28.455 183.005 28.785 183.255 ;
        RECT 28.955 182.845 29.205 183.445 ;
        RECT 29.375 183.425 29.585 184.245 ;
        RECT 29.815 183.570 30.075 184.075 ;
        RECT 30.255 183.865 30.585 184.245 ;
        RECT 30.765 183.695 30.935 184.075 ;
        RECT 27.135 181.865 27.315 182.625 ;
        RECT 27.495 181.695 27.825 182.455 ;
        RECT 27.995 181.865 28.265 182.770 ;
        RECT 28.475 181.695 28.705 182.835 ;
        RECT 28.875 181.865 29.205 182.845 ;
        RECT 29.375 181.695 29.585 182.835 ;
        RECT 29.815 182.770 29.995 183.570 ;
        RECT 30.270 183.525 30.935 183.695 ;
        RECT 30.270 183.270 30.440 183.525 ;
        RECT 32.115 183.445 32.425 184.245 ;
        RECT 32.630 183.445 33.325 184.075 ;
        RECT 33.495 183.700 38.840 184.245 ;
        RECT 30.165 182.940 30.440 183.270 ;
        RECT 30.665 182.975 31.005 183.345 ;
        RECT 32.125 183.005 32.460 183.275 ;
        RECT 30.270 182.795 30.440 182.940 ;
        RECT 32.630 182.845 32.800 183.445 ;
        RECT 32.970 183.005 33.305 183.255 ;
        RECT 35.080 182.870 35.420 183.700 ;
        RECT 39.015 183.475 41.605 184.245 ;
        RECT 41.775 183.520 42.065 184.245 ;
        RECT 42.235 183.485 42.945 184.075 ;
        RECT 43.455 183.715 43.785 184.075 ;
        RECT 43.985 183.885 44.315 184.245 ;
        RECT 44.485 183.715 44.815 184.075 ;
        RECT 43.455 183.505 44.815 183.715 ;
        RECT 44.995 183.570 45.255 184.075 ;
        RECT 45.435 183.865 45.765 184.245 ;
        RECT 45.945 183.695 46.115 184.075 ;
        RECT 29.815 181.865 30.085 182.770 ;
        RECT 30.270 182.625 30.945 182.795 ;
        RECT 30.255 181.695 30.585 182.455 ;
        RECT 30.765 181.865 30.945 182.625 ;
        RECT 32.115 181.695 32.395 182.835 ;
        RECT 32.565 181.865 32.895 182.845 ;
        RECT 33.065 181.695 33.325 182.835 ;
        RECT 36.900 182.130 37.250 183.380 ;
        RECT 39.015 182.955 40.225 183.475 ;
        RECT 40.395 182.785 41.605 183.305 ;
        RECT 33.495 181.695 38.840 182.130 ;
        RECT 39.015 181.695 41.605 182.785 ;
        RECT 41.775 181.695 42.065 182.860 ;
        RECT 42.235 182.515 42.440 183.485 ;
        RECT 42.610 182.715 42.940 183.255 ;
        RECT 43.115 183.005 43.610 183.335 ;
        RECT 43.930 183.005 44.305 183.335 ;
        RECT 44.515 183.005 44.825 183.335 ;
        RECT 43.115 182.715 43.440 183.005 ;
        RECT 43.635 182.515 43.965 182.735 ;
        RECT 42.235 182.285 43.965 182.515 ;
        RECT 42.235 181.865 42.935 182.285 ;
        RECT 43.135 181.695 43.465 182.055 ;
        RECT 43.635 181.885 43.965 182.285 ;
        RECT 44.135 182.035 44.305 183.005 ;
        RECT 44.995 182.770 45.175 183.570 ;
        RECT 45.450 183.525 46.115 183.695 ;
        RECT 46.375 183.570 46.635 184.075 ;
        RECT 46.815 183.865 47.145 184.245 ;
        RECT 47.325 183.695 47.495 184.075 ;
        RECT 45.450 183.270 45.620 183.525 ;
        RECT 45.345 182.940 45.620 183.270 ;
        RECT 45.845 182.975 46.185 183.345 ;
        RECT 45.450 182.795 45.620 182.940 ;
        RECT 44.485 181.695 44.815 182.755 ;
        RECT 44.995 181.865 45.265 182.770 ;
        RECT 45.450 182.625 46.125 182.795 ;
        RECT 45.435 181.695 45.765 182.455 ;
        RECT 45.945 181.865 46.125 182.625 ;
        RECT 46.375 182.770 46.555 183.570 ;
        RECT 46.830 183.525 47.495 183.695 ;
        RECT 47.845 183.695 48.015 184.075 ;
        RECT 48.195 183.865 48.525 184.245 ;
        RECT 47.845 183.525 48.510 183.695 ;
        RECT 48.705 183.570 48.965 184.075 ;
        RECT 46.830 183.270 47.000 183.525 ;
        RECT 46.725 182.940 47.000 183.270 ;
        RECT 47.225 182.975 47.565 183.345 ;
        RECT 47.775 182.975 48.115 183.345 ;
        RECT 48.340 183.270 48.510 183.525 ;
        RECT 46.830 182.795 47.000 182.940 ;
        RECT 48.340 182.940 48.615 183.270 ;
        RECT 48.340 182.795 48.510 182.940 ;
        RECT 46.375 181.865 46.645 182.770 ;
        RECT 46.830 182.625 47.505 182.795 ;
        RECT 46.815 181.695 47.145 182.455 ;
        RECT 47.325 181.865 47.505 182.625 ;
        RECT 47.835 182.625 48.510 182.795 ;
        RECT 48.785 182.770 48.965 183.570 ;
        RECT 47.835 181.865 48.015 182.625 ;
        RECT 48.195 181.695 48.525 182.455 ;
        RECT 48.695 181.865 48.965 182.770 ;
        RECT 49.135 183.570 49.395 184.075 ;
        RECT 49.575 183.865 49.905 184.245 ;
        RECT 50.085 183.695 50.255 184.075 ;
        RECT 49.135 182.770 49.315 183.570 ;
        RECT 49.590 183.525 50.255 183.695 ;
        RECT 50.515 183.570 50.775 184.075 ;
        RECT 50.955 183.865 51.285 184.245 ;
        RECT 51.465 183.695 51.635 184.075 ;
        RECT 49.590 183.270 49.760 183.525 ;
        RECT 49.485 182.940 49.760 183.270 ;
        RECT 49.985 182.975 50.325 183.345 ;
        RECT 49.590 182.795 49.760 182.940 ;
        RECT 49.135 181.865 49.405 182.770 ;
        RECT 49.590 182.625 50.265 182.795 ;
        RECT 49.575 181.695 49.905 182.455 ;
        RECT 50.085 181.865 50.265 182.625 ;
        RECT 50.515 182.770 50.695 183.570 ;
        RECT 50.970 183.525 51.635 183.695 ;
        RECT 50.970 183.270 51.140 183.525 ;
        RECT 51.900 183.480 52.355 184.245 ;
        RECT 52.630 183.865 53.930 184.075 ;
        RECT 54.185 183.885 54.515 184.245 ;
        RECT 53.760 183.715 53.930 183.865 ;
        RECT 54.685 183.745 54.945 184.075 ;
        RECT 50.865 182.940 51.140 183.270 ;
        RECT 51.365 182.975 51.705 183.345 ;
        RECT 52.830 183.255 53.050 183.655 ;
        RECT 51.895 183.055 52.385 183.255 ;
        RECT 52.575 183.045 53.050 183.255 ;
        RECT 53.295 183.255 53.505 183.655 ;
        RECT 53.760 183.590 54.515 183.715 ;
        RECT 53.760 183.545 54.605 183.590 ;
        RECT 54.335 183.425 54.605 183.545 ;
        RECT 53.295 183.045 53.625 183.255 ;
        RECT 53.795 182.985 54.205 183.290 ;
        RECT 50.970 182.795 51.140 182.940 ;
        RECT 51.900 182.815 53.075 182.875 ;
        RECT 54.435 182.850 54.605 183.425 ;
        RECT 54.405 182.815 54.605 182.850 ;
        RECT 50.515 181.865 50.785 182.770 ;
        RECT 50.970 182.625 51.645 182.795 ;
        RECT 50.955 181.695 51.285 182.455 ;
        RECT 51.465 181.865 51.645 182.625 ;
        RECT 51.900 182.705 54.605 182.815 ;
        RECT 51.900 182.085 52.155 182.705 ;
        RECT 52.745 182.645 54.545 182.705 ;
        RECT 52.745 182.615 53.075 182.645 ;
        RECT 54.775 182.545 54.945 183.745 ;
        RECT 52.405 182.445 52.590 182.535 ;
        RECT 53.180 182.445 54.015 182.455 ;
        RECT 52.405 182.245 54.015 182.445 ;
        RECT 52.405 182.205 52.635 182.245 ;
        RECT 51.900 181.865 52.235 182.085 ;
        RECT 53.240 181.695 53.595 182.075 ;
        RECT 53.765 181.865 54.015 182.245 ;
        RECT 54.265 181.695 54.515 182.475 ;
        RECT 54.685 181.865 54.945 182.545 ;
        RECT 55.115 183.425 55.800 184.065 ;
        RECT 55.970 183.425 56.140 184.245 ;
        RECT 56.310 183.595 56.640 184.060 ;
        RECT 56.810 183.775 56.980 184.245 ;
        RECT 57.240 183.855 58.425 184.025 ;
        RECT 58.595 183.685 58.925 184.075 ;
        RECT 57.625 183.595 58.010 183.685 ;
        RECT 56.310 183.425 58.010 183.595 ;
        RECT 58.415 183.505 58.925 183.685 ;
        RECT 59.255 183.745 59.515 184.075 ;
        RECT 59.685 183.885 60.015 184.245 ;
        RECT 60.270 183.865 61.570 184.075 ;
        RECT 55.115 182.455 55.365 183.425 ;
        RECT 55.535 183.045 55.870 183.255 ;
        RECT 56.040 183.045 56.490 183.255 ;
        RECT 56.680 183.045 57.165 183.255 ;
        RECT 55.700 182.875 55.870 183.045 ;
        RECT 56.790 182.885 57.165 183.045 ;
        RECT 57.355 183.005 57.735 183.255 ;
        RECT 57.915 183.045 58.245 183.255 ;
        RECT 55.700 182.705 56.620 182.875 ;
        RECT 55.115 181.865 55.780 182.455 ;
        RECT 55.950 181.695 56.280 182.535 ;
        RECT 56.450 182.455 56.620 182.705 ;
        RECT 56.790 182.715 57.185 182.885 ;
        RECT 56.790 182.625 57.165 182.715 ;
        RECT 57.355 182.625 57.675 183.005 ;
        RECT 58.415 182.875 58.585 183.505 ;
        RECT 58.755 183.045 59.085 183.335 ;
        RECT 57.845 182.705 58.930 182.875 ;
        RECT 57.845 182.455 58.015 182.705 ;
        RECT 56.450 182.285 58.015 182.455 ;
        RECT 56.790 181.865 57.595 182.285 ;
        RECT 58.185 181.695 58.435 182.535 ;
        RECT 58.630 181.865 58.930 182.705 ;
        RECT 59.255 182.545 59.425 183.745 ;
        RECT 60.270 183.715 60.440 183.865 ;
        RECT 59.685 183.590 60.440 183.715 ;
        RECT 59.595 183.545 60.440 183.590 ;
        RECT 59.595 183.425 59.865 183.545 ;
        RECT 59.595 182.850 59.765 183.425 ;
        RECT 59.995 182.985 60.405 183.290 ;
        RECT 60.695 183.255 60.905 183.655 ;
        RECT 60.575 183.045 60.905 183.255 ;
        RECT 61.150 183.255 61.370 183.655 ;
        RECT 61.845 183.480 62.300 184.245 ;
        RECT 61.150 183.045 61.625 183.255 ;
        RECT 61.815 183.055 62.305 183.255 ;
        RECT 59.595 182.815 59.795 182.850 ;
        RECT 61.125 182.815 62.300 182.875 ;
        RECT 59.595 182.705 62.300 182.815 ;
        RECT 59.655 182.645 61.455 182.705 ;
        RECT 61.125 182.615 61.455 182.645 ;
        RECT 59.255 181.865 59.515 182.545 ;
        RECT 59.685 181.695 59.935 182.475 ;
        RECT 60.185 182.445 61.020 182.455 ;
        RECT 61.610 182.445 61.795 182.535 ;
        RECT 60.185 182.245 61.795 182.445 ;
        RECT 60.185 181.865 60.435 182.245 ;
        RECT 61.565 182.205 61.795 182.245 ;
        RECT 62.045 182.085 62.300 182.705 ;
        RECT 60.605 181.695 60.960 182.075 ;
        RECT 61.965 181.865 62.300 182.085 ;
        RECT 63.410 181.875 63.690 184.065 ;
        RECT 63.890 183.875 64.620 184.245 ;
        RECT 65.200 183.705 65.630 184.065 ;
        RECT 63.890 183.515 65.630 183.705 ;
        RECT 63.890 183.005 64.150 183.515 ;
        RECT 63.880 181.695 64.165 182.835 ;
        RECT 64.360 182.715 64.620 183.335 ;
        RECT 64.815 182.715 65.240 183.335 ;
        RECT 65.410 183.285 65.630 183.515 ;
        RECT 65.800 183.465 66.045 184.245 ;
        RECT 65.410 182.985 65.955 183.285 ;
        RECT 66.245 183.165 66.475 184.065 ;
        RECT 64.430 182.345 65.455 182.545 ;
        RECT 64.430 181.875 64.600 182.345 ;
        RECT 64.775 181.695 65.105 182.175 ;
        RECT 65.275 181.875 65.455 182.345 ;
        RECT 65.625 181.875 65.955 182.985 ;
        RECT 66.135 182.485 66.475 183.165 ;
        RECT 66.655 182.665 66.885 184.005 ;
        RECT 67.535 183.520 67.825 184.245 ;
        RECT 68.445 183.765 68.615 184.245 ;
        RECT 68.785 183.595 69.115 184.070 ;
        RECT 69.285 183.765 69.455 184.245 ;
        RECT 69.625 183.595 69.955 184.070 ;
        RECT 70.125 183.765 70.295 184.245 ;
        RECT 70.465 183.595 70.795 184.070 ;
        RECT 70.965 183.765 71.135 184.245 ;
        RECT 71.305 183.595 71.635 184.070 ;
        RECT 71.805 183.765 71.975 184.245 ;
        RECT 72.145 183.595 72.475 184.070 ;
        RECT 72.645 183.765 72.815 184.245 ;
        RECT 72.985 183.595 73.315 184.070 ;
        RECT 67.995 183.425 71.635 183.595 ;
        RECT 71.805 183.425 73.315 183.595 ;
        RECT 73.505 183.425 73.835 184.070 ;
        RECT 74.005 183.425 74.175 184.245 ;
        RECT 74.440 183.595 74.710 183.805 ;
        RECT 74.930 183.785 75.260 184.245 ;
        RECT 75.770 183.785 76.520 184.075 ;
        RECT 74.440 183.425 75.775 183.595 ;
        RECT 67.995 182.885 68.380 183.425 ;
        RECT 71.805 183.255 71.975 183.425 ;
        RECT 73.505 183.255 73.675 183.425 ;
        RECT 75.605 183.255 75.775 183.425 ;
        RECT 68.590 183.055 71.975 183.255 ;
        RECT 72.145 183.055 73.675 183.255 ;
        RECT 73.845 183.055 74.265 183.255 ;
        RECT 71.805 182.885 71.975 183.055 ;
        RECT 66.135 182.285 66.885 182.485 ;
        RECT 66.125 181.695 66.475 182.105 ;
        RECT 66.645 181.895 66.885 182.285 ;
        RECT 67.535 181.695 67.825 182.860 ;
        RECT 67.995 182.715 71.635 182.885 ;
        RECT 71.805 182.715 73.315 182.885 ;
        RECT 68.445 181.695 68.615 182.495 ;
        RECT 68.785 181.865 69.115 182.715 ;
        RECT 69.285 181.695 69.455 182.495 ;
        RECT 69.625 181.865 69.955 182.715 ;
        RECT 70.125 181.695 70.295 182.495 ;
        RECT 70.465 181.865 70.795 182.715 ;
        RECT 70.965 181.695 71.135 182.495 ;
        RECT 71.305 181.865 71.635 182.715 ;
        RECT 71.805 181.695 71.975 182.545 ;
        RECT 72.145 181.865 72.475 182.715 ;
        RECT 72.645 181.695 72.815 182.545 ;
        RECT 72.985 181.865 73.315 182.715 ;
        RECT 73.505 182.785 73.675 183.055 ;
        RECT 74.440 183.015 74.790 183.255 ;
        RECT 74.960 183.015 75.435 183.255 ;
        RECT 75.605 183.005 75.980 183.255 ;
        RECT 73.505 181.865 73.835 182.785 ;
        RECT 74.005 181.695 74.175 182.885 ;
        RECT 75.605 182.835 75.775 183.005 ;
        RECT 74.440 182.665 75.775 182.835 ;
        RECT 74.440 182.505 74.720 182.665 ;
        RECT 76.150 182.495 76.520 183.785 ;
        RECT 76.825 183.765 77.125 184.245 ;
        RECT 77.295 183.595 77.555 184.050 ;
        RECT 77.725 183.765 77.985 184.245 ;
        RECT 78.165 183.595 78.425 184.050 ;
        RECT 78.595 183.765 78.845 184.245 ;
        RECT 79.025 183.595 79.285 184.050 ;
        RECT 79.455 183.765 79.705 184.245 ;
        RECT 79.885 183.595 80.145 184.050 ;
        RECT 80.315 183.765 80.560 184.245 ;
        RECT 80.730 183.595 81.005 184.050 ;
        RECT 81.175 183.765 81.420 184.245 ;
        RECT 81.590 183.595 81.850 184.050 ;
        RECT 82.020 183.765 82.280 184.245 ;
        RECT 82.450 183.595 82.710 184.050 ;
        RECT 82.880 183.765 83.140 184.245 ;
        RECT 83.310 183.595 83.570 184.050 ;
        RECT 83.740 183.685 84.000 184.245 ;
        RECT 76.825 183.425 83.570 183.595 ;
        RECT 76.825 182.835 77.990 183.425 ;
        RECT 84.170 183.255 84.420 184.065 ;
        RECT 84.600 183.720 84.860 184.245 ;
        RECT 85.030 183.255 85.280 184.065 ;
        RECT 85.460 183.735 85.765 184.245 ;
        RECT 78.160 183.005 85.280 183.255 ;
        RECT 85.450 183.005 85.765 183.565 ;
        RECT 85.935 183.495 87.145 184.245 ;
        RECT 76.825 182.610 83.570 182.835 ;
        RECT 74.930 181.695 75.180 182.495 ;
        RECT 75.350 182.325 76.520 182.495 ;
        RECT 75.350 181.865 75.680 182.325 ;
        RECT 75.850 181.695 76.065 182.155 ;
        RECT 76.825 181.695 77.095 182.440 ;
        RECT 77.265 181.870 77.555 182.610 ;
        RECT 78.165 182.595 83.570 182.610 ;
        RECT 77.725 181.700 77.980 182.425 ;
        RECT 78.165 181.870 78.425 182.595 ;
        RECT 78.595 181.700 78.840 182.425 ;
        RECT 79.025 181.870 79.285 182.595 ;
        RECT 79.455 181.700 79.700 182.425 ;
        RECT 79.885 181.870 80.145 182.595 ;
        RECT 80.315 181.700 80.560 182.425 ;
        RECT 80.730 181.870 80.990 182.595 ;
        RECT 81.160 181.700 81.420 182.425 ;
        RECT 81.590 181.870 81.850 182.595 ;
        RECT 82.020 181.700 82.280 182.425 ;
        RECT 82.450 181.870 82.710 182.595 ;
        RECT 82.880 181.700 83.140 182.425 ;
        RECT 83.310 181.870 83.570 182.595 ;
        RECT 83.740 181.700 84.000 182.495 ;
        RECT 84.170 181.870 84.420 183.005 ;
        RECT 77.725 181.695 84.000 181.700 ;
        RECT 84.600 181.695 84.860 182.505 ;
        RECT 85.035 181.865 85.280 183.005 ;
        RECT 85.935 182.785 86.455 183.325 ;
        RECT 86.625 182.955 87.145 183.495 ;
        RECT 85.460 181.695 85.755 182.505 ;
        RECT 85.935 181.695 87.145 182.785 ;
        RECT 15.930 181.525 87.230 181.695 ;
        RECT 16.015 180.435 17.225 181.525 ;
        RECT 16.015 179.725 16.535 180.265 ;
        RECT 16.705 179.895 17.225 180.435 ;
        RECT 18.500 180.555 18.890 180.730 ;
        RECT 19.375 180.725 19.705 181.525 ;
        RECT 19.875 180.735 20.410 181.355 ;
        RECT 18.500 180.385 19.925 180.555 ;
        RECT 16.015 178.975 17.225 179.725 ;
        RECT 18.375 179.655 18.730 180.215 ;
        RECT 18.900 179.485 19.070 180.385 ;
        RECT 19.240 179.655 19.505 180.215 ;
        RECT 19.755 179.885 19.925 180.385 ;
        RECT 20.095 179.715 20.410 180.735 ;
        RECT 20.615 180.570 20.885 181.525 ;
        RECT 18.480 178.975 18.720 179.485 ;
        RECT 18.900 179.155 19.180 179.485 ;
        RECT 19.410 178.975 19.625 179.485 ;
        RECT 19.795 179.145 20.410 179.715 ;
        RECT 21.070 180.470 21.375 181.255 ;
        RECT 21.555 181.055 22.240 181.525 ;
        RECT 21.550 180.535 22.245 180.845 ;
        RECT 21.070 179.665 21.245 180.470 ;
        RECT 22.420 180.365 22.705 181.310 ;
        RECT 22.905 181.075 23.235 181.525 ;
        RECT 23.405 180.905 23.575 181.335 ;
        RECT 21.845 180.215 22.705 180.365 ;
        RECT 21.415 180.195 22.705 180.215 ;
        RECT 22.895 180.675 23.575 180.905 ;
        RECT 23.925 180.905 24.095 181.335 ;
        RECT 24.265 181.075 24.595 181.525 ;
        RECT 23.925 180.675 24.600 180.905 ;
        RECT 21.415 179.835 22.405 180.195 ;
        RECT 22.895 180.025 23.130 180.675 ;
        RECT 20.615 178.975 20.885 179.610 ;
        RECT 21.070 179.145 21.305 179.665 ;
        RECT 22.235 179.500 22.405 179.835 ;
        RECT 22.575 179.695 23.130 180.025 ;
        RECT 22.915 179.545 23.130 179.695 ;
        RECT 23.300 180.335 23.605 180.505 ;
        RECT 23.300 179.655 23.600 180.335 ;
        RECT 23.895 179.655 24.195 180.505 ;
        RECT 24.365 180.025 24.600 180.675 ;
        RECT 24.770 180.365 25.055 181.310 ;
        RECT 25.235 181.055 25.920 181.525 ;
        RECT 25.230 180.535 25.925 180.845 ;
        RECT 26.100 180.470 26.405 181.255 ;
        RECT 24.770 180.215 25.630 180.365 ;
        RECT 24.770 180.195 26.055 180.215 ;
        RECT 24.365 179.695 24.900 180.025 ;
        RECT 25.070 179.835 26.055 180.195 ;
        RECT 24.365 179.545 24.585 179.695 ;
        RECT 21.475 178.975 21.875 179.470 ;
        RECT 22.235 179.305 22.635 179.500 ;
        RECT 22.465 179.160 22.635 179.305 ;
        RECT 22.915 179.170 23.155 179.545 ;
        RECT 23.325 178.975 23.655 179.480 ;
        RECT 23.840 178.975 24.175 179.480 ;
        RECT 24.345 179.170 24.585 179.545 ;
        RECT 25.070 179.500 25.240 179.835 ;
        RECT 26.230 179.665 26.405 180.470 ;
        RECT 27.065 180.915 27.395 181.345 ;
        RECT 27.575 181.085 27.770 181.525 ;
        RECT 27.940 180.915 28.270 181.345 ;
        RECT 27.065 180.745 28.270 180.915 ;
        RECT 27.065 180.415 27.960 180.745 ;
        RECT 28.440 180.575 28.715 181.345 ;
        RECT 28.130 180.385 28.715 180.575 ;
        RECT 27.070 179.885 27.365 180.215 ;
        RECT 27.545 179.885 27.960 180.215 ;
        RECT 24.865 179.305 25.240 179.500 ;
        RECT 24.865 179.160 25.035 179.305 ;
        RECT 25.600 178.975 25.995 179.470 ;
        RECT 26.165 179.145 26.405 179.665 ;
        RECT 27.065 178.975 27.365 179.705 ;
        RECT 27.545 179.265 27.775 179.885 ;
        RECT 28.130 179.715 28.305 180.385 ;
        RECT 28.895 180.360 29.185 181.525 ;
        RECT 30.285 180.465 30.615 181.315 ;
        RECT 30.285 180.335 30.505 180.465 ;
        RECT 30.785 180.385 31.035 181.525 ;
        RECT 31.225 180.885 31.475 181.305 ;
        RECT 31.705 181.055 32.035 181.525 ;
        RECT 32.265 180.885 32.515 181.305 ;
        RECT 31.225 180.715 32.515 180.885 ;
        RECT 32.695 180.885 33.025 181.315 ;
        RECT 32.695 180.715 33.150 180.885 ;
        RECT 27.975 179.535 28.305 179.715 ;
        RECT 28.475 179.565 28.715 180.215 ;
        RECT 30.285 179.700 30.475 180.335 ;
        RECT 31.215 180.215 31.430 180.545 ;
        RECT 30.645 179.885 30.955 180.215 ;
        RECT 31.125 179.885 31.430 180.215 ;
        RECT 31.605 179.885 31.890 180.545 ;
        RECT 32.085 179.885 32.350 180.545 ;
        RECT 32.565 179.885 32.810 180.545 ;
        RECT 30.785 179.715 30.955 179.885 ;
        RECT 32.980 179.715 33.150 180.715 ;
        RECT 33.500 180.385 33.820 181.525 ;
        RECT 34.000 180.215 34.195 181.265 ;
        RECT 34.375 180.675 34.705 181.355 ;
        RECT 34.905 180.725 35.160 181.525 ;
        RECT 35.355 180.685 35.610 181.355 ;
        RECT 35.780 180.765 36.110 181.525 ;
        RECT 36.280 180.925 36.530 181.355 ;
        RECT 36.700 181.105 37.055 181.525 ;
        RECT 37.245 181.185 38.415 181.355 ;
        RECT 37.245 181.145 37.575 181.185 ;
        RECT 37.685 180.925 37.915 181.015 ;
        RECT 36.280 180.685 37.915 180.925 ;
        RECT 38.085 180.685 38.415 181.185 ;
        RECT 35.355 180.675 35.565 180.685 ;
        RECT 34.375 180.395 34.725 180.675 ;
        RECT 33.560 180.165 33.820 180.215 ;
        RECT 33.555 179.995 33.820 180.165 ;
        RECT 33.560 179.885 33.820 179.995 ;
        RECT 34.000 179.885 34.385 180.215 ;
        RECT 34.555 180.015 34.725 180.395 ;
        RECT 34.915 180.185 35.160 180.545 ;
        RECT 34.555 179.845 35.075 180.015 ;
        RECT 27.975 179.155 28.200 179.535 ;
        RECT 28.370 178.975 28.700 179.365 ;
        RECT 28.895 178.975 29.185 179.700 ;
        RECT 30.285 179.190 30.615 179.700 ;
        RECT 30.785 179.545 33.150 179.715 ;
        RECT 30.785 178.975 31.115 179.375 ;
        RECT 32.165 179.205 32.495 179.545 ;
        RECT 33.500 179.505 34.715 179.675 ;
        RECT 32.665 178.975 32.995 179.375 ;
        RECT 33.500 179.155 33.790 179.505 ;
        RECT 33.985 178.975 34.315 179.335 ;
        RECT 34.485 179.200 34.715 179.505 ;
        RECT 34.905 179.280 35.075 179.845 ;
        RECT 35.355 179.555 35.525 180.675 ;
        RECT 38.585 180.515 38.755 181.355 ;
        RECT 35.695 180.345 38.755 180.515 ;
        RECT 39.020 180.805 39.355 181.315 ;
        RECT 35.695 179.795 35.865 180.345 ;
        RECT 36.095 179.965 36.460 180.165 ;
        RECT 36.630 179.965 36.960 180.165 ;
        RECT 35.695 179.625 36.495 179.795 ;
        RECT 35.355 179.475 35.540 179.555 ;
        RECT 35.355 179.145 35.610 179.475 ;
        RECT 35.825 178.975 36.155 179.455 ;
        RECT 36.325 179.395 36.495 179.625 ;
        RECT 36.675 179.565 36.960 179.965 ;
        RECT 37.230 179.965 37.705 180.165 ;
        RECT 37.875 179.965 38.320 180.165 ;
        RECT 38.490 179.965 38.840 180.175 ;
        RECT 37.230 179.565 37.510 179.965 ;
        RECT 37.690 179.625 38.755 179.795 ;
        RECT 37.690 179.395 37.860 179.625 ;
        RECT 36.325 179.145 37.860 179.395 ;
        RECT 38.085 178.975 38.415 179.455 ;
        RECT 38.585 179.145 38.755 179.625 ;
        RECT 39.020 179.450 39.275 180.805 ;
        RECT 39.605 180.725 39.935 181.525 ;
        RECT 40.180 180.935 40.465 181.355 ;
        RECT 40.720 181.105 41.050 181.525 ;
        RECT 41.275 181.185 42.435 181.355 ;
        RECT 41.275 180.935 41.605 181.185 ;
        RECT 40.180 180.765 41.605 180.935 ;
        RECT 41.835 180.555 42.005 181.015 ;
        RECT 42.265 180.685 42.435 181.185 ;
        RECT 39.635 180.385 42.005 180.555 ;
        RECT 39.635 180.215 39.805 180.385 ;
        RECT 42.255 180.335 42.465 180.505 ;
        RECT 42.695 180.415 42.955 181.355 ;
        RECT 43.125 181.125 43.455 181.525 ;
        RECT 44.600 181.260 44.855 181.355 ;
        RECT 43.715 181.090 44.855 181.260 ;
        RECT 45.025 181.145 45.355 181.315 ;
        RECT 43.715 180.865 43.885 181.090 ;
        RECT 43.125 180.695 43.885 180.865 ;
        RECT 44.600 180.955 44.855 181.090 ;
        RECT 42.255 180.215 42.460 180.335 ;
        RECT 39.500 179.885 39.805 180.215 ;
        RECT 40.000 180.165 40.250 180.215 ;
        RECT 39.995 179.995 40.250 180.165 ;
        RECT 40.000 179.885 40.250 179.995 ;
        RECT 39.635 179.715 39.805 179.885 ;
        RECT 40.460 179.825 40.730 180.215 ;
        RECT 40.920 180.165 41.210 180.215 ;
        RECT 40.915 179.995 41.210 180.165 ;
        RECT 39.635 179.545 40.195 179.715 ;
        RECT 40.455 179.655 40.730 179.825 ;
        RECT 40.460 179.555 40.730 179.655 ;
        RECT 40.920 179.555 41.210 179.995 ;
        RECT 41.380 179.550 41.800 180.215 ;
        RECT 42.110 179.885 42.460 180.215 ;
        RECT 42.695 179.700 42.870 180.415 ;
        RECT 43.125 180.215 43.295 180.695 ;
        RECT 44.150 180.605 44.320 180.795 ;
        RECT 44.600 180.785 45.010 180.955 ;
        RECT 43.040 179.885 43.295 180.215 ;
        RECT 43.520 179.885 43.850 180.505 ;
        RECT 44.150 180.435 44.670 180.605 ;
        RECT 44.020 179.885 44.310 180.265 ;
        RECT 44.500 179.715 44.670 180.435 ;
        RECT 39.020 179.190 39.355 179.450 ;
        RECT 40.025 179.375 40.195 179.545 ;
        RECT 39.525 178.975 39.855 179.375 ;
        RECT 40.025 179.205 41.640 179.375 ;
        RECT 42.185 178.975 42.515 179.695 ;
        RECT 42.695 179.145 42.955 179.700 ;
        RECT 43.790 179.545 44.670 179.715 ;
        RECT 44.840 179.760 45.010 180.785 ;
        RECT 45.185 180.895 45.355 181.145 ;
        RECT 45.525 181.065 45.775 181.525 ;
        RECT 45.945 180.895 46.125 181.355 ;
        RECT 45.185 180.725 46.125 180.895 ;
        RECT 46.840 180.725 47.095 181.525 ;
        RECT 47.295 180.675 47.625 181.355 ;
        RECT 45.210 180.245 45.690 180.545 ;
        RECT 44.840 179.590 45.190 179.760 ;
        RECT 45.430 179.655 45.690 180.245 ;
        RECT 45.890 179.655 46.150 180.545 ;
        RECT 46.840 180.185 47.085 180.545 ;
        RECT 47.275 180.395 47.625 180.675 ;
        RECT 47.275 180.015 47.445 180.395 ;
        RECT 47.805 180.215 48.000 181.265 ;
        RECT 48.180 180.385 48.500 181.525 ;
        RECT 48.695 180.470 49.000 181.255 ;
        RECT 49.180 181.055 49.865 181.525 ;
        RECT 49.175 180.535 49.870 180.845 ;
        RECT 46.925 179.845 47.445 180.015 ;
        RECT 47.615 179.885 48.000 180.215 ;
        RECT 48.180 180.165 48.440 180.215 ;
        RECT 48.180 179.995 48.445 180.165 ;
        RECT 48.180 179.885 48.440 179.995 ;
        RECT 46.925 179.825 47.095 179.845 ;
        RECT 46.895 179.655 47.095 179.825 ;
        RECT 43.125 178.975 43.555 179.420 ;
        RECT 43.790 179.145 43.960 179.545 ;
        RECT 44.130 178.975 44.850 179.375 ;
        RECT 45.020 179.145 45.190 179.590 ;
        RECT 45.765 178.975 46.165 179.485 ;
        RECT 46.925 179.280 47.095 179.655 ;
        RECT 47.285 179.505 48.500 179.675 ;
        RECT 47.285 179.200 47.515 179.505 ;
        RECT 47.685 178.975 48.015 179.335 ;
        RECT 48.210 179.155 48.500 179.505 ;
        RECT 48.695 179.665 48.870 180.470 ;
        RECT 50.045 180.365 50.330 181.310 ;
        RECT 50.505 181.075 50.835 181.525 ;
        RECT 51.005 180.905 51.175 181.335 ;
        RECT 49.470 180.215 50.330 180.365 ;
        RECT 49.045 180.195 50.330 180.215 ;
        RECT 50.500 180.675 51.175 180.905 ;
        RECT 51.525 180.905 51.695 181.335 ;
        RECT 51.865 181.075 52.195 181.525 ;
        RECT 51.525 180.675 52.200 180.905 ;
        RECT 49.045 179.835 50.030 180.195 ;
        RECT 50.500 180.025 50.735 180.675 ;
        RECT 48.695 179.145 48.935 179.665 ;
        RECT 49.860 179.500 50.030 179.835 ;
        RECT 50.200 179.695 50.735 180.025 ;
        RECT 50.515 179.545 50.735 179.695 ;
        RECT 50.905 179.655 51.205 180.505 ;
        RECT 51.495 179.655 51.795 180.505 ;
        RECT 51.965 180.025 52.200 180.675 ;
        RECT 52.370 180.365 52.655 181.310 ;
        RECT 52.835 181.055 53.520 181.525 ;
        RECT 52.830 180.535 53.525 180.845 ;
        RECT 53.700 180.470 54.005 181.255 ;
        RECT 52.370 180.215 53.230 180.365 ;
        RECT 52.370 180.195 53.655 180.215 ;
        RECT 51.965 179.695 52.500 180.025 ;
        RECT 52.670 179.835 53.655 180.195 ;
        RECT 51.965 179.545 52.185 179.695 ;
        RECT 49.105 178.975 49.500 179.470 ;
        RECT 49.860 179.305 50.235 179.500 ;
        RECT 50.065 179.160 50.235 179.305 ;
        RECT 50.515 179.170 50.755 179.545 ;
        RECT 50.925 178.975 51.260 179.480 ;
        RECT 51.440 178.975 51.775 179.480 ;
        RECT 51.945 179.170 52.185 179.545 ;
        RECT 52.670 179.500 52.840 179.835 ;
        RECT 53.830 179.665 54.005 180.470 ;
        RECT 54.655 180.360 54.945 181.525 ;
        RECT 55.120 181.135 55.455 181.355 ;
        RECT 56.460 181.145 56.815 181.525 ;
        RECT 55.120 180.515 55.375 181.135 ;
        RECT 55.625 180.975 55.855 181.015 ;
        RECT 56.985 180.975 57.235 181.355 ;
        RECT 55.625 180.775 57.235 180.975 ;
        RECT 55.625 180.685 55.810 180.775 ;
        RECT 56.400 180.765 57.235 180.775 ;
        RECT 57.485 180.745 57.735 181.525 ;
        RECT 57.905 180.675 58.165 181.355 ;
        RECT 55.965 180.575 56.295 180.605 ;
        RECT 55.965 180.515 57.765 180.575 ;
        RECT 55.120 180.405 57.825 180.515 ;
        RECT 55.120 180.345 56.295 180.405 ;
        RECT 57.625 180.370 57.825 180.405 ;
        RECT 55.115 179.965 55.605 180.165 ;
        RECT 55.795 179.965 56.270 180.175 ;
        RECT 52.465 179.305 52.840 179.500 ;
        RECT 52.465 179.160 52.635 179.305 ;
        RECT 53.200 178.975 53.595 179.470 ;
        RECT 53.765 179.145 54.005 179.665 ;
        RECT 54.655 178.975 54.945 179.700 ;
        RECT 55.120 178.975 55.575 179.740 ;
        RECT 56.050 179.565 56.270 179.965 ;
        RECT 56.515 179.965 56.845 180.175 ;
        RECT 56.515 179.565 56.725 179.965 ;
        RECT 57.015 179.930 57.425 180.235 ;
        RECT 57.655 179.795 57.825 180.370 ;
        RECT 57.555 179.675 57.825 179.795 ;
        RECT 56.980 179.630 57.825 179.675 ;
        RECT 56.980 179.505 57.735 179.630 ;
        RECT 56.980 179.355 57.150 179.505 ;
        RECT 57.995 179.475 58.165 180.675 ;
        RECT 59.265 181.185 60.435 181.355 ;
        RECT 59.265 180.515 59.595 181.185 ;
        RECT 60.105 181.145 60.435 181.185 ;
        RECT 60.605 181.145 60.980 181.525 ;
        RECT 59.765 180.975 59.995 181.015 ;
        RECT 59.765 180.925 60.380 180.975 ;
        RECT 61.125 180.925 61.295 181.055 ;
        RECT 59.765 180.725 61.295 180.925 ;
        RECT 61.530 180.745 61.795 181.525 ;
        RECT 59.765 180.685 60.645 180.725 ;
        RECT 62.105 180.595 62.275 181.355 ;
        RECT 62.490 180.765 62.820 181.525 ;
        RECT 60.785 180.515 61.845 180.555 ;
        RECT 59.265 180.385 61.845 180.515 ;
        RECT 62.105 180.425 62.820 180.595 ;
        RECT 62.990 180.450 63.245 181.355 ;
        RECT 59.265 180.335 61.010 180.385 ;
        RECT 59.295 179.655 59.745 180.165 ;
        RECT 59.935 179.965 60.410 180.165 ;
        RECT 60.160 179.565 60.410 179.965 ;
        RECT 60.660 179.965 61.010 180.165 ;
        RECT 60.660 179.565 60.870 179.965 ;
        RECT 61.180 179.885 61.505 180.215 ;
        RECT 61.675 179.715 61.845 180.385 ;
        RECT 62.015 179.875 62.370 180.245 ;
        RECT 62.650 180.215 62.820 180.425 ;
        RECT 62.650 179.885 62.905 180.215 ;
        RECT 61.115 179.545 61.845 179.715 ;
        RECT 62.650 179.695 62.820 179.885 ;
        RECT 63.075 179.720 63.245 180.450 ;
        RECT 63.420 180.375 63.680 181.525 ;
        RECT 63.855 180.385 64.195 181.355 ;
        RECT 64.365 180.385 64.535 181.525 ;
        RECT 64.805 180.725 65.055 181.525 ;
        RECT 65.700 180.555 66.030 181.355 ;
        RECT 66.330 180.725 66.660 181.525 ;
        RECT 66.830 180.555 67.160 181.355 ;
        RECT 64.725 180.385 67.160 180.555 ;
        RECT 67.575 180.385 67.805 181.525 ;
        RECT 55.850 179.145 57.150 179.355 ;
        RECT 57.405 178.975 57.735 179.335 ;
        RECT 57.905 179.145 58.165 179.475 ;
        RECT 59.265 178.975 59.715 179.485 ;
        RECT 61.115 179.395 61.295 179.545 ;
        RECT 59.990 179.145 61.295 179.395 ;
        RECT 62.105 179.525 62.820 179.695 ;
        RECT 61.475 178.975 61.805 179.375 ;
        RECT 62.105 179.145 62.275 179.525 ;
        RECT 62.490 178.975 62.820 179.355 ;
        RECT 62.990 179.145 63.245 179.720 ;
        RECT 63.420 178.975 63.680 179.815 ;
        RECT 63.855 179.775 64.030 180.385 ;
        RECT 64.725 180.135 64.895 180.385 ;
        RECT 64.200 179.965 64.895 180.135 ;
        RECT 65.070 179.965 65.490 180.165 ;
        RECT 65.660 179.965 65.990 180.165 ;
        RECT 66.160 179.965 66.490 180.165 ;
        RECT 63.855 179.145 64.195 179.775 ;
        RECT 64.365 178.975 64.615 179.775 ;
        RECT 64.805 179.625 66.030 179.795 ;
        RECT 64.805 179.145 65.135 179.625 ;
        RECT 65.305 178.975 65.530 179.435 ;
        RECT 65.700 179.145 66.030 179.625 ;
        RECT 66.660 179.755 66.830 180.385 ;
        RECT 67.975 180.375 68.305 181.355 ;
        RECT 68.475 180.385 68.685 181.525 ;
        RECT 68.925 180.715 69.220 181.525 ;
        RECT 67.015 179.965 67.365 180.215 ;
        RECT 67.555 179.965 67.885 180.215 ;
        RECT 66.660 179.145 67.160 179.755 ;
        RECT 67.575 178.975 67.805 179.795 ;
        RECT 68.055 179.775 68.305 180.375 ;
        RECT 69.400 180.215 69.645 181.355 ;
        RECT 69.820 180.715 70.080 181.525 ;
        RECT 70.680 181.520 76.955 181.525 ;
        RECT 70.260 180.215 70.510 181.350 ;
        RECT 70.680 180.725 70.940 181.520 ;
        RECT 71.110 180.625 71.370 181.350 ;
        RECT 71.540 180.795 71.800 181.520 ;
        RECT 71.970 180.625 72.230 181.350 ;
        RECT 72.400 180.795 72.660 181.520 ;
        RECT 72.830 180.625 73.090 181.350 ;
        RECT 73.260 180.795 73.520 181.520 ;
        RECT 73.690 180.625 73.950 181.350 ;
        RECT 74.120 180.795 74.365 181.520 ;
        RECT 74.535 180.625 74.795 181.350 ;
        RECT 74.980 180.795 75.225 181.520 ;
        RECT 75.395 180.625 75.655 181.350 ;
        RECT 75.840 180.795 76.085 181.520 ;
        RECT 76.255 180.625 76.515 181.350 ;
        RECT 76.700 180.795 76.955 181.520 ;
        RECT 71.110 180.610 76.515 180.625 ;
        RECT 77.125 180.610 77.415 181.350 ;
        RECT 77.585 180.780 77.855 181.525 ;
        RECT 71.110 180.385 77.855 180.610 ;
        RECT 67.975 179.145 68.305 179.775 ;
        RECT 68.475 178.975 68.685 179.795 ;
        RECT 68.915 179.655 69.230 180.215 ;
        RECT 69.400 179.965 76.520 180.215 ;
        RECT 68.915 178.975 69.220 179.485 ;
        RECT 69.400 179.155 69.650 179.965 ;
        RECT 69.820 178.975 70.080 179.500 ;
        RECT 70.260 179.155 70.510 179.965 ;
        RECT 76.690 179.795 77.855 180.385 ;
        RECT 78.120 180.555 78.395 181.355 ;
        RECT 78.565 180.725 78.895 181.525 ;
        RECT 79.065 181.185 80.205 181.355 ;
        RECT 79.065 180.555 79.235 181.185 ;
        RECT 78.120 180.345 79.235 180.555 ;
        RECT 79.405 180.555 79.735 181.015 ;
        RECT 79.905 180.725 80.205 181.185 ;
        RECT 79.405 180.335 80.165 180.555 ;
        RECT 80.415 180.360 80.705 181.525 ;
        RECT 80.880 180.525 81.135 181.525 ;
        RECT 78.120 179.965 78.840 180.165 ;
        RECT 79.010 179.965 79.780 180.165 ;
        RECT 79.950 179.795 80.165 180.335 ;
        RECT 71.110 179.625 77.855 179.795 ;
        RECT 70.680 178.975 70.940 179.535 ;
        RECT 71.110 179.170 71.370 179.625 ;
        RECT 71.540 178.975 71.800 179.455 ;
        RECT 71.970 179.170 72.230 179.625 ;
        RECT 72.400 178.975 72.660 179.455 ;
        RECT 72.830 179.170 73.090 179.625 ;
        RECT 73.260 178.975 73.505 179.455 ;
        RECT 73.675 179.170 73.950 179.625 ;
        RECT 74.120 178.975 74.365 179.455 ;
        RECT 74.535 179.170 74.795 179.625 ;
        RECT 74.975 178.975 75.225 179.455 ;
        RECT 75.395 179.170 75.655 179.625 ;
        RECT 75.835 178.975 76.085 179.455 ;
        RECT 76.255 179.170 76.515 179.625 ;
        RECT 76.695 178.975 76.955 179.455 ;
        RECT 77.125 179.170 77.385 179.625 ;
        RECT 77.555 178.975 77.855 179.455 ;
        RECT 78.120 178.975 78.395 179.795 ;
        RECT 78.565 179.625 80.165 179.795 ;
        RECT 78.565 179.615 79.735 179.625 ;
        RECT 78.565 179.145 78.895 179.615 ;
        RECT 79.065 178.975 79.235 179.445 ;
        RECT 79.405 179.145 79.735 179.615 ;
        RECT 79.905 178.975 80.195 179.445 ;
        RECT 80.415 178.975 80.705 179.700 ;
        RECT 80.895 178.975 81.135 179.775 ;
        RECT 81.320 179.145 81.565 181.355 ;
        RECT 81.735 181.075 82.585 181.525 ;
        RECT 82.755 180.895 83.015 181.355 ;
        RECT 81.895 180.675 83.015 180.895 ;
        RECT 83.195 180.845 83.400 180.875 ;
        RECT 83.195 180.675 83.405 180.845 ;
        RECT 81.895 180.220 82.065 180.675 ;
        RECT 81.735 179.730 82.065 180.220 ;
        RECT 82.235 179.900 82.645 180.505 ;
        RECT 83.195 180.290 83.400 180.675 ;
        RECT 83.585 180.540 83.910 181.525 ;
        RECT 84.185 180.595 84.355 181.355 ;
        RECT 84.570 180.765 84.900 181.525 ;
        RECT 84.185 180.425 84.900 180.595 ;
        RECT 85.070 180.450 85.325 181.355 ;
        RECT 82.815 179.915 83.400 180.290 ;
        RECT 83.655 179.885 83.915 180.340 ;
        RECT 84.095 179.875 84.450 180.245 ;
        RECT 84.730 180.215 84.900 180.425 ;
        RECT 84.730 179.885 84.985 180.215 ;
        RECT 81.735 179.525 82.585 179.730 ;
        RECT 81.735 178.975 82.065 179.355 ;
        RECT 82.255 179.145 82.585 179.525 ;
        RECT 82.755 179.525 83.910 179.715 ;
        RECT 84.730 179.695 84.900 179.885 ;
        RECT 85.155 179.720 85.325 180.450 ;
        RECT 85.500 180.375 85.760 181.525 ;
        RECT 85.935 180.435 87.145 181.525 ;
        RECT 85.935 179.895 86.455 180.435 ;
        RECT 82.755 179.355 82.965 179.525 ;
        RECT 83.635 179.385 83.910 179.525 ;
        RECT 84.185 179.525 84.900 179.695 ;
        RECT 83.135 178.975 83.465 179.355 ;
        RECT 84.185 179.145 84.355 179.525 ;
        RECT 84.570 178.975 84.900 179.355 ;
        RECT 85.070 179.145 85.325 179.720 ;
        RECT 85.500 178.975 85.760 179.815 ;
        RECT 86.625 179.725 87.145 180.265 ;
        RECT 85.935 178.975 87.145 179.725 ;
        RECT 15.930 178.805 87.230 178.975 ;
        RECT 16.015 178.055 17.225 178.805 ;
        RECT 17.485 178.255 17.655 178.635 ;
        RECT 17.835 178.425 18.165 178.805 ;
        RECT 17.485 178.085 18.150 178.255 ;
        RECT 18.345 178.130 18.605 178.635 ;
        RECT 16.015 177.515 16.535 178.055 ;
        RECT 16.705 177.345 17.225 177.885 ;
        RECT 17.415 177.535 17.755 177.905 ;
        RECT 17.980 177.830 18.150 178.085 ;
        RECT 17.980 177.500 18.255 177.830 ;
        RECT 17.980 177.355 18.150 177.500 ;
        RECT 16.015 176.255 17.225 177.345 ;
        RECT 17.475 177.185 18.150 177.355 ;
        RECT 18.425 177.330 18.605 178.130 ;
        RECT 19.700 178.155 19.970 178.365 ;
        RECT 20.190 178.345 20.520 178.805 ;
        RECT 21.030 178.345 21.780 178.635 ;
        RECT 19.700 177.985 21.035 178.155 ;
        RECT 20.865 177.815 21.035 177.985 ;
        RECT 19.700 177.575 20.050 177.815 ;
        RECT 20.220 177.575 20.695 177.815 ;
        RECT 20.865 177.565 21.240 177.815 ;
        RECT 20.865 177.395 21.035 177.565 ;
        RECT 17.475 176.425 17.655 177.185 ;
        RECT 17.835 176.255 18.165 177.015 ;
        RECT 18.335 176.425 18.605 177.330 ;
        RECT 19.700 177.225 21.035 177.395 ;
        RECT 19.700 177.065 19.980 177.225 ;
        RECT 21.410 177.055 21.780 178.345 ;
        RECT 22.000 177.965 22.260 178.805 ;
        RECT 22.435 178.060 22.690 178.635 ;
        RECT 22.860 178.425 23.190 178.805 ;
        RECT 23.405 178.255 23.575 178.635 ;
        RECT 22.860 178.085 23.575 178.255 ;
        RECT 23.835 178.130 24.095 178.635 ;
        RECT 24.275 178.425 24.605 178.805 ;
        RECT 24.785 178.255 24.955 178.635 ;
        RECT 20.190 176.255 20.440 177.055 ;
        RECT 20.610 176.885 21.780 177.055 ;
        RECT 20.610 176.425 20.940 176.885 ;
        RECT 21.110 176.255 21.325 176.715 ;
        RECT 22.000 176.255 22.260 177.405 ;
        RECT 22.435 177.330 22.605 178.060 ;
        RECT 22.860 177.895 23.030 178.085 ;
        RECT 22.775 177.565 23.030 177.895 ;
        RECT 22.860 177.355 23.030 177.565 ;
        RECT 23.310 177.535 23.665 177.905 ;
        RECT 22.435 176.425 22.690 177.330 ;
        RECT 22.860 177.185 23.575 177.355 ;
        RECT 22.860 176.255 23.190 177.015 ;
        RECT 23.405 176.425 23.575 177.185 ;
        RECT 23.835 177.330 24.005 178.130 ;
        RECT 24.290 178.085 24.955 178.255 ;
        RECT 25.305 178.255 25.475 178.635 ;
        RECT 25.655 178.425 25.985 178.805 ;
        RECT 25.305 178.085 25.970 178.255 ;
        RECT 26.165 178.130 26.425 178.635 ;
        RECT 24.290 177.830 24.460 178.085 ;
        RECT 24.175 177.500 24.460 177.830 ;
        RECT 24.695 177.535 25.025 177.905 ;
        RECT 25.235 177.535 25.565 177.905 ;
        RECT 25.800 177.830 25.970 178.085 ;
        RECT 24.290 177.355 24.460 177.500 ;
        RECT 25.800 177.500 26.085 177.830 ;
        RECT 25.800 177.355 25.970 177.500 ;
        RECT 23.835 176.425 24.105 177.330 ;
        RECT 24.290 177.185 24.955 177.355 ;
        RECT 24.275 176.255 24.605 177.015 ;
        RECT 24.785 176.425 24.955 177.185 ;
        RECT 25.305 177.185 25.970 177.355 ;
        RECT 26.255 177.330 26.425 178.130 ;
        RECT 26.595 178.035 30.105 178.805 ;
        RECT 26.595 177.515 28.245 178.035 ;
        RECT 31.195 178.005 31.505 178.805 ;
        RECT 31.710 178.005 32.405 178.635 ;
        RECT 32.575 178.260 37.920 178.805 ;
        RECT 31.710 177.955 31.885 178.005 ;
        RECT 28.415 177.345 30.105 177.865 ;
        RECT 31.205 177.565 31.540 177.835 ;
        RECT 31.710 177.405 31.880 177.955 ;
        RECT 32.050 177.565 32.385 177.815 ;
        RECT 34.160 177.430 34.500 178.260 ;
        RECT 38.095 178.035 41.605 178.805 ;
        RECT 41.775 178.080 42.065 178.805 ;
        RECT 42.320 178.305 42.815 178.635 ;
        RECT 25.305 176.425 25.475 177.185 ;
        RECT 25.655 176.255 25.985 177.015 ;
        RECT 26.155 176.425 26.425 177.330 ;
        RECT 26.595 176.255 30.105 177.345 ;
        RECT 31.195 176.255 31.475 177.395 ;
        RECT 31.645 176.425 31.975 177.405 ;
        RECT 32.145 176.255 32.405 177.395 ;
        RECT 35.980 176.690 36.330 177.940 ;
        RECT 38.095 177.515 39.745 178.035 ;
        RECT 39.915 177.345 41.605 177.865 ;
        RECT 32.575 176.255 37.920 176.690 ;
        RECT 38.095 176.255 41.605 177.345 ;
        RECT 41.775 176.255 42.065 177.420 ;
        RECT 42.235 176.815 42.475 178.125 ;
        RECT 42.645 177.395 42.815 178.305 ;
        RECT 43.035 177.565 43.385 178.530 ;
        RECT 43.565 177.565 43.865 178.535 ;
        RECT 44.045 177.565 44.325 178.535 ;
        RECT 44.505 178.005 44.775 178.805 ;
        RECT 44.945 178.085 45.285 178.595 ;
        RECT 45.480 178.415 45.810 178.805 ;
        RECT 45.980 178.245 46.205 178.625 ;
        RECT 44.520 177.565 44.850 177.815 ;
        RECT 44.520 177.395 44.835 177.565 ;
        RECT 42.645 177.225 44.835 177.395 ;
        RECT 42.240 176.255 42.575 176.635 ;
        RECT 42.745 176.425 42.995 177.225 ;
        RECT 43.215 176.255 43.545 176.975 ;
        RECT 43.730 176.425 43.980 177.225 ;
        RECT 44.445 176.255 44.775 177.055 ;
        RECT 45.025 176.685 45.285 178.085 ;
        RECT 45.465 177.565 45.705 178.215 ;
        RECT 45.875 178.065 46.205 178.245 ;
        RECT 45.875 177.395 46.050 178.065 ;
        RECT 46.405 177.895 46.635 178.515 ;
        RECT 46.815 178.075 47.115 178.805 ;
        RECT 47.755 178.005 48.450 178.635 ;
        RECT 48.655 178.005 48.965 178.805 ;
        RECT 49.135 178.130 49.395 178.635 ;
        RECT 49.575 178.425 49.905 178.805 ;
        RECT 50.085 178.255 50.255 178.635 ;
        RECT 46.220 177.565 46.635 177.895 ;
        RECT 46.815 177.565 47.110 177.895 ;
        RECT 47.775 177.565 48.110 177.815 ;
        RECT 48.280 177.405 48.450 178.005 ;
        RECT 48.620 177.565 48.955 177.835 ;
        RECT 44.945 176.425 45.285 176.685 ;
        RECT 45.465 177.205 46.050 177.395 ;
        RECT 45.465 176.435 45.740 177.205 ;
        RECT 46.220 177.035 47.115 177.365 ;
        RECT 45.910 176.865 47.115 177.035 ;
        RECT 45.910 176.435 46.240 176.865 ;
        RECT 46.410 176.255 46.605 176.695 ;
        RECT 46.785 176.435 47.115 176.865 ;
        RECT 47.755 176.255 48.015 177.395 ;
        RECT 48.185 176.425 48.515 177.405 ;
        RECT 48.685 176.255 48.965 177.395 ;
        RECT 49.135 177.330 49.305 178.130 ;
        RECT 49.590 178.085 50.255 178.255 ;
        RECT 50.515 178.130 50.775 178.635 ;
        RECT 50.955 178.425 51.285 178.805 ;
        RECT 51.465 178.255 51.635 178.635 ;
        RECT 49.590 177.830 49.760 178.085 ;
        RECT 49.475 177.500 49.760 177.830 ;
        RECT 49.995 177.535 50.325 177.905 ;
        RECT 49.590 177.355 49.760 177.500 ;
        RECT 49.135 176.425 49.405 177.330 ;
        RECT 49.590 177.185 50.255 177.355 ;
        RECT 49.575 176.255 49.905 177.015 ;
        RECT 50.085 176.425 50.255 177.185 ;
        RECT 50.515 177.330 50.695 178.130 ;
        RECT 50.970 178.085 51.635 178.255 ;
        RECT 50.970 177.830 51.140 178.085 ;
        RECT 51.895 178.005 52.590 178.635 ;
        RECT 52.795 178.005 53.105 178.805 ;
        RECT 53.275 178.130 53.535 178.635 ;
        RECT 53.715 178.425 54.045 178.805 ;
        RECT 54.225 178.255 54.395 178.635 ;
        RECT 50.865 177.500 51.140 177.830 ;
        RECT 51.365 177.535 51.705 177.905 ;
        RECT 51.915 177.565 52.250 177.815 ;
        RECT 50.970 177.355 51.140 177.500 ;
        RECT 52.420 177.445 52.590 178.005 ;
        RECT 52.760 177.565 53.095 177.835 ;
        RECT 52.415 177.405 52.590 177.445 ;
        RECT 50.515 176.425 50.785 177.330 ;
        RECT 50.970 177.185 51.645 177.355 ;
        RECT 50.955 176.255 51.285 177.015 ;
        RECT 51.465 176.425 51.645 177.185 ;
        RECT 51.895 176.255 52.155 177.395 ;
        RECT 52.325 176.425 52.655 177.405 ;
        RECT 52.825 176.255 53.105 177.395 ;
        RECT 53.275 177.330 53.455 178.130 ;
        RECT 53.730 178.085 54.395 178.255 ;
        RECT 53.730 177.830 53.900 178.085 ;
        RECT 53.625 177.500 53.900 177.830 ;
        RECT 54.125 177.535 54.465 177.905 ;
        RECT 53.730 177.355 53.900 177.500 ;
        RECT 53.275 176.425 53.545 177.330 ;
        RECT 53.730 177.185 54.405 177.355 ;
        RECT 53.715 176.255 54.045 177.015 ;
        RECT 54.225 176.425 54.405 177.185 ;
        RECT 54.670 176.435 54.950 178.625 ;
        RECT 55.150 178.435 55.880 178.805 ;
        RECT 56.460 178.265 56.890 178.625 ;
        RECT 55.150 178.075 56.890 178.265 ;
        RECT 55.150 177.565 55.410 178.075 ;
        RECT 55.140 176.255 55.425 177.395 ;
        RECT 55.620 177.275 55.880 177.895 ;
        RECT 56.075 177.275 56.500 177.895 ;
        RECT 56.670 177.845 56.890 178.075 ;
        RECT 57.060 178.025 57.305 178.805 ;
        RECT 56.670 177.545 57.215 177.845 ;
        RECT 57.505 177.725 57.735 178.625 ;
        RECT 55.690 176.905 56.715 177.105 ;
        RECT 55.690 176.435 55.860 176.905 ;
        RECT 56.035 176.255 56.365 176.735 ;
        RECT 56.535 176.435 56.715 176.905 ;
        RECT 56.885 176.435 57.215 177.545 ;
        RECT 57.395 177.045 57.735 177.725 ;
        RECT 57.915 177.225 58.145 178.565 ;
        RECT 58.335 178.005 59.030 178.635 ;
        RECT 59.235 178.005 59.545 178.805 ;
        RECT 59.725 178.295 60.175 178.805 ;
        RECT 60.450 178.385 61.755 178.635 ;
        RECT 61.935 178.405 62.265 178.805 ;
        RECT 61.575 178.235 61.755 178.385 ;
        RECT 58.355 177.565 58.690 177.815 ;
        RECT 58.860 177.405 59.030 178.005 ;
        RECT 59.200 177.565 59.535 177.835 ;
        RECT 59.755 177.615 60.205 178.125 ;
        RECT 60.620 177.815 60.870 178.215 ;
        RECT 60.395 177.615 60.870 177.815 ;
        RECT 61.120 177.815 61.330 178.215 ;
        RECT 61.575 178.065 62.305 178.235 ;
        RECT 61.120 177.615 61.470 177.815 ;
        RECT 61.640 177.565 61.965 177.895 ;
        RECT 57.395 176.845 58.145 177.045 ;
        RECT 57.385 176.255 57.735 176.665 ;
        RECT 57.905 176.455 58.145 176.845 ;
        RECT 58.335 176.255 58.595 177.395 ;
        RECT 58.765 176.425 59.095 177.405 ;
        RECT 59.725 177.395 61.470 177.445 ;
        RECT 62.135 177.395 62.305 178.065 ;
        RECT 59.265 176.255 59.545 177.395 ;
        RECT 59.725 177.265 62.305 177.395 ;
        RECT 59.725 176.595 60.055 177.265 ;
        RECT 61.245 177.225 62.305 177.265 ;
        RECT 62.935 178.080 63.195 178.635 ;
        RECT 63.365 178.360 63.795 178.805 ;
        RECT 64.030 178.235 64.200 178.635 ;
        RECT 64.370 178.405 65.090 178.805 ;
        RECT 62.935 177.365 63.110 178.080 ;
        RECT 64.030 178.065 64.910 178.235 ;
        RECT 65.260 178.190 65.430 178.635 ;
        RECT 66.005 178.295 66.405 178.805 ;
        RECT 63.280 177.565 63.535 177.895 ;
        RECT 60.225 177.055 61.105 177.095 ;
        RECT 60.225 176.855 61.755 177.055 ;
        RECT 60.225 176.805 60.840 176.855 ;
        RECT 60.225 176.765 60.455 176.805 ;
        RECT 61.585 176.725 61.755 176.855 ;
        RECT 60.565 176.595 60.895 176.635 ;
        RECT 59.725 176.425 60.895 176.595 ;
        RECT 61.065 176.255 61.440 176.635 ;
        RECT 61.990 176.255 62.255 177.035 ;
        RECT 62.935 176.425 63.195 177.365 ;
        RECT 63.365 177.085 63.535 177.565 ;
        RECT 63.760 177.275 64.090 177.895 ;
        RECT 64.260 177.515 64.550 177.895 ;
        RECT 64.740 177.345 64.910 178.065 ;
        RECT 64.390 177.175 64.910 177.345 ;
        RECT 65.080 178.020 65.430 178.190 ;
        RECT 63.365 176.915 64.125 177.085 ;
        RECT 64.390 176.985 64.560 177.175 ;
        RECT 65.080 176.995 65.250 178.020 ;
        RECT 65.670 177.535 65.930 178.125 ;
        RECT 65.450 177.235 65.930 177.535 ;
        RECT 66.130 177.235 66.390 178.125 ;
        RECT 67.535 178.080 67.825 178.805 ;
        RECT 67.995 178.305 68.255 178.635 ;
        RECT 68.425 178.445 68.755 178.805 ;
        RECT 69.010 178.425 70.310 178.635 ;
        RECT 63.955 176.690 64.125 176.915 ;
        RECT 64.840 176.825 65.250 176.995 ;
        RECT 65.425 176.885 66.365 177.055 ;
        RECT 64.840 176.690 65.095 176.825 ;
        RECT 63.365 176.255 63.695 176.655 ;
        RECT 63.955 176.520 65.095 176.690 ;
        RECT 65.425 176.635 65.595 176.885 ;
        RECT 64.840 176.425 65.095 176.520 ;
        RECT 65.265 176.465 65.595 176.635 ;
        RECT 65.765 176.255 66.015 176.715 ;
        RECT 66.185 176.425 66.365 176.885 ;
        RECT 67.535 176.255 67.825 177.420 ;
        RECT 67.995 177.105 68.165 178.305 ;
        RECT 69.010 178.275 69.180 178.425 ;
        RECT 68.425 178.150 69.180 178.275 ;
        RECT 68.335 178.105 69.180 178.150 ;
        RECT 68.335 177.985 68.605 178.105 ;
        RECT 68.335 177.410 68.505 177.985 ;
        RECT 68.735 177.545 69.145 177.850 ;
        RECT 69.435 177.815 69.645 178.215 ;
        RECT 69.315 177.605 69.645 177.815 ;
        RECT 69.890 177.815 70.110 178.215 ;
        RECT 70.585 178.040 71.040 178.805 ;
        RECT 71.700 178.050 71.935 178.380 ;
        RECT 72.105 178.065 72.435 178.805 ;
        RECT 72.670 178.425 73.865 178.635 ;
        RECT 69.890 177.605 70.365 177.815 ;
        RECT 70.555 177.615 71.045 177.815 ;
        RECT 68.335 177.375 68.535 177.410 ;
        RECT 69.865 177.375 71.040 177.435 ;
        RECT 68.335 177.265 71.040 177.375 ;
        RECT 68.395 177.205 70.195 177.265 ;
        RECT 69.865 177.175 70.195 177.205 ;
        RECT 67.995 176.425 68.255 177.105 ;
        RECT 68.425 176.255 68.675 177.035 ;
        RECT 68.925 177.005 69.760 177.015 ;
        RECT 70.350 177.005 70.535 177.095 ;
        RECT 68.925 176.805 70.535 177.005 ;
        RECT 68.925 176.425 69.175 176.805 ;
        RECT 70.305 176.765 70.535 176.805 ;
        RECT 70.785 176.645 71.040 177.265 ;
        RECT 71.700 177.395 71.870 178.050 ;
        RECT 72.670 177.985 72.945 178.425 ;
        RECT 73.115 178.085 73.445 178.255 ;
        RECT 73.120 177.985 73.445 178.085 ;
        RECT 73.615 178.195 73.865 178.425 ;
        RECT 74.035 178.365 74.205 178.805 ;
        RECT 74.375 178.195 74.725 178.635 ;
        RECT 75.815 178.295 76.120 178.805 ;
        RECT 73.615 177.985 74.725 178.195 ;
        RECT 72.045 177.565 72.390 177.895 ;
        RECT 72.620 177.395 72.950 177.815 ;
        RECT 71.700 177.225 72.950 177.395 ;
        RECT 71.700 177.030 72.000 177.225 ;
        RECT 73.120 177.055 73.400 177.985 ;
        RECT 73.580 177.615 74.725 177.815 ;
        RECT 73.580 177.445 73.770 177.615 ;
        RECT 75.815 177.565 76.130 178.125 ;
        RECT 76.300 177.815 76.550 178.625 ;
        RECT 76.720 178.280 76.980 178.805 ;
        RECT 77.160 177.815 77.410 178.625 ;
        RECT 77.580 178.245 77.840 178.805 ;
        RECT 78.010 178.155 78.270 178.610 ;
        RECT 78.440 178.325 78.700 178.805 ;
        RECT 78.870 178.155 79.130 178.610 ;
        RECT 79.300 178.325 79.560 178.805 ;
        RECT 79.730 178.155 79.990 178.610 ;
        RECT 80.160 178.325 80.405 178.805 ;
        RECT 80.575 178.155 80.850 178.610 ;
        RECT 81.020 178.325 81.265 178.805 ;
        RECT 81.435 178.155 81.695 178.610 ;
        RECT 81.875 178.325 82.125 178.805 ;
        RECT 82.295 178.155 82.555 178.610 ;
        RECT 82.735 178.325 82.985 178.805 ;
        RECT 83.155 178.155 83.415 178.610 ;
        RECT 83.595 178.325 83.855 178.805 ;
        RECT 84.025 178.155 84.285 178.610 ;
        RECT 84.455 178.325 84.755 178.805 ;
        RECT 78.010 177.985 84.755 178.155 ;
        RECT 85.935 178.055 87.145 178.805 ;
        RECT 76.300 177.565 83.420 177.815 ;
        RECT 73.575 177.275 73.770 177.445 ;
        RECT 74.035 177.395 74.205 177.445 ;
        RECT 73.580 177.235 73.770 177.275 ;
        RECT 73.950 177.055 74.225 177.395 ;
        RECT 69.345 176.255 69.700 176.635 ;
        RECT 70.705 176.425 71.040 176.645 ;
        RECT 72.170 176.255 72.425 177.055 ;
        RECT 72.625 176.885 74.225 177.055 ;
        RECT 72.625 176.425 72.955 176.885 ;
        RECT 73.125 176.255 73.700 176.715 ;
        RECT 73.870 176.425 74.225 176.885 ;
        RECT 74.395 176.255 74.725 177.395 ;
        RECT 75.825 176.255 76.120 177.065 ;
        RECT 76.300 176.425 76.545 177.565 ;
        RECT 76.720 176.255 76.980 177.065 ;
        RECT 77.160 176.430 77.410 177.565 ;
        RECT 83.590 177.395 84.755 177.985 ;
        RECT 78.010 177.170 84.755 177.395 ;
        RECT 85.935 177.345 86.455 177.885 ;
        RECT 86.625 177.515 87.145 178.055 ;
        RECT 78.010 177.155 83.415 177.170 ;
        RECT 77.580 176.260 77.840 177.055 ;
        RECT 78.010 176.430 78.270 177.155 ;
        RECT 78.440 176.260 78.700 176.985 ;
        RECT 78.870 176.430 79.130 177.155 ;
        RECT 79.300 176.260 79.560 176.985 ;
        RECT 79.730 176.430 79.990 177.155 ;
        RECT 80.160 176.260 80.420 176.985 ;
        RECT 80.590 176.430 80.850 177.155 ;
        RECT 81.020 176.260 81.265 176.985 ;
        RECT 81.435 176.430 81.695 177.155 ;
        RECT 81.880 176.260 82.125 176.985 ;
        RECT 82.295 176.430 82.555 177.155 ;
        RECT 82.740 176.260 82.985 176.985 ;
        RECT 83.155 176.430 83.415 177.155 ;
        RECT 83.600 176.260 83.855 176.985 ;
        RECT 84.025 176.430 84.315 177.170 ;
        RECT 77.580 176.255 83.855 176.260 ;
        RECT 84.485 176.255 84.755 177.000 ;
        RECT 85.935 176.255 87.145 177.345 ;
        RECT 15.930 176.085 87.230 176.255 ;
        RECT 16.015 174.995 17.225 176.085 ;
        RECT 16.015 174.285 16.535 174.825 ;
        RECT 16.705 174.455 17.225 174.995 ;
        RECT 16.015 173.535 17.225 174.285 ;
        RECT 18.315 173.815 18.595 175.915 ;
        RECT 18.785 175.325 19.570 176.085 ;
        RECT 19.965 175.255 20.350 175.915 ;
        RECT 19.965 175.155 20.375 175.255 ;
        RECT 18.765 174.945 20.375 175.155 ;
        RECT 20.675 175.065 20.875 175.855 ;
        RECT 18.765 174.345 19.040 174.945 ;
        RECT 20.545 174.895 20.875 175.065 ;
        RECT 21.045 174.905 21.365 176.085 ;
        RECT 21.535 175.650 26.880 176.085 ;
        RECT 20.545 174.775 20.725 174.895 ;
        RECT 19.210 174.525 19.565 174.775 ;
        RECT 19.760 174.725 20.225 174.775 ;
        RECT 19.755 174.555 20.225 174.725 ;
        RECT 19.760 174.525 20.225 174.555 ;
        RECT 20.395 174.525 20.725 174.775 ;
        RECT 20.900 174.525 21.365 174.725 ;
        RECT 18.765 174.165 20.015 174.345 ;
        RECT 19.650 174.095 20.015 174.165 ;
        RECT 20.185 174.145 21.365 174.315 ;
        RECT 18.825 173.535 18.995 173.995 ;
        RECT 20.185 173.925 20.515 174.145 ;
        RECT 19.265 173.745 20.515 173.925 ;
        RECT 20.685 173.535 20.855 173.975 ;
        RECT 21.025 173.730 21.365 174.145 ;
        RECT 23.120 174.080 23.460 174.910 ;
        RECT 24.940 174.400 25.290 175.650 ;
        RECT 27.055 174.995 28.725 176.085 ;
        RECT 27.055 174.305 27.805 174.825 ;
        RECT 27.975 174.475 28.725 174.995 ;
        RECT 28.895 174.920 29.185 176.085 ;
        RECT 29.375 175.195 29.635 175.905 ;
        RECT 29.805 175.375 30.135 176.085 ;
        RECT 30.305 175.195 30.535 175.905 ;
        RECT 29.375 174.955 30.535 175.195 ;
        RECT 30.715 175.175 30.985 175.905 ;
        RECT 31.165 175.355 31.505 176.085 ;
        RECT 30.715 174.955 31.485 175.175 ;
        RECT 29.365 174.445 29.665 174.775 ;
        RECT 29.845 174.465 30.370 174.775 ;
        RECT 30.550 174.465 31.015 174.775 ;
        RECT 21.535 173.535 26.880 174.080 ;
        RECT 27.055 173.535 28.725 174.305 ;
        RECT 28.895 173.535 29.185 174.260 ;
        RECT 29.375 173.535 29.665 174.265 ;
        RECT 29.845 173.825 30.075 174.465 ;
        RECT 31.195 174.285 31.485 174.955 ;
        RECT 30.255 174.085 31.485 174.285 ;
        RECT 30.255 173.715 30.565 174.085 ;
        RECT 30.745 173.535 31.415 173.905 ;
        RECT 31.675 173.715 31.935 175.905 ;
        RECT 32.115 174.995 35.625 176.085 ;
        RECT 32.115 174.305 33.765 174.825 ;
        RECT 33.935 174.475 35.625 174.995 ;
        RECT 36.255 174.945 36.515 176.085 ;
        RECT 36.685 174.935 37.015 175.915 ;
        RECT 37.185 174.945 37.465 176.085 ;
        RECT 37.635 175.650 42.980 176.085 ;
        RECT 43.155 175.650 48.500 176.085 ;
        RECT 36.275 174.525 36.610 174.775 ;
        RECT 36.780 174.335 36.950 174.935 ;
        RECT 37.120 174.505 37.455 174.775 ;
        RECT 32.115 173.535 35.625 174.305 ;
        RECT 36.255 173.705 36.950 174.335 ;
        RECT 37.155 173.535 37.465 174.335 ;
        RECT 39.220 174.080 39.560 174.910 ;
        RECT 41.040 174.400 41.390 175.650 ;
        RECT 44.740 174.080 45.080 174.910 ;
        RECT 46.560 174.400 46.910 175.650 ;
        RECT 49.605 175.135 49.880 175.905 ;
        RECT 50.050 175.475 50.380 175.905 ;
        RECT 50.550 175.645 50.745 176.085 ;
        RECT 50.925 175.475 51.255 175.905 ;
        RECT 50.050 175.305 51.255 175.475 ;
        RECT 49.605 174.945 50.190 175.135 ;
        RECT 50.360 174.975 51.255 175.305 ;
        RECT 52.365 175.135 52.640 175.905 ;
        RECT 52.810 175.475 53.140 175.905 ;
        RECT 53.310 175.645 53.505 176.085 ;
        RECT 53.685 175.475 54.015 175.905 ;
        RECT 52.810 175.305 54.015 175.475 ;
        RECT 52.365 174.945 52.950 175.135 ;
        RECT 53.120 174.975 54.015 175.305 ;
        RECT 49.605 174.125 49.845 174.775 ;
        RECT 50.015 174.275 50.190 174.945 ;
        RECT 50.360 174.445 50.775 174.775 ;
        RECT 50.955 174.445 51.250 174.775 ;
        RECT 50.015 174.095 50.345 174.275 ;
        RECT 37.635 173.535 42.980 174.080 ;
        RECT 43.155 173.535 48.500 174.080 ;
        RECT 49.620 173.535 49.950 173.925 ;
        RECT 50.120 173.715 50.345 174.095 ;
        RECT 50.545 173.825 50.775 174.445 ;
        RECT 50.955 173.535 51.255 174.265 ;
        RECT 52.365 174.125 52.605 174.775 ;
        RECT 52.775 174.275 52.950 174.945 ;
        RECT 54.655 174.920 54.945 176.085 ;
        RECT 55.575 175.010 55.845 175.915 ;
        RECT 56.015 175.325 56.345 176.085 ;
        RECT 56.525 175.155 56.705 175.915 ;
        RECT 53.120 174.445 53.535 174.775 ;
        RECT 53.715 174.445 54.010 174.775 ;
        RECT 52.775 174.095 53.105 174.275 ;
        RECT 52.380 173.535 52.710 173.925 ;
        RECT 52.880 173.715 53.105 174.095 ;
        RECT 53.305 173.825 53.535 174.445 ;
        RECT 53.715 173.535 54.015 174.265 ;
        RECT 54.655 173.535 54.945 174.260 ;
        RECT 55.575 174.210 55.755 175.010 ;
        RECT 56.030 174.985 56.705 175.155 ;
        RECT 56.030 174.840 56.200 174.985 ;
        RECT 56.995 174.945 57.225 176.085 ;
        RECT 57.395 174.935 57.725 175.915 ;
        RECT 57.895 174.945 58.105 176.085 ;
        RECT 58.335 174.945 58.615 176.085 ;
        RECT 58.785 174.935 59.115 175.915 ;
        RECT 59.285 174.945 59.545 176.085 ;
        RECT 59.715 175.235 59.975 175.915 ;
        RECT 60.145 175.305 60.395 176.085 ;
        RECT 60.645 175.535 60.895 175.915 ;
        RECT 61.065 175.705 61.420 176.085 ;
        RECT 62.425 175.695 62.760 175.915 ;
        RECT 62.025 175.535 62.255 175.575 ;
        RECT 60.645 175.335 62.255 175.535 ;
        RECT 60.645 175.325 61.480 175.335 ;
        RECT 62.070 175.245 62.255 175.335 ;
        RECT 55.925 174.510 56.200 174.840 ;
        RECT 56.030 174.255 56.200 174.510 ;
        RECT 56.425 174.435 56.765 174.805 ;
        RECT 56.975 174.525 57.305 174.775 ;
        RECT 55.575 173.705 55.835 174.210 ;
        RECT 56.030 174.085 56.695 174.255 ;
        RECT 56.015 173.535 56.345 173.915 ;
        RECT 56.525 173.705 56.695 174.085 ;
        RECT 56.995 173.535 57.225 174.355 ;
        RECT 57.475 174.335 57.725 174.935 ;
        RECT 58.345 174.505 58.680 174.775 ;
        RECT 57.395 173.705 57.725 174.335 ;
        RECT 57.895 173.535 58.105 174.355 ;
        RECT 58.850 174.335 59.020 174.935 ;
        RECT 59.190 174.525 59.525 174.775 ;
        RECT 58.335 173.535 58.645 174.335 ;
        RECT 58.850 173.705 59.545 174.335 ;
        RECT 59.715 174.035 59.885 175.235 ;
        RECT 61.585 175.135 61.915 175.165 ;
        RECT 60.115 175.075 61.915 175.135 ;
        RECT 62.505 175.075 62.760 175.695 ;
        RECT 60.055 174.965 62.760 175.075 ;
        RECT 60.055 174.930 60.255 174.965 ;
        RECT 60.055 174.355 60.225 174.930 ;
        RECT 61.585 174.905 62.760 174.965 ;
        RECT 63.395 175.010 63.665 175.915 ;
        RECT 63.835 175.325 64.165 176.085 ;
        RECT 64.345 175.155 64.525 175.915 ;
        RECT 60.455 174.490 60.865 174.795 ;
        RECT 61.035 174.525 61.365 174.735 ;
        RECT 60.055 174.235 60.325 174.355 ;
        RECT 60.055 174.190 60.900 174.235 ;
        RECT 60.145 174.065 60.900 174.190 ;
        RECT 61.155 174.125 61.365 174.525 ;
        RECT 61.610 174.525 62.085 174.735 ;
        RECT 62.275 174.525 62.765 174.725 ;
        RECT 61.610 174.125 61.830 174.525 ;
        RECT 59.715 173.705 59.975 174.035 ;
        RECT 60.730 173.915 60.900 174.065 ;
        RECT 60.145 173.535 60.475 173.895 ;
        RECT 60.730 173.705 62.030 173.915 ;
        RECT 62.305 173.535 62.760 174.300 ;
        RECT 63.395 174.210 63.575 175.010 ;
        RECT 63.850 174.985 64.525 175.155 ;
        RECT 63.850 174.840 64.020 174.985 ;
        RECT 64.785 174.945 65.115 176.085 ;
        RECT 65.645 175.115 65.975 175.900 ;
        RECT 65.295 174.945 65.975 175.115 ;
        RECT 66.195 174.945 66.425 176.085 ;
        RECT 63.745 174.510 64.020 174.840 ;
        RECT 63.850 174.255 64.020 174.510 ;
        RECT 64.245 174.435 64.585 174.805 ;
        RECT 64.775 174.525 65.125 174.775 ;
        RECT 65.295 174.345 65.465 174.945 ;
        RECT 66.595 174.935 66.925 175.915 ;
        RECT 67.095 174.945 67.305 176.085 ;
        RECT 67.640 175.285 67.895 176.085 ;
        RECT 68.065 175.115 68.395 175.915 ;
        RECT 68.565 175.285 68.735 176.085 ;
        RECT 68.905 175.115 69.235 175.915 ;
        RECT 67.535 174.945 69.235 175.115 ;
        RECT 69.405 174.945 69.665 176.085 ;
        RECT 70.040 175.645 70.370 176.085 ;
        RECT 70.540 175.475 70.775 175.915 ;
        RECT 70.960 175.705 71.290 176.085 ;
        RECT 71.500 175.475 71.845 175.915 ;
        RECT 69.835 175.235 71.845 175.475 ;
        RECT 65.635 174.525 65.985 174.775 ;
        RECT 66.175 174.525 66.505 174.775 ;
        RECT 63.395 173.705 63.655 174.210 ;
        RECT 63.850 174.085 64.515 174.255 ;
        RECT 63.835 173.535 64.165 173.915 ;
        RECT 64.345 173.705 64.515 174.085 ;
        RECT 64.785 173.535 65.055 174.345 ;
        RECT 65.225 173.705 65.555 174.345 ;
        RECT 65.725 173.535 65.965 174.345 ;
        RECT 66.195 173.535 66.425 174.355 ;
        RECT 66.675 174.335 66.925 174.935 ;
        RECT 67.535 174.355 67.815 174.945 ;
        RECT 67.985 174.525 68.735 174.775 ;
        RECT 68.905 174.525 69.665 174.775 ;
        RECT 66.595 173.705 66.925 174.335 ;
        RECT 67.095 173.535 67.305 174.355 ;
        RECT 67.535 174.105 68.395 174.355 ;
        RECT 69.835 174.335 70.065 175.235 ;
        RECT 72.020 175.065 72.365 175.820 ;
        RECT 72.535 175.245 72.865 176.085 ;
        RECT 73.075 175.245 73.405 176.085 ;
        RECT 73.575 175.065 73.920 175.820 ;
        RECT 74.095 175.475 74.440 175.915 ;
        RECT 74.650 175.705 74.980 176.085 ;
        RECT 75.165 175.475 75.400 175.915 ;
        RECT 75.570 175.645 75.900 176.085 ;
        RECT 74.095 175.235 76.105 175.475 ;
        RECT 70.235 174.525 70.565 175.065 ;
        RECT 68.565 174.165 69.665 174.335 ;
        RECT 67.645 173.915 67.975 173.935 ;
        RECT 68.565 173.915 68.815 174.165 ;
        RECT 67.645 173.705 68.815 173.915 ;
        RECT 68.985 173.535 69.155 173.995 ;
        RECT 69.325 173.705 69.665 174.165 ;
        RECT 69.835 173.705 70.440 174.335 ;
        RECT 70.775 173.705 71.105 175.065 ;
        RECT 71.275 174.445 71.565 175.065 ;
        RECT 71.735 174.445 72.365 175.065 ;
        RECT 72.535 174.455 72.865 175.065 ;
        RECT 73.075 174.455 73.405 175.065 ;
        RECT 73.575 174.445 74.205 175.065 ;
        RECT 74.375 174.445 74.665 175.065 ;
        RECT 71.500 174.075 72.865 174.275 ;
        RECT 71.500 173.705 71.845 174.075 ;
        RECT 72.035 173.535 72.365 173.905 ;
        RECT 72.535 173.705 72.865 174.075 ;
        RECT 73.075 174.075 74.440 174.275 ;
        RECT 73.075 173.705 73.405 174.075 ;
        RECT 73.575 173.535 73.905 173.905 ;
        RECT 74.095 173.705 74.440 174.075 ;
        RECT 74.835 173.705 75.165 175.065 ;
        RECT 75.375 174.525 75.705 175.065 ;
        RECT 75.875 174.335 76.105 175.235 ;
        RECT 76.735 174.945 77.065 176.085 ;
        RECT 77.235 175.455 77.590 175.915 ;
        RECT 77.760 175.625 78.335 176.085 ;
        RECT 78.505 175.455 78.835 175.915 ;
        RECT 77.235 175.285 78.835 175.455 ;
        RECT 79.035 175.285 79.290 176.085 ;
        RECT 77.235 174.945 77.510 175.285 ;
        RECT 77.690 174.725 77.880 175.105 ;
        RECT 76.735 174.525 77.880 174.725 ;
        RECT 78.060 174.355 78.340 175.285 ;
        RECT 79.460 175.115 79.760 175.310 ;
        RECT 78.510 174.945 79.760 175.115 ;
        RECT 78.510 174.525 78.840 174.945 ;
        RECT 79.070 174.445 79.415 174.775 ;
        RECT 75.500 173.705 76.105 174.335 ;
        RECT 76.735 174.145 77.845 174.355 ;
        RECT 76.735 173.705 77.085 174.145 ;
        RECT 77.255 173.535 77.425 173.975 ;
        RECT 77.595 173.915 77.845 174.145 ;
        RECT 78.015 174.255 78.340 174.355 ;
        RECT 78.015 174.085 78.345 174.255 ;
        RECT 78.515 173.915 78.790 174.355 ;
        RECT 79.590 174.290 79.760 174.945 ;
        RECT 80.415 174.920 80.705 176.085 ;
        RECT 80.875 174.945 81.205 176.085 ;
        RECT 81.375 175.455 81.730 175.915 ;
        RECT 81.900 175.625 82.475 176.085 ;
        RECT 82.645 175.455 82.975 175.915 ;
        RECT 81.375 175.285 82.975 175.455 ;
        RECT 83.175 175.285 83.430 176.085 ;
        RECT 81.375 174.945 81.650 175.285 ;
        RECT 81.830 174.725 82.020 175.105 ;
        RECT 80.875 174.555 82.025 174.725 ;
        RECT 80.875 174.525 82.020 174.555 ;
        RECT 82.200 174.355 82.480 175.285 ;
        RECT 83.600 175.115 83.900 175.310 ;
        RECT 82.650 174.945 83.900 175.115 ;
        RECT 84.185 175.155 84.355 175.915 ;
        RECT 84.570 175.325 84.900 176.085 ;
        RECT 84.185 174.985 84.900 175.155 ;
        RECT 85.070 175.010 85.325 175.915 ;
        RECT 82.650 174.525 82.980 174.945 ;
        RECT 83.210 174.445 83.555 174.775 ;
        RECT 77.595 173.705 78.790 173.915 ;
        RECT 79.025 173.535 79.355 174.275 ;
        RECT 79.525 173.960 79.760 174.290 ;
        RECT 80.415 173.535 80.705 174.260 ;
        RECT 80.875 174.145 81.985 174.355 ;
        RECT 80.875 173.705 81.225 174.145 ;
        RECT 81.395 173.535 81.565 173.975 ;
        RECT 81.735 173.915 81.985 174.145 ;
        RECT 82.155 174.255 82.480 174.355 ;
        RECT 82.155 174.085 82.485 174.255 ;
        RECT 82.655 173.915 82.930 174.355 ;
        RECT 83.730 174.290 83.900 174.945 ;
        RECT 84.095 174.435 84.450 174.805 ;
        RECT 84.730 174.775 84.900 174.985 ;
        RECT 84.730 174.445 84.985 174.775 ;
        RECT 81.735 173.705 82.930 173.915 ;
        RECT 83.165 173.535 83.495 174.275 ;
        RECT 83.665 173.960 83.900 174.290 ;
        RECT 84.730 174.255 84.900 174.445 ;
        RECT 85.155 174.280 85.325 175.010 ;
        RECT 85.500 174.935 85.760 176.085 ;
        RECT 85.935 174.995 87.145 176.085 ;
        RECT 85.935 174.455 86.455 174.995 ;
        RECT 84.185 174.085 84.900 174.255 ;
        RECT 84.185 173.705 84.355 174.085 ;
        RECT 84.570 173.535 84.900 173.915 ;
        RECT 85.070 173.705 85.325 174.280 ;
        RECT 85.500 173.535 85.760 174.375 ;
        RECT 86.625 174.285 87.145 174.825 ;
        RECT 85.935 173.535 87.145 174.285 ;
        RECT 15.930 173.365 87.230 173.535 ;
        RECT 16.015 172.615 17.225 173.365 ;
        RECT 16.015 172.075 16.535 172.615 ;
        RECT 17.395 172.595 19.065 173.365 ;
        RECT 19.700 172.625 19.955 173.195 ;
        RECT 20.125 172.965 20.455 173.365 ;
        RECT 20.880 172.830 21.410 173.195 ;
        RECT 21.600 173.025 21.875 173.195 ;
        RECT 21.595 172.855 21.875 173.025 ;
        RECT 20.880 172.795 21.055 172.830 ;
        RECT 20.125 172.625 21.055 172.795 ;
        RECT 16.705 171.905 17.225 172.445 ;
        RECT 17.395 172.075 18.145 172.595 ;
        RECT 18.315 171.905 19.065 172.425 ;
        RECT 16.015 170.815 17.225 171.905 ;
        RECT 17.395 170.815 19.065 171.905 ;
        RECT 19.700 171.955 19.870 172.625 ;
        RECT 20.125 172.455 20.295 172.625 ;
        RECT 20.040 172.125 20.295 172.455 ;
        RECT 20.520 172.125 20.715 172.455 ;
        RECT 19.700 170.985 20.035 171.955 ;
        RECT 20.205 170.815 20.375 171.955 ;
        RECT 20.545 171.155 20.715 172.125 ;
        RECT 20.885 171.495 21.055 172.625 ;
        RECT 21.225 171.835 21.395 172.635 ;
        RECT 21.600 172.035 21.875 172.855 ;
        RECT 22.045 171.835 22.235 173.195 ;
        RECT 22.415 172.830 22.925 173.365 ;
        RECT 23.145 172.555 23.390 173.160 ;
        RECT 23.835 172.595 26.425 173.365 ;
        RECT 26.605 172.635 26.905 173.365 ;
        RECT 22.435 172.385 23.665 172.555 ;
        RECT 21.225 171.665 22.235 171.835 ;
        RECT 22.405 171.820 23.155 172.010 ;
        RECT 20.885 171.325 22.010 171.495 ;
        RECT 22.405 171.155 22.575 171.820 ;
        RECT 23.325 171.575 23.665 172.385 ;
        RECT 23.835 172.075 25.045 172.595 ;
        RECT 27.085 172.455 27.315 173.075 ;
        RECT 27.515 172.805 27.740 173.185 ;
        RECT 27.910 172.975 28.240 173.365 ;
        RECT 27.515 172.625 27.845 172.805 ;
        RECT 25.215 171.905 26.425 172.425 ;
        RECT 26.610 172.125 26.905 172.455 ;
        RECT 27.085 172.125 27.500 172.455 ;
        RECT 27.670 171.955 27.845 172.625 ;
        RECT 28.015 172.125 28.255 172.775 ;
        RECT 28.470 172.625 29.085 173.195 ;
        RECT 29.255 172.855 29.470 173.365 ;
        RECT 29.700 172.855 29.980 173.185 ;
        RECT 30.160 172.855 30.400 173.365 ;
        RECT 20.545 170.985 22.575 171.155 ;
        RECT 22.745 170.815 22.915 171.575 ;
        RECT 23.150 171.165 23.665 171.575 ;
        RECT 23.835 170.815 26.425 171.905 ;
        RECT 26.605 171.595 27.500 171.925 ;
        RECT 27.670 171.765 28.255 171.955 ;
        RECT 26.605 171.425 27.810 171.595 ;
        RECT 26.605 170.995 26.935 171.425 ;
        RECT 27.115 170.815 27.310 171.255 ;
        RECT 27.480 170.995 27.810 171.425 ;
        RECT 27.980 170.995 28.255 171.765 ;
        RECT 28.470 171.605 28.785 172.625 ;
        RECT 28.955 171.955 29.125 172.455 ;
        RECT 29.375 172.125 29.640 172.685 ;
        RECT 29.810 171.955 29.980 172.855 ;
        RECT 30.735 172.755 31.075 173.170 ;
        RECT 31.245 172.925 31.415 173.365 ;
        RECT 31.585 172.975 32.835 173.155 ;
        RECT 31.585 172.755 31.915 172.975 ;
        RECT 33.105 172.905 33.275 173.365 ;
        RECT 30.150 172.125 30.505 172.685 ;
        RECT 30.735 172.585 31.915 172.755 ;
        RECT 32.085 172.735 32.450 172.805 ;
        RECT 32.085 172.555 33.335 172.735 ;
        RECT 30.735 172.175 31.200 172.375 ;
        RECT 31.375 172.125 31.705 172.375 ;
        RECT 31.875 172.345 32.340 172.375 ;
        RECT 31.875 172.175 32.345 172.345 ;
        RECT 31.875 172.125 32.340 172.175 ;
        RECT 32.535 172.125 32.890 172.375 ;
        RECT 31.375 172.005 31.555 172.125 ;
        RECT 28.955 171.785 30.380 171.955 ;
        RECT 28.470 170.985 29.005 171.605 ;
        RECT 29.175 170.815 29.505 171.615 ;
        RECT 29.990 171.610 30.380 171.785 ;
        RECT 30.735 170.815 31.055 171.995 ;
        RECT 31.225 171.835 31.555 172.005 ;
        RECT 33.060 171.955 33.335 172.555 ;
        RECT 31.225 171.045 31.425 171.835 ;
        RECT 31.725 171.745 33.335 171.955 ;
        RECT 31.725 171.645 32.135 171.745 ;
        RECT 31.750 170.985 32.135 171.645 ;
        RECT 32.530 170.815 33.315 171.575 ;
        RECT 33.505 170.985 33.785 173.085 ;
        RECT 34.880 172.625 35.135 173.195 ;
        RECT 35.305 172.965 35.635 173.365 ;
        RECT 36.060 172.830 36.590 173.195 ;
        RECT 36.060 172.795 36.235 172.830 ;
        RECT 35.305 172.625 36.235 172.795 ;
        RECT 34.880 171.955 35.050 172.625 ;
        RECT 35.305 172.455 35.475 172.625 ;
        RECT 35.220 172.125 35.475 172.455 ;
        RECT 35.700 172.125 35.895 172.455 ;
        RECT 34.880 170.985 35.215 171.955 ;
        RECT 35.385 170.815 35.555 171.955 ;
        RECT 35.725 171.155 35.895 172.125 ;
        RECT 36.065 171.495 36.235 172.625 ;
        RECT 36.405 171.835 36.575 172.635 ;
        RECT 36.780 172.345 37.055 173.195 ;
        RECT 36.775 172.175 37.055 172.345 ;
        RECT 36.780 172.035 37.055 172.175 ;
        RECT 37.225 171.835 37.415 173.195 ;
        RECT 37.595 172.830 38.105 173.365 ;
        RECT 38.325 172.555 38.570 173.160 ;
        RECT 39.015 172.595 41.605 173.365 ;
        RECT 41.775 172.640 42.065 173.365 ;
        RECT 42.245 172.635 42.545 173.365 ;
        RECT 37.615 172.385 38.845 172.555 ;
        RECT 36.405 171.665 37.415 171.835 ;
        RECT 37.585 171.820 38.335 172.010 ;
        RECT 36.065 171.325 37.190 171.495 ;
        RECT 37.585 171.155 37.755 171.820 ;
        RECT 38.505 171.575 38.845 172.385 ;
        RECT 39.015 172.075 40.225 172.595 ;
        RECT 42.725 172.455 42.955 173.075 ;
        RECT 43.155 172.805 43.380 173.185 ;
        RECT 43.550 172.975 43.880 173.365 ;
        RECT 43.155 172.625 43.485 172.805 ;
        RECT 40.395 171.905 41.605 172.425 ;
        RECT 42.250 172.125 42.545 172.455 ;
        RECT 42.725 172.125 43.140 172.455 ;
        RECT 35.725 170.985 37.755 171.155 ;
        RECT 37.925 170.815 38.095 171.575 ;
        RECT 38.330 171.165 38.845 171.575 ;
        RECT 39.015 170.815 41.605 171.905 ;
        RECT 41.775 170.815 42.065 171.980 ;
        RECT 43.310 171.955 43.485 172.625 ;
        RECT 43.655 172.125 43.895 172.775 ;
        RECT 42.245 171.595 43.140 171.925 ;
        RECT 43.310 171.765 43.895 171.955 ;
        RECT 42.245 171.425 43.450 171.595 ;
        RECT 42.245 170.995 42.575 171.425 ;
        RECT 42.755 170.815 42.950 171.255 ;
        RECT 43.120 170.995 43.450 171.425 ;
        RECT 43.620 170.995 43.895 171.765 ;
        RECT 44.545 170.995 44.805 173.185 ;
        RECT 45.065 172.995 45.735 173.365 ;
        RECT 45.915 172.815 46.225 173.185 ;
        RECT 44.995 172.615 46.225 172.815 ;
        RECT 44.995 171.945 45.285 172.615 ;
        RECT 46.405 172.435 46.635 173.075 ;
        RECT 46.815 172.635 47.105 173.365 ;
        RECT 47.295 172.595 49.885 173.365 ;
        RECT 50.080 172.975 50.410 173.365 ;
        RECT 50.580 172.805 50.805 173.185 ;
        RECT 45.465 172.125 45.930 172.435 ;
        RECT 46.110 172.125 46.635 172.435 ;
        RECT 46.815 172.125 47.115 172.455 ;
        RECT 47.295 172.075 48.505 172.595 ;
        RECT 44.995 171.725 45.765 171.945 ;
        RECT 44.975 170.815 45.315 171.545 ;
        RECT 45.495 170.995 45.765 171.725 ;
        RECT 45.945 171.705 47.105 171.945 ;
        RECT 48.675 171.905 49.885 172.425 ;
        RECT 50.065 172.125 50.305 172.775 ;
        RECT 50.475 172.625 50.805 172.805 ;
        RECT 50.475 171.955 50.650 172.625 ;
        RECT 51.005 172.455 51.235 173.075 ;
        RECT 51.415 172.635 51.715 173.365 ;
        RECT 52.840 172.975 53.170 173.365 ;
        RECT 53.340 172.805 53.565 173.185 ;
        RECT 50.820 172.125 51.235 172.455 ;
        RECT 51.415 172.125 51.710 172.455 ;
        RECT 52.825 172.125 53.065 172.775 ;
        RECT 53.235 172.625 53.565 172.805 ;
        RECT 53.235 171.955 53.410 172.625 ;
        RECT 53.765 172.455 53.995 173.075 ;
        RECT 54.175 172.635 54.475 173.365 ;
        RECT 55.575 172.690 55.835 173.195 ;
        RECT 56.015 172.985 56.345 173.365 ;
        RECT 56.525 172.815 56.695 173.195 ;
        RECT 53.580 172.125 53.995 172.455 ;
        RECT 54.175 172.125 54.470 172.455 ;
        RECT 45.945 170.995 46.175 171.705 ;
        RECT 46.345 170.815 46.675 171.525 ;
        RECT 46.845 170.995 47.105 171.705 ;
        RECT 47.295 170.815 49.885 171.905 ;
        RECT 50.065 171.765 50.650 171.955 ;
        RECT 50.065 170.995 50.340 171.765 ;
        RECT 50.820 171.595 51.715 171.925 ;
        RECT 50.510 171.425 51.715 171.595 ;
        RECT 50.510 170.995 50.840 171.425 ;
        RECT 51.010 170.815 51.205 171.255 ;
        RECT 51.385 170.995 51.715 171.425 ;
        RECT 52.825 171.765 53.410 171.955 ;
        RECT 52.825 170.995 53.100 171.765 ;
        RECT 53.580 171.595 54.475 171.925 ;
        RECT 53.270 171.425 54.475 171.595 ;
        RECT 53.270 170.995 53.600 171.425 ;
        RECT 53.770 170.815 53.965 171.255 ;
        RECT 54.145 170.995 54.475 171.425 ;
        RECT 55.575 171.890 55.755 172.690 ;
        RECT 56.030 172.645 56.695 172.815 ;
        RECT 56.030 172.390 56.200 172.645 ;
        RECT 55.925 172.060 56.200 172.390 ;
        RECT 56.425 172.095 56.765 172.465 ;
        RECT 56.030 171.915 56.200 172.060 ;
        RECT 55.575 170.985 55.845 171.890 ;
        RECT 56.030 171.745 56.705 171.915 ;
        RECT 56.015 170.815 56.345 171.575 ;
        RECT 56.525 170.985 56.705 171.745 ;
        RECT 56.970 170.995 57.250 173.185 ;
        RECT 57.450 172.995 58.180 173.365 ;
        RECT 58.760 172.825 59.190 173.185 ;
        RECT 57.450 172.635 59.190 172.825 ;
        RECT 57.450 172.125 57.710 172.635 ;
        RECT 57.440 170.815 57.725 171.955 ;
        RECT 57.920 171.835 58.180 172.455 ;
        RECT 58.375 171.835 58.800 172.455 ;
        RECT 58.970 172.405 59.190 172.635 ;
        RECT 59.360 172.585 59.605 173.365 ;
        RECT 58.970 172.105 59.515 172.405 ;
        RECT 59.805 172.285 60.035 173.185 ;
        RECT 57.990 171.465 59.015 171.665 ;
        RECT 57.990 170.995 58.160 171.465 ;
        RECT 58.335 170.815 58.665 171.295 ;
        RECT 58.835 170.995 59.015 171.465 ;
        RECT 59.185 170.995 59.515 172.105 ;
        RECT 59.695 171.605 60.035 172.285 ;
        RECT 60.215 171.785 60.445 173.125 ;
        RECT 60.725 172.815 60.895 173.195 ;
        RECT 61.075 172.985 61.405 173.365 ;
        RECT 60.725 172.645 61.390 172.815 ;
        RECT 61.585 172.690 61.845 173.195 ;
        RECT 60.655 172.095 60.985 172.465 ;
        RECT 61.220 172.390 61.390 172.645 ;
        RECT 61.220 172.060 61.505 172.390 ;
        RECT 61.220 171.915 61.390 172.060 ;
        RECT 60.725 171.745 61.390 171.915 ;
        RECT 61.675 171.890 61.845 172.690 ;
        RECT 59.695 171.405 60.445 171.605 ;
        RECT 59.685 170.815 60.035 171.225 ;
        RECT 60.205 171.015 60.445 171.405 ;
        RECT 60.725 170.985 60.895 171.745 ;
        RECT 61.075 170.815 61.405 171.575 ;
        RECT 61.575 170.985 61.845 171.890 ;
        RECT 62.015 172.690 62.275 173.195 ;
        RECT 62.455 172.985 62.785 173.365 ;
        RECT 62.965 172.815 63.135 173.195 ;
        RECT 62.015 171.890 62.185 172.690 ;
        RECT 62.470 172.645 63.135 172.815 ;
        RECT 63.485 172.815 63.655 173.195 ;
        RECT 63.835 172.985 64.165 173.365 ;
        RECT 63.485 172.645 64.150 172.815 ;
        RECT 64.345 172.690 64.605 173.195 ;
        RECT 62.470 172.390 62.640 172.645 ;
        RECT 62.355 172.060 62.640 172.390 ;
        RECT 62.875 172.095 63.205 172.465 ;
        RECT 63.415 172.095 63.755 172.465 ;
        RECT 63.980 172.390 64.150 172.645 ;
        RECT 62.470 171.915 62.640 172.060 ;
        RECT 63.980 172.060 64.255 172.390 ;
        RECT 63.980 171.915 64.150 172.060 ;
        RECT 62.015 170.985 62.285 171.890 ;
        RECT 62.470 171.745 63.135 171.915 ;
        RECT 62.455 170.815 62.785 171.575 ;
        RECT 62.965 170.985 63.135 171.745 ;
        RECT 63.475 171.745 64.150 171.915 ;
        RECT 64.425 171.890 64.605 172.690 ;
        RECT 63.475 170.985 63.655 171.745 ;
        RECT 63.835 170.815 64.165 171.575 ;
        RECT 64.335 170.985 64.605 171.890 ;
        RECT 64.775 172.690 65.035 173.195 ;
        RECT 65.215 172.985 65.545 173.365 ;
        RECT 65.725 172.815 65.895 173.195 ;
        RECT 64.775 171.890 64.955 172.690 ;
        RECT 65.230 172.645 65.895 172.815 ;
        RECT 66.245 172.815 66.415 173.195 ;
        RECT 66.595 172.985 66.925 173.365 ;
        RECT 66.245 172.645 66.910 172.815 ;
        RECT 67.105 172.690 67.365 173.195 ;
        RECT 65.230 172.390 65.400 172.645 ;
        RECT 65.125 172.060 65.400 172.390 ;
        RECT 65.625 172.095 65.965 172.465 ;
        RECT 66.175 172.095 66.505 172.465 ;
        RECT 66.740 172.390 66.910 172.645 ;
        RECT 65.230 171.915 65.400 172.060 ;
        RECT 66.740 172.060 67.025 172.390 ;
        RECT 66.740 171.915 66.910 172.060 ;
        RECT 64.775 170.985 65.045 171.890 ;
        RECT 65.230 171.745 65.905 171.915 ;
        RECT 65.215 170.815 65.545 171.575 ;
        RECT 65.725 170.985 65.905 171.745 ;
        RECT 66.245 171.745 66.910 171.915 ;
        RECT 67.195 171.890 67.365 172.690 ;
        RECT 67.535 172.640 67.825 173.365 ;
        RECT 68.545 172.815 68.715 173.195 ;
        RECT 68.895 172.985 69.225 173.365 ;
        RECT 68.545 172.645 69.210 172.815 ;
        RECT 69.405 172.690 69.665 173.195 ;
        RECT 68.475 172.095 68.815 172.465 ;
        RECT 69.040 172.390 69.210 172.645 ;
        RECT 69.040 172.060 69.315 172.390 ;
        RECT 66.245 170.985 66.415 171.745 ;
        RECT 66.595 170.815 66.925 171.575 ;
        RECT 67.095 170.985 67.365 171.890 ;
        RECT 67.535 170.815 67.825 171.980 ;
        RECT 69.040 171.915 69.210 172.060 ;
        RECT 68.535 171.745 69.210 171.915 ;
        RECT 69.485 171.890 69.665 172.690 ;
        RECT 69.895 172.545 70.105 173.365 ;
        RECT 70.275 172.565 70.605 173.195 ;
        RECT 70.275 171.965 70.525 172.565 ;
        RECT 70.775 172.545 71.005 173.365 ;
        RECT 71.370 172.715 71.700 173.180 ;
        RECT 71.870 172.895 72.040 173.365 ;
        RECT 72.210 172.715 72.540 173.195 ;
        RECT 71.370 172.545 72.540 172.715 ;
        RECT 70.695 172.125 71.025 172.375 ;
        RECT 71.215 172.165 71.860 172.375 ;
        RECT 72.030 172.165 72.600 172.375 ;
        RECT 72.770 171.995 72.940 173.195 ;
        RECT 73.480 172.795 73.650 173.000 ;
        RECT 68.535 170.985 68.715 171.745 ;
        RECT 68.895 170.815 69.225 171.575 ;
        RECT 69.395 170.985 69.665 171.890 ;
        RECT 69.895 170.815 70.105 171.955 ;
        RECT 70.275 170.985 70.605 171.965 ;
        RECT 70.775 170.815 71.005 171.955 ;
        RECT 71.430 170.815 71.760 171.915 ;
        RECT 72.235 171.585 72.940 171.995 ;
        RECT 73.110 172.625 73.650 172.795 ;
        RECT 73.930 172.625 74.100 173.365 ;
        RECT 74.365 172.625 74.725 173.000 ;
        RECT 74.985 172.815 75.155 173.195 ;
        RECT 75.370 172.985 75.700 173.365 ;
        RECT 74.985 172.645 75.700 172.815 ;
        RECT 73.110 171.925 73.280 172.625 ;
        RECT 73.450 172.125 73.780 172.455 ;
        RECT 73.950 172.125 74.300 172.455 ;
        RECT 73.110 171.755 73.735 171.925 ;
        RECT 73.950 171.585 74.215 172.125 ;
        RECT 74.470 171.970 74.725 172.625 ;
        RECT 74.895 172.095 75.250 172.465 ;
        RECT 75.530 172.455 75.700 172.645 ;
        RECT 75.870 172.620 76.125 173.195 ;
        RECT 75.530 172.125 75.785 172.455 ;
        RECT 72.235 171.415 74.215 171.585 ;
        RECT 72.235 170.985 72.560 171.415 ;
        RECT 72.730 170.815 73.060 171.235 ;
        RECT 73.805 170.815 74.215 171.245 ;
        RECT 74.385 170.985 74.725 171.970 ;
        RECT 75.530 171.915 75.700 172.125 ;
        RECT 74.985 171.745 75.700 171.915 ;
        RECT 75.955 171.890 76.125 172.620 ;
        RECT 76.300 172.525 76.560 173.365 ;
        RECT 76.735 172.855 77.040 173.365 ;
        RECT 76.735 172.125 77.050 172.685 ;
        RECT 77.220 172.375 77.470 173.185 ;
        RECT 77.640 172.840 77.900 173.365 ;
        RECT 78.080 172.375 78.330 173.185 ;
        RECT 78.500 172.805 78.760 173.365 ;
        RECT 78.930 172.715 79.190 173.170 ;
        RECT 79.360 172.885 79.620 173.365 ;
        RECT 79.790 172.715 80.050 173.170 ;
        RECT 80.220 172.885 80.480 173.365 ;
        RECT 80.650 172.715 80.910 173.170 ;
        RECT 81.080 172.885 81.325 173.365 ;
        RECT 81.495 172.715 81.770 173.170 ;
        RECT 81.940 172.885 82.185 173.365 ;
        RECT 82.355 172.715 82.615 173.170 ;
        RECT 82.795 172.885 83.045 173.365 ;
        RECT 83.215 172.715 83.475 173.170 ;
        RECT 83.655 172.885 83.905 173.365 ;
        RECT 84.075 172.715 84.335 173.170 ;
        RECT 84.515 172.885 84.775 173.365 ;
        RECT 84.945 172.715 85.205 173.170 ;
        RECT 85.375 172.885 85.675 173.365 ;
        RECT 78.930 172.545 85.675 172.715 ;
        RECT 85.935 172.615 87.145 173.365 ;
        RECT 77.220 172.125 84.340 172.375 ;
        RECT 74.985 170.985 75.155 171.745 ;
        RECT 75.370 170.815 75.700 171.575 ;
        RECT 75.870 170.985 76.125 171.890 ;
        RECT 76.300 170.815 76.560 171.965 ;
        RECT 76.745 170.815 77.040 171.625 ;
        RECT 77.220 170.985 77.465 172.125 ;
        RECT 77.640 170.815 77.900 171.625 ;
        RECT 78.080 170.990 78.330 172.125 ;
        RECT 84.510 171.955 85.675 172.545 ;
        RECT 78.930 171.730 85.675 171.955 ;
        RECT 85.935 171.905 86.455 172.445 ;
        RECT 86.625 172.075 87.145 172.615 ;
        RECT 78.930 171.715 84.335 171.730 ;
        RECT 78.500 170.820 78.760 171.615 ;
        RECT 78.930 170.990 79.190 171.715 ;
        RECT 79.360 170.820 79.620 171.545 ;
        RECT 79.790 170.990 80.050 171.715 ;
        RECT 80.220 170.820 80.480 171.545 ;
        RECT 80.650 170.990 80.910 171.715 ;
        RECT 81.080 170.820 81.340 171.545 ;
        RECT 81.510 170.990 81.770 171.715 ;
        RECT 81.940 170.820 82.185 171.545 ;
        RECT 82.355 170.990 82.615 171.715 ;
        RECT 82.800 170.820 83.045 171.545 ;
        RECT 83.215 170.990 83.475 171.715 ;
        RECT 83.660 170.820 83.905 171.545 ;
        RECT 84.075 170.990 84.335 171.715 ;
        RECT 84.520 170.820 84.775 171.545 ;
        RECT 84.945 170.990 85.235 171.730 ;
        RECT 78.500 170.815 84.775 170.820 ;
        RECT 85.405 170.815 85.675 171.560 ;
        RECT 85.935 170.815 87.145 171.905 ;
        RECT 15.930 170.645 87.230 170.815 ;
        RECT 16.015 169.555 17.225 170.645 ;
        RECT 17.395 169.555 19.065 170.645 ;
        RECT 16.015 168.845 16.535 169.385 ;
        RECT 16.705 169.015 17.225 169.555 ;
        RECT 17.395 168.865 18.145 169.385 ;
        RECT 18.315 169.035 19.065 169.555 ;
        RECT 19.240 169.505 19.575 170.475 ;
        RECT 19.745 169.505 19.915 170.645 ;
        RECT 20.085 170.305 22.115 170.475 ;
        RECT 16.015 168.095 17.225 168.845 ;
        RECT 17.395 168.095 19.065 168.865 ;
        RECT 19.240 168.835 19.410 169.505 ;
        RECT 20.085 169.335 20.255 170.305 ;
        RECT 19.580 169.005 19.835 169.335 ;
        RECT 20.060 169.005 20.255 169.335 ;
        RECT 20.425 169.965 21.550 170.135 ;
        RECT 19.665 168.835 19.835 169.005 ;
        RECT 20.425 168.835 20.595 169.965 ;
        RECT 19.240 168.265 19.495 168.835 ;
        RECT 19.665 168.665 20.595 168.835 ;
        RECT 20.765 169.625 21.775 169.795 ;
        RECT 20.765 168.825 20.935 169.625 ;
        RECT 20.420 168.630 20.595 168.665 ;
        RECT 19.665 168.095 19.995 168.495 ;
        RECT 20.420 168.265 20.950 168.630 ;
        RECT 21.140 168.605 21.415 169.425 ;
        RECT 21.135 168.435 21.415 168.605 ;
        RECT 21.140 168.265 21.415 168.435 ;
        RECT 21.585 168.265 21.775 169.625 ;
        RECT 21.945 169.640 22.115 170.305 ;
        RECT 22.285 169.885 22.455 170.645 ;
        RECT 22.690 169.885 23.205 170.295 ;
        RECT 21.945 169.450 22.695 169.640 ;
        RECT 22.865 169.075 23.205 169.885 ;
        RECT 23.375 169.555 25.965 170.645 ;
        RECT 21.975 168.905 23.205 169.075 ;
        RECT 21.955 168.095 22.465 168.630 ;
        RECT 22.685 168.300 22.930 168.905 ;
        RECT 23.375 168.865 24.585 169.385 ;
        RECT 24.755 169.035 25.965 169.555 ;
        RECT 26.145 170.035 26.475 170.465 ;
        RECT 26.655 170.205 26.850 170.645 ;
        RECT 27.020 170.035 27.350 170.465 ;
        RECT 26.145 169.865 27.350 170.035 ;
        RECT 26.145 169.535 27.040 169.865 ;
        RECT 27.520 169.695 27.795 170.465 ;
        RECT 27.210 169.505 27.795 169.695 ;
        RECT 26.150 169.005 26.445 169.335 ;
        RECT 26.625 169.005 27.040 169.335 ;
        RECT 23.375 168.095 25.965 168.865 ;
        RECT 26.145 168.095 26.445 168.825 ;
        RECT 26.625 168.385 26.855 169.005 ;
        RECT 27.210 168.835 27.385 169.505 ;
        RECT 28.895 169.480 29.185 170.645 ;
        RECT 29.390 169.855 29.925 170.475 ;
        RECT 27.055 168.655 27.385 168.835 ;
        RECT 27.555 168.685 27.795 169.335 ;
        RECT 29.390 168.835 29.705 169.855 ;
        RECT 30.095 169.845 30.425 170.645 ;
        RECT 31.665 170.035 31.995 170.465 ;
        RECT 32.175 170.205 32.370 170.645 ;
        RECT 32.540 170.035 32.870 170.465 ;
        RECT 31.665 169.865 32.870 170.035 ;
        RECT 30.910 169.675 31.300 169.850 ;
        RECT 29.875 169.505 31.300 169.675 ;
        RECT 31.665 169.535 32.560 169.865 ;
        RECT 33.040 169.695 33.315 170.465 ;
        RECT 32.730 169.505 33.315 169.695 ;
        RECT 34.420 169.505 34.755 170.475 ;
        RECT 34.925 169.505 35.095 170.645 ;
        RECT 35.265 170.305 37.295 170.475 ;
        RECT 29.875 169.005 30.045 169.505 ;
        RECT 27.055 168.275 27.280 168.655 ;
        RECT 27.450 168.095 27.780 168.485 ;
        RECT 28.895 168.095 29.185 168.820 ;
        RECT 29.390 168.265 30.005 168.835 ;
        RECT 30.295 168.775 30.560 169.335 ;
        RECT 30.730 168.605 30.900 169.505 ;
        RECT 31.070 168.775 31.425 169.335 ;
        RECT 31.670 169.005 31.965 169.335 ;
        RECT 32.145 169.005 32.560 169.335 ;
        RECT 30.175 168.095 30.390 168.605 ;
        RECT 30.620 168.275 30.900 168.605 ;
        RECT 31.080 168.095 31.320 168.605 ;
        RECT 31.665 168.095 31.965 168.825 ;
        RECT 32.145 168.385 32.375 169.005 ;
        RECT 32.730 168.835 32.905 169.505 ;
        RECT 32.575 168.655 32.905 168.835 ;
        RECT 33.075 168.685 33.315 169.335 ;
        RECT 34.420 168.835 34.590 169.505 ;
        RECT 35.265 169.335 35.435 170.305 ;
        RECT 34.760 169.005 35.015 169.335 ;
        RECT 35.240 169.005 35.435 169.335 ;
        RECT 35.605 169.965 36.730 170.135 ;
        RECT 34.845 168.835 35.015 169.005 ;
        RECT 35.605 168.835 35.775 169.965 ;
        RECT 32.575 168.275 32.800 168.655 ;
        RECT 32.970 168.095 33.300 168.485 ;
        RECT 34.420 168.265 34.675 168.835 ;
        RECT 34.845 168.665 35.775 168.835 ;
        RECT 35.945 169.625 36.955 169.795 ;
        RECT 35.945 168.825 36.115 169.625 ;
        RECT 35.600 168.630 35.775 168.665 ;
        RECT 34.845 168.095 35.175 168.495 ;
        RECT 35.600 168.265 36.130 168.630 ;
        RECT 36.320 168.605 36.595 169.425 ;
        RECT 36.315 168.435 36.595 168.605 ;
        RECT 36.320 168.265 36.595 168.435 ;
        RECT 36.765 168.265 36.955 169.625 ;
        RECT 37.125 169.640 37.295 170.305 ;
        RECT 37.465 169.885 37.635 170.645 ;
        RECT 37.870 169.885 38.385 170.295 ;
        RECT 37.125 169.450 37.875 169.640 ;
        RECT 38.045 169.075 38.385 169.885 ;
        RECT 38.595 169.505 38.825 170.645 ;
        RECT 38.995 169.495 39.325 170.475 ;
        RECT 39.495 169.505 39.705 170.645 ;
        RECT 39.935 169.505 40.195 170.645 ;
        RECT 40.365 169.495 40.695 170.475 ;
        RECT 40.865 169.505 41.145 170.645 ;
        RECT 42.245 170.035 42.575 170.465 ;
        RECT 42.755 170.205 42.950 170.645 ;
        RECT 43.120 170.035 43.450 170.465 ;
        RECT 42.245 169.865 43.450 170.035 ;
        RECT 42.245 169.535 43.140 169.865 ;
        RECT 43.620 169.695 43.895 170.465 ;
        RECT 43.310 169.505 43.895 169.695 ;
        RECT 44.115 169.505 44.345 170.645 ;
        RECT 38.575 169.085 38.905 169.335 ;
        RECT 37.155 168.905 38.385 169.075 ;
        RECT 37.135 168.095 37.645 168.630 ;
        RECT 37.865 168.300 38.110 168.905 ;
        RECT 38.595 168.095 38.825 168.915 ;
        RECT 39.075 168.895 39.325 169.495 ;
        RECT 39.955 169.085 40.290 169.335 ;
        RECT 38.995 168.265 39.325 168.895 ;
        RECT 39.495 168.095 39.705 168.915 ;
        RECT 40.460 168.895 40.630 169.495 ;
        RECT 40.800 169.065 41.135 169.335 ;
        RECT 42.250 169.005 42.545 169.335 ;
        RECT 42.725 169.005 43.140 169.335 ;
        RECT 39.935 168.265 40.630 168.895 ;
        RECT 40.835 168.095 41.145 168.895 ;
        RECT 42.245 168.095 42.545 168.825 ;
        RECT 42.725 168.385 42.955 169.005 ;
        RECT 43.310 168.835 43.485 169.505 ;
        RECT 44.515 169.495 44.845 170.475 ;
        RECT 45.015 169.505 45.225 170.645 ;
        RECT 45.455 169.555 46.665 170.645 ;
        RECT 43.155 168.655 43.485 168.835 ;
        RECT 43.655 168.685 43.895 169.335 ;
        RECT 44.095 169.085 44.425 169.335 ;
        RECT 43.155 168.275 43.380 168.655 ;
        RECT 43.550 168.095 43.880 168.485 ;
        RECT 44.115 168.095 44.345 168.915 ;
        RECT 44.595 168.895 44.845 169.495 ;
        RECT 44.515 168.265 44.845 168.895 ;
        RECT 45.015 168.095 45.225 168.915 ;
        RECT 45.455 168.845 45.975 169.385 ;
        RECT 46.145 169.015 46.665 169.555 ;
        RECT 46.835 169.505 47.095 170.645 ;
        RECT 47.265 169.495 47.595 170.475 ;
        RECT 47.765 169.505 48.045 170.645 ;
        RECT 48.215 170.210 53.560 170.645 ;
        RECT 46.855 169.085 47.190 169.335 ;
        RECT 47.360 168.895 47.530 169.495 ;
        RECT 47.700 169.065 48.035 169.335 ;
        RECT 45.455 168.095 46.665 168.845 ;
        RECT 46.835 168.265 47.530 168.895 ;
        RECT 47.735 168.095 48.045 168.895 ;
        RECT 49.800 168.640 50.140 169.470 ;
        RECT 51.620 168.960 51.970 170.210 ;
        RECT 54.655 169.480 54.945 170.645 ;
        RECT 55.115 169.505 55.390 170.475 ;
        RECT 55.600 169.845 55.880 170.645 ;
        RECT 56.050 170.135 57.665 170.465 ;
        RECT 56.050 169.795 57.225 169.965 ;
        RECT 56.050 169.675 56.220 169.795 ;
        RECT 55.560 169.505 56.220 169.675 ;
        RECT 48.215 168.095 53.560 168.640 ;
        RECT 54.655 168.095 54.945 168.820 ;
        RECT 55.115 168.770 55.285 169.505 ;
        RECT 55.560 169.335 55.730 169.505 ;
        RECT 56.480 169.335 56.725 169.625 ;
        RECT 56.895 169.505 57.225 169.795 ;
        RECT 57.485 169.335 57.655 169.895 ;
        RECT 57.905 169.505 58.165 170.645 ;
        RECT 58.335 169.555 60.005 170.645 ;
        RECT 55.455 169.005 55.730 169.335 ;
        RECT 55.900 169.005 56.725 169.335 ;
        RECT 56.940 169.005 57.655 169.335 ;
        RECT 57.825 169.085 58.160 169.335 ;
        RECT 55.560 168.835 55.730 169.005 ;
        RECT 57.405 168.915 57.655 169.005 ;
        RECT 55.115 168.425 55.390 168.770 ;
        RECT 55.560 168.665 57.225 168.835 ;
        RECT 55.580 168.095 55.955 168.495 ;
        RECT 56.125 168.315 56.295 168.665 ;
        RECT 56.465 168.095 56.795 168.495 ;
        RECT 56.965 168.265 57.225 168.665 ;
        RECT 57.405 168.495 57.735 168.915 ;
        RECT 57.905 168.095 58.165 168.915 ;
        RECT 58.335 168.865 59.085 169.385 ;
        RECT 59.255 169.035 60.005 169.555 ;
        RECT 60.640 169.695 60.905 170.465 ;
        RECT 61.075 169.925 61.405 170.645 ;
        RECT 61.595 170.105 61.855 170.465 ;
        RECT 62.025 170.275 62.355 170.645 ;
        RECT 62.525 170.105 62.785 170.465 ;
        RECT 61.595 169.875 62.785 170.105 ;
        RECT 63.355 169.695 63.645 170.465 ;
        RECT 58.335 168.095 60.005 168.865 ;
        RECT 60.640 168.275 60.975 169.695 ;
        RECT 61.150 169.515 63.645 169.695 ;
        RECT 63.875 169.805 64.130 170.475 ;
        RECT 64.300 169.885 64.630 170.645 ;
        RECT 64.800 170.045 65.050 170.475 ;
        RECT 65.220 170.225 65.575 170.645 ;
        RECT 65.765 170.305 66.935 170.475 ;
        RECT 65.765 170.265 66.095 170.305 ;
        RECT 66.205 170.045 66.435 170.135 ;
        RECT 64.800 169.805 66.435 170.045 ;
        RECT 66.605 169.805 66.935 170.305 ;
        RECT 63.875 169.795 64.085 169.805 ;
        RECT 61.150 168.825 61.375 169.515 ;
        RECT 61.575 169.005 61.855 169.335 ;
        RECT 62.035 169.005 62.610 169.335 ;
        RECT 62.790 169.005 63.225 169.335 ;
        RECT 63.405 169.005 63.675 169.335 ;
        RECT 61.150 168.635 63.635 168.825 ;
        RECT 61.155 168.095 61.900 168.465 ;
        RECT 62.465 168.275 62.720 168.635 ;
        RECT 62.900 168.095 63.230 168.465 ;
        RECT 63.410 168.275 63.635 168.635 ;
        RECT 63.875 168.675 64.045 169.795 ;
        RECT 67.105 169.635 67.275 170.475 ;
        RECT 64.215 169.465 67.275 169.635 ;
        RECT 67.545 170.035 67.875 170.465 ;
        RECT 68.055 170.205 68.250 170.645 ;
        RECT 68.420 170.035 68.750 170.465 ;
        RECT 67.545 169.865 68.750 170.035 ;
        RECT 67.545 169.535 68.440 169.865 ;
        RECT 68.920 169.695 69.195 170.465 ;
        RECT 70.305 169.845 70.635 170.645 ;
        RECT 70.815 170.305 72.245 170.475 ;
        RECT 68.610 169.505 69.195 169.695 ;
        RECT 70.815 169.675 71.065 170.305 ;
        RECT 70.295 169.505 71.065 169.675 ;
        RECT 64.215 168.915 64.385 169.465 ;
        RECT 64.615 169.085 64.980 169.285 ;
        RECT 65.150 169.085 65.480 169.285 ;
        RECT 64.215 168.745 65.015 168.915 ;
        RECT 63.875 168.595 64.060 168.675 ;
        RECT 63.875 168.265 64.130 168.595 ;
        RECT 64.345 168.095 64.675 168.575 ;
        RECT 64.845 168.515 65.015 168.745 ;
        RECT 65.195 168.685 65.480 169.085 ;
        RECT 65.750 169.085 66.225 169.285 ;
        RECT 66.395 169.085 66.840 169.285 ;
        RECT 67.010 169.085 67.360 169.295 ;
        RECT 65.750 168.685 66.030 169.085 ;
        RECT 67.550 169.005 67.845 169.335 ;
        RECT 68.025 169.005 68.440 169.335 ;
        RECT 66.210 168.745 67.275 168.915 ;
        RECT 66.210 168.515 66.380 168.745 ;
        RECT 64.845 168.265 66.380 168.515 ;
        RECT 66.605 168.095 66.935 168.575 ;
        RECT 67.105 168.265 67.275 168.745 ;
        RECT 67.545 168.095 67.845 168.825 ;
        RECT 68.025 168.385 68.255 169.005 ;
        RECT 68.610 168.835 68.785 169.505 ;
        RECT 68.455 168.655 68.785 168.835 ;
        RECT 68.955 168.685 69.195 169.335 ;
        RECT 70.295 168.835 70.465 169.505 ;
        RECT 70.635 169.005 71.040 169.335 ;
        RECT 71.255 169.005 71.505 170.135 ;
        RECT 71.705 169.335 71.905 170.135 ;
        RECT 72.075 169.625 72.245 170.305 ;
        RECT 72.415 169.795 72.730 170.645 ;
        RECT 72.905 169.845 73.345 170.475 ;
        RECT 72.075 169.455 72.865 169.625 ;
        RECT 71.705 169.005 71.950 169.335 ;
        RECT 72.135 169.005 72.525 169.285 ;
        RECT 72.695 169.005 72.865 169.455 ;
        RECT 73.035 168.835 73.345 169.845 ;
        RECT 74.505 169.675 74.865 169.850 ;
        RECT 75.450 169.845 75.620 170.645 ;
        RECT 75.790 170.015 76.120 170.475 ;
        RECT 76.290 170.185 76.460 170.645 ;
        RECT 75.790 169.845 76.565 170.015 ;
        RECT 74.505 169.505 75.965 169.675 ;
        RECT 74.500 169.285 74.695 169.335 ;
        RECT 74.495 169.115 74.695 169.285 ;
        RECT 68.455 168.275 68.680 168.655 ;
        RECT 68.850 168.095 69.180 168.485 ;
        RECT 70.295 168.265 70.785 168.835 ;
        RECT 70.955 168.665 72.115 168.835 ;
        RECT 70.955 168.265 71.185 168.665 ;
        RECT 71.355 168.095 71.775 168.495 ;
        RECT 71.945 168.265 72.115 168.665 ;
        RECT 72.285 168.095 72.735 168.835 ;
        RECT 72.905 168.275 73.345 168.835 ;
        RECT 74.500 168.775 74.695 169.115 ;
        RECT 74.865 168.605 75.045 169.505 ;
        RECT 75.215 168.775 75.625 169.335 ;
        RECT 75.795 169.005 75.965 169.505 ;
        RECT 76.135 168.835 76.565 169.845 ;
        RECT 76.790 169.775 77.075 170.645 ;
        RECT 77.245 170.015 77.505 170.475 ;
        RECT 77.680 170.185 77.935 170.645 ;
        RECT 78.105 170.015 78.365 170.475 ;
        RECT 77.245 169.845 78.365 170.015 ;
        RECT 78.535 169.845 78.845 170.645 ;
        RECT 77.245 169.595 77.505 169.845 ;
        RECT 79.015 169.675 79.325 170.475 ;
        RECT 75.870 168.665 76.565 168.835 ;
        RECT 76.750 169.425 77.505 169.595 ;
        RECT 78.295 169.505 79.325 169.675 ;
        RECT 76.750 168.915 77.155 169.425 ;
        RECT 78.295 169.255 78.465 169.505 ;
        RECT 77.325 169.085 78.465 169.255 ;
        RECT 76.750 168.745 78.400 168.915 ;
        RECT 78.635 168.765 78.985 169.335 ;
        RECT 74.455 168.095 74.695 168.605 ;
        RECT 74.865 168.265 75.155 168.605 ;
        RECT 75.385 168.095 75.700 168.605 ;
        RECT 75.870 168.395 76.040 168.665 ;
        RECT 76.210 168.095 76.540 168.495 ;
        RECT 76.795 168.095 77.075 168.575 ;
        RECT 77.245 168.355 77.505 168.745 ;
        RECT 77.680 168.095 77.935 168.575 ;
        RECT 78.105 168.355 78.400 168.745 ;
        RECT 79.155 168.595 79.325 169.505 ;
        RECT 80.415 169.480 80.705 170.645 ;
        RECT 80.915 170.305 82.055 170.475 ;
        RECT 80.915 169.845 81.215 170.305 ;
        RECT 81.385 169.675 81.715 170.135 ;
        RECT 80.955 169.625 81.715 169.675 ;
        RECT 80.935 169.455 81.715 169.625 ;
        RECT 81.885 169.675 82.055 170.305 ;
        RECT 82.225 169.845 82.555 170.645 ;
        RECT 82.725 169.675 83.000 170.475 ;
        RECT 81.885 169.465 83.000 169.675 ;
        RECT 83.175 169.675 83.485 170.475 ;
        RECT 83.655 169.845 83.965 170.645 ;
        RECT 84.135 170.015 84.395 170.475 ;
        RECT 84.565 170.185 84.820 170.645 ;
        RECT 84.995 170.015 85.255 170.475 ;
        RECT 84.135 169.845 85.255 170.015 ;
        RECT 83.175 169.505 84.205 169.675 ;
        RECT 80.955 168.915 81.170 169.455 ;
        RECT 81.340 169.085 82.110 169.285 ;
        RECT 82.280 169.085 83.000 169.285 ;
        RECT 78.580 168.095 78.855 168.575 ;
        RECT 79.025 168.265 79.325 168.595 ;
        RECT 80.415 168.095 80.705 168.820 ;
        RECT 80.955 168.745 82.555 168.915 ;
        RECT 81.385 168.735 82.555 168.745 ;
        RECT 80.925 168.095 81.215 168.565 ;
        RECT 81.385 168.265 81.715 168.735 ;
        RECT 81.885 168.095 82.055 168.565 ;
        RECT 82.225 168.265 82.555 168.735 ;
        RECT 82.725 168.095 83.000 168.915 ;
        RECT 83.175 168.595 83.345 169.505 ;
        RECT 83.515 168.765 83.865 169.335 ;
        RECT 84.035 169.255 84.205 169.505 ;
        RECT 84.995 169.595 85.255 169.845 ;
        RECT 85.425 169.775 85.710 170.645 ;
        RECT 84.995 169.425 85.750 169.595 ;
        RECT 84.035 169.085 85.175 169.255 ;
        RECT 85.345 168.915 85.750 169.425 ;
        RECT 85.935 169.555 87.145 170.645 ;
        RECT 85.935 169.015 86.455 169.555 ;
        RECT 84.100 168.745 85.750 168.915 ;
        RECT 86.625 168.845 87.145 169.385 ;
        RECT 83.175 168.265 83.475 168.595 ;
        RECT 83.645 168.095 83.920 168.575 ;
        RECT 84.100 168.355 84.395 168.745 ;
        RECT 84.565 168.095 84.820 168.575 ;
        RECT 84.995 168.355 85.255 168.745 ;
        RECT 85.425 168.095 85.705 168.575 ;
        RECT 85.935 168.095 87.145 168.845 ;
        RECT 15.930 167.925 87.230 168.095 ;
        RECT 16.015 167.175 17.225 167.925 ;
        RECT 16.015 166.635 16.535 167.175 ;
        RECT 17.395 167.155 19.985 167.925 ;
        RECT 16.705 166.465 17.225 167.005 ;
        RECT 17.395 166.635 18.605 167.155 ;
        RECT 20.430 167.115 20.675 167.720 ;
        RECT 20.895 167.390 21.405 167.925 ;
        RECT 18.775 166.465 19.985 166.985 ;
        RECT 16.015 165.375 17.225 166.465 ;
        RECT 17.395 165.375 19.985 166.465 ;
        RECT 20.155 166.945 21.385 167.115 ;
        RECT 20.155 166.135 20.495 166.945 ;
        RECT 20.665 166.380 21.415 166.570 ;
        RECT 20.155 165.725 20.670 166.135 ;
        RECT 20.905 165.375 21.075 166.135 ;
        RECT 21.245 165.715 21.415 166.380 ;
        RECT 21.585 166.395 21.775 167.755 ;
        RECT 21.945 166.905 22.220 167.755 ;
        RECT 22.410 167.390 22.940 167.755 ;
        RECT 23.365 167.525 23.695 167.925 ;
        RECT 22.765 167.355 22.940 167.390 ;
        RECT 21.945 166.735 22.225 166.905 ;
        RECT 21.945 166.595 22.220 166.735 ;
        RECT 22.425 166.395 22.595 167.195 ;
        RECT 21.585 166.225 22.595 166.395 ;
        RECT 22.765 167.185 23.695 167.355 ;
        RECT 23.865 167.185 24.120 167.755 ;
        RECT 22.765 166.055 22.935 167.185 ;
        RECT 23.525 167.015 23.695 167.185 ;
        RECT 21.810 165.885 22.935 166.055 ;
        RECT 23.105 166.685 23.300 167.015 ;
        RECT 23.525 166.685 23.780 167.015 ;
        RECT 23.105 165.715 23.275 166.685 ;
        RECT 23.950 166.515 24.120 167.185 ;
        RECT 24.295 167.315 24.635 167.730 ;
        RECT 24.805 167.485 24.975 167.925 ;
        RECT 25.145 167.535 26.395 167.715 ;
        RECT 25.145 167.315 25.475 167.535 ;
        RECT 26.665 167.465 26.835 167.925 ;
        RECT 24.295 167.145 25.475 167.315 ;
        RECT 25.645 167.295 26.010 167.365 ;
        RECT 25.645 167.115 26.895 167.295 ;
        RECT 24.295 166.735 24.760 166.935 ;
        RECT 24.935 166.685 25.265 166.935 ;
        RECT 25.435 166.905 25.900 166.935 ;
        RECT 25.435 166.735 25.905 166.905 ;
        RECT 25.435 166.685 25.900 166.735 ;
        RECT 26.095 166.685 26.450 166.935 ;
        RECT 24.935 166.565 25.115 166.685 ;
        RECT 21.245 165.545 23.275 165.715 ;
        RECT 23.445 165.375 23.615 166.515 ;
        RECT 23.785 165.545 24.120 166.515 ;
        RECT 24.295 165.375 24.615 166.555 ;
        RECT 24.785 166.395 25.115 166.565 ;
        RECT 26.620 166.515 26.895 167.115 ;
        RECT 24.785 165.605 24.985 166.395 ;
        RECT 25.285 166.305 26.895 166.515 ;
        RECT 25.285 166.205 25.695 166.305 ;
        RECT 25.310 165.545 25.695 166.205 ;
        RECT 26.090 165.375 26.875 166.135 ;
        RECT 27.065 165.545 27.345 167.645 ;
        RECT 27.515 167.380 32.860 167.925 ;
        RECT 33.035 167.380 38.380 167.925 ;
        RECT 29.100 166.550 29.440 167.380 ;
        RECT 30.920 165.810 31.270 167.060 ;
        RECT 34.620 166.550 34.960 167.380 ;
        RECT 38.555 167.155 41.145 167.925 ;
        RECT 41.775 167.200 42.065 167.925 ;
        RECT 42.235 167.155 44.825 167.925 ;
        RECT 45.455 167.185 45.795 167.755 ;
        RECT 45.990 167.260 46.160 167.925 ;
        RECT 46.440 167.585 46.660 167.630 ;
        RECT 46.435 167.415 46.660 167.585 ;
        RECT 46.830 167.445 47.275 167.615 ;
        RECT 46.440 167.275 46.660 167.415 ;
        RECT 36.440 165.810 36.790 167.060 ;
        RECT 38.555 166.635 39.765 167.155 ;
        RECT 39.935 166.465 41.145 166.985 ;
        RECT 42.235 166.635 43.445 167.155 ;
        RECT 27.515 165.375 32.860 165.810 ;
        RECT 33.035 165.375 38.380 165.810 ;
        RECT 38.555 165.375 41.145 166.465 ;
        RECT 41.775 165.375 42.065 166.540 ;
        RECT 43.615 166.465 44.825 166.985 ;
        RECT 42.235 165.375 44.825 166.465 ;
        RECT 45.455 166.215 45.630 167.185 ;
        RECT 46.440 167.105 46.935 167.275 ;
        RECT 45.800 166.565 45.970 167.015 ;
        RECT 46.140 166.735 46.590 166.935 ;
        RECT 46.760 166.910 46.935 167.105 ;
        RECT 47.105 166.655 47.275 167.445 ;
        RECT 47.445 167.320 47.695 167.690 ;
        RECT 47.525 166.935 47.695 167.320 ;
        RECT 47.865 167.285 48.115 167.690 ;
        RECT 48.285 167.455 48.455 167.925 ;
        RECT 48.625 167.285 48.965 167.690 ;
        RECT 47.865 167.105 48.965 167.285 ;
        RECT 49.135 167.155 50.805 167.925 ;
        RECT 50.985 167.200 51.315 167.710 ;
        RECT 51.485 167.525 51.815 167.925 ;
        RECT 52.865 167.355 53.195 167.695 ;
        RECT 53.365 167.525 53.695 167.925 ;
        RECT 47.525 166.765 47.720 166.935 ;
        RECT 45.800 166.395 46.195 166.565 ;
        RECT 47.105 166.515 47.380 166.655 ;
        RECT 45.455 165.545 45.715 166.215 ;
        RECT 46.025 166.125 46.195 166.395 ;
        RECT 46.365 166.295 47.380 166.515 ;
        RECT 47.550 166.515 47.720 166.765 ;
        RECT 47.890 166.685 48.450 166.935 ;
        RECT 47.550 166.125 48.105 166.515 ;
        RECT 46.025 165.955 48.105 166.125 ;
        RECT 45.885 165.375 46.215 165.775 ;
        RECT 47.085 165.375 47.485 165.775 ;
        RECT 47.775 165.720 48.105 165.955 ;
        RECT 48.275 165.585 48.450 166.685 ;
        RECT 48.620 166.365 48.965 166.935 ;
        RECT 49.135 166.635 49.885 167.155 ;
        RECT 50.055 166.465 50.805 166.985 ;
        RECT 48.620 165.375 48.965 166.195 ;
        RECT 49.135 165.375 50.805 166.465 ;
        RECT 50.985 166.435 51.175 167.200 ;
        RECT 51.485 167.185 53.850 167.355 ;
        RECT 51.485 167.015 51.655 167.185 ;
        RECT 51.345 166.685 51.655 167.015 ;
        RECT 51.825 166.685 52.130 167.015 ;
        RECT 50.985 165.585 51.315 166.435 ;
        RECT 51.485 165.375 51.735 166.515 ;
        RECT 51.915 166.355 52.130 166.685 ;
        RECT 52.305 166.355 52.590 167.015 ;
        RECT 52.785 166.355 53.050 167.015 ;
        RECT 53.265 166.355 53.510 167.015 ;
        RECT 53.680 166.185 53.850 167.185 ;
        RECT 54.400 167.145 54.900 167.755 ;
        RECT 54.195 166.685 54.545 166.935 ;
        RECT 54.730 166.515 54.900 167.145 ;
        RECT 55.530 167.275 55.860 167.755 ;
        RECT 56.030 167.465 56.255 167.925 ;
        RECT 56.425 167.275 56.755 167.755 ;
        RECT 55.530 167.105 56.755 167.275 ;
        RECT 56.945 167.125 57.195 167.925 ;
        RECT 57.365 167.125 57.705 167.755 ;
        RECT 58.040 167.415 58.280 167.925 ;
        RECT 58.460 167.415 58.740 167.745 ;
        RECT 58.970 167.415 59.185 167.925 ;
        RECT 55.070 166.735 55.400 166.935 ;
        RECT 55.570 166.735 55.900 166.935 ;
        RECT 56.070 166.735 56.490 166.935 ;
        RECT 56.665 166.765 57.360 166.935 ;
        RECT 56.665 166.515 56.835 166.765 ;
        RECT 57.530 166.515 57.705 167.125 ;
        RECT 57.935 166.685 58.290 167.245 ;
        RECT 58.460 166.515 58.630 167.415 ;
        RECT 58.800 166.685 59.065 167.245 ;
        RECT 59.355 167.185 59.970 167.755 ;
        RECT 59.315 166.515 59.485 167.015 ;
        RECT 51.925 166.015 53.215 166.185 ;
        RECT 51.925 165.595 52.175 166.015 ;
        RECT 52.405 165.375 52.735 165.845 ;
        RECT 52.965 165.595 53.215 166.015 ;
        RECT 53.395 166.015 53.850 166.185 ;
        RECT 54.400 166.345 56.835 166.515 ;
        RECT 53.395 165.585 53.725 166.015 ;
        RECT 54.400 165.545 54.730 166.345 ;
        RECT 54.900 165.375 55.230 166.175 ;
        RECT 55.530 165.545 55.860 166.345 ;
        RECT 56.505 165.375 56.755 166.175 ;
        RECT 57.025 165.375 57.195 166.515 ;
        RECT 57.365 165.545 57.705 166.515 ;
        RECT 58.060 166.345 59.485 166.515 ;
        RECT 58.060 166.170 58.450 166.345 ;
        RECT 58.935 165.375 59.265 166.175 ;
        RECT 59.655 166.165 59.970 167.185 ;
        RECT 60.175 167.125 60.870 167.755 ;
        RECT 61.075 167.125 61.385 167.925 ;
        RECT 61.555 167.155 64.145 167.925 ;
        RECT 64.340 167.535 64.670 167.925 ;
        RECT 64.840 167.365 65.065 167.745 ;
        RECT 60.195 166.685 60.530 166.935 ;
        RECT 60.700 166.565 60.870 167.125 ;
        RECT 61.040 166.685 61.375 166.955 ;
        RECT 61.555 166.635 62.765 167.155 ;
        RECT 60.695 166.525 60.870 166.565 ;
        RECT 59.435 165.545 59.970 166.165 ;
        RECT 60.175 165.375 60.435 166.515 ;
        RECT 60.605 165.545 60.935 166.525 ;
        RECT 61.105 165.375 61.385 166.515 ;
        RECT 62.935 166.465 64.145 166.985 ;
        RECT 64.325 166.685 64.565 167.335 ;
        RECT 64.735 167.185 65.065 167.365 ;
        RECT 64.735 166.515 64.910 167.185 ;
        RECT 65.265 167.015 65.495 167.635 ;
        RECT 65.675 167.195 65.975 167.925 ;
        RECT 66.245 167.375 66.415 167.755 ;
        RECT 66.595 167.545 66.925 167.925 ;
        RECT 66.245 167.205 66.910 167.375 ;
        RECT 67.105 167.250 67.365 167.755 ;
        RECT 65.080 166.685 65.495 167.015 ;
        RECT 65.675 166.685 65.970 167.015 ;
        RECT 66.175 166.655 66.515 167.025 ;
        RECT 66.740 166.950 66.910 167.205 ;
        RECT 61.555 165.375 64.145 166.465 ;
        RECT 64.325 166.325 64.910 166.515 ;
        RECT 66.740 166.620 67.015 166.950 ;
        RECT 64.325 165.555 64.600 166.325 ;
        RECT 65.080 166.155 65.975 166.485 ;
        RECT 66.740 166.475 66.910 166.620 ;
        RECT 64.770 165.985 65.975 166.155 ;
        RECT 64.770 165.555 65.100 165.985 ;
        RECT 65.270 165.375 65.465 165.815 ;
        RECT 65.645 165.555 65.975 165.985 ;
        RECT 66.235 166.305 66.910 166.475 ;
        RECT 67.185 166.450 67.365 167.250 ;
        RECT 67.535 167.200 67.825 167.925 ;
        RECT 69.005 167.375 69.175 167.755 ;
        RECT 69.355 167.545 69.685 167.925 ;
        RECT 69.005 167.205 69.670 167.375 ;
        RECT 69.865 167.250 70.125 167.755 ;
        RECT 68.935 166.655 69.265 167.025 ;
        RECT 69.500 166.950 69.670 167.205 ;
        RECT 69.500 166.620 69.785 166.950 ;
        RECT 66.235 165.545 66.415 166.305 ;
        RECT 66.595 165.375 66.925 166.135 ;
        RECT 67.095 165.545 67.365 166.450 ;
        RECT 67.535 165.375 67.825 166.540 ;
        RECT 69.500 166.475 69.670 166.620 ;
        RECT 69.005 166.305 69.670 166.475 ;
        RECT 69.955 166.450 70.125 167.250 ;
        RECT 70.385 167.375 70.555 167.755 ;
        RECT 70.735 167.545 71.065 167.925 ;
        RECT 70.385 167.205 71.050 167.375 ;
        RECT 71.245 167.250 71.505 167.755 ;
        RECT 70.315 166.655 70.645 167.025 ;
        RECT 70.880 166.950 71.050 167.205 ;
        RECT 70.880 166.620 71.165 166.950 ;
        RECT 70.880 166.475 71.050 166.620 ;
        RECT 69.005 165.545 69.175 166.305 ;
        RECT 69.355 165.375 69.685 166.135 ;
        RECT 69.855 165.545 70.125 166.450 ;
        RECT 70.385 166.305 71.050 166.475 ;
        RECT 71.335 166.450 71.505 167.250 ;
        RECT 70.385 165.545 70.555 166.305 ;
        RECT 70.735 165.375 71.065 166.135 ;
        RECT 71.235 165.545 71.505 166.450 ;
        RECT 71.675 167.185 72.035 167.560 ;
        RECT 72.300 167.185 72.470 167.925 ;
        RECT 72.750 167.355 72.920 167.560 ;
        RECT 72.750 167.185 73.290 167.355 ;
        RECT 71.675 166.530 71.930 167.185 ;
        RECT 72.100 166.685 72.450 167.015 ;
        RECT 72.620 166.685 72.950 167.015 ;
        RECT 71.675 165.545 72.015 166.530 ;
        RECT 72.185 166.145 72.450 166.685 ;
        RECT 73.120 166.485 73.290 167.185 ;
        RECT 72.665 166.315 73.290 166.485 ;
        RECT 73.460 166.555 73.630 167.755 ;
        RECT 73.860 167.275 74.190 167.755 ;
        RECT 74.360 167.455 74.530 167.925 ;
        RECT 74.700 167.275 75.030 167.740 ;
        RECT 73.860 167.105 75.030 167.275 ;
        RECT 75.370 167.355 75.625 167.705 ;
        RECT 75.795 167.525 76.125 167.925 ;
        RECT 76.295 167.355 76.465 167.705 ;
        RECT 76.635 167.525 77.015 167.925 ;
        RECT 75.370 167.185 77.035 167.355 ;
        RECT 77.205 167.250 77.480 167.595 ;
        RECT 78.580 167.420 78.915 167.925 ;
        RECT 79.085 167.355 79.325 167.730 ;
        RECT 79.605 167.595 79.775 167.740 ;
        RECT 79.605 167.400 79.980 167.595 ;
        RECT 80.340 167.430 80.735 167.925 ;
        RECT 76.865 167.015 77.035 167.185 ;
        RECT 73.800 166.725 74.370 166.935 ;
        RECT 74.540 166.725 75.185 166.935 ;
        RECT 75.355 166.685 75.700 167.015 ;
        RECT 75.870 166.685 76.695 167.015 ;
        RECT 76.865 166.685 77.140 167.015 ;
        RECT 73.460 166.145 74.165 166.555 ;
        RECT 72.185 165.975 74.165 166.145 ;
        RECT 72.185 165.375 72.595 165.805 ;
        RECT 73.340 165.375 73.670 165.795 ;
        RECT 73.840 165.545 74.165 165.975 ;
        RECT 74.640 165.375 74.970 166.475 ;
        RECT 75.375 166.225 75.700 166.515 ;
        RECT 75.870 166.395 76.065 166.685 ;
        RECT 76.865 166.515 77.035 166.685 ;
        RECT 77.310 166.515 77.480 167.250 ;
        RECT 76.375 166.345 77.035 166.515 ;
        RECT 76.375 166.225 76.545 166.345 ;
        RECT 75.375 166.055 76.545 166.225 ;
        RECT 75.355 165.595 76.545 165.885 ;
        RECT 76.715 165.375 76.995 166.175 ;
        RECT 77.205 165.545 77.480 166.515 ;
        RECT 78.635 166.395 78.935 167.245 ;
        RECT 79.105 167.205 79.325 167.355 ;
        RECT 79.105 166.875 79.640 167.205 ;
        RECT 79.810 167.065 79.980 167.400 ;
        RECT 80.905 167.235 81.145 167.755 ;
        RECT 81.335 167.265 81.610 167.925 ;
        RECT 81.780 167.295 82.030 167.755 ;
        RECT 82.205 167.430 82.535 167.925 ;
        RECT 79.105 166.225 79.340 166.875 ;
        RECT 79.810 166.705 80.795 167.065 ;
        RECT 78.665 165.995 79.340 166.225 ;
        RECT 79.510 166.685 80.795 166.705 ;
        RECT 79.510 166.535 80.370 166.685 ;
        RECT 78.665 165.565 78.835 165.995 ;
        RECT 79.005 165.375 79.335 165.825 ;
        RECT 79.510 165.590 79.795 166.535 ;
        RECT 80.970 166.430 81.145 167.235 ;
        RECT 81.780 167.085 81.950 167.295 ;
        RECT 82.715 167.260 82.945 167.705 ;
        RECT 81.335 166.565 81.950 167.085 ;
        RECT 82.120 166.585 82.350 167.015 ;
        RECT 82.535 166.765 82.945 167.260 ;
        RECT 83.115 167.440 83.905 167.705 ;
        RECT 83.115 166.585 83.370 167.440 ;
        RECT 84.185 167.375 84.355 167.755 ;
        RECT 84.570 167.545 84.900 167.925 ;
        RECT 83.540 166.765 83.925 167.245 ;
        RECT 84.185 167.205 84.900 167.375 ;
        RECT 84.095 166.655 84.450 167.025 ;
        RECT 84.730 167.015 84.900 167.205 ;
        RECT 85.070 167.180 85.325 167.755 ;
        RECT 84.730 166.685 84.985 167.015 ;
        RECT 79.970 166.055 80.665 166.365 ;
        RECT 79.975 165.375 80.660 165.845 ;
        RECT 80.840 165.645 81.145 166.430 ;
        RECT 81.335 165.375 81.595 166.385 ;
        RECT 81.765 166.215 81.935 166.565 ;
        RECT 82.120 166.415 83.910 166.585 ;
        RECT 84.730 166.475 84.900 166.685 ;
        RECT 81.765 165.545 82.040 166.215 ;
        RECT 82.240 165.375 82.455 166.220 ;
        RECT 82.680 166.120 82.930 166.415 ;
        RECT 83.155 166.055 83.485 166.245 ;
        RECT 82.640 165.545 83.115 165.885 ;
        RECT 83.295 165.880 83.485 166.055 ;
        RECT 83.655 166.050 83.910 166.415 ;
        RECT 84.185 166.305 84.900 166.475 ;
        RECT 85.155 166.450 85.325 167.180 ;
        RECT 85.500 167.085 85.760 167.925 ;
        RECT 85.935 167.175 87.145 167.925 ;
        RECT 83.295 165.375 83.925 165.880 ;
        RECT 84.185 165.545 84.355 166.305 ;
        RECT 84.570 165.375 84.900 166.135 ;
        RECT 85.070 165.545 85.325 166.450 ;
        RECT 85.500 165.375 85.760 166.525 ;
        RECT 85.935 166.465 86.455 167.005 ;
        RECT 86.625 166.635 87.145 167.175 ;
        RECT 85.935 165.375 87.145 166.465 ;
        RECT 15.930 165.205 87.230 165.375 ;
        RECT 16.015 164.115 17.225 165.205 ;
        RECT 17.395 164.115 19.985 165.205 ;
        RECT 16.015 163.405 16.535 163.945 ;
        RECT 16.705 163.575 17.225 164.115 ;
        RECT 17.395 163.425 18.605 163.945 ;
        RECT 18.775 163.595 19.985 164.115 ;
        RECT 20.155 164.445 20.670 164.855 ;
        RECT 20.905 164.445 21.075 165.205 ;
        RECT 21.245 164.865 23.275 165.035 ;
        RECT 20.155 163.635 20.495 164.445 ;
        RECT 21.245 164.200 21.415 164.865 ;
        RECT 21.810 164.525 22.935 164.695 ;
        RECT 20.665 164.010 21.415 164.200 ;
        RECT 21.585 164.185 22.595 164.355 ;
        RECT 20.155 163.465 21.385 163.635 ;
        RECT 16.015 162.655 17.225 163.405 ;
        RECT 17.395 162.655 19.985 163.425 ;
        RECT 20.430 162.860 20.675 163.465 ;
        RECT 20.895 162.655 21.405 163.190 ;
        RECT 21.585 162.825 21.775 164.185 ;
        RECT 21.945 163.845 22.220 163.985 ;
        RECT 21.945 163.675 22.225 163.845 ;
        RECT 21.945 162.825 22.220 163.675 ;
        RECT 22.425 163.385 22.595 164.185 ;
        RECT 22.765 163.395 22.935 164.525 ;
        RECT 23.105 163.895 23.275 164.865 ;
        RECT 23.445 164.065 23.615 165.205 ;
        RECT 23.785 164.065 24.120 165.035 ;
        RECT 24.295 164.115 26.885 165.205 ;
        RECT 23.105 163.565 23.300 163.895 ;
        RECT 23.525 163.565 23.780 163.895 ;
        RECT 23.525 163.395 23.695 163.565 ;
        RECT 23.950 163.395 24.120 164.065 ;
        RECT 22.765 163.225 23.695 163.395 ;
        RECT 22.765 163.190 22.940 163.225 ;
        RECT 22.410 162.825 22.940 163.190 ;
        RECT 23.365 162.655 23.695 163.055 ;
        RECT 23.865 162.825 24.120 163.395 ;
        RECT 24.295 163.425 25.505 163.945 ;
        RECT 25.675 163.595 26.885 164.115 ;
        RECT 27.515 164.065 27.775 165.205 ;
        RECT 27.945 164.055 28.275 165.035 ;
        RECT 28.445 164.065 28.725 165.205 ;
        RECT 27.535 163.645 27.870 163.895 ;
        RECT 28.040 163.455 28.210 164.055 ;
        RECT 28.895 164.040 29.185 165.205 ;
        RECT 29.355 164.025 29.675 165.205 ;
        RECT 29.845 164.185 30.045 164.975 ;
        RECT 30.370 164.375 30.755 165.035 ;
        RECT 31.150 164.445 31.935 165.205 ;
        RECT 30.345 164.275 30.755 164.375 ;
        RECT 29.845 164.015 30.175 164.185 ;
        RECT 30.345 164.065 31.955 164.275 ;
        RECT 29.995 163.895 30.175 164.015 ;
        RECT 28.380 163.625 28.715 163.895 ;
        RECT 29.355 163.645 29.820 163.845 ;
        RECT 29.995 163.645 30.325 163.895 ;
        RECT 30.495 163.845 30.960 163.895 ;
        RECT 30.495 163.675 30.965 163.845 ;
        RECT 30.495 163.645 30.960 163.675 ;
        RECT 31.155 163.645 31.510 163.895 ;
        RECT 31.680 163.465 31.955 164.065 ;
        RECT 24.295 162.655 26.885 163.425 ;
        RECT 27.515 162.825 28.210 163.455 ;
        RECT 28.415 162.655 28.725 163.455 ;
        RECT 28.895 162.655 29.185 163.380 ;
        RECT 29.355 163.265 30.535 163.435 ;
        RECT 29.355 162.850 29.695 163.265 ;
        RECT 29.865 162.655 30.035 163.095 ;
        RECT 30.205 163.045 30.535 163.265 ;
        RECT 30.705 163.285 31.955 163.465 ;
        RECT 30.705 163.215 31.070 163.285 ;
        RECT 30.205 162.865 31.455 163.045 ;
        RECT 31.725 162.655 31.895 163.115 ;
        RECT 32.125 162.935 32.405 165.035 ;
        RECT 33.040 164.065 33.375 165.035 ;
        RECT 33.545 164.065 33.715 165.205 ;
        RECT 33.885 164.865 35.915 165.035 ;
        RECT 33.040 163.395 33.210 164.065 ;
        RECT 33.885 163.895 34.055 164.865 ;
        RECT 33.380 163.565 33.635 163.895 ;
        RECT 33.860 163.565 34.055 163.895 ;
        RECT 34.225 164.525 35.350 164.695 ;
        RECT 33.465 163.395 33.635 163.565 ;
        RECT 34.225 163.395 34.395 164.525 ;
        RECT 33.040 162.825 33.295 163.395 ;
        RECT 33.465 163.225 34.395 163.395 ;
        RECT 34.565 164.185 35.575 164.355 ;
        RECT 34.565 163.385 34.735 164.185 ;
        RECT 34.220 163.190 34.395 163.225 ;
        RECT 33.465 162.655 33.795 163.055 ;
        RECT 34.220 162.825 34.750 163.190 ;
        RECT 34.940 163.165 35.215 163.985 ;
        RECT 34.935 162.995 35.215 163.165 ;
        RECT 34.940 162.825 35.215 162.995 ;
        RECT 35.385 162.825 35.575 164.185 ;
        RECT 35.745 164.200 35.915 164.865 ;
        RECT 36.085 164.445 36.255 165.205 ;
        RECT 36.490 164.445 37.005 164.855 ;
        RECT 35.745 164.010 36.495 164.200 ;
        RECT 36.665 163.635 37.005 164.445 ;
        RECT 37.175 164.065 37.435 165.205 ;
        RECT 37.605 164.055 37.935 165.035 ;
        RECT 38.105 164.065 38.385 165.205 ;
        RECT 38.555 164.115 41.145 165.205 ;
        RECT 37.195 163.645 37.530 163.895 ;
        RECT 35.775 163.465 37.005 163.635 ;
        RECT 35.755 162.655 36.265 163.190 ;
        RECT 36.485 162.860 36.730 163.465 ;
        RECT 37.700 163.455 37.870 164.055 ;
        RECT 38.040 163.625 38.375 163.895 ;
        RECT 37.175 162.825 37.870 163.455 ;
        RECT 38.075 162.655 38.385 163.455 ;
        RECT 38.555 163.425 39.765 163.945 ;
        RECT 39.935 163.595 41.145 164.115 ;
        RECT 41.320 164.255 41.585 165.025 ;
        RECT 41.755 164.485 42.085 165.205 ;
        RECT 42.275 164.665 42.535 165.025 ;
        RECT 42.705 164.835 43.035 165.205 ;
        RECT 43.205 164.665 43.465 165.025 ;
        RECT 42.275 164.435 43.465 164.665 ;
        RECT 44.035 164.255 44.325 165.025 ;
        RECT 44.535 164.770 49.880 165.205 ;
        RECT 38.555 162.655 41.145 163.425 ;
        RECT 41.320 162.835 41.655 164.255 ;
        RECT 41.830 164.075 44.325 164.255 ;
        RECT 41.830 163.385 42.055 164.075 ;
        RECT 42.255 163.565 42.535 163.895 ;
        RECT 42.715 163.565 43.290 163.895 ;
        RECT 43.470 163.565 43.905 163.895 ;
        RECT 44.085 163.565 44.355 163.895 ;
        RECT 41.830 163.195 44.315 163.385 ;
        RECT 46.120 163.200 46.460 164.030 ;
        RECT 47.940 163.520 48.290 164.770 ;
        RECT 50.055 164.115 53.565 165.205 ;
        RECT 50.055 163.425 51.705 163.945 ;
        RECT 51.875 163.595 53.565 164.115 ;
        RECT 54.655 164.040 54.945 165.205 ;
        RECT 55.115 164.065 55.390 165.035 ;
        RECT 55.600 164.405 55.880 165.205 ;
        RECT 56.050 164.695 57.665 165.025 ;
        RECT 56.050 164.355 57.225 164.525 ;
        RECT 56.050 164.235 56.220 164.355 ;
        RECT 55.560 164.065 56.220 164.235 ;
        RECT 41.835 162.655 42.580 163.025 ;
        RECT 43.145 162.835 43.400 163.195 ;
        RECT 43.580 162.655 43.910 163.025 ;
        RECT 44.090 162.835 44.315 163.195 ;
        RECT 44.535 162.655 49.880 163.200 ;
        RECT 50.055 162.655 53.565 163.425 ;
        RECT 54.655 162.655 54.945 163.380 ;
        RECT 55.115 163.330 55.285 164.065 ;
        RECT 55.560 163.895 55.730 164.065 ;
        RECT 56.480 163.895 56.725 164.185 ;
        RECT 56.895 164.065 57.225 164.355 ;
        RECT 57.485 163.895 57.655 164.455 ;
        RECT 57.905 164.065 58.165 165.205 ;
        RECT 58.335 164.770 63.680 165.205 ;
        RECT 55.455 163.565 55.730 163.895 ;
        RECT 55.900 163.565 56.725 163.895 ;
        RECT 56.940 163.565 57.655 163.895 ;
        RECT 57.825 163.645 58.160 163.895 ;
        RECT 55.560 163.395 55.730 163.565 ;
        RECT 57.405 163.475 57.655 163.565 ;
        RECT 55.115 162.985 55.390 163.330 ;
        RECT 55.560 163.225 57.225 163.395 ;
        RECT 55.580 162.655 55.955 163.055 ;
        RECT 56.125 162.875 56.295 163.225 ;
        RECT 56.465 162.655 56.795 163.055 ;
        RECT 56.965 162.825 57.225 163.225 ;
        RECT 57.405 163.055 57.735 163.475 ;
        RECT 57.905 162.655 58.165 163.475 ;
        RECT 59.920 163.200 60.260 164.030 ;
        RECT 61.740 163.520 62.090 164.770 ;
        RECT 63.855 164.115 67.365 165.205 ;
        RECT 67.535 164.115 68.745 165.205 ;
        RECT 63.855 163.425 65.505 163.945 ;
        RECT 65.675 163.595 67.365 164.115 ;
        RECT 58.335 162.655 63.680 163.200 ;
        RECT 63.855 162.655 67.365 163.425 ;
        RECT 67.535 163.405 68.055 163.945 ;
        RECT 68.225 163.575 68.745 164.115 ;
        RECT 67.535 162.655 68.745 163.405 ;
        RECT 68.915 162.825 69.665 165.035 ;
        RECT 69.835 164.650 70.440 165.205 ;
        RECT 70.615 164.695 71.095 165.035 ;
        RECT 71.265 164.660 71.520 165.205 ;
        RECT 69.835 164.550 70.450 164.650 ;
        RECT 70.265 164.525 70.450 164.550 ;
        RECT 69.835 163.930 70.095 164.380 ;
        RECT 70.265 164.280 70.595 164.525 ;
        RECT 70.765 164.205 71.520 164.455 ;
        RECT 71.690 164.335 71.965 165.035 ;
        RECT 70.750 164.170 71.520 164.205 ;
        RECT 70.735 164.160 71.520 164.170 ;
        RECT 70.730 164.145 71.625 164.160 ;
        RECT 70.710 164.130 71.625 164.145 ;
        RECT 70.690 164.120 71.625 164.130 ;
        RECT 70.665 164.110 71.625 164.120 ;
        RECT 70.595 164.080 71.625 164.110 ;
        RECT 70.575 164.050 71.625 164.080 ;
        RECT 70.555 164.020 71.625 164.050 ;
        RECT 70.525 163.995 71.625 164.020 ;
        RECT 70.490 163.960 71.625 163.995 ;
        RECT 70.460 163.955 71.625 163.960 ;
        RECT 70.460 163.950 70.850 163.955 ;
        RECT 70.460 163.940 70.825 163.950 ;
        RECT 70.460 163.935 70.810 163.940 ;
        RECT 70.460 163.930 70.795 163.935 ;
        RECT 69.835 163.925 70.795 163.930 ;
        RECT 69.835 163.915 70.785 163.925 ;
        RECT 69.835 163.910 70.775 163.915 ;
        RECT 69.835 163.900 70.765 163.910 ;
        RECT 69.835 163.890 70.760 163.900 ;
        RECT 69.835 163.885 70.755 163.890 ;
        RECT 69.835 163.870 70.745 163.885 ;
        RECT 69.835 163.855 70.740 163.870 ;
        RECT 69.835 163.830 70.730 163.855 ;
        RECT 69.835 163.760 70.725 163.830 ;
        RECT 69.835 163.205 70.385 163.590 ;
        RECT 70.555 163.035 70.725 163.760 ;
        RECT 69.835 162.865 70.725 163.035 ;
        RECT 70.895 163.360 71.225 163.785 ;
        RECT 71.395 163.560 71.625 163.955 ;
        RECT 70.895 162.875 71.115 163.360 ;
        RECT 71.795 163.305 71.965 164.335 ;
        RECT 72.145 164.065 72.475 165.205 ;
        RECT 73.005 164.235 73.335 165.020 ;
        RECT 72.655 164.065 73.335 164.235 ;
        RECT 74.055 164.275 74.235 165.035 ;
        RECT 74.415 164.445 74.745 165.205 ;
        RECT 74.055 164.105 74.730 164.275 ;
        RECT 74.915 164.130 75.185 165.035 ;
        RECT 75.355 164.695 76.545 164.985 ;
        RECT 72.135 163.645 72.485 163.895 ;
        RECT 72.655 163.465 72.825 164.065 ;
        RECT 74.560 163.960 74.730 164.105 ;
        RECT 72.995 163.645 73.345 163.895 ;
        RECT 73.995 163.555 74.335 163.925 ;
        RECT 74.560 163.630 74.835 163.960 ;
        RECT 71.285 162.655 71.535 163.195 ;
        RECT 71.705 162.825 71.965 163.305 ;
        RECT 72.145 162.655 72.415 163.465 ;
        RECT 72.585 162.825 72.915 163.465 ;
        RECT 73.085 162.655 73.325 163.465 ;
        RECT 74.560 163.375 74.730 163.630 ;
        RECT 74.065 163.205 74.730 163.375 ;
        RECT 75.005 163.330 75.185 164.130 ;
        RECT 75.375 164.355 76.545 164.525 ;
        RECT 76.715 164.405 76.995 165.205 ;
        RECT 75.375 164.065 75.700 164.355 ;
        RECT 76.375 164.235 76.545 164.355 ;
        RECT 75.870 163.895 76.065 164.185 ;
        RECT 76.375 164.065 77.035 164.235 ;
        RECT 77.205 164.065 77.480 165.035 ;
        RECT 78.155 164.865 79.295 165.035 ;
        RECT 78.155 164.405 78.455 164.865 ;
        RECT 78.625 164.235 78.955 164.695 ;
        RECT 78.195 164.185 78.955 164.235 ;
        RECT 76.865 163.895 77.035 164.065 ;
        RECT 75.355 163.565 75.700 163.895 ;
        RECT 75.870 163.565 76.695 163.895 ;
        RECT 76.865 163.565 77.140 163.895 ;
        RECT 76.865 163.395 77.035 163.565 ;
        RECT 74.065 162.825 74.235 163.205 ;
        RECT 74.415 162.655 74.745 163.035 ;
        RECT 74.925 162.825 75.185 163.330 ;
        RECT 75.370 163.225 77.035 163.395 ;
        RECT 77.310 163.330 77.480 164.065 ;
        RECT 78.175 164.015 78.955 164.185 ;
        RECT 79.125 164.235 79.295 164.865 ;
        RECT 79.465 164.405 79.795 165.205 ;
        RECT 79.965 164.235 80.240 165.035 ;
        RECT 79.125 164.025 80.240 164.235 ;
        RECT 80.415 164.040 80.705 165.205 ;
        RECT 80.915 164.065 81.145 165.205 ;
        RECT 81.315 164.055 81.645 165.035 ;
        RECT 81.815 164.065 82.025 165.205 ;
        RECT 82.385 164.865 84.435 165.035 ;
        RECT 82.385 164.365 82.635 164.865 ;
        RECT 82.805 164.195 83.015 164.695 ;
        RECT 83.225 164.365 83.435 164.865 ;
        RECT 83.765 164.195 84.015 164.695 ;
        RECT 84.185 164.365 84.435 164.865 ;
        RECT 84.605 164.195 84.855 165.035 ;
        RECT 85.025 164.365 85.275 165.205 ;
        RECT 85.445 164.195 85.700 165.035 ;
        RECT 75.370 162.875 75.625 163.225 ;
        RECT 75.795 162.655 76.125 163.055 ;
        RECT 76.295 162.875 76.465 163.225 ;
        RECT 76.635 162.655 77.015 163.055 ;
        RECT 77.205 162.985 77.480 163.330 ;
        RECT 78.195 163.475 78.410 164.015 ;
        RECT 78.580 163.645 79.350 163.845 ;
        RECT 79.520 163.645 80.240 163.845 ;
        RECT 80.895 163.645 81.225 163.895 ;
        RECT 78.195 163.305 79.795 163.475 ;
        RECT 78.625 163.295 79.795 163.305 ;
        RECT 78.165 162.655 78.455 163.125 ;
        RECT 78.625 162.825 78.955 163.295 ;
        RECT 79.125 162.655 79.295 163.125 ;
        RECT 79.465 162.825 79.795 163.295 ;
        RECT 79.965 162.655 80.240 163.475 ;
        RECT 80.415 162.655 80.705 163.380 ;
        RECT 80.915 162.655 81.145 163.475 ;
        RECT 81.395 163.455 81.645 164.055 ;
        RECT 82.255 164.025 83.015 164.195 ;
        RECT 82.255 163.475 82.715 164.025 ;
        RECT 83.210 163.855 83.475 164.195 ;
        RECT 83.765 164.025 85.700 164.195 ;
        RECT 85.935 164.115 87.145 165.205 ;
        RECT 82.885 163.645 83.475 163.855 ;
        RECT 83.665 163.645 84.715 163.855 ;
        RECT 84.885 163.645 85.715 163.855 ;
        RECT 85.935 163.575 86.455 164.115 ;
        RECT 81.315 162.825 81.645 163.455 ;
        RECT 81.815 162.655 82.025 163.475 ;
        RECT 82.255 163.295 85.315 163.475 ;
        RECT 82.305 162.655 82.595 163.125 ;
        RECT 82.765 162.825 83.095 163.295 ;
        RECT 83.265 162.655 83.975 163.125 ;
        RECT 84.145 162.825 84.475 163.295 ;
        RECT 84.645 162.655 84.815 163.125 ;
        RECT 84.985 162.825 85.315 163.295 ;
        RECT 85.485 162.655 85.760 163.475 ;
        RECT 86.625 163.405 87.145 163.945 ;
        RECT 85.935 162.655 87.145 163.405 ;
        RECT 15.930 162.485 87.230 162.655 ;
        RECT 16.015 161.735 17.225 162.485 ;
        RECT 16.015 161.195 16.535 161.735 ;
        RECT 17.400 161.645 17.660 162.485 ;
        RECT 17.835 161.740 18.090 162.315 ;
        RECT 18.260 162.105 18.590 162.485 ;
        RECT 18.805 161.935 18.975 162.315 ;
        RECT 18.260 161.765 18.975 161.935 ;
        RECT 19.235 161.985 19.495 162.315 ;
        RECT 19.705 162.005 19.980 162.485 ;
        RECT 16.705 161.025 17.225 161.565 ;
        RECT 16.015 159.935 17.225 161.025 ;
        RECT 17.400 159.935 17.660 161.085 ;
        RECT 17.835 161.010 18.005 161.740 ;
        RECT 18.260 161.575 18.430 161.765 ;
        RECT 18.175 161.245 18.430 161.575 ;
        RECT 18.260 161.035 18.430 161.245 ;
        RECT 18.710 161.215 19.065 161.585 ;
        RECT 19.235 161.075 19.405 161.985 ;
        RECT 20.190 161.915 20.395 162.315 ;
        RECT 20.565 162.085 20.900 162.485 ;
        RECT 19.575 161.245 19.935 161.825 ;
        RECT 20.190 161.745 20.875 161.915 ;
        RECT 20.115 161.075 20.365 161.575 ;
        RECT 17.835 160.105 18.090 161.010 ;
        RECT 18.260 160.865 18.975 161.035 ;
        RECT 18.260 159.935 18.590 160.695 ;
        RECT 18.805 160.105 18.975 160.865 ;
        RECT 19.235 160.905 20.365 161.075 ;
        RECT 19.235 160.135 19.505 160.905 ;
        RECT 20.535 160.715 20.875 161.745 ;
        RECT 19.675 159.935 20.005 160.715 ;
        RECT 20.210 160.540 20.875 160.715 ;
        RECT 21.075 161.810 21.335 162.315 ;
        RECT 21.515 162.105 21.845 162.485 ;
        RECT 22.025 161.935 22.195 162.315 ;
        RECT 22.455 161.940 27.800 162.485 ;
        RECT 21.075 161.010 21.245 161.810 ;
        RECT 21.530 161.765 22.195 161.935 ;
        RECT 21.530 161.510 21.700 161.765 ;
        RECT 21.415 161.180 21.700 161.510 ;
        RECT 21.935 161.215 22.265 161.585 ;
        RECT 21.530 161.035 21.700 161.180 ;
        RECT 24.040 161.110 24.380 161.940 ;
        RECT 28.495 161.665 28.705 162.485 ;
        RECT 28.875 161.685 29.205 162.315 ;
        RECT 20.210 160.135 20.395 160.540 ;
        RECT 20.565 159.935 20.900 160.360 ;
        RECT 21.075 160.105 21.345 161.010 ;
        RECT 21.530 160.865 22.195 161.035 ;
        RECT 21.515 159.935 21.845 160.695 ;
        RECT 22.025 160.105 22.195 160.865 ;
        RECT 25.860 160.370 26.210 161.620 ;
        RECT 28.875 161.085 29.125 161.685 ;
        RECT 29.375 161.665 29.605 162.485 ;
        RECT 30.015 161.855 30.345 162.215 ;
        RECT 30.975 162.025 31.225 162.485 ;
        RECT 31.395 162.025 31.945 162.315 ;
        RECT 30.015 161.665 31.405 161.855 ;
        RECT 31.235 161.575 31.405 161.665 ;
        RECT 29.295 161.245 29.625 161.495 ;
        RECT 29.815 161.245 30.505 161.495 ;
        RECT 30.735 161.245 31.065 161.495 ;
        RECT 31.235 161.245 31.525 161.575 ;
        RECT 22.455 159.935 27.800 160.370 ;
        RECT 28.495 159.935 28.705 161.075 ;
        RECT 28.875 160.105 29.205 161.085 ;
        RECT 29.375 159.935 29.605 161.075 ;
        RECT 29.815 160.805 30.130 161.245 ;
        RECT 31.235 160.995 31.405 161.245 ;
        RECT 30.465 160.825 31.405 160.995 ;
        RECT 30.015 159.935 30.295 160.605 ;
        RECT 30.465 160.275 30.765 160.825 ;
        RECT 31.695 160.655 31.945 162.025 ;
        RECT 32.115 161.685 32.405 162.485 ;
        RECT 32.580 161.745 32.835 162.315 ;
        RECT 33.005 162.085 33.335 162.485 ;
        RECT 33.760 161.950 34.290 162.315 ;
        RECT 33.760 161.915 33.935 161.950 ;
        RECT 33.005 161.745 33.935 161.915 ;
        RECT 32.580 161.075 32.750 161.745 ;
        RECT 33.005 161.575 33.175 161.745 ;
        RECT 32.920 161.245 33.175 161.575 ;
        RECT 33.400 161.245 33.595 161.575 ;
        RECT 30.975 159.935 31.305 160.655 ;
        RECT 31.495 160.105 31.945 160.655 ;
        RECT 32.115 159.935 32.405 161.075 ;
        RECT 32.580 160.105 32.915 161.075 ;
        RECT 33.085 159.935 33.255 161.075 ;
        RECT 33.425 160.275 33.595 161.245 ;
        RECT 33.765 160.615 33.935 161.745 ;
        RECT 34.105 160.955 34.275 161.755 ;
        RECT 34.480 161.465 34.755 162.315 ;
        RECT 34.475 161.295 34.755 161.465 ;
        RECT 34.480 161.155 34.755 161.295 ;
        RECT 34.925 160.955 35.115 162.315 ;
        RECT 35.295 161.950 35.805 162.485 ;
        RECT 36.025 161.675 36.270 162.280 ;
        RECT 36.715 161.715 38.385 162.485 ;
        RECT 38.720 161.975 38.960 162.485 ;
        RECT 39.140 161.975 39.420 162.305 ;
        RECT 39.650 161.975 39.865 162.485 ;
        RECT 35.315 161.505 36.545 161.675 ;
        RECT 34.105 160.785 35.115 160.955 ;
        RECT 35.285 160.940 36.035 161.130 ;
        RECT 33.765 160.445 34.890 160.615 ;
        RECT 35.285 160.275 35.455 160.940 ;
        RECT 36.205 160.695 36.545 161.505 ;
        RECT 36.715 161.195 37.465 161.715 ;
        RECT 37.635 161.025 38.385 161.545 ;
        RECT 38.615 161.245 38.970 161.805 ;
        RECT 39.140 161.075 39.310 161.975 ;
        RECT 39.480 161.245 39.745 161.805 ;
        RECT 40.035 161.745 40.650 162.315 ;
        RECT 41.775 161.760 42.065 162.485 ;
        RECT 39.995 161.075 40.165 161.575 ;
        RECT 33.425 160.105 35.455 160.275 ;
        RECT 35.625 159.935 35.795 160.695 ;
        RECT 36.030 160.285 36.545 160.695 ;
        RECT 36.715 159.935 38.385 161.025 ;
        RECT 38.740 160.905 40.165 161.075 ;
        RECT 38.740 160.730 39.130 160.905 ;
        RECT 39.615 159.935 39.945 160.735 ;
        RECT 40.335 160.725 40.650 161.745 ;
        RECT 42.235 161.665 42.920 162.305 ;
        RECT 43.090 161.665 43.260 162.485 ;
        RECT 43.430 161.835 43.760 162.300 ;
        RECT 43.930 162.015 44.100 162.485 ;
        RECT 44.360 162.095 45.545 162.265 ;
        RECT 45.715 161.925 46.045 162.315 ;
        RECT 44.745 161.835 45.130 161.925 ;
        RECT 43.430 161.665 45.130 161.835 ;
        RECT 45.535 161.745 46.045 161.925 ;
        RECT 46.385 161.765 46.715 162.485 ;
        RECT 47.260 162.085 48.875 162.255 ;
        RECT 49.045 162.085 49.375 162.485 ;
        RECT 48.705 161.915 48.875 162.085 ;
        RECT 49.545 162.010 49.880 162.270 ;
        RECT 40.115 160.105 40.650 160.725 ;
        RECT 41.775 159.935 42.065 161.100 ;
        RECT 42.235 160.695 42.485 161.665 ;
        RECT 42.655 161.285 42.990 161.495 ;
        RECT 43.160 161.285 43.610 161.495 ;
        RECT 43.800 161.285 44.285 161.495 ;
        RECT 42.820 161.115 42.990 161.285 ;
        RECT 43.910 161.125 44.285 161.285 ;
        RECT 44.475 161.245 44.855 161.495 ;
        RECT 45.035 161.285 45.365 161.495 ;
        RECT 42.820 160.945 43.740 161.115 ;
        RECT 42.235 160.105 42.900 160.695 ;
        RECT 43.070 159.935 43.400 160.775 ;
        RECT 43.570 160.695 43.740 160.945 ;
        RECT 43.910 160.955 44.305 161.125 ;
        RECT 43.910 160.865 44.285 160.955 ;
        RECT 44.475 160.865 44.795 161.245 ;
        RECT 45.535 161.115 45.705 161.745 ;
        RECT 45.875 161.285 46.205 161.575 ;
        RECT 46.440 161.465 46.790 161.575 ;
        RECT 46.435 161.295 46.790 161.465 ;
        RECT 46.440 161.245 46.790 161.295 ;
        RECT 47.100 161.245 47.520 161.910 ;
        RECT 47.690 161.805 47.980 161.905 ;
        RECT 48.170 161.805 48.440 161.905 ;
        RECT 47.690 161.635 47.985 161.805 ;
        RECT 48.170 161.635 48.445 161.805 ;
        RECT 48.705 161.745 49.265 161.915 ;
        RECT 47.690 161.245 47.980 161.635 ;
        RECT 48.170 161.245 48.440 161.635 ;
        RECT 49.095 161.575 49.265 161.745 ;
        RECT 48.650 161.465 48.900 161.575 ;
        RECT 48.650 161.295 48.905 161.465 ;
        RECT 48.650 161.245 48.900 161.295 ;
        RECT 49.095 161.245 49.400 161.575 ;
        RECT 44.965 160.945 46.050 161.115 ;
        RECT 46.440 160.955 46.645 161.245 ;
        RECT 49.095 161.075 49.265 161.245 ;
        RECT 44.965 160.695 45.135 160.945 ;
        RECT 43.570 160.525 45.135 160.695 ;
        RECT 43.910 160.105 44.715 160.525 ;
        RECT 45.305 159.935 45.555 160.775 ;
        RECT 45.750 160.105 46.050 160.945 ;
        RECT 46.895 160.905 49.265 161.075 ;
        RECT 46.465 160.275 46.635 160.775 ;
        RECT 46.895 160.445 47.065 160.905 ;
        RECT 47.295 160.525 48.720 160.695 ;
        RECT 47.295 160.275 47.625 160.525 ;
        RECT 46.465 160.105 47.625 160.275 ;
        RECT 47.850 159.935 48.180 160.355 ;
        RECT 48.435 160.105 48.720 160.525 ;
        RECT 48.965 159.935 49.295 160.735 ;
        RECT 49.625 160.655 49.880 162.010 ;
        RECT 50.060 161.720 50.515 162.485 ;
        RECT 50.790 162.105 52.090 162.315 ;
        RECT 52.345 162.125 52.675 162.485 ;
        RECT 51.920 161.955 52.090 162.105 ;
        RECT 52.845 161.985 53.105 162.315 ;
        RECT 52.875 161.975 53.105 161.985 ;
        RECT 50.990 161.495 51.210 161.895 ;
        RECT 50.055 161.295 50.545 161.495 ;
        RECT 50.735 161.285 51.210 161.495 ;
        RECT 51.455 161.495 51.665 161.895 ;
        RECT 51.920 161.830 52.675 161.955 ;
        RECT 51.920 161.785 52.765 161.830 ;
        RECT 52.495 161.665 52.765 161.785 ;
        RECT 51.455 161.285 51.785 161.495 ;
        RECT 51.955 161.225 52.365 161.530 ;
        RECT 49.545 160.145 49.880 160.655 ;
        RECT 50.060 161.055 51.235 161.115 ;
        RECT 52.595 161.090 52.765 161.665 ;
        RECT 52.565 161.055 52.765 161.090 ;
        RECT 50.060 160.945 52.765 161.055 ;
        RECT 50.060 160.325 50.315 160.945 ;
        RECT 50.905 160.885 52.705 160.945 ;
        RECT 50.905 160.855 51.235 160.885 ;
        RECT 52.935 160.785 53.105 161.975 ;
        RECT 53.275 161.940 58.620 162.485 ;
        RECT 54.860 161.110 55.200 161.940 ;
        RECT 58.805 161.890 59.055 162.315 ;
        RECT 59.225 162.060 59.555 162.485 ;
        RECT 59.725 162.065 60.815 162.315 ;
        RECT 61.005 162.065 62.095 162.315 ;
        RECT 59.725 161.890 59.895 162.065 ;
        RECT 58.805 161.720 59.895 161.890 ;
        RECT 60.065 161.725 61.755 161.895 ;
        RECT 61.925 161.890 62.095 162.065 ;
        RECT 62.265 162.060 62.595 162.485 ;
        RECT 62.765 161.890 63.085 162.315 ;
        RECT 50.565 160.685 50.750 160.775 ;
        RECT 51.340 160.685 52.175 160.695 ;
        RECT 50.565 160.485 52.175 160.685 ;
        RECT 50.565 160.445 50.795 160.485 ;
        RECT 50.060 160.105 50.395 160.325 ;
        RECT 51.400 159.935 51.755 160.315 ;
        RECT 51.925 160.105 52.175 160.485 ;
        RECT 52.425 159.935 52.675 160.715 ;
        RECT 52.845 160.105 53.105 160.785 ;
        RECT 56.680 160.370 57.030 161.620 ;
        RECT 58.860 161.465 59.490 161.495 ;
        RECT 59.780 161.465 60.410 161.495 ;
        RECT 58.855 161.295 59.490 161.465 ;
        RECT 59.775 161.295 60.410 161.465 ;
        RECT 60.580 161.085 60.870 161.725 ;
        RECT 61.925 161.720 63.085 161.890 ;
        RECT 63.415 161.755 63.705 162.485 ;
        RECT 61.155 161.295 61.810 161.495 ;
        RECT 62.100 161.465 63.210 161.495 ;
        RECT 62.075 161.295 63.210 161.465 ;
        RECT 63.405 161.245 63.705 161.575 ;
        RECT 63.885 161.555 64.115 162.195 ;
        RECT 64.295 161.935 64.605 162.305 ;
        RECT 64.785 162.115 65.455 162.485 ;
        RECT 64.295 161.735 65.525 161.935 ;
        RECT 63.885 161.245 64.410 161.555 ;
        RECT 64.590 161.245 65.055 161.555 ;
        RECT 58.805 160.915 60.870 161.085 ;
        RECT 53.275 159.935 58.620 160.370 ;
        RECT 58.805 160.105 59.055 160.915 ;
        RECT 59.225 160.275 59.475 160.745 ;
        RECT 59.645 160.445 59.975 160.915 ;
        RECT 60.145 160.275 60.315 160.745 ;
        RECT 60.485 160.445 60.870 160.915 ;
        RECT 61.085 160.915 63.015 161.085 ;
        RECT 65.235 161.065 65.525 161.735 ;
        RECT 61.085 160.275 61.335 160.915 ;
        RECT 59.225 160.105 61.335 160.275 ;
        RECT 61.505 159.935 61.675 160.745 ;
        RECT 61.845 160.105 62.175 160.915 ;
        RECT 62.345 159.935 62.515 160.745 ;
        RECT 62.685 160.105 63.015 160.915 ;
        RECT 63.415 160.825 64.575 161.065 ;
        RECT 63.415 160.115 63.675 160.825 ;
        RECT 63.845 159.935 64.175 160.645 ;
        RECT 64.345 160.115 64.575 160.825 ;
        RECT 64.755 160.845 65.525 161.065 ;
        RECT 64.755 160.115 65.025 160.845 ;
        RECT 65.205 159.935 65.545 160.665 ;
        RECT 65.715 160.115 65.975 162.305 ;
        RECT 66.155 161.735 67.365 162.485 ;
        RECT 67.535 161.760 67.825 162.485 ;
        RECT 66.155 161.195 66.675 161.735 ;
        RECT 66.845 161.025 67.365 161.565 ;
        RECT 66.155 159.935 67.365 161.025 ;
        RECT 67.535 159.935 67.825 161.100 ;
        RECT 67.995 160.105 68.275 162.205 ;
        RECT 68.505 162.025 68.675 162.485 ;
        RECT 68.945 162.095 70.195 162.275 ;
        RECT 69.330 161.855 69.695 161.925 ;
        RECT 68.445 161.675 69.695 161.855 ;
        RECT 69.865 161.875 70.195 162.095 ;
        RECT 70.365 162.045 70.535 162.485 ;
        RECT 70.705 161.875 71.045 162.290 ;
        RECT 71.215 162.105 72.105 162.275 ;
        RECT 69.865 161.705 71.045 161.875 ;
        RECT 68.445 161.075 68.720 161.675 ;
        RECT 71.215 161.550 71.765 161.935 ;
        RECT 68.890 161.245 69.245 161.495 ;
        RECT 69.440 161.465 69.905 161.495 ;
        RECT 69.435 161.295 69.905 161.465 ;
        RECT 69.440 161.245 69.905 161.295 ;
        RECT 70.075 161.245 70.405 161.495 ;
        RECT 70.580 161.295 71.045 161.495 ;
        RECT 71.935 161.380 72.105 162.105 ;
        RECT 71.215 161.310 72.105 161.380 ;
        RECT 72.275 161.780 72.495 162.265 ;
        RECT 72.665 161.945 72.915 162.485 ;
        RECT 73.085 161.835 73.345 162.315 ;
        RECT 73.515 162.105 74.405 162.275 ;
        RECT 72.275 161.355 72.605 161.780 ;
        RECT 70.225 161.125 70.405 161.245 ;
        RECT 71.215 161.285 72.110 161.310 ;
        RECT 71.215 161.270 72.120 161.285 ;
        RECT 71.215 161.255 72.125 161.270 ;
        RECT 71.215 161.250 72.135 161.255 ;
        RECT 71.215 161.240 72.140 161.250 ;
        RECT 71.215 161.230 72.145 161.240 ;
        RECT 71.215 161.225 72.155 161.230 ;
        RECT 71.215 161.215 72.165 161.225 ;
        RECT 71.215 161.210 72.175 161.215 ;
        RECT 68.445 160.865 70.055 161.075 ;
        RECT 70.225 160.955 70.555 161.125 ;
        RECT 69.645 160.765 70.055 160.865 ;
        RECT 68.465 159.935 69.250 160.695 ;
        RECT 69.645 160.105 70.030 160.765 ;
        RECT 70.355 160.165 70.555 160.955 ;
        RECT 70.725 159.935 71.045 161.115 ;
        RECT 71.215 160.760 71.475 161.210 ;
        RECT 71.840 161.205 72.175 161.210 ;
        RECT 71.840 161.200 72.190 161.205 ;
        RECT 71.840 161.190 72.205 161.200 ;
        RECT 71.840 161.185 72.230 161.190 ;
        RECT 72.775 161.185 73.005 161.580 ;
        RECT 71.840 161.180 73.005 161.185 ;
        RECT 71.870 161.145 73.005 161.180 ;
        RECT 71.905 161.120 73.005 161.145 ;
        RECT 71.935 161.090 73.005 161.120 ;
        RECT 71.955 161.060 73.005 161.090 ;
        RECT 71.975 161.030 73.005 161.060 ;
        RECT 72.045 161.020 73.005 161.030 ;
        RECT 72.070 161.010 73.005 161.020 ;
        RECT 72.090 160.995 73.005 161.010 ;
        RECT 72.110 160.980 73.005 160.995 ;
        RECT 72.115 160.970 72.900 160.980 ;
        RECT 72.130 160.935 72.900 160.970 ;
        RECT 71.645 160.615 71.975 160.860 ;
        RECT 72.145 160.685 72.900 160.935 ;
        RECT 73.175 160.805 73.345 161.835 ;
        RECT 73.515 161.550 74.065 161.935 ;
        RECT 74.235 161.380 74.405 162.105 ;
        RECT 71.645 160.590 71.830 160.615 ;
        RECT 71.215 160.490 71.830 160.590 ;
        RECT 71.215 159.935 71.820 160.490 ;
        RECT 71.995 160.105 72.475 160.445 ;
        RECT 72.645 159.935 72.900 160.480 ;
        RECT 73.070 160.105 73.345 160.805 ;
        RECT 73.515 161.310 74.405 161.380 ;
        RECT 74.575 161.780 74.795 162.265 ;
        RECT 74.965 161.945 75.215 162.485 ;
        RECT 75.385 161.835 75.645 162.315 ;
        RECT 76.735 161.975 77.040 162.485 ;
        RECT 74.575 161.355 74.905 161.780 ;
        RECT 73.515 161.285 74.410 161.310 ;
        RECT 73.515 161.270 74.420 161.285 ;
        RECT 73.515 161.255 74.425 161.270 ;
        RECT 73.515 161.250 74.435 161.255 ;
        RECT 73.515 161.240 74.440 161.250 ;
        RECT 73.515 161.230 74.445 161.240 ;
        RECT 73.515 161.225 74.455 161.230 ;
        RECT 73.515 161.215 74.465 161.225 ;
        RECT 73.515 161.210 74.475 161.215 ;
        RECT 73.515 160.760 73.775 161.210 ;
        RECT 74.140 161.205 74.475 161.210 ;
        RECT 74.140 161.200 74.490 161.205 ;
        RECT 74.140 161.190 74.505 161.200 ;
        RECT 74.140 161.185 74.530 161.190 ;
        RECT 75.075 161.185 75.305 161.580 ;
        RECT 74.140 161.180 75.305 161.185 ;
        RECT 74.170 161.145 75.305 161.180 ;
        RECT 74.205 161.120 75.305 161.145 ;
        RECT 74.235 161.090 75.305 161.120 ;
        RECT 74.255 161.060 75.305 161.090 ;
        RECT 74.275 161.030 75.305 161.060 ;
        RECT 74.345 161.020 75.305 161.030 ;
        RECT 74.370 161.010 75.305 161.020 ;
        RECT 74.390 160.995 75.305 161.010 ;
        RECT 74.410 160.980 75.305 160.995 ;
        RECT 74.415 160.970 75.200 160.980 ;
        RECT 74.430 160.935 75.200 160.970 ;
        RECT 73.945 160.615 74.275 160.860 ;
        RECT 74.445 160.685 75.200 160.935 ;
        RECT 75.475 160.805 75.645 161.835 ;
        RECT 76.735 161.245 77.050 161.805 ;
        RECT 77.220 161.495 77.470 162.305 ;
        RECT 77.640 161.960 77.900 162.485 ;
        RECT 78.080 161.495 78.330 162.305 ;
        RECT 78.500 161.925 78.760 162.485 ;
        RECT 78.930 161.835 79.190 162.290 ;
        RECT 79.360 162.005 79.620 162.485 ;
        RECT 79.790 161.835 80.050 162.290 ;
        RECT 80.220 162.005 80.480 162.485 ;
        RECT 80.650 161.835 80.910 162.290 ;
        RECT 81.080 162.005 81.325 162.485 ;
        RECT 81.495 161.835 81.770 162.290 ;
        RECT 81.940 162.005 82.185 162.485 ;
        RECT 82.355 161.835 82.615 162.290 ;
        RECT 82.795 162.005 83.045 162.485 ;
        RECT 83.215 161.835 83.475 162.290 ;
        RECT 83.655 162.005 83.905 162.485 ;
        RECT 84.075 161.835 84.335 162.290 ;
        RECT 84.515 162.005 84.775 162.485 ;
        RECT 84.945 161.835 85.205 162.290 ;
        RECT 85.375 162.005 85.675 162.485 ;
        RECT 78.930 161.665 85.675 161.835 ;
        RECT 85.935 161.735 87.145 162.485 ;
        RECT 77.220 161.245 84.340 161.495 ;
        RECT 73.945 160.590 74.130 160.615 ;
        RECT 73.515 160.490 74.130 160.590 ;
        RECT 73.515 159.935 74.120 160.490 ;
        RECT 74.295 160.105 74.775 160.445 ;
        RECT 74.945 159.935 75.200 160.480 ;
        RECT 75.370 160.105 75.645 160.805 ;
        RECT 76.745 159.935 77.040 160.745 ;
        RECT 77.220 160.105 77.465 161.245 ;
        RECT 77.640 159.935 77.900 160.745 ;
        RECT 78.080 160.110 78.330 161.245 ;
        RECT 84.510 161.075 85.675 161.665 ;
        RECT 78.930 160.850 85.675 161.075 ;
        RECT 85.935 161.025 86.455 161.565 ;
        RECT 86.625 161.195 87.145 161.735 ;
        RECT 78.930 160.835 84.335 160.850 ;
        RECT 78.500 159.940 78.760 160.735 ;
        RECT 78.930 160.110 79.190 160.835 ;
        RECT 79.360 159.940 79.620 160.665 ;
        RECT 79.790 160.110 80.050 160.835 ;
        RECT 80.220 159.940 80.480 160.665 ;
        RECT 80.650 160.110 80.910 160.835 ;
        RECT 81.080 159.940 81.340 160.665 ;
        RECT 81.510 160.110 81.770 160.835 ;
        RECT 81.940 159.940 82.185 160.665 ;
        RECT 82.355 160.110 82.615 160.835 ;
        RECT 82.800 159.940 83.045 160.665 ;
        RECT 83.215 160.110 83.475 160.835 ;
        RECT 83.660 159.940 83.905 160.665 ;
        RECT 84.075 160.110 84.335 160.835 ;
        RECT 84.520 159.940 84.775 160.665 ;
        RECT 84.945 160.110 85.235 160.850 ;
        RECT 78.500 159.935 84.775 159.940 ;
        RECT 85.405 159.935 85.675 160.680 ;
        RECT 85.935 159.935 87.145 161.025 ;
        RECT 15.930 159.765 87.230 159.935 ;
        RECT 16.015 158.675 17.225 159.765 ;
        RECT 16.015 157.965 16.535 158.505 ;
        RECT 16.705 158.135 17.225 158.675 ;
        RECT 18.320 158.625 18.640 159.765 ;
        RECT 18.820 158.455 19.015 159.505 ;
        RECT 19.195 158.915 19.525 159.595 ;
        RECT 19.725 158.965 19.980 159.765 ;
        RECT 20.245 159.145 20.415 159.575 ;
        RECT 20.585 159.315 20.915 159.765 ;
        RECT 20.245 158.915 20.925 159.145 ;
        RECT 19.195 158.635 19.545 158.915 ;
        RECT 18.380 158.405 18.640 158.455 ;
        RECT 18.375 158.235 18.640 158.405 ;
        RECT 18.380 158.125 18.640 158.235 ;
        RECT 18.820 158.125 19.205 158.455 ;
        RECT 19.375 158.255 19.545 158.635 ;
        RECT 19.735 158.425 19.980 158.785 ;
        RECT 19.375 158.085 19.895 158.255 ;
        RECT 16.015 157.215 17.225 157.965 ;
        RECT 18.320 157.745 19.535 157.915 ;
        RECT 18.320 157.395 18.610 157.745 ;
        RECT 18.805 157.215 19.135 157.575 ;
        RECT 19.305 157.440 19.535 157.745 ;
        RECT 19.725 157.520 19.895 158.085 ;
        RECT 20.220 158.065 20.520 158.745 ;
        RECT 20.215 157.895 20.520 158.065 ;
        RECT 20.690 158.265 20.925 158.915 ;
        RECT 21.115 158.605 21.400 159.550 ;
        RECT 21.580 159.295 22.265 159.765 ;
        RECT 21.575 158.775 22.270 159.085 ;
        RECT 22.445 158.710 22.750 159.495 ;
        RECT 22.935 158.810 23.205 159.765 ;
        RECT 23.380 158.965 23.635 159.765 ;
        RECT 23.835 158.915 24.165 159.595 ;
        RECT 21.115 158.455 21.975 158.605 ;
        RECT 21.115 158.435 22.405 158.455 ;
        RECT 20.690 157.935 21.245 158.265 ;
        RECT 21.415 158.075 22.405 158.435 ;
        RECT 20.690 157.785 20.905 157.935 ;
        RECT 20.165 157.215 20.495 157.720 ;
        RECT 20.665 157.410 20.905 157.785 ;
        RECT 21.415 157.740 21.585 158.075 ;
        RECT 22.575 157.905 22.750 158.710 ;
        RECT 23.380 158.425 23.625 158.785 ;
        RECT 23.815 158.635 24.165 158.915 ;
        RECT 23.815 158.255 23.985 158.635 ;
        RECT 24.345 158.455 24.540 159.505 ;
        RECT 24.720 158.625 25.040 159.765 ;
        RECT 25.215 158.675 28.725 159.765 ;
        RECT 21.185 157.545 21.585 157.740 ;
        RECT 21.185 157.400 21.355 157.545 ;
        RECT 21.945 157.215 22.345 157.710 ;
        RECT 22.515 157.385 22.750 157.905 ;
        RECT 23.465 158.085 23.985 158.255 ;
        RECT 24.155 158.125 24.540 158.455 ;
        RECT 24.720 158.405 24.980 158.455 ;
        RECT 24.720 158.235 24.985 158.405 ;
        RECT 24.720 158.125 24.980 158.235 ;
        RECT 22.935 157.215 23.205 157.850 ;
        RECT 23.465 157.520 23.635 158.085 ;
        RECT 25.215 157.985 26.865 158.505 ;
        RECT 27.035 158.155 28.725 158.675 ;
        RECT 28.895 158.600 29.185 159.765 ;
        RECT 29.360 158.615 29.620 159.765 ;
        RECT 29.795 158.690 30.050 159.595 ;
        RECT 30.220 159.005 30.550 159.765 ;
        RECT 30.765 158.835 30.935 159.595 ;
        RECT 23.825 157.745 25.040 157.915 ;
        RECT 23.825 157.440 24.055 157.745 ;
        RECT 24.225 157.215 24.555 157.575 ;
        RECT 24.750 157.395 25.040 157.745 ;
        RECT 25.215 157.215 28.725 157.985 ;
        RECT 28.895 157.215 29.185 157.940 ;
        RECT 29.360 157.215 29.620 158.055 ;
        RECT 29.795 157.960 29.965 158.690 ;
        RECT 30.220 158.665 30.935 158.835 ;
        RECT 31.195 158.675 34.705 159.765 ;
        RECT 35.995 159.095 36.275 159.765 ;
        RECT 36.445 158.875 36.745 159.425 ;
        RECT 36.945 159.045 37.275 159.765 ;
        RECT 37.465 159.045 37.925 159.595 ;
        RECT 38.095 159.330 43.440 159.765 ;
        RECT 30.220 158.455 30.390 158.665 ;
        RECT 30.135 158.125 30.390 158.455 ;
        RECT 29.795 157.385 30.050 157.960 ;
        RECT 30.220 157.935 30.390 158.125 ;
        RECT 30.670 158.115 31.025 158.485 ;
        RECT 31.195 157.985 32.845 158.505 ;
        RECT 33.015 158.155 34.705 158.675 ;
        RECT 35.810 158.455 36.075 158.815 ;
        RECT 36.445 158.705 37.385 158.875 ;
        RECT 37.215 158.455 37.385 158.705 ;
        RECT 35.810 158.205 36.485 158.455 ;
        RECT 36.705 158.205 37.045 158.455 ;
        RECT 37.215 158.125 37.505 158.455 ;
        RECT 37.215 158.035 37.385 158.125 ;
        RECT 30.220 157.765 30.935 157.935 ;
        RECT 30.220 157.215 30.550 157.595 ;
        RECT 30.765 157.385 30.935 157.765 ;
        RECT 31.195 157.215 34.705 157.985 ;
        RECT 35.995 157.845 37.385 158.035 ;
        RECT 35.995 157.485 36.325 157.845 ;
        RECT 37.675 157.675 37.925 159.045 ;
        RECT 39.680 157.760 40.020 158.590 ;
        RECT 41.500 158.080 41.850 159.330 ;
        RECT 43.615 158.675 45.285 159.765 ;
        RECT 43.615 157.985 44.365 158.505 ;
        RECT 44.535 158.155 45.285 158.675 ;
        RECT 45.455 158.160 45.735 159.595 ;
        RECT 45.905 158.990 46.615 159.765 ;
        RECT 46.785 158.820 47.115 159.595 ;
        RECT 45.965 158.605 47.115 158.820 ;
        RECT 36.945 157.215 37.195 157.675 ;
        RECT 37.365 157.385 37.925 157.675 ;
        RECT 38.095 157.215 43.440 157.760 ;
        RECT 43.615 157.215 45.285 157.985 ;
        RECT 45.455 157.385 45.795 158.160 ;
        RECT 45.965 158.035 46.250 158.605 ;
        RECT 46.435 158.205 46.905 158.435 ;
        RECT 47.310 158.405 47.525 159.520 ;
        RECT 47.705 159.045 48.035 159.765 ;
        RECT 47.815 158.405 48.045 158.745 ;
        RECT 48.215 158.675 49.885 159.765 ;
        RECT 50.145 159.145 50.315 159.575 ;
        RECT 50.485 159.315 50.815 159.765 ;
        RECT 50.145 158.915 50.825 159.145 ;
        RECT 47.075 158.225 47.525 158.405 ;
        RECT 47.075 158.205 47.405 158.225 ;
        RECT 47.715 158.205 48.045 158.405 ;
        RECT 45.965 157.845 46.675 158.035 ;
        RECT 46.375 157.705 46.675 157.845 ;
        RECT 46.865 157.845 48.045 158.035 ;
        RECT 46.865 157.765 47.195 157.845 ;
        RECT 46.375 157.695 46.690 157.705 ;
        RECT 46.375 157.685 46.700 157.695 ;
        RECT 46.375 157.680 46.710 157.685 ;
        RECT 45.965 157.215 46.135 157.675 ;
        RECT 46.375 157.670 46.715 157.680 ;
        RECT 46.375 157.665 46.720 157.670 ;
        RECT 46.375 157.655 46.725 157.665 ;
        RECT 46.375 157.650 46.730 157.655 ;
        RECT 46.375 157.385 46.735 157.650 ;
        RECT 47.365 157.215 47.535 157.675 ;
        RECT 47.705 157.385 48.045 157.845 ;
        RECT 48.215 157.985 48.965 158.505 ;
        RECT 49.135 158.155 49.885 158.675 ;
        RECT 50.120 158.405 50.420 158.745 ;
        RECT 50.115 158.235 50.420 158.405 ;
        RECT 48.215 157.215 49.885 157.985 ;
        RECT 50.120 157.895 50.420 158.235 ;
        RECT 50.590 158.265 50.825 158.915 ;
        RECT 51.015 158.605 51.300 159.550 ;
        RECT 51.480 159.295 52.165 159.765 ;
        RECT 51.475 158.775 52.170 159.085 ;
        RECT 52.345 158.710 52.650 159.495 ;
        RECT 52.835 158.810 53.105 159.765 ;
        RECT 51.015 158.455 51.875 158.605 ;
        RECT 51.015 158.435 52.305 158.455 ;
        RECT 50.590 157.935 51.145 158.265 ;
        RECT 51.315 158.075 52.305 158.435 ;
        RECT 50.590 157.785 50.805 157.935 ;
        RECT 50.065 157.215 50.395 157.720 ;
        RECT 50.565 157.410 50.805 157.785 ;
        RECT 51.315 157.740 51.485 158.075 ;
        RECT 52.475 157.905 52.650 158.710 ;
        RECT 53.275 158.675 54.485 159.765 ;
        RECT 51.085 157.545 51.485 157.740 ;
        RECT 51.085 157.400 51.255 157.545 ;
        RECT 51.845 157.215 52.245 157.710 ;
        RECT 52.415 157.385 52.650 157.905 ;
        RECT 53.275 157.965 53.795 158.505 ;
        RECT 53.965 158.135 54.485 158.675 ;
        RECT 54.655 158.600 54.945 159.765 ;
        RECT 55.555 158.625 55.895 159.765 ;
        RECT 56.065 159.085 56.235 159.595 ;
        RECT 56.445 159.265 56.695 159.765 ;
        RECT 56.905 159.385 58.165 159.595 ;
        RECT 56.905 159.085 57.155 159.385 ;
        RECT 56.065 158.915 57.155 159.085 ;
        RECT 57.385 158.915 57.735 159.215 ;
        RECT 57.905 158.965 58.165 159.385 ;
        RECT 56.065 158.875 56.235 158.915 ;
        RECT 56.995 158.555 57.395 158.745 ;
        RECT 55.500 158.145 55.915 158.455 ;
        RECT 56.085 158.125 56.445 158.455 ;
        RECT 56.655 158.205 57.020 158.385 ;
        RECT 52.835 157.215 53.105 157.850 ;
        RECT 53.275 157.215 54.485 157.965 ;
        RECT 54.655 157.215 54.945 157.940 ;
        RECT 55.555 157.215 55.895 157.935 ;
        RECT 56.085 157.545 56.285 158.125 ;
        RECT 56.655 157.895 56.845 158.205 ;
        RECT 57.225 158.125 57.395 158.555 ;
        RECT 57.565 157.935 57.735 158.915 ;
        RECT 58.335 158.675 60.005 159.765 ;
        RECT 57.905 158.125 58.165 158.455 ;
        RECT 56.545 157.475 56.845 157.895 ;
        RECT 57.085 157.765 57.735 157.935 ;
        RECT 58.335 157.985 59.085 158.505 ;
        RECT 59.255 158.155 60.005 158.675 ;
        RECT 60.645 159.155 60.975 159.585 ;
        RECT 61.155 159.325 61.350 159.765 ;
        RECT 61.520 159.155 61.850 159.585 ;
        RECT 60.645 158.985 61.850 159.155 ;
        RECT 60.645 158.655 61.540 158.985 ;
        RECT 62.020 158.815 62.295 159.585 ;
        RECT 62.940 159.255 64.595 159.545 ;
        RECT 61.710 158.625 62.295 158.815 ;
        RECT 62.940 158.915 64.530 159.085 ;
        RECT 64.765 158.965 65.045 159.765 ;
        RECT 62.940 158.625 63.260 158.915 ;
        RECT 64.360 158.795 64.530 158.915 ;
        RECT 60.650 158.125 60.945 158.455 ;
        RECT 61.125 158.125 61.540 158.455 ;
        RECT 57.085 157.725 57.335 157.765 ;
        RECT 57.015 157.555 57.335 157.725 ;
        RECT 57.085 157.425 57.335 157.555 ;
        RECT 57.825 157.215 58.155 157.595 ;
        RECT 58.335 157.215 60.005 157.985 ;
        RECT 60.645 157.215 60.945 157.945 ;
        RECT 61.125 157.505 61.355 158.125 ;
        RECT 61.710 157.955 61.885 158.625 ;
        RECT 63.455 158.575 64.170 158.745 ;
        RECT 64.360 158.625 65.085 158.795 ;
        RECT 65.255 158.625 65.525 159.595 ;
        RECT 65.695 158.675 68.285 159.765 ;
        RECT 68.915 159.210 69.520 159.765 ;
        RECT 69.695 159.255 70.175 159.595 ;
        RECT 70.345 159.220 70.600 159.765 ;
        RECT 68.915 159.110 69.530 159.210 ;
        RECT 69.345 159.085 69.530 159.110 ;
        RECT 61.555 157.775 61.885 157.955 ;
        RECT 62.055 157.805 62.295 158.455 ;
        RECT 62.940 157.885 63.290 158.455 ;
        RECT 63.460 158.125 64.170 158.575 ;
        RECT 64.915 158.455 65.085 158.625 ;
        RECT 64.340 158.125 64.745 158.455 ;
        RECT 64.915 158.125 65.185 158.455 ;
        RECT 64.915 157.955 65.085 158.125 ;
        RECT 63.475 157.785 65.085 157.955 ;
        RECT 65.355 157.890 65.525 158.625 ;
        RECT 61.555 157.395 61.780 157.775 ;
        RECT 61.950 157.215 62.280 157.605 ;
        RECT 62.945 157.215 63.275 157.715 ;
        RECT 63.475 157.435 63.645 157.785 ;
        RECT 63.845 157.215 64.175 157.615 ;
        RECT 64.345 157.435 64.515 157.785 ;
        RECT 64.685 157.215 65.065 157.615 ;
        RECT 65.255 157.545 65.525 157.890 ;
        RECT 65.695 157.985 66.905 158.505 ;
        RECT 67.075 158.155 68.285 158.675 ;
        RECT 68.915 158.490 69.175 158.940 ;
        RECT 69.345 158.840 69.675 159.085 ;
        RECT 69.845 158.765 70.600 159.015 ;
        RECT 70.770 158.895 71.045 159.595 ;
        RECT 69.830 158.730 70.600 158.765 ;
        RECT 69.815 158.720 70.600 158.730 ;
        RECT 69.810 158.705 70.705 158.720 ;
        RECT 69.790 158.690 70.705 158.705 ;
        RECT 69.770 158.680 70.705 158.690 ;
        RECT 69.745 158.670 70.705 158.680 ;
        RECT 69.675 158.640 70.705 158.670 ;
        RECT 69.655 158.610 70.705 158.640 ;
        RECT 69.635 158.580 70.705 158.610 ;
        RECT 69.605 158.555 70.705 158.580 ;
        RECT 69.570 158.520 70.705 158.555 ;
        RECT 69.540 158.515 70.705 158.520 ;
        RECT 69.540 158.510 69.930 158.515 ;
        RECT 69.540 158.500 69.905 158.510 ;
        RECT 69.540 158.495 69.890 158.500 ;
        RECT 69.540 158.490 69.875 158.495 ;
        RECT 68.915 158.485 69.875 158.490 ;
        RECT 68.915 158.475 69.865 158.485 ;
        RECT 68.915 158.470 69.855 158.475 ;
        RECT 68.915 158.460 69.845 158.470 ;
        RECT 68.915 158.450 69.840 158.460 ;
        RECT 68.915 158.445 69.835 158.450 ;
        RECT 68.915 158.430 69.825 158.445 ;
        RECT 68.915 158.415 69.820 158.430 ;
        RECT 68.915 158.390 69.810 158.415 ;
        RECT 68.915 158.320 69.805 158.390 ;
        RECT 65.695 157.215 68.285 157.985 ;
        RECT 68.915 157.765 69.465 158.150 ;
        RECT 69.635 157.595 69.805 158.320 ;
        RECT 68.915 157.425 69.805 157.595 ;
        RECT 69.975 157.920 70.305 158.345 ;
        RECT 70.475 158.120 70.705 158.515 ;
        RECT 69.975 157.435 70.195 157.920 ;
        RECT 70.875 157.865 71.045 158.895 ;
        RECT 71.225 158.625 71.555 159.765 ;
        RECT 72.085 158.795 72.415 159.580 ;
        RECT 71.735 158.625 72.415 158.795 ;
        RECT 72.595 158.675 76.105 159.765 ;
        RECT 71.215 158.205 71.565 158.455 ;
        RECT 71.735 158.025 71.905 158.625 ;
        RECT 72.075 158.205 72.425 158.455 ;
        RECT 70.365 157.215 70.615 157.755 ;
        RECT 70.785 157.385 71.045 157.865 ;
        RECT 71.225 157.215 71.495 158.025 ;
        RECT 71.665 157.385 71.995 158.025 ;
        RECT 72.165 157.215 72.405 158.025 ;
        RECT 72.595 157.985 74.245 158.505 ;
        RECT 74.415 158.155 76.105 158.675 ;
        RECT 77.275 158.835 77.455 159.595 ;
        RECT 77.635 159.005 77.965 159.765 ;
        RECT 77.275 158.665 77.950 158.835 ;
        RECT 78.135 158.690 78.405 159.595 ;
        RECT 78.580 159.340 78.915 159.765 ;
        RECT 79.085 159.160 79.270 159.565 ;
        RECT 77.780 158.520 77.950 158.665 ;
        RECT 77.215 158.115 77.555 158.485 ;
        RECT 77.780 158.190 78.055 158.520 ;
        RECT 72.595 157.215 76.105 157.985 ;
        RECT 77.780 157.935 77.950 158.190 ;
        RECT 77.285 157.765 77.950 157.935 ;
        RECT 78.225 157.890 78.405 158.690 ;
        RECT 77.285 157.385 77.455 157.765 ;
        RECT 77.635 157.215 77.965 157.595 ;
        RECT 78.145 157.385 78.405 157.890 ;
        RECT 78.605 158.985 79.270 159.160 ;
        RECT 79.475 158.985 79.805 159.765 ;
        RECT 78.605 157.955 78.945 158.985 ;
        RECT 79.975 158.795 80.245 159.565 ;
        RECT 79.115 158.625 80.245 158.795 ;
        RECT 79.115 158.125 79.365 158.625 ;
        RECT 78.605 157.785 79.290 157.955 ;
        RECT 79.545 157.875 79.905 158.455 ;
        RECT 78.580 157.215 78.915 157.615 ;
        RECT 79.085 157.385 79.290 157.785 ;
        RECT 80.075 157.715 80.245 158.625 ;
        RECT 80.415 158.600 80.705 159.765 ;
        RECT 81.425 159.185 81.595 159.595 ;
        RECT 81.765 159.385 82.095 159.765 ;
        RECT 82.740 159.385 83.410 159.765 ;
        RECT 83.645 159.215 83.815 159.595 ;
        RECT 83.985 159.385 84.325 159.765 ;
        RECT 84.495 159.215 84.665 159.595 ;
        RECT 85.005 159.385 85.335 159.765 ;
        RECT 85.505 159.215 85.765 159.595 ;
        RECT 81.425 159.015 83.175 159.185 ;
        RECT 81.400 158.405 81.580 158.765 ;
        RECT 81.395 158.235 81.580 158.405 ;
        RECT 81.400 158.125 81.580 158.235 ;
        RECT 79.500 157.215 79.775 157.695 ;
        RECT 79.985 157.385 80.245 157.715 ;
        RECT 80.415 157.215 80.705 157.940 ;
        RECT 81.750 157.935 81.920 159.015 ;
        RECT 82.240 158.675 82.570 158.845 ;
        RECT 81.425 157.765 81.920 157.935 ;
        RECT 81.425 157.385 81.595 157.765 ;
        RECT 81.765 157.215 82.095 157.595 ;
        RECT 82.265 157.385 82.490 158.675 ;
        RECT 83.005 158.455 83.175 159.015 ;
        RECT 83.485 159.045 84.665 159.215 ;
        RECT 84.835 159.045 85.765 159.215 ;
        RECT 82.665 157.935 82.835 158.455 ;
        RECT 83.005 158.125 83.315 158.455 ;
        RECT 83.485 157.935 83.655 159.045 ;
        RECT 84.835 158.875 85.005 159.045 ;
        RECT 83.825 158.705 85.005 158.875 ;
        RECT 83.825 158.530 83.995 158.705 ;
        RECT 84.155 158.235 84.425 158.405 ;
        RECT 82.665 157.765 83.655 157.935 ;
        RECT 82.660 157.215 82.990 157.595 ;
        RECT 83.260 157.385 83.430 157.765 ;
        RECT 84.160 157.550 84.425 158.235 ;
        RECT 84.600 157.555 84.905 158.535 ;
        RECT 85.075 157.895 85.425 158.435 ;
        RECT 85.595 157.715 85.765 159.045 ;
        RECT 85.935 158.675 87.145 159.765 ;
        RECT 85.935 158.135 86.455 158.675 ;
        RECT 86.625 157.965 87.145 158.505 ;
        RECT 85.085 157.215 85.335 157.715 ;
        RECT 85.505 157.385 85.765 157.715 ;
        RECT 85.935 157.215 87.145 157.965 ;
        RECT 15.930 157.045 87.230 157.215 ;
        RECT 16.015 156.295 17.225 157.045 ;
        RECT 17.395 156.475 17.830 156.875 ;
        RECT 18.000 156.645 18.385 157.045 ;
        RECT 17.395 156.305 18.385 156.475 ;
        RECT 18.555 156.305 18.980 156.875 ;
        RECT 19.170 156.475 19.425 156.875 ;
        RECT 19.595 156.645 19.980 157.045 ;
        RECT 19.170 156.305 19.980 156.475 ;
        RECT 20.150 156.305 20.395 156.875 ;
        RECT 20.585 156.475 20.840 156.875 ;
        RECT 21.010 156.645 21.395 157.045 ;
        RECT 20.585 156.305 21.395 156.475 ;
        RECT 21.565 156.305 21.825 156.875 ;
        RECT 23.000 156.475 23.175 156.875 ;
        RECT 23.345 156.665 23.675 157.045 ;
        RECT 23.920 156.545 24.150 156.875 ;
        RECT 23.000 156.305 23.630 156.475 ;
        RECT 16.015 155.755 16.535 156.295 ;
        RECT 18.050 156.135 18.385 156.305 ;
        RECT 18.630 156.135 18.980 156.305 ;
        RECT 19.630 156.135 19.980 156.305 ;
        RECT 20.225 156.135 20.395 156.305 ;
        RECT 21.045 156.135 21.395 156.305 ;
        RECT 16.705 155.585 17.225 156.125 ;
        RECT 16.015 154.495 17.225 155.585 ;
        RECT 17.395 155.430 17.880 156.135 ;
        RECT 18.050 155.805 18.460 156.135 ;
        RECT 18.050 155.260 18.385 155.805 ;
        RECT 18.630 155.635 19.460 156.135 ;
        RECT 17.395 155.090 18.385 155.260 ;
        RECT 18.555 155.455 19.460 155.635 ;
        RECT 19.630 155.805 20.055 156.135 ;
        RECT 17.395 154.665 17.830 155.090 ;
        RECT 18.000 154.495 18.385 154.920 ;
        RECT 18.555 154.665 18.980 155.455 ;
        RECT 19.630 155.285 19.980 155.805 ;
        RECT 20.225 155.635 20.875 156.135 ;
        RECT 19.150 155.090 19.980 155.285 ;
        RECT 20.150 155.455 20.875 155.635 ;
        RECT 21.045 155.805 21.470 156.135 ;
        RECT 19.150 154.665 19.425 155.090 ;
        RECT 19.595 154.495 19.980 154.920 ;
        RECT 20.150 154.665 20.395 155.455 ;
        RECT 21.045 155.285 21.395 155.805 ;
        RECT 21.640 155.635 21.825 156.305 ;
        RECT 23.460 156.135 23.630 156.305 ;
        RECT 20.585 155.090 21.395 155.285 ;
        RECT 20.585 154.665 20.840 155.090 ;
        RECT 21.010 154.495 21.395 154.920 ;
        RECT 21.565 154.665 21.825 155.635 ;
        RECT 22.915 155.455 23.280 156.135 ;
        RECT 23.460 155.805 23.810 156.135 ;
        RECT 23.460 155.285 23.630 155.805 ;
        RECT 23.000 155.115 23.630 155.285 ;
        RECT 23.980 155.255 24.150 156.545 ;
        RECT 24.350 155.435 24.630 156.710 ;
        RECT 24.855 155.685 25.125 156.710 ;
        RECT 25.585 156.665 25.915 157.045 ;
        RECT 26.085 156.790 26.420 156.835 ;
        RECT 24.815 155.515 25.125 155.685 ;
        RECT 24.855 155.435 25.125 155.515 ;
        RECT 25.315 155.435 25.655 156.465 ;
        RECT 26.085 156.325 26.425 156.790 ;
        RECT 25.825 155.805 26.085 156.135 ;
        RECT 25.825 155.255 25.995 155.805 ;
        RECT 26.255 155.635 26.425 156.325 ;
        RECT 23.000 154.665 23.175 155.115 ;
        RECT 23.980 155.085 25.995 155.255 ;
        RECT 23.345 154.495 23.675 154.935 ;
        RECT 23.980 154.665 24.150 155.085 ;
        RECT 24.385 154.495 25.055 154.905 ;
        RECT 25.270 154.665 25.440 155.085 ;
        RECT 25.640 154.495 25.970 154.905 ;
        RECT 26.165 154.665 26.425 155.635 ;
        RECT 26.595 156.545 26.855 156.875 ;
        RECT 27.165 156.665 27.495 157.045 ;
        RECT 27.675 156.705 29.155 156.875 ;
        RECT 26.595 155.845 26.765 156.545 ;
        RECT 27.675 156.375 28.075 156.705 ;
        RECT 27.115 156.185 27.325 156.365 ;
        RECT 27.115 156.015 27.735 156.185 ;
        RECT 27.905 155.895 28.075 156.375 ;
        RECT 28.265 156.205 28.815 156.535 ;
        RECT 26.595 155.675 27.725 155.845 ;
        RECT 27.905 155.725 28.475 155.895 ;
        RECT 26.595 154.995 26.765 155.675 ;
        RECT 27.555 155.555 27.725 155.675 ;
        RECT 26.935 155.175 27.285 155.505 ;
        RECT 27.555 155.385 28.135 155.555 ;
        RECT 28.305 155.215 28.475 155.725 ;
        RECT 27.735 155.045 28.475 155.215 ;
        RECT 28.645 155.215 28.815 156.205 ;
        RECT 28.985 155.805 29.155 156.705 ;
        RECT 29.405 156.135 29.590 156.715 ;
        RECT 29.860 156.135 30.055 156.710 ;
        RECT 30.265 156.665 30.595 157.045 ;
        RECT 29.405 155.805 29.635 156.135 ;
        RECT 29.860 155.805 30.115 156.135 ;
        RECT 29.405 155.495 29.590 155.805 ;
        RECT 29.860 155.495 30.055 155.805 ;
        RECT 30.425 155.215 30.595 156.135 ;
        RECT 28.645 155.045 30.595 155.215 ;
        RECT 26.595 154.665 26.855 154.995 ;
        RECT 27.165 154.495 27.495 154.875 ;
        RECT 27.735 154.665 27.925 155.045 ;
        RECT 28.175 154.495 28.505 154.875 ;
        RECT 28.715 154.665 28.885 155.045 ;
        RECT 29.080 154.495 29.410 154.875 ;
        RECT 29.670 154.665 29.840 155.045 ;
        RECT 30.265 154.495 30.595 154.875 ;
        RECT 30.765 154.665 31.025 156.875 ;
        RECT 31.195 156.275 33.785 157.045 ;
        RECT 34.110 156.395 34.440 156.860 ;
        RECT 34.610 156.575 34.780 157.045 ;
        RECT 34.950 156.395 35.280 156.875 ;
        RECT 31.195 155.755 32.405 156.275 ;
        RECT 34.110 156.225 35.280 156.395 ;
        RECT 32.575 155.585 33.785 156.105 ;
        RECT 33.955 155.845 34.600 156.055 ;
        RECT 34.770 155.845 35.340 156.055 ;
        RECT 35.510 155.675 35.680 156.875 ;
        RECT 36.220 156.475 36.390 156.680 ;
        RECT 31.195 154.495 33.785 155.585 ;
        RECT 34.170 154.495 34.500 155.595 ;
        RECT 34.975 155.265 35.680 155.675 ;
        RECT 35.850 156.305 36.390 156.475 ;
        RECT 36.670 156.305 36.840 157.045 ;
        RECT 37.105 156.305 37.465 156.680 ;
        RECT 35.850 155.605 36.020 156.305 ;
        RECT 36.190 155.805 36.520 156.135 ;
        RECT 36.690 155.805 37.040 156.135 ;
        RECT 35.850 155.435 36.475 155.605 ;
        RECT 36.690 155.265 36.955 155.805 ;
        RECT 37.210 155.650 37.465 156.305 ;
        RECT 37.635 156.275 41.145 157.045 ;
        RECT 41.775 156.320 42.065 157.045 ;
        RECT 37.635 155.755 39.285 156.275 ;
        RECT 34.975 155.095 36.955 155.265 ;
        RECT 34.975 154.665 35.300 155.095 ;
        RECT 35.470 154.495 35.800 154.915 ;
        RECT 36.545 154.495 36.955 154.925 ;
        RECT 37.125 154.665 37.465 155.650 ;
        RECT 39.455 155.585 41.145 156.105 ;
        RECT 37.635 154.495 41.145 155.585 ;
        RECT 41.775 154.495 42.065 155.660 ;
        RECT 42.240 155.445 42.575 156.865 ;
        RECT 42.755 156.675 43.500 157.045 ;
        RECT 44.065 156.505 44.320 156.865 ;
        RECT 44.500 156.675 44.830 157.045 ;
        RECT 45.010 156.505 45.235 156.865 ;
        RECT 42.750 156.315 45.235 156.505 ;
        RECT 42.750 155.625 42.975 156.315 ;
        RECT 43.175 155.805 43.455 156.135 ;
        RECT 43.635 155.805 44.210 156.135 ;
        RECT 44.390 155.805 44.825 156.135 ;
        RECT 45.005 155.805 45.275 156.135 ;
        RECT 42.750 155.445 45.245 155.625 ;
        RECT 42.240 154.675 42.505 155.445 ;
        RECT 42.675 154.495 43.005 155.215 ;
        RECT 43.195 155.035 44.385 155.265 ;
        RECT 43.195 154.675 43.455 155.035 ;
        RECT 43.625 154.495 43.955 154.865 ;
        RECT 44.125 154.675 44.385 155.035 ;
        RECT 44.955 154.675 45.245 155.445 ;
        RECT 45.465 154.675 45.725 156.865 ;
        RECT 45.985 156.675 46.655 157.045 ;
        RECT 46.835 156.495 47.145 156.865 ;
        RECT 45.915 156.295 47.145 156.495 ;
        RECT 45.915 155.625 46.205 156.295 ;
        RECT 47.325 156.115 47.555 156.755 ;
        RECT 47.735 156.315 48.025 157.045 ;
        RECT 48.215 156.275 49.885 157.045 ;
        RECT 46.385 155.805 46.850 156.115 ;
        RECT 47.030 155.805 47.555 156.115 ;
        RECT 47.735 155.805 48.035 156.135 ;
        RECT 48.215 155.755 48.965 156.275 ;
        RECT 50.065 156.235 50.335 157.045 ;
        RECT 50.505 156.235 50.835 156.875 ;
        RECT 51.005 156.235 51.245 157.045 ;
        RECT 51.435 156.500 56.780 157.045 ;
        RECT 45.915 155.405 46.685 155.625 ;
        RECT 45.895 154.495 46.235 155.225 ;
        RECT 46.415 154.675 46.685 155.405 ;
        RECT 46.865 155.385 48.025 155.625 ;
        RECT 49.135 155.585 49.885 156.105 ;
        RECT 50.055 155.805 50.405 156.055 ;
        RECT 50.575 155.635 50.745 156.235 ;
        RECT 50.915 155.805 51.265 156.055 ;
        RECT 53.020 155.670 53.360 156.500 ;
        RECT 56.955 156.275 60.465 157.045 ;
        RECT 60.635 156.295 61.845 157.045 ;
        RECT 46.865 154.675 47.095 155.385 ;
        RECT 47.265 154.495 47.595 155.205 ;
        RECT 47.765 154.675 48.025 155.385 ;
        RECT 48.215 154.495 49.885 155.585 ;
        RECT 50.065 154.495 50.395 155.635 ;
        RECT 50.575 155.465 51.255 155.635 ;
        RECT 50.925 154.680 51.255 155.465 ;
        RECT 54.840 154.930 55.190 156.180 ;
        RECT 56.955 155.755 58.605 156.275 ;
        RECT 58.775 155.585 60.465 156.105 ;
        RECT 60.635 155.755 61.155 156.295 ;
        RECT 62.075 156.225 62.285 157.045 ;
        RECT 62.455 156.245 62.785 156.875 ;
        RECT 61.325 155.585 61.845 156.125 ;
        RECT 62.455 155.645 62.705 156.245 ;
        RECT 62.955 156.225 63.185 157.045 ;
        RECT 63.395 156.275 66.905 157.045 ;
        RECT 67.535 156.320 67.825 157.045 ;
        RECT 68.015 156.315 68.305 157.045 ;
        RECT 62.875 155.805 63.205 156.055 ;
        RECT 63.395 155.755 65.045 156.275 ;
        RECT 51.435 154.495 56.780 154.930 ;
        RECT 56.955 154.495 60.465 155.585 ;
        RECT 60.635 154.495 61.845 155.585 ;
        RECT 62.075 154.495 62.285 155.635 ;
        RECT 62.455 154.665 62.785 155.645 ;
        RECT 62.955 154.495 63.185 155.635 ;
        RECT 65.215 155.585 66.905 156.105 ;
        RECT 68.005 155.805 68.305 156.135 ;
        RECT 68.485 156.115 68.715 156.755 ;
        RECT 68.895 156.495 69.205 156.865 ;
        RECT 69.385 156.675 70.055 157.045 ;
        RECT 68.895 156.295 70.125 156.495 ;
        RECT 68.485 155.805 69.010 156.115 ;
        RECT 69.190 155.805 69.655 156.115 ;
        RECT 63.395 154.495 66.905 155.585 ;
        RECT 67.535 154.495 67.825 155.660 ;
        RECT 69.835 155.625 70.125 156.295 ;
        RECT 68.015 155.385 69.175 155.625 ;
        RECT 68.015 154.675 68.275 155.385 ;
        RECT 68.445 154.495 68.775 155.205 ;
        RECT 68.945 154.675 69.175 155.385 ;
        RECT 69.355 155.405 70.125 155.625 ;
        RECT 69.355 154.675 69.625 155.405 ;
        RECT 69.805 154.495 70.145 155.225 ;
        RECT 70.315 154.675 70.575 156.865 ;
        RECT 70.755 156.585 71.315 156.875 ;
        RECT 71.485 156.585 71.735 157.045 ;
        RECT 70.755 155.215 71.005 156.585 ;
        RECT 72.355 156.415 72.685 156.775 ;
        RECT 73.055 156.500 78.400 157.045 ;
        RECT 71.295 156.225 72.685 156.415 ;
        RECT 71.295 156.135 71.465 156.225 ;
        RECT 71.175 155.805 71.465 156.135 ;
        RECT 71.635 155.805 71.975 156.055 ;
        RECT 72.195 155.805 72.870 156.055 ;
        RECT 71.295 155.555 71.465 155.805 ;
        RECT 71.295 155.385 72.235 155.555 ;
        RECT 72.605 155.445 72.870 155.805 ;
        RECT 74.640 155.670 74.980 156.500 ;
        RECT 79.495 156.370 79.755 156.875 ;
        RECT 79.935 156.665 80.265 157.045 ;
        RECT 80.445 156.495 80.615 156.875 ;
        RECT 70.755 154.665 71.215 155.215 ;
        RECT 71.405 154.495 71.735 155.215 ;
        RECT 71.935 154.835 72.235 155.385 ;
        RECT 72.405 154.495 72.685 155.165 ;
        RECT 76.460 154.930 76.810 156.180 ;
        RECT 79.495 155.570 79.675 156.370 ;
        RECT 79.950 156.325 80.615 156.495 ;
        RECT 80.965 156.495 81.135 156.875 ;
        RECT 81.315 156.665 81.645 157.045 ;
        RECT 80.965 156.325 81.630 156.495 ;
        RECT 81.825 156.370 82.085 156.875 ;
        RECT 79.950 156.070 80.120 156.325 ;
        RECT 79.845 155.740 80.120 156.070 ;
        RECT 80.345 155.775 80.685 156.145 ;
        RECT 80.895 155.775 81.235 156.145 ;
        RECT 81.460 156.070 81.630 156.325 ;
        RECT 79.950 155.595 80.120 155.740 ;
        RECT 81.460 155.740 81.735 156.070 ;
        RECT 81.460 155.595 81.630 155.740 ;
        RECT 73.055 154.495 78.400 154.930 ;
        RECT 79.495 154.665 79.765 155.570 ;
        RECT 79.950 155.425 80.625 155.595 ;
        RECT 79.935 154.495 80.265 155.255 ;
        RECT 80.445 154.665 80.625 155.425 ;
        RECT 80.955 155.425 81.630 155.595 ;
        RECT 81.905 155.570 82.085 156.370 ;
        RECT 82.260 156.205 82.520 157.045 ;
        RECT 82.695 156.300 82.950 156.875 ;
        RECT 83.120 156.665 83.450 157.045 ;
        RECT 83.665 156.495 83.835 156.875 ;
        RECT 83.120 156.325 83.835 156.495 ;
        RECT 84.185 156.495 84.355 156.875 ;
        RECT 84.570 156.665 84.900 157.045 ;
        RECT 84.185 156.325 84.900 156.495 ;
        RECT 80.955 154.665 81.135 155.425 ;
        RECT 81.315 154.495 81.645 155.255 ;
        RECT 81.815 154.665 82.085 155.570 ;
        RECT 82.260 154.495 82.520 155.645 ;
        RECT 82.695 155.570 82.865 156.300 ;
        RECT 83.120 156.135 83.290 156.325 ;
        RECT 83.035 155.805 83.290 156.135 ;
        RECT 83.120 155.595 83.290 155.805 ;
        RECT 83.570 155.775 83.925 156.145 ;
        RECT 84.095 155.775 84.450 156.145 ;
        RECT 84.730 156.135 84.900 156.325 ;
        RECT 85.070 156.300 85.325 156.875 ;
        RECT 84.730 155.805 84.985 156.135 ;
        RECT 84.730 155.595 84.900 155.805 ;
        RECT 82.695 154.665 82.950 155.570 ;
        RECT 83.120 155.425 83.835 155.595 ;
        RECT 83.120 154.495 83.450 155.255 ;
        RECT 83.665 154.665 83.835 155.425 ;
        RECT 84.185 155.425 84.900 155.595 ;
        RECT 85.155 155.570 85.325 156.300 ;
        RECT 85.500 156.205 85.760 157.045 ;
        RECT 85.935 156.295 87.145 157.045 ;
        RECT 84.185 154.665 84.355 155.425 ;
        RECT 84.570 154.495 84.900 155.255 ;
        RECT 85.070 154.665 85.325 155.570 ;
        RECT 85.500 154.495 85.760 155.645 ;
        RECT 85.935 155.585 86.455 156.125 ;
        RECT 86.625 155.755 87.145 156.295 ;
        RECT 85.935 154.495 87.145 155.585 ;
        RECT 15.930 154.325 87.230 154.495 ;
        RECT 16.015 153.235 17.225 154.325 ;
        RECT 16.015 152.525 16.535 153.065 ;
        RECT 16.705 152.695 17.225 153.235 ;
        RECT 17.395 153.185 17.685 154.325 ;
        RECT 17.855 153.605 18.305 154.155 ;
        RECT 18.495 153.605 18.825 154.325 ;
        RECT 16.015 151.775 17.225 152.525 ;
        RECT 17.395 151.775 17.685 152.575 ;
        RECT 17.855 152.235 18.105 153.605 ;
        RECT 19.035 153.435 19.335 153.985 ;
        RECT 19.505 153.655 19.785 154.325 ;
        RECT 20.245 153.705 20.415 154.135 ;
        RECT 20.585 153.875 20.915 154.325 ;
        RECT 20.245 153.475 20.920 153.705 ;
        RECT 18.395 153.265 19.335 153.435 ;
        RECT 18.395 153.015 18.565 153.265 ;
        RECT 19.670 153.015 19.985 153.455 ;
        RECT 18.275 152.685 18.565 153.015 ;
        RECT 18.735 152.765 19.065 153.015 ;
        RECT 19.295 152.765 19.985 153.015 ;
        RECT 18.395 152.595 18.565 152.685 ;
        RECT 18.395 152.405 19.785 152.595 ;
        RECT 20.215 152.455 20.515 153.305 ;
        RECT 20.685 152.825 20.920 153.475 ;
        RECT 21.090 153.165 21.375 154.110 ;
        RECT 21.555 153.855 22.240 154.325 ;
        RECT 21.550 153.335 22.245 153.645 ;
        RECT 22.420 153.270 22.725 154.055 ;
        RECT 21.090 153.015 21.950 153.165 ;
        RECT 21.090 152.995 22.375 153.015 ;
        RECT 20.685 152.495 21.220 152.825 ;
        RECT 21.390 152.635 22.375 152.995 ;
        RECT 17.855 151.945 18.405 152.235 ;
        RECT 18.575 151.775 18.825 152.235 ;
        RECT 19.455 152.045 19.785 152.405 ;
        RECT 20.685 152.345 20.905 152.495 ;
        RECT 20.160 151.775 20.495 152.280 ;
        RECT 20.665 151.970 20.905 152.345 ;
        RECT 21.390 152.300 21.560 152.635 ;
        RECT 22.550 152.465 22.725 153.270 ;
        RECT 22.915 153.235 24.585 154.325 ;
        RECT 25.215 153.815 25.475 154.325 ;
        RECT 21.185 152.105 21.560 152.300 ;
        RECT 21.185 151.960 21.355 152.105 ;
        RECT 21.920 151.775 22.315 152.270 ;
        RECT 22.485 151.945 22.725 152.465 ;
        RECT 22.915 152.545 23.665 153.065 ;
        RECT 23.835 152.715 24.585 153.235 ;
        RECT 25.215 152.765 25.555 153.645 ;
        RECT 25.725 152.935 25.895 154.155 ;
        RECT 26.135 153.820 26.750 154.325 ;
        RECT 26.135 153.285 26.385 153.650 ;
        RECT 26.555 153.645 26.750 153.820 ;
        RECT 26.920 153.815 27.395 154.155 ;
        RECT 27.565 153.780 27.780 154.325 ;
        RECT 26.555 153.455 26.885 153.645 ;
        RECT 27.105 153.285 27.820 153.580 ;
        RECT 27.990 153.455 28.265 154.155 ;
        RECT 26.135 153.115 27.925 153.285 ;
        RECT 25.725 152.685 26.520 152.935 ;
        RECT 25.725 152.595 25.975 152.685 ;
        RECT 22.915 151.775 24.585 152.545 ;
        RECT 25.215 151.775 25.475 152.595 ;
        RECT 25.645 152.175 25.975 152.595 ;
        RECT 26.690 152.260 26.945 153.115 ;
        RECT 26.155 151.995 26.945 152.260 ;
        RECT 27.115 152.415 27.525 152.935 ;
        RECT 27.695 152.685 27.925 153.115 ;
        RECT 28.095 152.425 28.265 153.455 ;
        RECT 28.895 153.160 29.185 154.325 ;
        RECT 29.355 153.815 29.615 154.325 ;
        RECT 29.355 152.765 29.695 153.645 ;
        RECT 29.865 152.935 30.035 154.155 ;
        RECT 30.275 153.820 30.890 154.325 ;
        RECT 30.275 153.285 30.525 153.650 ;
        RECT 30.695 153.645 30.890 153.820 ;
        RECT 31.060 153.815 31.535 154.155 ;
        RECT 31.705 153.780 31.920 154.325 ;
        RECT 30.695 153.455 31.025 153.645 ;
        RECT 31.245 153.285 31.960 153.580 ;
        RECT 32.130 153.455 32.405 154.155 ;
        RECT 30.275 153.115 32.065 153.285 ;
        RECT 29.865 152.685 30.660 152.935 ;
        RECT 29.865 152.595 30.115 152.685 ;
        RECT 27.115 151.995 27.315 152.415 ;
        RECT 27.505 151.775 27.835 152.235 ;
        RECT 28.005 151.945 28.265 152.425 ;
        RECT 28.895 151.775 29.185 152.500 ;
        RECT 29.355 151.775 29.615 152.595 ;
        RECT 29.785 152.175 30.115 152.595 ;
        RECT 30.830 152.260 31.085 153.115 ;
        RECT 30.295 151.995 31.085 152.260 ;
        RECT 31.255 152.415 31.665 152.935 ;
        RECT 31.835 152.685 32.065 153.115 ;
        RECT 32.235 152.425 32.405 153.455 ;
        RECT 33.560 153.355 33.830 154.150 ;
        RECT 34.010 153.525 34.225 154.325 ;
        RECT 34.405 153.355 34.690 154.150 ;
        RECT 33.560 153.185 34.690 153.355 ;
        RECT 33.540 152.715 34.040 152.980 ;
        RECT 34.260 152.685 34.645 153.015 ;
        RECT 34.870 152.685 35.150 154.155 ;
        RECT 35.330 152.740 35.660 154.155 ;
        RECT 35.830 152.980 36.035 154.155 ;
        RECT 36.205 153.335 36.415 154.150 ;
        RECT 36.655 153.505 36.985 154.325 ;
        RECT 36.205 153.155 36.855 153.335 ;
        RECT 37.160 153.310 37.415 154.150 ;
        RECT 37.640 153.900 37.975 154.325 ;
        RECT 38.145 153.720 38.330 154.125 ;
        RECT 35.830 152.740 36.260 152.980 ;
        RECT 34.260 152.535 34.565 152.685 ;
        RECT 31.255 151.995 31.455 152.415 ;
        RECT 31.645 151.775 31.975 152.235 ;
        RECT 32.145 151.945 32.405 152.425 ;
        RECT 33.595 151.775 33.835 152.450 ;
        RECT 34.010 151.975 34.565 152.535 ;
        RECT 36.635 152.515 36.855 153.155 ;
        RECT 34.745 152.345 36.855 152.515 ;
        RECT 34.745 151.950 34.950 152.345 ;
        RECT 35.635 152.340 36.855 152.345 ;
        RECT 35.120 151.775 35.465 152.175 ;
        RECT 35.635 151.950 35.965 152.340 ;
        RECT 36.240 151.775 36.915 152.160 ;
        RECT 37.085 151.945 37.415 153.310 ;
        RECT 37.665 153.545 38.330 153.720 ;
        RECT 38.535 153.545 38.865 154.325 ;
        RECT 37.665 152.515 38.005 153.545 ;
        RECT 39.035 153.355 39.305 154.125 ;
        RECT 38.175 153.185 39.305 153.355 ;
        RECT 39.485 153.185 39.815 154.325 ;
        RECT 40.345 153.355 40.675 154.140 ;
        RECT 41.515 153.655 41.795 154.325 ;
        RECT 41.965 153.435 42.265 153.985 ;
        RECT 42.465 153.605 42.795 154.325 ;
        RECT 42.985 153.605 43.445 154.155 ;
        RECT 39.995 153.185 40.675 153.355 ;
        RECT 38.175 152.685 38.425 153.185 ;
        RECT 37.665 152.345 38.350 152.515 ;
        RECT 38.605 152.435 38.965 153.015 ;
        RECT 37.640 151.775 37.975 152.175 ;
        RECT 38.145 151.945 38.350 152.345 ;
        RECT 39.135 152.275 39.305 153.185 ;
        RECT 39.475 152.765 39.825 153.015 ;
        RECT 39.995 152.585 40.165 153.185 ;
        RECT 41.330 153.015 41.595 153.375 ;
        RECT 41.965 153.265 42.905 153.435 ;
        RECT 42.735 153.015 42.905 153.265 ;
        RECT 40.335 152.765 40.685 153.015 ;
        RECT 41.330 152.765 42.005 153.015 ;
        RECT 42.225 152.765 42.565 153.015 ;
        RECT 42.735 152.685 43.025 153.015 ;
        RECT 42.735 152.595 42.905 152.685 ;
        RECT 38.560 151.775 38.835 152.255 ;
        RECT 39.045 151.945 39.305 152.275 ;
        RECT 39.485 151.775 39.755 152.585 ;
        RECT 39.925 151.945 40.255 152.585 ;
        RECT 40.425 151.775 40.665 152.585 ;
        RECT 41.515 152.405 42.905 152.595 ;
        RECT 41.515 152.045 41.845 152.405 ;
        RECT 43.195 152.235 43.445 153.605 ;
        RECT 44.110 153.525 44.360 154.325 ;
        RECT 44.530 153.695 44.860 154.155 ;
        RECT 45.030 153.865 45.245 154.325 ;
        RECT 44.530 153.525 45.700 153.695 ;
        RECT 43.620 153.355 43.900 153.515 ;
        RECT 43.620 153.185 44.955 153.355 ;
        RECT 44.785 153.015 44.955 153.185 ;
        RECT 43.620 152.765 43.970 153.005 ;
        RECT 44.140 152.765 44.615 153.005 ;
        RECT 44.785 152.765 45.160 153.015 ;
        RECT 44.785 152.595 44.955 152.765 ;
        RECT 42.465 151.775 42.715 152.235 ;
        RECT 42.885 151.945 43.445 152.235 ;
        RECT 43.620 152.425 44.955 152.595 ;
        RECT 43.620 152.215 43.890 152.425 ;
        RECT 45.330 152.235 45.700 153.525 ;
        RECT 45.915 153.235 47.585 154.325 ;
        RECT 44.110 151.775 44.440 152.235 ;
        RECT 44.950 151.945 45.700 152.235 ;
        RECT 45.915 152.545 46.665 153.065 ;
        RECT 46.835 152.715 47.585 153.235 ;
        RECT 48.215 153.475 48.555 154.115 ;
        RECT 48.725 153.865 48.970 154.325 ;
        RECT 49.145 153.695 49.395 154.155 ;
        RECT 49.585 153.945 50.255 154.325 ;
        RECT 50.455 153.695 50.705 154.155 ;
        RECT 49.145 153.525 50.705 153.695 ;
        RECT 45.915 151.775 47.585 152.545 ;
        RECT 48.215 152.360 48.385 153.475 ;
        RECT 51.465 153.355 51.635 154.155 ;
        RECT 48.695 153.185 51.635 153.355 ;
        RECT 51.985 153.395 52.155 154.155 ;
        RECT 52.370 153.565 52.700 154.325 ;
        RECT 51.985 153.225 52.700 153.395 ;
        RECT 52.870 153.250 53.125 154.155 ;
        RECT 48.695 153.015 48.865 153.185 ;
        RECT 48.555 152.685 48.865 153.015 ;
        RECT 49.035 152.685 49.370 153.015 ;
        RECT 48.695 152.515 48.865 152.685 ;
        RECT 48.215 151.945 48.525 152.360 ;
        RECT 48.695 152.345 49.390 152.515 ;
        RECT 49.640 152.440 49.835 153.015 ;
        RECT 50.095 152.685 50.440 153.015 ;
        RECT 50.750 152.685 51.225 153.015 ;
        RECT 51.480 152.685 51.665 153.015 ;
        RECT 50.095 152.455 50.285 152.685 ;
        RECT 51.895 152.675 52.250 153.045 ;
        RECT 52.530 153.015 52.700 153.225 ;
        RECT 52.530 152.685 52.785 153.015 ;
        RECT 48.720 151.775 49.050 152.155 ;
        RECT 49.220 152.115 49.390 152.345 ;
        RECT 50.455 152.345 51.635 152.515 ;
        RECT 52.530 152.495 52.700 152.685 ;
        RECT 52.955 152.520 53.125 153.250 ;
        RECT 53.300 153.175 53.560 154.325 ;
        RECT 54.655 153.160 54.945 154.325 ;
        RECT 50.455 152.115 50.625 152.345 ;
        RECT 49.220 151.945 50.625 152.115 ;
        RECT 50.895 151.775 51.225 152.175 ;
        RECT 51.465 151.945 51.635 152.345 ;
        RECT 51.985 152.325 52.700 152.495 ;
        RECT 51.985 151.945 52.155 152.325 ;
        RECT 52.370 151.775 52.700 152.155 ;
        RECT 52.870 151.945 53.125 152.520 ;
        RECT 53.300 151.775 53.560 152.615 ;
        RECT 54.655 151.775 54.945 152.500 ;
        RECT 55.115 152.055 55.395 154.155 ;
        RECT 55.585 153.565 56.370 154.325 ;
        RECT 56.765 153.495 57.150 154.155 ;
        RECT 56.765 153.395 57.175 153.495 ;
        RECT 55.565 153.185 57.175 153.395 ;
        RECT 57.475 153.305 57.675 154.095 ;
        RECT 55.565 152.585 55.840 153.185 ;
        RECT 57.345 153.135 57.675 153.305 ;
        RECT 57.845 153.145 58.165 154.325 ;
        RECT 58.335 153.725 58.595 154.145 ;
        RECT 58.765 153.895 59.095 154.325 ;
        RECT 59.785 153.895 60.530 154.065 ;
        RECT 58.335 153.555 60.190 153.725 ;
        RECT 57.345 153.015 57.525 153.135 ;
        RECT 56.010 152.765 56.365 153.015 ;
        RECT 56.560 152.965 57.025 153.015 ;
        RECT 56.555 152.795 57.025 152.965 ;
        RECT 56.560 152.765 57.025 152.795 ;
        RECT 57.195 152.765 57.525 153.015 ;
        RECT 57.700 152.765 58.165 152.965 ;
        RECT 55.565 152.405 56.815 152.585 ;
        RECT 56.450 152.335 56.815 152.405 ;
        RECT 56.985 152.385 58.165 152.555 ;
        RECT 55.625 151.775 55.795 152.235 ;
        RECT 56.985 152.165 57.315 152.385 ;
        RECT 56.065 151.985 57.315 152.165 ;
        RECT 57.485 151.775 57.655 152.215 ;
        RECT 57.825 151.970 58.165 152.385 ;
        RECT 58.335 152.515 58.510 153.555 ;
        RECT 58.680 152.685 59.030 153.385 ;
        RECT 59.245 153.215 59.850 153.385 ;
        RECT 59.200 152.685 59.490 153.015 ;
        RECT 59.660 152.935 59.850 153.215 ;
        RECT 60.020 153.275 60.190 153.555 ;
        RECT 60.360 153.645 60.530 153.895 ;
        RECT 60.755 153.815 61.395 154.145 ;
        RECT 60.360 153.475 61.395 153.645 ;
        RECT 61.565 153.525 61.845 154.325 ;
        RECT 61.225 153.355 61.395 153.475 ;
        RECT 60.020 153.105 60.670 153.275 ;
        RECT 61.225 153.185 61.885 153.355 ;
        RECT 62.055 153.185 62.330 154.155 ;
        RECT 59.660 152.765 60.105 152.935 ;
        RECT 59.660 152.515 59.850 152.765 ;
        RECT 60.500 152.685 60.670 153.105 ;
        RECT 61.715 153.015 61.885 153.185 ;
        RECT 60.890 152.685 61.545 153.015 ;
        RECT 61.715 152.685 61.990 153.015 ;
        RECT 61.715 152.515 61.885 152.685 ;
        RECT 58.335 152.140 58.655 152.515 ;
        RECT 58.910 151.775 59.080 152.515 ;
        RECT 59.330 152.345 59.850 152.515 ;
        RECT 60.275 152.345 61.885 152.515 ;
        RECT 62.160 152.450 62.330 153.185 ;
        RECT 62.500 153.130 62.670 154.325 ;
        RECT 62.935 153.185 63.195 154.325 ;
        RECT 63.365 153.175 63.695 154.155 ;
        RECT 63.865 153.185 64.145 154.325 ;
        RECT 64.315 153.235 65.525 154.325 ;
        RECT 62.955 152.765 63.290 153.015 ;
        RECT 59.330 152.140 59.500 152.345 ;
        RECT 59.745 151.775 60.100 152.175 ;
        RECT 60.275 151.995 60.445 152.345 ;
        RECT 60.645 151.775 60.975 152.175 ;
        RECT 61.145 151.995 61.315 152.345 ;
        RECT 61.485 151.775 61.865 152.175 ;
        RECT 62.055 152.105 62.330 152.450 ;
        RECT 62.500 151.775 62.670 152.715 ;
        RECT 63.460 152.575 63.630 153.175 ;
        RECT 63.800 152.745 64.135 153.015 ;
        RECT 62.935 151.945 63.630 152.575 ;
        RECT 63.835 151.775 64.145 152.575 ;
        RECT 64.315 152.525 64.835 153.065 ;
        RECT 65.005 152.695 65.525 153.235 ;
        RECT 65.715 153.435 65.975 154.145 ;
        RECT 66.145 153.615 66.475 154.325 ;
        RECT 66.645 153.435 66.875 154.145 ;
        RECT 65.715 153.195 66.875 153.435 ;
        RECT 67.055 153.415 67.325 154.145 ;
        RECT 67.505 153.595 67.845 154.325 ;
        RECT 67.055 153.195 67.825 153.415 ;
        RECT 65.705 152.685 66.005 153.015 ;
        RECT 66.185 152.705 66.710 153.015 ;
        RECT 66.890 152.705 67.355 153.015 ;
        RECT 64.315 151.775 65.525 152.525 ;
        RECT 65.715 151.775 66.005 152.505 ;
        RECT 66.185 152.065 66.415 152.705 ;
        RECT 67.535 152.525 67.825 153.195 ;
        RECT 66.595 152.325 67.825 152.525 ;
        RECT 66.595 151.955 66.905 152.325 ;
        RECT 67.085 151.775 67.755 152.145 ;
        RECT 68.015 151.955 68.275 154.145 ;
        RECT 68.465 153.715 68.795 154.145 ;
        RECT 68.975 153.885 69.170 154.325 ;
        RECT 69.340 153.715 69.670 154.145 ;
        RECT 68.465 153.545 69.670 153.715 ;
        RECT 68.465 153.215 69.360 153.545 ;
        RECT 69.840 153.375 70.115 154.145 ;
        RECT 70.295 153.890 75.640 154.325 ;
        RECT 69.530 153.185 70.115 153.375 ;
        RECT 68.470 152.685 68.765 153.015 ;
        RECT 68.945 152.685 69.360 153.015 ;
        RECT 68.465 151.775 68.765 152.505 ;
        RECT 68.945 152.065 69.175 152.685 ;
        RECT 69.530 152.515 69.705 153.185 ;
        RECT 69.375 152.335 69.705 152.515 ;
        RECT 69.875 152.365 70.115 153.015 ;
        RECT 69.375 151.955 69.600 152.335 ;
        RECT 71.880 152.320 72.220 153.150 ;
        RECT 73.700 152.640 74.050 153.890 ;
        RECT 75.815 153.235 79.325 154.325 ;
        RECT 75.815 152.545 77.465 153.065 ;
        RECT 77.635 152.715 79.325 153.235 ;
        RECT 80.415 153.160 80.705 154.325 ;
        RECT 80.875 153.235 82.545 154.325 ;
        RECT 80.875 152.545 81.625 153.065 ;
        RECT 81.795 152.715 82.545 153.235 ;
        RECT 82.795 153.395 82.975 154.155 ;
        RECT 83.155 153.565 83.485 154.325 ;
        RECT 82.795 153.225 83.470 153.395 ;
        RECT 83.655 153.250 83.925 154.155 ;
        RECT 83.300 153.080 83.470 153.225 ;
        RECT 82.735 152.675 83.075 153.045 ;
        RECT 83.300 152.750 83.575 153.080 ;
        RECT 69.770 151.775 70.100 152.165 ;
        RECT 70.295 151.775 75.640 152.320 ;
        RECT 75.815 151.775 79.325 152.545 ;
        RECT 80.415 151.775 80.705 152.500 ;
        RECT 80.875 151.775 82.545 152.545 ;
        RECT 83.300 152.495 83.470 152.750 ;
        RECT 82.805 152.325 83.470 152.495 ;
        RECT 83.745 152.450 83.925 153.250 ;
        RECT 82.805 151.945 82.975 152.325 ;
        RECT 83.155 151.775 83.485 152.155 ;
        RECT 83.665 151.945 83.925 152.450 ;
        RECT 84.095 153.355 84.365 154.125 ;
        RECT 84.535 153.545 84.865 154.325 ;
        RECT 85.070 153.720 85.255 154.125 ;
        RECT 85.425 153.900 85.760 154.325 ;
        RECT 85.070 153.545 85.735 153.720 ;
        RECT 84.095 153.185 85.225 153.355 ;
        RECT 84.095 152.275 84.265 153.185 ;
        RECT 84.435 152.435 84.795 153.015 ;
        RECT 84.975 152.685 85.225 153.185 ;
        RECT 85.395 152.515 85.735 153.545 ;
        RECT 85.935 153.235 87.145 154.325 ;
        RECT 85.935 152.695 86.455 153.235 ;
        RECT 86.625 152.525 87.145 153.065 ;
        RECT 85.050 152.345 85.735 152.515 ;
        RECT 84.095 151.945 84.355 152.275 ;
        RECT 84.565 151.775 84.840 152.255 ;
        RECT 85.050 151.945 85.255 152.345 ;
        RECT 85.425 151.775 85.760 152.175 ;
        RECT 85.935 151.775 87.145 152.525 ;
        RECT 15.930 151.605 87.230 151.775 ;
        RECT 16.015 150.855 17.225 151.605 ;
        RECT 16.015 150.315 16.535 150.855 ;
        RECT 17.400 150.765 17.660 151.605 ;
        RECT 17.835 150.860 18.090 151.435 ;
        RECT 18.260 151.225 18.590 151.605 ;
        RECT 18.805 151.055 18.975 151.435 ;
        RECT 18.260 150.885 18.975 151.055 ;
        RECT 16.705 150.145 17.225 150.685 ;
        RECT 16.015 149.055 17.225 150.145 ;
        RECT 17.400 149.055 17.660 150.205 ;
        RECT 17.835 150.130 18.005 150.860 ;
        RECT 18.260 150.695 18.430 150.885 ;
        RECT 19.275 150.785 19.505 151.605 ;
        RECT 19.675 150.805 20.005 151.435 ;
        RECT 18.175 150.365 18.430 150.695 ;
        RECT 18.260 150.155 18.430 150.365 ;
        RECT 18.710 150.335 19.065 150.705 ;
        RECT 19.255 150.365 19.585 150.615 ;
        RECT 19.755 150.205 20.005 150.805 ;
        RECT 20.175 150.785 20.385 151.605 ;
        RECT 20.615 150.930 20.875 151.435 ;
        RECT 21.055 151.225 21.385 151.605 ;
        RECT 21.565 151.055 21.735 151.435 ;
        RECT 21.995 151.060 27.340 151.605 ;
        RECT 27.515 151.060 32.860 151.605 ;
        RECT 33.060 151.215 33.390 151.605 ;
        RECT 17.835 149.225 18.090 150.130 ;
        RECT 18.260 149.985 18.975 150.155 ;
        RECT 18.260 149.055 18.590 149.815 ;
        RECT 18.805 149.225 18.975 149.985 ;
        RECT 19.275 149.055 19.505 150.195 ;
        RECT 19.675 149.225 20.005 150.205 ;
        RECT 20.175 149.055 20.385 150.195 ;
        RECT 20.615 150.130 20.785 150.930 ;
        RECT 21.070 150.885 21.735 151.055 ;
        RECT 21.070 150.630 21.240 150.885 ;
        RECT 20.955 150.300 21.240 150.630 ;
        RECT 21.475 150.335 21.805 150.705 ;
        RECT 21.070 150.155 21.240 150.300 ;
        RECT 23.580 150.230 23.920 151.060 ;
        RECT 20.615 149.225 20.885 150.130 ;
        RECT 21.070 149.985 21.735 150.155 ;
        RECT 21.055 149.055 21.385 149.815 ;
        RECT 21.565 149.225 21.735 149.985 ;
        RECT 25.400 149.490 25.750 150.740 ;
        RECT 29.100 150.230 29.440 151.060 ;
        RECT 33.560 151.045 33.785 151.425 ;
        RECT 30.920 149.490 31.270 150.740 ;
        RECT 33.045 150.365 33.285 151.015 ;
        RECT 33.455 150.865 33.785 151.045 ;
        RECT 33.455 150.195 33.630 150.865 ;
        RECT 33.985 150.695 34.215 151.315 ;
        RECT 34.395 150.875 34.695 151.605 ;
        RECT 34.965 151.055 35.135 151.435 ;
        RECT 35.350 151.225 35.680 151.605 ;
        RECT 34.965 150.885 35.680 151.055 ;
        RECT 33.800 150.365 34.215 150.695 ;
        RECT 34.395 150.365 34.690 150.695 ;
        RECT 34.875 150.335 35.230 150.705 ;
        RECT 35.510 150.695 35.680 150.885 ;
        RECT 35.850 150.860 36.105 151.435 ;
        RECT 35.510 150.365 35.765 150.695 ;
        RECT 33.045 150.005 33.630 150.195 ;
        RECT 21.995 149.055 27.340 149.490 ;
        RECT 27.515 149.055 32.860 149.490 ;
        RECT 33.045 149.235 33.320 150.005 ;
        RECT 33.800 149.835 34.695 150.165 ;
        RECT 35.510 150.155 35.680 150.365 ;
        RECT 33.490 149.665 34.695 149.835 ;
        RECT 33.490 149.235 33.820 149.665 ;
        RECT 33.990 149.055 34.185 149.495 ;
        RECT 34.365 149.235 34.695 149.665 ;
        RECT 34.965 149.985 35.680 150.155 ;
        RECT 35.935 150.130 36.105 150.860 ;
        RECT 36.280 150.765 36.540 151.605 ;
        RECT 36.715 150.835 40.225 151.605 ;
        RECT 40.395 150.855 41.605 151.605 ;
        RECT 41.775 150.880 42.065 151.605 ;
        RECT 42.235 151.060 47.580 151.605 ;
        RECT 36.715 150.315 38.365 150.835 ;
        RECT 34.965 149.225 35.135 149.985 ;
        RECT 35.350 149.055 35.680 149.815 ;
        RECT 35.850 149.225 36.105 150.130 ;
        RECT 36.280 149.055 36.540 150.205 ;
        RECT 38.535 150.145 40.225 150.665 ;
        RECT 40.395 150.315 40.915 150.855 ;
        RECT 41.085 150.145 41.605 150.685 ;
        RECT 43.820 150.230 44.160 151.060 ;
        RECT 48.215 151.020 48.525 151.435 ;
        RECT 48.720 151.225 49.050 151.605 ;
        RECT 49.220 151.265 50.625 151.435 ;
        RECT 49.220 151.035 49.390 151.265 ;
        RECT 36.715 149.055 40.225 150.145 ;
        RECT 40.395 149.055 41.605 150.145 ;
        RECT 41.775 149.055 42.065 150.220 ;
        RECT 45.640 149.490 45.990 150.740 ;
        RECT 48.215 149.905 48.385 151.020 ;
        RECT 48.695 150.865 49.390 151.035 ;
        RECT 50.455 151.035 50.625 151.265 ;
        RECT 50.895 151.205 51.225 151.605 ;
        RECT 51.465 151.035 51.635 151.435 ;
        RECT 48.695 150.695 48.865 150.865 ;
        RECT 48.555 150.365 48.865 150.695 ;
        RECT 49.035 150.365 49.370 150.695 ;
        RECT 49.640 150.365 49.835 150.940 ;
        RECT 50.095 150.695 50.285 150.925 ;
        RECT 50.455 150.865 51.635 151.035 ;
        RECT 51.930 150.865 52.545 151.435 ;
        RECT 52.715 151.095 52.930 151.605 ;
        RECT 53.160 151.095 53.440 151.425 ;
        RECT 53.620 151.095 53.860 151.605 ;
        RECT 50.095 150.365 50.440 150.695 ;
        RECT 50.750 150.365 51.225 150.695 ;
        RECT 51.480 150.365 51.665 150.695 ;
        RECT 48.695 150.195 48.865 150.365 ;
        RECT 48.695 150.025 51.635 150.195 ;
        RECT 42.235 149.055 47.580 149.490 ;
        RECT 48.215 149.265 48.555 149.905 ;
        RECT 49.145 149.685 50.705 149.855 ;
        RECT 48.725 149.055 48.970 149.515 ;
        RECT 49.145 149.225 49.395 149.685 ;
        RECT 49.585 149.055 50.255 149.435 ;
        RECT 50.455 149.225 50.705 149.685 ;
        RECT 51.465 149.225 51.635 150.025 ;
        RECT 51.930 149.845 52.245 150.865 ;
        RECT 52.415 150.195 52.585 150.695 ;
        RECT 52.835 150.365 53.100 150.925 ;
        RECT 53.270 150.195 53.440 151.095 ;
        RECT 53.610 150.365 53.965 150.925 ;
        RECT 54.215 150.795 54.455 151.605 ;
        RECT 54.625 150.795 54.955 151.435 ;
        RECT 55.125 150.795 55.395 151.605 ;
        RECT 54.195 150.365 54.545 150.615 ;
        RECT 54.715 150.195 54.885 150.795 ;
        RECT 55.055 150.365 55.405 150.615 ;
        RECT 52.415 150.025 53.840 150.195 ;
        RECT 51.930 149.225 52.465 149.845 ;
        RECT 52.635 149.055 52.965 149.855 ;
        RECT 53.450 149.850 53.840 150.025 ;
        RECT 54.205 150.025 54.885 150.195 ;
        RECT 54.205 149.240 54.535 150.025 ;
        RECT 55.065 149.055 55.395 150.195 ;
        RECT 55.575 149.225 55.855 151.325 ;
        RECT 56.085 151.145 56.255 151.605 ;
        RECT 56.525 151.215 57.775 151.395 ;
        RECT 56.910 150.975 57.275 151.045 ;
        RECT 56.025 150.795 57.275 150.975 ;
        RECT 57.445 150.995 57.775 151.215 ;
        RECT 57.945 151.165 58.115 151.605 ;
        RECT 58.285 150.995 58.625 151.410 ;
        RECT 57.445 150.825 58.625 150.995 ;
        RECT 58.795 150.805 59.105 151.605 ;
        RECT 59.310 150.805 60.005 151.435 ;
        RECT 60.175 151.060 65.520 151.605 ;
        RECT 56.025 150.195 56.300 150.795 ;
        RECT 56.470 150.365 56.825 150.615 ;
        RECT 57.020 150.585 57.485 150.615 ;
        RECT 57.015 150.415 57.485 150.585 ;
        RECT 57.020 150.365 57.485 150.415 ;
        RECT 57.655 150.365 57.985 150.615 ;
        RECT 58.160 150.415 58.625 150.615 ;
        RECT 58.805 150.365 59.140 150.635 ;
        RECT 57.805 150.245 57.985 150.365 ;
        RECT 56.025 149.985 57.635 150.195 ;
        RECT 57.805 150.075 58.135 150.245 ;
        RECT 57.225 149.885 57.635 149.985 ;
        RECT 56.045 149.055 56.830 149.815 ;
        RECT 57.225 149.225 57.610 149.885 ;
        RECT 57.935 149.285 58.135 150.075 ;
        RECT 58.305 149.055 58.625 150.235 ;
        RECT 59.310 150.205 59.480 150.805 ;
        RECT 59.650 150.365 59.985 150.615 ;
        RECT 61.760 150.230 62.100 151.060 ;
        RECT 65.705 150.875 66.005 151.605 ;
        RECT 58.795 149.055 59.075 150.195 ;
        RECT 59.245 149.225 59.575 150.205 ;
        RECT 59.745 149.055 60.005 150.195 ;
        RECT 63.580 149.490 63.930 150.740 ;
        RECT 66.185 150.695 66.415 151.315 ;
        RECT 66.615 151.045 66.840 151.425 ;
        RECT 67.010 151.215 67.340 151.605 ;
        RECT 66.615 150.865 66.945 151.045 ;
        RECT 65.710 150.365 66.005 150.695 ;
        RECT 66.185 150.365 66.600 150.695 ;
        RECT 66.770 150.195 66.945 150.865 ;
        RECT 67.115 150.365 67.355 151.015 ;
        RECT 67.535 150.880 67.825 151.605 ;
        RECT 67.995 151.060 73.340 151.605 ;
        RECT 73.515 151.060 78.860 151.605 ;
        RECT 79.035 151.060 84.380 151.605 ;
        RECT 69.580 150.230 69.920 151.060 ;
        RECT 65.705 149.835 66.600 150.165 ;
        RECT 66.770 150.005 67.355 150.195 ;
        RECT 65.705 149.665 66.910 149.835 ;
        RECT 60.175 149.055 65.520 149.490 ;
        RECT 65.705 149.235 66.035 149.665 ;
        RECT 66.215 149.055 66.410 149.495 ;
        RECT 66.580 149.235 66.910 149.665 ;
        RECT 67.080 149.235 67.355 150.005 ;
        RECT 67.535 149.055 67.825 150.220 ;
        RECT 71.400 149.490 71.750 150.740 ;
        RECT 75.100 150.230 75.440 151.060 ;
        RECT 76.920 149.490 77.270 150.740 ;
        RECT 80.620 150.230 80.960 151.060 ;
        RECT 84.555 150.930 84.815 151.435 ;
        RECT 84.995 151.225 85.325 151.605 ;
        RECT 85.505 151.055 85.675 151.435 ;
        RECT 82.440 149.490 82.790 150.740 ;
        RECT 84.555 150.130 84.725 150.930 ;
        RECT 85.010 150.885 85.675 151.055 ;
        RECT 85.010 150.630 85.180 150.885 ;
        RECT 85.935 150.855 87.145 151.605 ;
        RECT 84.895 150.300 85.180 150.630 ;
        RECT 85.415 150.335 85.745 150.705 ;
        RECT 85.010 150.155 85.180 150.300 ;
        RECT 67.995 149.055 73.340 149.490 ;
        RECT 73.515 149.055 78.860 149.490 ;
        RECT 79.035 149.055 84.380 149.490 ;
        RECT 84.555 149.225 84.825 150.130 ;
        RECT 85.010 149.985 85.675 150.155 ;
        RECT 84.995 149.055 85.325 149.815 ;
        RECT 85.505 149.225 85.675 149.985 ;
        RECT 85.935 150.145 86.455 150.685 ;
        RECT 86.625 150.315 87.145 150.855 ;
        RECT 85.935 149.055 87.145 150.145 ;
        RECT 15.930 148.885 87.230 149.055 ;
        RECT 16.015 147.795 17.225 148.885 ;
        RECT 17.395 148.450 22.740 148.885 ;
        RECT 22.915 148.450 28.260 148.885 ;
        RECT 16.015 147.085 16.535 147.625 ;
        RECT 16.705 147.255 17.225 147.795 ;
        RECT 16.015 146.335 17.225 147.085 ;
        RECT 18.980 146.880 19.320 147.710 ;
        RECT 20.800 147.200 21.150 148.450 ;
        RECT 24.500 146.880 24.840 147.710 ;
        RECT 26.320 147.200 26.670 148.450 ;
        RECT 28.895 147.720 29.185 148.885 ;
        RECT 29.355 147.795 31.025 148.885 ;
        RECT 29.355 147.105 30.105 147.625 ;
        RECT 30.275 147.275 31.025 147.795 ;
        RECT 31.655 147.745 31.935 148.885 ;
        RECT 32.105 147.735 32.435 148.715 ;
        RECT 32.605 147.745 32.865 148.885 ;
        RECT 33.040 148.045 33.360 148.885 ;
        RECT 33.530 147.865 33.730 148.655 ;
        RECT 34.055 147.955 34.440 148.715 ;
        RECT 34.835 148.125 35.635 148.885 ;
        RECT 32.170 147.695 32.345 147.735 ;
        RECT 31.665 147.305 32.000 147.575 ;
        RECT 32.170 147.135 32.340 147.695 ;
        RECT 32.510 147.325 32.845 147.575 ;
        RECT 33.040 147.525 33.360 147.865 ;
        RECT 33.530 147.695 33.885 147.865 ;
        RECT 34.055 147.745 35.655 147.955 ;
        RECT 33.705 147.575 33.885 147.695 ;
        RECT 33.040 147.325 33.535 147.525 ;
        RECT 33.705 147.325 34.035 147.575 ;
        RECT 34.205 147.325 34.670 147.575 ;
        RECT 34.840 147.325 35.195 147.575 ;
        RECT 35.375 147.145 35.655 147.745 ;
        RECT 17.395 146.335 22.740 146.880 ;
        RECT 22.915 146.335 28.260 146.880 ;
        RECT 28.895 146.335 29.185 147.060 ;
        RECT 29.355 146.335 31.025 147.105 ;
        RECT 31.655 146.335 31.965 147.135 ;
        RECT 32.170 146.505 32.865 147.135 ;
        RECT 33.040 147.075 34.070 147.115 ;
        RECT 33.040 146.945 34.240 147.075 ;
        RECT 33.040 146.530 33.375 146.945 ;
        RECT 33.545 146.335 33.715 146.775 ;
        RECT 33.900 146.725 34.240 146.945 ;
        RECT 34.415 146.965 35.655 147.145 ;
        RECT 34.415 146.895 34.780 146.965 ;
        RECT 33.900 146.545 35.165 146.725 ;
        RECT 35.425 146.335 35.605 146.795 ;
        RECT 35.825 146.615 36.040 148.715 ;
        RECT 36.265 147.695 36.515 148.885 ;
        RECT 36.715 147.745 37.100 148.705 ;
        RECT 37.315 148.085 37.605 148.885 ;
        RECT 37.775 148.545 39.140 148.715 ;
        RECT 37.775 147.915 37.945 148.545 ;
        RECT 37.270 147.745 37.945 147.915 ;
        RECT 36.275 146.335 36.445 147.135 ;
        RECT 36.715 147.075 36.890 147.745 ;
        RECT 37.270 147.575 37.440 147.745 ;
        RECT 38.115 147.575 38.440 148.375 ;
        RECT 38.810 148.335 39.140 148.545 ;
        RECT 38.810 148.085 39.765 148.335 ;
        RECT 37.075 147.325 37.440 147.575 ;
        RECT 37.635 147.325 37.885 147.575 ;
        RECT 37.075 147.245 37.265 147.325 ;
        RECT 37.635 147.245 37.805 147.325 ;
        RECT 38.095 147.245 38.440 147.575 ;
        RECT 38.610 147.245 38.885 147.910 ;
        RECT 39.070 147.245 39.425 147.910 ;
        RECT 39.595 147.075 39.765 148.085 ;
        RECT 39.935 147.745 40.225 148.885 ;
        RECT 40.395 147.795 42.985 148.885 ;
        RECT 39.950 147.245 40.225 147.575 ;
        RECT 36.715 146.505 37.225 147.075 ;
        RECT 37.770 146.905 39.170 147.075 ;
        RECT 37.395 146.335 37.565 146.895 ;
        RECT 37.770 146.505 38.100 146.905 ;
        RECT 38.275 146.335 38.605 146.735 ;
        RECT 38.840 146.715 39.170 146.905 ;
        RECT 39.340 146.885 39.765 147.075 ;
        RECT 40.395 147.105 41.605 147.625 ;
        RECT 41.775 147.275 42.985 147.795 ;
        RECT 43.155 147.745 43.485 148.885 ;
        RECT 43.655 148.255 44.010 148.715 ;
        RECT 44.180 148.425 44.755 148.885 ;
        RECT 44.925 148.255 45.255 148.715 ;
        RECT 43.655 148.085 45.255 148.255 ;
        RECT 45.455 148.085 45.710 148.885 ;
        RECT 46.375 148.450 51.720 148.885 ;
        RECT 43.655 147.745 43.930 148.085 ;
        RECT 44.110 147.525 44.300 147.905 ;
        RECT 43.155 147.325 44.300 147.525 ;
        RECT 44.480 147.155 44.760 148.085 ;
        RECT 45.880 147.915 46.180 148.110 ;
        RECT 44.930 147.745 46.180 147.915 ;
        RECT 44.930 147.325 45.260 147.745 ;
        RECT 45.490 147.245 45.835 147.575 ;
        RECT 39.935 146.715 40.225 146.985 ;
        RECT 38.840 146.505 40.225 146.715 ;
        RECT 40.395 146.335 42.985 147.105 ;
        RECT 43.155 146.945 44.265 147.155 ;
        RECT 43.155 146.505 43.505 146.945 ;
        RECT 43.675 146.335 43.845 146.775 ;
        RECT 44.015 146.715 44.265 146.945 ;
        RECT 44.435 147.055 44.760 147.155 ;
        RECT 44.435 146.885 44.765 147.055 ;
        RECT 44.935 146.715 45.210 147.155 ;
        RECT 46.010 147.090 46.180 147.745 ;
        RECT 44.015 146.505 45.210 146.715 ;
        RECT 45.445 146.335 45.775 147.075 ;
        RECT 45.945 146.760 46.180 147.090 ;
        RECT 47.960 146.880 48.300 147.710 ;
        RECT 49.780 147.200 50.130 148.450 ;
        RECT 51.895 147.795 54.485 148.885 ;
        RECT 51.895 147.105 53.105 147.625 ;
        RECT 53.275 147.275 54.485 147.795 ;
        RECT 54.655 147.720 54.945 148.885 ;
        RECT 55.575 148.285 55.835 148.705 ;
        RECT 56.005 148.455 56.335 148.885 ;
        RECT 57.000 148.455 57.745 148.625 ;
        RECT 57.970 148.545 58.610 148.705 ;
        RECT 55.575 148.115 57.405 148.285 ;
        RECT 46.375 146.335 51.720 146.880 ;
        RECT 51.895 146.335 54.485 147.105 ;
        RECT 55.575 147.075 55.745 148.115 ;
        RECT 55.915 147.245 56.265 147.945 ;
        RECT 56.480 147.775 57.065 147.945 ;
        RECT 56.435 147.245 56.725 147.575 ;
        RECT 56.895 147.495 57.065 147.775 ;
        RECT 57.235 147.835 57.405 148.115 ;
        RECT 57.575 148.205 57.745 148.455 ;
        RECT 57.935 148.375 58.610 148.545 ;
        RECT 57.575 148.035 58.610 148.205 ;
        RECT 58.780 148.085 59.060 148.885 ;
        RECT 58.440 147.915 58.610 148.035 ;
        RECT 57.235 147.665 57.885 147.835 ;
        RECT 58.440 147.745 59.100 147.915 ;
        RECT 59.270 147.745 59.545 148.715 ;
        RECT 59.805 147.955 59.975 148.715 ;
        RECT 60.190 148.125 60.520 148.885 ;
        RECT 59.805 147.785 60.520 147.955 ;
        RECT 60.690 147.810 60.945 148.715 ;
        RECT 56.895 147.325 57.320 147.495 ;
        RECT 56.895 147.075 57.065 147.325 ;
        RECT 57.715 147.245 57.885 147.665 ;
        RECT 58.930 147.575 59.100 147.745 ;
        RECT 58.105 147.245 58.760 147.575 ;
        RECT 58.930 147.245 59.205 147.575 ;
        RECT 58.930 147.075 59.100 147.245 ;
        RECT 54.655 146.335 54.945 147.060 ;
        RECT 55.575 146.700 55.890 147.075 ;
        RECT 56.145 146.335 56.315 147.075 ;
        RECT 56.565 146.905 57.065 147.075 ;
        RECT 57.505 146.905 59.100 147.075 ;
        RECT 59.375 147.010 59.545 147.745 ;
        RECT 59.715 147.235 60.070 147.605 ;
        RECT 60.350 147.575 60.520 147.785 ;
        RECT 60.350 147.245 60.605 147.575 ;
        RECT 60.350 147.055 60.520 147.245 ;
        RECT 60.775 147.080 60.945 147.810 ;
        RECT 61.120 147.735 61.380 148.885 ;
        RECT 61.560 148.315 61.880 148.715 ;
        RECT 61.560 147.865 61.730 148.315 ;
        RECT 62.050 148.085 62.360 148.885 ;
        RECT 62.530 148.255 62.860 148.715 ;
        RECT 63.030 148.425 63.200 148.885 ;
        RECT 63.370 148.255 63.700 148.715 ;
        RECT 63.870 148.425 64.120 148.885 ;
        RECT 64.310 148.425 64.560 148.885 ;
        RECT 62.530 148.205 63.700 148.255 ;
        RECT 64.730 148.255 64.980 148.715 ;
        RECT 65.230 148.425 65.520 148.885 ;
        RECT 65.695 148.450 71.040 148.885 ;
        RECT 71.215 148.450 76.560 148.885 ;
        RECT 64.730 148.205 65.520 148.255 ;
        RECT 62.530 148.035 65.520 148.205 ;
        RECT 61.560 147.695 65.120 147.865 ;
        RECT 56.565 146.700 56.735 146.905 ;
        RECT 56.960 146.335 57.335 146.735 ;
        RECT 57.505 146.555 57.675 146.905 ;
        RECT 57.860 146.335 58.190 146.735 ;
        RECT 58.360 146.555 58.530 146.905 ;
        RECT 58.700 146.335 59.080 146.735 ;
        RECT 59.270 146.665 59.545 147.010 ;
        RECT 59.805 146.885 60.520 147.055 ;
        RECT 59.805 146.505 59.975 146.885 ;
        RECT 60.190 146.335 60.520 146.715 ;
        RECT 60.690 146.505 60.945 147.080 ;
        RECT 61.120 146.335 61.380 147.175 ;
        RECT 61.560 146.905 61.730 147.695 ;
        RECT 61.900 147.325 62.250 147.525 ;
        RECT 62.530 147.325 63.210 147.525 ;
        RECT 63.420 147.325 64.610 147.525 ;
        RECT 64.790 147.325 65.120 147.695 ;
        RECT 65.320 147.155 65.520 148.035 ;
        RECT 61.560 146.505 61.880 146.905 ;
        RECT 62.050 146.335 62.360 147.155 ;
        RECT 62.530 146.965 64.220 147.155 ;
        RECT 62.530 146.505 62.860 146.965 ;
        RECT 63.470 146.885 64.220 146.965 ;
        RECT 63.030 146.335 63.280 146.795 ;
        RECT 64.390 146.715 64.560 147.155 ;
        RECT 64.730 146.885 65.520 147.155 ;
        RECT 67.280 146.880 67.620 147.710 ;
        RECT 69.100 147.200 69.450 148.450 ;
        RECT 72.800 146.880 73.140 147.710 ;
        RECT 74.620 147.200 74.970 148.450 ;
        RECT 76.735 147.795 80.245 148.885 ;
        RECT 76.735 147.105 78.385 147.625 ;
        RECT 78.555 147.275 80.245 147.795 ;
        RECT 80.415 147.720 80.705 148.885 ;
        RECT 80.875 147.795 83.465 148.885 ;
        RECT 84.100 148.460 84.435 148.885 ;
        RECT 84.605 148.280 84.790 148.685 ;
        RECT 80.875 147.105 82.085 147.625 ;
        RECT 82.255 147.275 83.465 147.795 ;
        RECT 84.125 148.105 84.790 148.280 ;
        RECT 84.995 148.105 85.325 148.885 ;
        RECT 63.470 146.505 65.520 146.715 ;
        RECT 65.695 146.335 71.040 146.880 ;
        RECT 71.215 146.335 76.560 146.880 ;
        RECT 76.735 146.335 80.245 147.105 ;
        RECT 80.415 146.335 80.705 147.060 ;
        RECT 80.875 146.335 83.465 147.105 ;
        RECT 84.125 147.075 84.465 148.105 ;
        RECT 85.495 147.915 85.765 148.685 ;
        RECT 84.635 147.745 85.765 147.915 ;
        RECT 84.635 147.245 84.885 147.745 ;
        RECT 84.125 146.905 84.810 147.075 ;
        RECT 85.065 146.995 85.425 147.575 ;
        RECT 84.100 146.335 84.435 146.735 ;
        RECT 84.605 146.505 84.810 146.905 ;
        RECT 85.595 146.835 85.765 147.745 ;
        RECT 85.935 147.795 87.145 148.885 ;
        RECT 85.935 147.255 86.455 147.795 ;
        RECT 86.625 147.085 87.145 147.625 ;
        RECT 85.020 146.335 85.295 146.815 ;
        RECT 85.505 146.505 85.765 146.835 ;
        RECT 85.935 146.335 87.145 147.085 ;
        RECT 15.930 146.165 87.230 146.335 ;
        RECT 16.015 145.415 17.225 146.165 ;
        RECT 17.395 145.620 22.740 146.165 ;
        RECT 22.915 145.620 28.260 146.165 ;
        RECT 28.435 145.620 33.780 146.165 ;
        RECT 34.045 145.825 34.215 145.860 ;
        RECT 34.015 145.655 34.215 145.825 ;
        RECT 16.015 144.875 16.535 145.415 ;
        RECT 16.705 144.705 17.225 145.245 ;
        RECT 18.980 144.790 19.320 145.620 ;
        RECT 16.015 143.615 17.225 144.705 ;
        RECT 20.800 144.050 21.150 145.300 ;
        RECT 24.500 144.790 24.840 145.620 ;
        RECT 26.320 144.050 26.670 145.300 ;
        RECT 30.020 144.790 30.360 145.620 ;
        RECT 31.840 144.050 32.190 145.300 ;
        RECT 34.045 145.295 34.215 145.655 ;
        RECT 34.405 145.635 34.635 145.940 ;
        RECT 34.805 145.805 35.135 146.165 ;
        RECT 35.330 145.635 35.620 145.985 ;
        RECT 34.405 145.465 35.620 145.635 ;
        RECT 35.795 145.705 36.355 145.995 ;
        RECT 36.525 145.705 36.775 146.165 ;
        RECT 34.045 145.125 34.565 145.295 ;
        RECT 33.960 144.595 34.205 144.955 ;
        RECT 34.395 144.745 34.565 145.125 ;
        RECT 34.735 144.925 35.120 145.255 ;
        RECT 35.300 145.145 35.560 145.255 ;
        RECT 35.300 144.975 35.565 145.145 ;
        RECT 35.300 144.925 35.560 144.975 ;
        RECT 34.395 144.465 34.745 144.745 ;
        RECT 17.395 143.615 22.740 144.050 ;
        RECT 22.915 143.615 28.260 144.050 ;
        RECT 28.435 143.615 33.780 144.050 ;
        RECT 33.960 143.615 34.215 144.415 ;
        RECT 34.415 143.785 34.745 144.465 ;
        RECT 34.925 143.875 35.120 144.925 ;
        RECT 35.300 143.615 35.620 144.755 ;
        RECT 35.795 144.335 36.045 145.705 ;
        RECT 37.395 145.535 37.725 145.895 ;
        RECT 39.035 145.655 39.275 146.165 ;
        RECT 39.445 145.655 39.735 145.995 ;
        RECT 39.965 145.655 40.280 146.165 ;
        RECT 36.335 145.345 37.725 145.535 ;
        RECT 36.335 145.255 36.505 145.345 ;
        RECT 36.215 144.925 36.505 145.255 ;
        RECT 36.675 144.925 37.015 145.175 ;
        RECT 37.235 144.925 37.910 145.175 ;
        RECT 39.080 145.145 39.275 145.485 ;
        RECT 39.075 144.975 39.275 145.145 ;
        RECT 39.080 144.925 39.275 144.975 ;
        RECT 36.335 144.675 36.505 144.925 ;
        RECT 36.335 144.505 37.275 144.675 ;
        RECT 37.645 144.565 37.910 144.925 ;
        RECT 39.445 144.755 39.625 145.655 ;
        RECT 40.450 145.595 40.620 145.865 ;
        RECT 40.790 145.765 41.120 146.165 ;
        RECT 39.795 144.925 40.205 145.485 ;
        RECT 40.450 145.425 41.145 145.595 ;
        RECT 41.775 145.440 42.065 146.165 ;
        RECT 42.240 145.765 42.575 146.165 ;
        RECT 42.745 145.595 42.950 145.995 ;
        RECT 43.160 145.685 43.435 146.165 ;
        RECT 43.645 145.665 43.905 145.995 ;
        RECT 40.375 144.755 40.545 145.255 ;
        RECT 39.085 144.585 40.545 144.755 ;
        RECT 35.795 143.785 36.255 144.335 ;
        RECT 36.445 143.615 36.775 144.335 ;
        RECT 36.975 143.955 37.275 144.505 ;
        RECT 39.085 144.410 39.445 144.585 ;
        RECT 40.715 144.415 41.145 145.425 ;
        RECT 42.265 145.425 42.950 145.595 ;
        RECT 37.445 143.615 37.725 144.285 ;
        RECT 40.030 143.615 40.200 144.415 ;
        RECT 40.370 144.245 41.145 144.415 ;
        RECT 40.370 143.785 40.700 144.245 ;
        RECT 40.870 143.615 41.040 144.075 ;
        RECT 41.775 143.615 42.065 144.780 ;
        RECT 42.265 144.395 42.605 145.425 ;
        RECT 42.775 144.755 43.025 145.255 ;
        RECT 43.205 144.925 43.565 145.505 ;
        RECT 43.735 144.755 43.905 145.665 ;
        RECT 44.165 145.615 44.335 145.995 ;
        RECT 44.515 145.785 44.845 146.165 ;
        RECT 44.165 145.445 44.830 145.615 ;
        RECT 45.025 145.490 45.285 145.995 ;
        RECT 45.455 145.620 50.800 146.165 ;
        RECT 50.975 145.620 56.320 146.165 ;
        RECT 44.095 144.895 44.425 145.265 ;
        RECT 44.660 145.190 44.830 145.445 ;
        RECT 42.775 144.585 43.905 144.755 ;
        RECT 44.660 144.860 44.945 145.190 ;
        RECT 44.660 144.715 44.830 144.860 ;
        RECT 42.265 144.220 42.930 144.395 ;
        RECT 42.240 143.615 42.575 144.040 ;
        RECT 42.745 143.815 42.930 144.220 ;
        RECT 43.135 143.615 43.465 144.395 ;
        RECT 43.635 143.815 43.905 144.585 ;
        RECT 44.165 144.545 44.830 144.715 ;
        RECT 45.115 144.690 45.285 145.490 ;
        RECT 47.040 144.790 47.380 145.620 ;
        RECT 44.165 143.785 44.335 144.545 ;
        RECT 44.515 143.615 44.845 144.375 ;
        RECT 45.015 143.785 45.285 144.690 ;
        RECT 48.860 144.050 49.210 145.300 ;
        RECT 52.560 144.790 52.900 145.620 ;
        RECT 56.495 145.395 60.005 146.165 ;
        RECT 60.640 145.785 62.690 145.995 ;
        RECT 54.380 144.050 54.730 145.300 ;
        RECT 56.495 144.875 58.145 145.395 ;
        RECT 60.640 145.345 61.430 145.615 ;
        RECT 61.600 145.345 61.770 145.785 ;
        RECT 62.880 145.705 63.130 146.165 ;
        RECT 61.940 145.535 62.690 145.615 ;
        RECT 63.300 145.535 63.630 145.995 ;
        RECT 61.940 145.345 63.630 145.535 ;
        RECT 63.800 145.345 64.110 146.165 ;
        RECT 64.280 145.595 64.600 145.995 ;
        RECT 60.640 145.315 60.865 145.345 ;
        RECT 58.315 144.705 60.005 145.225 ;
        RECT 45.455 143.615 50.800 144.050 ;
        RECT 50.975 143.615 56.320 144.050 ;
        RECT 56.495 143.615 60.005 144.705 ;
        RECT 60.640 144.465 60.840 145.315 ;
        RECT 61.040 144.805 61.370 145.175 ;
        RECT 61.550 144.975 62.740 145.175 ;
        RECT 62.950 144.975 63.630 145.175 ;
        RECT 63.910 144.975 64.260 145.175 ;
        RECT 64.430 144.805 64.600 145.595 ;
        RECT 64.775 145.395 67.365 146.165 ;
        RECT 67.535 145.440 67.825 146.165 ;
        RECT 67.995 145.620 73.340 146.165 ;
        RECT 73.515 145.620 78.860 146.165 ;
        RECT 79.035 145.620 84.380 146.165 ;
        RECT 64.775 144.875 65.985 145.395 ;
        RECT 61.040 144.635 64.600 144.805 ;
        RECT 66.155 144.705 67.365 145.225 ;
        RECT 69.580 144.790 69.920 145.620 ;
        RECT 60.640 144.295 63.630 144.465 ;
        RECT 60.640 144.245 61.430 144.295 ;
        RECT 60.640 143.615 60.930 144.075 ;
        RECT 61.180 143.785 61.430 144.245 ;
        RECT 62.460 144.245 63.630 144.295 ;
        RECT 61.600 143.615 61.850 144.075 ;
        RECT 62.040 143.615 62.290 144.075 ;
        RECT 62.460 143.785 62.790 144.245 ;
        RECT 62.960 143.615 63.130 144.075 ;
        RECT 63.300 143.785 63.630 144.245 ;
        RECT 63.800 143.615 64.110 144.415 ;
        RECT 64.430 144.185 64.600 144.635 ;
        RECT 64.280 143.785 64.600 144.185 ;
        RECT 64.775 143.615 67.365 144.705 ;
        RECT 67.535 143.615 67.825 144.780 ;
        RECT 71.400 144.050 71.750 145.300 ;
        RECT 75.100 144.790 75.440 145.620 ;
        RECT 76.920 144.050 77.270 145.300 ;
        RECT 80.620 144.790 80.960 145.620 ;
        RECT 84.735 145.505 85.075 146.165 ;
        RECT 82.440 144.050 82.790 145.300 ;
        RECT 67.995 143.615 73.340 144.050 ;
        RECT 73.515 143.615 78.860 144.050 ;
        RECT 79.035 143.615 84.380 144.050 ;
        RECT 84.555 143.785 85.075 145.335 ;
        RECT 85.245 144.510 85.765 145.995 ;
        RECT 85.935 145.415 87.145 146.165 ;
        RECT 85.935 144.705 86.455 145.245 ;
        RECT 86.625 144.875 87.145 145.415 ;
        RECT 85.245 143.615 85.575 144.340 ;
        RECT 85.935 143.615 87.145 144.705 ;
        RECT 15.930 143.445 87.230 143.615 ;
        RECT 16.015 142.355 17.225 143.445 ;
        RECT 17.395 143.010 22.740 143.445 ;
        RECT 16.015 141.645 16.535 142.185 ;
        RECT 16.705 141.815 17.225 142.355 ;
        RECT 16.015 140.895 17.225 141.645 ;
        RECT 18.980 141.440 19.320 142.270 ;
        RECT 20.800 141.760 21.150 143.010 ;
        RECT 23.835 141.725 24.355 143.275 ;
        RECT 24.525 142.720 24.855 143.445 ;
        RECT 17.395 140.895 22.740 141.440 ;
        RECT 24.015 140.895 24.355 141.555 ;
        RECT 24.525 141.065 25.045 142.550 ;
        RECT 25.215 142.355 28.725 143.445 ;
        RECT 25.215 141.665 26.865 142.185 ;
        RECT 27.035 141.835 28.725 142.355 ;
        RECT 28.895 142.280 29.185 143.445 ;
        RECT 29.355 142.355 32.865 143.445 ;
        RECT 29.355 141.665 31.005 142.185 ;
        RECT 31.175 141.835 32.865 142.355 ;
        RECT 33.495 142.370 33.765 143.275 ;
        RECT 33.935 142.685 34.265 143.445 ;
        RECT 34.445 142.515 34.615 143.275 ;
        RECT 25.215 140.895 28.725 141.665 ;
        RECT 28.895 140.895 29.185 141.620 ;
        RECT 29.355 140.895 32.865 141.665 ;
        RECT 33.495 141.570 33.665 142.370 ;
        RECT 33.950 142.345 34.615 142.515 ;
        RECT 34.875 142.355 36.545 143.445 ;
        RECT 33.950 142.200 34.120 142.345 ;
        RECT 33.835 141.870 34.120 142.200 ;
        RECT 33.950 141.615 34.120 141.870 ;
        RECT 34.355 141.795 34.685 142.165 ;
        RECT 34.875 141.665 35.625 142.185 ;
        RECT 35.795 141.835 36.545 142.355 ;
        RECT 36.805 142.515 36.975 143.275 ;
        RECT 37.190 142.685 37.520 143.445 ;
        RECT 36.805 142.345 37.520 142.515 ;
        RECT 37.690 142.370 37.945 143.275 ;
        RECT 36.715 141.795 37.070 142.165 ;
        RECT 37.350 142.135 37.520 142.345 ;
        RECT 37.350 141.805 37.605 142.135 ;
        RECT 33.495 141.065 33.755 141.570 ;
        RECT 33.950 141.445 34.615 141.615 ;
        RECT 33.935 140.895 34.265 141.275 ;
        RECT 34.445 141.065 34.615 141.445 ;
        RECT 34.875 140.895 36.545 141.665 ;
        RECT 37.350 141.615 37.520 141.805 ;
        RECT 37.775 141.640 37.945 142.370 ;
        RECT 38.120 142.295 38.380 143.445 ;
        RECT 38.555 142.305 38.815 143.445 ;
        RECT 38.985 142.295 39.315 143.275 ;
        RECT 39.485 142.305 39.765 143.445 ;
        RECT 40.015 142.515 40.195 143.275 ;
        RECT 40.375 142.685 40.705 143.445 ;
        RECT 40.015 142.345 40.690 142.515 ;
        RECT 40.875 142.370 41.145 143.275 ;
        RECT 38.575 141.885 38.910 142.135 ;
        RECT 36.805 141.445 37.520 141.615 ;
        RECT 36.805 141.065 36.975 141.445 ;
        RECT 37.190 140.895 37.520 141.275 ;
        RECT 37.690 141.065 37.945 141.640 ;
        RECT 38.120 140.895 38.380 141.735 ;
        RECT 39.080 141.695 39.250 142.295 ;
        RECT 40.520 142.200 40.690 142.345 ;
        RECT 39.420 141.865 39.755 142.135 ;
        RECT 39.955 141.795 40.295 142.165 ;
        RECT 40.520 141.870 40.795 142.200 ;
        RECT 38.555 141.065 39.250 141.695 ;
        RECT 39.455 140.895 39.765 141.695 ;
        RECT 40.520 141.615 40.690 141.870 ;
        RECT 40.025 141.445 40.690 141.615 ;
        RECT 40.965 141.570 41.145 142.370 ;
        RECT 41.775 142.280 42.065 143.445 ;
        RECT 43.155 142.475 43.425 143.245 ;
        RECT 43.595 142.665 43.925 143.445 ;
        RECT 44.130 142.840 44.315 143.245 ;
        RECT 44.485 143.020 44.820 143.445 ;
        RECT 44.130 142.665 44.795 142.840 ;
        RECT 43.155 142.305 44.285 142.475 ;
        RECT 40.025 141.065 40.195 141.445 ;
        RECT 40.375 140.895 40.705 141.275 ;
        RECT 40.885 141.065 41.145 141.570 ;
        RECT 41.775 140.895 42.065 141.620 ;
        RECT 43.155 141.395 43.325 142.305 ;
        RECT 43.495 141.555 43.855 142.135 ;
        RECT 44.035 141.805 44.285 142.305 ;
        RECT 44.455 141.635 44.795 142.665 ;
        RECT 44.995 142.355 46.205 143.445 ;
        RECT 44.110 141.465 44.795 141.635 ;
        RECT 44.995 141.645 45.515 142.185 ;
        RECT 45.685 141.815 46.205 142.355 ;
        RECT 46.465 142.515 46.635 143.275 ;
        RECT 46.850 142.685 47.180 143.445 ;
        RECT 46.465 142.345 47.180 142.515 ;
        RECT 47.350 142.370 47.605 143.275 ;
        RECT 46.375 141.795 46.730 142.165 ;
        RECT 47.010 142.135 47.180 142.345 ;
        RECT 47.010 141.805 47.265 142.135 ;
        RECT 43.155 141.065 43.415 141.395 ;
        RECT 43.625 140.895 43.900 141.375 ;
        RECT 44.110 141.065 44.315 141.465 ;
        RECT 44.485 140.895 44.820 141.295 ;
        RECT 44.995 140.895 46.205 141.645 ;
        RECT 47.010 141.615 47.180 141.805 ;
        RECT 47.435 141.640 47.605 142.370 ;
        RECT 47.780 142.295 48.040 143.445 ;
        RECT 48.215 143.010 53.560 143.445 ;
        RECT 46.465 141.445 47.180 141.615 ;
        RECT 46.465 141.065 46.635 141.445 ;
        RECT 46.850 140.895 47.180 141.275 ;
        RECT 47.350 141.065 47.605 141.640 ;
        RECT 47.780 140.895 48.040 141.735 ;
        RECT 49.800 141.440 50.140 142.270 ;
        RECT 51.620 141.760 51.970 143.010 ;
        RECT 54.655 142.280 54.945 143.445 ;
        RECT 55.115 143.010 60.460 143.445 ;
        RECT 60.635 143.010 65.980 143.445 ;
        RECT 48.215 140.895 53.560 141.440 ;
        RECT 54.655 140.895 54.945 141.620 ;
        RECT 56.700 141.440 57.040 142.270 ;
        RECT 58.520 141.760 58.870 143.010 ;
        RECT 62.220 141.440 62.560 142.270 ;
        RECT 64.040 141.760 64.390 143.010 ;
        RECT 66.155 142.355 67.365 143.445 ;
        RECT 66.155 141.645 66.675 142.185 ;
        RECT 66.845 141.815 67.365 142.355 ;
        RECT 67.535 142.280 67.825 143.445 ;
        RECT 67.995 143.010 73.340 143.445 ;
        RECT 73.515 143.010 78.860 143.445 ;
        RECT 55.115 140.895 60.460 141.440 ;
        RECT 60.635 140.895 65.980 141.440 ;
        RECT 66.155 140.895 67.365 141.645 ;
        RECT 67.535 140.895 67.825 141.620 ;
        RECT 69.580 141.440 69.920 142.270 ;
        RECT 71.400 141.760 71.750 143.010 ;
        RECT 75.100 141.440 75.440 142.270 ;
        RECT 76.920 141.760 77.270 143.010 ;
        RECT 79.035 142.355 80.245 143.445 ;
        RECT 79.035 141.645 79.555 142.185 ;
        RECT 79.725 141.815 80.245 142.355 ;
        RECT 80.415 142.280 80.705 143.445 ;
        RECT 80.875 142.355 84.385 143.445 ;
        RECT 84.555 142.355 85.765 143.445 ;
        RECT 80.875 141.665 82.525 142.185 ;
        RECT 82.695 141.835 84.385 142.355 ;
        RECT 67.995 140.895 73.340 141.440 ;
        RECT 73.515 140.895 78.860 141.440 ;
        RECT 79.035 140.895 80.245 141.645 ;
        RECT 80.415 140.895 80.705 141.620 ;
        RECT 80.875 140.895 84.385 141.665 ;
        RECT 84.555 141.645 85.075 142.185 ;
        RECT 85.245 141.815 85.765 142.355 ;
        RECT 85.935 142.355 87.145 143.445 ;
        RECT 85.935 141.815 86.455 142.355 ;
        RECT 86.625 141.645 87.145 142.185 ;
        RECT 84.555 140.895 85.765 141.645 ;
        RECT 85.935 140.895 87.145 141.645 ;
        RECT 15.930 140.725 87.230 140.895 ;
      LAYER met1 ;
        RECT 19.680 215.850 20.000 215.910 ;
        RECT 39.460 215.850 39.780 215.910 ;
        RECT 19.680 215.710 39.780 215.850 ;
        RECT 19.680 215.650 20.000 215.710 ;
        RECT 39.460 215.650 39.780 215.710 ;
        RECT 22.440 214.830 22.760 214.890 ;
        RECT 78.100 214.830 78.420 214.890 ;
        RECT 22.440 214.690 78.420 214.830 ;
        RECT 22.440 214.630 22.760 214.690 ;
        RECT 78.100 214.630 78.420 214.690 ;
        RECT 24.280 214.490 24.600 214.550 ;
        RECT 30.260 214.490 30.580 214.550 ;
        RECT 79.480 214.490 79.800 214.550 ;
        RECT 24.280 214.350 79.800 214.490 ;
        RECT 24.280 214.290 24.600 214.350 ;
        RECT 30.260 214.290 30.580 214.350 ;
        RECT 79.480 214.290 79.800 214.350 ;
        RECT 22.900 214.150 23.220 214.210 ;
        RECT 52.340 214.150 52.660 214.210 ;
        RECT 22.900 214.010 52.660 214.150 ;
        RECT 22.900 213.950 23.220 214.010 ;
        RECT 52.340 213.950 52.660 214.010 ;
        RECT 17.380 213.810 17.700 213.870 ;
        RECT 29.800 213.810 30.120 213.870 ;
        RECT 17.380 213.670 30.120 213.810 ;
        RECT 17.380 213.610 17.700 213.670 ;
        RECT 29.800 213.610 30.120 213.670 ;
        RECT 34.400 213.810 34.720 213.870 ;
        RECT 56.940 213.810 57.260 213.870 ;
        RECT 34.400 213.670 57.260 213.810 ;
        RECT 34.400 213.610 34.720 213.670 ;
        RECT 56.940 213.610 57.260 213.670 ;
        RECT 14.620 213.130 14.940 213.190 ;
        RECT 20.140 213.130 20.460 213.190 ;
        RECT 14.620 212.990 20.460 213.130 ;
        RECT 14.620 212.930 14.940 212.990 ;
        RECT 20.140 212.930 20.460 212.990 ;
        RECT 33.020 213.130 33.340 213.190 ;
        RECT 39.920 213.130 40.240 213.190 ;
        RECT 33.020 212.990 40.240 213.130 ;
        RECT 33.020 212.930 33.340 212.990 ;
        RECT 39.920 212.930 40.240 212.990 ;
        RECT 57.400 213.130 57.720 213.190 ;
        RECT 80.400 213.130 80.720 213.190 ;
        RECT 57.400 212.990 80.720 213.130 ;
        RECT 57.400 212.930 57.720 212.990 ;
        RECT 80.400 212.930 80.720 212.990 ;
        RECT 27.500 212.790 27.820 212.850 ;
        RECT 59.240 212.790 59.560 212.850 ;
        RECT 27.500 212.650 59.560 212.790 ;
        RECT 27.500 212.590 27.820 212.650 ;
        RECT 59.240 212.590 59.560 212.650 ;
        RECT 28.880 212.450 29.200 212.510 ;
        RECT 69.360 212.450 69.680 212.510 ;
        RECT 28.880 212.310 69.680 212.450 ;
        RECT 28.880 212.250 29.200 212.310 ;
        RECT 69.360 212.250 69.680 212.310 ;
        RECT 21.980 212.110 22.300 212.170 ;
        RECT 39.460 212.110 39.780 212.170 ;
        RECT 21.980 211.970 39.780 212.110 ;
        RECT 21.980 211.910 22.300 211.970 ;
        RECT 39.460 211.910 39.780 211.970 ;
        RECT 15.930 211.290 87.230 211.770 ;
        RECT 19.680 210.890 20.000 211.150 ;
        RECT 22.900 210.890 23.220 211.150 ;
        RECT 27.040 211.090 27.360 211.150 ;
        RECT 60.620 211.090 60.940 211.150 ;
        RECT 65.220 211.090 65.540 211.150 ;
        RECT 23.910 210.950 27.360 211.090 ;
        RECT 17.855 210.750 18.145 210.795 ;
        RECT 23.910 210.750 24.050 210.950 ;
        RECT 27.040 210.890 27.360 210.950 ;
        RECT 30.350 210.950 65.540 211.090 ;
        RECT 17.855 210.610 18.990 210.750 ;
        RECT 17.855 210.565 18.145 210.610 ;
        RECT 18.850 210.470 18.990 210.610 ;
        RECT 22.070 210.610 24.050 210.750 ;
        RECT 18.315 210.225 18.605 210.455 ;
        RECT 18.390 210.070 18.530 210.225 ;
        RECT 18.760 210.210 19.080 210.470 ;
        RECT 22.070 210.455 22.210 210.610 ;
        RECT 24.280 210.550 24.600 210.810 ;
        RECT 21.995 210.225 22.285 210.455 ;
        RECT 23.820 210.210 24.140 210.470 ;
        RECT 25.200 210.210 25.520 210.470 ;
        RECT 27.500 210.210 27.820 210.470 ;
        RECT 28.420 210.210 28.740 210.470 ;
        RECT 30.350 210.455 30.490 210.950 ;
        RECT 60.620 210.890 60.940 210.950 ;
        RECT 65.220 210.890 65.540 210.950 ;
        RECT 65.770 210.950 72.580 211.090 ;
        RECT 34.860 210.750 35.180 210.810 ;
        RECT 43.155 210.750 43.445 210.795 ;
        RECT 31.270 210.610 43.445 210.750 ;
        RECT 31.270 210.455 31.410 210.610 ;
        RECT 34.860 210.550 35.180 210.610 ;
        RECT 43.155 210.565 43.445 210.610 ;
        RECT 51.895 210.750 52.185 210.795 ;
        RECT 54.640 210.750 54.960 210.810 ;
        RECT 51.895 210.610 54.960 210.750 ;
        RECT 51.895 210.565 52.185 210.610 ;
        RECT 54.640 210.550 54.960 210.610 ;
        RECT 63.840 210.750 64.160 210.810 ;
        RECT 65.770 210.750 65.910 210.950 ;
        RECT 63.840 210.610 65.910 210.750 ;
        RECT 69.360 210.750 69.680 210.810 ;
        RECT 71.200 210.750 71.520 210.810 ;
        RECT 69.360 210.610 71.520 210.750 ;
        RECT 72.440 210.750 72.580 210.950 ;
        RECT 79.480 210.890 79.800 211.150 ;
        RECT 72.440 210.610 82.930 210.750 ;
        RECT 63.840 210.550 64.160 210.610 ;
        RECT 69.360 210.550 69.680 210.610 ;
        RECT 71.200 210.550 71.520 210.610 ;
        RECT 30.275 210.225 30.565 210.455 ;
        RECT 31.195 210.225 31.485 210.455 ;
        RECT 32.575 210.225 32.865 210.455 ;
        RECT 34.400 210.410 34.720 210.470 ;
        RECT 35.335 210.410 35.625 210.455 ;
        RECT 34.400 210.270 35.625 210.410 ;
        RECT 28.880 210.070 29.200 210.130 ;
        RECT 18.390 209.930 29.200 210.070 ;
        RECT 28.880 209.870 29.200 209.930 ;
        RECT 29.800 210.070 30.120 210.130 ;
        RECT 29.800 209.930 31.410 210.070 ;
        RECT 29.800 209.870 30.120 209.930 ;
        RECT 21.075 209.730 21.365 209.775 ;
        RECT 29.340 209.730 29.660 209.790 ;
        RECT 21.075 209.590 29.660 209.730 ;
        RECT 21.075 209.545 21.365 209.590 ;
        RECT 29.340 209.530 29.660 209.590 ;
        RECT 30.720 209.530 31.040 209.790 ;
        RECT 31.270 209.730 31.410 209.930 ;
        RECT 31.640 209.870 31.960 210.130 ;
        RECT 32.650 209.730 32.790 210.225 ;
        RECT 34.400 210.210 34.720 210.270 ;
        RECT 35.335 210.225 35.625 210.270 ;
        RECT 35.780 210.210 36.100 210.470 ;
        RECT 36.240 210.210 36.560 210.470 ;
        RECT 37.620 210.210 37.940 210.470 ;
        RECT 38.375 210.225 38.665 210.455 ;
        RECT 33.020 210.070 33.340 210.130 ;
        RECT 36.700 210.070 37.020 210.130 ;
        RECT 33.020 209.930 37.020 210.070 ;
        RECT 33.020 209.870 33.340 209.930 ;
        RECT 31.270 209.590 32.790 209.730 ;
        RECT 33.480 209.530 33.800 209.790 ;
        RECT 34.490 209.775 34.630 209.930 ;
        RECT 36.700 209.870 37.020 209.930 ;
        RECT 34.415 209.545 34.705 209.775 ;
        RECT 38.450 209.730 38.590 210.225 ;
        RECT 39.460 210.210 39.780 210.470 ;
        RECT 40.380 210.210 40.700 210.470 ;
        RECT 52.355 210.410 52.645 210.455 ;
        RECT 52.800 210.410 53.120 210.470 ;
        RECT 52.355 210.270 53.120 210.410 ;
        RECT 52.355 210.225 52.645 210.270 ;
        RECT 52.800 210.210 53.120 210.270 ;
        RECT 53.275 210.410 53.565 210.455 ;
        RECT 58.780 210.410 59.100 210.470 ;
        RECT 53.275 210.270 59.100 210.410 ;
        RECT 53.275 210.225 53.565 210.270 ;
        RECT 58.780 210.210 59.100 210.270 ;
        RECT 67.060 210.210 67.380 210.470 ;
        RECT 67.520 210.410 67.840 210.470 ;
        RECT 67.995 210.410 68.285 210.455 ;
        RECT 67.520 210.270 68.285 210.410 ;
        RECT 67.520 210.210 67.840 210.270 ;
        RECT 67.995 210.225 68.285 210.270 ;
        RECT 68.440 210.210 68.760 210.470 ;
        RECT 69.835 210.410 70.125 210.455 ;
        RECT 73.040 210.410 73.360 210.470 ;
        RECT 69.835 210.270 73.360 210.410 ;
        RECT 69.835 210.225 70.125 210.270 ;
        RECT 73.040 210.210 73.360 210.270 ;
        RECT 79.020 210.210 79.340 210.470 ;
        RECT 82.790 210.455 82.930 210.610 ;
        RECT 82.715 210.225 83.005 210.455 ;
        RECT 85.460 210.210 85.780 210.470 ;
        RECT 39.000 209.870 39.320 210.130 ;
        RECT 55.560 209.870 55.880 210.130 ;
        RECT 56.020 209.870 56.340 210.130 ;
        RECT 56.480 209.870 56.800 210.130 ;
        RECT 56.955 209.885 57.245 210.115 ;
        RECT 57.875 210.070 58.165 210.115 ;
        RECT 57.875 209.930 78.330 210.070 ;
        RECT 57.875 209.885 58.165 209.930 ;
        RECT 34.950 209.590 38.590 209.730 ;
        RECT 41.315 209.730 41.605 209.775 ;
        RECT 47.740 209.730 48.060 209.790 ;
        RECT 57.030 209.730 57.170 209.885 ;
        RECT 41.315 209.590 48.060 209.730 ;
        RECT 26.120 209.190 26.440 209.450 ;
        RECT 27.960 209.190 28.280 209.450 ;
        RECT 28.420 209.390 28.740 209.450 ;
        RECT 34.950 209.390 35.090 209.590 ;
        RECT 41.315 209.545 41.605 209.590 ;
        RECT 47.740 209.530 48.060 209.590 ;
        RECT 48.290 209.590 57.170 209.730 ;
        RECT 60.635 209.730 60.925 209.775 ;
        RECT 73.040 209.730 73.360 209.790 ;
        RECT 60.635 209.590 73.360 209.730 ;
        RECT 28.420 209.250 35.090 209.390 ;
        RECT 28.420 209.190 28.740 209.250 ;
        RECT 37.160 209.190 37.480 209.450 ;
        RECT 38.540 209.390 38.860 209.450 ;
        RECT 48.290 209.390 48.430 209.590 ;
        RECT 60.635 209.545 60.925 209.590 ;
        RECT 73.040 209.530 73.360 209.590 ;
        RECT 38.540 209.250 48.430 209.390 ;
        RECT 38.540 209.190 38.860 209.250 ;
        RECT 53.720 209.190 54.040 209.450 ;
        RECT 66.140 209.390 66.460 209.450 ;
        RECT 69.375 209.390 69.665 209.435 ;
        RECT 66.140 209.250 69.665 209.390 ;
        RECT 78.190 209.390 78.330 209.930 ;
        RECT 78.560 209.870 78.880 210.130 ;
        RECT 80.860 209.870 81.180 210.130 ;
        RECT 83.175 210.070 83.465 210.115 ;
        RECT 85.000 210.070 85.320 210.130 ;
        RECT 83.175 209.930 85.320 210.070 ;
        RECT 83.175 209.885 83.465 209.930 ;
        RECT 85.000 209.870 85.320 209.930 ;
        RECT 79.940 209.730 80.260 209.790 ;
        RECT 84.555 209.730 84.845 209.775 ;
        RECT 79.940 209.590 84.845 209.730 ;
        RECT 79.940 209.530 80.260 209.590 ;
        RECT 84.555 209.545 84.845 209.590 ;
        RECT 82.240 209.390 82.560 209.450 ;
        RECT 78.190 209.250 82.560 209.390 ;
        RECT 66.140 209.190 66.460 209.250 ;
        RECT 69.375 209.205 69.665 209.250 ;
        RECT 82.240 209.190 82.560 209.250 ;
        RECT 83.160 209.390 83.480 209.450 ;
        RECT 84.095 209.390 84.385 209.435 ;
        RECT 83.160 209.250 84.385 209.390 ;
        RECT 83.160 209.190 83.480 209.250 ;
        RECT 84.095 209.205 84.385 209.250 ;
        RECT 15.930 208.570 87.230 209.050 ;
        RECT 15.540 208.370 15.860 208.430 ;
        RECT 21.075 208.370 21.365 208.415 ;
        RECT 15.540 208.230 21.365 208.370 ;
        RECT 15.540 208.170 15.860 208.230 ;
        RECT 21.075 208.185 21.365 208.230 ;
        RECT 24.740 208.370 25.060 208.430 ;
        RECT 26.595 208.370 26.885 208.415 ;
        RECT 24.740 208.230 26.885 208.370 ;
        RECT 24.740 208.170 25.060 208.230 ;
        RECT 26.595 208.185 26.885 208.230 ;
        RECT 27.040 208.370 27.360 208.430 ;
        RECT 29.340 208.370 29.660 208.430 ;
        RECT 33.020 208.370 33.340 208.430 ;
        RECT 27.040 208.230 29.660 208.370 ;
        RECT 27.040 208.170 27.360 208.230 ;
        RECT 29.340 208.170 29.660 208.230 ;
        RECT 30.910 208.230 33.340 208.370 ;
        RECT 19.680 208.030 20.000 208.090 ;
        RECT 23.360 208.030 23.680 208.090 ;
        RECT 27.500 208.030 27.820 208.090 ;
        RECT 30.910 208.030 31.050 208.230 ;
        RECT 33.020 208.170 33.340 208.230 ;
        RECT 65.220 208.370 65.540 208.430 ;
        RECT 68.915 208.370 69.205 208.415 ;
        RECT 65.220 208.230 69.205 208.370 ;
        RECT 65.220 208.170 65.540 208.230 ;
        RECT 68.915 208.185 69.205 208.230 ;
        RECT 70.740 208.370 71.060 208.430 ;
        RECT 70.740 208.230 81.090 208.370 ;
        RECT 70.740 208.170 71.060 208.230 ;
        RECT 39.475 208.030 39.765 208.075 ;
        RECT 40.380 208.030 40.700 208.090 ;
        RECT 47.280 208.030 47.600 208.090 ;
        RECT 19.680 207.890 23.130 208.030 ;
        RECT 19.680 207.830 20.000 207.890 ;
        RECT 20.155 207.690 20.445 207.735 ;
        RECT 22.990 207.690 23.130 207.890 ;
        RECT 23.360 207.890 31.050 208.030 ;
        RECT 31.270 207.890 38.590 208.030 ;
        RECT 23.360 207.830 23.680 207.890 ;
        RECT 27.500 207.830 27.820 207.890 ;
        RECT 28.420 207.690 28.740 207.750 ;
        RECT 20.155 207.550 22.670 207.690 ;
        RECT 22.990 207.550 28.740 207.690 ;
        RECT 20.155 207.505 20.445 207.550 ;
        RECT 19.220 207.150 19.540 207.410 ;
        RECT 21.995 207.165 22.285 207.395 ;
        RECT 22.530 207.350 22.670 207.550 ;
        RECT 28.420 207.490 28.740 207.550 ;
        RECT 22.915 207.350 23.205 207.395 ;
        RECT 22.530 207.210 23.205 207.350 ;
        RECT 22.915 207.165 23.205 207.210 ;
        RECT 23.375 207.350 23.665 207.395 ;
        RECT 24.280 207.350 24.600 207.410 ;
        RECT 23.375 207.210 24.600 207.350 ;
        RECT 23.375 207.165 23.665 207.210 ;
        RECT 15.080 207.010 15.400 207.070 ;
        RECT 22.070 207.010 22.210 207.165 ;
        RECT 15.080 206.870 22.210 207.010 ;
        RECT 22.990 207.010 23.130 207.165 ;
        RECT 24.280 207.150 24.600 207.210 ;
        RECT 24.755 207.350 25.045 207.395 ;
        RECT 26.120 207.350 26.440 207.410 ;
        RECT 24.755 207.210 26.440 207.350 ;
        RECT 24.755 207.165 25.045 207.210 ;
        RECT 26.120 207.150 26.440 207.210 ;
        RECT 27.960 207.150 28.280 207.410 ;
        RECT 31.270 207.395 31.410 207.890 ;
        RECT 32.100 207.690 32.420 207.750 ;
        RECT 36.700 207.690 37.020 207.750 ;
        RECT 38.450 207.690 38.590 207.890 ;
        RECT 39.475 207.890 47.600 208.030 ;
        RECT 39.475 207.845 39.765 207.890 ;
        RECT 40.380 207.830 40.700 207.890 ;
        RECT 47.280 207.830 47.600 207.890 ;
        RECT 52.340 208.030 52.660 208.090 ;
        RECT 56.480 208.030 56.800 208.090 ;
        RECT 75.340 208.030 75.660 208.090 ;
        RECT 78.575 208.030 78.865 208.075 ;
        RECT 52.340 207.890 75.660 208.030 ;
        RECT 52.340 207.830 52.660 207.890 ;
        RECT 56.480 207.830 56.800 207.890 ;
        RECT 75.340 207.830 75.660 207.890 ;
        RECT 76.350 207.890 78.865 208.030 ;
        RECT 57.875 207.690 58.165 207.735 ;
        RECT 58.320 207.690 58.640 207.750 ;
        RECT 67.980 207.690 68.300 207.750 ;
        RECT 32.100 207.550 35.550 207.690 ;
        RECT 32.100 207.490 32.420 207.550 ;
        RECT 35.410 207.410 35.550 207.550 ;
        RECT 36.700 207.550 38.305 207.690 ;
        RECT 38.450 207.550 52.110 207.690 ;
        RECT 36.700 207.490 37.020 207.550 ;
        RECT 31.195 207.165 31.485 207.395 ;
        RECT 25.200 207.010 25.520 207.070 ;
        RECT 22.990 206.870 25.520 207.010 ;
        RECT 15.080 206.810 15.400 206.870 ;
        RECT 25.200 206.810 25.520 206.870 ;
        RECT 25.660 207.010 25.980 207.070 ;
        RECT 26.825 207.010 27.115 207.055 ;
        RECT 31.270 207.010 31.410 207.165 ;
        RECT 31.640 207.150 31.960 207.410 ;
        RECT 32.575 207.165 32.865 207.395 ;
        RECT 33.035 207.350 33.325 207.395 ;
        RECT 33.955 207.350 34.245 207.395 ;
        RECT 33.035 207.210 34.245 207.350 ;
        RECT 33.035 207.165 33.325 207.210 ;
        RECT 33.955 207.165 34.245 207.210 ;
        RECT 25.660 206.870 31.410 207.010 ;
        RECT 32.650 207.010 32.790 207.165 ;
        RECT 35.320 207.150 35.640 207.410 ;
        RECT 35.780 207.150 36.100 207.410 ;
        RECT 37.620 207.150 37.940 207.410 ;
        RECT 38.165 207.350 38.305 207.550 ;
        RECT 41.300 207.350 41.620 207.410 ;
        RECT 38.165 207.210 41.620 207.350 ;
        RECT 41.300 207.150 41.620 207.210 ;
        RECT 44.980 207.350 45.300 207.410 ;
        RECT 45.915 207.350 46.205 207.395 ;
        RECT 44.980 207.210 46.205 207.350 ;
        RECT 44.980 207.150 45.300 207.210 ;
        RECT 45.915 207.165 46.205 207.210 ;
        RECT 46.375 207.165 46.665 207.395 ;
        RECT 34.400 207.010 34.720 207.070 ;
        RECT 32.650 206.870 34.720 207.010 ;
        RECT 25.660 206.810 25.980 206.870 ;
        RECT 26.825 206.825 27.115 206.870 ;
        RECT 34.400 206.810 34.720 206.870 ;
        RECT 36.715 207.010 37.005 207.055 ;
        RECT 37.710 207.010 37.850 207.150 ;
        RECT 39.460 207.010 39.780 207.070 ;
        RECT 36.715 206.870 39.780 207.010 ;
        RECT 36.715 206.825 37.005 206.870 ;
        RECT 39.460 206.810 39.780 206.870 ;
        RECT 45.440 207.010 45.760 207.070 ;
        RECT 46.450 207.010 46.590 207.165 ;
        RECT 46.820 207.150 47.140 207.410 ;
        RECT 47.740 207.150 48.060 207.410 ;
        RECT 48.775 207.395 48.915 207.550 ;
        RECT 51.970 207.410 52.110 207.550 ;
        RECT 57.875 207.550 58.640 207.690 ;
        RECT 57.875 207.505 58.165 207.550 ;
        RECT 58.320 207.490 58.640 207.550 ;
        RECT 58.870 207.550 68.300 207.690 ;
        RECT 48.700 207.165 48.990 207.395 ;
        RECT 50.500 207.150 50.820 207.410 ;
        RECT 50.960 207.150 51.280 207.410 ;
        RECT 51.880 207.150 52.200 207.410 ;
        RECT 52.355 207.350 52.645 207.395 ;
        RECT 58.870 207.350 59.010 207.550 ;
        RECT 67.980 207.490 68.300 207.550 ;
        RECT 73.975 207.690 74.265 207.735 ;
        RECT 76.350 207.690 76.490 207.890 ;
        RECT 78.575 207.845 78.865 207.890 ;
        RECT 73.975 207.550 76.490 207.690 ;
        RECT 73.975 207.505 74.265 207.550 ;
        RECT 77.180 207.490 77.500 207.750 ;
        RECT 80.950 207.735 81.090 208.230 ;
        RECT 84.095 208.030 84.385 208.075 ;
        RECT 81.410 207.890 84.385 208.030 ;
        RECT 77.655 207.690 77.945 207.735 ;
        RECT 77.655 207.550 80.630 207.690 ;
        RECT 77.655 207.505 77.945 207.550 ;
        RECT 52.355 207.210 59.010 207.350 ;
        RECT 52.355 207.165 52.645 207.210 ;
        RECT 59.240 207.150 59.560 207.410 ;
        RECT 65.680 207.350 66.000 207.410 ;
        RECT 71.675 207.350 71.965 207.395 ;
        RECT 65.680 207.210 71.965 207.350 ;
        RECT 65.680 207.150 66.000 207.210 ;
        RECT 71.675 207.165 71.965 207.210 ;
        RECT 73.500 207.150 73.820 207.410 ;
        RECT 75.340 207.150 75.660 207.410 ;
        RECT 79.940 207.150 80.260 207.410 ;
        RECT 80.490 207.350 80.630 207.550 ;
        RECT 80.875 207.505 81.165 207.735 ;
        RECT 81.410 207.350 81.550 207.890 ;
        RECT 84.095 207.845 84.385 207.890 ;
        RECT 83.160 207.490 83.480 207.750 ;
        RECT 80.490 207.210 81.550 207.350 ;
        RECT 82.700 207.150 83.020 207.410 ;
        RECT 85.460 207.150 85.780 207.410 ;
        RECT 45.440 206.870 46.590 207.010 ;
        RECT 45.440 206.810 45.760 206.870 ;
        RECT 48.200 206.810 48.520 207.070 ;
        RECT 49.120 207.010 49.440 207.070 ;
        RECT 55.575 207.010 55.865 207.055 ;
        RECT 58.780 207.010 59.100 207.070 ;
        RECT 61.540 207.010 61.860 207.070 ;
        RECT 49.120 206.870 53.950 207.010 ;
        RECT 49.120 206.810 49.440 206.870 ;
        RECT 16.000 206.670 16.320 206.730 ;
        RECT 18.315 206.670 18.605 206.715 ;
        RECT 16.000 206.530 18.605 206.670 ;
        RECT 16.000 206.470 16.320 206.530 ;
        RECT 18.315 206.485 18.605 206.530 ;
        RECT 19.220 206.670 19.540 206.730 ;
        RECT 23.360 206.670 23.680 206.730 ;
        RECT 19.220 206.530 23.680 206.670 ;
        RECT 19.220 206.470 19.540 206.530 ;
        RECT 23.360 206.470 23.680 206.530 ;
        RECT 24.295 206.670 24.585 206.715 ;
        RECT 28.880 206.670 29.200 206.730 ;
        RECT 24.295 206.530 29.200 206.670 ;
        RECT 24.295 206.485 24.585 206.530 ;
        RECT 28.880 206.470 29.200 206.530 ;
        RECT 30.275 206.670 30.565 206.715 ;
        RECT 30.720 206.670 31.040 206.730 ;
        RECT 30.275 206.530 31.040 206.670 ;
        RECT 30.275 206.485 30.565 206.530 ;
        RECT 30.720 206.470 31.040 206.530 ;
        RECT 33.020 206.670 33.340 206.730 ;
        RECT 34.875 206.670 35.165 206.715 ;
        RECT 42.220 206.670 42.540 206.730 ;
        RECT 33.020 206.530 42.540 206.670 ;
        RECT 33.020 206.470 33.340 206.530 ;
        RECT 34.875 206.485 35.165 206.530 ;
        RECT 42.220 206.470 42.540 206.530 ;
        RECT 46.360 206.670 46.680 206.730 ;
        RECT 49.595 206.670 49.885 206.715 ;
        RECT 46.360 206.530 49.885 206.670 ;
        RECT 46.360 206.470 46.680 206.530 ;
        RECT 49.595 206.485 49.885 206.530 ;
        RECT 53.260 206.470 53.580 206.730 ;
        RECT 53.810 206.670 53.950 206.870 ;
        RECT 55.575 206.870 61.860 207.010 ;
        RECT 55.575 206.825 55.865 206.870 ;
        RECT 58.780 206.810 59.100 206.870 ;
        RECT 61.540 206.810 61.860 206.870 ;
        RECT 62.475 206.825 62.765 207.055 ;
        RECT 68.900 207.010 69.220 207.070 ;
        RECT 74.895 207.010 75.185 207.055 ;
        RECT 83.620 207.010 83.940 207.070 ;
        RECT 68.900 206.870 75.185 207.010 ;
        RECT 62.550 206.670 62.690 206.825 ;
        RECT 68.900 206.810 69.220 206.870 ;
        RECT 74.895 206.825 75.185 206.870 ;
        RECT 75.430 206.870 83.940 207.010 ;
        RECT 53.810 206.530 62.690 206.670 ;
        RECT 69.360 206.670 69.680 206.730 ;
        RECT 75.430 206.670 75.570 206.870 ;
        RECT 83.620 206.810 83.940 206.870 ;
        RECT 69.360 206.530 75.570 206.670 ;
        RECT 69.360 206.470 69.680 206.530 ;
        RECT 79.480 206.470 79.800 206.730 ;
        RECT 84.080 206.670 84.400 206.730 ;
        RECT 84.555 206.670 84.845 206.715 ;
        RECT 84.080 206.530 84.845 206.670 ;
        RECT 84.080 206.470 84.400 206.530 ;
        RECT 84.555 206.485 84.845 206.530 ;
        RECT 15.930 205.850 87.230 206.330 ;
        RECT 16.460 205.650 16.780 205.710 ;
        RECT 17.855 205.650 18.145 205.695 ;
        RECT 16.460 205.510 18.145 205.650 ;
        RECT 16.460 205.450 16.780 205.510 ;
        RECT 17.855 205.465 18.145 205.510 ;
        RECT 19.680 205.450 20.000 205.710 ;
        RECT 23.820 205.650 24.140 205.710 ;
        RECT 20.690 205.510 24.140 205.650 ;
        RECT 18.300 204.970 18.620 205.030 ;
        RECT 18.775 204.970 19.065 205.015 ;
        RECT 18.300 204.830 19.065 204.970 ;
        RECT 18.300 204.770 18.620 204.830 ;
        RECT 18.775 204.785 19.065 204.830 ;
        RECT 19.220 204.770 19.540 205.030 ;
        RECT 20.690 205.015 20.830 205.510 ;
        RECT 23.820 205.450 24.140 205.510 ;
        RECT 25.660 205.450 25.980 205.710 ;
        RECT 55.560 205.650 55.880 205.710 ;
        RECT 67.060 205.650 67.380 205.710 ;
        RECT 26.195 205.510 55.880 205.650 ;
        RECT 21.075 205.310 21.365 205.355 ;
        RECT 26.195 205.310 26.335 205.510 ;
        RECT 55.560 205.450 55.880 205.510 ;
        RECT 56.110 205.510 67.380 205.650 ;
        RECT 21.075 205.170 26.335 205.310 ;
        RECT 21.075 205.125 21.365 205.170 ;
        RECT 26.595 205.125 26.885 205.355 ;
        RECT 28.420 205.310 28.740 205.370 ;
        RECT 32.100 205.310 32.420 205.370 ;
        RECT 28.420 205.170 32.420 205.310 ;
        RECT 20.155 204.785 20.445 205.015 ;
        RECT 20.615 204.785 20.905 205.015 ;
        RECT 20.230 204.630 20.370 204.785 ;
        RECT 21.520 204.770 21.840 205.030 ;
        RECT 21.980 204.770 22.300 205.030 ;
        RECT 23.370 204.785 23.660 205.015 ;
        RECT 23.835 204.970 24.125 205.015 ;
        RECT 24.280 204.970 24.600 205.030 ;
        RECT 25.660 204.970 25.980 205.030 ;
        RECT 23.835 204.830 24.600 204.970 ;
        RECT 23.835 204.785 24.125 204.830 ;
        RECT 23.445 204.630 23.585 204.785 ;
        RECT 24.280 204.770 24.600 204.830 ;
        RECT 24.830 204.830 25.980 204.970 ;
        RECT 24.830 204.630 24.970 204.830 ;
        RECT 25.660 204.770 25.980 204.830 ;
        RECT 26.120 204.970 26.440 205.030 ;
        RECT 26.670 204.970 26.810 205.125 ;
        RECT 28.420 205.110 28.740 205.170 ;
        RECT 32.100 205.110 32.420 205.170 ;
        RECT 32.560 205.310 32.880 205.370 ;
        RECT 43.155 205.310 43.445 205.355 ;
        RECT 32.560 205.170 43.445 205.310 ;
        RECT 32.560 205.110 32.880 205.170 ;
        RECT 43.155 205.125 43.445 205.170 ;
        RECT 44.980 205.310 45.300 205.370 ;
        RECT 51.420 205.310 51.740 205.370 ;
        RECT 44.980 205.170 51.740 205.310 ;
        RECT 44.980 205.110 45.300 205.170 ;
        RECT 51.420 205.110 51.740 205.170 ;
        RECT 26.120 204.830 26.810 204.970 ;
        RECT 26.120 204.770 26.440 204.830 ;
        RECT 27.975 204.785 28.265 205.015 ;
        RECT 28.880 204.970 29.200 205.030 ;
        RECT 31.180 204.970 31.500 205.030 ;
        RECT 28.880 204.830 31.500 204.970 ;
        RECT 20.230 204.490 24.970 204.630 ;
        RECT 25.200 204.630 25.520 204.690 ;
        RECT 27.055 204.630 27.345 204.675 ;
        RECT 25.200 204.490 27.345 204.630 ;
        RECT 28.050 204.630 28.190 204.785 ;
        RECT 28.880 204.770 29.200 204.830 ;
        RECT 31.180 204.770 31.500 204.830 ;
        RECT 31.655 204.970 31.945 205.015 ;
        RECT 34.860 204.970 35.180 205.030 ;
        RECT 31.655 204.830 35.180 204.970 ;
        RECT 31.655 204.785 31.945 204.830 ;
        RECT 34.860 204.770 35.180 204.830 ;
        RECT 41.315 204.970 41.605 205.015 ;
        RECT 49.120 204.970 49.440 205.030 ;
        RECT 41.315 204.830 49.440 204.970 ;
        RECT 41.315 204.785 41.605 204.830 ;
        RECT 49.120 204.770 49.440 204.830 ;
        RECT 49.580 204.970 49.900 205.030 ;
        RECT 56.110 204.970 56.250 205.510 ;
        RECT 67.060 205.450 67.380 205.510 ;
        RECT 67.980 205.450 68.300 205.710 ;
        RECT 69.360 205.650 69.680 205.710 ;
        RECT 83.635 205.650 83.925 205.695 ;
        RECT 68.530 205.510 69.680 205.650 ;
        RECT 56.480 205.310 56.800 205.370 ;
        RECT 65.220 205.310 65.540 205.370 ;
        RECT 68.530 205.310 68.670 205.510 ;
        RECT 69.360 205.450 69.680 205.510 ;
        RECT 79.110 205.510 83.925 205.650 ;
        RECT 79.110 205.310 79.250 205.510 ;
        RECT 83.635 205.465 83.925 205.510 ;
        RECT 84.080 205.650 84.400 205.710 ;
        RECT 84.555 205.650 84.845 205.695 ;
        RECT 84.080 205.510 84.845 205.650 ;
        RECT 84.080 205.450 84.400 205.510 ;
        RECT 84.555 205.465 84.845 205.510 ;
        RECT 56.480 205.170 65.540 205.310 ;
        RECT 56.480 205.110 56.800 205.170 ;
        RECT 65.220 205.110 65.540 205.170 ;
        RECT 66.230 205.170 68.670 205.310 ;
        RECT 69.450 205.170 79.250 205.310 ;
        RECT 83.085 205.310 83.375 205.355 ;
        RECT 83.085 205.170 85.690 205.310 ;
        RECT 49.580 204.830 56.250 204.970 ;
        RECT 58.780 204.970 59.100 205.030 ;
        RECT 61.095 204.970 61.385 205.015 ;
        RECT 58.780 204.830 61.385 204.970 ;
        RECT 49.580 204.770 49.900 204.830 ;
        RECT 58.780 204.770 59.100 204.830 ;
        RECT 61.095 204.785 61.385 204.830 ;
        RECT 61.555 204.785 61.845 205.015 ;
        RECT 62.475 204.785 62.765 205.015 ;
        RECT 29.800 204.630 30.120 204.690 ;
        RECT 33.940 204.630 34.260 204.690 ;
        RECT 28.050 204.490 34.260 204.630 ;
        RECT 25.200 204.430 25.520 204.490 ;
        RECT 27.055 204.445 27.345 204.490 ;
        RECT 27.130 204.290 27.270 204.445 ;
        RECT 29.800 204.430 30.120 204.490 ;
        RECT 33.940 204.430 34.260 204.490 ;
        RECT 35.320 204.630 35.640 204.690 ;
        RECT 40.380 204.630 40.700 204.690 ;
        RECT 35.320 204.490 40.700 204.630 ;
        RECT 35.320 204.430 35.640 204.490 ;
        RECT 40.380 204.430 40.700 204.490 ;
        RECT 51.420 204.630 51.740 204.690 ;
        RECT 58.320 204.630 58.640 204.690 ;
        RECT 51.420 204.490 58.640 204.630 ;
        RECT 51.420 204.430 51.740 204.490 ;
        RECT 58.320 204.430 58.640 204.490 ;
        RECT 59.240 204.630 59.560 204.690 ;
        RECT 61.630 204.630 61.770 204.785 ;
        RECT 59.240 204.490 61.770 204.630 ;
        RECT 59.240 204.430 59.560 204.490 ;
        RECT 62.000 204.430 62.320 204.690 ;
        RECT 62.550 204.630 62.690 204.785 ;
        RECT 62.920 204.770 63.240 205.030 ;
        RECT 64.315 204.970 64.605 205.015 ;
        RECT 65.680 204.970 66.000 205.030 ;
        RECT 66.230 205.015 66.370 205.170 ;
        RECT 64.315 204.830 66.000 204.970 ;
        RECT 64.315 204.785 64.605 204.830 ;
        RECT 65.680 204.770 66.000 204.830 ;
        RECT 66.155 204.785 66.445 205.015 ;
        RECT 69.450 204.690 69.590 205.170 ;
        RECT 83.085 205.125 83.375 205.170 ;
        RECT 71.660 204.770 71.980 205.030 ;
        RECT 72.120 204.970 72.440 205.030 ;
        RECT 72.120 204.770 72.580 204.970 ;
        RECT 81.780 204.770 82.100 205.030 ;
        RECT 82.255 204.785 82.545 205.015 ;
        RECT 83.620 204.970 83.940 205.030 ;
        RECT 84.095 204.970 84.385 205.015 ;
        RECT 83.620 204.830 84.385 204.970 ;
        RECT 63.380 204.630 63.700 204.690 ;
        RECT 62.550 204.490 63.700 204.630 ;
        RECT 63.380 204.430 63.700 204.490 ;
        RECT 64.760 204.430 65.080 204.690 ;
        RECT 67.060 204.630 67.380 204.690 ;
        RECT 68.440 204.630 68.760 204.690 ;
        RECT 67.060 204.490 68.760 204.630 ;
        RECT 67.060 204.430 67.380 204.490 ;
        RECT 68.440 204.430 68.760 204.490 ;
        RECT 68.900 204.430 69.220 204.690 ;
        RECT 69.360 204.430 69.680 204.690 ;
        RECT 71.215 204.630 71.505 204.675 ;
        RECT 72.440 204.630 72.580 204.770 ;
        RECT 78.560 204.630 78.880 204.690 ;
        RECT 82.330 204.630 82.470 204.785 ;
        RECT 83.620 204.770 83.940 204.830 ;
        RECT 84.095 204.785 84.385 204.830 ;
        RECT 71.215 204.490 78.330 204.630 ;
        RECT 71.215 204.445 71.505 204.490 ;
        RECT 27.960 204.290 28.280 204.350 ;
        RECT 27.130 204.150 28.280 204.290 ;
        RECT 27.960 204.090 28.280 204.150 ;
        RECT 31.180 204.290 31.500 204.350 ;
        RECT 36.700 204.290 37.020 204.350 ;
        RECT 31.180 204.150 37.020 204.290 ;
        RECT 31.180 204.090 31.500 204.150 ;
        RECT 36.700 204.090 37.020 204.150 ;
        RECT 37.160 204.290 37.480 204.350 ;
        RECT 59.700 204.290 60.020 204.350 ;
        RECT 72.135 204.290 72.425 204.335 ;
        RECT 37.160 204.150 58.780 204.290 ;
        RECT 37.160 204.090 37.480 204.150 ;
        RECT 23.820 203.950 24.140 204.010 ;
        RECT 24.755 203.950 25.045 203.995 ;
        RECT 23.820 203.810 25.045 203.950 ;
        RECT 23.820 203.750 24.140 203.810 ;
        RECT 24.755 203.765 25.045 203.810 ;
        RECT 25.675 203.950 25.965 203.995 ;
        RECT 26.120 203.950 26.440 204.010 ;
        RECT 25.675 203.810 26.440 203.950 ;
        RECT 25.675 203.765 25.965 203.810 ;
        RECT 26.120 203.750 26.440 203.810 ;
        RECT 27.500 203.950 27.820 204.010 ;
        RECT 28.420 203.950 28.740 204.010 ;
        RECT 27.500 203.810 28.740 203.950 ;
        RECT 27.500 203.750 27.820 203.810 ;
        RECT 28.420 203.750 28.740 203.810 ;
        RECT 28.880 203.750 29.200 204.010 ;
        RECT 34.860 203.950 35.180 204.010 ;
        RECT 39.000 203.950 39.320 204.010 ;
        RECT 48.200 203.950 48.520 204.010 ;
        RECT 34.860 203.810 48.520 203.950 ;
        RECT 34.860 203.750 35.180 203.810 ;
        RECT 39.000 203.750 39.320 203.810 ;
        RECT 48.200 203.750 48.520 203.810 ;
        RECT 54.640 203.750 54.960 204.010 ;
        RECT 58.640 203.950 58.780 204.150 ;
        RECT 59.700 204.150 72.425 204.290 ;
        RECT 78.190 204.290 78.330 204.490 ;
        RECT 78.560 204.490 82.470 204.630 ;
        RECT 78.560 204.430 78.880 204.490 ;
        RECT 85.550 204.290 85.690 205.170 ;
        RECT 78.190 204.150 85.690 204.290 ;
        RECT 59.700 204.090 60.020 204.150 ;
        RECT 72.135 204.105 72.425 204.150 ;
        RECT 64.300 203.950 64.620 204.010 ;
        RECT 71.660 203.950 71.980 204.010 ;
        RECT 58.640 203.810 71.980 203.950 ;
        RECT 64.300 203.750 64.620 203.810 ;
        RECT 71.660 203.750 71.980 203.810 ;
        RECT 74.420 203.750 74.740 204.010 ;
        RECT 15.930 203.130 87.230 203.610 ;
        RECT 22.440 202.930 22.760 202.990 ;
        RECT 23.375 202.930 23.665 202.975 ;
        RECT 35.320 202.930 35.640 202.990 ;
        RECT 22.440 202.790 23.665 202.930 ;
        RECT 22.440 202.730 22.760 202.790 ;
        RECT 23.375 202.745 23.665 202.790 ;
        RECT 28.510 202.790 35.640 202.930 ;
        RECT 15.540 202.590 15.860 202.650 ;
        RECT 20.615 202.590 20.905 202.635 ;
        RECT 15.540 202.450 20.905 202.590 ;
        RECT 15.540 202.390 15.860 202.450 ;
        RECT 20.615 202.405 20.905 202.450 ;
        RECT 24.295 202.250 24.585 202.295 ;
        RECT 27.500 202.250 27.820 202.310 ;
        RECT 28.510 202.250 28.650 202.790 ;
        RECT 35.320 202.730 35.640 202.790 ;
        RECT 35.780 202.930 36.100 202.990 ;
        RECT 37.620 202.930 37.940 202.990 ;
        RECT 35.780 202.790 37.940 202.930 ;
        RECT 35.780 202.730 36.100 202.790 ;
        RECT 37.620 202.730 37.940 202.790 ;
        RECT 38.555 202.930 38.845 202.975 ;
        RECT 73.960 202.930 74.280 202.990 ;
        RECT 38.555 202.790 74.280 202.930 ;
        RECT 38.555 202.745 38.845 202.790 ;
        RECT 73.960 202.730 74.280 202.790 ;
        RECT 29.340 202.390 29.660 202.650 ;
        RECT 31.180 202.590 31.500 202.650 ;
        RECT 44.520 202.590 44.840 202.650 ;
        RECT 31.180 202.450 44.840 202.590 ;
        RECT 31.180 202.390 31.500 202.450 ;
        RECT 44.520 202.390 44.840 202.450 ;
        RECT 47.755 202.590 48.045 202.635 ;
        RECT 49.120 202.590 49.440 202.650 ;
        RECT 47.755 202.450 49.440 202.590 ;
        RECT 47.755 202.405 48.045 202.450 ;
        RECT 49.120 202.390 49.440 202.450 ;
        RECT 56.480 202.390 56.800 202.650 ;
        RECT 56.940 202.590 57.260 202.650 ;
        RECT 76.275 202.590 76.565 202.635 ;
        RECT 56.940 202.450 76.565 202.590 ;
        RECT 56.940 202.390 57.260 202.450 ;
        RECT 76.275 202.405 76.565 202.450 ;
        RECT 77.640 202.590 77.960 202.650 ;
        RECT 85.015 202.590 85.305 202.635 ;
        RECT 77.640 202.450 85.305 202.590 ;
        RECT 77.640 202.390 77.960 202.450 ;
        RECT 85.015 202.405 85.305 202.450 ;
        RECT 19.770 202.110 24.585 202.250 ;
        RECT 19.770 201.970 19.910 202.110 ;
        RECT 24.295 202.065 24.585 202.110 ;
        RECT 25.290 202.110 27.820 202.250 ;
        RECT 18.315 201.910 18.605 201.955 ;
        RECT 19.680 201.910 20.000 201.970 ;
        RECT 18.315 201.770 20.000 201.910 ;
        RECT 18.315 201.725 18.605 201.770 ;
        RECT 19.680 201.710 20.000 201.770 ;
        RECT 21.520 201.710 21.840 201.970 ;
        RECT 22.900 201.710 23.220 201.970 ;
        RECT 23.360 201.910 23.680 201.970 ;
        RECT 25.290 201.955 25.430 202.110 ;
        RECT 27.500 202.050 27.820 202.110 ;
        RECT 28.050 202.110 28.650 202.250 ;
        RECT 29.800 202.250 30.120 202.310 ;
        RECT 43.140 202.250 43.460 202.310 ;
        RECT 56.570 202.250 56.710 202.390 ;
        RECT 29.800 202.110 43.460 202.250 ;
        RECT 28.050 201.955 28.190 202.110 ;
        RECT 29.800 202.050 30.120 202.110 ;
        RECT 43.140 202.050 43.460 202.110 ;
        RECT 55.650 202.110 56.710 202.250 ;
        RECT 58.335 202.250 58.625 202.295 ;
        RECT 70.740 202.250 71.060 202.310 ;
        RECT 58.335 202.110 71.060 202.250 ;
        RECT 23.835 201.910 24.125 201.955 ;
        RECT 23.360 201.770 24.125 201.910 ;
        RECT 23.360 201.710 23.680 201.770 ;
        RECT 23.835 201.725 24.125 201.770 ;
        RECT 25.215 201.725 25.505 201.955 ;
        RECT 26.595 201.910 26.885 201.955 ;
        RECT 25.750 201.770 26.885 201.910 ;
        RECT 24.280 201.570 24.600 201.630 ;
        RECT 25.750 201.570 25.890 201.770 ;
        RECT 26.595 201.725 26.885 201.770 ;
        RECT 27.975 201.725 28.265 201.955 ;
        RECT 28.435 201.910 28.725 201.955 ;
        RECT 28.435 201.770 30.030 201.910 ;
        RECT 28.435 201.725 28.725 201.770 ;
        RECT 24.280 201.430 25.890 201.570 ;
        RECT 26.135 201.570 26.425 201.615 ;
        RECT 29.340 201.570 29.660 201.630 ;
        RECT 26.135 201.430 29.660 201.570 ;
        RECT 29.890 201.570 30.030 201.770 ;
        RECT 30.260 201.710 30.580 201.970 ;
        RECT 30.735 201.910 31.025 201.955 ;
        RECT 31.640 201.910 31.960 201.970 ;
        RECT 30.735 201.770 31.960 201.910 ;
        RECT 30.735 201.725 31.025 201.770 ;
        RECT 31.640 201.710 31.960 201.770 ;
        RECT 32.100 201.710 32.420 201.970 ;
        RECT 52.340 201.910 52.660 201.970 ;
        RECT 32.650 201.770 52.660 201.910 ;
        RECT 32.650 201.570 32.790 201.770 ;
        RECT 52.340 201.710 52.660 201.770 ;
        RECT 53.260 201.910 53.580 201.970 ;
        RECT 55.115 201.910 55.405 201.955 ;
        RECT 55.650 201.910 55.790 202.110 ;
        RECT 58.335 202.065 58.625 202.110 ;
        RECT 70.740 202.050 71.060 202.110 ;
        RECT 53.260 201.770 55.790 201.910 ;
        RECT 53.260 201.710 53.580 201.770 ;
        RECT 55.115 201.725 55.405 201.770 ;
        RECT 56.020 201.710 56.340 201.970 ;
        RECT 56.480 201.710 56.800 201.970 ;
        RECT 57.415 201.725 57.705 201.955 ;
        RECT 57.860 201.910 58.180 201.970 ;
        RECT 59.255 201.910 59.545 201.955 ;
        RECT 57.860 201.770 59.545 201.910 ;
        RECT 29.890 201.430 32.790 201.570 ;
        RECT 33.955 201.570 34.245 201.615 ;
        RECT 36.240 201.570 36.560 201.630 ;
        RECT 33.955 201.430 36.560 201.570 ;
        RECT 24.280 201.370 24.600 201.430 ;
        RECT 26.135 201.385 26.425 201.430 ;
        RECT 29.340 201.370 29.660 201.430 ;
        RECT 33.955 201.385 34.245 201.430 ;
        RECT 36.240 201.370 36.560 201.430 ;
        RECT 36.700 201.570 37.020 201.630 ;
        RECT 44.520 201.570 44.840 201.630 ;
        RECT 36.700 201.430 44.840 201.570 ;
        RECT 36.700 201.370 37.020 201.430 ;
        RECT 44.520 201.370 44.840 201.430 ;
        RECT 44.980 201.370 45.300 201.630 ;
        RECT 51.420 201.570 51.740 201.630 ;
        RECT 54.195 201.570 54.485 201.615 ;
        RECT 51.420 201.430 54.485 201.570 ;
        RECT 51.420 201.370 51.740 201.430 ;
        RECT 54.195 201.385 54.485 201.430 ;
        RECT 19.235 201.230 19.525 201.275 ;
        RECT 20.140 201.230 20.460 201.290 ;
        RECT 19.235 201.090 20.460 201.230 ;
        RECT 19.235 201.045 19.525 201.090 ;
        RECT 20.140 201.030 20.460 201.090 ;
        RECT 23.360 201.230 23.680 201.290 ;
        RECT 24.740 201.230 25.060 201.290 ;
        RECT 23.360 201.090 25.060 201.230 ;
        RECT 23.360 201.030 23.680 201.090 ;
        RECT 24.740 201.030 25.060 201.090 ;
        RECT 25.200 201.230 25.520 201.290 ;
        RECT 26.595 201.230 26.885 201.275 ;
        RECT 25.200 201.090 26.885 201.230 ;
        RECT 25.200 201.030 25.520 201.090 ;
        RECT 26.595 201.045 26.885 201.090 ;
        RECT 27.515 201.230 27.805 201.275 ;
        RECT 30.260 201.230 30.580 201.290 ;
        RECT 27.515 201.090 30.580 201.230 ;
        RECT 27.515 201.045 27.805 201.090 ;
        RECT 30.260 201.030 30.580 201.090 ;
        RECT 31.195 201.230 31.485 201.275 ;
        RECT 31.640 201.230 31.960 201.290 ;
        RECT 31.195 201.090 31.960 201.230 ;
        RECT 31.195 201.045 31.485 201.090 ;
        RECT 31.640 201.030 31.960 201.090 ;
        RECT 33.035 201.230 33.325 201.275 ;
        RECT 39.460 201.230 39.780 201.290 ;
        RECT 33.035 201.090 39.780 201.230 ;
        RECT 33.035 201.045 33.325 201.090 ;
        RECT 39.460 201.030 39.780 201.090 ;
        RECT 43.600 201.230 43.920 201.290 ;
        RECT 57.490 201.230 57.630 201.725 ;
        RECT 57.860 201.710 58.180 201.770 ;
        RECT 59.255 201.725 59.545 201.770 ;
        RECT 60.175 201.910 60.465 201.955 ;
        RECT 61.080 201.910 61.400 201.970 ;
        RECT 79.035 201.910 79.325 201.955 ;
        RECT 79.480 201.910 79.800 201.970 ;
        RECT 60.175 201.770 70.510 201.910 ;
        RECT 60.175 201.725 60.465 201.770 ;
        RECT 61.080 201.710 61.400 201.770 ;
        RECT 58.320 201.570 58.640 201.630 ;
        RECT 60.635 201.570 60.925 201.615 ;
        RECT 69.835 201.570 70.125 201.615 ;
        RECT 58.320 201.430 60.925 201.570 ;
        RECT 58.320 201.370 58.640 201.430 ;
        RECT 60.635 201.385 60.925 201.430 ;
        RECT 61.170 201.430 70.125 201.570 ;
        RECT 70.370 201.570 70.510 201.770 ;
        RECT 79.035 201.770 79.800 201.910 ;
        RECT 79.035 201.725 79.325 201.770 ;
        RECT 79.110 201.570 79.250 201.725 ;
        RECT 79.480 201.710 79.800 201.770 ;
        RECT 80.400 201.910 80.720 201.970 ;
        RECT 80.875 201.910 81.165 201.955 ;
        RECT 80.400 201.770 81.165 201.910 ;
        RECT 80.400 201.710 80.720 201.770 ;
        RECT 80.875 201.725 81.165 201.770 ;
        RECT 81.320 201.910 81.640 201.970 ;
        RECT 83.175 201.910 83.465 201.955 ;
        RECT 84.095 201.910 84.385 201.955 ;
        RECT 81.320 201.770 83.465 201.910 ;
        RECT 81.320 201.710 81.640 201.770 ;
        RECT 83.175 201.725 83.465 201.770 ;
        RECT 83.710 201.770 84.385 201.910 ;
        RECT 70.370 201.430 79.250 201.570 ;
        RECT 43.600 201.090 57.630 201.230 ;
        RECT 59.240 201.230 59.560 201.290 ;
        RECT 59.715 201.230 60.005 201.275 ;
        RECT 59.240 201.090 60.005 201.230 ;
        RECT 43.600 201.030 43.920 201.090 ;
        RECT 59.240 201.030 59.560 201.090 ;
        RECT 59.715 201.045 60.005 201.090 ;
        RECT 60.160 201.230 60.480 201.290 ;
        RECT 61.170 201.230 61.310 201.430 ;
        RECT 69.835 201.385 70.125 201.430 ;
        RECT 82.240 201.370 82.560 201.630 ;
        RECT 60.160 201.090 61.310 201.230 ;
        RECT 61.540 201.230 61.860 201.290 ;
        RECT 67.075 201.230 67.365 201.275 ;
        RECT 61.540 201.090 67.365 201.230 ;
        RECT 60.160 201.030 60.480 201.090 ;
        RECT 61.540 201.030 61.860 201.090 ;
        RECT 67.075 201.045 67.365 201.090 ;
        RECT 79.955 201.230 80.245 201.275 ;
        RECT 83.710 201.230 83.850 201.770 ;
        RECT 84.095 201.725 84.385 201.770 ;
        RECT 79.955 201.090 83.850 201.230 ;
        RECT 79.955 201.045 80.245 201.090 ;
        RECT 15.930 200.410 87.230 200.890 ;
        RECT 20.155 200.210 20.445 200.255 ;
        RECT 20.600 200.210 20.920 200.270 ;
        RECT 20.155 200.070 20.920 200.210 ;
        RECT 20.155 200.025 20.445 200.070 ;
        RECT 20.600 200.010 20.920 200.070 ;
        RECT 21.060 200.210 21.380 200.270 ;
        RECT 21.535 200.210 21.825 200.255 ;
        RECT 21.060 200.070 21.825 200.210 ;
        RECT 21.060 200.010 21.380 200.070 ;
        RECT 21.535 200.025 21.825 200.070 ;
        RECT 28.435 200.210 28.725 200.255 ;
        RECT 29.800 200.210 30.120 200.270 ;
        RECT 28.435 200.070 30.120 200.210 ;
        RECT 28.435 200.025 28.725 200.070 ;
        RECT 29.800 200.010 30.120 200.070 ;
        RECT 33.480 200.210 33.800 200.270 ;
        RECT 33.480 200.070 35.550 200.210 ;
        RECT 33.480 200.010 33.800 200.070 ;
        RECT 18.760 199.330 19.080 199.590 ;
        RECT 20.690 199.575 20.830 200.010 ;
        RECT 22.440 199.870 22.760 199.930 ;
        RECT 23.835 199.870 24.125 199.915 ;
        RECT 22.440 199.730 24.125 199.870 ;
        RECT 22.440 199.670 22.760 199.730 ;
        RECT 23.835 199.685 24.125 199.730 ;
        RECT 25.200 199.870 25.520 199.930 ;
        RECT 25.200 199.730 26.350 199.870 ;
        RECT 25.200 199.670 25.520 199.730 ;
        RECT 20.615 199.345 20.905 199.575 ;
        RECT 22.900 199.330 23.220 199.590 ;
        RECT 23.360 199.330 23.680 199.590 ;
        RECT 24.280 199.575 24.600 199.590 ;
        RECT 24.280 199.530 24.815 199.575 ;
        RECT 25.675 199.530 25.965 199.575 ;
        RECT 24.280 199.390 25.965 199.530 ;
        RECT 26.210 199.530 26.350 199.730 ;
        RECT 29.340 199.670 29.660 199.930 ;
        RECT 35.410 199.915 35.550 200.070 ;
        RECT 37.160 200.010 37.480 200.270 ;
        RECT 38.540 200.010 38.860 200.270 ;
        RECT 39.000 200.210 39.320 200.270 ;
        RECT 45.915 200.210 46.205 200.255 ;
        RECT 46.820 200.210 47.140 200.270 ;
        RECT 53.260 200.210 53.580 200.270 ;
        RECT 39.000 200.070 45.670 200.210 ;
        RECT 39.000 200.010 39.320 200.070 ;
        RECT 29.930 199.730 35.090 199.870 ;
        RECT 26.595 199.530 26.885 199.575 ;
        RECT 26.210 199.390 26.885 199.530 ;
        RECT 24.280 199.345 24.815 199.390 ;
        RECT 25.675 199.345 25.965 199.390 ;
        RECT 26.595 199.345 26.885 199.390 ;
        RECT 27.975 199.530 28.265 199.575 ;
        RECT 29.930 199.530 30.070 199.730 ;
        RECT 30.810 199.575 30.950 199.730 ;
        RECT 34.950 199.590 35.090 199.730 ;
        RECT 35.335 199.685 35.625 199.915 ;
        RECT 36.240 199.870 36.560 199.930 ;
        RECT 45.530 199.870 45.670 200.070 ;
        RECT 45.915 200.070 47.140 200.210 ;
        RECT 45.915 200.025 46.205 200.070 ;
        RECT 46.820 200.010 47.140 200.070 ;
        RECT 47.370 200.070 53.580 200.210 ;
        RECT 47.370 199.870 47.510 200.070 ;
        RECT 53.260 200.010 53.580 200.070 ;
        RECT 54.640 200.210 54.960 200.270 ;
        RECT 66.155 200.210 66.445 200.255 ;
        RECT 67.060 200.210 67.380 200.270 ;
        RECT 54.640 200.070 64.990 200.210 ;
        RECT 54.640 200.010 54.960 200.070 ;
        RECT 50.055 199.870 50.345 199.915 ;
        RECT 50.960 199.870 51.280 199.930 ;
        RECT 36.240 199.730 45.210 199.870 ;
        RECT 45.530 199.730 47.510 199.870 ;
        RECT 36.240 199.670 36.560 199.730 ;
        RECT 27.975 199.390 30.070 199.530 ;
        RECT 27.975 199.345 28.265 199.390 ;
        RECT 30.275 199.345 30.565 199.575 ;
        RECT 30.735 199.345 31.025 199.575 ;
        RECT 31.180 199.530 31.500 199.590 ;
        RECT 31.655 199.530 31.945 199.575 ;
        RECT 31.180 199.390 31.945 199.530 ;
        RECT 24.280 199.330 24.600 199.345 ;
        RECT 21.980 198.990 22.300 199.250 ;
        RECT 25.200 198.990 25.520 199.250 ;
        RECT 26.120 199.190 26.440 199.250 ;
        RECT 27.515 199.190 27.805 199.235 ;
        RECT 26.120 199.050 27.805 199.190 ;
        RECT 26.120 198.990 26.440 199.050 ;
        RECT 27.515 199.005 27.805 199.050 ;
        RECT 29.340 199.190 29.660 199.250 ;
        RECT 30.350 199.190 30.490 199.345 ;
        RECT 31.180 199.330 31.500 199.390 ;
        RECT 31.655 199.345 31.945 199.390 ;
        RECT 32.100 199.330 32.420 199.590 ;
        RECT 32.575 199.530 32.865 199.575 ;
        RECT 32.575 199.390 34.700 199.530 ;
        RECT 32.575 199.345 32.865 199.390 ;
        RECT 29.340 199.050 30.490 199.190 ;
        RECT 27.590 198.850 27.730 199.005 ;
        RECT 29.340 198.990 29.660 199.050 ;
        RECT 32.650 198.850 32.790 199.345 ;
        RECT 34.560 199.190 34.700 199.390 ;
        RECT 34.860 199.330 35.180 199.590 ;
        RECT 35.795 199.345 36.085 199.575 ;
        RECT 35.870 199.190 36.010 199.345 ;
        RECT 36.700 199.330 37.020 199.590 ;
        RECT 37.250 199.575 37.390 199.730 ;
        RECT 37.175 199.345 37.465 199.575 ;
        RECT 38.095 199.530 38.385 199.575 ;
        RECT 39.000 199.530 39.320 199.590 ;
        RECT 38.095 199.390 39.320 199.530 ;
        RECT 38.095 199.345 38.385 199.390 ;
        RECT 39.000 199.330 39.320 199.390 ;
        RECT 39.460 199.330 39.780 199.590 ;
        RECT 39.935 199.530 40.225 199.575 ;
        RECT 41.760 199.530 42.080 199.590 ;
        RECT 39.935 199.390 42.080 199.530 ;
        RECT 39.935 199.345 40.225 199.390 ;
        RECT 41.760 199.330 42.080 199.390 ;
        RECT 42.220 199.530 42.540 199.590 ;
        RECT 42.695 199.530 42.985 199.575 ;
        RECT 42.220 199.390 42.985 199.530 ;
        RECT 42.220 199.330 42.540 199.390 ;
        RECT 42.695 199.345 42.985 199.390 ;
        RECT 43.140 199.330 43.460 199.590 ;
        RECT 45.070 199.575 45.210 199.730 ;
        RECT 44.995 199.345 45.285 199.575 ;
        RECT 46.835 199.530 47.125 199.575 ;
        RECT 47.370 199.530 47.510 199.730 ;
        RECT 48.290 199.730 49.335 199.870 ;
        RECT 46.835 199.390 47.510 199.530 ;
        RECT 46.835 199.345 47.125 199.390 ;
        RECT 47.740 199.330 48.060 199.590 ;
        RECT 48.290 199.575 48.430 199.730 ;
        RECT 48.215 199.345 48.505 199.575 ;
        RECT 48.680 199.295 48.970 199.525 ;
        RECT 38.540 199.190 38.860 199.250 ;
        RECT 34.560 199.050 38.860 199.190 ;
        RECT 38.540 198.990 38.860 199.050 ;
        RECT 40.380 198.990 40.700 199.250 ;
        RECT 40.840 198.990 41.160 199.250 ;
        RECT 27.590 198.710 32.790 198.850 ;
        RECT 33.495 198.850 33.785 198.895 ;
        RECT 37.620 198.850 37.940 198.910 ;
        RECT 48.755 198.850 48.895 199.295 ;
        RECT 33.495 198.710 35.090 198.850 ;
        RECT 33.495 198.665 33.785 198.710 ;
        RECT 17.840 198.310 18.160 198.570 ;
        RECT 29.800 198.510 30.120 198.570 ;
        RECT 33.955 198.510 34.245 198.555 ;
        RECT 29.800 198.370 34.245 198.510 ;
        RECT 34.950 198.510 35.090 198.710 ;
        RECT 37.620 198.710 48.895 198.850 ;
        RECT 37.620 198.650 37.940 198.710 ;
        RECT 36.240 198.510 36.560 198.570 ;
        RECT 34.950 198.370 36.560 198.510 ;
        RECT 29.800 198.310 30.120 198.370 ;
        RECT 33.955 198.325 34.245 198.370 ;
        RECT 36.240 198.310 36.560 198.370 ;
        RECT 40.380 198.510 40.700 198.570 ;
        RECT 44.995 198.510 45.285 198.555 ;
        RECT 49.195 198.510 49.335 199.730 ;
        RECT 50.055 199.730 51.280 199.870 ;
        RECT 50.055 199.685 50.345 199.730 ;
        RECT 50.960 199.670 51.280 199.730 ;
        RECT 56.020 199.870 56.340 199.930 ;
        RECT 64.315 199.870 64.605 199.915 ;
        RECT 56.020 199.730 64.605 199.870 ;
        RECT 64.850 199.870 64.990 200.070 ;
        RECT 66.155 200.070 67.380 200.210 ;
        RECT 66.155 200.025 66.445 200.070 ;
        RECT 67.060 200.010 67.380 200.070 ;
        RECT 67.980 200.210 68.300 200.270 ;
        RECT 74.435 200.210 74.725 200.255 ;
        RECT 67.980 200.070 74.725 200.210 ;
        RECT 67.980 200.010 68.300 200.070 ;
        RECT 74.435 200.025 74.725 200.070 ;
        RECT 78.560 200.210 78.880 200.270 ;
        RECT 82.240 200.210 82.560 200.270 ;
        RECT 78.560 200.070 82.560 200.210 ;
        RECT 78.560 200.010 78.880 200.070 ;
        RECT 82.240 200.010 82.560 200.070 ;
        RECT 84.555 200.210 84.845 200.255 ;
        RECT 87.300 200.210 87.620 200.270 ;
        RECT 84.555 200.070 87.620 200.210 ;
        RECT 84.555 200.025 84.845 200.070 ;
        RECT 87.300 200.010 87.620 200.070 ;
        RECT 69.820 199.870 70.140 199.930 ;
        RECT 64.850 199.730 68.210 199.870 ;
        RECT 56.020 199.670 56.340 199.730 ;
        RECT 64.315 199.685 64.605 199.730 ;
        RECT 50.515 199.530 50.805 199.575 ;
        RECT 53.720 199.530 54.040 199.590 ;
        RECT 50.515 199.390 54.040 199.530 ;
        RECT 50.515 199.345 50.805 199.390 ;
        RECT 53.720 199.330 54.040 199.390 ;
        RECT 59.700 199.330 60.020 199.590 ;
        RECT 60.620 199.330 60.940 199.590 ;
        RECT 61.540 199.330 61.860 199.590 ;
        RECT 62.935 199.530 63.225 199.575 ;
        RECT 65.235 199.530 65.525 199.575 ;
        RECT 62.935 199.390 65.525 199.530 ;
        RECT 62.935 199.345 63.225 199.390 ;
        RECT 65.235 199.345 65.525 199.390 ;
        RECT 66.615 199.530 66.905 199.575 ;
        RECT 67.520 199.530 67.840 199.590 ;
        RECT 68.070 199.575 68.210 199.730 ;
        RECT 69.820 199.730 79.710 199.870 ;
        RECT 69.820 199.670 70.140 199.730 ;
        RECT 66.615 199.390 67.840 199.530 ;
        RECT 66.615 199.345 66.905 199.390 ;
        RECT 58.320 199.190 58.640 199.250 ;
        RECT 60.160 199.190 60.480 199.250 ;
        RECT 58.320 199.050 60.480 199.190 ;
        RECT 58.320 198.990 58.640 199.050 ;
        RECT 60.160 198.990 60.480 199.050 ;
        RECT 61.095 199.005 61.385 199.235 ;
        RECT 62.015 199.005 62.305 199.235 ;
        RECT 54.640 198.850 54.960 198.910 ;
        RECT 60.620 198.850 60.940 198.910 ;
        RECT 61.170 198.850 61.310 199.005 ;
        RECT 54.640 198.710 57.170 198.850 ;
        RECT 54.640 198.650 54.960 198.710 ;
        RECT 40.380 198.370 49.335 198.510 ;
        RECT 52.340 198.510 52.660 198.570 ;
        RECT 56.480 198.510 56.800 198.570 ;
        RECT 52.340 198.370 56.800 198.510 ;
        RECT 57.030 198.510 57.170 198.710 ;
        RECT 60.620 198.710 61.310 198.850 ;
        RECT 61.540 198.850 61.860 198.910 ;
        RECT 62.090 198.850 62.230 199.005 ;
        RECT 61.540 198.710 62.230 198.850 ;
        RECT 60.620 198.650 60.940 198.710 ;
        RECT 61.540 198.650 61.860 198.710 ;
        RECT 66.690 198.510 66.830 199.345 ;
        RECT 67.520 199.330 67.840 199.390 ;
        RECT 67.995 199.345 68.285 199.575 ;
        RECT 68.440 199.530 68.760 199.590 ;
        RECT 77.195 199.530 77.485 199.575 ;
        RECT 68.440 199.390 77.485 199.530 ;
        RECT 68.440 199.330 68.760 199.390 ;
        RECT 77.195 199.345 77.485 199.390 ;
        RECT 78.560 199.330 78.880 199.590 ;
        RECT 79.020 199.330 79.340 199.590 ;
        RECT 79.570 199.575 79.710 199.730 ;
        RECT 80.030 199.730 83.850 199.870 ;
        RECT 80.030 199.575 80.170 199.730 ;
        RECT 83.710 199.590 83.850 199.730 ;
        RECT 79.495 199.345 79.785 199.575 ;
        RECT 79.955 199.345 80.245 199.575 ;
        RECT 82.240 199.330 82.560 199.590 ;
        RECT 83.620 199.330 83.940 199.590 ;
        RECT 85.475 199.530 85.765 199.575 ;
        RECT 85.920 199.530 86.240 199.590 ;
        RECT 85.475 199.390 86.240 199.530 ;
        RECT 85.475 199.345 85.765 199.390 ;
        RECT 85.920 199.330 86.240 199.390 ;
        RECT 76.720 199.190 77.040 199.250 ;
        RECT 81.335 199.190 81.625 199.235 ;
        RECT 83.175 199.190 83.465 199.235 ;
        RECT 76.720 199.050 81.625 199.190 ;
        RECT 76.720 198.990 77.040 199.050 ;
        RECT 81.335 199.005 81.625 199.050 ;
        RECT 81.870 199.050 83.465 199.190 ;
        RECT 79.020 198.850 79.340 198.910 ;
        RECT 81.870 198.850 82.010 199.050 ;
        RECT 83.175 199.005 83.465 199.050 ;
        RECT 79.020 198.710 82.010 198.850 ;
        RECT 79.020 198.650 79.340 198.710 ;
        RECT 82.735 198.665 83.025 198.895 ;
        RECT 57.030 198.370 66.830 198.510 ;
        RECT 78.100 198.510 78.420 198.570 ;
        RECT 82.790 198.510 82.930 198.665 ;
        RECT 78.100 198.370 82.930 198.510 ;
        RECT 40.380 198.310 40.700 198.370 ;
        RECT 44.995 198.325 45.285 198.370 ;
        RECT 52.340 198.310 52.660 198.370 ;
        RECT 56.480 198.310 56.800 198.370 ;
        RECT 78.100 198.310 78.420 198.370 ;
        RECT 15.930 197.690 87.230 198.170 ;
        RECT 22.455 197.490 22.745 197.535 ;
        RECT 22.900 197.490 23.220 197.550 ;
        RECT 22.455 197.350 23.220 197.490 ;
        RECT 22.455 197.305 22.745 197.350 ;
        RECT 22.900 197.290 23.220 197.350 ;
        RECT 27.040 197.490 27.360 197.550 ;
        RECT 27.515 197.490 27.805 197.535 ;
        RECT 27.040 197.350 27.805 197.490 ;
        RECT 27.040 197.290 27.360 197.350 ;
        RECT 27.515 197.305 27.805 197.350 ;
        RECT 28.420 197.490 28.740 197.550 ;
        RECT 29.815 197.490 30.105 197.535 ;
        RECT 28.420 197.350 30.105 197.490 ;
        RECT 28.420 197.290 28.740 197.350 ;
        RECT 29.815 197.305 30.105 197.350 ;
        RECT 31.655 197.490 31.945 197.535 ;
        RECT 42.220 197.490 42.540 197.550 ;
        RECT 31.655 197.350 42.540 197.490 ;
        RECT 31.655 197.305 31.945 197.350 ;
        RECT 42.220 197.290 42.540 197.350 ;
        RECT 47.740 197.490 48.060 197.550 ;
        RECT 50.055 197.490 50.345 197.535 ;
        RECT 47.740 197.350 50.345 197.490 ;
        RECT 47.740 197.290 48.060 197.350 ;
        RECT 50.055 197.305 50.345 197.350 ;
        RECT 52.340 197.490 52.660 197.550 ;
        RECT 57.860 197.490 58.180 197.550 ;
        RECT 78.560 197.490 78.880 197.550 ;
        RECT 52.340 197.350 58.180 197.490 ;
        RECT 52.340 197.290 52.660 197.350 ;
        RECT 57.860 197.290 58.180 197.350 ;
        RECT 63.930 197.350 78.880 197.490 ;
        RECT 23.360 197.150 23.680 197.210 ;
        RECT 29.340 197.150 29.660 197.210 ;
        RECT 31.180 197.150 31.500 197.210 ;
        RECT 33.940 197.150 34.260 197.210 ;
        RECT 23.360 197.010 24.970 197.150 ;
        RECT 23.360 196.950 23.680 197.010 ;
        RECT 20.140 196.610 20.460 196.870 ;
        RECT 24.280 196.810 24.600 196.870 ;
        RECT 24.140 196.610 24.600 196.810 ;
        RECT 19.235 196.335 19.525 196.565 ;
        RECT 19.680 196.470 20.000 196.530 ;
        RECT 21.535 196.470 21.825 196.515 ;
        RECT 19.310 196.190 19.450 196.335 ;
        RECT 19.680 196.330 21.825 196.470 ;
        RECT 19.680 196.270 20.000 196.330 ;
        RECT 21.535 196.285 21.825 196.330 ;
        RECT 22.900 196.270 23.220 196.530 ;
        RECT 23.705 196.470 23.995 196.515 ;
        RECT 24.140 196.470 24.280 196.610 ;
        RECT 24.830 196.515 24.970 197.010 ;
        RECT 29.340 197.010 31.500 197.150 ;
        RECT 29.340 196.950 29.660 197.010 ;
        RECT 31.180 196.950 31.500 197.010 ;
        RECT 32.190 197.010 34.260 197.150 ;
        RECT 32.190 196.855 32.330 197.010 ;
        RECT 33.940 196.950 34.260 197.010 ;
        RECT 36.700 196.950 37.020 197.210 ;
        RECT 39.935 197.150 40.225 197.195 ;
        RECT 44.980 197.150 45.300 197.210 ;
        RECT 39.935 197.010 45.300 197.150 ;
        RECT 39.935 196.965 40.225 197.010 ;
        RECT 44.980 196.950 45.300 197.010 ;
        RECT 48.200 197.150 48.520 197.210 ;
        RECT 48.200 197.010 52.570 197.150 ;
        RECT 48.200 196.950 48.520 197.010 ;
        RECT 25.290 196.670 31.870 196.810 ;
        RECT 25.290 196.530 25.430 196.670 ;
        RECT 23.705 196.330 24.280 196.470 ;
        RECT 23.705 196.285 23.995 196.330 ;
        RECT 24.755 196.285 25.045 196.515 ;
        RECT 19.220 195.930 19.540 196.190 ;
        RECT 20.600 195.930 20.920 196.190 ;
        RECT 24.290 195.945 24.580 196.175 ;
        RECT 24.830 196.130 24.970 196.285 ;
        RECT 25.200 196.270 25.520 196.530 ;
        RECT 26.120 196.270 26.440 196.530 ;
        RECT 28.420 196.270 28.740 196.530 ;
        RECT 29.355 196.285 29.645 196.515 ;
        RECT 30.275 196.285 30.565 196.515 ;
        RECT 30.735 196.470 31.025 196.515 ;
        RECT 31.180 196.470 31.500 196.530 ;
        RECT 30.735 196.330 31.500 196.470 ;
        RECT 31.730 196.470 31.870 196.670 ;
        RECT 32.115 196.625 32.405 196.855 ;
        RECT 36.790 196.810 36.930 196.950 ;
        RECT 34.030 196.670 36.930 196.810 ;
        RECT 39.460 196.810 39.780 196.870 ;
        RECT 42.220 196.810 42.540 196.870 ;
        RECT 39.460 196.670 42.540 196.810 ;
        RECT 32.575 196.470 32.865 196.515 ;
        RECT 31.730 196.330 32.865 196.470 ;
        RECT 30.735 196.285 31.025 196.330 ;
        RECT 26.210 196.130 26.350 196.270 ;
        RECT 24.830 195.990 26.350 196.130 ;
        RECT 27.040 196.130 27.360 196.190 ;
        RECT 29.430 196.130 29.570 196.285 ;
        RECT 27.040 195.990 29.570 196.130 ;
        RECT 30.350 196.130 30.490 196.285 ;
        RECT 31.180 196.270 31.500 196.330 ;
        RECT 32.575 196.285 32.865 196.330 ;
        RECT 33.020 196.470 33.340 196.530 ;
        RECT 34.030 196.515 34.170 196.670 ;
        RECT 39.460 196.610 39.780 196.670 ;
        RECT 42.220 196.610 42.540 196.670 ;
        RECT 47.280 196.810 47.600 196.870 ;
        RECT 52.430 196.855 52.570 197.010 ;
        RECT 51.435 196.810 51.725 196.855 ;
        RECT 47.280 196.670 51.725 196.810 ;
        RECT 47.280 196.610 47.600 196.670 ;
        RECT 51.435 196.625 51.725 196.670 ;
        RECT 52.355 196.625 52.645 196.855 ;
        RECT 60.620 196.810 60.940 196.870 ;
        RECT 52.890 196.670 60.940 196.810 ;
        RECT 33.495 196.470 33.785 196.515 ;
        RECT 33.020 196.330 33.785 196.470 ;
        RECT 33.020 196.270 33.340 196.330 ;
        RECT 33.495 196.285 33.785 196.330 ;
        RECT 33.955 196.285 34.245 196.515 ;
        RECT 34.400 196.270 34.720 196.530 ;
        RECT 35.335 196.470 35.625 196.515 ;
        RECT 36.700 196.470 37.020 196.530 ;
        RECT 35.335 196.330 37.020 196.470 ;
        RECT 35.335 196.285 35.625 196.330 ;
        RECT 36.700 196.270 37.020 196.330 ;
        RECT 37.175 196.470 37.465 196.515 ;
        RECT 37.620 196.470 37.940 196.530 ;
        RECT 37.175 196.330 37.940 196.470 ;
        RECT 37.175 196.285 37.465 196.330 ;
        RECT 37.620 196.270 37.940 196.330 ;
        RECT 39.015 196.470 39.305 196.515 ;
        RECT 41.300 196.470 41.620 196.530 ;
        RECT 39.015 196.330 41.620 196.470 ;
        RECT 39.015 196.285 39.305 196.330 ;
        RECT 41.300 196.270 41.620 196.330 ;
        RECT 43.140 196.470 43.460 196.530 ;
        RECT 45.440 196.470 45.760 196.530 ;
        RECT 50.975 196.470 51.265 196.515 ;
        RECT 43.140 196.330 45.760 196.470 ;
        RECT 43.140 196.270 43.460 196.330 ;
        RECT 45.440 196.270 45.760 196.330 ;
        RECT 45.990 196.330 51.265 196.470 ;
        RECT 38.095 196.130 38.385 196.175 ;
        RECT 30.350 195.990 38.385 196.130 ;
        RECT 18.315 195.790 18.605 195.835 ;
        RECT 24.370 195.790 24.510 195.945 ;
        RECT 27.040 195.930 27.360 195.990 ;
        RECT 38.095 195.945 38.385 195.990 ;
        RECT 38.540 196.130 38.860 196.190 ;
        RECT 45.990 196.130 46.130 196.330 ;
        RECT 50.975 196.285 51.265 196.330 ;
        RECT 51.895 196.470 52.185 196.515 ;
        RECT 52.890 196.470 53.030 196.670 ;
        RECT 60.620 196.610 60.940 196.670 ;
        RECT 51.895 196.330 53.030 196.470 ;
        RECT 53.260 196.470 53.580 196.530 ;
        RECT 59.700 196.470 60.020 196.530 ;
        RECT 63.930 196.515 64.070 197.350 ;
        RECT 78.560 197.290 78.880 197.350 ;
        RECT 84.095 197.490 84.385 197.535 ;
        RECT 85.000 197.490 85.320 197.550 ;
        RECT 84.095 197.350 85.320 197.490 ;
        RECT 84.095 197.305 84.385 197.350 ;
        RECT 85.000 197.290 85.320 197.350 ;
        RECT 73.515 197.150 73.805 197.195 ;
        RECT 82.700 197.150 83.020 197.210 ;
        RECT 73.515 197.010 83.020 197.150 ;
        RECT 73.515 196.965 73.805 197.010 ;
        RECT 82.700 196.950 83.020 197.010 ;
        RECT 68.440 196.810 68.760 196.870 ;
        RECT 69.820 196.810 70.140 196.870 ;
        RECT 76.720 196.810 77.040 196.870 ;
        RECT 65.770 196.670 68.760 196.810 ;
        RECT 53.260 196.330 60.020 196.470 ;
        RECT 51.895 196.285 52.185 196.330 ;
        RECT 38.540 195.990 46.130 196.130 ;
        RECT 24.740 195.790 25.060 195.850 ;
        RECT 18.315 195.650 25.060 195.790 ;
        RECT 18.315 195.605 18.605 195.650 ;
        RECT 24.740 195.590 25.060 195.650 ;
        RECT 25.200 195.790 25.520 195.850 ;
        RECT 26.135 195.790 26.425 195.835 ;
        RECT 25.200 195.650 26.425 195.790 ;
        RECT 25.200 195.590 25.520 195.650 ;
        RECT 26.135 195.605 26.425 195.650 ;
        RECT 28.420 195.790 28.740 195.850 ;
        RECT 31.180 195.790 31.500 195.850 ;
        RECT 28.420 195.650 31.500 195.790 ;
        RECT 28.420 195.590 28.740 195.650 ;
        RECT 31.180 195.590 31.500 195.650 ;
        RECT 31.640 195.790 31.960 195.850 ;
        RECT 35.780 195.790 36.100 195.850 ;
        RECT 31.640 195.650 36.100 195.790 ;
        RECT 31.640 195.590 31.960 195.650 ;
        RECT 35.780 195.590 36.100 195.650 ;
        RECT 36.255 195.790 36.545 195.835 ;
        RECT 37.620 195.790 37.940 195.850 ;
        RECT 36.255 195.650 37.940 195.790 ;
        RECT 38.170 195.790 38.310 195.945 ;
        RECT 38.540 195.930 38.860 195.990 ;
        RECT 49.135 195.945 49.425 196.175 ;
        RECT 49.580 196.130 49.900 196.190 ;
        RECT 51.970 196.130 52.110 196.285 ;
        RECT 53.260 196.270 53.580 196.330 ;
        RECT 59.700 196.270 60.020 196.330 ;
        RECT 63.855 196.285 64.145 196.515 ;
        RECT 64.315 196.470 64.605 196.515 ;
        RECT 65.770 196.470 65.910 196.670 ;
        RECT 68.440 196.610 68.760 196.670 ;
        RECT 68.990 196.670 70.140 196.810 ;
        RECT 68.990 196.515 69.130 196.670 ;
        RECT 69.820 196.610 70.140 196.670 ;
        RECT 70.370 196.670 77.040 196.810 ;
        RECT 64.315 196.330 65.910 196.470 ;
        RECT 64.315 196.285 64.605 196.330 ;
        RECT 68.915 196.285 69.205 196.515 ;
        RECT 69.360 196.270 69.680 196.530 ;
        RECT 70.370 196.515 70.510 196.670 ;
        RECT 76.720 196.610 77.040 196.670 ;
        RECT 70.295 196.285 70.585 196.515 ;
        RECT 70.740 196.270 71.060 196.530 ;
        RECT 80.400 196.270 80.720 196.530 ;
        RECT 80.860 196.470 81.180 196.530 ;
        RECT 82.715 196.470 83.005 196.515 ;
        RECT 80.860 196.330 83.005 196.470 ;
        RECT 80.860 196.270 81.180 196.330 ;
        RECT 82.715 196.285 83.005 196.330 ;
        RECT 83.160 196.270 83.480 196.530 ;
        RECT 84.540 196.270 84.860 196.530 ;
        RECT 49.580 195.990 52.110 196.130 ;
        RECT 39.000 195.790 39.320 195.850 ;
        RECT 41.760 195.790 42.080 195.850 ;
        RECT 38.170 195.650 42.080 195.790 ;
        RECT 36.255 195.605 36.545 195.650 ;
        RECT 37.620 195.590 37.940 195.650 ;
        RECT 39.000 195.590 39.320 195.650 ;
        RECT 41.760 195.590 42.080 195.650 ;
        RECT 42.220 195.790 42.540 195.850 ;
        RECT 42.695 195.790 42.985 195.835 ;
        RECT 44.060 195.790 44.380 195.850 ;
        RECT 42.220 195.650 44.380 195.790 ;
        RECT 42.220 195.590 42.540 195.650 ;
        RECT 42.695 195.605 42.985 195.650 ;
        RECT 44.060 195.590 44.380 195.650 ;
        RECT 44.520 195.790 44.840 195.850 ;
        RECT 47.740 195.790 48.060 195.850 ;
        RECT 44.520 195.650 48.060 195.790 ;
        RECT 49.210 195.790 49.350 195.945 ;
        RECT 49.580 195.930 49.900 195.990 ;
        RECT 55.115 195.945 55.405 196.175 ;
        RECT 64.390 195.990 65.910 196.130 ;
        RECT 55.190 195.790 55.330 195.945 ;
        RECT 64.390 195.850 64.530 195.990 ;
        RECT 62.000 195.790 62.320 195.850 ;
        RECT 49.210 195.650 62.320 195.790 ;
        RECT 44.520 195.590 44.840 195.650 ;
        RECT 47.740 195.590 48.060 195.650 ;
        RECT 62.000 195.590 62.320 195.650 ;
        RECT 64.300 195.590 64.620 195.850 ;
        RECT 65.220 195.590 65.540 195.850 ;
        RECT 65.770 195.835 65.910 195.990 ;
        RECT 66.140 195.930 66.460 196.190 ;
        RECT 67.075 196.130 67.365 196.175 ;
        RECT 67.075 195.990 72.580 196.130 ;
        RECT 67.075 195.945 67.365 195.990 ;
        RECT 65.695 195.605 65.985 195.835 ;
        RECT 66.600 195.790 66.920 195.850 ;
        RECT 67.995 195.790 68.285 195.835 ;
        RECT 66.600 195.650 68.285 195.790 ;
        RECT 72.440 195.790 72.580 195.990 ;
        RECT 79.940 195.930 80.260 196.190 ;
        RECT 80.490 196.130 80.630 196.270 ;
        RECT 80.490 195.990 81.090 196.130 ;
        RECT 80.400 195.790 80.720 195.850 ;
        RECT 80.950 195.835 81.090 195.990 ;
        RECT 72.440 195.650 80.720 195.790 ;
        RECT 66.600 195.590 66.920 195.650 ;
        RECT 67.995 195.605 68.285 195.650 ;
        RECT 80.400 195.590 80.720 195.650 ;
        RECT 80.875 195.605 81.165 195.835 ;
        RECT 85.000 195.590 85.320 195.850 ;
        RECT 15.930 194.970 87.230 195.450 ;
        RECT 18.760 194.770 19.080 194.830 ;
        RECT 20.615 194.770 20.905 194.815 ;
        RECT 18.760 194.630 20.905 194.770 ;
        RECT 18.760 194.570 19.080 194.630 ;
        RECT 20.615 194.585 20.905 194.630 ;
        RECT 21.060 194.770 21.380 194.830 ;
        RECT 22.455 194.770 22.745 194.815 ;
        RECT 23.360 194.770 23.680 194.830 ;
        RECT 21.060 194.630 23.680 194.770 ;
        RECT 21.060 194.570 21.380 194.630 ;
        RECT 22.455 194.585 22.745 194.630 ;
        RECT 23.360 194.570 23.680 194.630 ;
        RECT 25.660 194.770 25.980 194.830 ;
        RECT 26.595 194.770 26.885 194.815 ;
        RECT 34.860 194.770 35.180 194.830 ;
        RECT 25.660 194.630 26.885 194.770 ;
        RECT 25.660 194.570 25.980 194.630 ;
        RECT 26.595 194.585 26.885 194.630 ;
        RECT 27.590 194.630 31.410 194.770 ;
        RECT 15.080 194.430 15.400 194.490 ;
        RECT 27.590 194.430 27.730 194.630 ;
        RECT 15.080 194.290 19.450 194.430 ;
        RECT 15.080 194.230 15.400 194.290 ;
        RECT 18.760 193.890 19.080 194.150 ;
        RECT 19.310 194.135 19.450 194.290 ;
        RECT 25.750 194.290 27.730 194.430 ;
        RECT 19.235 193.905 19.525 194.135 ;
        RECT 21.535 194.090 21.825 194.135 ;
        RECT 22.440 194.090 22.760 194.150 ;
        RECT 21.535 193.950 22.760 194.090 ;
        RECT 21.535 193.905 21.825 193.950 ;
        RECT 17.840 193.750 18.160 193.810 ;
        RECT 21.610 193.750 21.750 193.905 ;
        RECT 22.440 193.890 22.760 193.950 ;
        RECT 22.915 193.905 23.205 194.135 ;
        RECT 24.755 194.090 25.045 194.135 ;
        RECT 25.200 194.090 25.520 194.150 ;
        RECT 25.750 194.135 25.890 194.290 ;
        RECT 28.420 194.230 28.740 194.490 ;
        RECT 24.755 193.950 25.520 194.090 ;
        RECT 24.755 193.905 25.045 193.950 ;
        RECT 17.840 193.610 21.750 193.750 ;
        RECT 17.840 193.550 18.160 193.610 ;
        RECT 22.990 193.410 23.130 193.905 ;
        RECT 25.200 193.890 25.520 193.950 ;
        RECT 25.675 193.905 25.965 194.135 ;
        RECT 26.135 193.905 26.425 194.135 ;
        RECT 26.580 194.090 26.900 194.150 ;
        RECT 27.515 194.090 27.805 194.135 ;
        RECT 26.580 193.950 27.805 194.090 ;
        RECT 23.360 193.750 23.680 193.810 ;
        RECT 25.750 193.750 25.890 193.905 ;
        RECT 23.360 193.610 25.890 193.750 ;
        RECT 26.210 193.750 26.350 193.905 ;
        RECT 26.580 193.890 26.900 193.950 ;
        RECT 27.515 193.905 27.805 193.950 ;
        RECT 29.340 193.890 29.660 194.150 ;
        RECT 29.800 194.090 30.120 194.150 ;
        RECT 31.270 194.135 31.410 194.630 ;
        RECT 31.730 194.630 35.180 194.770 ;
        RECT 31.730 194.490 31.870 194.630 ;
        RECT 34.860 194.570 35.180 194.630 ;
        RECT 38.095 194.585 38.385 194.815 ;
        RECT 40.855 194.770 41.145 194.815 ;
        RECT 43.140 194.770 43.460 194.830 ;
        RECT 48.200 194.770 48.520 194.830 ;
        RECT 40.855 194.630 43.460 194.770 ;
        RECT 40.855 194.585 41.145 194.630 ;
        RECT 31.640 194.230 31.960 194.490 ;
        RECT 32.115 194.430 32.405 194.475 ;
        RECT 37.620 194.430 37.940 194.490 ;
        RECT 32.115 194.290 37.940 194.430 ;
        RECT 38.170 194.430 38.310 194.585 ;
        RECT 43.140 194.570 43.460 194.630 ;
        RECT 43.690 194.630 48.520 194.770 ;
        RECT 43.690 194.475 43.830 194.630 ;
        RECT 48.200 194.570 48.520 194.630 ;
        RECT 50.975 194.770 51.265 194.815 ;
        RECT 51.880 194.770 52.200 194.830 ;
        RECT 50.975 194.630 52.200 194.770 ;
        RECT 50.975 194.585 51.265 194.630 ;
        RECT 51.880 194.570 52.200 194.630 ;
        RECT 60.635 194.585 60.925 194.815 ;
        RECT 65.680 194.770 66.000 194.830 ;
        RECT 68.915 194.770 69.205 194.815 ;
        RECT 84.540 194.770 84.860 194.830 ;
        RECT 65.680 194.630 69.205 194.770 ;
        RECT 38.170 194.290 43.370 194.430 ;
        RECT 32.115 194.245 32.405 194.290 ;
        RECT 37.620 194.230 37.940 194.290 ;
        RECT 43.230 194.150 43.370 194.290 ;
        RECT 43.615 194.245 43.905 194.475 ;
        RECT 44.075 194.430 44.365 194.475 ;
        RECT 44.520 194.430 44.840 194.490 ;
        RECT 44.075 194.290 44.840 194.430 ;
        RECT 44.075 194.245 44.365 194.290 ;
        RECT 44.520 194.230 44.840 194.290 ;
        RECT 45.440 194.430 45.760 194.490 ;
        RECT 49.580 194.430 49.900 194.490 ;
        RECT 45.440 194.290 49.900 194.430 ;
        RECT 45.440 194.230 45.760 194.290 ;
        RECT 49.580 194.230 49.900 194.290 ;
        RECT 57.860 194.430 58.180 194.490 ;
        RECT 60.710 194.430 60.850 194.585 ;
        RECT 65.680 194.570 66.000 194.630 ;
        RECT 68.915 194.585 69.205 194.630 ;
        RECT 72.440 194.630 84.860 194.770 ;
        RECT 72.440 194.430 72.580 194.630 ;
        RECT 84.540 194.570 84.860 194.630 ;
        RECT 85.000 194.430 85.320 194.490 ;
        RECT 57.860 194.290 72.580 194.430 ;
        RECT 74.050 194.290 85.320 194.430 ;
        RECT 57.860 194.230 58.180 194.290 ;
        RECT 30.735 194.090 31.025 194.135 ;
        RECT 29.800 193.950 31.025 194.090 ;
        RECT 29.800 193.890 30.120 193.950 ;
        RECT 30.735 193.905 31.025 193.950 ;
        RECT 31.195 194.090 31.485 194.135 ;
        RECT 33.480 194.090 33.800 194.150 ;
        RECT 31.195 193.950 33.800 194.090 ;
        RECT 31.195 193.905 31.485 193.950 ;
        RECT 33.480 193.890 33.800 193.950 ;
        RECT 33.940 194.090 34.260 194.150 ;
        RECT 34.415 194.090 34.705 194.135 ;
        RECT 33.940 193.950 34.705 194.090 ;
        RECT 33.940 193.890 34.260 193.950 ;
        RECT 34.415 193.905 34.705 193.950 ;
        RECT 29.890 193.750 30.030 193.890 ;
        RECT 26.210 193.610 30.030 193.750 ;
        RECT 34.490 193.750 34.630 193.905 ;
        RECT 35.320 193.890 35.640 194.150 ;
        RECT 38.555 194.090 38.845 194.135 ;
        RECT 40.840 194.090 41.160 194.150 ;
        RECT 38.555 193.950 41.160 194.090 ;
        RECT 38.555 193.905 38.845 193.950 ;
        RECT 40.840 193.890 41.160 193.950 ;
        RECT 43.140 193.890 43.460 194.150 ;
        RECT 44.980 193.890 45.300 194.150 ;
        RECT 46.375 194.110 46.665 194.135 ;
        RECT 45.990 193.970 46.665 194.110 ;
        RECT 35.780 193.750 36.100 193.810 ;
        RECT 34.490 193.610 36.100 193.750 ;
        RECT 23.360 193.550 23.680 193.610 ;
        RECT 35.780 193.550 36.100 193.610 ;
        RECT 37.160 193.750 37.480 193.810 ;
        RECT 39.935 193.750 40.225 193.795 ;
        RECT 42.220 193.750 42.540 193.810 ;
        RECT 37.160 193.610 37.850 193.750 ;
        RECT 37.160 193.550 37.480 193.610 ;
        RECT 26.580 193.410 26.900 193.470 ;
        RECT 22.990 193.270 26.900 193.410 ;
        RECT 26.580 193.210 26.900 193.270 ;
        RECT 29.800 193.410 30.120 193.470 ;
        RECT 30.275 193.410 30.565 193.455 ;
        RECT 29.800 193.270 30.565 193.410 ;
        RECT 29.800 193.210 30.120 193.270 ;
        RECT 30.275 193.225 30.565 193.270 ;
        RECT 32.115 193.410 32.405 193.455 ;
        RECT 33.940 193.410 34.260 193.470 ;
        RECT 32.115 193.270 34.260 193.410 ;
        RECT 32.115 193.225 32.405 193.270 ;
        RECT 33.940 193.210 34.260 193.270 ;
        RECT 34.860 193.410 35.180 193.470 ;
        RECT 37.710 193.455 37.850 193.610 ;
        RECT 39.935 193.610 42.540 193.750 ;
        RECT 45.990 193.750 46.130 193.970 ;
        RECT 46.375 193.905 46.665 193.970 ;
        RECT 46.835 194.090 47.125 194.135 ;
        RECT 47.740 194.090 48.060 194.150 ;
        RECT 46.835 193.950 48.060 194.090 ;
        RECT 46.835 193.905 47.125 193.950 ;
        RECT 47.740 193.890 48.060 193.950 ;
        RECT 48.200 193.890 48.520 194.150 ;
        RECT 57.400 193.890 57.720 194.150 ;
        RECT 67.075 194.090 67.365 194.135 ;
        RECT 68.900 194.090 69.220 194.150 ;
        RECT 74.050 194.135 74.190 194.290 ;
        RECT 85.000 194.230 85.320 194.290 ;
        RECT 67.075 193.950 69.220 194.090 ;
        RECT 67.075 193.905 67.365 193.950 ;
        RECT 68.900 193.890 69.220 193.950 ;
        RECT 69.450 193.950 70.510 194.090 ;
        RECT 56.020 193.750 56.340 193.810 ;
        RECT 45.990 193.610 56.340 193.750 ;
        RECT 39.935 193.565 40.225 193.610 ;
        RECT 42.220 193.550 42.540 193.610 ;
        RECT 56.020 193.550 56.340 193.610 ;
        RECT 65.680 193.750 66.000 193.810 ;
        RECT 67.980 193.750 68.300 193.810 ;
        RECT 65.680 193.610 68.300 193.750 ;
        RECT 65.680 193.550 66.000 193.610 ;
        RECT 67.980 193.550 68.300 193.610 ;
        RECT 34.860 193.270 37.390 193.410 ;
        RECT 34.860 193.210 35.180 193.270 ;
        RECT 14.620 193.070 14.940 193.130 ;
        RECT 17.855 193.070 18.145 193.115 ;
        RECT 14.620 192.930 18.145 193.070 ;
        RECT 14.620 192.870 14.940 192.930 ;
        RECT 17.855 192.885 18.145 192.930 ;
        RECT 19.220 193.070 19.540 193.130 ;
        RECT 20.155 193.070 20.445 193.115 ;
        RECT 20.600 193.070 20.920 193.130 ;
        RECT 19.220 192.930 20.920 193.070 ;
        RECT 19.220 192.870 19.540 192.930 ;
        RECT 20.155 192.885 20.445 192.930 ;
        RECT 20.600 192.870 20.920 192.930 ;
        RECT 23.835 193.070 24.125 193.115 ;
        RECT 24.280 193.070 24.600 193.130 ;
        RECT 23.835 192.930 24.600 193.070 ;
        RECT 23.835 192.885 24.125 192.930 ;
        RECT 24.280 192.870 24.600 192.930 ;
        RECT 26.120 193.070 26.440 193.130 ;
        RECT 33.495 193.070 33.785 193.115 ;
        RECT 36.240 193.070 36.560 193.130 ;
        RECT 26.120 192.930 36.560 193.070 ;
        RECT 37.250 193.070 37.390 193.270 ;
        RECT 37.635 193.225 37.925 193.455 ;
        RECT 39.015 193.410 39.305 193.455 ;
        RECT 39.460 193.410 39.780 193.470 ;
        RECT 45.440 193.410 45.760 193.470 ;
        RECT 39.015 193.270 39.780 193.410 ;
        RECT 39.015 193.225 39.305 193.270 ;
        RECT 39.460 193.210 39.780 193.270 ;
        RECT 41.390 193.270 45.760 193.410 ;
        RECT 41.390 193.070 41.530 193.270 ;
        RECT 45.440 193.210 45.760 193.270 ;
        RECT 47.755 193.410 48.045 193.455 ;
        RECT 69.450 193.410 69.590 193.950 ;
        RECT 69.835 193.565 70.125 193.795 ;
        RECT 47.755 193.270 69.590 193.410 ;
        RECT 47.755 193.225 48.045 193.270 ;
        RECT 37.250 192.930 41.530 193.070 ;
        RECT 41.760 193.070 42.080 193.130 ;
        RECT 42.235 193.070 42.525 193.115 ;
        RECT 41.760 192.930 42.525 193.070 ;
        RECT 26.120 192.870 26.440 192.930 ;
        RECT 33.495 192.885 33.785 192.930 ;
        RECT 36.240 192.870 36.560 192.930 ;
        RECT 41.760 192.870 42.080 192.930 ;
        RECT 42.235 192.885 42.525 192.930 ;
        RECT 48.200 193.070 48.520 193.130 ;
        RECT 54.640 193.070 54.960 193.130 ;
        RECT 48.200 192.930 54.960 193.070 ;
        RECT 48.200 192.870 48.520 192.930 ;
        RECT 54.640 192.870 54.960 192.930 ;
        RECT 55.560 193.070 55.880 193.130 ;
        RECT 58.780 193.070 59.100 193.130 ;
        RECT 55.560 192.930 59.100 193.070 ;
        RECT 55.560 192.870 55.880 192.930 ;
        RECT 58.780 192.870 59.100 192.930 ;
        RECT 59.700 193.070 60.020 193.130 ;
        RECT 69.910 193.070 70.050 193.565 ;
        RECT 70.370 193.410 70.510 193.950 ;
        RECT 73.975 193.905 74.265 194.135 ;
        RECT 74.420 193.890 74.740 194.150 ;
        RECT 75.340 193.890 75.660 194.150 ;
        RECT 85.460 193.890 85.780 194.150 ;
        RECT 72.580 193.750 72.900 193.810 ;
        RECT 73.055 193.750 73.345 193.795 ;
        RECT 72.580 193.610 73.345 193.750 ;
        RECT 72.580 193.550 72.900 193.610 ;
        RECT 73.055 193.565 73.345 193.610 ;
        RECT 73.515 193.750 73.805 193.795 ;
        RECT 73.515 193.610 73.915 193.750 ;
        RECT 73.515 193.565 73.805 193.610 ;
        RECT 73.590 193.410 73.730 193.565 ;
        RECT 77.640 193.410 77.960 193.470 ;
        RECT 70.370 193.270 77.960 193.410 ;
        RECT 77.640 193.210 77.960 193.270 ;
        RECT 79.035 193.410 79.325 193.455 ;
        RECT 79.480 193.410 79.800 193.470 ;
        RECT 79.035 193.270 79.800 193.410 ;
        RECT 79.035 193.225 79.325 193.270 ;
        RECT 79.480 193.210 79.800 193.270 ;
        RECT 79.940 193.410 80.260 193.470 ;
        RECT 82.240 193.410 82.560 193.470 ;
        RECT 79.940 193.270 82.560 193.410 ;
        RECT 79.940 193.210 80.260 193.270 ;
        RECT 82.240 193.210 82.560 193.270 ;
        RECT 59.700 192.930 70.050 193.070 ;
        RECT 70.755 193.070 71.045 193.115 ;
        RECT 71.200 193.070 71.520 193.130 ;
        RECT 70.755 192.930 71.520 193.070 ;
        RECT 59.700 192.870 60.020 192.930 ;
        RECT 70.755 192.885 71.045 192.930 ;
        RECT 71.200 192.870 71.520 192.930 ;
        RECT 72.120 192.870 72.440 193.130 ;
        RECT 15.930 192.250 87.230 192.730 ;
        RECT 21.075 192.050 21.365 192.095 ;
        RECT 21.520 192.050 21.840 192.110 ;
        RECT 21.075 191.910 21.840 192.050 ;
        RECT 21.075 191.865 21.365 191.910 ;
        RECT 21.520 191.850 21.840 191.910 ;
        RECT 27.040 192.050 27.360 192.110 ;
        RECT 39.460 192.050 39.780 192.110 ;
        RECT 27.040 191.910 39.780 192.050 ;
        RECT 27.040 191.850 27.360 191.910 ;
        RECT 39.460 191.850 39.780 191.910 ;
        RECT 40.380 191.850 40.700 192.110 ;
        RECT 41.300 192.050 41.620 192.110 ;
        RECT 48.200 192.050 48.520 192.110 ;
        RECT 41.300 191.910 48.520 192.050 ;
        RECT 41.300 191.850 41.620 191.910 ;
        RECT 48.200 191.850 48.520 191.910 ;
        RECT 50.500 191.850 50.820 192.110 ;
        RECT 51.880 192.050 52.200 192.110 ;
        RECT 53.260 192.050 53.580 192.110 ;
        RECT 51.880 191.910 53.580 192.050 ;
        RECT 51.880 191.850 52.200 191.910 ;
        RECT 53.260 191.850 53.580 191.910 ;
        RECT 54.195 192.050 54.485 192.095 ;
        RECT 54.640 192.050 54.960 192.110 ;
        RECT 54.195 191.910 54.960 192.050 ;
        RECT 54.195 191.865 54.485 191.910 ;
        RECT 54.640 191.850 54.960 191.910 ;
        RECT 55.560 192.050 55.880 192.110 ;
        RECT 58.335 192.050 58.625 192.095 ;
        RECT 69.360 192.050 69.680 192.110 ;
        RECT 55.560 191.910 58.625 192.050 ;
        RECT 55.560 191.850 55.880 191.910 ;
        RECT 58.335 191.865 58.625 191.910 ;
        RECT 59.790 191.910 69.680 192.050 ;
        RECT 17.380 191.710 17.700 191.770 ;
        RECT 23.375 191.710 23.665 191.755 ;
        RECT 17.380 191.570 23.665 191.710 ;
        RECT 17.380 191.510 17.700 191.570 ;
        RECT 23.375 191.525 23.665 191.570 ;
        RECT 23.820 191.710 24.140 191.770 ;
        RECT 26.595 191.710 26.885 191.755 ;
        RECT 35.320 191.710 35.640 191.770 ;
        RECT 35.795 191.710 36.085 191.755 ;
        RECT 23.820 191.570 35.090 191.710 ;
        RECT 23.820 191.510 24.140 191.570 ;
        RECT 26.595 191.525 26.885 191.570 ;
        RECT 22.900 191.370 23.220 191.430 ;
        RECT 19.310 191.230 23.220 191.370 ;
        RECT 18.760 190.830 19.080 191.090 ;
        RECT 19.310 191.075 19.450 191.230 ;
        RECT 22.900 191.170 23.220 191.230 ;
        RECT 29.340 191.370 29.660 191.430 ;
        RECT 31.180 191.370 31.500 191.430 ;
        RECT 29.340 191.230 31.500 191.370 ;
        RECT 29.340 191.170 29.660 191.230 ;
        RECT 31.180 191.170 31.500 191.230 ;
        RECT 32.560 191.370 32.880 191.430 ;
        RECT 33.495 191.370 33.785 191.415 ;
        RECT 33.940 191.370 34.260 191.430 ;
        RECT 32.560 191.230 34.260 191.370 ;
        RECT 34.950 191.370 35.090 191.570 ;
        RECT 35.320 191.570 36.085 191.710 ;
        RECT 35.320 191.510 35.640 191.570 ;
        RECT 35.795 191.525 36.085 191.570 ;
        RECT 36.700 191.510 37.020 191.770 ;
        RECT 37.160 191.710 37.480 191.770 ;
        RECT 37.635 191.710 37.925 191.755 ;
        RECT 37.160 191.570 37.925 191.710 ;
        RECT 37.160 191.510 37.480 191.570 ;
        RECT 37.635 191.525 37.925 191.570 ;
        RECT 42.680 191.710 43.000 191.770 ;
        RECT 44.980 191.710 45.300 191.770 ;
        RECT 48.660 191.710 48.980 191.770 ;
        RECT 42.680 191.570 45.300 191.710 ;
        RECT 42.680 191.510 43.000 191.570 ;
        RECT 44.980 191.510 45.300 191.570 ;
        RECT 45.990 191.570 48.980 191.710 ;
        RECT 34.950 191.230 36.010 191.370 ;
        RECT 32.560 191.170 32.880 191.230 ;
        RECT 33.495 191.185 33.785 191.230 ;
        RECT 33.940 191.170 34.260 191.230 ;
        RECT 19.235 190.845 19.525 191.075 ;
        RECT 20.140 191.030 20.460 191.090 ;
        RECT 20.615 191.030 20.905 191.075 ;
        RECT 21.060 191.030 21.380 191.090 ;
        RECT 20.140 190.890 21.380 191.030 ;
        RECT 20.140 190.830 20.460 190.890 ;
        RECT 20.615 190.845 20.905 190.890 ;
        RECT 21.060 190.830 21.380 190.890 ;
        RECT 21.995 191.030 22.285 191.075 ;
        RECT 26.580 191.030 26.900 191.090 ;
        RECT 21.995 190.890 26.900 191.030 ;
        RECT 21.995 190.845 22.285 190.890 ;
        RECT 26.580 190.830 26.900 190.890 ;
        RECT 27.515 190.845 27.805 191.075 ;
        RECT 18.850 190.690 18.990 190.830 ;
        RECT 23.835 190.690 24.125 190.735 ;
        RECT 18.850 190.550 19.910 190.690 ;
        RECT 18.315 190.350 18.605 190.395 ;
        RECT 18.760 190.350 19.080 190.410 ;
        RECT 19.770 190.395 19.910 190.550 ;
        RECT 22.990 190.550 24.125 190.690 ;
        RECT 18.315 190.210 19.080 190.350 ;
        RECT 18.315 190.165 18.605 190.210 ;
        RECT 18.760 190.150 19.080 190.210 ;
        RECT 19.695 190.165 19.985 190.395 ;
        RECT 22.440 190.350 22.760 190.410 ;
        RECT 22.990 190.350 23.130 190.550 ;
        RECT 23.835 190.505 24.125 190.550 ;
        RECT 24.280 190.690 24.600 190.750 ;
        RECT 24.755 190.690 25.045 190.735 ;
        RECT 24.280 190.550 25.045 190.690 ;
        RECT 27.590 190.690 27.730 190.845 ;
        RECT 34.860 190.830 35.180 191.090 ;
        RECT 27.960 190.690 28.280 190.750 ;
        RECT 27.590 190.550 28.280 190.690 ;
        RECT 35.870 190.690 36.010 191.230 ;
        RECT 36.255 191.030 36.545 191.075 ;
        RECT 36.790 191.030 36.930 191.510 ;
        RECT 36.255 190.890 36.930 191.030 ;
        RECT 36.255 190.845 36.545 190.890 ;
        RECT 37.620 190.830 37.940 191.090 ;
        RECT 41.300 191.030 41.620 191.090 ;
        RECT 45.990 191.030 46.130 191.570 ;
        RECT 48.660 191.510 48.980 191.570 ;
        RECT 49.120 191.510 49.440 191.770 ;
        RECT 49.210 191.370 49.350 191.510 ;
        RECT 50.590 191.415 50.730 191.850 ;
        RECT 47.370 191.230 49.350 191.370 ;
        RECT 41.300 190.890 46.130 191.030 ;
        RECT 41.300 190.830 41.620 190.890 ;
        RECT 46.820 190.830 47.140 191.090 ;
        RECT 47.370 191.075 47.510 191.230 ;
        RECT 50.515 191.185 50.805 191.415 ;
        RECT 47.295 190.845 47.585 191.075 ;
        RECT 48.215 190.845 48.505 191.075 ;
        RECT 44.520 190.690 44.840 190.750 ;
        RECT 35.870 190.550 44.840 190.690 ;
        RECT 24.280 190.490 24.600 190.550 ;
        RECT 24.755 190.505 25.045 190.550 ;
        RECT 27.960 190.490 28.280 190.550 ;
        RECT 44.520 190.490 44.840 190.550 ;
        RECT 48.290 190.410 48.430 190.845 ;
        RECT 48.660 190.830 48.980 191.090 ;
        RECT 49.220 191.030 49.510 191.075 ;
        RECT 49.220 190.890 49.810 191.030 ;
        RECT 49.220 190.845 49.510 190.890 ;
        RECT 49.670 190.690 49.810 190.890 ;
        RECT 50.960 190.830 51.280 191.090 ;
        RECT 51.970 191.075 52.110 191.850 ;
        RECT 58.780 191.710 59.100 191.770 ;
        RECT 52.890 191.570 59.100 191.710 ;
        RECT 52.890 191.075 53.030 191.570 ;
        RECT 58.780 191.510 59.100 191.570 ;
        RECT 59.790 191.370 59.930 191.910 ;
        RECT 69.360 191.850 69.680 191.910 ;
        RECT 81.320 192.050 81.640 192.110 ;
        RECT 82.240 192.050 82.560 192.110 ;
        RECT 81.320 191.910 82.560 192.050 ;
        RECT 81.320 191.850 81.640 191.910 ;
        RECT 82.240 191.850 82.560 191.910 ;
        RECT 83.160 192.050 83.480 192.110 ;
        RECT 84.555 192.050 84.845 192.095 ;
        RECT 83.160 191.910 84.845 192.050 ;
        RECT 83.160 191.850 83.480 191.910 ;
        RECT 84.555 191.865 84.845 191.910 ;
        RECT 76.720 191.710 77.040 191.770 ;
        RECT 76.720 191.570 85.690 191.710 ;
        RECT 76.720 191.510 77.040 191.570 ;
        RECT 54.730 191.230 59.930 191.370 ;
        RECT 60.175 191.410 60.465 191.415 ;
        RECT 60.175 191.370 61.310 191.410 ;
        RECT 66.140 191.370 66.460 191.430 ;
        RECT 75.340 191.370 75.660 191.430 ;
        RECT 79.020 191.370 79.340 191.430 ;
        RECT 60.175 191.270 79.340 191.370 ;
        RECT 51.765 190.890 52.110 191.075 ;
        RECT 51.765 190.845 52.055 190.890 ;
        RECT 52.815 190.845 53.105 191.075 ;
        RECT 53.275 191.030 53.565 191.075 ;
        RECT 54.180 191.030 54.500 191.090 ;
        RECT 53.275 190.890 54.500 191.030 ;
        RECT 53.275 190.845 53.565 190.890 ;
        RECT 54.180 190.830 54.500 190.890 ;
        RECT 50.500 190.690 50.820 190.750 ;
        RECT 49.670 190.550 50.820 190.690 ;
        RECT 50.500 190.490 50.820 190.550 ;
        RECT 52.340 190.490 52.660 190.750 ;
        RECT 22.440 190.210 23.130 190.350 ;
        RECT 25.675 190.350 25.965 190.395 ;
        RECT 26.120 190.350 26.440 190.410 ;
        RECT 25.675 190.210 26.440 190.350 ;
        RECT 22.440 190.150 22.760 190.210 ;
        RECT 25.675 190.165 25.965 190.210 ;
        RECT 26.120 190.150 26.440 190.210 ;
        RECT 27.040 190.350 27.360 190.410 ;
        RECT 30.275 190.350 30.565 190.395 ;
        RECT 27.040 190.210 30.565 190.350 ;
        RECT 27.040 190.150 27.360 190.210 ;
        RECT 30.275 190.165 30.565 190.210 ;
        RECT 32.100 190.150 32.420 190.410 ;
        RECT 32.575 190.350 32.865 190.395 ;
        RECT 33.020 190.350 33.340 190.410 ;
        RECT 32.575 190.210 33.340 190.350 ;
        RECT 32.575 190.165 32.865 190.210 ;
        RECT 33.020 190.150 33.340 190.210 ;
        RECT 33.480 190.350 33.800 190.410 ;
        RECT 36.715 190.350 37.005 190.395 ;
        RECT 33.480 190.210 37.005 190.350 ;
        RECT 33.480 190.150 33.800 190.210 ;
        RECT 36.715 190.165 37.005 190.210 ;
        RECT 48.200 190.150 48.520 190.410 ;
        RECT 49.120 190.350 49.440 190.410 ;
        RECT 54.730 190.350 54.870 191.230 ;
        RECT 60.175 191.185 60.465 191.270 ;
        RECT 61.170 191.230 79.340 191.270 ;
        RECT 66.140 191.170 66.460 191.230 ;
        RECT 75.340 191.170 75.660 191.230 ;
        RECT 79.020 191.170 79.340 191.230 ;
        RECT 80.860 191.370 81.180 191.430 ;
        RECT 84.095 191.370 84.385 191.415 ;
        RECT 80.860 191.230 84.385 191.370 ;
        RECT 80.860 191.170 81.180 191.230 ;
        RECT 84.095 191.185 84.385 191.230 ;
        RECT 56.940 190.830 57.260 191.090 ;
        RECT 58.795 191.030 59.085 191.075 ;
        RECT 59.240 191.030 59.560 191.090 ;
        RECT 58.795 190.890 59.560 191.030 ;
        RECT 58.795 190.845 59.085 190.890 ;
        RECT 49.120 190.210 54.870 190.350 ;
        RECT 58.870 190.350 59.010 190.845 ;
        RECT 59.240 190.830 59.560 190.890 ;
        RECT 59.700 190.830 60.020 191.090 ;
        RECT 60.815 190.900 61.105 191.045 ;
        RECT 60.815 190.815 61.310 190.900 ;
        RECT 61.540 190.830 61.860 191.090 ;
        RECT 62.000 190.830 62.320 191.090 ;
        RECT 69.360 191.030 69.680 191.090 ;
        RECT 70.755 191.030 71.045 191.075 ;
        RECT 80.400 191.030 80.720 191.090 ;
        RECT 82.255 191.030 82.545 191.075 ;
        RECT 69.360 190.890 76.030 191.030 ;
        RECT 69.360 190.830 69.680 190.890 ;
        RECT 70.755 190.845 71.045 190.890 ;
        RECT 60.890 190.760 61.310 190.815 ;
        RECT 61.170 190.690 61.310 190.760 ;
        RECT 75.340 190.690 75.660 190.750 ;
        RECT 61.170 190.550 75.660 190.690 ;
        RECT 75.340 190.490 75.660 190.550 ;
        RECT 67.520 190.350 67.840 190.410 ;
        RECT 58.870 190.210 67.840 190.350 ;
        RECT 49.120 190.150 49.440 190.210 ;
        RECT 67.520 190.150 67.840 190.210 ;
        RECT 68.900 190.350 69.220 190.410 ;
        RECT 72.595 190.350 72.885 190.395 ;
        RECT 68.900 190.210 72.885 190.350 ;
        RECT 75.890 190.350 76.030 190.890 ;
        RECT 80.400 190.890 82.545 191.030 ;
        RECT 80.400 190.830 80.720 190.890 ;
        RECT 82.255 190.845 82.545 190.890 ;
        RECT 85.000 190.830 85.320 191.090 ;
        RECT 85.550 191.075 85.690 191.570 ;
        RECT 85.475 190.845 85.765 191.075 ;
        RECT 79.940 190.490 80.260 190.750 ;
        RECT 80.875 190.690 81.165 190.735 ;
        RECT 80.875 190.550 82.010 190.690 ;
        RECT 80.875 190.505 81.165 190.550 ;
        RECT 81.335 190.350 81.625 190.395 ;
        RECT 75.890 190.210 81.625 190.350 ;
        RECT 81.870 190.350 82.010 190.550 ;
        RECT 83.160 190.490 83.480 190.750 ;
        RECT 84.540 190.350 84.860 190.410 ;
        RECT 81.870 190.210 84.860 190.350 ;
        RECT 68.900 190.150 69.220 190.210 ;
        RECT 72.595 190.165 72.885 190.210 ;
        RECT 81.335 190.165 81.625 190.210 ;
        RECT 84.540 190.150 84.860 190.210 ;
        RECT 15.930 189.530 87.230 190.010 ;
        RECT 14.620 189.330 14.940 189.390 ;
        RECT 17.855 189.330 18.145 189.375 ;
        RECT 21.980 189.330 22.300 189.390 ;
        RECT 14.620 189.190 18.145 189.330 ;
        RECT 14.620 189.130 14.940 189.190 ;
        RECT 17.855 189.145 18.145 189.190 ;
        RECT 19.310 189.190 22.300 189.330 ;
        RECT 18.760 188.450 19.080 188.710 ;
        RECT 19.310 188.695 19.450 189.190 ;
        RECT 21.980 189.130 22.300 189.190 ;
        RECT 23.820 189.330 24.140 189.390 ;
        RECT 25.675 189.330 25.965 189.375 ;
        RECT 35.780 189.330 36.100 189.390 ;
        RECT 41.300 189.330 41.620 189.390 ;
        RECT 23.820 189.190 25.965 189.330 ;
        RECT 23.820 189.130 24.140 189.190 ;
        RECT 25.675 189.145 25.965 189.190 ;
        RECT 28.510 189.190 35.550 189.330 ;
        RECT 19.695 188.990 19.985 189.035 ;
        RECT 21.520 188.990 21.840 189.050 ;
        RECT 23.375 188.990 23.665 189.035 ;
        RECT 28.510 188.990 28.650 189.190 ;
        RECT 19.695 188.850 21.290 188.990 ;
        RECT 19.695 188.805 19.985 188.850 ;
        RECT 21.150 188.695 21.290 188.850 ;
        RECT 21.520 188.850 23.130 188.990 ;
        RECT 21.520 188.790 21.840 188.850 ;
        RECT 19.235 188.465 19.525 188.695 ;
        RECT 20.155 188.650 20.445 188.695 ;
        RECT 20.155 188.510 20.830 188.650 ;
        RECT 20.155 188.465 20.445 188.510 ;
        RECT 20.690 187.970 20.830 188.510 ;
        RECT 21.075 188.465 21.365 188.695 ;
        RECT 21.980 188.450 22.300 188.710 ;
        RECT 22.440 188.450 22.760 188.710 ;
        RECT 22.990 188.650 23.130 188.850 ;
        RECT 23.375 188.850 28.650 188.990 ;
        RECT 33.035 188.990 33.325 189.035 ;
        RECT 35.410 188.990 35.550 189.190 ;
        RECT 35.780 189.190 41.620 189.330 ;
        RECT 35.780 189.130 36.100 189.190 ;
        RECT 41.300 189.130 41.620 189.190 ;
        RECT 41.760 189.330 42.080 189.390 ;
        RECT 42.695 189.330 42.985 189.375 ;
        RECT 41.760 189.190 42.985 189.330 ;
        RECT 41.760 189.130 42.080 189.190 ;
        RECT 42.695 189.145 42.985 189.190 ;
        RECT 44.060 189.130 44.380 189.390 ;
        RECT 46.820 189.130 47.140 189.390 ;
        RECT 49.120 189.130 49.440 189.390 ;
        RECT 62.920 189.330 63.240 189.390 ;
        RECT 52.890 189.190 63.240 189.330 ;
        RECT 49.210 188.990 49.350 189.130 ;
        RECT 33.035 188.850 34.630 188.990 ;
        RECT 35.410 188.850 46.630 188.990 ;
        RECT 23.375 188.805 23.665 188.850 ;
        RECT 33.035 188.805 33.325 188.850 ;
        RECT 25.380 188.650 25.670 188.695 ;
        RECT 22.990 188.510 25.670 188.650 ;
        RECT 25.380 188.465 25.670 188.510 ;
        RECT 26.120 188.650 26.440 188.710 ;
        RECT 27.515 188.650 27.805 188.695 ;
        RECT 26.120 188.510 27.805 188.650 ;
        RECT 26.120 188.450 26.440 188.510 ;
        RECT 27.515 188.465 27.805 188.510 ;
        RECT 27.960 188.450 28.280 188.710 ;
        RECT 28.420 188.450 28.740 188.710 ;
        RECT 29.355 188.465 29.645 188.695 ;
        RECT 29.815 188.650 30.105 188.695 ;
        RECT 31.180 188.650 31.500 188.710 ;
        RECT 29.815 188.510 31.500 188.650 ;
        RECT 29.815 188.465 30.105 188.510 ;
        RECT 21.535 188.310 21.825 188.355 ;
        RECT 22.900 188.310 23.220 188.370 ;
        RECT 21.535 188.170 23.220 188.310 ;
        RECT 21.535 188.125 21.825 188.170 ;
        RECT 22.900 188.110 23.220 188.170 ;
        RECT 24.280 188.310 24.600 188.370 ;
        RECT 29.430 188.310 29.570 188.465 ;
        RECT 24.280 188.170 29.570 188.310 ;
        RECT 24.280 188.110 24.600 188.170 ;
        RECT 23.360 187.970 23.680 188.030 ;
        RECT 20.690 187.830 23.680 187.970 ;
        RECT 23.360 187.770 23.680 187.830 ;
        RECT 28.435 187.970 28.725 188.015 ;
        RECT 29.890 187.970 30.030 188.465 ;
        RECT 31.180 188.450 31.500 188.510 ;
        RECT 32.560 188.650 32.880 188.710 ;
        RECT 34.490 188.650 34.630 188.850 ;
        RECT 35.320 188.650 35.640 188.710 ;
        RECT 37.175 188.650 37.465 188.695 ;
        RECT 32.560 188.640 33.710 188.650 ;
        RECT 32.560 188.510 34.170 188.640 ;
        RECT 34.490 188.510 37.465 188.650 ;
        RECT 32.560 188.450 32.880 188.510 ;
        RECT 33.570 188.500 34.170 188.510 ;
        RECT 30.260 188.310 30.580 188.370 ;
        RECT 34.030 188.355 34.170 188.500 ;
        RECT 35.320 188.450 35.640 188.510 ;
        RECT 37.175 188.465 37.465 188.510 ;
        RECT 37.635 188.650 37.925 188.695 ;
        RECT 39.920 188.650 40.240 188.710 ;
        RECT 43.140 188.650 43.460 188.710 ;
        RECT 37.635 188.510 39.690 188.650 ;
        RECT 37.635 188.465 37.925 188.510 ;
        RECT 30.260 188.170 31.870 188.310 ;
        RECT 30.260 188.110 30.580 188.170 ;
        RECT 28.435 187.830 30.030 187.970 ;
        RECT 31.730 187.970 31.870 188.170 ;
        RECT 33.495 188.125 33.785 188.355 ;
        RECT 33.955 188.125 34.245 188.355 ;
        RECT 37.710 188.310 37.850 188.465 ;
        RECT 34.490 188.170 37.850 188.310 ;
        RECT 33.570 187.970 33.710 188.125 ;
        RECT 34.490 187.970 34.630 188.170 ;
        RECT 38.095 188.125 38.385 188.355 ;
        RECT 31.730 187.830 33.250 187.970 ;
        RECT 33.570 187.830 34.630 187.970 ;
        RECT 37.160 187.970 37.480 188.030 ;
        RECT 38.170 187.970 38.310 188.125 ;
        RECT 37.160 187.830 38.310 187.970 ;
        RECT 39.550 187.970 39.690 188.510 ;
        RECT 39.920 188.510 43.460 188.650 ;
        RECT 39.920 188.450 40.240 188.510 ;
        RECT 43.140 188.450 43.460 188.510 ;
        RECT 41.300 188.310 41.620 188.370 ;
        RECT 43.615 188.310 43.905 188.355 ;
        RECT 41.300 188.170 43.905 188.310 ;
        RECT 41.300 188.110 41.620 188.170 ;
        RECT 43.615 188.125 43.905 188.170 ;
        RECT 44.520 188.310 44.840 188.370 ;
        RECT 44.995 188.310 45.285 188.355 ;
        RECT 44.520 188.170 45.285 188.310 ;
        RECT 46.490 188.310 46.630 188.850 ;
        RECT 48.290 188.850 49.350 188.990 ;
        RECT 50.500 188.990 50.820 189.050 ;
        RECT 52.890 189.035 53.030 189.190 ;
        RECT 62.920 189.130 63.240 189.190 ;
        RECT 69.360 189.130 69.680 189.390 ;
        RECT 74.880 189.330 75.200 189.390 ;
        RECT 83.160 189.330 83.480 189.390 ;
        RECT 74.880 189.190 83.480 189.330 ;
        RECT 74.880 189.130 75.200 189.190 ;
        RECT 83.160 189.130 83.480 189.190 ;
        RECT 50.500 188.850 51.650 188.990 ;
        RECT 46.835 188.650 47.125 188.695 ;
        RECT 47.280 188.650 47.600 188.710 ;
        RECT 46.835 188.510 47.600 188.650 ;
        RECT 46.835 188.465 47.125 188.510 ;
        RECT 47.280 188.450 47.600 188.510 ;
        RECT 47.740 188.450 48.060 188.710 ;
        RECT 48.290 188.695 48.430 188.850 ;
        RECT 50.500 188.790 50.820 188.850 ;
        RECT 48.215 188.465 48.505 188.695 ;
        RECT 48.955 188.465 49.245 188.695 ;
        RECT 50.975 188.465 51.265 188.695 ;
        RECT 49.030 188.310 49.170 188.465 ;
        RECT 46.490 188.170 49.170 188.310 ;
        RECT 44.520 188.110 44.840 188.170 ;
        RECT 44.995 188.125 45.285 188.170 ;
        RECT 49.595 188.125 49.885 188.355 ;
        RECT 41.760 187.970 42.080 188.030 ;
        RECT 39.550 187.830 42.080 187.970 ;
        RECT 28.435 187.785 28.725 187.830 ;
        RECT 24.755 187.630 25.045 187.675 ;
        RECT 25.660 187.630 25.980 187.690 ;
        RECT 24.755 187.490 25.980 187.630 ;
        RECT 24.755 187.445 25.045 187.490 ;
        RECT 25.660 187.430 25.980 187.490 ;
        RECT 29.800 187.630 30.120 187.690 ;
        RECT 30.275 187.630 30.565 187.675 ;
        RECT 29.800 187.490 30.565 187.630 ;
        RECT 29.800 187.430 30.120 187.490 ;
        RECT 30.275 187.445 30.565 187.490 ;
        RECT 31.195 187.630 31.485 187.675 ;
        RECT 31.640 187.630 31.960 187.690 ;
        RECT 31.195 187.490 31.960 187.630 ;
        RECT 33.110 187.630 33.250 187.830 ;
        RECT 37.160 187.770 37.480 187.830 ;
        RECT 41.760 187.770 42.080 187.830 ;
        RECT 46.415 187.970 46.705 188.015 ;
        RECT 47.740 187.970 48.060 188.030 ;
        RECT 49.670 187.970 49.810 188.125 ;
        RECT 50.040 188.110 50.360 188.370 ;
        RECT 50.500 188.310 50.820 188.370 ;
        RECT 51.050 188.310 51.190 188.465 ;
        RECT 50.500 188.170 51.190 188.310 ;
        RECT 51.510 188.310 51.650 188.850 ;
        RECT 52.815 188.805 53.105 189.035 ;
        RECT 53.260 188.990 53.580 189.050 ;
        RECT 56.940 188.990 57.260 189.050 ;
        RECT 53.260 188.850 57.260 188.990 ;
        RECT 53.260 188.790 53.580 188.850 ;
        RECT 56.940 188.790 57.260 188.850 ;
        RECT 57.415 188.990 57.705 189.035 ;
        RECT 57.860 188.990 58.180 189.050 ;
        RECT 57.415 188.850 58.180 188.990 ;
        RECT 57.415 188.805 57.705 188.850 ;
        RECT 57.860 188.790 58.180 188.850 ;
        RECT 67.075 188.990 67.365 189.035 ;
        RECT 73.040 188.990 73.360 189.050 ;
        RECT 67.075 188.850 73.360 188.990 ;
        RECT 67.075 188.805 67.365 188.850 ;
        RECT 73.040 188.790 73.360 188.850 ;
        RECT 84.080 188.990 84.400 189.050 ;
        RECT 85.015 188.990 85.305 189.035 ;
        RECT 84.080 188.850 85.305 188.990 ;
        RECT 84.080 188.790 84.400 188.850 ;
        RECT 85.015 188.805 85.305 188.850 ;
        RECT 51.895 188.650 52.185 188.695 ;
        RECT 52.355 188.650 52.645 188.695 ;
        RECT 51.895 188.510 52.645 188.650 ;
        RECT 51.895 188.465 52.185 188.510 ;
        RECT 52.355 188.465 52.645 188.510 ;
        RECT 54.195 188.650 54.485 188.695 ;
        RECT 55.100 188.650 55.420 188.710 ;
        RECT 69.065 188.650 69.355 188.695 ;
        RECT 54.195 188.510 55.420 188.650 ;
        RECT 54.195 188.465 54.485 188.510 ;
        RECT 55.100 188.450 55.420 188.510 ;
        RECT 63.470 188.510 69.355 188.650 ;
        RECT 63.470 188.370 63.610 188.510 ;
        RECT 69.065 188.465 69.355 188.510 ;
        RECT 71.675 188.650 71.965 188.695 ;
        RECT 72.120 188.650 72.440 188.710 ;
        RECT 71.675 188.510 72.440 188.650 ;
        RECT 71.675 188.465 71.965 188.510 ;
        RECT 72.120 188.450 72.440 188.510 ;
        RECT 73.515 188.465 73.805 188.695 ;
        RECT 73.960 188.650 74.280 188.710 ;
        RECT 75.800 188.650 76.120 188.710 ;
        RECT 73.960 188.510 76.120 188.650 ;
        RECT 53.275 188.310 53.565 188.355 ;
        RECT 54.640 188.310 54.960 188.370 ;
        RECT 51.510 188.170 54.960 188.310 ;
        RECT 50.500 188.110 50.820 188.170 ;
        RECT 53.275 188.125 53.565 188.170 ;
        RECT 54.640 188.110 54.960 188.170 ;
        RECT 56.020 188.310 56.340 188.370 ;
        RECT 57.860 188.310 58.180 188.370 ;
        RECT 56.020 188.170 58.180 188.310 ;
        RECT 56.020 188.110 56.340 188.170 ;
        RECT 57.860 188.110 58.180 188.170 ;
        RECT 63.380 188.110 63.700 188.370 ;
        RECT 71.200 188.310 71.520 188.370 ;
        RECT 73.590 188.310 73.730 188.465 ;
        RECT 73.960 188.450 74.280 188.510 ;
        RECT 75.800 188.450 76.120 188.510 ;
        RECT 83.160 188.650 83.480 188.710 ;
        RECT 83.635 188.650 83.925 188.695 ;
        RECT 83.160 188.510 83.925 188.650 ;
        RECT 83.160 188.450 83.480 188.510 ;
        RECT 83.635 188.465 83.925 188.510 ;
        RECT 84.095 188.310 84.385 188.355 ;
        RECT 71.200 188.170 84.385 188.310 ;
        RECT 71.200 188.110 71.520 188.170 ;
        RECT 84.095 188.125 84.385 188.170 ;
        RECT 46.415 187.830 49.810 187.970 ;
        RECT 51.420 187.970 51.740 188.030 ;
        RECT 68.455 187.970 68.745 188.015 ;
        RECT 51.420 187.830 68.745 187.970 ;
        RECT 46.415 187.785 46.705 187.830 ;
        RECT 47.740 187.770 48.060 187.830 ;
        RECT 51.420 187.770 51.740 187.830 ;
        RECT 68.455 187.785 68.745 187.830 ;
        RECT 35.335 187.630 35.625 187.675 ;
        RECT 33.110 187.490 35.625 187.630 ;
        RECT 31.195 187.445 31.485 187.490 ;
        RECT 31.640 187.430 31.960 187.490 ;
        RECT 35.335 187.445 35.625 187.490 ;
        RECT 39.460 187.630 39.780 187.690 ;
        RECT 40.855 187.630 41.145 187.675 ;
        RECT 39.460 187.490 41.145 187.630 ;
        RECT 39.460 187.430 39.780 187.490 ;
        RECT 40.855 187.445 41.145 187.490 ;
        RECT 43.140 187.630 43.460 187.690 ;
        RECT 45.455 187.630 45.745 187.675 ;
        RECT 43.140 187.490 45.745 187.630 ;
        RECT 43.140 187.430 43.460 187.490 ;
        RECT 45.455 187.445 45.745 187.490 ;
        RECT 50.960 187.630 51.280 187.690 ;
        RECT 59.240 187.630 59.560 187.690 ;
        RECT 50.960 187.490 59.560 187.630 ;
        RECT 50.960 187.430 51.280 187.490 ;
        RECT 59.240 187.430 59.560 187.490 ;
        RECT 60.620 187.430 60.940 187.690 ;
        RECT 62.460 187.630 62.780 187.690 ;
        RECT 71.215 187.630 71.505 187.675 ;
        RECT 62.460 187.490 71.505 187.630 ;
        RECT 62.460 187.430 62.780 187.490 ;
        RECT 71.215 187.445 71.505 187.490 ;
        RECT 72.580 187.430 72.900 187.690 ;
        RECT 77.195 187.630 77.485 187.675 ;
        RECT 82.240 187.630 82.560 187.690 ;
        RECT 77.195 187.490 82.560 187.630 ;
        RECT 77.195 187.445 77.485 187.490 ;
        RECT 82.240 187.430 82.560 187.490 ;
        RECT 15.930 186.810 87.230 187.290 ;
        RECT 18.315 186.610 18.605 186.655 ;
        RECT 19.680 186.610 20.000 186.670 ;
        RECT 27.040 186.610 27.360 186.670 ;
        RECT 18.315 186.470 20.000 186.610 ;
        RECT 18.315 186.425 18.605 186.470 ;
        RECT 19.680 186.410 20.000 186.470 ;
        RECT 21.610 186.470 27.360 186.610 ;
        RECT 21.610 186.315 21.750 186.470 ;
        RECT 27.040 186.410 27.360 186.470 ;
        RECT 29.355 186.610 29.645 186.655 ;
        RECT 29.800 186.610 30.120 186.670 ;
        RECT 29.355 186.470 30.120 186.610 ;
        RECT 29.355 186.425 29.645 186.470 ;
        RECT 29.800 186.410 30.120 186.470 ;
        RECT 30.735 186.610 31.025 186.655 ;
        RECT 31.180 186.610 31.500 186.670 ;
        RECT 30.735 186.470 31.500 186.610 ;
        RECT 30.735 186.425 31.025 186.470 ;
        RECT 31.180 186.410 31.500 186.470 ;
        RECT 33.020 186.610 33.340 186.670 ;
        RECT 35.320 186.610 35.640 186.670 ;
        RECT 33.020 186.470 35.640 186.610 ;
        RECT 33.020 186.410 33.340 186.470 ;
        RECT 35.320 186.410 35.640 186.470 ;
        RECT 35.780 186.410 36.100 186.670 ;
        RECT 36.715 186.610 37.005 186.655 ;
        RECT 38.080 186.610 38.400 186.670 ;
        RECT 36.715 186.470 38.400 186.610 ;
        RECT 36.715 186.425 37.005 186.470 ;
        RECT 38.080 186.410 38.400 186.470 ;
        RECT 41.300 186.410 41.620 186.670 ;
        RECT 47.295 186.610 47.585 186.655 ;
        RECT 48.200 186.610 48.520 186.670 ;
        RECT 43.690 186.470 47.050 186.610 ;
        RECT 21.535 186.085 21.825 186.315 ;
        RECT 21.980 186.070 22.300 186.330 ;
        RECT 24.295 186.270 24.585 186.315 ;
        RECT 25.200 186.270 25.520 186.330 ;
        RECT 24.295 186.130 25.520 186.270 ;
        RECT 24.295 186.085 24.585 186.130 ;
        RECT 25.200 186.070 25.520 186.130 ;
        RECT 25.660 186.270 25.980 186.330 ;
        RECT 28.880 186.270 29.200 186.330 ;
        RECT 25.660 186.130 28.650 186.270 ;
        RECT 25.660 186.070 25.980 186.130 ;
        RECT 19.695 185.930 19.985 185.975 ;
        RECT 19.695 185.790 21.290 185.930 ;
        RECT 19.695 185.745 19.985 185.790 ;
        RECT 17.380 185.390 17.700 185.650 ;
        RECT 19.235 185.405 19.525 185.635 ;
        RECT 20.155 185.590 20.445 185.635 ;
        RECT 20.600 185.590 20.920 185.650 ;
        RECT 21.150 185.635 21.290 185.790 ;
        RECT 23.360 185.730 23.680 185.990 ;
        RECT 26.120 185.930 26.440 185.990 ;
        RECT 27.515 185.930 27.805 185.975 ;
        RECT 26.120 185.790 27.805 185.930 ;
        RECT 28.510 185.930 28.650 186.130 ;
        RECT 28.880 186.130 37.850 186.270 ;
        RECT 28.880 186.070 29.200 186.130 ;
        RECT 33.955 185.930 34.245 185.975 ;
        RECT 37.160 185.930 37.480 185.990 ;
        RECT 28.510 185.790 33.710 185.930 ;
        RECT 26.120 185.730 26.440 185.790 ;
        RECT 27.515 185.745 27.805 185.790 ;
        RECT 20.155 185.450 20.920 185.590 ;
        RECT 20.155 185.405 20.445 185.450 ;
        RECT 19.310 185.250 19.450 185.405 ;
        RECT 20.600 185.390 20.920 185.450 ;
        RECT 21.075 185.405 21.365 185.635 ;
        RECT 22.440 185.390 22.760 185.650 ;
        RECT 23.450 185.590 23.590 185.730 ;
        RECT 24.920 185.590 25.210 185.635 ;
        RECT 23.450 185.450 25.210 185.590 ;
        RECT 24.920 185.405 25.210 185.450 ;
        RECT 27.055 185.590 27.345 185.635 ;
        RECT 29.800 185.590 30.120 185.650 ;
        RECT 27.055 185.450 30.120 185.590 ;
        RECT 27.055 185.405 27.345 185.450 ;
        RECT 29.800 185.390 30.120 185.450 ;
        RECT 30.275 185.590 30.565 185.635 ;
        RECT 32.100 185.590 32.420 185.650 ;
        RECT 30.275 185.450 32.420 185.590 ;
        RECT 33.570 185.590 33.710 185.790 ;
        RECT 33.955 185.790 37.480 185.930 ;
        RECT 33.955 185.745 34.245 185.790 ;
        RECT 37.160 185.730 37.480 185.790 ;
        RECT 37.710 185.715 37.850 186.130 ;
        RECT 42.220 186.070 42.540 186.330 ;
        RECT 34.875 185.590 35.165 185.635 ;
        RECT 35.780 185.590 36.100 185.650 ;
        RECT 33.570 185.450 34.700 185.590 ;
        RECT 30.275 185.405 30.565 185.450 ;
        RECT 32.100 185.390 32.420 185.450 ;
        RECT 21.980 185.250 22.300 185.310 ;
        RECT 19.310 185.110 22.300 185.250 ;
        RECT 21.980 185.050 22.300 185.110 ;
        RECT 23.375 185.250 23.665 185.295 ;
        RECT 32.575 185.250 32.865 185.295 ;
        RECT 33.480 185.250 33.800 185.310 ;
        RECT 23.375 185.110 28.190 185.250 ;
        RECT 23.375 185.065 23.665 185.110 ;
        RECT 23.820 184.910 24.140 184.970 ;
        RECT 25.215 184.910 25.505 184.955 ;
        RECT 23.820 184.770 25.505 184.910 ;
        RECT 23.820 184.710 24.140 184.770 ;
        RECT 25.215 184.725 25.505 184.770 ;
        RECT 26.120 184.910 26.440 184.970 ;
        RECT 27.500 184.910 27.820 184.970 ;
        RECT 26.120 184.770 27.820 184.910 ;
        RECT 28.050 184.910 28.190 185.110 ;
        RECT 32.575 185.110 33.800 185.250 ;
        RECT 34.560 185.250 34.700 185.450 ;
        RECT 34.875 185.450 36.100 185.590 ;
        RECT 37.635 185.485 37.925 185.715 ;
        RECT 34.875 185.405 35.165 185.450 ;
        RECT 35.780 185.390 36.100 185.450 ;
        RECT 39.000 185.390 39.320 185.650 ;
        RECT 39.460 185.390 39.780 185.650 ;
        RECT 40.395 185.590 40.685 185.635 ;
        RECT 40.840 185.590 41.160 185.650 ;
        RECT 40.395 185.450 41.160 185.590 ;
        RECT 40.395 185.405 40.685 185.450 ;
        RECT 40.840 185.390 41.160 185.450 ;
        RECT 43.155 185.590 43.445 185.635 ;
        RECT 43.690 185.590 43.830 186.470 ;
        RECT 44.060 186.270 44.380 186.330 ;
        RECT 46.910 186.270 47.050 186.470 ;
        RECT 47.295 186.470 48.520 186.610 ;
        RECT 47.295 186.425 47.585 186.470 ;
        RECT 48.200 186.410 48.520 186.470 ;
        RECT 51.895 186.610 52.185 186.655 ;
        RECT 52.800 186.610 53.120 186.670 ;
        RECT 51.895 186.470 53.120 186.610 ;
        RECT 51.895 186.425 52.185 186.470 ;
        RECT 52.800 186.410 53.120 186.470 ;
        RECT 53.735 186.610 54.025 186.655 ;
        RECT 54.640 186.610 54.960 186.670 ;
        RECT 63.380 186.610 63.700 186.670 ;
        RECT 53.735 186.470 63.700 186.610 ;
        RECT 53.735 186.425 54.025 186.470 ;
        RECT 54.640 186.410 54.960 186.470 ;
        RECT 63.380 186.410 63.700 186.470 ;
        RECT 65.220 186.610 65.540 186.670 ;
        RECT 70.740 186.610 71.060 186.670 ;
        RECT 65.220 186.470 67.750 186.610 ;
        RECT 65.220 186.410 65.540 186.470 ;
        RECT 47.740 186.270 48.060 186.330 ;
        RECT 50.500 186.270 50.820 186.330 ;
        RECT 57.400 186.270 57.720 186.330 ;
        RECT 67.610 186.270 67.750 186.470 ;
        RECT 70.740 186.470 78.330 186.610 ;
        RECT 70.740 186.410 71.060 186.470 ;
        RECT 73.040 186.270 73.360 186.330 ;
        RECT 77.640 186.270 77.960 186.330 ;
        RECT 44.060 186.130 46.130 186.270 ;
        RECT 46.910 186.130 48.060 186.270 ;
        RECT 44.060 186.070 44.380 186.130 ;
        RECT 45.440 185.635 45.760 185.660 ;
        RECT 45.990 185.635 46.130 186.130 ;
        RECT 47.740 186.070 48.060 186.130 ;
        RECT 49.195 186.130 50.820 186.270 ;
        RECT 49.195 185.930 49.335 186.130 ;
        RECT 50.500 186.070 50.820 186.130 ;
        RECT 51.970 186.130 57.170 186.270 ;
        RECT 47.370 185.790 49.335 185.930 ;
        RECT 43.155 185.450 43.830 185.590 ;
        RECT 43.155 185.405 43.445 185.450 ;
        RECT 44.075 185.405 44.365 185.635 ;
        RECT 44.535 185.405 44.825 185.635 ;
        RECT 45.175 185.405 45.760 185.635 ;
        RECT 45.915 185.405 46.205 185.635 ;
        RECT 44.150 185.250 44.290 185.405 ;
        RECT 34.560 185.110 44.290 185.250 ;
        RECT 44.610 185.250 44.750 185.405 ;
        RECT 45.440 185.400 45.760 185.405 ;
        RECT 47.370 185.250 47.510 185.790 ;
        RECT 48.200 185.390 48.520 185.650 ;
        RECT 48.675 185.405 48.965 185.635 ;
        RECT 49.195 185.590 49.335 185.790 ;
        RECT 49.580 185.730 49.900 185.990 ;
        RECT 50.055 185.590 50.345 185.635 ;
        RECT 49.195 185.450 50.345 185.590 ;
        RECT 50.055 185.405 50.345 185.450 ;
        RECT 44.610 185.110 47.510 185.250 ;
        RECT 47.740 185.250 48.060 185.310 ;
        RECT 48.750 185.250 48.890 185.405 ;
        RECT 50.500 185.390 50.820 185.650 ;
        RECT 50.960 185.390 51.280 185.650 ;
        RECT 51.970 185.635 52.110 186.130 ;
        RECT 52.340 185.930 52.660 185.990 ;
        RECT 57.030 185.930 57.170 186.130 ;
        RECT 57.400 186.130 67.290 186.270 ;
        RECT 67.610 186.130 77.960 186.270 ;
        RECT 57.400 186.070 57.720 186.130 ;
        RECT 63.840 185.930 64.160 185.990 ;
        RECT 52.340 185.790 53.030 185.930 ;
        RECT 57.030 185.790 64.160 185.930 ;
        RECT 52.340 185.730 52.660 185.790 ;
        RECT 52.890 185.635 53.030 185.790 ;
        RECT 63.840 185.730 64.160 185.790 ;
        RECT 51.895 185.405 52.185 185.635 ;
        RECT 52.815 185.405 53.105 185.635 ;
        RECT 54.195 185.590 54.485 185.635 ;
        RECT 58.780 185.590 59.100 185.650 ;
        RECT 54.195 185.450 59.100 185.590 ;
        RECT 54.195 185.405 54.485 185.450 ;
        RECT 58.780 185.390 59.100 185.450 ;
        RECT 65.680 185.590 66.000 185.650 ;
        RECT 67.150 185.635 67.290 186.130 ;
        RECT 73.040 186.070 73.360 186.130 ;
        RECT 77.640 186.070 77.960 186.130 ;
        RECT 75.340 185.930 75.660 185.990 ;
        RECT 78.190 185.930 78.330 186.470 ;
        RECT 83.160 186.410 83.480 186.670 ;
        RECT 75.340 185.790 77.410 185.930 ;
        RECT 78.190 185.790 84.310 185.930 ;
        RECT 75.340 185.730 75.660 185.790 ;
        RECT 66.155 185.590 66.445 185.635 ;
        RECT 65.680 185.450 66.445 185.590 ;
        RECT 65.680 185.390 66.000 185.450 ;
        RECT 66.155 185.405 66.445 185.450 ;
        RECT 67.075 185.405 67.365 185.635 ;
        RECT 72.580 185.590 72.900 185.650 ;
        RECT 77.270 185.635 77.410 185.790 ;
        RECT 72.440 185.390 72.900 185.590 ;
        RECT 76.275 185.405 76.565 185.635 ;
        RECT 77.195 185.405 77.485 185.635 ;
        RECT 63.855 185.250 64.145 185.295 ;
        RECT 72.440 185.250 72.580 185.390 ;
        RECT 47.740 185.110 63.610 185.250 ;
        RECT 32.575 185.065 32.865 185.110 ;
        RECT 33.480 185.050 33.800 185.110 ;
        RECT 30.260 184.910 30.580 184.970 ;
        RECT 28.050 184.770 30.580 184.910 ;
        RECT 26.120 184.710 26.440 184.770 ;
        RECT 27.500 184.710 27.820 184.770 ;
        RECT 30.260 184.710 30.580 184.770 ;
        RECT 33.035 184.910 33.325 184.955 ;
        RECT 34.400 184.910 34.720 184.970 ;
        RECT 33.035 184.770 34.720 184.910 ;
        RECT 33.035 184.725 33.325 184.770 ;
        RECT 34.400 184.710 34.720 184.770 ;
        RECT 34.860 184.910 35.180 184.970 ;
        RECT 37.620 184.910 37.940 184.970 ;
        RECT 34.860 184.770 37.940 184.910 ;
        RECT 34.860 184.710 35.180 184.770 ;
        RECT 37.620 184.710 37.940 184.770 ;
        RECT 41.760 184.910 42.080 184.970 ;
        RECT 44.610 184.910 44.750 185.110 ;
        RECT 47.740 185.050 48.060 185.110 ;
        RECT 41.760 184.770 44.750 184.910 ;
        RECT 51.420 184.910 51.740 184.970 ;
        RECT 53.720 184.910 54.040 184.970 ;
        RECT 51.420 184.770 54.040 184.910 ;
        RECT 41.760 184.710 42.080 184.770 ;
        RECT 51.420 184.710 51.740 184.770 ;
        RECT 53.720 184.710 54.040 184.770 ;
        RECT 56.940 184.910 57.260 184.970 ;
        RECT 62.000 184.910 62.320 184.970 ;
        RECT 56.940 184.770 62.320 184.910 ;
        RECT 63.470 184.910 63.610 185.110 ;
        RECT 63.855 185.110 72.580 185.250 ;
        RECT 76.350 185.250 76.490 185.405 ;
        RECT 77.640 185.390 77.960 185.650 ;
        RECT 78.100 185.390 78.420 185.650 ;
        RECT 80.860 185.590 81.180 185.650 ;
        RECT 84.170 185.635 84.310 185.790 ;
        RECT 81.335 185.590 81.625 185.635 ;
        RECT 80.860 185.450 81.625 185.590 ;
        RECT 80.860 185.390 81.180 185.450 ;
        RECT 81.335 185.405 81.625 185.450 ;
        RECT 83.635 185.405 83.925 185.635 ;
        RECT 84.095 185.405 84.385 185.635 ;
        RECT 79.495 185.250 79.785 185.295 ;
        RECT 83.160 185.250 83.480 185.310 ;
        RECT 76.350 185.110 78.330 185.250 ;
        RECT 63.855 185.065 64.145 185.110 ;
        RECT 78.190 184.970 78.330 185.110 ;
        RECT 79.495 185.110 83.480 185.250 ;
        RECT 83.710 185.250 83.850 185.405 ;
        RECT 85.000 185.390 85.320 185.650 ;
        RECT 86.380 185.250 86.700 185.310 ;
        RECT 87.300 185.250 87.620 185.310 ;
        RECT 83.710 185.110 87.620 185.250 ;
        RECT 79.495 185.065 79.785 185.110 ;
        RECT 83.160 185.050 83.480 185.110 ;
        RECT 86.380 185.050 86.700 185.110 ;
        RECT 87.300 185.050 87.620 185.110 ;
        RECT 68.440 184.910 68.760 184.970 ;
        RECT 63.470 184.770 68.760 184.910 ;
        RECT 56.940 184.710 57.260 184.770 ;
        RECT 62.000 184.710 62.320 184.770 ;
        RECT 68.440 184.710 68.760 184.770 ;
        RECT 73.960 184.910 74.280 184.970 ;
        RECT 74.435 184.910 74.725 184.955 ;
        RECT 73.960 184.770 74.725 184.910 ;
        RECT 73.960 184.710 74.280 184.770 ;
        RECT 74.435 184.725 74.725 184.770 ;
        RECT 78.100 184.710 78.420 184.970 ;
        RECT 79.020 184.910 79.340 184.970 ;
        RECT 81.780 184.910 82.100 184.970 ;
        RECT 84.555 184.910 84.845 184.955 ;
        RECT 79.020 184.770 84.845 184.910 ;
        RECT 79.020 184.710 79.340 184.770 ;
        RECT 81.780 184.710 82.100 184.770 ;
        RECT 84.555 184.725 84.845 184.770 ;
        RECT 15.930 184.090 87.230 184.570 ;
        RECT 16.460 183.890 16.780 183.950 ;
        RECT 19.695 183.890 19.985 183.935 ;
        RECT 16.460 183.750 19.985 183.890 ;
        RECT 16.460 183.690 16.780 183.750 ;
        RECT 19.695 183.705 19.985 183.750 ;
        RECT 22.440 183.890 22.760 183.950 ;
        RECT 23.375 183.890 23.665 183.935 ;
        RECT 22.440 183.750 23.665 183.890 ;
        RECT 22.440 183.690 22.760 183.750 ;
        RECT 23.375 183.705 23.665 183.750 ;
        RECT 24.295 183.890 24.585 183.935 ;
        RECT 25.660 183.890 25.980 183.950 ;
        RECT 24.295 183.750 25.980 183.890 ;
        RECT 24.295 183.705 24.585 183.750 ;
        RECT 25.660 183.690 25.980 183.750 ;
        RECT 26.595 183.705 26.885 183.935 ;
        RECT 18.760 183.550 19.080 183.610 ;
        RECT 21.535 183.550 21.825 183.595 ;
        RECT 18.760 183.410 21.825 183.550 ;
        RECT 26.670 183.550 26.810 183.705 ;
        RECT 27.960 183.690 28.280 183.950 ;
        RECT 28.420 183.890 28.740 183.950 ;
        RECT 28.895 183.890 29.185 183.935 ;
        RECT 28.420 183.750 29.185 183.890 ;
        RECT 28.420 183.690 28.740 183.750 ;
        RECT 28.895 183.705 29.185 183.750 ;
        RECT 33.020 183.690 33.340 183.950 ;
        RECT 33.940 183.890 34.260 183.950 ;
        RECT 34.860 183.890 35.180 183.950 ;
        RECT 33.940 183.750 35.180 183.890 ;
        RECT 33.940 183.690 34.260 183.750 ;
        RECT 34.860 183.690 35.180 183.750 ;
        RECT 39.000 183.890 39.320 183.950 ;
        RECT 42.235 183.890 42.525 183.935 ;
        RECT 39.000 183.750 42.525 183.890 ;
        RECT 39.000 183.690 39.320 183.750 ;
        RECT 42.235 183.705 42.525 183.750 ;
        RECT 44.980 183.690 45.300 183.950 ;
        RECT 45.900 183.890 46.220 183.950 ;
        RECT 46.375 183.890 46.665 183.935 ;
        RECT 45.900 183.750 46.665 183.890 ;
        RECT 45.900 183.690 46.220 183.750 ;
        RECT 46.375 183.705 46.665 183.750 ;
        RECT 48.675 183.890 48.965 183.935 ;
        RECT 51.880 183.890 52.200 183.950 ;
        RECT 48.675 183.750 52.200 183.890 ;
        RECT 48.675 183.705 48.965 183.750 ;
        RECT 51.880 183.690 52.200 183.750 ;
        RECT 57.860 183.890 58.180 183.950 ;
        RECT 58.780 183.890 59.100 183.950 ;
        RECT 57.860 183.750 59.100 183.890 ;
        RECT 57.860 183.690 58.180 183.750 ;
        RECT 58.780 183.690 59.100 183.750 ;
        RECT 59.240 183.690 59.560 183.950 ;
        RECT 60.160 183.890 60.480 183.950 ;
        RECT 61.540 183.890 61.860 183.950 ;
        RECT 63.395 183.890 63.685 183.935 ;
        RECT 60.160 183.750 60.850 183.890 ;
        RECT 60.160 183.690 60.480 183.750 ;
        RECT 29.340 183.550 29.660 183.610 ;
        RECT 26.670 183.410 29.660 183.550 ;
        RECT 18.760 183.350 19.080 183.410 ;
        RECT 21.535 183.365 21.825 183.410 ;
        RECT 29.340 183.350 29.660 183.410 ;
        RECT 31.640 183.550 31.960 183.610 ;
        RECT 43.140 183.550 43.460 183.610 ;
        RECT 52.815 183.550 53.105 183.595 ;
        RECT 54.640 183.550 54.960 183.610 ;
        RECT 59.330 183.550 59.470 183.690 ;
        RECT 60.710 183.595 60.850 183.750 ;
        RECT 61.540 183.750 63.685 183.890 ;
        RECT 61.540 183.690 61.860 183.750 ;
        RECT 63.395 183.705 63.685 183.750 ;
        RECT 66.140 183.890 66.460 183.950 ;
        RECT 66.615 183.890 66.905 183.935 ;
        RECT 66.140 183.750 66.905 183.890 ;
        RECT 66.140 183.690 66.460 183.750 ;
        RECT 66.615 183.705 66.905 183.750 ;
        RECT 71.660 183.890 71.980 183.950 ;
        RECT 76.275 183.890 76.565 183.935 ;
        RECT 85.000 183.890 85.320 183.950 ;
        RECT 71.660 183.750 85.320 183.890 ;
        RECT 71.660 183.690 71.980 183.750 ;
        RECT 76.275 183.705 76.565 183.750 ;
        RECT 85.000 183.690 85.320 183.750 ;
        RECT 31.640 183.410 43.460 183.550 ;
        RECT 31.640 183.350 31.960 183.410 ;
        RECT 43.140 183.350 43.460 183.410 ;
        RECT 44.150 183.410 52.110 183.550 ;
        RECT 16.000 183.210 16.320 183.270 ;
        RECT 19.235 183.210 19.525 183.255 ;
        RECT 16.000 183.070 19.525 183.210 ;
        RECT 16.000 183.010 16.320 183.070 ;
        RECT 19.235 183.025 19.525 183.070 ;
        RECT 20.600 183.010 20.920 183.270 ;
        RECT 22.900 183.010 23.220 183.270 ;
        RECT 23.820 183.010 24.140 183.270 ;
        RECT 24.740 183.210 25.060 183.270 ;
        RECT 25.215 183.210 25.505 183.255 ;
        RECT 24.740 183.070 25.505 183.210 ;
        RECT 24.740 183.010 25.060 183.070 ;
        RECT 25.215 183.025 25.505 183.070 ;
        RECT 25.660 183.010 25.980 183.270 ;
        RECT 27.040 183.010 27.360 183.270 ;
        RECT 28.435 183.025 28.725 183.255 ;
        RECT 19.680 182.870 20.000 182.930 ;
        RECT 28.510 182.870 28.650 183.025 ;
        RECT 30.720 183.010 31.040 183.270 ;
        RECT 32.115 183.025 32.405 183.255 ;
        RECT 33.035 183.210 33.325 183.255 ;
        RECT 38.540 183.210 38.860 183.270 ;
        RECT 33.035 183.070 38.860 183.210 ;
        RECT 33.035 183.025 33.325 183.070 ;
        RECT 19.680 182.730 28.650 182.870 ;
        RECT 32.190 182.870 32.330 183.025 ;
        RECT 38.540 183.010 38.860 183.070 ;
        RECT 41.760 183.210 42.080 183.270 ;
        RECT 44.150 183.210 44.290 183.410 ;
        RECT 51.970 183.270 52.110 183.410 ;
        RECT 52.815 183.410 56.250 183.550 ;
        RECT 52.815 183.365 53.105 183.410 ;
        RECT 54.640 183.350 54.960 183.410 ;
        RECT 41.760 183.070 44.290 183.210 ;
        RECT 41.760 183.010 42.080 183.070 ;
        RECT 44.520 183.010 44.840 183.270 ;
        RECT 45.915 183.210 46.205 183.255 ;
        RECT 46.360 183.210 46.680 183.270 ;
        RECT 45.915 183.070 46.680 183.210 ;
        RECT 45.915 183.025 46.205 183.070 ;
        RECT 46.360 183.010 46.680 183.070 ;
        RECT 47.280 183.010 47.600 183.270 ;
        RECT 47.755 183.025 48.045 183.255 ;
        RECT 50.055 183.210 50.345 183.255 ;
        RECT 50.960 183.210 51.280 183.270 ;
        RECT 50.055 183.070 51.280 183.210 ;
        RECT 50.055 183.025 50.345 183.070 ;
        RECT 33.940 182.870 34.260 182.930 ;
        RECT 42.695 182.870 42.985 182.915 ;
        RECT 32.190 182.730 42.985 182.870 ;
        RECT 19.680 182.670 20.000 182.730 ;
        RECT 33.940 182.670 34.260 182.730 ;
        RECT 42.695 182.685 42.985 182.730 ;
        RECT 43.155 182.685 43.445 182.915 ;
        RECT 47.830 182.870 47.970 183.025 ;
        RECT 50.960 183.010 51.280 183.070 ;
        RECT 51.420 183.010 51.740 183.270 ;
        RECT 51.880 183.010 52.200 183.270 ;
        RECT 52.340 183.210 52.660 183.270 ;
        RECT 53.275 183.210 53.565 183.255 ;
        RECT 52.340 183.070 53.565 183.210 ;
        RECT 52.340 183.010 52.660 183.070 ;
        RECT 53.275 183.025 53.565 183.070 ;
        RECT 53.720 183.010 54.040 183.270 ;
        RECT 56.110 183.255 56.250 183.410 ;
        RECT 56.570 183.410 59.470 183.550 ;
        RECT 56.035 183.025 56.325 183.255 ;
        RECT 50.500 182.870 50.820 182.930 ;
        RECT 55.115 182.870 55.405 182.915 ;
        RECT 47.830 182.730 50.270 182.870 ;
        RECT 16.920 182.530 17.240 182.590 ;
        RECT 29.815 182.530 30.105 182.575 ;
        RECT 16.920 182.390 30.105 182.530 ;
        RECT 16.920 182.330 17.240 182.390 ;
        RECT 29.815 182.345 30.105 182.390 ;
        RECT 30.260 182.530 30.580 182.590 ;
        RECT 41.760 182.530 42.080 182.590 ;
        RECT 43.230 182.530 43.370 182.685 ;
        RECT 30.260 182.390 42.080 182.530 ;
        RECT 30.260 182.330 30.580 182.390 ;
        RECT 41.760 182.330 42.080 182.390 ;
        RECT 42.310 182.390 43.370 182.530 ;
        RECT 43.600 182.530 43.920 182.590 ;
        RECT 49.135 182.530 49.425 182.575 ;
        RECT 43.600 182.390 49.425 182.530 ;
        RECT 50.130 182.530 50.270 182.730 ;
        RECT 50.500 182.730 55.405 182.870 ;
        RECT 50.500 182.670 50.820 182.730 ;
        RECT 55.115 182.685 55.405 182.730 ;
        RECT 56.570 182.530 56.710 183.410 ;
        RECT 60.635 183.365 60.925 183.595 ;
        RECT 72.580 183.550 72.900 183.610 ;
        RECT 82.240 183.550 82.560 183.610 ;
        RECT 85.475 183.550 85.765 183.595 ;
        RECT 72.580 183.410 74.650 183.550 ;
        RECT 72.580 183.350 72.900 183.410 ;
        RECT 57.875 183.025 58.165 183.255 ;
        RECT 58.795 183.210 59.085 183.255 ;
        RECT 59.240 183.210 59.560 183.270 ;
        RECT 58.795 183.070 59.560 183.210 ;
        RECT 58.795 183.025 59.085 183.070 ;
        RECT 56.955 182.685 57.245 182.915 ;
        RECT 50.130 182.390 56.710 182.530 ;
        RECT 57.030 182.530 57.170 182.685 ;
        RECT 57.400 182.670 57.720 182.930 ;
        RECT 57.950 182.870 58.090 183.025 ;
        RECT 59.240 183.010 59.560 183.070 ;
        RECT 60.175 183.025 60.465 183.255 ;
        RECT 61.095 183.210 61.385 183.255 ;
        RECT 61.540 183.210 61.860 183.270 ;
        RECT 61.095 183.070 61.860 183.210 ;
        RECT 61.095 183.025 61.385 183.070 ;
        RECT 59.700 182.870 60.020 182.930 ;
        RECT 57.950 182.730 60.020 182.870 ;
        RECT 60.250 182.870 60.390 183.025 ;
        RECT 61.540 183.010 61.860 183.070 ;
        RECT 62.015 183.210 62.305 183.255 ;
        RECT 62.460 183.210 62.780 183.270 ;
        RECT 62.015 183.070 62.780 183.210 ;
        RECT 62.015 183.025 62.305 183.070 ;
        RECT 62.460 183.010 62.780 183.070 ;
        RECT 63.380 183.210 63.700 183.270 ;
        RECT 64.775 183.210 65.065 183.255 ;
        RECT 63.380 183.070 65.065 183.210 ;
        RECT 63.380 183.010 63.700 183.070 ;
        RECT 64.775 183.025 65.065 183.070 ;
        RECT 73.960 183.010 74.280 183.270 ;
        RECT 74.510 183.255 74.650 183.410 ;
        RECT 82.240 183.410 85.765 183.550 ;
        RECT 82.240 183.350 82.560 183.410 ;
        RECT 85.475 183.365 85.765 183.410 ;
        RECT 74.435 183.025 74.725 183.255 ;
        RECT 74.880 183.010 75.200 183.270 ;
        RECT 60.250 182.730 63.150 182.870 ;
        RECT 59.700 182.670 60.020 182.730 ;
        RECT 59.790 182.530 59.930 182.670 ;
        RECT 63.010 182.590 63.150 182.730 ;
        RECT 64.315 182.685 64.605 182.915 ;
        RECT 74.050 182.870 74.190 183.010 ;
        RECT 84.080 182.870 84.400 182.930 ;
        RECT 74.050 182.730 84.400 182.870 ;
        RECT 62.460 182.530 62.780 182.590 ;
        RECT 57.030 182.390 58.230 182.530 ;
        RECT 59.790 182.390 62.780 182.530 ;
        RECT 42.310 182.250 42.450 182.390 ;
        RECT 43.600 182.330 43.920 182.390 ;
        RECT 49.135 182.345 49.425 182.390 ;
        RECT 18.300 181.990 18.620 182.250 ;
        RECT 21.995 182.190 22.285 182.235 ;
        RECT 22.900 182.190 23.220 182.250 ;
        RECT 24.280 182.190 24.600 182.250 ;
        RECT 21.995 182.050 24.600 182.190 ;
        RECT 21.995 182.005 22.285 182.050 ;
        RECT 22.900 181.990 23.220 182.050 ;
        RECT 24.280 181.990 24.600 182.050 ;
        RECT 27.040 182.190 27.360 182.250 ;
        RECT 42.220 182.190 42.540 182.250 ;
        RECT 27.040 182.050 42.540 182.190 ;
        RECT 27.040 181.990 27.360 182.050 ;
        RECT 42.220 181.990 42.540 182.050 ;
        RECT 42.680 182.190 43.000 182.250 ;
        RECT 44.075 182.190 44.365 182.235 ;
        RECT 42.680 182.050 44.365 182.190 ;
        RECT 42.680 181.990 43.000 182.050 ;
        RECT 44.075 182.005 44.365 182.050 ;
        RECT 48.200 182.190 48.520 182.250 ;
        RECT 50.500 182.190 50.820 182.250 ;
        RECT 48.200 182.050 50.820 182.190 ;
        RECT 48.200 181.990 48.520 182.050 ;
        RECT 50.500 181.990 50.820 182.050 ;
        RECT 53.720 182.190 54.040 182.250 ;
        RECT 54.655 182.190 54.945 182.235 ;
        RECT 53.720 182.050 54.945 182.190 ;
        RECT 58.090 182.190 58.230 182.390 ;
        RECT 62.460 182.330 62.780 182.390 ;
        RECT 62.920 182.330 63.240 182.590 ;
        RECT 64.390 182.530 64.530 182.685 ;
        RECT 84.080 182.670 84.400 182.730 ;
        RECT 67.060 182.530 67.380 182.590 ;
        RECT 79.020 182.530 79.340 182.590 ;
        RECT 64.390 182.390 67.380 182.530 ;
        RECT 67.060 182.330 67.380 182.390 ;
        RECT 72.440 182.390 79.340 182.530 ;
        RECT 58.780 182.190 59.100 182.250 ;
        RECT 58.090 182.050 59.100 182.190 ;
        RECT 53.720 181.990 54.040 182.050 ;
        RECT 54.655 182.005 54.945 182.050 ;
        RECT 58.780 181.990 59.100 182.050 ;
        RECT 59.255 182.190 59.545 182.235 ;
        RECT 59.700 182.190 60.020 182.250 ;
        RECT 59.255 182.050 60.020 182.190 ;
        RECT 59.255 182.005 59.545 182.050 ;
        RECT 59.700 181.990 60.020 182.050 ;
        RECT 64.760 182.190 65.080 182.250 ;
        RECT 72.440 182.190 72.580 182.390 ;
        RECT 79.020 182.330 79.340 182.390 ;
        RECT 64.760 182.050 72.580 182.190 ;
        RECT 64.760 181.990 65.080 182.050 ;
        RECT 78.100 181.990 78.420 182.250 ;
        RECT 15.930 181.370 87.230 181.850 ;
        RECT 21.060 180.970 21.380 181.230 ;
        RECT 24.740 181.170 25.060 181.230 ;
        RECT 27.040 181.170 27.360 181.230 ;
        RECT 24.740 181.030 27.360 181.170 ;
        RECT 24.740 180.970 25.060 181.030 ;
        RECT 27.040 180.970 27.360 181.030 ;
        RECT 28.435 181.170 28.725 181.215 ;
        RECT 30.720 181.170 31.040 181.230 ;
        RECT 39.015 181.170 39.305 181.215 ;
        RECT 28.435 181.030 31.040 181.170 ;
        RECT 28.435 180.985 28.725 181.030 ;
        RECT 30.720 180.970 31.040 181.030 ;
        RECT 32.650 181.030 39.305 181.170 ;
        RECT 21.995 180.830 22.285 180.875 ;
        RECT 24.280 180.830 24.600 180.890 ;
        RECT 25.200 180.830 25.520 180.890 ;
        RECT 21.995 180.690 23.170 180.830 ;
        RECT 21.995 180.645 22.285 180.690 ;
        RECT 19.235 180.150 19.525 180.195 ;
        RECT 20.140 180.150 20.460 180.210 ;
        RECT 19.235 180.010 20.460 180.150 ;
        RECT 23.030 180.150 23.170 180.690 ;
        RECT 24.140 180.690 25.520 180.830 ;
        RECT 24.140 180.630 24.600 180.690 ;
        RECT 25.200 180.630 25.520 180.690 ;
        RECT 26.120 180.630 26.440 180.890 ;
        RECT 23.375 180.490 23.665 180.535 ;
        RECT 24.140 180.490 24.280 180.630 ;
        RECT 23.375 180.350 24.280 180.490 ;
        RECT 24.740 180.490 25.060 180.550 ;
        RECT 28.420 180.490 28.740 180.550 ;
        RECT 32.650 180.535 32.790 181.030 ;
        RECT 39.015 180.985 39.305 181.030 ;
        RECT 42.680 180.970 43.000 181.230 ;
        RECT 47.740 180.970 48.060 181.230 ;
        RECT 52.340 181.170 52.660 181.230 ;
        RECT 53.735 181.170 54.025 181.215 ;
        RECT 49.215 181.030 54.025 181.170 ;
        RECT 34.400 180.630 34.720 180.890 ;
        RECT 35.335 180.830 35.625 180.875 ;
        RECT 41.760 180.830 42.080 180.890 ;
        RECT 49.215 180.830 49.355 181.030 ;
        RECT 52.340 180.970 52.660 181.030 ;
        RECT 53.735 180.985 54.025 181.030 ;
        RECT 56.020 181.170 56.340 181.230 ;
        RECT 62.000 181.170 62.320 181.230 ;
        RECT 62.935 181.170 63.225 181.215 ;
        RECT 56.020 181.030 60.850 181.170 ;
        RECT 35.335 180.690 42.080 180.830 ;
        RECT 35.335 180.645 35.625 180.690 ;
        RECT 41.760 180.630 42.080 180.690 ;
        RECT 42.310 180.690 49.355 180.830 ;
        RECT 42.310 180.535 42.450 180.690 ;
        RECT 49.595 180.645 49.885 180.875 ;
        RECT 52.815 180.830 53.105 180.875 ;
        RECT 51.970 180.690 53.105 180.830 ;
        RECT 24.740 180.350 28.740 180.490 ;
        RECT 23.375 180.305 23.665 180.350 ;
        RECT 24.740 180.290 25.060 180.350 ;
        RECT 28.420 180.290 28.740 180.350 ;
        RECT 30.275 180.305 30.565 180.535 ;
        RECT 32.575 180.305 32.865 180.535 ;
        RECT 34.875 180.490 35.165 180.535 ;
        RECT 42.235 180.490 42.525 180.535 ;
        RECT 34.875 180.350 42.525 180.490 ;
        RECT 34.875 180.305 35.165 180.350 ;
        RECT 42.235 180.305 42.525 180.350 ;
        RECT 43.140 180.490 43.460 180.550 ;
        RECT 45.455 180.490 45.745 180.535 ;
        RECT 45.900 180.490 46.220 180.550 ;
        RECT 43.140 180.350 46.220 180.490 ;
        RECT 23.820 180.150 24.140 180.210 ;
        RECT 23.030 180.010 24.140 180.150 ;
        RECT 19.235 179.965 19.525 180.010 ;
        RECT 20.140 179.950 20.460 180.010 ;
        RECT 23.820 179.950 24.140 180.010 ;
        RECT 27.055 180.150 27.345 180.195 ;
        RECT 30.350 180.150 30.490 180.305 ;
        RECT 43.140 180.290 43.460 180.350 ;
        RECT 45.455 180.305 45.745 180.350 ;
        RECT 45.900 180.290 46.220 180.350 ;
        RECT 46.835 180.490 47.125 180.535 ;
        RECT 49.120 180.490 49.440 180.550 ;
        RECT 49.670 180.490 49.810 180.645 ;
        RECT 51.435 180.490 51.725 180.535 ;
        RECT 46.835 180.350 48.890 180.490 ;
        RECT 46.835 180.305 47.125 180.350 ;
        RECT 27.055 180.010 30.490 180.150 ;
        RECT 27.055 179.965 27.345 180.010 ;
        RECT 31.180 179.950 31.500 180.210 ;
        RECT 31.640 179.950 31.960 180.210 ;
        RECT 32.100 179.950 32.420 180.210 ;
        RECT 33.495 179.965 33.785 180.195 ;
        RECT 33.955 180.150 34.245 180.195 ;
        RECT 35.320 180.150 35.640 180.210 ;
        RECT 33.955 180.010 35.640 180.150 ;
        RECT 33.955 179.965 34.245 180.010 ;
        RECT 18.315 179.810 18.605 179.855 ;
        RECT 22.440 179.810 22.760 179.870 ;
        RECT 18.315 179.670 22.760 179.810 ;
        RECT 18.315 179.625 18.605 179.670 ;
        RECT 19.770 179.530 19.910 179.670 ;
        RECT 22.440 179.610 22.760 179.670 ;
        RECT 28.435 179.810 28.725 179.855 ;
        RECT 33.020 179.810 33.340 179.870 ;
        RECT 28.435 179.670 33.340 179.810 ;
        RECT 28.435 179.625 28.725 179.670 ;
        RECT 33.020 179.610 33.340 179.670 ;
        RECT 19.680 179.270 20.000 179.530 ;
        RECT 20.140 179.270 20.460 179.530 ;
        RECT 27.040 179.470 27.360 179.530 ;
        RECT 27.515 179.470 27.805 179.515 ;
        RECT 27.040 179.330 27.805 179.470 ;
        RECT 33.570 179.470 33.710 179.965 ;
        RECT 35.320 179.950 35.640 180.010 ;
        RECT 35.780 180.200 36.100 180.210 ;
        RECT 35.780 180.195 36.240 180.200 ;
        RECT 35.780 179.965 36.325 180.195 ;
        RECT 35.780 179.950 36.100 179.965 ;
        RECT 36.700 179.950 37.020 180.210 ;
        RECT 38.080 180.150 38.400 180.210 ;
        RECT 37.885 180.010 38.400 180.150 ;
        RECT 38.080 179.950 38.400 180.010 ;
        RECT 38.540 179.950 38.860 180.210 ;
        RECT 39.920 179.950 40.240 180.210 ;
        RECT 40.840 179.950 41.160 180.210 ;
        RECT 41.760 180.195 42.080 180.210 ;
        RECT 41.545 179.965 42.080 180.195 ;
        RECT 41.760 179.950 42.080 179.965 ;
        RECT 42.680 180.150 43.000 180.210 ;
        RECT 43.615 180.150 43.905 180.195 ;
        RECT 42.680 180.010 43.905 180.150 ;
        RECT 42.680 179.950 43.000 180.010 ;
        RECT 43.615 179.965 43.905 180.010 ;
        RECT 44.075 179.965 44.365 180.195 ;
        RECT 47.740 180.150 48.060 180.210 ;
        RECT 48.215 180.150 48.505 180.195 ;
        RECT 47.740 180.010 48.505 180.150 ;
        RECT 37.175 179.810 37.465 179.855 ;
        RECT 37.175 179.670 37.850 179.810 ;
        RECT 37.175 179.625 37.465 179.670 ;
        RECT 37.710 179.530 37.850 179.670 ;
        RECT 36.700 179.470 37.020 179.530 ;
        RECT 33.570 179.330 37.020 179.470 ;
        RECT 27.040 179.270 27.360 179.330 ;
        RECT 27.515 179.285 27.805 179.330 ;
        RECT 36.700 179.270 37.020 179.330 ;
        RECT 37.620 179.270 37.940 179.530 ;
        RECT 38.170 179.470 38.310 179.950 ;
        RECT 40.380 179.610 40.700 179.870 ;
        RECT 43.140 179.470 43.460 179.530 ;
        RECT 38.170 179.330 43.460 179.470 ;
        RECT 44.150 179.470 44.290 179.965 ;
        RECT 47.740 179.950 48.060 180.010 ;
        RECT 48.215 179.965 48.505 180.010 ;
        RECT 45.915 179.810 46.205 179.855 ;
        RECT 46.360 179.810 46.680 179.870 ;
        RECT 45.915 179.670 46.680 179.810 ;
        RECT 45.915 179.625 46.205 179.670 ;
        RECT 46.360 179.610 46.680 179.670 ;
        RECT 46.835 179.810 47.125 179.855 ;
        RECT 47.280 179.810 47.600 179.870 ;
        RECT 46.835 179.670 47.600 179.810 ;
        RECT 46.835 179.625 47.125 179.670 ;
        RECT 47.280 179.610 47.600 179.670 ;
        RECT 44.520 179.470 44.840 179.530 ;
        RECT 48.750 179.515 48.890 180.350 ;
        RECT 49.120 180.350 51.725 180.490 ;
        RECT 49.120 180.290 49.440 180.350 ;
        RECT 51.435 180.305 51.725 180.350 ;
        RECT 49.580 180.150 49.900 180.210 ;
        RECT 50.500 180.150 50.820 180.210 ;
        RECT 51.970 180.150 52.110 180.690 ;
        RECT 52.815 180.645 53.105 180.690 ;
        RECT 53.810 180.490 53.950 180.985 ;
        RECT 56.020 180.970 56.340 181.030 ;
        RECT 57.400 180.830 57.720 180.890 ;
        RECT 57.030 180.690 57.720 180.830 ;
        RECT 57.030 180.490 57.170 180.690 ;
        RECT 57.400 180.630 57.720 180.690 ;
        RECT 57.875 180.645 58.165 180.875 ;
        RECT 58.320 180.830 58.640 180.890 ;
        RECT 59.255 180.830 59.545 180.875 ;
        RECT 58.320 180.690 59.545 180.830 ;
        RECT 60.710 180.830 60.850 181.030 ;
        RECT 62.000 181.030 63.225 181.170 ;
        RECT 62.000 180.970 62.320 181.030 ;
        RECT 62.935 180.985 63.225 181.030 ;
        RECT 63.840 180.970 64.160 181.230 ;
        RECT 69.360 181.170 69.680 181.230 ;
        RECT 81.335 181.170 81.625 181.215 ;
        RECT 69.360 181.030 81.625 181.170 ;
        RECT 69.360 180.970 69.680 181.030 ;
        RECT 81.335 180.985 81.625 181.030 ;
        RECT 70.740 180.830 71.060 180.890 ;
        RECT 60.710 180.690 62.230 180.830 ;
        RECT 57.950 180.490 58.090 180.645 ;
        RECT 58.320 180.630 58.640 180.690 ;
        RECT 59.255 180.645 59.545 180.690 ;
        RECT 61.540 180.490 61.860 180.550 ;
        RECT 53.810 180.350 57.170 180.490 ;
        RECT 54.640 180.150 54.960 180.210 ;
        RECT 57.030 180.195 57.170 180.350 ;
        RECT 57.490 180.350 58.090 180.490 ;
        RECT 58.410 180.350 61.860 180.490 ;
        RECT 57.490 180.210 57.630 180.350 ;
        RECT 55.115 180.150 55.405 180.195 ;
        RECT 49.580 180.010 50.820 180.150 ;
        RECT 49.580 179.950 49.900 180.010 ;
        RECT 50.500 179.950 50.820 180.010 ;
        RECT 51.050 180.010 52.110 180.150 ;
        RECT 52.430 180.010 55.405 180.150 ;
        RECT 51.050 179.870 51.190 180.010 ;
        RECT 50.960 179.610 51.280 179.870 ;
        RECT 44.150 179.330 44.840 179.470 ;
        RECT 43.140 179.270 43.460 179.330 ;
        RECT 44.520 179.270 44.840 179.330 ;
        RECT 48.675 179.470 48.965 179.515 ;
        RECT 52.430 179.470 52.570 180.010 ;
        RECT 54.640 179.950 54.960 180.010 ;
        RECT 55.115 179.965 55.405 180.010 ;
        RECT 56.955 179.965 57.245 180.195 ;
        RECT 57.400 179.950 57.720 180.210 ;
        RECT 52.800 179.810 53.120 179.870 ;
        RECT 56.035 179.810 56.325 179.855 ;
        RECT 52.800 179.670 56.325 179.810 ;
        RECT 52.800 179.610 53.120 179.670 ;
        RECT 56.035 179.625 56.325 179.670 ;
        RECT 48.675 179.330 52.570 179.470 ;
        RECT 56.110 179.470 56.250 179.625 ;
        RECT 56.480 179.610 56.800 179.870 ;
        RECT 58.410 179.470 58.550 180.350 ;
        RECT 61.540 180.290 61.860 180.350 ;
        RECT 59.240 179.950 59.560 180.210 ;
        RECT 59.700 180.150 60.020 180.210 ;
        RECT 61.080 180.195 61.400 180.210 ;
        RECT 62.090 180.195 62.230 180.690 ;
        RECT 66.230 180.690 71.060 180.830 ;
        RECT 64.760 180.490 65.080 180.550 ;
        RECT 66.230 180.490 66.370 180.690 ;
        RECT 70.740 180.630 71.060 180.690 ;
        RECT 75.340 180.630 75.660 180.890 ;
        RECT 78.560 180.830 78.880 180.890 ;
        RECT 79.495 180.830 79.785 180.875 ;
        RECT 78.560 180.690 79.785 180.830 ;
        RECT 78.560 180.630 78.880 180.690 ;
        RECT 79.495 180.645 79.785 180.690 ;
        RECT 81.780 180.830 82.100 180.890 ;
        RECT 81.780 180.690 82.930 180.830 ;
        RECT 81.780 180.630 82.100 180.690 ;
        RECT 64.760 180.350 66.370 180.490 ;
        RECT 64.760 180.290 65.080 180.350 ;
        RECT 60.635 180.150 60.925 180.195 ;
        RECT 59.700 180.010 60.925 180.150 ;
        RECT 59.700 179.950 60.020 180.010 ;
        RECT 60.635 179.965 60.925 180.010 ;
        RECT 61.080 179.965 61.410 180.195 ;
        RECT 62.015 179.965 62.305 180.195 ;
        RECT 63.380 180.150 63.700 180.210 ;
        RECT 66.230 180.195 66.370 180.350 ;
        RECT 67.150 180.350 82.470 180.490 ;
        RECT 67.150 180.210 67.290 180.350 ;
        RECT 82.330 180.210 82.470 180.350 ;
        RECT 65.235 180.150 65.525 180.195 ;
        RECT 63.380 180.010 65.525 180.150 ;
        RECT 61.080 179.950 61.400 179.965 ;
        RECT 63.380 179.950 63.700 180.010 ;
        RECT 65.235 179.965 65.525 180.010 ;
        RECT 65.695 179.965 65.985 180.195 ;
        RECT 66.155 179.965 66.445 180.195 ;
        RECT 60.160 179.610 60.480 179.870 ;
        RECT 65.770 179.810 65.910 179.965 ;
        RECT 67.060 179.950 67.380 180.210 ;
        RECT 67.520 179.950 67.840 180.210 ;
        RECT 68.900 179.950 69.220 180.210 ;
        RECT 71.660 180.150 71.980 180.210 ;
        RECT 70.370 180.010 71.980 180.150 ;
        RECT 70.370 179.810 70.510 180.010 ;
        RECT 71.660 179.950 71.980 180.010 ;
        RECT 72.120 180.150 72.440 180.210 ;
        RECT 75.800 180.150 76.120 180.210 ;
        RECT 78.115 180.150 78.405 180.195 ;
        RECT 72.120 180.010 78.405 180.150 ;
        RECT 72.120 179.950 72.440 180.010 ;
        RECT 75.800 179.950 76.120 180.010 ;
        RECT 78.115 179.965 78.405 180.010 ;
        RECT 79.020 179.950 79.340 180.210 ;
        RECT 82.240 179.950 82.560 180.210 ;
        RECT 82.790 180.150 82.930 180.690 ;
        RECT 83.160 180.630 83.480 180.890 ;
        RECT 83.635 180.150 83.925 180.195 ;
        RECT 82.790 180.010 83.925 180.150 ;
        RECT 83.635 179.965 83.925 180.010 ;
        RECT 84.095 179.965 84.385 180.195 ;
        RECT 65.770 179.670 70.510 179.810 ;
        RECT 70.740 179.810 71.060 179.870 ;
        RECT 84.170 179.810 84.310 179.965 ;
        RECT 70.740 179.670 84.310 179.810 ;
        RECT 67.150 179.530 67.290 179.670 ;
        RECT 70.740 179.610 71.060 179.670 ;
        RECT 56.110 179.330 58.550 179.470 ;
        RECT 48.675 179.285 48.965 179.330 ;
        RECT 67.060 179.270 67.380 179.530 ;
        RECT 67.995 179.470 68.285 179.515 ;
        RECT 68.440 179.470 68.760 179.530 ;
        RECT 67.995 179.330 68.760 179.470 ;
        RECT 67.995 179.285 68.285 179.330 ;
        RECT 68.440 179.270 68.760 179.330 ;
        RECT 85.000 179.270 85.320 179.530 ;
        RECT 15.930 178.650 87.230 179.130 ;
        RECT 23.835 178.265 24.125 178.495 ;
        RECT 31.180 178.450 31.500 178.510 ;
        RECT 38.080 178.450 38.400 178.510 ;
        RECT 44.075 178.450 44.365 178.495 ;
        RECT 31.180 178.310 44.365 178.450 ;
        RECT 15.540 178.110 15.860 178.170 ;
        RECT 23.910 178.110 24.050 178.265 ;
        RECT 31.180 178.250 31.500 178.310 ;
        RECT 38.080 178.250 38.400 178.310 ;
        RECT 44.075 178.265 44.365 178.310 ;
        RECT 44.980 178.250 45.300 178.510 ;
        RECT 46.360 178.300 46.680 178.510 ;
        RECT 49.135 178.450 49.425 178.495 ;
        RECT 50.960 178.450 51.280 178.510 ;
        RECT 46.910 178.310 47.510 178.450 ;
        RECT 46.910 178.300 47.050 178.310 ;
        RECT 46.360 178.250 47.050 178.300 ;
        RECT 15.540 177.970 24.050 178.110 ;
        RECT 31.655 178.110 31.945 178.155 ;
        RECT 33.480 178.110 33.800 178.170 ;
        RECT 31.655 177.970 33.800 178.110 ;
        RECT 15.540 177.910 15.860 177.970 ;
        RECT 31.655 177.925 31.945 177.970 ;
        RECT 33.480 177.910 33.800 177.970 ;
        RECT 40.380 178.110 40.700 178.170 ;
        RECT 46.455 178.160 47.050 178.250 ;
        RECT 47.370 178.110 47.510 178.310 ;
        RECT 49.135 178.310 51.280 178.450 ;
        RECT 49.135 178.265 49.425 178.310 ;
        RECT 50.960 178.250 51.280 178.310 ;
        RECT 61.080 178.450 61.400 178.510 ;
        RECT 62.935 178.450 63.225 178.495 ;
        RECT 61.080 178.310 63.225 178.450 ;
        RECT 61.080 178.250 61.400 178.310 ;
        RECT 57.860 178.110 58.180 178.170 ;
        RECT 59.715 178.110 60.005 178.155 ;
        RECT 40.380 177.970 43.830 178.110 ;
        RECT 47.370 177.970 54.870 178.110 ;
        RECT 40.380 177.910 40.700 177.970 ;
        RECT 43.690 177.830 43.830 177.970 ;
        RECT 17.380 177.570 17.700 177.830 ;
        RECT 19.680 177.570 20.000 177.830 ;
        RECT 20.465 177.770 20.755 177.815 ;
        RECT 22.440 177.770 22.760 177.830 ;
        RECT 20.465 177.630 22.760 177.770 ;
        RECT 20.465 177.585 20.755 177.630 ;
        RECT 22.440 177.570 22.760 177.630 ;
        RECT 22.900 177.770 23.220 177.830 ;
        RECT 23.375 177.770 23.665 177.815 ;
        RECT 22.900 177.630 23.665 177.770 ;
        RECT 22.900 177.570 23.220 177.630 ;
        RECT 23.375 177.585 23.665 177.630 ;
        RECT 24.740 177.570 25.060 177.830 ;
        RECT 25.215 177.585 25.505 177.815 ;
        RECT 31.195 177.585 31.485 177.815 ;
        RECT 32.100 177.770 32.420 177.830 ;
        RECT 37.620 177.770 37.940 177.830 ;
        RECT 32.100 177.630 37.940 177.770 ;
        RECT 15.080 177.430 15.400 177.490 ;
        RECT 25.290 177.430 25.430 177.585 ;
        RECT 15.080 177.290 25.430 177.430 ;
        RECT 31.270 177.430 31.410 177.585 ;
        RECT 32.100 177.570 32.420 177.630 ;
        RECT 37.620 177.570 37.940 177.630 ;
        RECT 43.155 177.585 43.445 177.815 ;
        RECT 31.640 177.430 31.960 177.490 ;
        RECT 33.940 177.430 34.260 177.490 ;
        RECT 31.270 177.290 34.260 177.430 ;
        RECT 15.080 177.230 15.400 177.290 ;
        RECT 31.640 177.230 31.960 177.290 ;
        RECT 33.940 177.230 34.260 177.290 ;
        RECT 42.680 177.430 43.000 177.490 ;
        RECT 43.230 177.430 43.370 177.585 ;
        RECT 43.600 177.570 43.920 177.830 ;
        RECT 44.980 177.770 45.300 177.830 ;
        RECT 45.455 177.770 45.745 177.815 ;
        RECT 44.980 177.630 45.745 177.770 ;
        RECT 46.820 177.690 47.140 177.950 ;
        RECT 44.980 177.570 45.300 177.630 ;
        RECT 45.455 177.585 45.745 177.630 ;
        RECT 46.835 177.585 47.125 177.690 ;
        RECT 47.755 177.585 48.045 177.815 ;
        RECT 48.200 177.770 48.520 177.830 ;
        RECT 48.675 177.770 48.965 177.815 ;
        RECT 48.200 177.630 48.965 177.770 ;
        RECT 42.680 177.290 43.370 177.430 ;
        RECT 43.690 177.290 47.055 177.430 ;
        RECT 42.680 177.230 43.000 177.290 ;
        RECT 43.690 177.150 43.830 177.290 ;
        RECT 21.520 176.890 21.840 177.150 ;
        RECT 26.120 176.890 26.440 177.150 ;
        RECT 42.235 177.090 42.525 177.135 ;
        RECT 43.600 177.090 43.920 177.150 ;
        RECT 42.235 176.950 43.920 177.090 ;
        RECT 42.235 176.905 42.525 176.950 ;
        RECT 43.600 176.890 43.920 176.950 ;
        RECT 18.300 176.550 18.620 176.810 ;
        RECT 22.440 176.550 22.760 176.810 ;
        RECT 36.700 176.750 37.020 176.810 ;
        RECT 38.540 176.750 38.860 176.810 ;
        RECT 36.700 176.610 38.860 176.750 ;
        RECT 36.700 176.550 37.020 176.610 ;
        RECT 38.540 176.550 38.860 176.610 ;
        RECT 44.520 176.750 44.840 176.810 ;
        RECT 45.455 176.750 45.745 176.795 ;
        RECT 44.520 176.610 45.745 176.750 ;
        RECT 46.915 176.750 47.055 177.290 ;
        RECT 47.280 177.090 47.600 177.150 ;
        RECT 47.830 177.090 47.970 177.585 ;
        RECT 48.200 177.570 48.520 177.630 ;
        RECT 48.675 177.585 48.965 177.630 ;
        RECT 50.055 177.770 50.345 177.815 ;
        RECT 50.960 177.770 51.280 177.830 ;
        RECT 50.055 177.630 51.280 177.770 ;
        RECT 50.055 177.585 50.345 177.630 ;
        RECT 50.960 177.570 51.280 177.630 ;
        RECT 51.420 177.570 51.740 177.830 ;
        RECT 51.880 177.570 52.200 177.830 ;
        RECT 52.815 177.770 53.105 177.815 ;
        RECT 53.720 177.770 54.040 177.830 ;
        RECT 52.815 177.630 54.040 177.770 ;
        RECT 52.815 177.585 53.105 177.630 ;
        RECT 53.720 177.570 54.040 177.630 ;
        RECT 54.180 177.570 54.500 177.830 ;
        RECT 54.730 177.770 54.870 177.970 ;
        RECT 57.860 177.970 60.005 178.110 ;
        RECT 57.860 177.910 58.180 177.970 ;
        RECT 59.715 177.925 60.005 177.970 ;
        RECT 61.630 177.925 61.770 178.310 ;
        RECT 62.935 178.265 63.225 178.310 ;
        RECT 68.900 178.450 69.220 178.510 ;
        RECT 76.260 178.450 76.580 178.510 ;
        RECT 68.900 178.310 76.580 178.450 ;
        RECT 68.900 178.250 69.220 178.310 ;
        RECT 62.460 178.110 62.780 178.170 ;
        RECT 67.060 178.110 67.380 178.170 ;
        RECT 69.910 178.155 70.050 178.310 ;
        RECT 76.260 178.250 76.580 178.310 ;
        RECT 79.020 178.450 79.340 178.510 ;
        RECT 82.240 178.450 82.560 178.510 ;
        RECT 79.020 178.310 82.560 178.450 ;
        RECT 79.020 178.250 79.340 178.310 ;
        RECT 82.240 178.250 82.560 178.310 ;
        RECT 69.375 178.110 69.665 178.155 ;
        RECT 62.460 177.970 66.830 178.110 ;
        RECT 58.335 177.770 58.625 177.815 ;
        RECT 58.780 177.770 59.100 177.830 ;
        RECT 54.730 177.630 57.630 177.770 ;
        RECT 52.355 177.430 52.645 177.475 ;
        RECT 48.750 177.290 52.645 177.430 ;
        RECT 48.750 177.150 48.890 177.290 ;
        RECT 52.355 177.245 52.645 177.290 ;
        RECT 55.575 177.245 55.865 177.475 ;
        RECT 56.035 177.430 56.325 177.475 ;
        RECT 56.940 177.430 57.260 177.490 ;
        RECT 56.035 177.290 57.260 177.430 ;
        RECT 57.490 177.430 57.630 177.630 ;
        RECT 58.335 177.630 59.100 177.770 ;
        RECT 58.335 177.585 58.625 177.630 ;
        RECT 58.780 177.570 59.100 177.630 ;
        RECT 59.240 177.570 59.560 177.830 ;
        RECT 60.160 177.770 60.480 177.830 ;
        RECT 60.635 177.770 60.925 177.815 ;
        RECT 60.160 177.630 60.925 177.770 ;
        RECT 60.160 177.570 60.480 177.630 ;
        RECT 60.635 177.585 60.925 177.630 ;
        RECT 57.875 177.430 58.165 177.475 ;
        RECT 57.490 177.290 60.390 177.430 ;
        RECT 56.035 177.245 56.325 177.290 ;
        RECT 47.280 176.950 47.970 177.090 ;
        RECT 47.280 176.890 47.600 176.950 ;
        RECT 48.200 176.890 48.520 177.150 ;
        RECT 48.660 176.890 48.980 177.150 ;
        RECT 50.515 177.090 50.805 177.135 ;
        RECT 52.800 177.090 53.120 177.150 ;
        RECT 50.515 176.950 53.120 177.090 ;
        RECT 50.515 176.905 50.805 176.950 ;
        RECT 52.800 176.890 53.120 176.950 ;
        RECT 53.275 177.090 53.565 177.135 ;
        RECT 55.650 177.090 55.790 177.245 ;
        RECT 56.940 177.230 57.260 177.290 ;
        RECT 57.875 177.245 58.165 177.290 ;
        RECT 59.715 177.090 60.005 177.135 ;
        RECT 53.275 176.950 55.330 177.090 ;
        RECT 55.650 176.950 60.005 177.090 ;
        RECT 53.275 176.905 53.565 176.950 ;
        RECT 49.120 176.750 49.440 176.810 ;
        RECT 46.915 176.610 49.440 176.750 ;
        RECT 44.520 176.550 44.840 176.610 ;
        RECT 45.455 176.565 45.745 176.610 ;
        RECT 49.120 176.550 49.440 176.610 ;
        RECT 53.720 176.750 54.040 176.810 ;
        RECT 54.655 176.750 54.945 176.795 ;
        RECT 53.720 176.610 54.945 176.750 ;
        RECT 55.190 176.750 55.330 176.950 ;
        RECT 59.715 176.905 60.005 176.950 ;
        RECT 56.020 176.750 56.340 176.810 ;
        RECT 55.190 176.610 56.340 176.750 ;
        RECT 53.720 176.550 54.040 176.610 ;
        RECT 54.655 176.565 54.945 176.610 ;
        RECT 56.020 176.550 56.340 176.610 ;
        RECT 56.940 176.750 57.260 176.810 ;
        RECT 58.795 176.750 59.085 176.795 ;
        RECT 56.940 176.610 59.085 176.750 ;
        RECT 56.940 176.550 57.260 176.610 ;
        RECT 58.795 176.565 59.085 176.610 ;
        RECT 59.240 176.750 59.560 176.810 ;
        RECT 60.250 176.750 60.390 177.290 ;
        RECT 60.710 177.090 60.850 177.585 ;
        RECT 61.080 177.570 61.400 177.830 ;
        RECT 61.580 177.695 61.870 177.925 ;
        RECT 62.460 177.910 62.780 177.970 ;
        RECT 64.315 177.770 64.605 177.815 ;
        RECT 62.550 177.630 64.605 177.770 ;
        RECT 62.550 177.490 62.690 177.630 ;
        RECT 64.315 177.585 64.605 177.630 ;
        RECT 65.220 177.770 65.540 177.830 ;
        RECT 65.695 177.770 65.985 177.815 ;
        RECT 65.220 177.630 65.985 177.770 ;
        RECT 65.220 177.570 65.540 177.630 ;
        RECT 65.695 177.585 65.985 177.630 ;
        RECT 62.460 177.230 62.780 177.490 ;
        RECT 63.380 177.430 63.700 177.490 ;
        RECT 63.855 177.430 64.145 177.475 ;
        RECT 63.380 177.290 64.145 177.430 ;
        RECT 63.380 177.230 63.700 177.290 ;
        RECT 63.855 177.245 64.145 177.290 ;
        RECT 64.760 177.430 65.080 177.490 ;
        RECT 66.155 177.430 66.445 177.475 ;
        RECT 64.760 177.290 66.445 177.430 ;
        RECT 66.690 177.430 66.830 177.970 ;
        RECT 67.060 177.970 69.665 178.110 ;
        RECT 67.060 177.910 67.380 177.970 ;
        RECT 69.375 177.925 69.665 177.970 ;
        RECT 69.835 177.925 70.125 178.155 ;
        RECT 75.815 178.110 76.105 178.155 ;
        RECT 79.480 178.110 79.800 178.170 ;
        RECT 75.815 177.970 79.800 178.110 ;
        RECT 75.815 177.925 76.105 177.970 ;
        RECT 79.480 177.910 79.800 177.970 ;
        RECT 68.900 177.570 69.220 177.830 ;
        RECT 70.755 177.585 71.045 177.815 ;
        RECT 72.135 177.770 72.425 177.815 ;
        RECT 73.040 177.770 73.360 177.830 ;
        RECT 74.880 177.770 75.200 177.830 ;
        RECT 72.135 177.630 75.200 177.770 ;
        RECT 72.135 177.585 72.425 177.630 ;
        RECT 70.830 177.430 70.970 177.585 ;
        RECT 73.040 177.570 73.360 177.630 ;
        RECT 74.880 177.570 75.200 177.630 ;
        RECT 72.580 177.430 72.900 177.490 ;
        RECT 73.515 177.430 73.805 177.475 ;
        RECT 66.690 177.290 72.350 177.430 ;
        RECT 64.760 177.230 65.080 177.290 ;
        RECT 66.155 177.245 66.445 177.290 ;
        RECT 67.995 177.090 68.285 177.135 ;
        RECT 60.710 176.950 68.285 177.090 ;
        RECT 67.995 176.905 68.285 176.950 ;
        RECT 69.360 177.090 69.680 177.150 ;
        RECT 71.200 177.090 71.520 177.150 ;
        RECT 69.360 176.950 71.520 177.090 ;
        RECT 72.210 177.090 72.350 177.290 ;
        RECT 72.580 177.290 73.805 177.430 ;
        RECT 72.580 177.230 72.900 177.290 ;
        RECT 73.515 177.245 73.805 177.290 ;
        RECT 73.960 177.430 74.280 177.490 ;
        RECT 77.180 177.430 77.500 177.490 ;
        RECT 73.960 177.290 77.500 177.430 ;
        RECT 73.960 177.230 74.280 177.290 ;
        RECT 77.180 177.230 77.500 177.290 ;
        RECT 81.780 177.090 82.100 177.150 ;
        RECT 72.210 176.950 82.100 177.090 ;
        RECT 69.360 176.890 69.680 176.950 ;
        RECT 71.200 176.890 71.520 176.950 ;
        RECT 81.780 176.890 82.100 176.950 ;
        RECT 59.240 176.610 60.390 176.750 ;
        RECT 61.540 176.750 61.860 176.810 ;
        RECT 62.460 176.750 62.780 176.810 ;
        RECT 61.540 176.610 62.780 176.750 ;
        RECT 59.240 176.550 59.560 176.610 ;
        RECT 61.540 176.550 61.860 176.610 ;
        RECT 62.460 176.550 62.780 176.610 ;
        RECT 63.380 176.750 63.700 176.810 ;
        RECT 64.760 176.750 65.080 176.810 ;
        RECT 63.380 176.610 65.080 176.750 ;
        RECT 63.380 176.550 63.700 176.610 ;
        RECT 64.760 176.550 65.080 176.610 ;
        RECT 68.900 176.750 69.220 176.810 ;
        RECT 73.960 176.750 74.280 176.810 ;
        RECT 68.900 176.610 74.280 176.750 ;
        RECT 68.900 176.550 69.220 176.610 ;
        RECT 73.960 176.550 74.280 176.610 ;
        RECT 80.860 176.750 81.180 176.810 ;
        RECT 82.240 176.750 82.560 176.810 ;
        RECT 80.860 176.610 82.560 176.750 ;
        RECT 80.860 176.550 81.180 176.610 ;
        RECT 82.240 176.550 82.560 176.610 ;
        RECT 15.930 175.930 87.230 176.410 ;
        RECT 31.655 175.730 31.945 175.775 ;
        RECT 39.460 175.730 39.780 175.790 ;
        RECT 53.260 175.730 53.580 175.790 ;
        RECT 59.715 175.730 60.005 175.775 ;
        RECT 61.080 175.730 61.400 175.790 ;
        RECT 31.655 175.590 39.780 175.730 ;
        RECT 31.655 175.545 31.945 175.590 ;
        RECT 39.460 175.530 39.780 175.590 ;
        RECT 49.030 175.590 53.580 175.730 ;
        RECT 32.100 175.390 32.420 175.450 ;
        RECT 19.770 175.250 32.420 175.390 ;
        RECT 17.840 175.050 18.160 175.110 ;
        RECT 19.770 175.050 19.910 175.250 ;
        RECT 32.100 175.190 32.420 175.250 ;
        RECT 37.160 175.390 37.480 175.450 ;
        RECT 49.030 175.390 49.170 175.590 ;
        RECT 53.260 175.530 53.580 175.590 ;
        RECT 53.810 175.590 56.710 175.730 ;
        RECT 37.160 175.250 49.170 175.390 ;
        RECT 49.595 175.390 49.885 175.435 ;
        RECT 50.960 175.390 51.280 175.450 ;
        RECT 49.595 175.250 51.280 175.390 ;
        RECT 37.160 175.190 37.480 175.250 ;
        RECT 49.595 175.205 49.885 175.250 ;
        RECT 50.960 175.190 51.280 175.250 ;
        RECT 52.355 175.205 52.645 175.435 ;
        RECT 52.800 175.390 53.120 175.450 ;
        RECT 53.810 175.390 53.950 175.590 ;
        RECT 52.800 175.250 53.950 175.390 ;
        RECT 55.575 175.390 55.865 175.435 ;
        RECT 56.020 175.390 56.340 175.450 ;
        RECT 55.575 175.250 56.340 175.390 ;
        RECT 56.570 175.390 56.710 175.590 ;
        RECT 59.715 175.590 61.400 175.730 ;
        RECT 59.715 175.545 60.005 175.590 ;
        RECT 61.080 175.530 61.400 175.590 ;
        RECT 62.460 175.730 62.780 175.790 ;
        RECT 63.395 175.730 63.685 175.775 ;
        RECT 62.460 175.590 63.685 175.730 ;
        RECT 62.460 175.530 62.780 175.590 ;
        RECT 63.395 175.545 63.685 175.590 ;
        RECT 65.695 175.730 65.985 175.775 ;
        RECT 67.980 175.730 68.300 175.790 ;
        RECT 71.200 175.730 71.520 175.790 ;
        RECT 65.695 175.590 68.300 175.730 ;
        RECT 65.695 175.545 65.985 175.590 ;
        RECT 67.980 175.530 68.300 175.590 ;
        RECT 68.990 175.590 71.520 175.730 ;
        RECT 56.570 175.250 66.370 175.390 ;
        RECT 17.840 174.910 19.910 175.050 ;
        RECT 17.840 174.850 18.160 174.910 ;
        RECT 19.220 174.510 19.540 174.770 ;
        RECT 19.770 174.755 19.910 174.910 ;
        RECT 20.600 174.850 20.920 175.110 ;
        RECT 22.440 175.050 22.760 175.110 ;
        RECT 41.300 175.050 41.620 175.110 ;
        RECT 52.430 175.050 52.570 175.205 ;
        RECT 52.800 175.190 53.120 175.250 ;
        RECT 55.575 175.205 55.865 175.250 ;
        RECT 56.020 175.190 56.340 175.250 ;
        RECT 22.440 174.910 41.620 175.050 ;
        RECT 22.440 174.850 22.760 174.910 ;
        RECT 41.300 174.850 41.620 174.910 ;
        RECT 49.670 174.910 52.570 175.050 ;
        RECT 53.260 175.050 53.580 175.110 ;
        RECT 61.080 175.050 61.400 175.110 ;
        RECT 53.260 174.910 57.170 175.050 ;
        RECT 19.695 174.525 19.985 174.755 ;
        RECT 21.075 174.710 21.365 174.755 ;
        RECT 25.660 174.710 25.980 174.770 ;
        RECT 21.075 174.570 25.980 174.710 ;
        RECT 21.075 174.525 21.365 174.570 ;
        RECT 25.660 174.510 25.980 174.570 ;
        RECT 26.580 174.510 26.900 174.770 ;
        RECT 29.340 174.510 29.660 174.770 ;
        RECT 30.735 174.525 31.025 174.755 ;
        RECT 33.940 174.710 34.260 174.770 ;
        RECT 36.255 174.710 36.545 174.755 ;
        RECT 33.940 174.570 36.545 174.710 ;
        RECT 26.670 174.370 26.810 174.510 ;
        RECT 30.810 174.370 30.950 174.525 ;
        RECT 33.940 174.510 34.260 174.570 ;
        RECT 36.255 174.525 36.545 174.570 ;
        RECT 37.175 174.710 37.465 174.755 ;
        RECT 39.920 174.710 40.240 174.770 ;
        RECT 49.670 174.755 49.810 174.910 ;
        RECT 53.260 174.850 53.580 174.910 ;
        RECT 37.175 174.570 40.240 174.710 ;
        RECT 37.175 174.525 37.465 174.570 ;
        RECT 39.920 174.510 40.240 174.570 ;
        RECT 49.595 174.525 49.885 174.755 ;
        RECT 50.960 174.510 51.280 174.770 ;
        RECT 53.720 174.510 54.040 174.770 ;
        RECT 57.030 174.755 57.170 174.910 ;
        RECT 59.330 174.910 61.400 175.050 ;
        RECT 56.495 174.710 56.785 174.755 ;
        RECT 56.110 174.570 56.785 174.710 ;
        RECT 26.670 174.230 30.950 174.370 ;
        RECT 52.340 174.170 52.660 174.430 ;
        RECT 54.180 174.170 54.500 174.430 ;
        RECT 56.110 174.370 56.250 174.570 ;
        RECT 56.495 174.525 56.785 174.570 ;
        RECT 56.955 174.525 57.245 174.755 ;
        RECT 57.415 174.525 57.705 174.755 ;
        RECT 57.860 174.710 58.180 174.770 ;
        RECT 59.330 174.755 59.470 174.910 ;
        RECT 61.080 174.850 61.400 174.910 ;
        RECT 61.540 175.050 61.860 175.110 ;
        RECT 61.540 174.910 64.070 175.050 ;
        RECT 61.540 174.850 61.860 174.910 ;
        RECT 58.335 174.710 58.625 174.755 ;
        RECT 57.860 174.570 58.625 174.710 ;
        RECT 57.490 174.370 57.630 174.525 ;
        RECT 57.860 174.510 58.180 174.570 ;
        RECT 58.335 174.525 58.625 174.570 ;
        RECT 59.255 174.525 59.545 174.755 ;
        RECT 60.160 174.710 60.480 174.770 ;
        RECT 60.635 174.710 60.925 174.755 ;
        RECT 60.160 174.570 60.925 174.710 ;
        RECT 60.160 174.510 60.480 174.570 ;
        RECT 60.635 174.525 60.925 174.570 ;
        RECT 62.000 174.510 62.320 174.770 ;
        RECT 62.460 174.510 62.780 174.770 ;
        RECT 56.110 174.230 56.710 174.370 ;
        RECT 57.490 174.230 58.090 174.370 ;
        RECT 18.315 174.030 18.605 174.075 ;
        RECT 26.580 174.030 26.900 174.090 ;
        RECT 18.315 173.890 26.900 174.030 ;
        RECT 18.315 173.845 18.605 173.890 ;
        RECT 26.580 173.830 26.900 173.890 ;
        RECT 28.420 174.030 28.740 174.090 ;
        RECT 29.815 174.030 30.105 174.075 ;
        RECT 28.420 173.890 30.105 174.030 ;
        RECT 28.420 173.830 28.740 173.890 ;
        RECT 29.815 173.845 30.105 173.890 ;
        RECT 36.700 173.830 37.020 174.090 ;
        RECT 42.220 174.030 42.540 174.090 ;
        RECT 49.580 174.030 49.900 174.090 ;
        RECT 50.515 174.030 50.805 174.075 ;
        RECT 42.220 173.890 50.805 174.030 ;
        RECT 42.220 173.830 42.540 173.890 ;
        RECT 49.580 173.830 49.900 173.890 ;
        RECT 50.515 173.845 50.805 173.890 ;
        RECT 51.420 174.030 51.740 174.090 ;
        RECT 51.880 174.030 52.200 174.090 ;
        RECT 51.420 173.890 52.200 174.030 ;
        RECT 51.420 173.830 51.740 173.890 ;
        RECT 51.880 173.830 52.200 173.890 ;
        RECT 53.260 173.830 53.580 174.090 ;
        RECT 54.270 174.030 54.410 174.170 ;
        RECT 56.020 174.030 56.340 174.090 ;
        RECT 54.270 173.890 56.340 174.030 ;
        RECT 56.570 174.030 56.710 174.230 ;
        RECT 57.950 174.090 58.090 174.230 ;
        RECT 61.080 174.170 61.400 174.430 ;
        RECT 61.555 174.370 61.845 174.415 ;
        RECT 62.090 174.370 62.230 174.510 ;
        RECT 61.555 174.230 62.230 174.370 ;
        RECT 63.930 174.370 64.070 174.910 ;
        RECT 64.315 174.770 64.605 174.835 ;
        RECT 64.300 174.510 64.620 174.770 ;
        RECT 64.760 174.510 65.080 174.770 ;
        RECT 65.680 174.510 66.000 174.770 ;
        RECT 66.230 174.755 66.370 175.250 ;
        RECT 67.520 174.850 67.840 175.110 ;
        RECT 68.990 175.050 69.130 175.590 ;
        RECT 71.200 175.530 71.520 175.590 ;
        RECT 72.120 175.530 72.440 175.790 ;
        RECT 72.580 175.730 72.900 175.790 ;
        RECT 75.340 175.730 75.660 175.790 ;
        RECT 72.580 175.590 75.660 175.730 ;
        RECT 72.580 175.530 72.900 175.590 ;
        RECT 75.340 175.530 75.660 175.590 ;
        RECT 78.575 175.730 78.865 175.775 ;
        RECT 79.940 175.730 80.260 175.790 ;
        RECT 78.575 175.590 80.260 175.730 ;
        RECT 78.575 175.545 78.865 175.590 ;
        RECT 79.940 175.530 80.260 175.590 ;
        RECT 81.335 175.730 81.625 175.775 ;
        RECT 81.780 175.730 82.100 175.790 ;
        RECT 81.335 175.590 82.100 175.730 ;
        RECT 81.335 175.545 81.625 175.590 ;
        RECT 81.780 175.530 82.100 175.590 ;
        RECT 83.620 175.730 83.940 175.790 ;
        RECT 86.840 175.730 87.160 175.790 ;
        RECT 83.620 175.590 87.160 175.730 ;
        RECT 83.620 175.530 83.940 175.590 ;
        RECT 86.840 175.530 87.160 175.590 ;
        RECT 69.820 175.190 70.140 175.450 ;
        RECT 72.670 175.390 72.810 175.530 ;
        RECT 76.720 175.390 77.040 175.450 ;
        RECT 71.750 175.250 72.810 175.390 ;
        RECT 73.130 175.250 77.040 175.390 ;
        RECT 68.530 174.910 69.130 175.050 ;
        RECT 71.215 175.050 71.505 175.095 ;
        RECT 71.750 175.050 71.890 175.250 ;
        RECT 72.580 175.095 72.900 175.110 ;
        RECT 73.130 175.095 73.270 175.250 ;
        RECT 76.720 175.190 77.040 175.250 ;
        RECT 77.180 175.390 77.500 175.450 ;
        RECT 77.180 175.250 84.310 175.390 ;
        RECT 77.180 175.190 77.500 175.250 ;
        RECT 71.215 174.910 71.890 175.050 ;
        RECT 68.530 174.755 68.670 174.910 ;
        RECT 71.215 174.865 71.505 174.910 ;
        RECT 72.555 174.865 72.900 175.095 ;
        RECT 73.055 174.865 73.345 175.095 ;
        RECT 82.240 175.050 82.560 175.110 ;
        RECT 83.620 175.050 83.940 175.110 ;
        RECT 76.810 174.910 82.560 175.050 ;
        RECT 72.580 174.850 72.900 174.865 ;
        RECT 66.155 174.525 66.445 174.755 ;
        RECT 68.455 174.525 68.745 174.755 ;
        RECT 69.360 174.510 69.680 174.770 ;
        RECT 70.295 174.525 70.585 174.755 ;
        RECT 66.615 174.370 66.905 174.415 ;
        RECT 70.370 174.370 70.510 174.525 ;
        RECT 73.960 174.510 74.280 174.770 ;
        RECT 74.420 174.510 74.740 174.770 ;
        RECT 75.355 174.525 75.645 174.755 ;
        RECT 75.800 174.710 76.120 174.770 ;
        RECT 76.810 174.755 76.950 174.910 ;
        RECT 82.240 174.850 82.560 174.910 ;
        RECT 82.790 174.910 83.940 175.050 ;
        RECT 76.735 174.710 77.025 174.755 ;
        RECT 75.800 174.570 77.025 174.710 ;
        RECT 75.430 174.370 75.570 174.525 ;
        RECT 75.800 174.510 76.120 174.570 ;
        RECT 76.735 174.525 77.025 174.570 ;
        RECT 79.035 174.525 79.325 174.755 ;
        RECT 81.795 174.710 82.085 174.755 ;
        RECT 82.790 174.710 82.930 174.910 ;
        RECT 83.620 174.850 83.940 174.910 ;
        RECT 81.795 174.570 82.930 174.710 ;
        RECT 81.795 174.525 82.085 174.570 ;
        RECT 63.930 174.230 75.570 174.370 ;
        RECT 79.110 174.370 79.250 174.525 ;
        RECT 83.160 174.510 83.480 174.770 ;
        RECT 84.170 174.755 84.310 175.250 ;
        RECT 84.095 174.525 84.385 174.755 ;
        RECT 86.380 174.370 86.700 174.430 ;
        RECT 79.110 174.230 86.700 174.370 ;
        RECT 61.555 174.185 61.845 174.230 ;
        RECT 66.615 174.185 66.905 174.230 ;
        RECT 86.380 174.170 86.700 174.230 ;
        RECT 57.400 174.030 57.720 174.090 ;
        RECT 56.570 173.890 57.720 174.030 ;
        RECT 56.020 173.830 56.340 173.890 ;
        RECT 57.400 173.830 57.720 173.890 ;
        RECT 57.860 173.830 58.180 174.090 ;
        RECT 58.780 173.830 59.100 174.090 ;
        RECT 59.700 174.030 60.020 174.090 ;
        RECT 64.760 174.030 65.080 174.090 ;
        RECT 59.700 173.890 65.080 174.030 ;
        RECT 59.700 173.830 60.020 173.890 ;
        RECT 64.760 173.830 65.080 173.890 ;
        RECT 67.980 174.030 68.300 174.090 ;
        RECT 70.755 174.030 71.045 174.075 ;
        RECT 74.895 174.030 75.185 174.075 ;
        RECT 67.980 173.890 75.185 174.030 ;
        RECT 67.980 173.830 68.300 173.890 ;
        RECT 70.755 173.845 71.045 173.890 ;
        RECT 74.895 173.845 75.185 173.890 ;
        RECT 75.815 174.030 76.105 174.075 ;
        RECT 84.540 174.030 84.860 174.090 ;
        RECT 75.815 173.890 84.860 174.030 ;
        RECT 75.815 173.845 76.105 173.890 ;
        RECT 84.540 173.830 84.860 173.890 ;
        RECT 85.000 173.830 85.320 174.090 ;
        RECT 15.930 173.210 87.230 173.690 ;
        RECT 19.695 173.010 19.985 173.055 ;
        RECT 20.600 173.010 20.920 173.070 ;
        RECT 19.695 172.870 20.920 173.010 ;
        RECT 19.695 172.825 19.985 172.870 ;
        RECT 20.600 172.810 20.920 172.870 ;
        RECT 21.520 172.810 21.840 173.070 ;
        RECT 27.055 173.010 27.345 173.055 ;
        RECT 28.420 173.010 28.740 173.070 ;
        RECT 27.055 172.870 28.740 173.010 ;
        RECT 27.055 172.825 27.345 172.870 ;
        RECT 28.420 172.810 28.740 172.870 ;
        RECT 29.340 173.010 29.660 173.070 ;
        RECT 33.495 173.010 33.785 173.055 ;
        RECT 29.340 172.870 33.785 173.010 ;
        RECT 29.340 172.810 29.660 172.870 ;
        RECT 33.495 172.825 33.785 172.870 ;
        RECT 36.700 173.010 37.020 173.070 ;
        RECT 37.175 173.010 37.465 173.055 ;
        RECT 36.700 172.870 37.465 173.010 ;
        RECT 36.700 172.810 37.020 172.870 ;
        RECT 37.175 172.825 37.465 172.870 ;
        RECT 42.220 173.010 42.540 173.070 ;
        RECT 42.695 173.010 42.985 173.055 ;
        RECT 42.220 172.870 42.985 173.010 ;
        RECT 42.220 172.810 42.540 172.870 ;
        RECT 42.695 172.825 42.985 172.870 ;
        RECT 44.060 173.010 44.380 173.070 ;
        RECT 44.535 173.010 44.825 173.055 ;
        RECT 54.640 173.010 54.960 173.070 ;
        RECT 44.060 172.870 44.825 173.010 ;
        RECT 44.060 172.810 44.380 172.870 ;
        RECT 44.535 172.825 44.825 172.870 ;
        RECT 45.990 172.870 54.960 173.010 ;
        RECT 25.660 172.670 25.980 172.730 ;
        RECT 43.615 172.670 43.905 172.715 ;
        RECT 25.660 172.530 31.050 172.670 ;
        RECT 25.660 172.470 25.980 172.530 ;
        RECT 26.580 172.130 26.900 172.390 ;
        RECT 27.040 172.330 27.360 172.390 ;
        RECT 27.975 172.330 28.265 172.375 ;
        RECT 27.040 172.190 28.265 172.330 ;
        RECT 27.040 172.130 27.360 172.190 ;
        RECT 27.975 172.145 28.265 172.190 ;
        RECT 29.340 172.130 29.660 172.390 ;
        RECT 30.165 172.130 30.485 172.390 ;
        RECT 30.910 172.375 31.050 172.530 ;
        RECT 35.870 172.530 43.905 172.670 ;
        RECT 30.735 172.190 31.050 172.375 ;
        RECT 30.735 172.145 31.025 172.190 ;
        RECT 32.100 172.130 32.420 172.390 ;
        RECT 32.575 172.330 32.865 172.375 ;
        RECT 34.860 172.330 35.180 172.390 ;
        RECT 32.575 172.190 35.180 172.330 ;
        RECT 32.575 172.145 32.865 172.190 ;
        RECT 34.860 172.130 35.180 172.190 ;
        RECT 21.980 171.790 22.300 172.050 ;
        RECT 22.440 171.790 22.760 172.050 ;
        RECT 35.870 171.990 36.010 172.530 ;
        RECT 43.615 172.485 43.905 172.530 ;
        RECT 36.715 172.330 37.005 172.375 ;
        RECT 39.000 172.330 39.320 172.390 ;
        RECT 36.715 172.190 39.320 172.330 ;
        RECT 36.715 172.145 37.005 172.190 ;
        RECT 39.000 172.130 39.320 172.190 ;
        RECT 41.300 172.330 41.620 172.390 ;
        RECT 42.235 172.330 42.525 172.375 ;
        RECT 41.300 172.190 42.525 172.330 ;
        RECT 41.300 172.130 41.620 172.190 ;
        RECT 42.235 172.145 42.525 172.190 ;
        RECT 44.980 172.330 45.300 172.390 ;
        RECT 45.455 172.330 45.745 172.375 ;
        RECT 44.980 172.190 45.745 172.330 ;
        RECT 44.980 172.130 45.300 172.190 ;
        RECT 45.455 172.145 45.745 172.190 ;
        RECT 28.050 171.850 36.010 171.990 ;
        RECT 37.160 171.990 37.480 172.050 ;
        RECT 37.635 171.990 37.925 172.035 ;
        RECT 37.160 171.850 37.925 171.990 ;
        RECT 28.050 171.695 28.190 171.850 ;
        RECT 37.160 171.790 37.480 171.850 ;
        RECT 37.635 171.805 37.925 171.850 ;
        RECT 38.080 171.990 38.400 172.050 ;
        RECT 44.520 171.990 44.840 172.050 ;
        RECT 38.080 171.850 44.840 171.990 ;
        RECT 38.080 171.790 38.400 171.850 ;
        RECT 44.520 171.790 44.840 171.850 ;
        RECT 27.975 171.465 28.265 171.695 ;
        RECT 31.195 171.650 31.485 171.695 ;
        RECT 34.875 171.650 35.165 171.695 ;
        RECT 31.195 171.510 35.165 171.650 ;
        RECT 31.195 171.465 31.485 171.510 ;
        RECT 34.875 171.465 35.165 171.510 ;
        RECT 43.615 171.650 43.905 171.695 ;
        RECT 45.990 171.650 46.130 172.870 ;
        RECT 54.640 172.810 54.960 172.870 ;
        RECT 55.560 172.810 55.880 173.070 ;
        RECT 56.020 173.010 56.340 173.070 ;
        RECT 62.015 173.010 62.305 173.055 ;
        RECT 66.140 173.010 66.460 173.070 ;
        RECT 56.020 172.870 62.305 173.010 ;
        RECT 56.020 172.810 56.340 172.870 ;
        RECT 62.015 172.825 62.305 172.870 ;
        RECT 63.010 172.870 66.460 173.010 ;
        RECT 46.375 172.670 46.665 172.715 ;
        RECT 50.500 172.670 50.820 172.730 ;
        RECT 46.375 172.530 50.820 172.670 ;
        RECT 46.375 172.485 46.665 172.530 ;
        RECT 50.500 172.470 50.820 172.530 ;
        RECT 50.975 172.670 51.265 172.715 ;
        RECT 51.880 172.670 52.200 172.730 ;
        RECT 50.975 172.530 52.200 172.670 ;
        RECT 50.975 172.485 51.265 172.530 ;
        RECT 51.880 172.470 52.200 172.530 ;
        RECT 52.340 172.670 52.660 172.730 ;
        RECT 52.815 172.670 53.105 172.715 ;
        RECT 52.340 172.530 53.105 172.670 ;
        RECT 52.340 172.470 52.660 172.530 ;
        RECT 52.815 172.485 53.105 172.530 ;
        RECT 46.820 172.130 47.140 172.390 ;
        RECT 50.055 172.145 50.345 172.375 ;
        RECT 50.130 171.990 50.270 172.145 ;
        RECT 51.420 172.130 51.740 172.390 ;
        RECT 53.720 172.130 54.040 172.390 ;
        RECT 54.195 172.145 54.485 172.375 ;
        RECT 54.270 171.990 54.410 172.145 ;
        RECT 56.480 172.130 56.800 172.390 ;
        RECT 57.860 172.130 58.180 172.390 ;
        RECT 58.335 172.330 58.625 172.375 ;
        RECT 58.780 172.330 59.100 172.390 ;
        RECT 58.335 172.190 59.100 172.330 ;
        RECT 58.335 172.145 58.625 172.190 ;
        RECT 58.780 172.130 59.100 172.190 ;
        RECT 60.635 172.330 60.925 172.375 ;
        RECT 61.540 172.330 61.860 172.390 ;
        RECT 63.010 172.375 63.150 172.870 ;
        RECT 66.140 172.810 66.460 172.870 ;
        RECT 67.075 172.825 67.365 173.055 ;
        RECT 69.375 173.010 69.665 173.055 ;
        RECT 80.400 173.010 80.720 173.070 ;
        RECT 69.375 172.870 80.720 173.010 ;
        RECT 69.375 172.825 69.665 172.870 ;
        RECT 66.600 172.670 66.920 172.730 ;
        RECT 63.470 172.530 66.920 172.670 ;
        RECT 67.150 172.670 67.290 172.825 ;
        RECT 80.400 172.810 80.720 172.870 ;
        RECT 81.320 173.010 81.640 173.070 ;
        RECT 83.175 173.010 83.465 173.055 ;
        RECT 81.320 172.870 83.465 173.010 ;
        RECT 81.320 172.810 81.640 172.870 ;
        RECT 83.175 172.825 83.465 172.870 ;
        RECT 69.820 172.670 70.140 172.730 ;
        RECT 75.800 172.670 76.120 172.730 ;
        RECT 67.150 172.530 70.140 172.670 ;
        RECT 63.470 172.375 63.610 172.530 ;
        RECT 66.600 172.470 66.920 172.530 ;
        RECT 69.820 172.470 70.140 172.530 ;
        RECT 70.830 172.530 76.120 172.670 ;
        RECT 60.635 172.190 61.860 172.330 ;
        RECT 60.635 172.145 60.925 172.190 ;
        RECT 61.540 172.130 61.860 172.190 ;
        RECT 62.935 172.145 63.225 172.375 ;
        RECT 63.395 172.145 63.685 172.375 ;
        RECT 65.680 172.130 66.000 172.390 ;
        RECT 66.155 172.330 66.445 172.375 ;
        RECT 67.520 172.330 67.840 172.390 ;
        RECT 66.155 172.190 67.840 172.330 ;
        RECT 66.155 172.145 66.445 172.190 ;
        RECT 67.520 172.130 67.840 172.190 ;
        RECT 68.440 172.130 68.760 172.390 ;
        RECT 70.830 172.375 70.970 172.530 ;
        RECT 75.800 172.470 76.120 172.530 ;
        RECT 70.755 172.145 71.045 172.375 ;
        RECT 71.200 172.130 71.520 172.390 ;
        RECT 71.660 172.330 71.980 172.390 ;
        RECT 72.135 172.330 72.425 172.375 ;
        RECT 71.660 172.190 72.425 172.330 ;
        RECT 71.660 172.130 71.980 172.190 ;
        RECT 72.135 172.145 72.425 172.190 ;
        RECT 73.515 172.330 73.805 172.375 ;
        RECT 74.420 172.330 74.740 172.390 ;
        RECT 73.515 172.190 74.740 172.330 ;
        RECT 73.515 172.145 73.805 172.190 ;
        RECT 74.420 172.130 74.740 172.190 ;
        RECT 74.895 172.350 75.185 172.375 ;
        RECT 74.895 172.210 75.570 172.350 ;
        RECT 74.895 172.145 75.185 172.210 ;
        RECT 56.955 171.990 57.245 172.035 ;
        RECT 50.130 171.850 53.030 171.990 ;
        RECT 54.270 171.850 57.245 171.990 ;
        RECT 43.615 171.510 46.130 171.650 ;
        RECT 46.450 171.510 49.810 171.650 ;
        RECT 43.615 171.465 43.905 171.510 ;
        RECT 32.100 171.310 32.420 171.370 ;
        RECT 35.320 171.310 35.640 171.370 ;
        RECT 32.100 171.170 35.640 171.310 ;
        RECT 32.100 171.110 32.420 171.170 ;
        RECT 35.320 171.110 35.640 171.170 ;
        RECT 37.620 171.310 37.940 171.370 ;
        RECT 44.060 171.310 44.380 171.370 ;
        RECT 37.620 171.170 44.380 171.310 ;
        RECT 37.620 171.110 37.940 171.170 ;
        RECT 44.060 171.110 44.380 171.170 ;
        RECT 44.520 171.310 44.840 171.370 ;
        RECT 46.450 171.310 46.590 171.510 ;
        RECT 44.520 171.170 46.590 171.310 ;
        RECT 49.670 171.310 49.810 171.510 ;
        RECT 50.040 171.450 50.360 171.710 ;
        RECT 52.890 171.695 53.030 171.850 ;
        RECT 56.955 171.805 57.245 171.850 ;
        RECT 59.240 171.990 59.560 172.050 ;
        RECT 60.175 171.990 60.465 172.035 ;
        RECT 75.430 171.990 75.570 172.210 ;
        RECT 76.260 172.330 76.580 172.390 ;
        RECT 76.735 172.330 77.025 172.375 ;
        RECT 76.260 172.190 77.025 172.330 ;
        RECT 76.260 172.130 76.580 172.190 ;
        RECT 76.735 172.145 77.025 172.190 ;
        RECT 59.240 171.850 60.465 171.990 ;
        RECT 59.240 171.790 59.560 171.850 ;
        RECT 60.175 171.805 60.465 171.850 ;
        RECT 61.630 171.850 75.570 171.990 ;
        RECT 52.815 171.465 53.105 171.695 ;
        RECT 59.700 171.650 60.020 171.710 ;
        RECT 61.630 171.695 61.770 171.850 ;
        RECT 53.350 171.510 60.020 171.650 ;
        RECT 53.350 171.310 53.490 171.510 ;
        RECT 59.700 171.450 60.020 171.510 ;
        RECT 61.555 171.465 61.845 171.695 ;
        RECT 62.460 171.650 62.780 171.710 ;
        RECT 63.840 171.650 64.160 171.710 ;
        RECT 62.460 171.510 64.160 171.650 ;
        RECT 62.460 171.450 62.780 171.510 ;
        RECT 63.840 171.450 64.160 171.510 ;
        RECT 64.760 171.450 65.080 171.710 ;
        RECT 73.500 171.650 73.820 171.710 ;
        RECT 65.310 171.510 73.820 171.650 ;
        RECT 49.670 171.170 53.490 171.310 ;
        RECT 64.315 171.310 64.605 171.355 ;
        RECT 65.310 171.310 65.450 171.510 ;
        RECT 73.500 171.450 73.820 171.510 ;
        RECT 73.960 171.650 74.280 171.710 ;
        RECT 74.435 171.650 74.725 171.695 ;
        RECT 73.960 171.510 74.725 171.650 ;
        RECT 73.960 171.450 74.280 171.510 ;
        RECT 74.435 171.465 74.725 171.510 ;
        RECT 75.800 171.450 76.120 171.710 ;
        RECT 64.315 171.170 65.450 171.310 ;
        RECT 44.520 171.110 44.840 171.170 ;
        RECT 64.315 171.125 64.605 171.170 ;
        RECT 15.930 170.490 87.230 170.970 ;
        RECT 19.220 170.090 19.540 170.350 ;
        RECT 31.180 170.290 31.500 170.350 ;
        RECT 24.140 170.150 31.500 170.290 ;
        RECT 21.520 169.410 21.840 169.670 ;
        RECT 21.995 169.610 22.285 169.655 ;
        RECT 22.440 169.610 22.760 169.670 ;
        RECT 24.140 169.610 24.280 170.150 ;
        RECT 31.180 170.090 31.500 170.150 ;
        RECT 33.035 170.290 33.325 170.335 ;
        RECT 33.480 170.290 33.800 170.350 ;
        RECT 33.035 170.150 33.800 170.290 ;
        RECT 33.035 170.105 33.325 170.150 ;
        RECT 33.480 170.090 33.800 170.150 ;
        RECT 34.415 170.290 34.705 170.335 ;
        RECT 34.860 170.290 35.180 170.350 ;
        RECT 34.415 170.150 35.180 170.290 ;
        RECT 34.415 170.105 34.705 170.150 ;
        RECT 34.860 170.090 35.180 170.150 ;
        RECT 35.780 170.290 36.100 170.350 ;
        RECT 40.840 170.290 41.160 170.350 ;
        RECT 44.520 170.290 44.840 170.350 ;
        RECT 35.780 170.150 44.840 170.290 ;
        RECT 35.780 170.090 36.100 170.150 ;
        RECT 40.840 170.090 41.160 170.150 ;
        RECT 44.520 170.090 44.840 170.150 ;
        RECT 46.820 170.290 47.140 170.350 ;
        RECT 47.295 170.290 47.585 170.335 ;
        RECT 46.820 170.150 47.585 170.290 ;
        RECT 46.820 170.090 47.140 170.150 ;
        RECT 47.295 170.105 47.585 170.150 ;
        RECT 56.020 170.090 56.340 170.350 ;
        RECT 62.920 170.290 63.240 170.350 ;
        RECT 73.055 170.290 73.345 170.335 ;
        RECT 62.920 170.150 73.345 170.290 ;
        RECT 62.920 170.090 63.240 170.150 ;
        RECT 73.055 170.105 73.345 170.150 ;
        RECT 27.515 169.950 27.805 169.995 ;
        RECT 28.880 169.950 29.200 170.010 ;
        RECT 27.515 169.810 29.200 169.950 ;
        RECT 27.515 169.765 27.805 169.810 ;
        RECT 28.880 169.750 29.200 169.810 ;
        RECT 29.340 169.950 29.660 170.010 ;
        RECT 29.340 169.810 38.310 169.950 ;
        RECT 29.340 169.750 29.660 169.810 ;
        RECT 21.995 169.470 24.280 169.610 ;
        RECT 21.995 169.425 22.285 169.470 ;
        RECT 21.060 169.270 21.380 169.330 ;
        RECT 22.070 169.270 22.210 169.425 ;
        RECT 22.440 169.410 22.760 169.470 ;
        RECT 36.700 169.410 37.020 169.670 ;
        RECT 37.620 169.410 37.940 169.670 ;
        RECT 21.060 169.130 22.210 169.270 ;
        RECT 26.135 169.270 26.425 169.315 ;
        RECT 27.040 169.270 27.360 169.330 ;
        RECT 26.135 169.130 27.360 169.270 ;
        RECT 21.060 169.070 21.380 169.130 ;
        RECT 26.135 169.085 26.425 169.130 ;
        RECT 27.040 169.070 27.360 169.130 ;
        RECT 27.500 169.070 27.820 169.330 ;
        RECT 29.340 169.270 29.660 169.330 ;
        RECT 30.275 169.270 30.565 169.315 ;
        RECT 29.340 169.130 30.565 169.270 ;
        RECT 29.340 169.070 29.660 169.130 ;
        RECT 30.275 169.085 30.565 169.130 ;
        RECT 31.180 169.070 31.500 169.330 ;
        RECT 31.655 169.270 31.945 169.315 ;
        RECT 33.480 169.270 33.800 169.330 ;
        RECT 31.655 169.130 33.800 169.270 ;
        RECT 31.655 169.085 31.945 169.130 ;
        RECT 33.480 169.070 33.800 169.130 ;
        RECT 38.170 169.280 38.310 169.810 ;
        RECT 38.540 169.750 38.860 170.010 ;
        RECT 40.380 169.950 40.700 170.010 ;
        RECT 43.615 169.950 43.905 169.995 ;
        RECT 48.660 169.950 48.980 170.010 ;
        RECT 40.380 169.810 41.530 169.950 ;
        RECT 40.380 169.750 40.700 169.810 ;
        RECT 38.630 169.610 38.770 169.750 ;
        RECT 38.630 169.470 40.150 169.610 ;
        RECT 40.010 169.325 40.150 169.470 ;
        RECT 38.515 169.280 38.805 169.325 ;
        RECT 38.170 169.095 38.805 169.280 ;
        RECT 39.935 169.095 40.225 169.325 ;
        RECT 38.170 169.080 38.770 169.095 ;
        RECT 27.590 168.930 27.730 169.070 ;
        RECT 30.720 168.930 31.040 168.990 ;
        RECT 33.035 168.930 33.325 168.975 ;
        RECT 27.590 168.790 33.325 168.930 ;
        RECT 30.720 168.730 31.040 168.790 ;
        RECT 33.035 168.745 33.325 168.790 ;
        RECT 19.220 168.590 19.540 168.650 ;
        RECT 21.075 168.590 21.365 168.635 ;
        RECT 21.980 168.590 22.300 168.650 ;
        RECT 19.220 168.450 22.300 168.590 ;
        RECT 19.220 168.390 19.540 168.450 ;
        RECT 21.075 168.405 21.365 168.450 ;
        RECT 21.980 168.390 22.300 168.450 ;
        RECT 26.595 168.590 26.885 168.635 ;
        RECT 29.355 168.590 29.645 168.635 ;
        RECT 32.115 168.590 32.405 168.635 ;
        RECT 26.595 168.450 32.405 168.590 ;
        RECT 26.595 168.405 26.885 168.450 ;
        RECT 29.355 168.405 29.645 168.450 ;
        RECT 32.115 168.405 32.405 168.450 ;
        RECT 35.780 168.590 36.100 168.650 ;
        RECT 36.255 168.590 36.545 168.635 ;
        RECT 35.780 168.450 36.545 168.590 ;
        RECT 38.630 168.590 38.770 169.080 ;
        RECT 40.840 169.070 41.160 169.330 ;
        RECT 39.015 168.930 39.305 168.975 ;
        RECT 41.390 168.930 41.530 169.810 ;
        RECT 43.615 169.810 48.980 169.950 ;
        RECT 43.615 169.765 43.905 169.810 ;
        RECT 48.660 169.750 48.980 169.810 ;
        RECT 50.960 169.950 51.280 170.010 ;
        RECT 63.855 169.950 64.145 169.995 ;
        RECT 50.960 169.810 64.145 169.950 ;
        RECT 50.960 169.750 51.280 169.810 ;
        RECT 63.855 169.765 64.145 169.810 ;
        RECT 64.760 169.750 65.080 170.010 ;
        RECT 68.915 169.950 69.205 169.995 ;
        RECT 67.150 169.810 69.205 169.950 ;
        RECT 41.760 169.610 42.080 169.670 ;
        RECT 59.700 169.610 60.020 169.670 ;
        RECT 61.080 169.610 61.400 169.670 ;
        RECT 41.760 169.470 47.050 169.610 ;
        RECT 41.760 169.410 42.080 169.470 ;
        RECT 42.220 169.070 42.540 169.330 ;
        RECT 42.770 169.315 42.910 169.470 ;
        RECT 42.695 169.085 42.985 169.315 ;
        RECT 44.060 169.070 44.380 169.330 ;
        RECT 46.910 169.315 47.050 169.470 ;
        RECT 59.700 169.470 62.230 169.610 ;
        RECT 59.700 169.410 60.020 169.470 ;
        RECT 61.080 169.410 61.400 169.470 ;
        RECT 46.835 169.085 47.125 169.315 ;
        RECT 47.755 169.270 48.045 169.315 ;
        RECT 48.200 169.270 48.520 169.330 ;
        RECT 56.480 169.270 56.800 169.330 ;
        RECT 47.755 169.130 48.520 169.270 ;
        RECT 47.755 169.085 48.045 169.130 ;
        RECT 48.200 169.070 48.520 169.130 ;
        RECT 48.750 169.130 56.800 169.270 ;
        RECT 43.615 168.930 43.905 168.975 ;
        RECT 39.015 168.790 40.610 168.930 ;
        RECT 41.390 168.790 43.905 168.930 ;
        RECT 39.015 168.745 39.305 168.790 ;
        RECT 39.935 168.590 40.225 168.635 ;
        RECT 38.630 168.450 40.225 168.590 ;
        RECT 40.470 168.590 40.610 168.790 ;
        RECT 43.615 168.745 43.905 168.790 ;
        RECT 43.140 168.590 43.460 168.650 ;
        RECT 40.470 168.450 43.460 168.590 ;
        RECT 44.150 168.590 44.290 169.070 ;
        RECT 44.535 168.930 44.825 168.975 ;
        RECT 44.980 168.930 45.300 168.990 ;
        RECT 48.750 168.930 48.890 169.130 ;
        RECT 56.480 169.070 56.800 169.130 ;
        RECT 57.860 169.070 58.180 169.330 ;
        RECT 62.090 169.315 62.230 169.470 ;
        RECT 61.555 169.085 61.845 169.315 ;
        RECT 62.015 169.085 62.305 169.315 ;
        RECT 44.535 168.790 48.890 168.930 ;
        RECT 51.420 168.930 51.740 168.990 ;
        RECT 60.635 168.930 60.925 168.975 ;
        RECT 51.420 168.790 60.925 168.930 ;
        RECT 61.630 168.930 61.770 169.085 ;
        RECT 62.920 169.070 63.240 169.330 ;
        RECT 63.380 169.070 63.700 169.330 ;
        RECT 64.850 169.315 64.990 169.750 ;
        RECT 64.750 169.085 65.040 169.315 ;
        RECT 65.220 169.070 65.540 169.330 ;
        RECT 66.600 169.270 66.920 169.330 ;
        RECT 67.150 169.315 67.290 169.810 ;
        RECT 68.915 169.765 69.205 169.810 ;
        RECT 71.200 169.950 71.520 170.010 ;
        RECT 71.675 169.950 71.965 169.995 ;
        RECT 75.340 169.950 75.660 170.010 ;
        RECT 71.200 169.810 75.660 169.950 ;
        RECT 71.200 169.750 71.520 169.810 ;
        RECT 71.675 169.765 71.965 169.810 ;
        RECT 75.340 169.750 75.660 169.810 ;
        RECT 76.260 169.750 76.580 170.010 ;
        RECT 68.440 169.610 68.760 169.670 ;
        RECT 80.875 169.610 81.165 169.655 ;
        RECT 82.700 169.610 83.020 169.670 ;
        RECT 68.440 169.470 81.165 169.610 ;
        RECT 68.440 169.410 68.760 169.470 ;
        RECT 80.875 169.425 81.165 169.470 ;
        RECT 81.870 169.470 83.020 169.610 ;
        RECT 66.405 169.130 66.920 169.270 ;
        RECT 66.600 169.070 66.920 169.130 ;
        RECT 67.075 169.085 67.365 169.315 ;
        RECT 67.520 169.120 67.840 169.380 ;
        RECT 69.820 169.270 70.140 169.330 ;
        RECT 70.755 169.270 71.045 169.315 ;
        RECT 69.820 169.130 71.045 169.270 ;
        RECT 69.820 169.070 70.140 169.130 ;
        RECT 70.755 169.085 71.045 169.130 ;
        RECT 71.215 169.270 71.505 169.315 ;
        RECT 71.660 169.270 71.980 169.330 ;
        RECT 71.215 169.130 71.980 169.270 ;
        RECT 71.215 169.085 71.505 169.130 ;
        RECT 71.660 169.070 71.980 169.130 ;
        RECT 72.135 169.270 72.425 169.315 ;
        RECT 72.580 169.270 72.900 169.330 ;
        RECT 72.135 169.130 72.900 169.270 ;
        RECT 72.135 169.085 72.425 169.130 ;
        RECT 72.580 169.070 72.900 169.130 ;
        RECT 74.420 169.270 74.740 169.330 ;
        RECT 81.870 169.315 82.010 169.470 ;
        RECT 82.700 169.410 83.020 169.470 ;
        RECT 74.420 169.130 79.250 169.270 ;
        RECT 74.420 169.070 74.740 169.130 ;
        RECT 65.695 168.930 65.985 168.975 ;
        RECT 61.630 168.790 68.670 168.930 ;
        RECT 44.535 168.745 44.825 168.790 ;
        RECT 44.980 168.730 45.300 168.790 ;
        RECT 51.420 168.730 51.740 168.790 ;
        RECT 60.635 168.745 60.925 168.790 ;
        RECT 65.695 168.745 65.985 168.790 ;
        RECT 50.960 168.590 51.280 168.650 ;
        RECT 44.150 168.450 51.280 168.590 ;
        RECT 35.780 168.390 36.100 168.450 ;
        RECT 36.255 168.405 36.545 168.450 ;
        RECT 39.935 168.405 40.225 168.450 ;
        RECT 43.140 168.390 43.460 168.450 ;
        RECT 50.960 168.390 51.280 168.450 ;
        RECT 52.800 168.590 53.120 168.650 ;
        RECT 55.115 168.590 55.405 168.635 ;
        RECT 52.800 168.450 55.405 168.590 ;
        RECT 52.800 168.390 53.120 168.450 ;
        RECT 55.115 168.405 55.405 168.450 ;
        RECT 64.760 168.590 65.080 168.650 ;
        RECT 67.995 168.590 68.285 168.635 ;
        RECT 64.760 168.450 68.285 168.590 ;
        RECT 68.530 168.590 68.670 168.790 ;
        RECT 68.900 168.730 69.220 168.990 ;
        RECT 75.355 168.930 75.645 168.975 ;
        RECT 75.800 168.930 76.120 168.990 ;
        RECT 75.355 168.790 76.120 168.930 ;
        RECT 75.355 168.745 75.645 168.790 ;
        RECT 75.800 168.730 76.120 168.790 ;
        RECT 78.100 168.930 78.420 168.990 ;
        RECT 78.575 168.930 78.865 168.975 ;
        RECT 78.100 168.790 78.865 168.930 ;
        RECT 79.110 168.930 79.250 169.130 ;
        RECT 81.795 169.085 82.085 169.315 ;
        RECT 82.240 169.070 82.560 169.330 ;
        RECT 83.635 168.930 83.925 168.975 ;
        RECT 79.110 168.790 83.925 168.930 ;
        RECT 78.100 168.730 78.420 168.790 ;
        RECT 78.575 168.745 78.865 168.790 ;
        RECT 83.635 168.745 83.925 168.790 ;
        RECT 73.500 168.590 73.820 168.650 ;
        RECT 68.530 168.450 73.820 168.590 ;
        RECT 64.760 168.390 65.080 168.450 ;
        RECT 67.995 168.405 68.285 168.450 ;
        RECT 73.500 168.390 73.820 168.450 ;
        RECT 15.930 167.770 87.230 168.250 ;
        RECT 20.140 167.570 20.460 167.630 ;
        RECT 21.535 167.570 21.825 167.615 ;
        RECT 20.140 167.430 21.825 167.570 ;
        RECT 20.140 167.370 20.460 167.430 ;
        RECT 21.535 167.385 21.825 167.430 ;
        RECT 27.040 167.370 27.360 167.630 ;
        RECT 31.180 167.570 31.500 167.630 ;
        RECT 37.620 167.570 37.940 167.630 ;
        RECT 31.180 167.430 37.940 167.570 ;
        RECT 31.180 167.370 31.500 167.430 ;
        RECT 37.620 167.370 37.940 167.430 ;
        RECT 45.440 167.370 45.760 167.630 ;
        RECT 46.360 167.370 46.680 167.630 ;
        RECT 50.500 167.570 50.820 167.630 ;
        RECT 50.975 167.570 51.265 167.615 ;
        RECT 53.260 167.570 53.580 167.630 ;
        RECT 59.715 167.570 60.005 167.615 ;
        RECT 66.140 167.570 66.460 167.630 ;
        RECT 50.500 167.430 51.265 167.570 ;
        RECT 50.500 167.370 50.820 167.430 ;
        RECT 50.975 167.385 51.265 167.430 ;
        RECT 51.970 167.430 60.005 167.570 ;
        RECT 36.700 167.230 37.020 167.290 ;
        RECT 24.370 167.090 37.020 167.230 ;
        RECT 21.520 166.890 21.840 166.950 ;
        RECT 24.370 166.935 24.510 167.090 ;
        RECT 36.700 167.030 37.020 167.090 ;
        RECT 21.995 166.890 22.285 166.935 ;
        RECT 21.520 166.750 22.285 166.890 ;
        RECT 21.520 166.690 21.840 166.750 ;
        RECT 21.995 166.705 22.285 166.750 ;
        RECT 24.295 166.705 24.585 166.935 ;
        RECT 25.660 166.690 25.980 166.950 ;
        RECT 26.120 166.690 26.440 166.950 ;
        RECT 41.760 166.890 42.080 166.950 ;
        RECT 51.970 166.935 52.110 167.430 ;
        RECT 53.260 167.370 53.580 167.430 ;
        RECT 59.715 167.385 60.005 167.430 ;
        RECT 64.390 167.430 66.460 167.570 ;
        RECT 52.340 167.230 52.660 167.290 ;
        RECT 58.780 167.230 59.100 167.290 ;
        RECT 64.390 167.275 64.530 167.430 ;
        RECT 66.140 167.370 66.460 167.430 ;
        RECT 67.075 167.570 67.365 167.615 ;
        RECT 81.780 167.570 82.100 167.630 ;
        RECT 67.075 167.430 82.100 167.570 ;
        RECT 67.075 167.385 67.365 167.430 ;
        RECT 81.780 167.370 82.100 167.430 ;
        RECT 82.715 167.570 83.005 167.615 ;
        RECT 84.080 167.570 84.400 167.630 ;
        RECT 82.715 167.430 84.400 167.570 ;
        RECT 82.715 167.385 83.005 167.430 ;
        RECT 84.080 167.370 84.400 167.430 ;
        RECT 52.340 167.090 53.490 167.230 ;
        RECT 52.340 167.030 52.660 167.090 ;
        RECT 46.080 166.890 46.370 166.935 ;
        RECT 41.760 166.750 46.370 166.890 ;
        RECT 41.760 166.690 42.080 166.750 ;
        RECT 46.080 166.705 46.370 166.750 ;
        RECT 51.895 166.705 52.185 166.935 ;
        RECT 52.800 166.690 53.120 166.950 ;
        RECT 53.350 166.935 53.490 167.090 ;
        RECT 55.650 167.090 57.170 167.230 ;
        RECT 53.275 166.705 53.565 166.935 ;
        RECT 53.720 166.890 54.040 166.950 ;
        RECT 54.195 166.890 54.485 166.935 ;
        RECT 53.720 166.750 54.485 166.890 ;
        RECT 53.720 166.690 54.040 166.750 ;
        RECT 54.195 166.705 54.485 166.750 ;
        RECT 55.100 166.690 55.420 166.950 ;
        RECT 55.650 166.935 55.790 167.090 ;
        RECT 57.030 166.950 57.170 167.090 ;
        RECT 58.780 167.090 61.310 167.230 ;
        RECT 58.780 167.030 59.100 167.090 ;
        RECT 55.575 166.705 55.865 166.935 ;
        RECT 56.020 166.690 56.340 166.950 ;
        RECT 56.940 166.890 57.260 166.950 ;
        RECT 57.875 166.890 58.165 166.935 ;
        RECT 56.940 166.750 58.165 166.890 ;
        RECT 56.940 166.690 57.260 166.750 ;
        RECT 57.875 166.705 58.165 166.750 ;
        RECT 58.320 166.890 58.640 166.950 ;
        RECT 61.170 166.935 61.310 167.090 ;
        RECT 64.315 167.045 64.605 167.275 ;
        RECT 64.760 167.230 65.080 167.290 ;
        RECT 65.235 167.230 65.525 167.275 ;
        RECT 64.760 167.090 65.525 167.230 ;
        RECT 64.760 167.030 65.080 167.090 ;
        RECT 65.235 167.045 65.525 167.090 ;
        RECT 67.980 167.230 68.300 167.290 ;
        RECT 71.200 167.230 71.520 167.290 ;
        RECT 75.800 167.230 76.120 167.290 ;
        RECT 83.635 167.230 83.925 167.275 ;
        RECT 85.460 167.230 85.780 167.290 ;
        RECT 67.980 167.090 70.510 167.230 ;
        RECT 60.175 166.890 60.465 166.935 ;
        RECT 58.320 166.750 60.465 166.890 ;
        RECT 58.320 166.690 58.640 166.750 ;
        RECT 60.175 166.705 60.465 166.750 ;
        RECT 61.095 166.705 61.385 166.935 ;
        RECT 65.675 166.815 65.965 167.045 ;
        RECT 67.980 167.030 68.300 167.090 ;
        RECT 21.060 166.350 21.380 166.610 ;
        RECT 30.720 166.550 31.040 166.610 ;
        RECT 48.675 166.550 48.965 166.595 ;
        RECT 51.420 166.550 51.740 166.610 ;
        RECT 30.720 166.410 51.740 166.550 ;
        RECT 30.720 166.350 31.040 166.410 ;
        RECT 48.675 166.365 48.965 166.410 ;
        RECT 51.420 166.350 51.740 166.410 ;
        RECT 52.355 166.550 52.645 166.595 ;
        RECT 54.640 166.550 54.960 166.610 ;
        RECT 52.355 166.410 54.960 166.550 ;
        RECT 56.110 166.550 56.250 166.690 ;
        RECT 65.770 166.610 65.910 166.815 ;
        RECT 66.155 166.705 66.445 166.935 ;
        RECT 68.915 166.890 69.205 166.935 ;
        RECT 69.820 166.890 70.140 166.950 ;
        RECT 70.370 166.935 70.510 167.090 ;
        RECT 71.200 167.090 75.570 167.230 ;
        RECT 71.200 167.030 71.520 167.090 ;
        RECT 68.915 166.750 70.140 166.890 ;
        RECT 68.915 166.705 69.205 166.750 ;
        RECT 60.635 166.550 60.925 166.595 ;
        RECT 56.110 166.410 60.925 166.550 ;
        RECT 52.355 166.365 52.645 166.410 ;
        RECT 54.640 166.350 54.960 166.410 ;
        RECT 60.635 166.365 60.925 166.410 ;
        RECT 65.680 166.350 66.000 166.610 ;
        RECT 66.230 166.550 66.370 166.705 ;
        RECT 69.820 166.690 70.140 166.750 ;
        RECT 70.295 166.705 70.585 166.935 ;
        RECT 71.675 166.890 71.965 166.935 ;
        RECT 72.120 166.890 72.440 166.950 ;
        RECT 71.675 166.750 72.440 166.890 ;
        RECT 71.675 166.705 71.965 166.750 ;
        RECT 72.120 166.690 72.440 166.750 ;
        RECT 72.595 166.890 72.885 166.935 ;
        RECT 73.040 166.890 73.360 166.950 ;
        RECT 72.595 166.750 73.360 166.890 ;
        RECT 72.595 166.705 72.885 166.750 ;
        RECT 73.040 166.690 73.360 166.750 ;
        RECT 73.960 166.690 74.280 166.950 ;
        RECT 74.420 166.890 74.740 166.950 ;
        RECT 75.430 166.935 75.570 167.090 ;
        RECT 75.800 167.090 85.780 167.230 ;
        RECT 75.800 167.030 76.120 167.090 ;
        RECT 83.635 167.045 83.925 167.090 ;
        RECT 85.460 167.030 85.780 167.090 ;
        RECT 74.895 166.890 75.185 166.935 ;
        RECT 74.420 166.750 75.185 166.890 ;
        RECT 74.420 166.690 74.740 166.750 ;
        RECT 74.895 166.705 75.185 166.750 ;
        RECT 75.355 166.705 75.645 166.935 ;
        RECT 76.260 166.690 76.580 166.950 ;
        RECT 84.095 166.890 84.385 166.935 ;
        RECT 80.030 166.750 84.385 166.890 ;
        RECT 80.030 166.610 80.170 166.750 ;
        RECT 84.095 166.705 84.385 166.750 ;
        RECT 78.100 166.550 78.420 166.610 ;
        RECT 66.230 166.410 78.420 166.550 ;
        RECT 78.100 166.350 78.420 166.410 ;
        RECT 78.560 166.350 78.880 166.610 ;
        RECT 79.940 166.350 80.260 166.610 ;
        RECT 80.860 166.550 81.180 166.610 ;
        RECT 82.240 166.550 82.560 166.610 ;
        RECT 80.860 166.410 82.560 166.550 ;
        RECT 80.860 166.350 81.180 166.410 ;
        RECT 82.240 166.350 82.560 166.410 ;
        RECT 48.215 166.210 48.505 166.255 ;
        RECT 57.415 166.210 57.705 166.255 ;
        RECT 48.215 166.070 57.705 166.210 ;
        RECT 48.215 166.025 48.505 166.070 ;
        RECT 57.415 166.025 57.705 166.070 ;
        RECT 63.380 166.210 63.700 166.270 ;
        RECT 64.315 166.210 64.605 166.255 ;
        RECT 63.380 166.070 64.605 166.210 ;
        RECT 65.770 166.210 65.910 166.350 ;
        RECT 67.520 166.210 67.840 166.270 ;
        RECT 65.770 166.070 67.840 166.210 ;
        RECT 63.380 166.010 63.700 166.070 ;
        RECT 64.315 166.025 64.605 166.070 ;
        RECT 67.520 166.010 67.840 166.070 ;
        RECT 69.820 166.010 70.140 166.270 ;
        RECT 70.740 166.210 71.060 166.270 ;
        RECT 71.215 166.210 71.505 166.255 ;
        RECT 70.740 166.070 71.505 166.210 ;
        RECT 70.740 166.010 71.060 166.070 ;
        RECT 71.215 166.025 71.505 166.070 ;
        RECT 72.580 166.210 72.900 166.270 ;
        RECT 76.260 166.210 76.580 166.270 ;
        RECT 72.580 166.070 76.580 166.210 ;
        RECT 72.580 166.010 72.900 166.070 ;
        RECT 76.260 166.010 76.580 166.070 ;
        RECT 77.180 166.010 77.500 166.270 ;
        RECT 80.415 166.210 80.705 166.255 ;
        RECT 83.160 166.210 83.480 166.270 ;
        RECT 85.015 166.210 85.305 166.255 ;
        RECT 80.415 166.070 85.305 166.210 ;
        RECT 80.415 166.025 80.705 166.070 ;
        RECT 83.160 166.010 83.480 166.070 ;
        RECT 85.015 166.025 85.305 166.070 ;
        RECT 23.835 165.870 24.125 165.915 ;
        RECT 24.755 165.870 25.045 165.915 ;
        RECT 23.835 165.730 25.045 165.870 ;
        RECT 23.835 165.685 24.125 165.730 ;
        RECT 24.755 165.685 25.045 165.730 ;
        RECT 27.960 165.870 28.280 165.930 ;
        RECT 48.660 165.870 48.980 165.930 ;
        RECT 27.960 165.730 48.980 165.870 ;
        RECT 27.960 165.670 28.280 165.730 ;
        RECT 48.660 165.670 48.980 165.730 ;
        RECT 73.040 165.870 73.360 165.930 ;
        RECT 75.340 165.870 75.660 165.930 ;
        RECT 73.040 165.730 75.660 165.870 ;
        RECT 73.040 165.670 73.360 165.730 ;
        RECT 75.340 165.670 75.660 165.730 ;
        RECT 79.480 165.870 79.800 165.930 ;
        RECT 80.860 165.870 81.180 165.930 ;
        RECT 79.480 165.730 81.180 165.870 ;
        RECT 79.480 165.670 79.800 165.730 ;
        RECT 80.860 165.670 81.180 165.730 ;
        RECT 81.780 165.670 82.100 165.930 ;
        RECT 82.240 165.870 82.560 165.930 ;
        RECT 82.715 165.870 83.005 165.915 ;
        RECT 84.540 165.870 84.860 165.930 ;
        RECT 82.240 165.730 84.860 165.870 ;
        RECT 82.240 165.670 82.560 165.730 ;
        RECT 82.715 165.685 83.005 165.730 ;
        RECT 84.540 165.670 84.860 165.730 ;
        RECT 15.930 165.050 87.230 165.530 ;
        RECT 25.660 164.850 25.980 164.910 ;
        RECT 27.975 164.850 28.265 164.895 ;
        RECT 25.660 164.710 28.265 164.850 ;
        RECT 25.660 164.650 25.980 164.710 ;
        RECT 27.975 164.665 28.265 164.710 ;
        RECT 32.115 164.850 32.405 164.895 ;
        RECT 33.480 164.850 33.800 164.910 ;
        RECT 32.115 164.710 33.800 164.850 ;
        RECT 32.115 164.665 32.405 164.710 ;
        RECT 21.060 163.970 21.380 164.230 ;
        RECT 28.050 164.170 28.190 164.665 ;
        RECT 33.480 164.650 33.800 164.710 ;
        RECT 41.300 164.650 41.620 164.910 ;
        RECT 43.140 164.850 43.460 164.910 ;
        RECT 45.440 164.850 45.760 164.910 ;
        RECT 43.140 164.710 45.760 164.850 ;
        RECT 43.140 164.650 43.460 164.710 ;
        RECT 45.440 164.650 45.760 164.710 ;
        RECT 53.720 164.850 54.040 164.910 ;
        RECT 55.115 164.850 55.405 164.895 ;
        RECT 53.720 164.710 55.405 164.850 ;
        RECT 53.720 164.650 54.040 164.710 ;
        RECT 55.115 164.665 55.405 164.710 ;
        RECT 57.415 164.850 57.705 164.895 ;
        RECT 58.320 164.850 58.640 164.910 ;
        RECT 57.415 164.710 58.640 164.850 ;
        RECT 57.415 164.665 57.705 164.710 ;
        RECT 58.320 164.650 58.640 164.710 ;
        RECT 69.375 164.850 69.665 164.895 ;
        RECT 70.280 164.850 70.600 164.910 ;
        RECT 69.375 164.710 70.600 164.850 ;
        RECT 69.375 164.665 69.665 164.710 ;
        RECT 70.280 164.650 70.600 164.710 ;
        RECT 70.740 164.850 71.060 164.910 ;
        RECT 72.580 164.850 72.900 164.910 ;
        RECT 73.055 164.850 73.345 164.895 ;
        RECT 70.740 164.710 72.350 164.850 ;
        RECT 70.740 164.650 71.060 164.710 ;
        RECT 33.035 164.325 33.325 164.555 ;
        RECT 29.815 164.170 30.105 164.215 ;
        RECT 33.110 164.170 33.250 164.325 ;
        RECT 28.050 164.030 29.570 164.170 ;
        RECT 20.140 163.830 20.460 163.890 ;
        RECT 21.995 163.830 22.285 163.875 ;
        RECT 20.140 163.690 22.285 163.830 ;
        RECT 20.140 163.630 20.460 163.690 ;
        RECT 21.995 163.645 22.285 163.690 ;
        RECT 27.515 163.645 27.805 163.875 ;
        RECT 27.590 163.490 27.730 163.645 ;
        RECT 28.420 163.630 28.740 163.890 ;
        RECT 29.430 163.875 29.570 164.030 ;
        RECT 29.815 164.030 33.250 164.170 ;
        RECT 36.255 164.170 36.545 164.215 ;
        RECT 36.700 164.170 37.020 164.230 ;
        RECT 36.255 164.030 37.020 164.170 ;
        RECT 29.815 163.985 30.105 164.030 ;
        RECT 36.255 163.985 36.545 164.030 ;
        RECT 36.700 163.970 37.020 164.030 ;
        RECT 40.380 164.170 40.700 164.230 ;
        RECT 46.820 164.170 47.140 164.230 ;
        RECT 40.380 164.030 47.140 164.170 ;
        RECT 40.380 163.970 40.700 164.030 ;
        RECT 29.355 163.645 29.645 163.875 ;
        RECT 30.735 163.645 31.025 163.875 ;
        RECT 31.195 163.830 31.485 163.875 ;
        RECT 32.560 163.830 32.880 163.890 ;
        RECT 31.195 163.690 32.880 163.830 ;
        RECT 31.195 163.645 31.485 163.690 ;
        RECT 29.800 163.490 30.120 163.550 ;
        RECT 27.590 163.350 30.120 163.490 ;
        RECT 30.810 163.490 30.950 163.645 ;
        RECT 32.560 163.630 32.880 163.690 ;
        RECT 33.480 163.830 33.800 163.890 ;
        RECT 37.175 163.830 37.465 163.875 ;
        RECT 33.480 163.690 37.465 163.830 ;
        RECT 33.480 163.630 33.800 163.690 ;
        RECT 37.175 163.645 37.465 163.690 ;
        RECT 38.080 163.630 38.400 163.890 ;
        RECT 42.770 163.875 42.910 164.030 ;
        RECT 46.820 163.970 47.140 164.030 ;
        RECT 56.480 163.970 56.800 164.230 ;
        RECT 63.840 164.170 64.160 164.230 ;
        RECT 57.490 164.030 64.160 164.170 ;
        RECT 42.235 163.645 42.525 163.875 ;
        RECT 42.695 163.645 42.985 163.875 ;
        RECT 36.240 163.490 36.560 163.550 ;
        RECT 30.810 163.350 36.560 163.490 ;
        RECT 42.310 163.490 42.450 163.645 ;
        RECT 43.600 163.630 43.920 163.890 ;
        RECT 44.075 163.830 44.365 163.875 ;
        RECT 49.580 163.830 49.900 163.890 ;
        RECT 44.075 163.690 49.900 163.830 ;
        RECT 44.075 163.645 44.365 163.690 ;
        RECT 49.580 163.630 49.900 163.690 ;
        RECT 51.880 163.830 52.200 163.890 ;
        RECT 57.490 163.830 57.630 164.030 ;
        RECT 63.840 163.970 64.160 164.030 ;
        RECT 51.880 163.690 57.630 163.830 ;
        RECT 51.880 163.630 52.200 163.690 ;
        RECT 57.860 163.630 58.180 163.890 ;
        RECT 72.210 163.875 72.350 164.710 ;
        RECT 72.580 164.710 73.345 164.850 ;
        RECT 72.580 164.650 72.900 164.710 ;
        RECT 73.055 164.665 73.345 164.710 ;
        RECT 73.960 164.850 74.280 164.910 ;
        RECT 75.340 164.850 75.660 164.910 ;
        RECT 73.960 164.710 75.660 164.850 ;
        RECT 73.960 164.650 74.280 164.710 ;
        RECT 75.340 164.650 75.660 164.710 ;
        RECT 73.500 164.510 73.820 164.570 ;
        RECT 77.195 164.510 77.485 164.555 ;
        RECT 73.500 164.370 77.485 164.510 ;
        RECT 73.500 164.310 73.820 164.370 ;
        RECT 77.195 164.325 77.485 164.370 ;
        RECT 74.420 164.170 74.740 164.230 ;
        RECT 75.815 164.170 76.105 164.215 ;
        RECT 74.420 164.030 76.105 164.170 ;
        RECT 74.420 163.970 74.740 164.030 ;
        RECT 75.815 163.985 76.105 164.030 ;
        RECT 78.100 163.970 78.420 164.230 ;
        RECT 79.110 164.030 83.390 164.170 ;
        RECT 72.135 163.645 72.425 163.875 ;
        RECT 72.580 163.830 72.900 163.890 ;
        RECT 73.055 163.830 73.345 163.875 ;
        RECT 72.580 163.690 73.345 163.830 ;
        RECT 72.580 163.630 72.900 163.690 ;
        RECT 73.055 163.645 73.345 163.690 ;
        RECT 73.960 163.630 74.280 163.890 ;
        RECT 52.800 163.490 53.120 163.550 ;
        RECT 42.310 163.350 61.770 163.490 ;
        RECT 29.800 163.290 30.120 163.350 ;
        RECT 36.240 163.290 36.560 163.350 ;
        RECT 52.800 163.290 53.120 163.350 ;
        RECT 61.630 163.210 61.770 163.350 ;
        RECT 69.820 163.290 70.140 163.550 ;
        RECT 74.510 163.490 74.650 163.970 ;
        RECT 75.355 163.830 75.645 163.875 ;
        RECT 76.720 163.830 77.040 163.890 ;
        RECT 79.110 163.875 79.250 164.030 ;
        RECT 83.250 163.890 83.390 164.030 ;
        RECT 75.355 163.690 77.040 163.830 ;
        RECT 75.355 163.645 75.645 163.690 ;
        RECT 76.720 163.630 77.040 163.690 ;
        RECT 79.035 163.645 79.325 163.875 ;
        RECT 79.955 163.830 80.245 163.875 ;
        RECT 80.400 163.830 80.720 163.890 ;
        RECT 79.955 163.690 80.720 163.830 ;
        RECT 79.955 163.645 80.245 163.690 ;
        RECT 80.400 163.630 80.720 163.690 ;
        RECT 80.875 163.830 81.165 163.875 ;
        RECT 82.700 163.830 83.020 163.890 ;
        RECT 80.875 163.690 83.020 163.830 ;
        RECT 80.875 163.645 81.165 163.690 ;
        RECT 82.700 163.630 83.020 163.690 ;
        RECT 83.160 163.630 83.480 163.890 ;
        RECT 84.095 163.830 84.385 163.875 ;
        RECT 84.540 163.830 84.860 163.890 ;
        RECT 84.095 163.690 84.860 163.830 ;
        RECT 84.095 163.645 84.385 163.690 ;
        RECT 84.540 163.630 84.860 163.690 ;
        RECT 85.015 163.645 85.305 163.875 ;
        RECT 71.750 163.350 74.650 163.490 ;
        RECT 78.560 163.490 78.880 163.550 ;
        RECT 85.090 163.490 85.230 163.645 ;
        RECT 78.560 163.350 85.230 163.490 ;
        RECT 21.520 162.950 21.840 163.210 ;
        RECT 23.835 163.150 24.125 163.195 ;
        RECT 26.120 163.150 26.440 163.210 ;
        RECT 23.835 163.010 26.440 163.150 ;
        RECT 23.835 162.965 24.125 163.010 ;
        RECT 26.120 162.950 26.440 163.010 ;
        RECT 33.940 163.150 34.260 163.210 ;
        RECT 34.875 163.150 35.165 163.195 ;
        RECT 33.940 163.010 35.165 163.150 ;
        RECT 33.940 162.950 34.260 163.010 ;
        RECT 34.875 162.965 35.165 163.010 ;
        RECT 35.335 163.150 35.625 163.195 ;
        RECT 36.700 163.150 37.020 163.210 ;
        RECT 37.175 163.150 37.465 163.195 ;
        RECT 35.335 163.010 37.465 163.150 ;
        RECT 35.335 162.965 35.625 163.010 ;
        RECT 36.700 162.950 37.020 163.010 ;
        RECT 37.175 162.965 37.465 163.010 ;
        RECT 47.740 163.150 48.060 163.210 ;
        RECT 50.040 163.150 50.360 163.210 ;
        RECT 51.420 163.150 51.740 163.210 ;
        RECT 61.080 163.150 61.400 163.210 ;
        RECT 47.740 163.010 61.400 163.150 ;
        RECT 47.740 162.950 48.060 163.010 ;
        RECT 50.040 162.950 50.360 163.010 ;
        RECT 51.420 162.950 51.740 163.010 ;
        RECT 61.080 162.950 61.400 163.010 ;
        RECT 61.540 163.150 61.860 163.210 ;
        RECT 71.750 163.195 71.890 163.350 ;
        RECT 78.560 163.290 78.880 163.350 ;
        RECT 70.835 163.150 71.125 163.195 ;
        RECT 61.540 163.010 71.125 163.150 ;
        RECT 61.540 162.950 61.860 163.010 ;
        RECT 70.835 162.965 71.125 163.010 ;
        RECT 71.675 162.965 71.965 163.195 ;
        RECT 74.880 162.950 75.200 163.210 ;
        RECT 79.020 163.150 79.340 163.210 ;
        RECT 82.715 163.150 83.005 163.195 ;
        RECT 79.020 163.010 83.005 163.150 ;
        RECT 79.020 162.950 79.340 163.010 ;
        RECT 82.715 162.965 83.005 163.010 ;
        RECT 15.930 162.330 87.230 162.810 ;
        RECT 20.600 162.130 20.920 162.190 ;
        RECT 22.440 162.130 22.760 162.190 ;
        RECT 20.600 161.990 32.330 162.130 ;
        RECT 20.600 161.930 20.920 161.990 ;
        RECT 22.440 161.930 22.760 161.990 ;
        RECT 28.420 161.790 28.740 161.850 ;
        RECT 32.190 161.790 32.330 161.990 ;
        RECT 32.560 161.930 32.880 162.190 ;
        RECT 34.875 162.130 35.165 162.175 ;
        RECT 36.700 162.130 37.020 162.190 ;
        RECT 34.875 161.990 37.020 162.130 ;
        RECT 34.875 161.945 35.165 161.990 ;
        RECT 36.700 161.930 37.020 161.990 ;
        RECT 42.235 162.130 42.525 162.175 ;
        RECT 43.600 162.130 43.920 162.190 ;
        RECT 42.235 161.990 43.920 162.130 ;
        RECT 42.235 161.945 42.525 161.990 ;
        RECT 43.600 161.930 43.920 161.990 ;
        RECT 44.060 162.130 44.380 162.190 ;
        RECT 44.060 161.990 48.430 162.130 ;
        RECT 44.060 161.930 44.380 161.990 ;
        RECT 37.620 161.790 37.940 161.850 ;
        RECT 38.555 161.790 38.845 161.835 ;
        RECT 45.440 161.790 45.760 161.850 ;
        RECT 28.420 161.650 30.950 161.790 ;
        RECT 32.190 161.650 37.390 161.790 ;
        RECT 28.420 161.590 28.740 161.650 ;
        RECT 18.775 161.265 19.065 161.495 ;
        RECT 18.850 161.110 18.990 161.265 ;
        RECT 19.680 161.250 20.000 161.510 ;
        RECT 28.970 161.495 29.110 161.650 ;
        RECT 21.995 161.450 22.285 161.495 ;
        RECT 28.895 161.450 29.185 161.495 ;
        RECT 21.995 161.310 29.185 161.450 ;
        RECT 21.995 161.265 22.285 161.310 ;
        RECT 28.895 161.265 29.185 161.310 ;
        RECT 29.340 161.250 29.660 161.510 ;
        RECT 29.800 161.450 30.120 161.510 ;
        RECT 30.810 161.495 30.950 161.650 ;
        RECT 30.275 161.450 30.565 161.495 ;
        RECT 29.800 161.310 30.565 161.450 ;
        RECT 29.800 161.250 30.120 161.310 ;
        RECT 30.275 161.265 30.565 161.310 ;
        RECT 30.735 161.265 31.025 161.495 ;
        RECT 33.940 161.450 34.260 161.510 ;
        RECT 34.415 161.450 34.705 161.495 ;
        RECT 36.240 161.450 36.560 161.510 ;
        RECT 33.940 161.310 36.560 161.450 ;
        RECT 37.250 161.450 37.390 161.650 ;
        RECT 37.620 161.650 44.750 161.790 ;
        RECT 37.620 161.590 37.940 161.650 ;
        RECT 38.555 161.605 38.845 161.650 ;
        RECT 39.475 161.450 39.765 161.495 ;
        RECT 40.380 161.450 40.700 161.510 ;
        RECT 37.250 161.310 39.230 161.450 ;
        RECT 30.350 161.110 30.490 161.265 ;
        RECT 33.940 161.250 34.260 161.310 ;
        RECT 34.415 161.265 34.705 161.310 ;
        RECT 36.240 161.250 36.560 161.310 ;
        RECT 35.795 161.110 36.085 161.155 ;
        RECT 36.700 161.110 37.020 161.170 ;
        RECT 38.080 161.110 38.400 161.170 ;
        RECT 18.850 160.970 21.290 161.110 ;
        RECT 30.350 160.970 32.330 161.110 ;
        RECT 17.840 160.570 18.160 160.830 ;
        RECT 21.150 160.815 21.290 160.970 ;
        RECT 21.075 160.585 21.365 160.815 ;
        RECT 32.190 160.770 32.330 160.970 ;
        RECT 35.795 160.970 38.400 161.110 ;
        RECT 39.090 161.110 39.230 161.310 ;
        RECT 39.475 161.310 40.700 161.450 ;
        RECT 39.475 161.265 39.765 161.310 ;
        RECT 40.380 161.250 40.700 161.310 ;
        RECT 40.840 161.450 41.160 161.510 ;
        RECT 44.610 161.495 44.750 161.650 ;
        RECT 45.440 161.650 46.590 161.790 ;
        RECT 45.440 161.590 45.760 161.650 ;
        RECT 43.155 161.450 43.445 161.495 ;
        RECT 40.840 161.310 43.445 161.450 ;
        RECT 40.840 161.250 41.160 161.310 ;
        RECT 43.155 161.265 43.445 161.310 ;
        RECT 44.535 161.265 44.825 161.495 ;
        RECT 44.980 161.250 45.300 161.510 ;
        RECT 45.900 161.450 46.220 161.510 ;
        RECT 46.450 161.495 46.590 161.650 ;
        RECT 47.740 161.590 48.060 161.850 ;
        RECT 48.290 161.835 48.430 161.990 ;
        RECT 49.580 161.930 49.900 162.190 ;
        RECT 50.590 161.990 52.570 162.130 ;
        RECT 48.215 161.790 48.505 161.835 ;
        RECT 50.590 161.790 50.730 161.990 ;
        RECT 48.215 161.650 50.730 161.790 ;
        RECT 48.215 161.605 48.505 161.650 ;
        RECT 50.960 161.590 51.280 161.850 ;
        RECT 51.420 161.590 51.740 161.850 ;
        RECT 52.430 161.790 52.570 161.990 ;
        RECT 52.800 161.930 53.120 162.190 ;
        RECT 54.180 162.130 54.500 162.190 ;
        RECT 61.080 162.130 61.400 162.190 ;
        RECT 63.855 162.130 64.145 162.175 ;
        RECT 54.180 161.990 60.850 162.130 ;
        RECT 54.180 161.930 54.500 161.990 ;
        RECT 58.320 161.790 58.640 161.850 ;
        RECT 60.710 161.790 60.850 161.990 ;
        RECT 61.080 161.990 64.145 162.130 ;
        RECT 61.080 161.930 61.400 161.990 ;
        RECT 63.855 161.945 64.145 161.990 ;
        RECT 65.680 162.130 66.000 162.190 ;
        RECT 67.995 162.130 68.285 162.175 ;
        RECT 65.680 161.990 68.285 162.130 ;
        RECT 65.680 161.930 66.000 161.990 ;
        RECT 67.995 161.945 68.285 161.990 ;
        RECT 73.040 161.930 73.360 162.190 ;
        RECT 75.340 161.930 75.660 162.190 ;
        RECT 83.160 161.930 83.480 162.190 ;
        RECT 62.460 161.790 62.780 161.850 ;
        RECT 69.820 161.790 70.140 161.850 ;
        RECT 71.200 161.790 71.520 161.850 ;
        RECT 52.430 161.650 58.640 161.790 ;
        RECT 58.320 161.590 58.640 161.650 ;
        RECT 58.870 161.650 60.390 161.790 ;
        RECT 60.710 161.650 62.230 161.790 ;
        RECT 45.530 161.310 46.220 161.450 ;
        RECT 43.600 161.110 43.920 161.170 ;
        RECT 44.075 161.110 44.365 161.155 ;
        RECT 45.530 161.110 45.670 161.310 ;
        RECT 45.900 161.250 46.220 161.310 ;
        RECT 46.375 161.265 46.665 161.495 ;
        RECT 47.065 161.265 47.355 161.495 ;
        RECT 48.675 161.450 48.965 161.495 ;
        RECT 50.055 161.450 50.345 161.495 ;
        RECT 48.675 161.310 50.345 161.450 ;
        RECT 48.675 161.265 48.965 161.310 ;
        RECT 50.055 161.265 50.345 161.310 ;
        RECT 51.895 161.450 52.185 161.495 ;
        RECT 54.180 161.450 54.500 161.510 ;
        RECT 58.870 161.495 59.010 161.650 ;
        RECT 51.895 161.310 54.500 161.450 ;
        RECT 51.895 161.265 52.185 161.310 ;
        RECT 47.140 161.110 47.280 161.265 ;
        RECT 39.090 160.970 44.365 161.110 ;
        RECT 35.795 160.925 36.085 160.970 ;
        RECT 36.700 160.910 37.020 160.970 ;
        RECT 38.080 160.910 38.400 160.970 ;
        RECT 43.600 160.910 43.920 160.970 ;
        RECT 44.075 160.925 44.365 160.970 ;
        RECT 45.070 160.970 45.670 161.110 ;
        RECT 46.155 160.970 47.280 161.110 ;
        RECT 47.740 161.110 48.060 161.170 ;
        RECT 48.750 161.110 48.890 161.265 ;
        RECT 47.740 160.970 48.890 161.110 ;
        RECT 50.130 161.110 50.270 161.265 ;
        RECT 54.180 161.250 54.500 161.310 ;
        RECT 58.795 161.265 59.085 161.495 ;
        RECT 59.715 161.265 60.005 161.495 ;
        RECT 56.020 161.110 56.340 161.170 ;
        RECT 58.870 161.110 59.010 161.265 ;
        RECT 50.130 160.970 59.010 161.110 ;
        RECT 38.540 160.770 38.860 160.830 ;
        RECT 32.190 160.630 38.860 160.770 ;
        RECT 38.540 160.570 38.860 160.630 ;
        RECT 40.395 160.770 40.685 160.815 ;
        RECT 41.300 160.770 41.620 160.830 ;
        RECT 40.395 160.630 41.620 160.770 ;
        RECT 40.395 160.585 40.685 160.630 ;
        RECT 41.300 160.570 41.620 160.630 ;
        RECT 20.140 160.230 20.460 160.490 ;
        RECT 31.655 160.430 31.945 160.475 ;
        RECT 45.070 160.430 45.210 160.970 ;
        RECT 46.155 160.830 46.295 160.970 ;
        RECT 47.740 160.910 48.060 160.970 ;
        RECT 56.020 160.910 56.340 160.970 ;
        RECT 45.900 160.630 46.295 160.830 ;
        RECT 50.960 160.770 51.280 160.830 ;
        RECT 53.260 160.770 53.580 160.830 ;
        RECT 56.480 160.770 56.800 160.830 ;
        RECT 59.790 160.770 59.930 161.265 ;
        RECT 60.250 161.170 60.390 161.650 ;
        RECT 61.080 161.250 61.400 161.510 ;
        RECT 62.090 161.495 62.230 161.650 ;
        RECT 62.460 161.650 64.990 161.790 ;
        RECT 62.460 161.590 62.780 161.650 ;
        RECT 64.850 161.495 64.990 161.650 ;
        RECT 69.820 161.650 71.520 161.790 ;
        RECT 69.820 161.590 70.140 161.650 ;
        RECT 62.015 161.265 62.305 161.495 ;
        RECT 63.395 161.450 63.685 161.495 ;
        RECT 62.550 161.310 63.685 161.450 ;
        RECT 60.160 161.110 60.480 161.170 ;
        RECT 62.550 161.110 62.690 161.310 ;
        RECT 63.395 161.265 63.685 161.310 ;
        RECT 64.775 161.265 65.065 161.495 ;
        RECT 68.440 161.450 68.760 161.510 ;
        RECT 68.915 161.450 69.205 161.495 ;
        RECT 68.440 161.310 69.205 161.450 ;
        RECT 68.440 161.250 68.760 161.310 ;
        RECT 68.915 161.265 69.205 161.310 ;
        RECT 69.375 161.450 69.665 161.495 ;
        RECT 70.280 161.450 70.600 161.510 ;
        RECT 70.830 161.495 70.970 161.650 ;
        RECT 71.200 161.590 71.520 161.650 ;
        RECT 69.375 161.310 70.600 161.450 ;
        RECT 69.375 161.265 69.665 161.310 ;
        RECT 70.280 161.250 70.600 161.310 ;
        RECT 70.755 161.265 71.045 161.495 ;
        RECT 72.365 161.450 72.655 161.665 ;
        RECT 73.500 161.590 73.820 161.850 ;
        RECT 74.420 161.835 74.740 161.850 ;
        RECT 74.420 161.605 74.805 161.835 ;
        RECT 76.735 161.790 77.025 161.835 ;
        RECT 81.320 161.790 81.640 161.850 ;
        RECT 76.735 161.650 81.640 161.790 ;
        RECT 76.735 161.605 77.025 161.650 ;
        RECT 74.420 161.590 74.740 161.605 ;
        RECT 81.320 161.590 81.640 161.650 ;
        RECT 71.290 161.435 72.655 161.450 ;
        RECT 71.290 161.310 72.580 161.435 ;
        RECT 60.160 160.970 62.690 161.110 ;
        RECT 62.920 161.110 63.240 161.170 ;
        RECT 65.695 161.110 65.985 161.155 ;
        RECT 71.290 161.110 71.430 161.310 ;
        RECT 62.920 160.970 71.430 161.110 ;
        RECT 60.160 160.910 60.480 160.970 ;
        RECT 62.920 160.910 63.240 160.970 ;
        RECT 65.695 160.925 65.985 160.970 ;
        RECT 50.960 160.630 59.930 160.770 ;
        RECT 60.635 160.770 60.925 160.815 ;
        RECT 69.820 160.770 70.140 160.830 ;
        RECT 70.295 160.770 70.585 160.815 ;
        RECT 72.580 160.770 72.900 160.830 ;
        RECT 60.635 160.630 74.650 160.770 ;
        RECT 45.900 160.570 46.220 160.630 ;
        RECT 50.960 160.570 51.280 160.630 ;
        RECT 53.260 160.570 53.580 160.630 ;
        RECT 56.480 160.570 56.800 160.630 ;
        RECT 60.635 160.585 60.925 160.630 ;
        RECT 69.820 160.570 70.140 160.630 ;
        RECT 70.295 160.585 70.585 160.630 ;
        RECT 72.580 160.570 72.900 160.630 ;
        RECT 31.655 160.290 45.210 160.430 ;
        RECT 45.440 160.430 45.760 160.490 ;
        RECT 47.280 160.430 47.600 160.490 ;
        RECT 45.440 160.290 47.600 160.430 ;
        RECT 31.655 160.245 31.945 160.290 ;
        RECT 45.440 160.230 45.760 160.290 ;
        RECT 47.280 160.230 47.600 160.290 ;
        RECT 48.660 160.430 48.980 160.490 ;
        RECT 51.880 160.430 52.200 160.490 ;
        RECT 48.660 160.290 52.200 160.430 ;
        RECT 48.660 160.230 48.980 160.290 ;
        RECT 51.880 160.230 52.200 160.290 ;
        RECT 58.320 160.430 58.640 160.490 ;
        RECT 66.600 160.430 66.920 160.490 ;
        RECT 69.360 160.430 69.680 160.490 ;
        RECT 58.320 160.290 69.680 160.430 ;
        RECT 58.320 160.230 58.640 160.290 ;
        RECT 66.600 160.230 66.920 160.290 ;
        RECT 69.360 160.230 69.680 160.290 ;
        RECT 70.740 160.430 71.060 160.490 ;
        RECT 74.510 160.475 74.650 160.630 ;
        RECT 72.135 160.430 72.425 160.475 ;
        RECT 70.740 160.290 72.425 160.430 ;
        RECT 70.740 160.230 71.060 160.290 ;
        RECT 72.135 160.245 72.425 160.290 ;
        RECT 74.435 160.245 74.725 160.475 ;
        RECT 15.930 159.610 87.230 160.090 ;
        RECT 19.220 159.210 19.540 159.470 ;
        RECT 21.520 159.410 21.840 159.470 ;
        RECT 23.835 159.410 24.125 159.455 ;
        RECT 21.520 159.270 24.125 159.410 ;
        RECT 21.520 159.210 21.840 159.270 ;
        RECT 23.835 159.225 24.125 159.270 ;
        RECT 24.280 159.210 24.600 159.470 ;
        RECT 27.040 159.410 27.360 159.470 ;
        RECT 29.800 159.410 30.120 159.470 ;
        RECT 27.040 159.270 30.120 159.410 ;
        RECT 27.040 159.210 27.360 159.270 ;
        RECT 29.800 159.210 30.120 159.270 ;
        RECT 37.620 159.210 37.940 159.470 ;
        RECT 43.600 159.410 43.920 159.470 ;
        RECT 47.295 159.410 47.585 159.455 ;
        RECT 43.600 159.270 53.030 159.410 ;
        RECT 43.600 159.210 43.920 159.270 ;
        RECT 47.295 159.225 47.585 159.270 ;
        RECT 20.140 159.070 20.460 159.130 ;
        RECT 21.995 159.070 22.285 159.115 ;
        RECT 25.200 159.070 25.520 159.130 ;
        RECT 18.390 158.930 25.520 159.070 ;
        RECT 18.390 158.435 18.530 158.930 ;
        RECT 20.140 158.870 20.460 158.930 ;
        RECT 21.995 158.885 22.285 158.930 ;
        RECT 25.200 158.870 25.520 158.930 ;
        RECT 34.400 159.070 34.720 159.130 ;
        RECT 36.240 159.070 36.560 159.130 ;
        RECT 45.900 159.070 46.220 159.130 ;
        RECT 34.400 158.930 36.010 159.070 ;
        RECT 34.400 158.870 34.720 158.930 ;
        RECT 19.695 158.545 19.985 158.775 ;
        RECT 22.440 158.730 22.760 158.790 ;
        RECT 35.870 158.775 36.010 158.930 ;
        RECT 36.240 158.930 46.220 159.070 ;
        RECT 36.240 158.870 36.560 158.930 ;
        RECT 45.900 158.870 46.220 158.930 ;
        RECT 51.420 158.870 51.740 159.130 ;
        RECT 52.355 159.070 52.645 159.115 ;
        RECT 51.970 158.930 52.645 159.070 ;
        RECT 52.890 159.070 53.030 159.270 ;
        RECT 63.380 159.210 63.700 159.470 ;
        RECT 64.760 159.410 65.080 159.470 ;
        RECT 65.235 159.410 65.525 159.455 ;
        RECT 64.760 159.270 65.525 159.410 ;
        RECT 64.760 159.210 65.080 159.270 ;
        RECT 65.235 159.225 65.525 159.270 ;
        RECT 69.820 159.210 70.140 159.470 ;
        RECT 70.755 159.410 71.045 159.455 ;
        RECT 71.660 159.410 71.980 159.470 ;
        RECT 70.755 159.270 71.980 159.410 ;
        RECT 70.755 159.225 71.045 159.270 ;
        RECT 71.660 159.210 71.980 159.270 ;
        RECT 72.135 159.410 72.425 159.455 ;
        RECT 76.720 159.410 77.040 159.470 ;
        RECT 72.135 159.270 77.040 159.410 ;
        RECT 72.135 159.225 72.425 159.270 ;
        RECT 76.720 159.210 77.040 159.270 ;
        RECT 78.100 159.210 78.420 159.470 ;
        RECT 62.015 159.070 62.305 159.115 ;
        RECT 68.440 159.070 68.760 159.130 ;
        RECT 52.890 158.930 57.630 159.070 ;
        RECT 23.375 158.730 23.665 158.775 ;
        RECT 35.795 158.730 36.085 158.775 ;
        RECT 37.620 158.730 37.940 158.790 ;
        RECT 51.970 158.730 52.110 158.930 ;
        RECT 52.355 158.885 52.645 158.930 ;
        RECT 53.260 158.730 53.580 158.790 ;
        RECT 56.955 158.730 57.245 158.775 ;
        RECT 22.440 158.590 23.665 158.730 ;
        RECT 18.315 158.205 18.605 158.435 ;
        RECT 18.775 158.205 19.065 158.435 ;
        RECT 19.770 158.390 19.910 158.545 ;
        RECT 22.440 158.530 22.760 158.590 ;
        RECT 23.375 158.545 23.665 158.590 ;
        RECT 24.370 158.590 35.550 158.730 ;
        RECT 24.370 158.390 24.510 158.590 ;
        RECT 19.770 158.250 24.510 158.390 ;
        RECT 24.755 158.390 25.045 158.435 ;
        RECT 25.200 158.390 25.520 158.450 ;
        RECT 24.755 158.250 25.520 158.390 ;
        RECT 24.755 158.205 25.045 158.250 ;
        RECT 18.850 158.050 18.990 158.205 ;
        RECT 25.200 158.190 25.520 158.250 ;
        RECT 30.735 158.390 31.025 158.435 ;
        RECT 34.400 158.390 34.720 158.450 ;
        RECT 30.735 158.250 34.720 158.390 ;
        RECT 35.410 158.390 35.550 158.590 ;
        RECT 35.795 158.590 37.940 158.730 ;
        RECT 35.795 158.545 36.085 158.590 ;
        RECT 37.620 158.530 37.940 158.590 ;
        RECT 46.910 158.590 51.190 158.730 ;
        RECT 51.970 158.590 53.580 158.730 ;
        RECT 46.910 158.450 47.050 158.590 ;
        RECT 36.715 158.390 37.005 158.435 ;
        RECT 40.840 158.390 41.160 158.450 ;
        RECT 35.410 158.250 41.160 158.390 ;
        RECT 30.735 158.205 31.025 158.250 ;
        RECT 34.400 158.190 34.720 158.250 ;
        RECT 36.715 158.205 37.005 158.250 ;
        RECT 40.840 158.190 41.160 158.250 ;
        RECT 46.375 158.390 46.665 158.435 ;
        RECT 46.820 158.390 47.140 158.450 ;
        RECT 46.375 158.250 47.140 158.390 ;
        RECT 46.375 158.205 46.665 158.250 ;
        RECT 46.820 158.190 47.140 158.250 ;
        RECT 47.755 158.390 48.045 158.435 ;
        RECT 48.660 158.390 48.980 158.450 ;
        RECT 47.755 158.250 48.980 158.390 ;
        RECT 47.755 158.205 48.045 158.250 ;
        RECT 48.660 158.190 48.980 158.250 ;
        RECT 50.040 158.190 50.360 158.450 ;
        RECT 51.050 158.390 51.190 158.590 ;
        RECT 53.260 158.530 53.580 158.590 ;
        RECT 55.190 158.590 57.245 158.730 ;
        RECT 55.190 158.390 55.330 158.590 ;
        RECT 56.955 158.545 57.245 158.590 ;
        RECT 51.050 158.250 55.330 158.390 ;
        RECT 55.575 158.390 55.865 158.435 ;
        RECT 56.020 158.390 56.340 158.450 ;
        RECT 55.575 158.250 56.340 158.390 ;
        RECT 55.575 158.205 55.865 158.250 ;
        RECT 56.020 158.190 56.340 158.250 ;
        RECT 20.155 158.050 20.445 158.095 ;
        RECT 24.280 158.050 24.600 158.110 ;
        RECT 18.850 157.910 24.600 158.050 ;
        RECT 40.930 158.050 41.070 158.190 ;
        RECT 57.030 158.050 57.170 158.545 ;
        RECT 57.490 158.390 57.630 158.930 ;
        RECT 62.015 158.930 68.760 159.070 ;
        RECT 62.015 158.885 62.305 158.930 ;
        RECT 68.440 158.870 68.760 158.930 ;
        RECT 68.990 158.930 78.790 159.070 ;
        RECT 61.540 158.730 61.860 158.790 ;
        RECT 63.395 158.730 63.685 158.775 ;
        RECT 61.540 158.590 63.685 158.730 ;
        RECT 61.540 158.530 61.860 158.590 ;
        RECT 63.395 158.545 63.685 158.590 ;
        RECT 63.840 158.730 64.160 158.790 ;
        RECT 68.990 158.730 69.130 158.930 ;
        RECT 78.650 158.775 78.790 158.930 ;
        RECT 63.840 158.590 69.130 158.730 ;
        RECT 78.575 158.730 78.865 158.775 ;
        RECT 78.575 158.590 84.770 158.730 ;
        RECT 63.840 158.530 64.160 158.590 ;
        RECT 78.575 158.545 78.865 158.590 ;
        RECT 84.630 158.450 84.770 158.590 ;
        RECT 57.875 158.390 58.165 158.435 ;
        RECT 59.700 158.390 60.020 158.450 ;
        RECT 57.490 158.250 60.020 158.390 ;
        RECT 57.875 158.205 58.165 158.250 ;
        RECT 59.700 158.190 60.020 158.250 ;
        RECT 60.160 158.390 60.480 158.450 ;
        RECT 60.635 158.390 60.925 158.435 ;
        RECT 60.160 158.250 60.925 158.390 ;
        RECT 60.160 158.190 60.480 158.250 ;
        RECT 60.635 158.205 60.925 158.250 ;
        RECT 61.080 158.190 61.400 158.450 ;
        RECT 62.920 158.190 63.240 158.450 ;
        RECT 64.315 158.205 64.605 158.435 ;
        RECT 67.980 158.390 68.300 158.450 ;
        RECT 71.200 158.390 71.520 158.450 ;
        RECT 67.980 158.250 71.520 158.390 ;
        RECT 62.015 158.050 62.305 158.095 ;
        RECT 62.460 158.050 62.780 158.110 ;
        RECT 64.390 158.050 64.530 158.205 ;
        RECT 67.980 158.190 68.300 158.250 ;
        RECT 71.200 158.190 71.520 158.250 ;
        RECT 72.135 158.390 72.425 158.435 ;
        RECT 74.420 158.390 74.740 158.450 ;
        RECT 72.135 158.250 74.740 158.390 ;
        RECT 72.135 158.205 72.425 158.250 ;
        RECT 68.915 158.050 69.205 158.095 ;
        RECT 72.210 158.050 72.350 158.205 ;
        RECT 74.420 158.190 74.740 158.250 ;
        RECT 77.195 158.390 77.485 158.435 ;
        RECT 79.020 158.390 79.340 158.450 ;
        RECT 77.195 158.250 79.340 158.390 ;
        RECT 77.195 158.205 77.485 158.250 ;
        RECT 79.020 158.190 79.340 158.250 ;
        RECT 81.335 158.205 81.625 158.435 ;
        RECT 40.930 157.910 52.110 158.050 ;
        RECT 57.030 157.910 62.780 158.050 ;
        RECT 20.155 157.865 20.445 157.910 ;
        RECT 24.280 157.850 24.600 157.910 ;
        RECT 22.455 157.710 22.745 157.755 ;
        RECT 28.880 157.710 29.200 157.770 ;
        RECT 22.455 157.570 29.200 157.710 ;
        RECT 22.455 157.525 22.745 157.570 ;
        RECT 28.880 157.510 29.200 157.570 ;
        RECT 45.440 157.510 45.760 157.770 ;
        RECT 51.970 157.710 52.110 157.910 ;
        RECT 62.015 157.865 62.305 157.910 ;
        RECT 62.460 157.850 62.780 157.910 ;
        RECT 63.010 157.910 69.205 158.050 ;
        RECT 63.010 157.770 63.150 157.910 ;
        RECT 68.915 157.865 69.205 157.910 ;
        RECT 70.370 157.910 72.350 158.050 ;
        RECT 79.495 158.050 79.785 158.095 ;
        RECT 79.940 158.050 80.260 158.110 ;
        RECT 79.495 157.910 80.260 158.050 ;
        RECT 56.035 157.710 56.325 157.755 ;
        RECT 51.970 157.570 56.325 157.710 ;
        RECT 56.035 157.525 56.325 157.570 ;
        RECT 56.480 157.510 56.800 157.770 ;
        RECT 56.940 157.510 57.260 157.770 ;
        RECT 62.920 157.510 63.240 157.770 ;
        RECT 68.440 157.710 68.760 157.770 ;
        RECT 69.915 157.710 70.205 157.755 ;
        RECT 70.370 157.710 70.510 157.910 ;
        RECT 79.495 157.865 79.785 157.910 ;
        RECT 79.940 157.850 80.260 157.910 ;
        RECT 68.440 157.570 70.510 157.710 ;
        RECT 79.020 157.710 79.340 157.770 ;
        RECT 81.410 157.710 81.550 158.205 ;
        RECT 84.080 158.190 84.400 158.450 ;
        RECT 84.540 158.390 84.860 158.450 ;
        RECT 85.015 158.390 85.305 158.435 ;
        RECT 84.540 158.250 85.305 158.390 ;
        RECT 84.540 158.190 84.860 158.250 ;
        RECT 85.015 158.205 85.305 158.250 ;
        RECT 79.020 157.570 81.550 157.710 ;
        RECT 82.255 157.710 82.545 157.755 ;
        RECT 82.700 157.710 83.020 157.770 ;
        RECT 82.255 157.570 83.020 157.710 ;
        RECT 68.440 157.510 68.760 157.570 ;
        RECT 69.915 157.525 70.205 157.570 ;
        RECT 79.020 157.510 79.340 157.570 ;
        RECT 82.255 157.525 82.545 157.570 ;
        RECT 82.700 157.510 83.020 157.570 ;
        RECT 84.555 157.710 84.845 157.755 ;
        RECT 85.460 157.710 85.780 157.770 ;
        RECT 84.555 157.570 85.780 157.710 ;
        RECT 84.555 157.525 84.845 157.570 ;
        RECT 85.460 157.510 85.780 157.570 ;
        RECT 15.930 156.890 87.230 157.370 ;
        RECT 23.360 156.690 23.680 156.750 ;
        RECT 24.295 156.690 24.585 156.735 ;
        RECT 23.360 156.550 24.585 156.690 ;
        RECT 23.360 156.490 23.680 156.550 ;
        RECT 24.295 156.505 24.585 156.550 ;
        RECT 26.135 156.690 26.425 156.735 ;
        RECT 40.380 156.690 40.700 156.750 ;
        RECT 26.135 156.550 40.700 156.690 ;
        RECT 26.135 156.505 26.425 156.550 ;
        RECT 40.380 156.490 40.700 156.550 ;
        RECT 42.220 156.490 42.540 156.750 ;
        RECT 57.860 156.690 58.180 156.750 ;
        RECT 44.150 156.550 58.180 156.690 ;
        RECT 27.040 156.150 27.360 156.410 ;
        RECT 27.500 156.350 27.820 156.410 ;
        RECT 37.175 156.350 37.465 156.395 ;
        RECT 44.150 156.350 44.290 156.550 ;
        RECT 57.860 156.490 58.180 156.550 ;
        RECT 68.900 156.690 69.220 156.750 ;
        RECT 68.900 156.550 70.050 156.690 ;
        RECT 68.900 156.490 69.220 156.550 ;
        RECT 45.440 156.350 45.760 156.410 ;
        RECT 27.500 156.210 36.470 156.350 ;
        RECT 27.500 156.150 27.820 156.210 ;
        RECT 27.590 155.870 30.030 156.010 ;
        RECT 17.380 155.470 17.700 155.730 ;
        RECT 18.775 155.670 19.065 155.715 ;
        RECT 22.915 155.670 23.205 155.715 ;
        RECT 18.775 155.530 23.205 155.670 ;
        RECT 18.775 155.485 19.065 155.530 ;
        RECT 22.915 155.485 23.205 155.530 ;
        RECT 22.990 155.330 23.130 155.485 ;
        RECT 24.740 155.470 25.060 155.730 ;
        RECT 25.200 155.715 25.520 155.730 ;
        RECT 25.200 155.670 25.630 155.715 ;
        RECT 27.590 155.670 27.730 155.870 ;
        RECT 29.890 155.730 30.030 155.870 ;
        RECT 33.940 155.810 34.260 156.070 ;
        RECT 34.860 155.810 35.180 156.070 ;
        RECT 36.330 156.055 36.470 156.210 ;
        RECT 37.175 156.210 44.290 156.350 ;
        RECT 44.610 156.210 45.760 156.350 ;
        RECT 37.175 156.165 37.465 156.210 ;
        RECT 36.255 156.010 36.545 156.055 ;
        RECT 37.620 156.010 37.940 156.070 ;
        RECT 36.255 155.870 37.940 156.010 ;
        RECT 36.255 155.825 36.545 155.870 ;
        RECT 37.620 155.810 37.940 155.870 ;
        RECT 43.155 155.825 43.445 156.055 ;
        RECT 43.615 156.010 43.905 156.055 ;
        RECT 44.060 156.010 44.380 156.070 ;
        RECT 44.610 156.055 44.750 156.210 ;
        RECT 45.440 156.150 45.760 156.210 ;
        RECT 45.900 156.350 46.220 156.410 ;
        RECT 50.500 156.350 50.820 156.410 ;
        RECT 62.475 156.350 62.765 156.395 ;
        RECT 45.900 156.210 50.270 156.350 ;
        RECT 45.900 156.150 46.220 156.210 ;
        RECT 43.615 155.870 44.380 156.010 ;
        RECT 43.615 155.825 43.905 155.870 ;
        RECT 25.200 155.530 27.730 155.670 ;
        RECT 25.200 155.485 25.630 155.530 ;
        RECT 25.200 155.470 25.520 155.485 ;
        RECT 29.340 155.470 29.660 155.730 ;
        RECT 29.800 155.470 30.120 155.730 ;
        RECT 43.230 155.670 43.370 155.825 ;
        RECT 44.060 155.810 44.380 155.870 ;
        RECT 44.535 155.825 44.825 156.055 ;
        RECT 44.980 155.810 45.300 156.070 ;
        RECT 46.375 156.010 46.665 156.055 ;
        RECT 46.820 156.010 47.140 156.070 ;
        RECT 46.375 155.870 47.140 156.010 ;
        RECT 46.375 155.825 46.665 155.870 ;
        RECT 45.455 155.670 45.745 155.715 ;
        RECT 43.230 155.530 45.745 155.670 ;
        RECT 45.455 155.485 45.745 155.530 ;
        RECT 24.280 155.330 24.600 155.390 ;
        RECT 27.040 155.330 27.360 155.390 ;
        RECT 22.990 155.190 27.360 155.330 ;
        RECT 29.430 155.330 29.570 155.470 ;
        RECT 30.735 155.330 31.025 155.375 ;
        RECT 46.450 155.330 46.590 155.825 ;
        RECT 46.820 155.810 47.140 155.870 ;
        RECT 47.280 155.810 47.600 156.070 ;
        RECT 47.740 155.810 48.060 156.070 ;
        RECT 50.130 156.055 50.270 156.210 ;
        RECT 50.500 156.210 62.765 156.350 ;
        RECT 50.500 156.150 50.820 156.210 ;
        RECT 62.475 156.165 62.765 156.210 ;
        RECT 50.055 155.825 50.345 156.055 ;
        RECT 50.975 156.010 51.265 156.055 ;
        RECT 51.880 156.010 52.200 156.070 ;
        RECT 50.975 155.870 52.200 156.010 ;
        RECT 50.975 155.825 51.265 155.870 ;
        RECT 50.130 155.670 50.270 155.825 ;
        RECT 51.880 155.810 52.200 155.870 ;
        RECT 62.935 155.825 63.225 156.055 ;
        RECT 67.520 156.010 67.840 156.070 ;
        RECT 67.995 156.010 68.285 156.055 ;
        RECT 67.520 155.870 68.285 156.010 ;
        RECT 51.420 155.670 51.740 155.730 ;
        RECT 50.130 155.530 51.740 155.670 ;
        RECT 63.010 155.670 63.150 155.825 ;
        RECT 67.520 155.810 67.840 155.870 ;
        RECT 67.995 155.825 68.285 155.870 ;
        RECT 68.455 156.010 68.745 156.055 ;
        RECT 68.900 156.010 69.220 156.070 ;
        RECT 68.455 155.870 69.220 156.010 ;
        RECT 68.455 155.825 68.745 155.870 ;
        RECT 68.530 155.670 68.670 155.825 ;
        RECT 68.900 155.810 69.220 155.870 ;
        RECT 69.375 155.825 69.665 156.055 ;
        RECT 69.910 156.010 70.050 156.550 ;
        RECT 70.280 156.490 70.600 156.750 ;
        RECT 81.795 156.690 82.085 156.735 ;
        RECT 82.240 156.690 82.560 156.750 ;
        RECT 81.795 156.550 82.560 156.690 ;
        RECT 81.795 156.505 82.085 156.550 ;
        RECT 82.240 156.490 82.560 156.550 ;
        RECT 82.715 156.505 83.005 156.735 ;
        RECT 79.020 156.350 79.340 156.410 ;
        RECT 82.790 156.350 82.930 156.505 ;
        RECT 85.000 156.490 85.320 156.750 ;
        RECT 84.540 156.350 84.860 156.410 ;
        RECT 86.840 156.350 87.160 156.410 ;
        RECT 72.210 156.210 82.930 156.350 ;
        RECT 83.710 156.210 87.160 156.350 ;
        RECT 71.675 156.010 71.965 156.055 ;
        RECT 69.910 155.870 71.965 156.010 ;
        RECT 71.675 155.825 71.965 155.870 ;
        RECT 69.450 155.670 69.590 155.825 ;
        RECT 69.820 155.670 70.140 155.730 ;
        RECT 63.010 155.530 68.670 155.670 ;
        RECT 68.990 155.530 70.140 155.670 ;
        RECT 51.420 155.470 51.740 155.530 ;
        RECT 52.800 155.330 53.120 155.390 ;
        RECT 29.430 155.190 30.030 155.330 ;
        RECT 24.280 155.130 24.600 155.190 ;
        RECT 27.040 155.130 27.360 155.190 ;
        RECT 29.890 154.990 30.030 155.190 ;
        RECT 30.735 155.190 46.590 155.330 ;
        RECT 46.910 155.190 53.120 155.330 ;
        RECT 30.735 155.145 31.025 155.190 ;
        RECT 41.760 154.990 42.080 155.050 ;
        RECT 46.910 154.990 47.050 155.190 ;
        RECT 52.800 155.130 53.120 155.190 ;
        RECT 53.260 155.330 53.580 155.390 ;
        RECT 57.860 155.330 58.180 155.390 ;
        RECT 66.140 155.330 66.460 155.390 ;
        RECT 68.990 155.330 69.130 155.530 ;
        RECT 69.820 155.470 70.140 155.530 ;
        RECT 53.260 155.190 69.130 155.330 ;
        RECT 69.360 155.330 69.680 155.390 ;
        RECT 70.755 155.330 71.045 155.375 ;
        RECT 69.360 155.190 71.045 155.330 ;
        RECT 53.260 155.130 53.580 155.190 ;
        RECT 57.860 155.130 58.180 155.190 ;
        RECT 66.140 155.130 66.460 155.190 ;
        RECT 69.360 155.130 69.680 155.190 ;
        RECT 70.755 155.145 71.045 155.190 ;
        RECT 29.890 154.850 47.050 154.990 ;
        RECT 41.760 154.790 42.080 154.850 ;
        RECT 50.960 154.790 51.280 155.050 ;
        RECT 51.420 154.990 51.740 155.050 ;
        RECT 53.350 154.990 53.490 155.130 ;
        RECT 51.420 154.850 53.490 154.990 ;
        RECT 58.780 154.990 59.100 155.050 ;
        RECT 72.210 154.990 72.350 156.210 ;
        RECT 79.020 156.150 79.340 156.210 ;
        RECT 80.400 155.810 80.720 156.070 ;
        RECT 80.875 156.010 81.165 156.055 ;
        RECT 81.780 156.010 82.100 156.070 ;
        RECT 83.710 156.055 83.850 156.210 ;
        RECT 84.540 156.150 84.860 156.210 ;
        RECT 86.840 156.150 87.160 156.210 ;
        RECT 80.875 155.870 82.100 156.010 ;
        RECT 80.875 155.825 81.165 155.870 ;
        RECT 81.780 155.810 82.100 155.870 ;
        RECT 83.635 155.825 83.925 156.055 ;
        RECT 84.095 155.825 84.385 156.055 ;
        RECT 72.595 155.485 72.885 155.715 ;
        RECT 81.320 155.670 81.640 155.730 ;
        RECT 84.170 155.670 84.310 155.825 ;
        RECT 81.320 155.530 84.310 155.670 ;
        RECT 72.670 155.330 72.810 155.485 ;
        RECT 81.320 155.470 81.640 155.530 ;
        RECT 85.460 155.330 85.780 155.390 ;
        RECT 72.670 155.190 85.780 155.330 ;
        RECT 85.460 155.130 85.780 155.190 ;
        RECT 58.780 154.850 72.350 154.990 ;
        RECT 51.420 154.790 51.740 154.850 ;
        RECT 58.780 154.790 59.100 154.850 ;
        RECT 79.480 154.790 79.800 155.050 ;
        RECT 15.930 154.170 87.230 154.650 ;
        RECT 22.455 153.970 22.745 154.015 ;
        RECT 22.900 153.970 23.220 154.030 ;
        RECT 22.455 153.830 23.220 153.970 ;
        RECT 22.455 153.785 22.745 153.830 ;
        RECT 22.900 153.770 23.220 153.830 ;
        RECT 23.360 153.970 23.680 154.030 ;
        RECT 27.055 153.970 27.345 154.015 ;
        RECT 30.260 153.970 30.580 154.030 ;
        RECT 31.195 153.970 31.485 154.015 ;
        RECT 23.360 153.830 27.345 153.970 ;
        RECT 23.360 153.770 23.680 153.830 ;
        RECT 27.055 153.785 27.345 153.830 ;
        RECT 27.590 153.830 31.485 153.970 ;
        RECT 21.995 153.630 22.285 153.675 ;
        RECT 24.280 153.630 24.600 153.690 ;
        RECT 21.995 153.490 24.600 153.630 ;
        RECT 21.995 153.445 22.285 153.490 ;
        RECT 22.070 153.290 22.210 153.445 ;
        RECT 24.280 153.430 24.600 153.490 ;
        RECT 24.740 153.630 25.060 153.690 ;
        RECT 25.215 153.630 25.505 153.675 ;
        RECT 27.590 153.630 27.730 153.830 ;
        RECT 30.260 153.770 30.580 153.830 ;
        RECT 31.195 153.785 31.485 153.830 ;
        RECT 34.860 153.970 35.180 154.030 ;
        RECT 43.155 153.970 43.445 154.015 ;
        RECT 44.980 153.970 45.300 154.030 ;
        RECT 34.860 153.830 42.450 153.970 ;
        RECT 34.860 153.770 35.180 153.830 ;
        RECT 24.740 153.490 27.730 153.630 ;
        RECT 32.115 153.630 32.405 153.675 ;
        RECT 33.940 153.630 34.260 153.690 ;
        RECT 32.115 153.490 35.090 153.630 ;
        RECT 24.740 153.430 25.060 153.490 ;
        RECT 25.215 153.445 25.505 153.490 ;
        RECT 32.115 153.445 32.405 153.490 ;
        RECT 33.940 153.430 34.260 153.490 ;
        RECT 18.850 153.150 22.210 153.290 ;
        RECT 29.430 153.150 34.630 153.290 ;
        RECT 18.850 152.995 18.990 153.150 ;
        RECT 18.775 152.765 19.065 152.995 ;
        RECT 19.695 152.765 19.985 152.995 ;
        RECT 23.360 152.950 23.680 153.010 ;
        RECT 29.430 152.995 29.570 153.150 ;
        RECT 29.355 152.950 29.645 152.995 ;
        RECT 23.360 152.810 29.645 152.950 ;
        RECT 19.220 152.610 19.540 152.670 ;
        RECT 19.770 152.610 19.910 152.765 ;
        RECT 23.360 152.750 23.680 152.810 ;
        RECT 29.355 152.765 29.645 152.810 ;
        RECT 33.480 152.750 33.800 153.010 ;
        RECT 33.940 152.950 34.260 153.010 ;
        RECT 34.490 152.995 34.630 153.150 ;
        RECT 34.415 152.950 34.705 152.995 ;
        RECT 33.940 152.810 34.705 152.950 ;
        RECT 34.950 152.950 35.090 153.490 ;
        RECT 35.335 153.290 35.625 153.335 ;
        RECT 35.335 153.150 40.610 153.290 ;
        RECT 35.335 153.105 35.625 153.150 ;
        RECT 40.470 153.010 40.610 153.150 ;
        RECT 35.795 152.950 36.085 152.995 ;
        RECT 39.475 152.950 39.765 152.995 ;
        RECT 34.950 152.810 39.765 152.950 ;
        RECT 33.940 152.750 34.260 152.810 ;
        RECT 34.415 152.765 34.705 152.810 ;
        RECT 35.795 152.765 36.085 152.810 ;
        RECT 39.475 152.765 39.765 152.810 ;
        RECT 20.155 152.610 20.445 152.655 ;
        RECT 25.200 152.610 25.520 152.670 ;
        RECT 19.220 152.470 25.520 152.610 ;
        RECT 19.220 152.410 19.540 152.470 ;
        RECT 20.155 152.425 20.445 152.470 ;
        RECT 25.200 152.410 25.520 152.470 ;
        RECT 27.040 152.410 27.360 152.670 ;
        RECT 29.800 152.610 30.120 152.670 ;
        RECT 31.195 152.610 31.485 152.655 ;
        RECT 29.800 152.470 31.485 152.610 ;
        RECT 34.490 152.610 34.630 152.765 ;
        RECT 40.380 152.750 40.700 153.010 ;
        RECT 41.760 152.750 42.080 153.010 ;
        RECT 42.310 152.995 42.450 153.830 ;
        RECT 43.155 153.830 45.300 153.970 ;
        RECT 43.155 153.785 43.445 153.830 ;
        RECT 44.980 153.770 45.300 153.830 ;
        RECT 46.360 153.970 46.680 154.030 ;
        RECT 48.215 153.970 48.505 154.015 ;
        RECT 46.360 153.830 48.505 153.970 ;
        RECT 46.360 153.770 46.680 153.830 ;
        RECT 48.215 153.785 48.505 153.830 ;
        RECT 52.815 153.970 53.105 154.015 ;
        RECT 53.260 153.970 53.580 154.030 ;
        RECT 52.815 153.830 53.580 153.970 ;
        RECT 52.815 153.785 53.105 153.830 ;
        RECT 53.260 153.770 53.580 153.830 ;
        RECT 55.100 153.770 55.420 154.030 ;
        RECT 56.480 153.970 56.800 154.030 ;
        RECT 57.415 153.970 57.705 154.015 ;
        RECT 56.480 153.830 57.705 153.970 ;
        RECT 56.480 153.770 56.800 153.830 ;
        RECT 57.415 153.785 57.705 153.830 ;
        RECT 61.095 153.970 61.385 154.015 ;
        RECT 63.840 153.970 64.160 154.030 ;
        RECT 61.095 153.830 64.160 153.970 ;
        RECT 61.095 153.785 61.385 153.830 ;
        RECT 63.840 153.770 64.160 153.830 ;
        RECT 67.980 153.770 68.300 154.030 ;
        RECT 83.620 153.770 83.940 154.030 ;
        RECT 45.455 153.630 45.745 153.675 ;
        RECT 49.120 153.630 49.440 153.690 ;
        RECT 52.340 153.630 52.660 153.690 ;
        RECT 45.455 153.490 52.660 153.630 ;
        RECT 45.455 153.445 45.745 153.490 ;
        RECT 49.120 153.430 49.440 153.490 ;
        RECT 52.340 153.430 52.660 153.490 ;
        RECT 53.720 153.630 54.040 153.690 ;
        RECT 53.720 153.490 59.470 153.630 ;
        RECT 53.720 153.430 54.040 153.490 ;
        RECT 50.040 153.290 50.360 153.350 ;
        RECT 43.690 153.150 50.360 153.290 ;
        RECT 42.235 152.765 42.525 152.995 ;
        RECT 43.140 152.950 43.460 153.010 ;
        RECT 43.690 152.995 43.830 153.150 ;
        RECT 50.040 153.090 50.360 153.150 ;
        RECT 51.510 153.150 58.550 153.290 ;
        RECT 44.520 152.995 44.840 153.010 ;
        RECT 43.615 152.950 43.905 152.995 ;
        RECT 43.140 152.810 43.905 152.950 ;
        RECT 43.140 152.750 43.460 152.810 ;
        RECT 43.615 152.765 43.905 152.810 ;
        RECT 44.385 152.765 44.840 152.995 ;
        RECT 49.135 152.950 49.425 152.995 ;
        RECT 49.135 152.810 50.730 152.950 ;
        RECT 49.135 152.765 49.425 152.810 ;
        RECT 44.520 152.750 44.840 152.765 ;
        RECT 34.490 152.470 38.310 152.610 ;
        RECT 29.800 152.410 30.120 152.470 ;
        RECT 31.195 152.425 31.485 152.470 ;
        RECT 17.855 152.270 18.145 152.315 ;
        RECT 27.500 152.270 27.820 152.330 ;
        RECT 17.855 152.130 27.820 152.270 ;
        RECT 17.855 152.085 18.145 152.130 ;
        RECT 27.500 152.070 27.820 152.130 ;
        RECT 27.975 152.270 28.265 152.315 ;
        RECT 33.020 152.270 33.340 152.330 ;
        RECT 34.860 152.270 35.180 152.330 ;
        RECT 27.975 152.130 35.180 152.270 ;
        RECT 27.975 152.085 28.265 152.130 ;
        RECT 33.020 152.070 33.340 152.130 ;
        RECT 34.860 152.070 35.180 152.130 ;
        RECT 37.175 152.270 37.465 152.315 ;
        RECT 37.620 152.270 37.940 152.330 ;
        RECT 38.170 152.315 38.310 152.470 ;
        RECT 38.540 152.410 38.860 152.670 ;
        RECT 44.610 152.610 44.750 152.750 ;
        RECT 49.580 152.610 49.900 152.670 ;
        RECT 44.610 152.470 49.900 152.610 ;
        RECT 49.580 152.410 49.900 152.470 ;
        RECT 50.040 152.410 50.360 152.670 ;
        RECT 50.590 152.610 50.730 152.810 ;
        RECT 50.960 152.750 51.280 153.010 ;
        RECT 51.510 152.995 51.650 153.150 ;
        RECT 51.435 152.765 51.725 152.995 ;
        RECT 51.895 152.960 52.185 152.995 ;
        RECT 51.895 152.950 52.570 152.960 ;
        RECT 52.800 152.950 53.120 153.010 ;
        RECT 51.895 152.820 53.120 152.950 ;
        RECT 51.895 152.765 52.185 152.820 ;
        RECT 52.430 152.810 53.120 152.820 ;
        RECT 52.800 152.750 53.120 152.810 ;
        RECT 56.020 152.750 56.340 153.010 ;
        RECT 56.495 152.950 56.785 152.995 ;
        RECT 56.940 152.950 57.260 153.010 ;
        RECT 56.495 152.810 57.260 152.950 ;
        RECT 56.495 152.765 56.785 152.810 ;
        RECT 55.100 152.610 55.420 152.670 ;
        RECT 56.570 152.610 56.710 152.765 ;
        RECT 56.940 152.750 57.260 152.810 ;
        RECT 57.860 152.750 58.180 153.010 ;
        RECT 50.590 152.470 51.880 152.610 ;
        RECT 37.175 152.130 37.940 152.270 ;
        RECT 37.175 152.085 37.465 152.130 ;
        RECT 37.620 152.070 37.940 152.130 ;
        RECT 38.095 152.085 38.385 152.315 ;
        RECT 39.920 152.070 40.240 152.330 ;
        RECT 51.740 152.270 51.880 152.470 ;
        RECT 55.100 152.470 56.710 152.610 ;
        RECT 58.410 152.610 58.550 153.150 ;
        RECT 58.780 152.750 59.100 153.010 ;
        RECT 59.330 152.995 59.470 153.490 ;
        RECT 62.015 153.445 62.305 153.675 ;
        RECT 63.380 153.630 63.700 153.690 ;
        RECT 69.835 153.630 70.125 153.675 ;
        RECT 73.500 153.630 73.820 153.690 ;
        RECT 63.380 153.490 73.820 153.630 ;
        RECT 62.090 153.290 62.230 153.445 ;
        RECT 63.380 153.430 63.700 153.490 ;
        RECT 69.835 153.445 70.125 153.490 ;
        RECT 73.500 153.430 73.820 153.490 ;
        RECT 85.460 153.430 85.780 153.690 ;
        RECT 62.090 153.150 69.130 153.290 ;
        RECT 59.255 152.765 59.545 152.995 ;
        RECT 61.080 152.750 61.400 153.010 ;
        RECT 63.010 152.995 63.150 153.150 ;
        RECT 68.990 153.010 69.130 153.150 ;
        RECT 62.935 152.765 63.225 152.995 ;
        RECT 63.905 152.950 64.195 152.995 ;
        RECT 63.905 152.810 64.530 152.950 ;
        RECT 63.905 152.765 64.195 152.810 ;
        RECT 62.460 152.610 62.780 152.670 ;
        RECT 58.410 152.470 62.780 152.610 ;
        RECT 64.390 152.610 64.530 152.810 ;
        RECT 65.680 152.750 66.000 153.010 ;
        RECT 67.060 152.750 67.380 153.010 ;
        RECT 67.520 152.950 67.840 153.010 ;
        RECT 68.455 152.950 68.745 152.995 ;
        RECT 67.520 152.810 68.745 152.950 ;
        RECT 67.520 152.750 67.840 152.810 ;
        RECT 68.455 152.765 68.745 152.810 ;
        RECT 68.900 152.750 69.220 153.010 ;
        RECT 69.820 152.750 70.140 153.010 ;
        RECT 82.700 152.750 83.020 153.010 ;
        RECT 64.760 152.610 65.080 152.670 ;
        RECT 67.610 152.610 67.750 152.750 ;
        RECT 64.390 152.470 67.750 152.610 ;
        RECT 79.480 152.610 79.800 152.670 ;
        RECT 84.555 152.610 84.845 152.655 ;
        RECT 79.480 152.470 84.845 152.610 ;
        RECT 55.100 152.410 55.420 152.470 ;
        RECT 62.460 152.410 62.780 152.470 ;
        RECT 64.760 152.410 65.080 152.470 ;
        RECT 79.480 152.410 79.800 152.470 ;
        RECT 84.555 152.425 84.845 152.470 ;
        RECT 53.720 152.270 54.040 152.330 ;
        RECT 62.935 152.270 63.225 152.315 ;
        RECT 51.740 152.130 63.225 152.270 ;
        RECT 53.720 152.070 54.040 152.130 ;
        RECT 62.935 152.085 63.225 152.130 ;
        RECT 66.140 152.070 66.460 152.330 ;
        RECT 15.930 151.450 87.230 151.930 ;
        RECT 33.940 151.050 34.260 151.310 ;
        RECT 35.795 151.250 36.085 151.295 ;
        RECT 47.740 151.250 48.060 151.310 ;
        RECT 63.380 151.250 63.700 151.310 ;
        RECT 34.490 151.110 48.060 151.250 ;
        RECT 33.020 150.710 33.340 150.970 ;
        RECT 33.480 150.910 33.800 150.970 ;
        RECT 34.490 150.910 34.630 151.110 ;
        RECT 35.795 151.065 36.085 151.110 ;
        RECT 47.740 151.050 48.060 151.110 ;
        RECT 51.510 151.110 63.700 151.250 ;
        RECT 33.480 150.770 34.630 150.910 ;
        RECT 33.480 150.710 33.800 150.770 ;
        RECT 18.775 150.385 19.065 150.615 ;
        RECT 18.850 150.230 18.990 150.385 ;
        RECT 19.220 150.370 19.540 150.630 ;
        RECT 34.490 150.615 34.630 150.770 ;
        RECT 49.580 150.710 49.900 150.970 ;
        RECT 19.695 150.570 19.985 150.615 ;
        RECT 21.535 150.570 21.825 150.615 ;
        RECT 19.695 150.430 21.825 150.570 ;
        RECT 19.695 150.385 19.985 150.430 ;
        RECT 21.535 150.385 21.825 150.430 ;
        RECT 34.415 150.385 34.705 150.615 ;
        RECT 34.875 150.385 35.165 150.615 ;
        RECT 49.135 150.385 49.425 150.615 ;
        RECT 22.900 150.230 23.220 150.290 ;
        RECT 34.950 150.230 35.090 150.385 ;
        RECT 18.850 150.090 20.830 150.230 ;
        RECT 17.840 149.690 18.160 149.950 ;
        RECT 20.690 149.935 20.830 150.090 ;
        RECT 22.900 150.090 35.090 150.230 ;
        RECT 22.900 150.030 23.220 150.090 ;
        RECT 20.615 149.705 20.905 149.935 ;
        RECT 48.200 149.690 48.520 149.950 ;
        RECT 33.035 149.550 33.325 149.595 ;
        RECT 33.480 149.550 33.800 149.610 ;
        RECT 33.035 149.410 33.800 149.550 ;
        RECT 49.210 149.550 49.350 150.385 ;
        RECT 50.040 150.370 50.360 150.630 ;
        RECT 51.510 150.615 51.650 151.110 ;
        RECT 63.380 151.050 63.700 151.110 ;
        RECT 63.930 151.110 67.290 151.250 ;
        RECT 54.640 150.910 54.960 150.970 ;
        RECT 55.575 150.910 55.865 150.955 ;
        RECT 57.860 150.910 58.180 150.970 ;
        RECT 63.930 150.910 64.070 151.110 ;
        RECT 67.150 150.970 67.290 151.110 ;
        RECT 66.140 150.910 66.460 150.970 ;
        RECT 51.970 150.770 54.410 150.910 ;
        RECT 51.970 150.630 52.110 150.770 ;
        RECT 50.975 150.385 51.265 150.615 ;
        RECT 51.435 150.385 51.725 150.615 ;
        RECT 51.050 150.230 51.190 150.385 ;
        RECT 51.880 150.370 52.200 150.630 ;
        RECT 52.800 150.370 53.120 150.630 ;
        RECT 53.720 150.370 54.040 150.630 ;
        RECT 54.270 150.615 54.410 150.770 ;
        RECT 54.640 150.770 55.865 150.910 ;
        RECT 54.640 150.710 54.960 150.770 ;
        RECT 55.575 150.725 55.865 150.770 ;
        RECT 57.030 150.770 58.180 150.910 ;
        RECT 54.195 150.385 54.485 150.615 ;
        RECT 55.100 150.370 55.420 150.630 ;
        RECT 56.020 150.570 56.340 150.630 ;
        RECT 57.030 150.615 57.170 150.770 ;
        RECT 57.860 150.710 58.180 150.770 ;
        RECT 58.410 150.770 64.070 150.910 ;
        RECT 65.310 150.770 66.460 150.910 ;
        RECT 56.495 150.570 56.785 150.615 ;
        RECT 56.020 150.430 56.785 150.570 ;
        RECT 56.020 150.370 56.340 150.430 ;
        RECT 56.495 150.385 56.785 150.430 ;
        RECT 56.955 150.385 57.245 150.615 ;
        RECT 57.400 150.570 57.720 150.630 ;
        RECT 58.410 150.615 58.550 150.770 ;
        RECT 58.335 150.570 58.625 150.615 ;
        RECT 57.400 150.430 58.625 150.570 ;
        RECT 54.655 150.230 54.945 150.275 ;
        RECT 51.050 150.090 54.945 150.230 ;
        RECT 56.570 150.230 56.710 150.385 ;
        RECT 57.400 150.370 57.720 150.430 ;
        RECT 58.335 150.385 58.625 150.430 ;
        RECT 58.795 150.385 59.085 150.615 ;
        RECT 59.700 150.570 60.020 150.630 ;
        RECT 65.310 150.570 65.450 150.770 ;
        RECT 66.140 150.710 66.460 150.770 ;
        RECT 67.060 150.710 67.380 150.970 ;
        RECT 59.700 150.430 65.450 150.570 ;
        RECT 57.860 150.230 58.180 150.290 ;
        RECT 58.870 150.230 59.010 150.385 ;
        RECT 59.700 150.370 60.020 150.430 ;
        RECT 65.680 150.370 66.000 150.630 ;
        RECT 85.460 150.370 85.780 150.630 ;
        RECT 65.770 150.230 65.910 150.370 ;
        RECT 56.570 150.090 65.910 150.230 ;
        RECT 54.655 150.045 54.945 150.090 ;
        RECT 57.860 150.030 58.180 150.090 ;
        RECT 59.255 149.890 59.545 149.935 ;
        RECT 56.110 149.750 59.545 149.890 ;
        RECT 52.800 149.550 53.120 149.610 ;
        RECT 56.110 149.550 56.250 149.750 ;
        RECT 59.255 149.705 59.545 149.750 ;
        RECT 62.460 149.890 62.780 149.950 ;
        RECT 67.075 149.890 67.365 149.935 ;
        RECT 62.460 149.750 67.365 149.890 ;
        RECT 62.460 149.690 62.780 149.750 ;
        RECT 67.075 149.705 67.365 149.750 ;
        RECT 79.940 149.890 80.260 149.950 ;
        RECT 84.555 149.890 84.845 149.935 ;
        RECT 79.940 149.750 84.845 149.890 ;
        RECT 79.940 149.690 80.260 149.750 ;
        RECT 84.555 149.705 84.845 149.750 ;
        RECT 49.210 149.410 56.250 149.550 ;
        RECT 56.480 149.550 56.800 149.610 ;
        RECT 57.875 149.550 58.165 149.595 ;
        RECT 64.760 149.550 65.080 149.610 ;
        RECT 56.480 149.410 65.080 149.550 ;
        RECT 33.035 149.365 33.325 149.410 ;
        RECT 33.480 149.350 33.800 149.410 ;
        RECT 52.800 149.350 53.120 149.410 ;
        RECT 56.480 149.350 56.800 149.410 ;
        RECT 57.875 149.365 58.165 149.410 ;
        RECT 64.760 149.350 65.080 149.410 ;
        RECT 15.930 148.730 87.230 149.210 ;
        RECT 33.480 148.330 33.800 148.590 ;
        RECT 36.715 148.530 37.005 148.575 ;
        RECT 37.160 148.530 37.480 148.590 ;
        RECT 36.715 148.390 37.480 148.530 ;
        RECT 36.715 148.345 37.005 148.390 ;
        RECT 37.160 148.330 37.480 148.390 ;
        RECT 39.000 148.530 39.320 148.590 ;
        RECT 44.995 148.530 45.285 148.575 ;
        RECT 55.100 148.530 55.420 148.590 ;
        RECT 39.000 148.390 55.420 148.530 ;
        RECT 39.000 148.330 39.320 148.390 ;
        RECT 44.995 148.345 45.285 148.390 ;
        RECT 55.100 148.330 55.420 148.390 ;
        RECT 57.875 148.530 58.165 148.575 ;
        RECT 58.780 148.530 59.100 148.590 ;
        RECT 57.875 148.390 59.100 148.530 ;
        RECT 57.875 148.345 58.165 148.390 ;
        RECT 58.780 148.330 59.100 148.390 ;
        RECT 59.255 148.530 59.545 148.575 ;
        RECT 59.700 148.530 60.020 148.590 ;
        RECT 59.255 148.390 60.020 148.530 ;
        RECT 59.255 148.345 59.545 148.390 ;
        RECT 59.700 148.330 60.020 148.390 ;
        RECT 60.635 148.530 60.925 148.575 ;
        RECT 61.080 148.530 61.400 148.590 ;
        RECT 60.635 148.390 61.400 148.530 ;
        RECT 60.635 148.345 60.925 148.390 ;
        RECT 32.115 147.850 32.405 147.895 ;
        RECT 35.795 147.850 36.085 147.895 ;
        RECT 36.700 147.850 37.020 147.910 ;
        RECT 32.115 147.710 34.630 147.850 ;
        RECT 32.115 147.665 32.405 147.710 ;
        RECT 31.640 147.310 31.960 147.570 ;
        RECT 34.490 147.555 34.630 147.710 ;
        RECT 35.795 147.710 37.020 147.850 ;
        RECT 35.795 147.665 36.085 147.710 ;
        RECT 36.700 147.650 37.020 147.710 ;
        RECT 55.560 147.850 55.880 147.910 ;
        RECT 56.035 147.850 56.325 147.895 ;
        RECT 60.710 147.850 60.850 148.345 ;
        RECT 61.080 148.330 61.400 148.390 ;
        RECT 84.540 148.330 84.860 148.590 ;
        RECT 64.760 147.990 65.080 148.250 ;
        RECT 55.560 147.710 56.325 147.850 ;
        RECT 55.560 147.650 55.880 147.710 ;
        RECT 56.035 147.665 56.325 147.710 ;
        RECT 58.410 147.710 62.690 147.850 ;
        RECT 32.575 147.325 32.865 147.555 ;
        RECT 33.035 147.325 33.325 147.555 ;
        RECT 34.415 147.325 34.705 147.555 ;
        RECT 34.875 147.510 35.165 147.555 ;
        RECT 37.620 147.510 37.940 147.570 ;
        RECT 34.875 147.370 37.940 147.510 ;
        RECT 34.875 147.325 35.165 147.370 ;
        RECT 32.650 146.830 32.790 147.325 ;
        RECT 33.110 147.170 33.250 147.325 ;
        RECT 37.620 147.310 37.940 147.370 ;
        RECT 38.080 147.310 38.400 147.570 ;
        RECT 38.540 147.310 38.860 147.570 ;
        RECT 39.015 147.325 39.305 147.555 ;
        RECT 33.940 147.170 34.260 147.230 ;
        RECT 39.090 147.170 39.230 147.325 ;
        RECT 39.920 147.310 40.240 147.570 ;
        RECT 43.140 147.310 43.460 147.570 ;
        RECT 44.520 147.510 44.840 147.570 ;
        RECT 45.455 147.510 45.745 147.555 ;
        RECT 44.520 147.370 45.745 147.510 ;
        RECT 44.520 147.310 44.840 147.370 ;
        RECT 45.455 147.325 45.745 147.370 ;
        RECT 53.260 147.510 53.580 147.570 ;
        RECT 58.410 147.555 58.550 147.710 ;
        RECT 56.495 147.510 56.785 147.555 ;
        RECT 53.260 147.370 56.785 147.510 ;
        RECT 53.260 147.310 53.580 147.370 ;
        RECT 56.495 147.325 56.785 147.370 ;
        RECT 58.335 147.325 58.625 147.555 ;
        RECT 59.240 147.510 59.560 147.570 ;
        RECT 62.550 147.555 62.690 147.710 ;
        RECT 59.715 147.510 60.005 147.555 ;
        RECT 59.240 147.370 60.005 147.510 ;
        RECT 59.240 147.310 59.560 147.370 ;
        RECT 59.715 147.325 60.005 147.370 ;
        RECT 62.015 147.325 62.305 147.555 ;
        RECT 62.475 147.510 62.765 147.555 ;
        RECT 62.920 147.510 63.240 147.570 ;
        RECT 62.475 147.370 63.240 147.510 ;
        RECT 62.475 147.325 62.765 147.370 ;
        RECT 33.110 147.030 39.230 147.170 ;
        RECT 58.780 147.170 59.100 147.230 ;
        RECT 62.090 147.170 62.230 147.325 ;
        RECT 62.920 147.310 63.240 147.370 ;
        RECT 63.840 147.310 64.160 147.570 ;
        RECT 58.780 147.030 62.230 147.170 ;
        RECT 33.940 146.970 34.260 147.030 ;
        RECT 58.780 146.970 59.100 147.030 ;
        RECT 85.000 146.970 85.320 147.230 ;
        RECT 38.080 146.830 38.400 146.890 ;
        RECT 32.650 146.690 38.400 146.830 ;
        RECT 38.080 146.630 38.400 146.690 ;
        RECT 15.930 146.010 87.230 146.490 ;
        RECT 33.940 145.610 34.260 145.870 ;
        RECT 43.140 145.810 43.460 145.870 ;
        RECT 40.010 145.670 43.460 145.810 ;
        RECT 31.640 145.470 31.960 145.530 ;
        RECT 35.795 145.470 36.085 145.515 ;
        RECT 38.540 145.470 38.860 145.530 ;
        RECT 40.010 145.515 40.150 145.670 ;
        RECT 43.140 145.610 43.460 145.670 ;
        RECT 31.640 145.330 38.860 145.470 ;
        RECT 31.640 145.270 31.960 145.330 ;
        RECT 35.795 145.285 36.085 145.330 ;
        RECT 38.540 145.270 38.860 145.330 ;
        RECT 39.935 145.285 40.225 145.515 ;
        RECT 42.235 145.470 42.525 145.515 ;
        RECT 44.520 145.470 44.840 145.530 ;
        RECT 42.235 145.330 44.840 145.470 ;
        RECT 42.235 145.285 42.525 145.330 ;
        RECT 26.580 145.130 26.900 145.190 ;
        RECT 35.335 145.130 35.625 145.175 ;
        RECT 26.580 144.990 35.625 145.130 ;
        RECT 26.580 144.930 26.900 144.990 ;
        RECT 35.335 144.945 35.625 144.990 ;
        RECT 36.715 145.130 37.005 145.175 ;
        RECT 39.015 145.130 39.305 145.175 ;
        RECT 42.310 145.130 42.450 145.285 ;
        RECT 44.520 145.270 44.840 145.330 ;
        RECT 57.860 145.470 58.180 145.530 ;
        RECT 60.635 145.470 60.925 145.515 ;
        RECT 57.860 145.330 60.925 145.470 ;
        RECT 57.860 145.270 58.180 145.330 ;
        RECT 60.635 145.285 60.925 145.330 ;
        RECT 36.715 144.990 42.450 145.130 ;
        RECT 42.680 145.130 43.000 145.190 ;
        RECT 43.155 145.130 43.445 145.175 ;
        RECT 42.680 144.990 43.445 145.130 ;
        RECT 36.715 144.945 37.005 144.990 ;
        RECT 39.015 144.945 39.305 144.990 ;
        RECT 33.480 144.790 33.800 144.850 ;
        RECT 33.955 144.790 34.245 144.835 ;
        RECT 33.480 144.650 34.245 144.790 ;
        RECT 35.410 144.790 35.550 144.945 ;
        RECT 42.680 144.930 43.000 144.990 ;
        RECT 43.155 144.945 43.445 144.990 ;
        RECT 44.075 145.130 44.365 145.175 ;
        RECT 47.280 145.130 47.600 145.190 ;
        RECT 44.075 144.990 47.600 145.130 ;
        RECT 44.075 144.945 44.365 144.990 ;
        RECT 47.280 144.930 47.600 144.990 ;
        RECT 61.555 144.945 61.845 145.175 ;
        RECT 37.635 144.790 37.925 144.835 ;
        RECT 58.780 144.790 59.100 144.850 ;
        RECT 61.630 144.790 61.770 144.945 ;
        RECT 62.920 144.930 63.240 145.190 ;
        RECT 63.840 144.930 64.160 145.190 ;
        RECT 35.410 144.650 61.770 144.790 ;
        RECT 33.480 144.590 33.800 144.650 ;
        RECT 33.955 144.605 34.245 144.650 ;
        RECT 37.635 144.605 37.925 144.650 ;
        RECT 34.030 144.450 34.170 144.605 ;
        RECT 58.780 144.590 59.100 144.650 ;
        RECT 85.460 144.590 85.780 144.850 ;
        RECT 40.855 144.450 41.145 144.495 ;
        RECT 55.560 144.450 55.880 144.510 ;
        RECT 34.030 144.310 41.145 144.450 ;
        RECT 40.855 144.265 41.145 144.310 ;
        RECT 44.610 144.310 55.880 144.450 ;
        RECT 34.875 144.110 35.165 144.155 ;
        RECT 40.380 144.110 40.700 144.170 ;
        RECT 44.610 144.110 44.750 144.310 ;
        RECT 55.560 144.250 55.880 144.310 ;
        RECT 34.875 143.970 44.750 144.110 ;
        RECT 44.995 144.110 45.285 144.155 ;
        RECT 46.360 144.110 46.680 144.170 ;
        RECT 44.995 143.970 46.680 144.110 ;
        RECT 34.875 143.925 35.165 143.970 ;
        RECT 40.380 143.910 40.700 143.970 ;
        RECT 44.995 143.925 45.285 143.970 ;
        RECT 46.360 143.910 46.680 143.970 ;
        RECT 15.930 143.290 87.230 143.770 ;
        RECT 33.495 143.090 33.785 143.135 ;
        RECT 34.400 143.090 34.720 143.150 ;
        RECT 33.495 142.950 34.720 143.090 ;
        RECT 33.495 142.905 33.785 142.950 ;
        RECT 34.400 142.890 34.720 142.950 ;
        RECT 38.080 143.090 38.400 143.150 ;
        RECT 39.015 143.090 39.305 143.135 ;
        RECT 38.080 142.950 39.305 143.090 ;
        RECT 38.080 142.890 38.400 142.950 ;
        RECT 39.015 142.905 39.305 142.950 ;
        RECT 40.855 143.090 41.145 143.135 ;
        RECT 42.680 143.090 43.000 143.150 ;
        RECT 40.855 142.950 43.000 143.090 ;
        RECT 40.855 142.905 41.145 142.950 ;
        RECT 42.680 142.890 43.000 142.950 ;
        RECT 43.140 143.090 43.460 143.150 ;
        RECT 44.075 143.090 44.365 143.135 ;
        RECT 43.140 142.950 44.365 143.090 ;
        RECT 43.140 142.890 43.460 142.950 ;
        RECT 44.075 142.905 44.365 142.950 ;
        RECT 37.635 142.750 37.925 142.795 ;
        RECT 41.760 142.750 42.080 142.810 ;
        RECT 37.635 142.610 42.080 142.750 ;
        RECT 37.635 142.565 37.925 142.610 ;
        RECT 41.760 142.550 42.080 142.610 ;
        RECT 40.380 142.410 40.700 142.470 ;
        RECT 38.630 142.270 40.700 142.410 ;
        RECT 23.360 142.070 23.680 142.130 ;
        RECT 23.835 142.070 24.125 142.115 ;
        RECT 23.360 141.930 24.125 142.070 ;
        RECT 23.360 141.870 23.680 141.930 ;
        RECT 23.835 141.885 24.125 141.930 ;
        RECT 33.020 142.070 33.340 142.130 ;
        RECT 34.415 142.070 34.705 142.115 ;
        RECT 33.020 141.930 34.705 142.070 ;
        RECT 33.020 141.870 33.340 141.930 ;
        RECT 34.415 141.885 34.705 141.930 ;
        RECT 36.700 141.870 37.020 142.130 ;
        RECT 38.630 142.115 38.770 142.270 ;
        RECT 40.380 142.210 40.700 142.270 ;
        RECT 38.555 141.885 38.845 142.115 ;
        RECT 39.475 141.885 39.765 142.115 ;
        RECT 39.550 141.730 39.690 141.885 ;
        RECT 39.920 141.870 40.240 142.130 ;
        RECT 43.140 142.070 43.460 142.130 ;
        RECT 40.470 141.930 43.460 142.070 ;
        RECT 40.470 141.730 40.610 141.930 ;
        RECT 43.140 141.870 43.460 141.930 ;
        RECT 46.360 141.870 46.680 142.130 ;
        RECT 39.550 141.590 40.610 141.730 ;
        RECT 42.680 141.730 43.000 141.790 ;
        RECT 43.615 141.730 43.905 141.775 ;
        RECT 42.680 141.590 43.905 141.730 ;
        RECT 42.680 141.530 43.000 141.590 ;
        RECT 43.615 141.545 43.905 141.590 ;
        RECT 45.900 141.390 46.220 141.450 ;
        RECT 47.295 141.390 47.585 141.435 ;
        RECT 45.900 141.250 47.585 141.390 ;
        RECT 45.900 141.190 46.220 141.250 ;
        RECT 47.295 141.205 47.585 141.250 ;
        RECT 15.930 140.570 87.230 141.050 ;
      LAYER met2 ;
        RECT 10.500 219.000 10.780 223.000 ;
        RECT 13.720 219.000 14.000 223.000 ;
        RECT 16.940 219.000 17.220 223.000 ;
        RECT 20.160 219.000 20.440 223.000 ;
        RECT 23.380 219.000 23.660 223.000 ;
        RECT 26.600 219.000 26.880 223.000 ;
        RECT 29.820 219.000 30.100 223.000 ;
        RECT 33.040 219.000 33.320 223.000 ;
        RECT 36.260 219.000 36.540 223.000 ;
        RECT 36.790 219.280 38.310 219.420 ;
        RECT 10.570 216.135 10.710 219.000 ;
        RECT 10.500 215.765 10.780 216.135 ;
        RECT 13.790 182.815 13.930 219.000 ;
        RECT 14.650 212.900 14.910 213.220 ;
        RECT 14.710 193.580 14.850 212.900 ;
        RECT 15.560 211.685 15.840 212.055 ;
        RECT 15.630 208.460 15.770 211.685 ;
        RECT 17.010 209.900 17.150 219.000 ;
        RECT 19.710 215.620 19.970 215.940 ;
        RECT 17.410 213.580 17.670 213.900 ;
        RECT 16.550 209.760 17.150 209.900 ;
        RECT 15.570 208.140 15.830 208.460 ;
        RECT 15.110 206.780 15.370 207.100 ;
        RECT 15.170 199.700 15.310 206.780 ;
        RECT 16.030 206.440 16.290 206.760 ;
        RECT 15.570 202.360 15.830 202.680 ;
        RECT 15.630 201.855 15.770 202.360 ;
        RECT 15.560 201.485 15.840 201.855 ;
        RECT 15.170 199.560 15.770 199.700 ;
        RECT 15.100 194.685 15.380 195.055 ;
        RECT 15.170 194.520 15.310 194.685 ;
        RECT 15.110 194.200 15.370 194.520 ;
        RECT 14.710 193.440 15.310 193.580 ;
        RECT 14.650 192.840 14.910 193.160 ;
        RECT 14.710 192.335 14.850 192.840 ;
        RECT 14.640 191.965 14.920 192.335 ;
        RECT 14.640 189.245 14.920 189.615 ;
        RECT 14.650 189.100 14.910 189.245 ;
        RECT 13.720 182.445 14.000 182.815 ;
        RECT 15.170 177.520 15.310 193.440 ;
        RECT 15.630 178.200 15.770 199.560 ;
        RECT 16.090 183.300 16.230 206.440 ;
        RECT 16.550 205.740 16.690 209.760 ;
        RECT 16.940 208.285 17.220 208.655 ;
        RECT 16.490 205.420 16.750 205.740 ;
        RECT 16.480 204.885 16.760 205.255 ;
        RECT 16.550 183.980 16.690 204.885 ;
        RECT 16.490 183.660 16.750 183.980 ;
        RECT 16.030 182.980 16.290 183.300 ;
        RECT 17.010 182.620 17.150 208.285 ;
        RECT 17.470 191.800 17.610 213.580 ;
        RECT 18.780 212.365 19.060 212.735 ;
        RECT 18.850 210.500 18.990 212.365 ;
        RECT 19.770 211.180 19.910 215.620 ;
        RECT 20.230 213.220 20.370 219.000 ;
        RECT 20.620 218.485 20.900 218.855 ;
        RECT 20.170 212.900 20.430 213.220 ;
        RECT 19.710 210.860 19.970 211.180 ;
        RECT 18.790 210.180 19.050 210.500 ;
        RECT 19.710 207.800 19.970 208.120 ;
        RECT 19.250 207.295 19.510 207.440 ;
        RECT 19.240 206.925 19.520 207.295 ;
        RECT 19.250 206.440 19.510 206.760 ;
        RECT 19.310 205.060 19.450 206.440 ;
        RECT 19.770 205.740 19.910 207.800 ;
        RECT 19.710 205.420 19.970 205.740 ;
        RECT 18.330 204.740 18.590 205.060 ;
        RECT 19.250 204.740 19.510 205.060 ;
        RECT 17.870 198.455 18.130 198.600 ;
        RECT 17.860 198.085 18.140 198.455 ;
        RECT 17.870 193.520 18.130 193.840 ;
        RECT 17.410 191.480 17.670 191.800 ;
        RECT 17.410 185.360 17.670 185.680 ;
        RECT 17.470 184.855 17.610 185.360 ;
        RECT 17.400 184.485 17.680 184.855 ;
        RECT 16.950 182.300 17.210 182.620 ;
        RECT 15.570 177.880 15.830 178.200 ;
        RECT 17.400 177.685 17.680 178.055 ;
        RECT 17.410 177.540 17.670 177.685 ;
        RECT 15.110 177.200 15.370 177.520 ;
        RECT 17.930 175.140 18.070 193.520 ;
        RECT 18.390 182.280 18.530 204.740 ;
        RECT 19.710 201.680 19.970 202.000 ;
        RECT 18.790 199.300 19.050 199.620 ;
        RECT 18.850 194.860 18.990 199.300 ;
        RECT 19.770 196.560 19.910 201.680 ;
        RECT 20.170 201.000 20.430 201.320 ;
        RECT 20.230 196.900 20.370 201.000 ;
        RECT 20.690 200.300 20.830 218.485 ;
        RECT 22.470 214.600 22.730 214.920 ;
        RECT 22.010 211.880 22.270 212.200 ;
        RECT 21.080 211.005 21.360 211.375 ;
        RECT 21.150 200.300 21.290 211.005 ;
        RECT 22.070 205.060 22.210 211.880 ;
        RECT 21.550 204.740 21.810 205.060 ;
        RECT 22.010 204.740 22.270 205.060 ;
        RECT 21.610 203.215 21.750 204.740 ;
        RECT 21.540 202.845 21.820 203.215 ;
        RECT 22.530 203.020 22.670 214.600 ;
        RECT 22.930 213.920 23.190 214.240 ;
        RECT 22.990 211.180 23.130 213.920 ;
        RECT 23.450 213.415 23.590 219.000 ;
        RECT 24.310 214.260 24.570 214.580 ;
        RECT 23.380 213.045 23.660 213.415 ;
        RECT 22.930 210.860 23.190 211.180 ;
        RECT 24.370 210.840 24.510 214.260 ;
        RECT 24.310 210.520 24.570 210.840 ;
        RECT 23.850 210.180 24.110 210.500 ;
        RECT 23.910 210.015 24.050 210.180 ;
        RECT 23.840 209.645 24.120 210.015 ;
        RECT 23.390 207.800 23.650 208.120 ;
        RECT 23.450 206.760 23.590 207.800 ;
        RECT 24.370 207.440 24.510 210.520 ;
        RECT 25.230 210.180 25.490 210.500 ;
        RECT 24.770 208.140 25.030 208.460 ;
        RECT 24.310 207.120 24.570 207.440 ;
        RECT 23.390 206.440 23.650 206.760 ;
        RECT 23.840 206.245 24.120 206.615 ;
        RECT 23.380 205.565 23.660 205.935 ;
        RECT 23.910 205.740 24.050 206.245 ;
        RECT 22.470 202.700 22.730 203.020 ;
        RECT 23.450 202.000 23.590 205.565 ;
        RECT 23.850 205.420 24.110 205.740 ;
        RECT 24.310 204.740 24.570 205.060 ;
        RECT 23.850 203.720 24.110 204.040 ;
        RECT 21.550 201.680 21.810 202.000 ;
        RECT 22.930 201.855 23.190 202.000 ;
        RECT 20.630 199.980 20.890 200.300 ;
        RECT 21.090 199.980 21.350 200.300 ;
        RECT 20.170 196.580 20.430 196.900 ;
        RECT 19.710 196.240 19.970 196.560 ;
        RECT 19.250 195.900 19.510 196.220 ;
        RECT 18.790 194.540 19.050 194.860 ;
        RECT 18.790 193.860 19.050 194.180 ;
        RECT 18.850 191.120 18.990 193.860 ;
        RECT 19.310 193.160 19.450 195.900 ;
        RECT 19.250 192.840 19.510 193.160 ;
        RECT 18.790 190.800 19.050 191.120 ;
        RECT 18.790 190.120 19.050 190.440 ;
        RECT 18.850 188.740 18.990 190.120 ;
        RECT 18.790 188.420 19.050 188.740 ;
        RECT 18.790 183.320 19.050 183.640 ;
        RECT 18.330 181.960 18.590 182.280 ;
        RECT 18.850 181.340 18.990 183.320 ;
        RECT 19.310 182.870 19.450 192.840 ;
        RECT 19.770 186.700 19.910 196.240 ;
        RECT 20.230 191.540 20.370 196.580 ;
        RECT 20.630 195.900 20.890 196.220 ;
        RECT 20.690 193.160 20.830 195.900 ;
        RECT 21.090 194.540 21.350 194.860 ;
        RECT 20.630 192.840 20.890 193.160 ;
        RECT 20.230 191.400 20.830 191.540 ;
        RECT 20.170 190.800 20.430 191.120 ;
        RECT 19.710 186.380 19.970 186.700 ;
        RECT 19.710 182.870 19.970 182.960 ;
        RECT 19.310 182.730 19.970 182.870 ;
        RECT 19.710 182.640 19.970 182.730 ;
        RECT 18.390 181.200 18.990 181.340 ;
        RECT 18.390 176.840 18.530 181.200 ;
        RECT 20.230 180.240 20.370 190.800 ;
        RECT 20.690 189.615 20.830 191.400 ;
        RECT 21.150 191.120 21.290 194.540 ;
        RECT 21.610 192.140 21.750 201.680 ;
        RECT 22.920 201.485 23.200 201.855 ;
        RECT 23.390 201.680 23.650 202.000 ;
        RECT 23.390 201.000 23.650 201.320 ;
        RECT 22.470 199.640 22.730 199.960 ;
        RECT 22.010 198.960 22.270 199.280 ;
        RECT 21.550 191.820 21.810 192.140 ;
        RECT 21.090 190.800 21.350 191.120 ;
        RECT 20.620 189.245 20.900 189.615 ;
        RECT 22.070 189.420 22.210 198.960 ;
        RECT 22.530 196.470 22.670 199.640 ;
        RECT 23.450 199.620 23.590 201.000 ;
        RECT 22.930 199.300 23.190 199.620 ;
        RECT 23.390 199.300 23.650 199.620 ;
        RECT 22.990 197.580 23.130 199.300 ;
        RECT 22.930 197.260 23.190 197.580 ;
        RECT 23.450 197.240 23.590 199.300 ;
        RECT 23.390 196.920 23.650 197.240 ;
        RECT 22.930 196.470 23.190 196.560 ;
        RECT 22.530 196.330 23.190 196.470 ;
        RECT 22.930 196.240 23.190 196.330 ;
        RECT 22.460 195.365 22.740 195.735 ;
        RECT 22.530 194.180 22.670 195.365 ;
        RECT 22.470 193.860 22.730 194.180 ;
        RECT 22.990 193.750 23.130 196.240 ;
        RECT 23.380 194.685 23.660 195.055 ;
        RECT 23.390 194.540 23.650 194.685 ;
        RECT 23.390 193.750 23.650 193.840 ;
        RECT 22.990 193.610 23.650 193.750 ;
        RECT 22.990 191.460 23.130 193.610 ;
        RECT 23.390 193.520 23.650 193.610 ;
        RECT 23.910 193.580 24.050 203.720 ;
        RECT 24.370 203.215 24.510 204.740 ;
        RECT 24.300 202.845 24.580 203.215 ;
        RECT 24.310 201.340 24.570 201.660 ;
        RECT 24.370 201.175 24.510 201.340 ;
        RECT 24.830 201.320 24.970 208.140 ;
        RECT 25.290 207.100 25.430 210.180 ;
        RECT 26.150 209.160 26.410 209.480 ;
        RECT 26.210 207.975 26.350 209.160 ;
        RECT 26.140 207.605 26.420 207.975 ;
        RECT 26.150 207.120 26.410 207.440 ;
        RECT 25.230 206.780 25.490 207.100 ;
        RECT 25.690 206.780 25.950 207.100 ;
        RECT 25.290 204.720 25.430 206.780 ;
        RECT 25.750 205.740 25.890 206.780 ;
        RECT 25.690 205.420 25.950 205.740 ;
        RECT 25.680 204.885 25.960 205.255 ;
        RECT 26.210 205.060 26.350 207.120 ;
        RECT 25.690 204.740 25.950 204.885 ;
        RECT 26.150 204.740 26.410 205.060 ;
        RECT 25.230 204.400 25.490 204.720 ;
        RECT 26.210 204.460 26.350 204.740 ;
        RECT 25.750 204.320 26.350 204.460 ;
        RECT 25.220 203.525 25.500 203.895 ;
        RECT 25.290 201.320 25.430 203.525 ;
        RECT 24.300 200.805 24.580 201.175 ;
        RECT 24.770 201.000 25.030 201.320 ;
        RECT 25.230 201.000 25.490 201.320 ;
        RECT 25.750 200.495 25.890 204.320 ;
        RECT 26.150 203.720 26.410 204.040 ;
        RECT 25.680 200.125 25.960 200.495 ;
        RECT 25.230 199.870 25.490 199.960 ;
        RECT 25.230 199.730 25.890 199.870 ;
        RECT 25.230 199.640 25.490 199.730 ;
        RECT 24.310 199.300 24.570 199.620 ;
        RECT 24.370 196.900 24.510 199.300 ;
        RECT 25.230 198.960 25.490 199.280 ;
        RECT 24.760 197.405 25.040 197.775 ;
        RECT 24.310 196.580 24.570 196.900 ;
        RECT 24.830 195.880 24.970 197.405 ;
        RECT 25.290 196.560 25.430 198.960 ;
        RECT 25.750 197.775 25.890 199.730 ;
        RECT 26.210 199.280 26.350 203.720 ;
        RECT 26.150 198.960 26.410 199.280 ;
        RECT 25.680 197.405 25.960 197.775 ;
        RECT 25.230 196.470 25.490 196.560 ;
        RECT 25.230 196.330 25.890 196.470 ;
        RECT 25.230 196.240 25.490 196.330 ;
        RECT 24.770 195.560 25.030 195.880 ;
        RECT 25.230 195.560 25.490 195.880 ;
        RECT 25.290 194.180 25.430 195.560 ;
        RECT 25.750 194.860 25.890 196.330 ;
        RECT 26.150 196.240 26.410 196.560 ;
        RECT 26.670 196.415 26.810 219.000 ;
        RECT 29.360 213.725 29.640 214.095 ;
        RECT 29.890 213.900 30.030 219.000 ;
        RECT 30.290 214.260 30.550 214.580 ;
        RECT 27.980 213.045 28.260 213.415 ;
        RECT 27.530 212.560 27.790 212.880 ;
        RECT 27.070 210.860 27.330 211.180 ;
        RECT 27.130 208.460 27.270 210.860 ;
        RECT 27.590 210.500 27.730 212.560 ;
        RECT 27.530 210.180 27.790 210.500 ;
        RECT 28.050 209.480 28.190 213.045 ;
        RECT 28.910 212.220 29.170 212.540 ;
        RECT 28.440 210.325 28.720 210.695 ;
        RECT 28.450 210.180 28.710 210.325 ;
        RECT 28.970 210.160 29.110 212.220 ;
        RECT 28.910 209.840 29.170 210.160 ;
        RECT 29.430 209.820 29.570 213.725 ;
        RECT 29.830 213.580 30.090 213.900 ;
        RECT 29.830 209.840 30.090 210.160 ;
        RECT 29.370 209.500 29.630 209.820 ;
        RECT 27.990 209.160 28.250 209.480 ;
        RECT 28.450 209.160 28.710 209.480 ;
        RECT 27.070 208.140 27.330 208.460 ;
        RECT 27.530 207.800 27.790 208.120 ;
        RECT 27.060 206.925 27.340 207.295 ;
        RECT 27.130 197.580 27.270 206.925 ;
        RECT 27.590 204.040 27.730 207.800 ;
        RECT 28.510 207.780 28.650 209.160 ;
        RECT 29.370 208.140 29.630 208.460 ;
        RECT 28.450 207.460 28.710 207.780 ;
        RECT 27.990 207.120 28.250 207.440 ;
        RECT 28.050 206.615 28.190 207.120 ;
        RECT 27.980 206.245 28.260 206.615 ;
        RECT 28.910 206.440 29.170 206.760 ;
        RECT 28.450 205.255 28.710 205.400 ;
        RECT 28.440 204.885 28.720 205.255 ;
        RECT 28.970 205.060 29.110 206.440 ;
        RECT 28.910 204.740 29.170 205.060 ;
        RECT 27.990 204.060 28.250 204.380 ;
        RECT 27.530 203.720 27.790 204.040 ;
        RECT 27.530 202.020 27.790 202.340 ;
        RECT 27.070 197.260 27.330 197.580 ;
        RECT 25.690 194.540 25.950 194.860 ;
        RECT 25.230 193.860 25.490 194.180 ;
        RECT 23.910 193.440 24.970 193.580 ;
        RECT 24.310 192.840 24.570 193.160 ;
        RECT 23.850 191.710 24.110 191.800 ;
        RECT 23.450 191.570 24.110 191.710 ;
        RECT 22.930 191.140 23.190 191.460 ;
        RECT 22.920 190.605 23.200 190.975 ;
        RECT 22.470 190.120 22.730 190.440 ;
        RECT 22.010 189.100 22.270 189.420 ;
        RECT 21.550 188.990 21.810 189.080 ;
        RECT 20.690 188.850 21.810 188.990 ;
        RECT 20.690 185.680 20.830 188.850 ;
        RECT 21.550 188.760 21.810 188.850 ;
        RECT 22.070 188.740 22.210 189.100 ;
        RECT 22.530 188.740 22.670 190.120 ;
        RECT 22.010 188.420 22.270 188.740 ;
        RECT 22.470 188.420 22.730 188.740 ;
        RECT 22.070 186.360 22.210 188.420 ;
        RECT 22.010 186.040 22.270 186.360 ;
        RECT 20.630 185.590 20.890 185.680 ;
        RECT 20.630 185.450 21.290 185.590 ;
        RECT 20.630 185.360 20.890 185.450 ;
        RECT 20.620 183.125 20.900 183.495 ;
        RECT 20.630 182.980 20.890 183.125 ;
        RECT 21.150 181.260 21.290 185.450 ;
        RECT 22.070 185.340 22.210 186.040 ;
        RECT 22.530 185.680 22.670 188.420 ;
        RECT 22.990 188.400 23.130 190.605 ;
        RECT 22.930 188.080 23.190 188.400 ;
        RECT 23.450 188.060 23.590 191.570 ;
        RECT 23.850 191.480 24.110 191.570 ;
        RECT 24.370 190.780 24.510 192.840 ;
        RECT 24.310 190.690 24.570 190.780 ;
        RECT 23.910 190.550 24.570 190.690 ;
        RECT 23.910 189.420 24.050 190.550 ;
        RECT 24.310 190.460 24.570 190.550 ;
        RECT 23.850 189.100 24.110 189.420 ;
        RECT 24.300 189.245 24.580 189.615 ;
        RECT 23.390 187.740 23.650 188.060 ;
        RECT 23.450 186.020 23.590 187.740 ;
        RECT 23.390 185.700 23.650 186.020 ;
        RECT 22.470 185.360 22.730 185.680 ;
        RECT 22.010 185.020 22.270 185.340 ;
        RECT 22.530 183.980 22.670 185.360 ;
        RECT 23.910 185.000 24.050 189.100 ;
        RECT 24.370 188.400 24.510 189.245 ;
        RECT 24.310 188.080 24.570 188.400 ;
        RECT 23.850 184.680 24.110 185.000 ;
        RECT 22.470 183.660 22.730 183.980 ;
        RECT 23.840 183.805 24.120 184.175 ;
        RECT 21.090 180.940 21.350 181.260 ;
        RECT 20.170 179.920 20.430 180.240 ;
        RECT 19.710 179.240 19.970 179.560 ;
        RECT 20.170 179.240 20.430 179.560 ;
        RECT 19.770 177.860 19.910 179.240 ;
        RECT 19.710 177.540 19.970 177.860 ;
        RECT 18.330 176.520 18.590 176.840 ;
        RECT 17.870 174.820 18.130 175.140 ;
        RECT 18.390 171.935 18.530 176.520 ;
        RECT 19.250 174.480 19.510 174.800 ;
        RECT 18.320 171.565 18.600 171.935 ;
        RECT 19.310 170.380 19.450 174.480 ;
        RECT 19.250 170.060 19.510 170.380 ;
        RECT 19.250 168.360 19.510 168.680 ;
        RECT 17.860 160.685 18.140 161.055 ;
        RECT 17.870 160.540 18.130 160.685 ;
        RECT 19.310 159.500 19.450 168.360 ;
        RECT 20.230 167.660 20.370 179.240 ;
        RECT 20.630 174.820 20.890 175.140 ;
        RECT 20.690 173.100 20.830 174.820 ;
        RECT 20.630 172.780 20.890 173.100 ;
        RECT 21.150 172.500 21.290 180.940 ;
        RECT 22.530 179.900 22.670 183.660 ;
        RECT 23.910 183.300 24.050 183.805 ;
        RECT 22.930 182.980 23.190 183.300 ;
        RECT 23.850 182.980 24.110 183.300 ;
        RECT 22.990 182.280 23.130 182.980 ;
        RECT 22.930 181.960 23.190 182.280 ;
        RECT 23.910 180.240 24.050 182.980 ;
        RECT 24.370 182.700 24.510 188.080 ;
        RECT 24.830 183.300 24.970 193.440 ;
        RECT 26.210 193.160 26.350 196.240 ;
        RECT 26.600 196.045 26.880 196.415 ;
        RECT 27.070 195.900 27.330 196.220 ;
        RECT 26.610 193.860 26.870 194.180 ;
        RECT 26.670 193.500 26.810 193.860 ;
        RECT 26.610 193.180 26.870 193.500 ;
        RECT 26.150 192.840 26.410 193.160 ;
        RECT 26.670 191.655 26.810 193.180 ;
        RECT 27.130 192.140 27.270 195.900 ;
        RECT 27.070 191.820 27.330 192.140 ;
        RECT 26.600 191.285 26.880 191.655 ;
        RECT 26.610 191.030 26.870 191.120 ;
        RECT 27.130 191.030 27.270 191.820 ;
        RECT 27.590 191.370 27.730 202.020 ;
        RECT 28.050 192.335 28.190 204.060 ;
        RECT 28.450 203.720 28.710 204.040 ;
        RECT 28.910 203.720 29.170 204.040 ;
        RECT 28.510 197.580 28.650 203.720 ;
        RECT 28.450 197.260 28.710 197.580 ;
        RECT 28.440 196.725 28.720 197.095 ;
        RECT 28.510 196.560 28.650 196.725 ;
        RECT 28.450 196.240 28.710 196.560 ;
        RECT 28.450 195.560 28.710 195.880 ;
        RECT 28.510 194.520 28.650 195.560 ;
        RECT 28.450 194.200 28.710 194.520 ;
        RECT 27.980 191.965 28.260 192.335 ;
        RECT 27.590 191.230 28.650 191.370 ;
        RECT 26.610 190.890 27.270 191.030 ;
        RECT 26.610 190.800 26.870 190.890 ;
        RECT 26.150 190.120 26.410 190.440 ;
        RECT 26.210 188.740 26.350 190.120 ;
        RECT 26.150 188.420 26.410 188.740 ;
        RECT 25.690 187.400 25.950 187.720 ;
        RECT 25.750 186.360 25.890 187.400 ;
        RECT 25.230 186.215 25.490 186.360 ;
        RECT 25.220 185.845 25.500 186.215 ;
        RECT 25.690 186.040 25.950 186.360 ;
        RECT 26.210 186.020 26.350 188.420 ;
        RECT 26.150 185.700 26.410 186.020 ;
        RECT 25.680 185.165 25.960 185.535 ;
        RECT 25.750 183.980 25.890 185.165 ;
        RECT 26.150 184.680 26.410 185.000 ;
        RECT 25.690 183.660 25.950 183.980 ;
        RECT 24.770 182.980 25.030 183.300 ;
        RECT 25.690 182.980 25.950 183.300 ;
        RECT 25.750 182.815 25.890 182.980 ;
        RECT 24.370 182.560 24.970 182.700 ;
        RECT 24.310 181.960 24.570 182.280 ;
        RECT 24.370 180.920 24.510 181.960 ;
        RECT 24.830 181.260 24.970 182.560 ;
        RECT 25.680 182.445 25.960 182.815 ;
        RECT 25.680 181.765 25.960 182.135 ;
        RECT 24.770 180.940 25.030 181.260 ;
        RECT 24.310 180.600 24.570 180.920 ;
        RECT 25.230 180.600 25.490 180.920 ;
        RECT 24.770 180.260 25.030 180.580 ;
        RECT 23.850 179.920 24.110 180.240 ;
        RECT 22.470 179.580 22.730 179.900 ;
        RECT 23.910 178.300 24.050 179.920 ;
        RECT 23.450 178.160 24.050 178.300 ;
        RECT 22.470 177.540 22.730 177.860 ;
        RECT 22.930 177.540 23.190 177.860 ;
        RECT 21.550 176.860 21.810 177.180 ;
        RECT 21.610 173.100 21.750 176.860 ;
        RECT 22.530 176.840 22.670 177.540 ;
        RECT 22.470 176.520 22.730 176.840 ;
        RECT 22.530 175.140 22.670 176.520 ;
        RECT 22.470 174.820 22.730 175.140 ;
        RECT 21.550 172.780 21.810 173.100 ;
        RECT 20.690 172.360 21.290 172.500 ;
        RECT 20.170 167.340 20.430 167.660 ;
        RECT 20.230 163.920 20.370 167.340 ;
        RECT 20.170 163.600 20.430 163.920 ;
        RECT 20.690 162.220 20.830 172.360 ;
        RECT 21.610 169.700 21.750 172.780 ;
        RECT 22.010 171.760 22.270 172.080 ;
        RECT 22.470 171.760 22.730 172.080 ;
        RECT 21.550 169.380 21.810 169.700 ;
        RECT 21.090 169.040 21.350 169.360 ;
        RECT 21.150 166.640 21.290 169.040 ;
        RECT 22.070 168.680 22.210 171.760 ;
        RECT 22.530 169.700 22.670 171.760 ;
        RECT 22.470 169.380 22.730 169.700 ;
        RECT 22.010 168.360 22.270 168.680 ;
        RECT 21.550 166.660 21.810 166.980 ;
        RECT 21.090 166.320 21.350 166.640 ;
        RECT 21.150 164.260 21.290 166.320 ;
        RECT 21.090 163.940 21.350 164.260 ;
        RECT 21.610 163.240 21.750 166.660 ;
        RECT 21.550 162.920 21.810 163.240 ;
        RECT 20.630 161.900 20.890 162.220 ;
        RECT 19.710 161.220 19.970 161.540 ;
        RECT 19.250 159.180 19.510 159.500 ;
        RECT 19.770 157.655 19.910 161.220 ;
        RECT 20.170 160.200 20.430 160.520 ;
        RECT 20.230 159.160 20.370 160.200 ;
        RECT 21.610 159.500 21.750 162.920 ;
        RECT 22.470 161.900 22.730 162.220 ;
        RECT 21.550 159.180 21.810 159.500 ;
        RECT 20.170 158.840 20.430 159.160 ;
        RECT 22.530 158.820 22.670 161.900 ;
        RECT 22.470 158.500 22.730 158.820 ;
        RECT 19.700 157.285 19.980 157.655 ;
        RECT 17.410 155.440 17.670 155.760 ;
        RECT 17.470 154.935 17.610 155.440 ;
        RECT 17.400 154.565 17.680 154.935 ;
        RECT 22.990 154.060 23.130 177.540 ;
        RECT 23.450 156.780 23.590 178.160 ;
        RECT 24.830 177.860 24.970 180.260 ;
        RECT 24.770 177.540 25.030 177.860 ;
        RECT 25.290 167.175 25.430 180.600 ;
        RECT 25.750 175.220 25.890 181.765 ;
        RECT 26.210 180.920 26.350 184.680 ;
        RECT 26.150 180.600 26.410 180.920 ;
        RECT 26.140 179.725 26.420 180.095 ;
        RECT 26.210 177.180 26.350 179.725 ;
        RECT 26.150 176.860 26.410 177.180 ;
        RECT 25.750 175.080 26.350 175.220 ;
        RECT 25.690 174.480 25.950 174.800 ;
        RECT 25.750 172.760 25.890 174.480 ;
        RECT 25.690 172.440 25.950 172.760 ;
        RECT 25.220 166.805 25.500 167.175 ;
        RECT 25.750 166.980 25.890 172.440 ;
        RECT 26.210 167.740 26.350 175.080 ;
        RECT 26.670 174.800 26.810 190.800 ;
        RECT 27.990 190.460 28.250 190.780 ;
        RECT 27.070 190.120 27.330 190.440 ;
        RECT 27.130 186.700 27.270 190.120 ;
        RECT 28.050 189.330 28.190 190.460 ;
        RECT 27.590 189.190 28.190 189.330 ;
        RECT 27.070 186.380 27.330 186.700 ;
        RECT 27.590 185.000 27.730 189.190 ;
        RECT 28.510 188.740 28.650 191.230 ;
        RECT 27.990 188.420 28.250 188.740 ;
        RECT 28.450 188.420 28.710 188.740 ;
        RECT 28.050 186.215 28.190 188.420 ;
        RECT 27.980 185.845 28.260 186.215 ;
        RECT 27.060 184.485 27.340 184.855 ;
        RECT 27.530 184.680 27.790 185.000 ;
        RECT 27.130 183.300 27.270 184.485 ;
        RECT 27.070 182.980 27.330 183.300 ;
        RECT 27.070 181.960 27.330 182.280 ;
        RECT 27.130 181.260 27.270 181.960 ;
        RECT 27.070 180.940 27.330 181.260 ;
        RECT 27.130 179.560 27.270 180.940 ;
        RECT 27.070 179.240 27.330 179.560 ;
        RECT 26.610 174.710 26.870 174.800 ;
        RECT 26.610 174.570 27.270 174.710 ;
        RECT 26.610 174.480 26.870 174.570 ;
        RECT 26.610 173.800 26.870 174.120 ;
        RECT 26.670 172.420 26.810 173.800 ;
        RECT 27.130 172.420 27.270 174.570 ;
        RECT 27.590 173.180 27.730 184.680 ;
        RECT 27.980 183.805 28.260 184.175 ;
        RECT 28.510 183.980 28.650 188.420 ;
        RECT 28.970 186.360 29.110 203.720 ;
        RECT 29.430 202.680 29.570 208.140 ;
        RECT 29.890 204.720 30.030 209.840 ;
        RECT 29.830 204.400 30.090 204.720 ;
        RECT 29.820 202.845 30.100 203.215 ;
        RECT 29.370 202.360 29.630 202.680 ;
        RECT 29.890 202.340 30.030 202.845 ;
        RECT 29.830 202.020 30.090 202.340 ;
        RECT 29.370 201.340 29.630 201.660 ;
        RECT 29.430 199.960 29.570 201.340 ;
        RECT 29.890 200.300 30.030 202.020 ;
        RECT 30.350 202.000 30.490 214.260 ;
        RECT 33.110 213.220 33.250 219.000 ;
        RECT 36.330 218.740 36.470 219.000 ;
        RECT 36.790 218.740 36.930 219.280 ;
        RECT 36.330 218.600 36.930 218.740 ;
        RECT 34.430 213.580 34.690 213.900 ;
        RECT 33.050 212.900 33.310 213.220 ;
        RECT 33.040 211.005 33.320 211.375 ;
        RECT 33.110 210.160 33.250 211.005 ;
        RECT 34.490 210.500 34.630 213.580 ;
        RECT 37.640 212.365 37.920 212.735 ;
        RECT 34.780 211.345 36.320 211.715 ;
        RECT 36.720 211.090 37.000 211.375 ;
        RECT 35.410 211.005 37.000 211.090 ;
        RECT 35.410 210.950 36.930 211.005 ;
        RECT 34.890 210.520 35.150 210.840 ;
        RECT 34.430 210.180 34.690 210.500 ;
        RECT 31.670 210.015 31.930 210.160 ;
        RECT 30.750 209.500 31.010 209.820 ;
        RECT 31.660 209.645 31.940 210.015 ;
        RECT 33.050 209.840 33.310 210.160 ;
        RECT 33.510 209.500 33.770 209.820 ;
        RECT 30.810 208.370 30.950 209.500 ;
        RECT 31.480 208.625 33.020 208.995 ;
        RECT 30.810 208.230 32.790 208.370 ;
        RECT 32.130 207.460 32.390 207.780 ;
        RECT 31.670 207.120 31.930 207.440 ;
        RECT 30.750 206.440 31.010 206.760 ;
        RECT 30.810 202.535 30.950 206.440 ;
        RECT 31.210 204.740 31.470 205.060 ;
        RECT 31.270 204.380 31.410 204.740 ;
        RECT 31.730 204.575 31.870 207.120 ;
        RECT 32.190 205.400 32.330 207.460 ;
        RECT 32.650 205.400 32.790 208.230 ;
        RECT 33.050 208.140 33.310 208.460 ;
        RECT 33.110 206.760 33.250 208.140 ;
        RECT 33.050 206.440 33.310 206.760 ;
        RECT 32.130 205.080 32.390 205.400 ;
        RECT 32.590 205.080 32.850 205.400 ;
        RECT 31.210 204.060 31.470 204.380 ;
        RECT 31.660 204.205 31.940 204.575 ;
        RECT 31.480 203.185 33.020 203.555 ;
        RECT 30.740 202.165 31.020 202.535 ;
        RECT 31.210 202.360 31.470 202.680 ;
        RECT 30.290 201.680 30.550 202.000 ;
        RECT 30.290 201.230 30.550 201.320 ;
        RECT 31.270 201.230 31.410 202.360 ;
        RECT 31.660 202.165 31.940 202.535 ;
        RECT 31.730 202.000 31.870 202.165 ;
        RECT 31.670 201.680 31.930 202.000 ;
        RECT 32.130 201.680 32.390 202.000 ;
        RECT 33.570 201.855 33.710 209.500 ;
        RECT 34.950 208.540 35.090 210.520 ;
        RECT 35.410 210.015 35.550 210.950 ;
        RECT 37.710 210.500 37.850 212.365 ;
        RECT 35.810 210.180 36.070 210.500 ;
        RECT 36.270 210.180 36.530 210.500 ;
        RECT 37.650 210.180 37.910 210.500 ;
        RECT 35.340 209.645 35.620 210.015 ;
        RECT 35.870 209.335 36.010 210.180 ;
        RECT 36.330 210.015 36.470 210.180 ;
        RECT 36.260 209.645 36.540 210.015 ;
        RECT 36.730 209.840 36.990 210.160 ;
        RECT 35.800 208.965 36.080 209.335 ;
        RECT 34.950 208.400 36.010 208.540 ;
        RECT 34.030 207.550 35.090 207.690 ;
        RECT 35.340 207.605 35.620 207.975 ;
        RECT 34.030 205.935 34.170 207.550 ;
        RECT 34.430 206.780 34.690 207.100 ;
        RECT 33.960 205.565 34.240 205.935 ;
        RECT 33.970 204.400 34.230 204.720 ;
        RECT 34.030 203.215 34.170 204.400 ;
        RECT 34.490 203.895 34.630 206.780 ;
        RECT 34.950 206.670 35.090 207.550 ;
        RECT 35.410 207.440 35.550 207.605 ;
        RECT 35.870 207.440 36.010 208.400 ;
        RECT 36.790 207.780 36.930 209.840 ;
        RECT 37.190 209.160 37.450 209.480 ;
        RECT 36.730 207.460 36.990 207.780 ;
        RECT 35.350 207.120 35.610 207.440 ;
        RECT 35.810 207.120 36.070 207.440 ;
        RECT 34.950 206.530 36.930 206.670 ;
        RECT 37.250 206.615 37.390 209.160 ;
        RECT 37.710 207.440 37.850 210.180 ;
        RECT 37.650 207.120 37.910 207.440 ;
        RECT 34.780 205.905 36.320 206.275 ;
        RECT 36.790 205.935 36.930 206.530 ;
        RECT 37.180 206.245 37.460 206.615 ;
        RECT 36.720 205.565 37.000 205.935 ;
        RECT 34.890 204.740 35.150 205.060 ;
        RECT 34.950 204.040 35.090 204.740 ;
        RECT 35.350 204.400 35.610 204.720 ;
        RECT 34.420 203.525 34.700 203.895 ;
        RECT 34.890 203.720 35.150 204.040 ;
        RECT 33.960 202.845 34.240 203.215 ;
        RECT 35.410 203.020 35.550 204.400 ;
        RECT 36.730 204.060 36.990 204.380 ;
        RECT 37.190 204.060 37.450 204.380 ;
        RECT 35.350 202.700 35.610 203.020 ;
        RECT 35.810 202.700 36.070 203.020 ;
        RECT 36.260 202.845 36.540 203.215 ;
        RECT 35.870 202.250 36.010 202.700 ;
        RECT 34.030 202.110 36.010 202.250 ;
        RECT 30.290 201.090 31.410 201.230 ;
        RECT 30.290 201.000 30.550 201.090 ;
        RECT 31.670 201.000 31.930 201.320 ;
        RECT 31.730 200.380 31.870 201.000 ;
        RECT 32.190 200.495 32.330 201.680 ;
        RECT 33.500 201.485 33.780 201.855 ;
        RECT 34.030 201.175 34.170 202.110 ;
        RECT 36.330 201.660 36.470 202.845 ;
        RECT 36.790 201.660 36.930 204.060 ;
        RECT 36.270 201.340 36.530 201.660 ;
        RECT 36.730 201.340 36.990 201.660 ;
        RECT 33.960 200.805 34.240 201.175 ;
        RECT 29.830 199.980 30.090 200.300 ;
        RECT 31.270 200.240 31.870 200.380 ;
        RECT 31.270 200.210 31.410 200.240 ;
        RECT 30.810 200.070 31.410 200.210 ;
        RECT 32.120 200.125 32.400 200.495 ;
        RECT 34.780 200.465 36.320 200.835 ;
        RECT 29.370 199.815 29.630 199.960 ;
        RECT 29.360 199.445 29.640 199.815 ;
        RECT 29.370 198.960 29.630 199.280 ;
        RECT 29.430 197.240 29.570 198.960 ;
        RECT 30.810 198.850 30.950 200.070 ;
        RECT 33.510 199.980 33.770 200.300 ;
        RECT 36.720 200.125 37.000 200.495 ;
        RECT 37.250 200.300 37.390 204.060 ;
        RECT 37.650 202.700 37.910 203.020 ;
        RECT 37.710 201.175 37.850 202.700 ;
        RECT 37.640 200.805 37.920 201.175 ;
        RECT 31.200 199.445 31.480 199.815 ;
        RECT 31.210 199.300 31.470 199.445 ;
        RECT 32.130 199.300 32.390 199.620 ;
        RECT 30.255 198.710 30.950 198.850 ;
        RECT 29.830 198.280 30.090 198.600 ;
        RECT 29.370 196.920 29.630 197.240 ;
        RECT 29.360 196.045 29.640 196.415 ;
        RECT 29.430 194.180 29.570 196.045 ;
        RECT 29.890 194.180 30.030 198.280 ;
        RECT 30.255 197.660 30.395 198.710 ;
        RECT 32.190 198.510 32.330 199.300 ;
        RECT 33.570 198.510 33.710 199.980 ;
        RECT 36.270 199.870 36.530 199.960 ;
        RECT 35.870 199.730 36.530 199.870 ;
        RECT 34.890 199.300 35.150 199.620 ;
        RECT 32.190 198.370 33.710 198.510 ;
        RECT 31.480 197.745 33.020 198.115 ;
        RECT 30.255 197.520 30.490 197.660 ;
        RECT 29.370 193.860 29.630 194.180 ;
        RECT 29.830 193.860 30.090 194.180 ;
        RECT 29.360 193.325 29.640 193.695 ;
        RECT 29.830 193.410 30.090 193.500 ;
        RECT 30.350 193.410 30.490 197.520 ;
        RECT 31.210 197.150 31.470 197.240 ;
        RECT 31.210 197.010 32.330 197.150 ;
        RECT 31.210 196.920 31.470 197.010 ;
        RECT 31.210 196.240 31.470 196.560 ;
        RECT 31.270 195.880 31.410 196.240 ;
        RECT 31.210 195.560 31.470 195.880 ;
        RECT 31.670 195.560 31.930 195.880 ;
        RECT 31.270 194.375 31.410 195.560 ;
        RECT 31.730 195.055 31.870 195.560 ;
        RECT 31.660 194.685 31.940 195.055 ;
        RECT 31.670 194.430 31.930 194.520 ;
        RECT 32.190 194.430 32.330 197.010 ;
        RECT 33.050 196.470 33.310 196.560 ;
        RECT 33.570 196.470 33.710 198.370 ;
        RECT 33.960 197.405 34.240 197.775 ;
        RECT 34.030 197.240 34.170 197.405 ;
        RECT 33.970 196.920 34.230 197.240 ;
        RECT 34.430 196.470 34.690 196.560 ;
        RECT 33.050 196.330 33.710 196.470 ;
        RECT 34.030 196.330 34.690 196.470 ;
        RECT 33.050 196.240 33.310 196.330 ;
        RECT 31.200 194.005 31.480 194.375 ;
        RECT 31.670 194.290 32.330 194.430 ;
        RECT 31.670 194.200 31.930 194.290 ;
        RECT 33.110 193.695 33.250 196.240 ;
        RECT 34.030 194.180 34.170 196.330 ;
        RECT 34.430 196.240 34.690 196.330 ;
        RECT 34.950 195.790 35.090 199.300 ;
        RECT 35.870 195.880 36.010 199.730 ;
        RECT 36.270 199.640 36.530 199.730 ;
        RECT 36.790 199.620 36.930 200.125 ;
        RECT 37.190 199.980 37.450 200.300 ;
        RECT 36.730 199.300 36.990 199.620 ;
        RECT 36.270 198.280 36.530 198.600 ;
        RECT 34.490 195.650 35.090 195.790 ;
        RECT 33.510 193.860 33.770 194.180 ;
        RECT 33.970 193.860 34.230 194.180 ;
        RECT 29.430 191.460 29.570 193.325 ;
        RECT 29.830 193.270 30.490 193.410 ;
        RECT 33.040 193.325 33.320 193.695 ;
        RECT 29.830 193.180 30.090 193.270 ;
        RECT 29.370 191.140 29.630 191.460 ;
        RECT 29.890 189.615 30.030 193.180 ;
        RECT 30.740 192.645 31.020 193.015 ;
        RECT 30.280 191.965 30.560 192.335 ;
        RECT 29.820 189.245 30.100 189.615 ;
        RECT 30.350 188.990 30.490 191.965 ;
        RECT 29.430 188.850 30.490 188.990 ;
        RECT 28.910 186.040 29.170 186.360 ;
        RECT 27.990 183.660 28.250 183.805 ;
        RECT 28.450 183.660 28.710 183.980 ;
        RECT 28.510 180.580 28.650 183.660 ;
        RECT 29.430 183.640 29.570 188.850 ;
        RECT 29.820 187.885 30.100 188.255 ;
        RECT 30.290 188.080 30.550 188.400 ;
        RECT 29.890 187.720 30.030 187.885 ;
        RECT 29.830 187.400 30.090 187.720 ;
        RECT 29.820 186.525 30.100 186.895 ;
        RECT 29.830 186.380 30.090 186.525 ;
        RECT 29.830 185.590 30.090 185.680 ;
        RECT 30.350 185.590 30.490 188.080 ;
        RECT 29.830 185.450 30.490 185.590 ;
        RECT 29.830 185.360 30.090 185.450 ;
        RECT 30.290 184.680 30.550 185.000 ;
        RECT 30.350 184.175 30.490 184.680 ;
        RECT 30.280 183.805 30.560 184.175 ;
        RECT 29.370 183.320 29.630 183.640 ;
        RECT 30.810 183.300 30.950 192.645 ;
        RECT 31.480 192.305 33.020 192.675 ;
        RECT 31.210 191.140 31.470 191.460 ;
        RECT 32.590 191.140 32.850 191.460 ;
        RECT 31.270 188.740 31.410 191.140 ;
        RECT 31.660 190.605 31.940 190.975 ;
        RECT 31.210 188.420 31.470 188.740 ;
        RECT 31.730 187.720 31.870 190.605 ;
        RECT 32.130 190.295 32.390 190.440 ;
        RECT 32.120 189.925 32.400 190.295 ;
        RECT 32.650 188.740 32.790 191.140 ;
        RECT 33.570 190.440 33.710 193.860 ;
        RECT 33.970 193.180 34.230 193.500 ;
        RECT 34.030 191.460 34.170 193.180 ;
        RECT 33.970 191.140 34.230 191.460 ;
        RECT 33.050 190.120 33.310 190.440 ;
        RECT 33.510 190.120 33.770 190.440 ;
        RECT 33.110 189.615 33.250 190.120 ;
        RECT 33.040 189.245 33.320 189.615 ;
        RECT 32.590 188.420 32.850 188.740 ;
        RECT 31.670 187.400 31.930 187.720 ;
        RECT 33.570 187.630 33.710 190.120 ;
        RECT 33.960 189.245 34.240 189.615 ;
        RECT 34.490 189.330 34.630 195.650 ;
        RECT 35.810 195.560 36.070 195.880 ;
        RECT 36.330 195.790 36.470 198.280 ;
        RECT 36.790 197.240 36.930 199.300 ;
        RECT 37.250 197.775 37.390 199.980 ;
        RECT 37.650 198.620 37.910 198.940 ;
        RECT 37.180 197.405 37.460 197.775 ;
        RECT 36.730 196.920 36.990 197.240 ;
        RECT 37.710 196.560 37.850 198.620 ;
        RECT 36.730 196.300 36.990 196.560 ;
        RECT 37.650 196.415 37.910 196.560 ;
        RECT 36.730 196.240 37.390 196.300 ;
        RECT 36.790 196.160 37.390 196.240 ;
        RECT 36.330 195.650 36.930 195.790 ;
        RECT 34.780 195.025 36.320 195.395 ;
        RECT 34.890 194.540 35.150 194.860 ;
        RECT 34.950 193.500 35.090 194.540 ;
        RECT 35.350 193.860 35.610 194.180 ;
        RECT 34.890 193.180 35.150 193.500 ;
        RECT 35.410 193.015 35.550 193.860 ;
        RECT 35.810 193.520 36.070 193.840 ;
        RECT 35.340 192.645 35.620 193.015 ;
        RECT 35.340 191.965 35.620 192.335 ;
        RECT 35.410 191.800 35.550 191.965 ;
        RECT 34.880 191.285 35.160 191.655 ;
        RECT 35.350 191.480 35.610 191.800 ;
        RECT 34.950 191.120 35.090 191.285 ;
        RECT 34.890 190.800 35.150 191.120 ;
        RECT 35.870 190.975 36.010 193.520 ;
        RECT 36.270 192.840 36.530 193.160 ;
        RECT 36.330 191.030 36.470 192.840 ;
        RECT 36.790 191.800 36.930 195.650 ;
        RECT 37.250 193.840 37.390 196.160 ;
        RECT 37.640 196.045 37.920 196.415 ;
        RECT 37.650 195.560 37.910 195.880 ;
        RECT 37.710 194.520 37.850 195.560 ;
        RECT 37.650 194.200 37.910 194.520 ;
        RECT 37.190 193.695 37.450 193.840 ;
        RECT 37.180 193.325 37.460 193.695 ;
        RECT 36.730 191.480 36.990 191.800 ;
        RECT 37.190 191.480 37.450 191.800 ;
        RECT 35.800 190.605 36.080 190.975 ;
        RECT 36.330 190.890 36.930 191.030 ;
        RECT 34.780 189.585 36.320 189.955 ;
        RECT 34.030 188.140 34.170 189.245 ;
        RECT 34.490 189.190 35.090 189.330 ;
        RECT 34.030 188.000 34.630 188.140 ;
        RECT 33.570 187.490 34.170 187.630 ;
        RECT 31.480 186.865 33.020 187.235 ;
        RECT 31.210 186.380 31.470 186.700 ;
        RECT 33.050 186.380 33.310 186.700 ;
        RECT 31.270 186.215 31.410 186.380 ;
        RECT 31.200 185.845 31.480 186.215 ;
        RECT 32.120 185.845 32.400 186.215 ;
        RECT 32.190 185.680 32.330 185.845 ;
        RECT 31.660 185.165 31.940 185.535 ;
        RECT 32.130 185.360 32.390 185.680 ;
        RECT 31.730 183.640 31.870 185.165 ;
        RECT 33.110 183.980 33.250 186.380 ;
        RECT 33.510 185.020 33.770 185.340 ;
        RECT 33.570 184.855 33.710 185.020 ;
        RECT 33.500 184.485 33.780 184.855 ;
        RECT 33.050 183.660 33.310 183.980 ;
        RECT 31.670 183.320 31.930 183.640 ;
        RECT 30.750 182.980 31.010 183.300 ;
        RECT 29.820 182.530 30.100 182.815 ;
        RECT 30.290 182.530 30.550 182.620 ;
        RECT 29.820 182.445 30.550 182.530 ;
        RECT 30.740 182.445 31.020 182.815 ;
        RECT 29.890 182.390 30.550 182.445 ;
        RECT 28.450 180.260 28.710 180.580 ;
        RECT 29.370 174.480 29.630 174.800 ;
        RECT 28.450 173.800 28.710 174.120 ;
        RECT 27.590 173.040 28.190 173.180 ;
        RECT 28.510 173.100 28.650 173.800 ;
        RECT 29.430 173.100 29.570 174.480 ;
        RECT 26.610 172.100 26.870 172.420 ;
        RECT 27.070 172.330 27.330 172.420 ;
        RECT 27.070 172.190 27.730 172.330 ;
        RECT 27.070 172.100 27.330 172.190 ;
        RECT 27.590 169.360 27.730 172.190 ;
        RECT 27.070 169.040 27.330 169.360 ;
        RECT 27.530 169.040 27.790 169.360 ;
        RECT 26.210 167.600 26.810 167.740 ;
        RECT 27.130 167.660 27.270 169.040 ;
        RECT 25.690 166.660 25.950 166.980 ;
        RECT 26.150 166.660 26.410 166.980 ;
        RECT 25.750 164.940 25.890 166.660 ;
        RECT 25.690 164.620 25.950 164.940 ;
        RECT 26.210 163.240 26.350 166.660 ;
        RECT 26.150 162.920 26.410 163.240 ;
        RECT 24.310 159.180 24.570 159.500 ;
        RECT 24.370 158.140 24.510 159.180 ;
        RECT 25.230 158.840 25.490 159.160 ;
        RECT 25.290 158.480 25.430 158.840 ;
        RECT 25.230 158.160 25.490 158.480 ;
        RECT 24.310 157.820 24.570 158.140 ;
        RECT 23.390 156.460 23.650 156.780 ;
        RECT 23.450 154.060 23.590 156.460 ;
        RECT 24.370 155.420 24.510 157.820 ;
        RECT 25.290 155.760 25.430 158.160 ;
        RECT 24.770 155.440 25.030 155.760 ;
        RECT 25.230 155.440 25.490 155.760 ;
        RECT 24.310 155.100 24.570 155.420 ;
        RECT 22.930 153.740 23.190 154.060 ;
        RECT 23.390 153.740 23.650 154.060 ;
        RECT 19.250 152.380 19.510 152.700 ;
        RECT 19.310 150.660 19.450 152.380 ;
        RECT 19.250 150.340 19.510 150.660 ;
        RECT 22.990 150.320 23.130 153.740 ;
        RECT 23.450 153.040 23.590 153.740 ;
        RECT 24.370 153.720 24.510 155.100 ;
        RECT 24.830 153.720 24.970 155.440 ;
        RECT 24.310 153.400 24.570 153.720 ;
        RECT 24.770 153.400 25.030 153.720 ;
        RECT 23.390 152.720 23.650 153.040 ;
        RECT 25.290 152.700 25.430 155.440 ;
        RECT 25.230 152.380 25.490 152.700 ;
        RECT 17.860 149.805 18.140 150.175 ;
        RECT 22.930 150.000 23.190 150.320 ;
        RECT 17.870 149.660 18.130 149.805 ;
        RECT 26.670 145.220 26.810 167.600 ;
        RECT 27.070 167.340 27.330 167.660 ;
        RECT 28.050 165.960 28.190 173.040 ;
        RECT 28.450 172.780 28.710 173.100 ;
        RECT 29.370 172.780 29.630 173.100 ;
        RECT 29.370 172.100 29.630 172.420 ;
        RECT 29.430 170.040 29.570 172.100 ;
        RECT 28.910 169.895 29.170 170.040 ;
        RECT 28.900 169.525 29.180 169.895 ;
        RECT 29.370 169.720 29.630 170.040 ;
        RECT 29.430 169.360 29.570 169.720 ;
        RECT 29.370 169.040 29.630 169.360 ;
        RECT 27.990 165.640 28.250 165.960 ;
        RECT 29.890 164.170 30.030 182.390 ;
        RECT 30.290 182.300 30.550 182.390 ;
        RECT 30.810 181.260 30.950 182.445 ;
        RECT 31.480 181.425 33.020 181.795 ;
        RECT 30.750 180.940 31.010 181.260 ;
        RECT 31.210 179.920 31.470 180.240 ;
        RECT 31.670 179.920 31.930 180.240 ;
        RECT 32.130 179.920 32.390 180.240 ;
        RECT 31.270 178.540 31.410 179.920 ;
        RECT 31.210 178.220 31.470 178.540 ;
        RECT 31.730 177.520 31.870 179.920 ;
        RECT 32.190 177.860 32.330 179.920 ;
        RECT 33.050 179.580 33.310 179.900 ;
        RECT 32.130 177.540 32.390 177.860 ;
        RECT 31.670 177.200 31.930 177.520 ;
        RECT 33.110 177.430 33.250 179.580 ;
        RECT 33.570 178.200 33.710 184.485 ;
        RECT 34.030 183.980 34.170 187.490 ;
        RECT 34.490 185.000 34.630 188.000 ;
        RECT 34.950 185.000 35.090 189.190 ;
        RECT 35.810 189.100 36.070 189.420 ;
        RECT 35.350 188.420 35.610 188.740 ;
        RECT 35.410 186.700 35.550 188.420 ;
        RECT 35.870 186.700 36.010 189.100 ;
        RECT 35.350 186.380 35.610 186.700 ;
        RECT 35.810 186.380 36.070 186.700 ;
        RECT 35.800 185.845 36.080 186.215 ;
        RECT 35.870 185.680 36.010 185.845 ;
        RECT 35.810 185.360 36.070 185.680 ;
        RECT 34.430 184.680 34.690 185.000 ;
        RECT 34.890 184.680 35.150 185.000 ;
        RECT 33.970 183.660 34.230 183.980 ;
        RECT 33.970 182.640 34.230 182.960 ;
        RECT 33.510 177.880 33.770 178.200 ;
        RECT 34.030 177.520 34.170 182.640 ;
        RECT 34.490 180.920 34.630 184.680 ;
        RECT 34.780 184.145 36.320 184.515 ;
        RECT 34.890 183.660 35.150 183.980 ;
        RECT 36.790 183.890 36.930 190.890 ;
        RECT 37.250 188.060 37.390 191.480 ;
        RECT 37.710 191.120 37.850 194.200 ;
        RECT 37.650 190.800 37.910 191.120 ;
        RECT 37.640 188.565 37.920 188.935 ;
        RECT 37.190 187.740 37.450 188.060 ;
        RECT 37.250 186.020 37.390 187.740 ;
        RECT 37.190 185.700 37.450 186.020 ;
        RECT 37.710 185.420 37.850 188.565 ;
        RECT 38.170 186.700 38.310 219.280 ;
        RECT 39.480 219.000 39.760 223.000 ;
        RECT 42.700 219.000 42.980 223.000 ;
        RECT 45.920 219.000 46.200 223.000 ;
        RECT 49.140 219.000 49.420 223.000 ;
        RECT 52.360 219.000 52.640 223.000 ;
        RECT 55.580 219.000 55.860 223.000 ;
        RECT 58.800 219.000 59.080 223.000 ;
        RECT 62.020 219.000 62.300 223.000 ;
        RECT 65.240 219.000 65.520 223.000 ;
        RECT 68.460 219.000 68.740 223.000 ;
        RECT 68.990 219.280 70.510 219.420 ;
        RECT 39.550 215.940 39.690 219.000 ;
        RECT 39.490 215.620 39.750 215.940 ;
        RECT 39.950 212.900 40.210 213.220 ;
        RECT 39.490 211.880 39.750 212.200 ;
        RECT 39.550 210.500 39.690 211.880 ;
        RECT 39.490 210.180 39.750 210.500 ;
        RECT 39.030 209.840 39.290 210.160 ;
        RECT 38.570 209.160 38.830 209.480 ;
        RECT 38.630 200.300 38.770 209.160 ;
        RECT 39.090 204.040 39.230 209.840 ;
        RECT 39.490 206.780 39.750 207.100 ;
        RECT 39.030 203.720 39.290 204.040 ;
        RECT 39.550 203.100 39.690 206.780 ;
        RECT 39.090 202.960 39.690 203.100 ;
        RECT 39.090 200.300 39.230 202.960 ;
        RECT 39.490 201.000 39.750 201.320 ;
        RECT 38.570 199.980 38.830 200.300 ;
        RECT 39.030 199.980 39.290 200.300 ;
        RECT 39.550 199.620 39.690 201.000 ;
        RECT 39.030 199.300 39.290 199.620 ;
        RECT 39.490 199.300 39.750 199.620 ;
        RECT 38.570 198.960 38.830 199.280 ;
        RECT 38.630 197.775 38.770 198.960 ;
        RECT 38.560 197.405 38.840 197.775 ;
        RECT 38.570 195.900 38.830 196.220 ;
        RECT 38.110 186.380 38.370 186.700 ;
        RECT 35.870 183.750 36.930 183.890 ;
        RECT 37.250 185.280 37.850 185.420 ;
        RECT 34.430 180.600 34.690 180.920 ;
        RECT 34.950 180.150 35.090 183.660 ;
        RECT 35.340 181.085 35.620 181.455 ;
        RECT 35.410 180.240 35.550 181.085 ;
        RECT 35.870 180.240 36.010 183.750 ;
        RECT 36.720 181.085 37.000 181.455 ;
        RECT 36.790 180.240 36.930 181.085 ;
        RECT 34.490 180.010 35.090 180.150 ;
        RECT 33.110 177.290 33.710 177.430 ;
        RECT 31.480 175.985 33.020 176.355 ;
        RECT 32.130 175.160 32.390 175.480 ;
        RECT 30.280 172.420 30.560 172.615 ;
        RECT 32.190 172.420 32.330 175.160 ;
        RECT 30.195 172.245 30.560 172.420 ;
        RECT 30.195 172.190 30.490 172.245 ;
        RECT 30.195 172.100 30.455 172.190 ;
        RECT 32.130 172.100 32.390 172.420 ;
        RECT 32.190 171.400 32.330 172.100 ;
        RECT 32.130 171.080 32.390 171.400 ;
        RECT 31.480 170.545 33.020 170.915 ;
        RECT 33.570 170.380 33.710 177.290 ;
        RECT 33.970 177.200 34.230 177.520 ;
        RECT 34.030 174.800 34.170 177.200 ;
        RECT 33.970 174.480 34.230 174.800 ;
        RECT 31.210 170.060 31.470 170.380 ;
        RECT 33.510 170.060 33.770 170.380 ;
        RECT 31.270 169.360 31.410 170.060 ;
        RECT 31.210 169.040 31.470 169.360 ;
        RECT 33.510 169.040 33.770 169.360 ;
        RECT 30.750 168.700 31.010 169.020 ;
        RECT 30.280 166.805 30.560 167.175 ;
        RECT 28.970 164.030 30.030 164.170 ;
        RECT 28.450 163.600 28.710 163.920 ;
        RECT 28.510 161.880 28.650 163.600 ;
        RECT 28.450 161.560 28.710 161.880 ;
        RECT 27.070 159.180 27.330 159.500 ;
        RECT 27.130 156.440 27.270 159.180 ;
        RECT 28.970 157.800 29.110 164.030 ;
        RECT 29.830 163.260 30.090 163.580 ;
        RECT 29.890 161.540 30.030 163.260 ;
        RECT 29.370 161.220 29.630 161.540 ;
        RECT 29.830 161.220 30.090 161.540 ;
        RECT 28.910 157.480 29.170 157.800 ;
        RECT 27.070 156.120 27.330 156.440 ;
        RECT 27.530 156.120 27.790 156.440 ;
        RECT 27.070 155.100 27.330 155.420 ;
        RECT 27.130 152.700 27.270 155.100 ;
        RECT 27.070 152.380 27.330 152.700 ;
        RECT 27.590 152.360 27.730 156.120 ;
        RECT 29.430 155.760 29.570 161.220 ;
        RECT 29.890 159.500 30.030 161.220 ;
        RECT 29.830 159.180 30.090 159.500 ;
        RECT 29.370 155.440 29.630 155.760 ;
        RECT 29.830 155.440 30.090 155.760 ;
        RECT 29.890 152.700 30.030 155.440 ;
        RECT 30.350 154.060 30.490 166.805 ;
        RECT 30.810 166.640 30.950 168.700 ;
        RECT 31.270 167.660 31.410 169.040 ;
        RECT 31.210 167.340 31.470 167.660 ;
        RECT 30.750 166.320 31.010 166.640 ;
        RECT 31.480 165.105 33.020 165.475 ;
        RECT 33.570 164.940 33.710 169.040 ;
        RECT 33.510 164.620 33.770 164.940 ;
        RECT 32.590 163.600 32.850 163.920 ;
        RECT 33.510 163.830 33.770 163.920 ;
        RECT 34.030 163.830 34.170 174.480 ;
        RECT 33.510 163.690 34.170 163.830 ;
        RECT 33.510 163.600 33.770 163.690 ;
        RECT 32.650 162.220 32.790 163.600 ;
        RECT 32.590 161.900 32.850 162.220 ;
        RECT 31.480 159.665 33.020 160.035 ;
        RECT 31.480 154.225 33.020 154.595 ;
        RECT 30.290 153.740 30.550 154.060 ;
        RECT 33.570 153.970 33.710 163.600 ;
        RECT 33.970 162.920 34.230 163.240 ;
        RECT 34.030 161.540 34.170 162.920 ;
        RECT 33.970 161.220 34.230 161.540 ;
        RECT 34.490 159.160 34.630 180.010 ;
        RECT 35.350 179.920 35.610 180.240 ;
        RECT 35.810 179.920 36.070 180.240 ;
        RECT 36.730 179.920 36.990 180.240 ;
        RECT 36.730 179.240 36.990 179.560 ;
        RECT 34.780 178.705 36.320 179.075 ;
        RECT 36.790 178.735 36.930 179.240 ;
        RECT 36.720 178.365 37.000 178.735 ;
        RECT 36.790 176.840 36.930 178.365 ;
        RECT 36.730 176.520 36.990 176.840 ;
        RECT 37.250 175.480 37.390 185.280 ;
        RECT 37.650 184.680 37.910 185.000 ;
        RECT 37.710 179.560 37.850 184.680 ;
        RECT 38.630 183.300 38.770 195.900 ;
        RECT 39.090 195.880 39.230 199.300 ;
        RECT 39.480 198.765 39.760 199.135 ;
        RECT 39.550 196.900 39.690 198.765 ;
        RECT 39.490 196.580 39.750 196.900 ;
        RECT 39.030 195.560 39.290 195.880 ;
        RECT 40.010 194.090 40.150 212.900 ;
        RECT 40.410 210.180 40.670 210.500 ;
        RECT 40.470 208.120 40.610 210.180 ;
        RECT 41.780 209.645 42.060 210.015 ;
        RECT 40.860 208.965 41.140 209.335 ;
        RECT 40.410 207.800 40.670 208.120 ;
        RECT 40.410 204.575 40.670 204.720 ;
        RECT 40.400 204.205 40.680 204.575 ;
        RECT 40.400 203.100 40.680 203.215 ;
        RECT 40.930 203.100 41.070 208.965 ;
        RECT 41.330 207.120 41.590 207.440 ;
        RECT 40.400 202.960 41.070 203.100 ;
        RECT 40.400 202.845 40.680 202.960 ;
        RECT 40.470 199.280 40.610 202.845 ;
        RECT 40.410 198.960 40.670 199.280 ;
        RECT 40.870 199.135 41.130 199.280 ;
        RECT 40.860 198.765 41.140 199.135 ;
        RECT 40.410 198.280 40.670 198.600 ;
        RECT 41.390 198.510 41.530 207.120 ;
        RECT 41.850 199.620 41.990 209.645 ;
        RECT 42.250 206.440 42.510 206.760 ;
        RECT 42.310 199.620 42.450 206.440 ;
        RECT 41.790 199.300 42.050 199.620 ;
        RECT 42.250 199.300 42.510 199.620 ;
        RECT 40.930 198.370 41.530 198.510 ;
        RECT 39.090 193.950 40.150 194.090 ;
        RECT 39.090 186.895 39.230 193.950 ;
        RECT 39.490 193.410 39.750 193.500 ;
        RECT 39.490 193.270 40.150 193.410 ;
        RECT 39.490 193.180 39.750 193.270 ;
        RECT 39.490 191.820 39.750 192.140 ;
        RECT 39.550 187.720 39.690 191.820 ;
        RECT 40.010 189.330 40.150 193.270 ;
        RECT 40.470 192.140 40.610 198.280 ;
        RECT 40.930 195.735 41.070 198.370 ;
        RECT 41.330 196.240 41.590 196.560 ;
        RECT 41.850 196.415 41.990 199.300 ;
        RECT 42.240 198.765 42.520 199.135 ;
        RECT 42.310 197.580 42.450 198.765 ;
        RECT 42.250 197.260 42.510 197.580 ;
        RECT 42.250 196.580 42.510 196.900 ;
        RECT 40.860 195.365 41.140 195.735 ;
        RECT 40.870 193.860 41.130 194.180 ;
        RECT 40.410 191.820 40.670 192.140 ;
        RECT 40.930 189.615 41.070 193.860 ;
        RECT 41.390 192.140 41.530 196.240 ;
        RECT 41.780 196.045 42.060 196.415 ;
        RECT 42.310 195.880 42.450 196.580 ;
        RECT 41.790 195.560 42.050 195.880 ;
        RECT 42.250 195.560 42.510 195.880 ;
        RECT 41.850 193.160 41.990 195.560 ;
        RECT 42.250 193.520 42.510 193.840 ;
        RECT 41.790 192.840 42.050 193.160 ;
        RECT 41.330 191.820 41.590 192.140 ;
        RECT 41.330 190.800 41.590 191.120 ;
        RECT 40.010 189.190 40.610 189.330 ;
        RECT 40.860 189.245 41.140 189.615 ;
        RECT 41.390 189.420 41.530 190.800 ;
        RECT 41.780 189.925 42.060 190.295 ;
        RECT 41.850 189.420 41.990 189.925 ;
        RECT 39.950 188.420 40.210 188.740 ;
        RECT 40.010 188.255 40.150 188.420 ;
        RECT 39.940 187.885 40.220 188.255 ;
        RECT 39.490 187.400 39.750 187.720 ;
        RECT 39.020 186.525 39.300 186.895 ;
        RECT 39.030 185.360 39.290 185.680 ;
        RECT 39.490 185.360 39.750 185.680 ;
        RECT 39.090 183.980 39.230 185.360 ;
        RECT 39.030 183.660 39.290 183.980 ;
        RECT 38.570 182.980 38.830 183.300 ;
        RECT 38.630 180.660 38.770 182.980 ;
        RECT 39.020 181.085 39.300 181.455 ;
        RECT 38.170 180.520 38.770 180.660 ;
        RECT 38.170 180.240 38.310 180.520 ;
        RECT 38.110 179.920 38.370 180.240 ;
        RECT 38.570 179.920 38.830 180.240 ;
        RECT 37.650 179.470 37.910 179.560 ;
        RECT 37.650 179.330 38.310 179.470 ;
        RECT 37.650 179.240 37.910 179.330 ;
        RECT 38.170 178.540 38.310 179.330 ;
        RECT 38.110 178.220 38.370 178.540 ;
        RECT 37.650 177.540 37.910 177.860 ;
        RECT 37.190 175.160 37.450 175.480 ;
        RECT 36.730 173.800 36.990 174.120 ;
        RECT 34.780 173.265 36.320 173.635 ;
        RECT 36.790 173.100 36.930 173.800 ;
        RECT 36.730 172.780 36.990 173.100 ;
        RECT 34.890 172.100 35.150 172.420 ;
        RECT 34.950 170.380 35.090 172.100 ;
        RECT 35.350 171.080 35.610 171.400 ;
        RECT 34.890 170.060 35.150 170.380 ;
        RECT 35.410 169.215 35.550 171.080 ;
        RECT 35.810 170.060 36.070 170.380 ;
        RECT 35.340 168.845 35.620 169.215 ;
        RECT 35.870 168.680 36.010 170.060 ;
        RECT 36.790 169.700 36.930 172.780 ;
        RECT 37.180 172.245 37.460 172.615 ;
        RECT 37.250 172.080 37.390 172.245 ;
        RECT 37.190 171.760 37.450 172.080 ;
        RECT 36.730 169.380 36.990 169.700 ;
        RECT 36.720 168.845 37.000 169.215 ;
        RECT 35.810 168.360 36.070 168.680 ;
        RECT 34.780 167.825 36.320 168.195 ;
        RECT 36.790 167.320 36.930 168.845 ;
        RECT 36.730 167.000 36.990 167.320 ;
        RECT 36.790 164.850 36.930 167.000 ;
        RECT 36.330 164.710 36.930 164.850 ;
        RECT 36.330 163.580 36.470 164.710 ;
        RECT 36.730 164.170 36.990 164.260 ;
        RECT 37.250 164.170 37.390 171.760 ;
        RECT 37.710 171.400 37.850 177.540 ;
        RECT 38.170 172.080 38.310 178.220 ;
        RECT 38.630 178.055 38.770 179.920 ;
        RECT 38.560 177.685 38.840 178.055 ;
        RECT 38.570 176.520 38.830 176.840 ;
        RECT 38.110 171.760 38.370 172.080 ;
        RECT 37.650 171.080 37.910 171.400 ;
        RECT 37.650 169.380 37.910 169.700 ;
        RECT 37.710 167.660 37.850 169.380 ;
        RECT 37.650 167.340 37.910 167.660 ;
        RECT 36.730 164.030 37.390 164.170 ;
        RECT 36.730 163.940 36.990 164.030 ;
        RECT 36.270 163.260 36.530 163.580 ;
        RECT 36.730 162.920 36.990 163.240 ;
        RECT 34.780 162.385 36.320 162.755 ;
        RECT 36.790 162.220 36.930 162.920 ;
        RECT 36.730 161.900 36.990 162.220 ;
        RECT 36.270 161.220 36.530 161.540 ;
        RECT 36.330 159.160 36.470 161.220 ;
        RECT 36.730 160.880 36.990 161.200 ;
        RECT 34.430 158.840 34.690 159.160 ;
        RECT 36.270 158.840 36.530 159.160 ;
        RECT 34.430 158.160 34.690 158.480 ;
        RECT 33.970 155.780 34.230 156.100 ;
        RECT 32.650 153.830 33.710 153.970 ;
        RECT 29.830 152.380 30.090 152.700 ;
        RECT 27.530 152.040 27.790 152.360 ;
        RECT 32.650 150.230 32.790 153.830 ;
        RECT 34.030 153.720 34.170 155.780 ;
        RECT 33.970 153.400 34.230 153.720 ;
        RECT 33.510 152.720 33.770 153.040 ;
        RECT 33.970 152.720 34.230 153.040 ;
        RECT 33.050 152.040 33.310 152.360 ;
        RECT 33.110 151.000 33.250 152.040 ;
        RECT 33.570 151.000 33.710 152.720 ;
        RECT 34.030 151.340 34.170 152.720 ;
        RECT 33.970 151.020 34.230 151.340 ;
        RECT 33.050 150.680 33.310 151.000 ;
        RECT 33.510 150.680 33.770 151.000 ;
        RECT 32.650 150.090 34.170 150.230 ;
        RECT 33.510 149.320 33.770 149.640 ;
        RECT 31.480 148.785 33.020 149.155 ;
        RECT 33.570 148.620 33.710 149.320 ;
        RECT 33.510 148.300 33.770 148.620 ;
        RECT 34.030 148.020 34.170 150.090 ;
        RECT 33.570 147.880 34.170 148.020 ;
        RECT 31.670 147.280 31.930 147.600 ;
        RECT 31.730 145.560 31.870 147.280 ;
        RECT 31.670 145.240 31.930 145.560 ;
        RECT 26.610 144.900 26.870 145.220 ;
        RECT 33.570 144.880 33.710 147.880 ;
        RECT 33.970 146.940 34.230 147.260 ;
        RECT 34.030 145.900 34.170 146.940 ;
        RECT 33.970 145.580 34.230 145.900 ;
        RECT 33.510 144.560 33.770 144.880 ;
        RECT 31.480 143.345 33.020 143.715 ;
        RECT 34.490 143.180 34.630 158.160 ;
        RECT 34.780 156.945 36.320 157.315 ;
        RECT 34.890 155.780 35.150 156.100 ;
        RECT 34.950 154.060 35.090 155.780 ;
        RECT 34.890 153.740 35.150 154.060 ;
        RECT 34.950 152.360 35.090 153.740 ;
        RECT 34.890 152.040 35.150 152.360 ;
        RECT 34.780 151.505 36.320 151.875 ;
        RECT 36.790 147.940 36.930 160.880 ;
        RECT 37.250 148.620 37.390 164.030 ;
        RECT 37.710 162.300 37.850 167.340 ;
        RECT 38.170 163.920 38.310 171.760 ;
        RECT 38.630 170.040 38.770 176.520 ;
        RECT 39.090 174.030 39.230 181.085 ;
        RECT 39.550 175.820 39.690 185.360 ;
        RECT 40.470 182.815 40.610 189.190 ;
        RECT 40.930 185.680 41.070 189.245 ;
        RECT 41.330 189.100 41.590 189.420 ;
        RECT 41.790 189.100 42.050 189.420 ;
        RECT 41.330 188.080 41.590 188.400 ;
        RECT 41.390 186.700 41.530 188.080 ;
        RECT 41.790 187.740 42.050 188.060 ;
        RECT 41.330 186.380 41.590 186.700 ;
        RECT 40.870 185.360 41.130 185.680 ;
        RECT 41.850 185.590 41.990 187.740 ;
        RECT 42.310 186.360 42.450 193.520 ;
        RECT 42.770 191.800 42.910 219.000 ;
        RECT 44.080 208.285 44.360 208.655 ;
        RECT 43.170 202.020 43.430 202.340 ;
        RECT 43.230 199.620 43.370 202.020 ;
        RECT 43.630 201.000 43.890 201.320 ;
        RECT 43.170 199.300 43.430 199.620 ;
        RECT 43.170 196.240 43.430 196.560 ;
        RECT 43.230 194.860 43.370 196.240 ;
        RECT 43.170 194.540 43.430 194.860 ;
        RECT 43.170 193.860 43.430 194.180 ;
        RECT 42.710 191.480 42.970 191.800 ;
        RECT 43.230 189.330 43.370 193.860 ;
        RECT 42.770 189.190 43.370 189.330 ;
        RECT 42.250 186.040 42.510 186.360 ;
        RECT 41.320 185.165 41.600 185.535 ;
        RECT 41.850 185.450 42.450 185.590 ;
        RECT 40.400 182.445 40.680 182.815 ;
        RECT 39.940 180.405 40.220 180.775 ;
        RECT 40.010 180.240 40.150 180.405 ;
        RECT 39.950 179.920 40.210 180.240 ;
        RECT 40.870 180.095 41.130 180.240 ;
        RECT 39.490 175.500 39.750 175.820 ;
        RECT 40.010 174.800 40.150 179.920 ;
        RECT 40.410 179.580 40.670 179.900 ;
        RECT 40.860 179.725 41.140 180.095 ;
        RECT 40.470 178.200 40.610 179.580 ;
        RECT 40.410 177.880 40.670 178.200 ;
        RECT 39.950 174.480 40.210 174.800 ;
        RECT 39.090 173.890 40.150 174.030 ;
        RECT 39.030 172.100 39.290 172.420 ;
        RECT 38.570 169.720 38.830 170.040 ;
        RECT 38.110 163.600 38.370 163.920 ;
        RECT 37.710 162.160 38.310 162.300 ;
        RECT 37.650 161.560 37.910 161.880 ;
        RECT 37.710 159.500 37.850 161.560 ;
        RECT 38.170 161.200 38.310 162.160 ;
        RECT 38.110 160.880 38.370 161.200 ;
        RECT 38.630 160.860 38.770 169.720 ;
        RECT 38.570 160.540 38.830 160.860 ;
        RECT 37.650 159.180 37.910 159.500 ;
        RECT 37.650 158.500 37.910 158.820 ;
        RECT 37.710 156.100 37.850 158.500 ;
        RECT 37.650 155.780 37.910 156.100 ;
        RECT 38.560 152.525 38.840 152.895 ;
        RECT 38.570 152.380 38.830 152.525 ;
        RECT 37.650 152.040 37.910 152.360 ;
        RECT 37.190 148.300 37.450 148.620 ;
        RECT 36.730 147.620 36.990 147.940 ;
        RECT 37.710 147.600 37.850 152.040 ;
        RECT 39.090 148.620 39.230 172.100 ;
        RECT 40.010 169.270 40.150 173.890 ;
        RECT 40.930 170.380 41.070 179.725 ;
        RECT 41.390 175.140 41.530 185.165 ;
        RECT 41.790 184.855 42.050 185.000 ;
        RECT 41.780 184.485 42.060 184.855 ;
        RECT 41.790 182.980 42.050 183.300 ;
        RECT 41.850 182.620 41.990 182.980 ;
        RECT 42.310 182.815 42.450 185.450 ;
        RECT 42.770 184.175 42.910 189.190 ;
        RECT 43.170 188.650 43.430 188.740 ;
        RECT 43.690 188.650 43.830 201.000 ;
        RECT 44.150 196.415 44.290 208.285 ;
        RECT 45.010 207.120 45.270 207.440 ;
        RECT 45.070 205.400 45.210 207.120 ;
        RECT 45.470 206.780 45.730 207.100 ;
        RECT 45.010 205.080 45.270 205.400 ;
        RECT 44.540 203.525 44.820 203.895 ;
        RECT 44.610 202.680 44.750 203.525 ;
        RECT 44.550 202.360 44.810 202.680 ;
        RECT 44.550 201.340 44.810 201.660 ;
        RECT 45.010 201.340 45.270 201.660 ;
        RECT 44.080 196.045 44.360 196.415 ;
        RECT 44.610 195.880 44.750 201.340 ;
        RECT 45.070 199.815 45.210 201.340 ;
        RECT 45.000 199.445 45.280 199.815 ;
        RECT 45.010 196.920 45.270 197.240 ;
        RECT 44.090 195.560 44.350 195.880 ;
        RECT 44.550 195.560 44.810 195.880 ;
        RECT 44.150 189.420 44.290 195.560 ;
        RECT 44.610 194.520 44.750 195.560 ;
        RECT 45.070 195.055 45.210 196.920 ;
        RECT 45.530 196.560 45.670 206.780 ;
        RECT 45.470 196.240 45.730 196.560 ;
        RECT 45.000 194.685 45.280 195.055 ;
        RECT 44.550 194.200 44.810 194.520 ;
        RECT 45.470 194.200 45.730 194.520 ;
        RECT 45.010 193.860 45.270 194.180 ;
        RECT 45.070 192.100 45.210 193.860 ;
        RECT 45.530 193.500 45.670 194.200 ;
        RECT 45.470 193.180 45.730 193.500 ;
        RECT 44.610 191.960 45.210 192.100 ;
        RECT 45.460 191.965 45.740 192.335 ;
        RECT 44.610 190.780 44.750 191.960 ;
        RECT 45.010 191.480 45.270 191.800 ;
        RECT 44.550 190.460 44.810 190.780 ;
        RECT 44.090 189.100 44.350 189.420 ;
        RECT 43.170 188.510 43.830 188.650 ;
        RECT 43.170 188.420 43.430 188.510 ;
        RECT 43.170 187.400 43.430 187.720 ;
        RECT 42.700 183.805 42.980 184.175 ;
        RECT 43.230 183.640 43.370 187.400 ;
        RECT 43.620 186.525 43.900 186.895 ;
        RECT 43.170 183.320 43.430 183.640 ;
        RECT 41.790 182.300 42.050 182.620 ;
        RECT 42.240 182.445 42.520 182.815 ;
        RECT 43.690 182.620 43.830 186.525 ;
        RECT 44.150 186.360 44.290 189.100 ;
        RECT 44.610 188.935 44.750 190.460 ;
        RECT 44.540 188.565 44.820 188.935 ;
        RECT 44.550 188.080 44.810 188.400 ;
        RECT 44.090 186.040 44.350 186.360 ;
        RECT 44.610 183.890 44.750 188.080 ;
        RECT 45.070 183.980 45.210 191.480 ;
        RECT 45.530 186.215 45.670 191.965 ;
        RECT 45.460 185.845 45.740 186.215 ;
        RECT 45.470 185.370 45.730 185.690 ;
        RECT 44.150 183.750 44.750 183.890 ;
        RECT 43.630 182.300 43.890 182.620 ;
        RECT 42.250 181.960 42.510 182.280 ;
        RECT 42.710 181.960 42.970 182.280 ;
        RECT 41.790 180.600 42.050 180.920 ;
        RECT 41.850 180.240 41.990 180.600 ;
        RECT 41.790 179.920 42.050 180.240 ;
        RECT 41.330 174.820 41.590 175.140 ;
        RECT 42.310 174.120 42.450 181.960 ;
        RECT 42.770 181.260 42.910 181.960 ;
        RECT 42.710 180.940 42.970 181.260 ;
        RECT 43.170 180.260 43.430 180.580 ;
        RECT 42.710 179.920 42.970 180.240 ;
        RECT 42.770 177.520 42.910 179.920 ;
        RECT 43.230 179.560 43.370 180.260 ;
        RECT 43.170 179.240 43.430 179.560 ;
        RECT 44.150 178.620 44.290 183.750 ;
        RECT 45.010 183.660 45.270 183.980 ;
        RECT 44.550 182.980 44.810 183.300 ;
        RECT 44.610 179.980 44.750 182.980 ;
        RECT 44.610 179.840 45.210 179.980 ;
        RECT 44.550 179.240 44.810 179.560 ;
        RECT 43.690 178.480 44.290 178.620 ;
        RECT 43.690 178.300 43.830 178.480 ;
        RECT 43.690 178.160 44.290 178.300 ;
        RECT 43.630 177.770 43.890 177.860 ;
        RECT 43.230 177.630 43.890 177.770 ;
        RECT 42.710 177.200 42.970 177.520 ;
        RECT 42.250 173.800 42.510 174.120 ;
        RECT 42.310 173.100 42.450 173.800 ;
        RECT 42.250 172.780 42.510 173.100 ;
        RECT 41.330 172.100 41.590 172.420 ;
        RECT 40.870 170.060 41.130 170.380 ;
        RECT 40.410 169.895 40.670 170.040 ;
        RECT 40.400 169.525 40.680 169.895 ;
        RECT 40.870 169.270 41.130 169.360 ;
        RECT 40.010 169.130 41.130 169.270 ;
        RECT 40.870 169.040 41.130 169.130 ;
        RECT 40.410 163.940 40.670 164.260 ;
        RECT 40.470 163.150 40.610 163.940 ;
        RECT 40.930 163.660 41.070 169.040 ;
        RECT 41.390 164.940 41.530 172.100 ;
        RECT 42.310 169.780 42.450 172.780 ;
        RECT 41.850 169.700 42.450 169.780 ;
        RECT 41.790 169.640 42.450 169.700 ;
        RECT 41.790 169.380 42.050 169.640 ;
        RECT 41.850 166.980 41.990 169.380 ;
        RECT 42.250 169.040 42.510 169.360 ;
        RECT 41.790 166.660 42.050 166.980 ;
        RECT 41.330 164.620 41.590 164.940 ;
        RECT 40.930 163.520 41.990 163.660 ;
        RECT 40.470 163.010 41.070 163.150 ;
        RECT 40.930 161.540 41.070 163.010 ;
        RECT 40.410 161.220 40.670 161.540 ;
        RECT 40.870 161.220 41.130 161.540 ;
        RECT 40.470 156.780 40.610 161.220 ;
        RECT 40.930 158.480 41.070 161.220 ;
        RECT 41.320 160.685 41.600 161.055 ;
        RECT 41.330 160.540 41.590 160.685 ;
        RECT 40.870 158.160 41.130 158.480 ;
        RECT 40.410 156.460 40.670 156.780 ;
        RECT 40.470 153.040 40.610 156.460 ;
        RECT 41.850 155.080 41.990 163.520 ;
        RECT 42.310 156.780 42.450 169.040 ;
        RECT 42.250 156.460 42.510 156.780 ;
        RECT 41.790 154.760 42.050 155.080 ;
        RECT 41.850 153.040 41.990 154.760 ;
        RECT 40.410 152.720 40.670 153.040 ;
        RECT 41.790 152.720 42.050 153.040 ;
        RECT 39.950 152.040 40.210 152.360 ;
        RECT 39.030 148.300 39.290 148.620 ;
        RECT 40.010 147.600 40.150 152.040 ;
        RECT 37.650 147.280 37.910 147.600 ;
        RECT 38.110 147.280 38.370 147.600 ;
        RECT 38.570 147.280 38.830 147.600 ;
        RECT 39.950 147.280 40.210 147.600 ;
        RECT 38.170 146.920 38.310 147.280 ;
        RECT 38.110 146.600 38.370 146.920 ;
        RECT 34.780 146.065 36.320 146.435 ;
        RECT 38.170 143.180 38.310 146.600 ;
        RECT 38.630 145.560 38.770 147.280 ;
        RECT 38.570 145.240 38.830 145.560 ;
        RECT 40.410 143.880 40.670 144.200 ;
        RECT 34.430 142.860 34.690 143.180 ;
        RECT 38.110 142.860 38.370 143.180 ;
        RECT 40.470 142.500 40.610 143.880 ;
        RECT 41.850 142.840 41.990 152.720 ;
        RECT 42.770 145.220 42.910 177.200 ;
        RECT 43.230 168.680 43.370 177.630 ;
        RECT 43.630 177.540 43.890 177.630 ;
        RECT 43.630 176.860 43.890 177.180 ;
        RECT 43.170 168.360 43.430 168.680 ;
        RECT 43.230 164.940 43.370 168.360 ;
        RECT 43.170 164.620 43.430 164.940 ;
        RECT 43.690 164.340 43.830 176.860 ;
        RECT 44.150 173.100 44.290 178.160 ;
        RECT 44.610 176.840 44.750 179.240 ;
        RECT 45.070 178.540 45.210 179.840 ;
        RECT 45.010 178.220 45.270 178.540 ;
        RECT 45.000 177.685 45.280 178.055 ;
        RECT 45.010 177.540 45.270 177.685 ;
        RECT 44.550 176.520 44.810 176.840 ;
        RECT 45.070 175.900 45.210 177.540 ;
        RECT 44.610 175.760 45.210 175.900 ;
        RECT 44.090 172.780 44.350 173.100 ;
        RECT 44.610 172.615 44.750 175.760 ;
        RECT 45.000 172.925 45.280 173.295 ;
        RECT 44.540 172.245 44.820 172.615 ;
        RECT 45.070 172.420 45.210 172.925 ;
        RECT 45.010 172.100 45.270 172.420 ;
        RECT 44.550 171.760 44.810 172.080 ;
        RECT 44.610 171.400 44.750 171.760 ;
        RECT 44.090 171.080 44.350 171.400 ;
        RECT 44.550 171.080 44.810 171.400 ;
        RECT 45.070 171.255 45.210 172.100 ;
        RECT 44.150 169.360 44.290 171.080 ;
        RECT 45.000 170.885 45.280 171.255 ;
        RECT 44.550 170.060 44.810 170.380 ;
        RECT 44.090 169.040 44.350 169.360 ;
        RECT 43.230 164.200 43.830 164.340 ;
        RECT 43.230 153.040 43.370 164.200 ;
        RECT 43.630 163.600 43.890 163.920 ;
        RECT 43.690 162.220 43.830 163.600 ;
        RECT 43.630 161.900 43.890 162.220 ;
        RECT 44.090 161.900 44.350 162.220 ;
        RECT 43.630 160.880 43.890 161.200 ;
        RECT 43.690 159.500 43.830 160.880 ;
        RECT 43.630 159.180 43.890 159.500 ;
        RECT 44.150 156.100 44.290 161.900 ;
        RECT 44.090 155.780 44.350 156.100 ;
        RECT 44.610 153.040 44.750 170.060 ;
        RECT 45.000 168.845 45.280 169.215 ;
        RECT 45.010 168.700 45.270 168.845 ;
        RECT 45.530 167.660 45.670 185.370 ;
        RECT 45.990 183.980 46.130 219.000 ;
        RECT 49.210 214.095 49.350 219.000 ;
        RECT 52.430 214.240 52.570 219.000 ;
        RECT 49.140 213.725 49.420 214.095 ;
        RECT 52.370 213.920 52.630 214.240 ;
        RECT 54.200 212.365 54.480 212.735 ;
        RECT 52.830 210.180 53.090 210.500 ;
        RECT 47.770 209.500 48.030 209.820 ;
        RECT 47.310 207.800 47.570 208.120 ;
        RECT 46.850 207.120 47.110 207.440 ;
        RECT 46.390 206.440 46.650 206.760 ;
        RECT 45.930 183.660 46.190 183.980 ;
        RECT 46.450 183.300 46.590 206.440 ;
        RECT 46.910 200.300 47.050 207.120 ;
        RECT 46.850 199.980 47.110 200.300 ;
        RECT 46.840 198.085 47.120 198.455 ;
        RECT 46.910 191.120 47.050 198.085 ;
        RECT 47.370 196.900 47.510 207.800 ;
        RECT 47.830 207.440 47.970 209.500 ;
        RECT 52.370 207.800 52.630 208.120 ;
        RECT 47.770 207.120 48.030 207.440 ;
        RECT 50.530 207.120 50.790 207.440 ;
        RECT 50.990 207.120 51.250 207.440 ;
        RECT 51.910 207.120 52.170 207.440 ;
        RECT 48.230 207.010 48.490 207.100 ;
        RECT 48.230 206.870 48.890 207.010 ;
        RECT 48.230 206.780 48.490 206.870 ;
        RECT 48.230 203.720 48.490 204.040 ;
        RECT 47.770 199.300 48.030 199.620 ;
        RECT 47.830 197.580 47.970 199.300 ;
        RECT 47.770 197.260 48.030 197.580 ;
        RECT 48.290 197.240 48.430 203.720 ;
        RECT 48.230 196.920 48.490 197.240 ;
        RECT 47.310 196.580 47.570 196.900 ;
        RECT 48.220 196.045 48.500 196.415 ;
        RECT 47.770 195.560 48.030 195.880 ;
        RECT 47.300 194.005 47.580 194.375 ;
        RECT 47.830 194.180 47.970 195.560 ;
        RECT 48.290 194.860 48.430 196.045 ;
        RECT 48.230 194.540 48.490 194.860 ;
        RECT 48.290 194.180 48.430 194.540 ;
        RECT 46.850 190.800 47.110 191.120 ;
        RECT 46.840 189.245 47.120 189.615 ;
        RECT 46.850 189.100 47.110 189.245 ;
        RECT 47.370 188.935 47.510 194.005 ;
        RECT 47.770 193.860 48.030 194.180 ;
        RECT 48.230 193.860 48.490 194.180 ;
        RECT 48.230 192.840 48.490 193.160 ;
        RECT 48.290 192.140 48.430 192.840 ;
        RECT 48.230 191.820 48.490 192.140 ;
        RECT 48.290 190.860 48.430 191.820 ;
        RECT 48.750 191.800 48.890 206.870 ;
        RECT 49.150 206.780 49.410 207.100 ;
        RECT 49.210 205.060 49.350 206.780 ;
        RECT 49.150 204.740 49.410 205.060 ;
        RECT 49.610 204.740 49.870 205.060 ;
        RECT 49.210 202.680 49.350 204.740 ;
        RECT 49.150 202.360 49.410 202.680 ;
        RECT 49.670 200.495 49.810 204.740 ;
        RECT 50.060 202.165 50.340 202.535 ;
        RECT 49.600 200.125 49.880 200.495 ;
        RECT 49.610 195.900 49.870 196.220 ;
        RECT 49.670 194.520 49.810 195.900 ;
        RECT 49.610 194.200 49.870 194.520 ;
        RECT 48.690 191.480 48.950 191.800 ;
        RECT 49.150 191.480 49.410 191.800 ;
        RECT 50.130 191.540 50.270 202.165 ;
        RECT 50.590 192.140 50.730 207.120 ;
        RECT 51.050 199.960 51.190 207.120 ;
        RECT 51.450 205.080 51.710 205.400 ;
        RECT 51.510 204.720 51.650 205.080 ;
        RECT 51.450 204.400 51.710 204.720 ;
        RECT 51.450 201.340 51.710 201.660 ;
        RECT 50.990 199.640 51.250 199.960 ;
        RECT 50.980 197.405 51.260 197.775 ;
        RECT 51.050 192.165 51.190 197.405 ;
        RECT 50.530 191.820 50.790 192.140 ;
        RECT 50.980 191.795 51.260 192.165 ;
        RECT 47.830 190.720 48.430 190.860 ;
        RECT 48.690 190.800 48.950 191.120 ;
        RECT 47.300 188.565 47.580 188.935 ;
        RECT 47.830 188.740 47.970 190.720 ;
        RECT 48.230 190.120 48.490 190.440 ;
        RECT 47.310 188.420 47.570 188.565 ;
        RECT 47.770 188.420 48.030 188.740 ;
        RECT 47.370 185.535 47.510 188.420 ;
        RECT 47.770 187.740 48.030 188.060 ;
        RECT 47.830 186.360 47.970 187.740 ;
        RECT 48.290 186.700 48.430 190.120 ;
        RECT 48.230 186.380 48.490 186.700 ;
        RECT 47.770 186.040 48.030 186.360 ;
        RECT 47.300 185.165 47.580 185.535 ;
        RECT 47.830 185.340 47.970 186.040 ;
        RECT 48.230 185.360 48.490 185.680 ;
        RECT 47.770 185.020 48.030 185.340 ;
        RECT 47.300 184.485 47.580 184.855 ;
        RECT 48.290 184.740 48.430 185.360 ;
        RECT 47.830 184.600 48.430 184.740 ;
        RECT 47.370 183.300 47.510 184.485 ;
        RECT 46.390 182.980 46.650 183.300 ;
        RECT 47.310 182.980 47.570 183.300 ;
        RECT 47.300 182.445 47.580 182.815 ;
        RECT 45.930 180.260 46.190 180.580 ;
        RECT 46.380 180.405 46.660 180.775 ;
        RECT 45.470 167.340 45.730 167.660 ;
        RECT 45.470 164.620 45.730 164.940 ;
        RECT 45.530 161.880 45.670 164.620 ;
        RECT 45.470 161.560 45.730 161.880 ;
        RECT 45.990 161.735 46.130 180.260 ;
        RECT 46.450 179.900 46.590 180.405 ;
        RECT 47.370 179.900 47.510 182.445 ;
        RECT 47.830 182.135 47.970 184.600 ;
        RECT 47.760 181.765 48.040 182.135 ;
        RECT 48.230 181.960 48.490 182.280 ;
        RECT 47.760 181.085 48.040 181.455 ;
        RECT 47.770 180.940 48.030 181.085 ;
        RECT 47.770 179.920 48.030 180.240 ;
        RECT 46.390 179.580 46.650 179.900 ;
        RECT 47.310 179.580 47.570 179.900 ;
        RECT 46.840 179.045 47.120 179.415 ;
        RECT 46.380 178.365 46.660 178.735 ;
        RECT 46.390 178.220 46.650 178.365 ;
        RECT 46.910 177.980 47.050 179.045 ;
        RECT 46.850 177.660 47.110 177.980 ;
        RECT 47.310 176.860 47.570 177.180 ;
        RECT 47.370 175.335 47.510 176.860 ;
        RECT 47.300 174.965 47.580 175.335 ;
        RECT 46.380 173.605 46.660 173.975 ;
        RECT 46.450 168.420 46.590 173.605 ;
        RECT 46.850 172.100 47.110 172.420 ;
        RECT 46.910 170.380 47.050 172.100 ;
        RECT 46.850 170.060 47.110 170.380 ;
        RECT 46.450 168.280 47.050 168.420 ;
        RECT 46.390 167.340 46.650 167.660 ;
        RECT 45.010 161.220 45.270 161.540 ;
        RECT 45.070 159.695 45.210 161.220 ;
        RECT 45.530 160.520 45.670 161.560 ;
        RECT 45.920 161.365 46.200 161.735 ;
        RECT 45.930 161.220 46.190 161.365 ;
        RECT 45.920 160.685 46.200 161.055 ;
        RECT 45.930 160.540 46.190 160.685 ;
        RECT 45.470 160.200 45.730 160.520 ;
        RECT 45.000 159.325 45.280 159.695 ;
        RECT 45.930 158.840 46.190 159.160 ;
        RECT 45.470 157.480 45.730 157.800 ;
        RECT 45.530 156.440 45.670 157.480 ;
        RECT 45.990 156.440 46.130 158.840 ;
        RECT 45.470 156.120 45.730 156.440 ;
        RECT 45.930 156.120 46.190 156.440 ;
        RECT 45.010 155.780 45.270 156.100 ;
        RECT 45.070 154.060 45.210 155.780 ;
        RECT 46.450 154.060 46.590 167.340 ;
        RECT 46.910 164.260 47.050 168.280 ;
        RECT 46.850 163.940 47.110 164.260 ;
        RECT 47.830 163.240 47.970 179.920 ;
        RECT 48.290 177.860 48.430 181.960 ;
        RECT 48.750 178.735 48.890 190.800 ;
        RECT 49.210 190.440 49.350 191.480 ;
        RECT 49.670 191.400 50.270 191.540 ;
        RECT 49.150 190.120 49.410 190.440 ;
        RECT 49.210 189.420 49.350 190.120 ;
        RECT 49.670 189.615 49.810 191.400 ;
        RECT 50.990 190.800 51.250 191.120 ;
        RECT 50.530 190.460 50.790 190.780 ;
        RECT 50.590 190.295 50.730 190.460 ;
        RECT 50.520 189.925 50.800 190.295 ;
        RECT 49.150 189.100 49.410 189.420 ;
        RECT 49.600 189.245 49.880 189.615 ;
        RECT 50.590 189.080 50.730 189.925 ;
        RECT 50.530 188.760 50.790 189.080 ;
        RECT 50.070 188.080 50.330 188.400 ;
        RECT 50.530 188.080 50.790 188.400 ;
        RECT 51.050 188.255 51.190 190.800 ;
        RECT 49.610 185.700 49.870 186.020 ;
        RECT 49.150 180.260 49.410 180.580 ;
        RECT 48.680 178.365 48.960 178.735 ;
        RECT 48.230 177.540 48.490 177.860 ;
        RECT 48.220 177.005 48.500 177.375 ;
        RECT 48.230 176.860 48.490 177.005 ;
        RECT 48.690 176.860 48.950 177.180 ;
        RECT 48.750 176.695 48.890 176.860 ;
        RECT 49.210 176.840 49.350 180.260 ;
        RECT 49.670 180.240 49.810 185.700 ;
        RECT 49.610 179.920 49.870 180.240 ;
        RECT 48.680 176.325 48.960 176.695 ;
        RECT 49.150 176.520 49.410 176.840 ;
        RECT 50.130 175.390 50.270 188.080 ;
        RECT 50.590 186.360 50.730 188.080 ;
        RECT 50.980 187.885 51.260 188.255 ;
        RECT 51.510 188.060 51.650 201.340 ;
        RECT 51.970 194.860 52.110 207.120 ;
        RECT 52.430 202.000 52.570 207.800 ;
        RECT 52.370 201.680 52.630 202.000 ;
        RECT 52.430 198.600 52.570 201.680 ;
        RECT 52.370 198.280 52.630 198.600 ;
        RECT 52.370 197.260 52.630 197.580 ;
        RECT 51.910 194.540 52.170 194.860 ;
        RECT 51.900 192.645 52.180 193.015 ;
        RECT 51.970 192.140 52.110 192.645 ;
        RECT 51.910 191.820 52.170 192.140 ;
        RECT 51.900 191.285 52.180 191.655 ;
        RECT 51.450 187.740 51.710 188.060 ;
        RECT 50.990 187.400 51.250 187.720 ;
        RECT 50.530 186.040 50.790 186.360 ;
        RECT 51.050 185.680 51.190 187.400 ;
        RECT 50.530 185.360 50.790 185.680 ;
        RECT 50.990 185.360 51.250 185.680 ;
        RECT 50.590 182.960 50.730 185.360 ;
        RECT 50.980 184.485 51.260 184.855 ;
        RECT 51.450 184.680 51.710 185.000 ;
        RECT 51.050 183.300 51.190 184.485 ;
        RECT 51.510 183.300 51.650 184.680 ;
        RECT 51.970 183.980 52.110 191.285 ;
        RECT 52.430 190.780 52.570 197.260 ;
        RECT 52.370 190.460 52.630 190.780 ;
        RECT 52.430 186.020 52.570 190.460 ;
        RECT 52.890 186.700 53.030 210.180 ;
        RECT 53.750 209.160 54.010 209.480 ;
        RECT 53.290 206.615 53.550 206.760 ;
        RECT 53.280 206.245 53.560 206.615 ;
        RECT 53.290 201.680 53.550 202.000 ;
        RECT 53.350 200.300 53.490 201.680 ;
        RECT 53.290 199.980 53.550 200.300 ;
        RECT 53.810 199.620 53.950 209.160 ;
        RECT 53.750 199.300 54.010 199.620 ;
        RECT 53.290 196.240 53.550 196.560 ;
        RECT 53.350 195.055 53.490 196.240 ;
        RECT 53.280 194.685 53.560 195.055 ;
        RECT 53.290 191.820 53.550 192.140 ;
        RECT 54.270 192.100 54.410 212.365 ;
        RECT 55.650 212.055 55.790 219.000 ;
        RECT 56.970 213.580 57.230 213.900 ;
        RECT 55.580 211.685 55.860 212.055 ;
        RECT 54.670 210.520 54.930 210.840 ;
        RECT 54.730 204.040 54.870 210.520 ;
        RECT 55.590 209.840 55.850 210.160 ;
        RECT 56.050 209.840 56.310 210.160 ;
        RECT 56.510 209.840 56.770 210.160 ;
        RECT 55.120 205.565 55.400 205.935 ;
        RECT 55.650 205.740 55.790 209.840 ;
        RECT 56.110 209.335 56.250 209.840 ;
        RECT 56.040 208.965 56.320 209.335 ;
        RECT 56.570 208.120 56.710 209.840 ;
        RECT 56.510 207.800 56.770 208.120 ;
        RECT 54.670 203.720 54.930 204.040 ;
        RECT 54.730 200.300 54.870 203.720 ;
        RECT 54.670 199.980 54.930 200.300 ;
        RECT 54.670 198.620 54.930 198.940 ;
        RECT 54.730 193.160 54.870 198.620 ;
        RECT 54.670 192.840 54.930 193.160 ;
        RECT 54.730 192.140 54.870 192.840 ;
        RECT 53.810 191.960 54.410 192.100 ;
        RECT 53.350 189.080 53.490 191.820 ;
        RECT 53.290 188.760 53.550 189.080 ;
        RECT 53.280 187.885 53.560 188.255 ;
        RECT 52.830 186.380 53.090 186.700 ;
        RECT 52.370 185.700 52.630 186.020 ;
        RECT 52.820 185.165 53.100 185.535 ;
        RECT 51.910 183.660 52.170 183.980 ;
        RECT 50.990 182.980 51.250 183.300 ;
        RECT 51.450 182.980 51.710 183.300 ;
        RECT 51.910 182.980 52.170 183.300 ;
        RECT 52.370 182.980 52.630 183.300 ;
        RECT 50.530 182.640 50.790 182.960 ;
        RECT 50.530 182.135 50.790 182.280 ;
        RECT 50.520 181.765 50.800 182.135 ;
        RECT 50.530 179.920 50.790 180.240 ;
        RECT 50.590 175.900 50.730 179.920 ;
        RECT 50.980 179.725 51.260 180.095 ;
        RECT 50.990 179.580 51.250 179.725 ;
        RECT 51.970 178.735 52.110 182.980 ;
        RECT 52.430 181.260 52.570 182.980 ;
        RECT 52.890 182.815 53.030 185.165 ;
        RECT 52.820 182.445 53.100 182.815 ;
        RECT 52.370 180.940 52.630 181.260 ;
        RECT 52.890 179.900 53.030 182.445 ;
        RECT 52.830 179.580 53.090 179.900 ;
        RECT 50.980 178.365 51.260 178.735 ;
        RECT 51.900 178.365 52.180 178.735 ;
        RECT 50.990 178.220 51.250 178.365 ;
        RECT 50.990 177.540 51.250 177.860 ;
        RECT 51.450 177.540 51.710 177.860 ;
        RECT 51.900 177.685 52.180 178.055 ;
        RECT 51.910 177.540 52.170 177.685 ;
        RECT 51.050 177.375 51.190 177.540 ;
        RECT 50.980 177.005 51.260 177.375 ;
        RECT 50.590 175.760 51.190 175.900 ;
        RECT 51.050 175.480 51.190 175.760 ;
        RECT 50.130 175.250 50.730 175.390 ;
        RECT 49.140 173.605 49.420 173.975 ;
        RECT 49.610 173.800 49.870 174.120 ;
        RECT 50.590 174.030 50.730 175.250 ;
        RECT 50.990 175.160 51.250 175.480 ;
        RECT 50.990 174.480 51.250 174.800 ;
        RECT 51.510 174.655 51.650 177.540 ;
        RECT 53.350 177.260 53.490 187.885 ;
        RECT 53.810 185.000 53.950 191.960 ;
        RECT 54.670 191.820 54.930 192.140 ;
        RECT 55.190 191.540 55.330 205.565 ;
        RECT 55.590 205.420 55.850 205.740 ;
        RECT 55.650 200.495 55.790 205.420 ;
        RECT 56.510 205.080 56.770 205.400 ;
        RECT 56.570 202.680 56.710 205.080 ;
        RECT 57.030 204.575 57.170 213.580 ;
        RECT 58.870 213.300 59.010 219.000 ;
        RECT 62.090 216.135 62.230 219.000 ;
        RECT 62.020 215.765 62.300 216.135 ;
        RECT 65.310 215.455 65.450 219.000 ;
        RECT 68.530 218.740 68.670 219.000 ;
        RECT 68.990 218.740 69.130 219.280 ;
        RECT 68.530 218.600 69.130 218.740 ;
        RECT 65.240 215.085 65.520 215.455 ;
        RECT 66.620 215.085 66.900 215.455 ;
        RECT 57.430 212.900 57.690 213.220 ;
        RECT 58.410 213.160 59.010 213.300 ;
        RECT 56.960 204.205 57.240 204.575 ;
        RECT 56.510 202.360 56.770 202.680 ;
        RECT 56.970 202.360 57.230 202.680 ;
        RECT 56.050 201.680 56.310 202.000 ;
        RECT 56.510 201.680 56.770 202.000 ;
        RECT 55.580 200.125 55.860 200.495 ;
        RECT 56.110 199.960 56.250 201.680 ;
        RECT 56.050 199.640 56.310 199.960 ;
        RECT 56.570 199.135 56.710 201.680 ;
        RECT 56.500 198.765 56.780 199.135 ;
        RECT 56.510 198.280 56.770 198.600 ;
        RECT 56.050 193.520 56.310 193.840 ;
        RECT 55.590 192.840 55.850 193.160 ;
        RECT 55.650 192.140 55.790 192.840 ;
        RECT 55.590 191.820 55.850 192.140 ;
        RECT 55.190 191.400 55.790 191.540 ;
        RECT 54.210 190.800 54.470 191.120 ;
        RECT 54.270 187.575 54.410 190.800 ;
        RECT 55.130 188.420 55.390 188.740 ;
        RECT 54.670 188.080 54.930 188.400 ;
        RECT 54.200 187.205 54.480 187.575 ;
        RECT 54.730 186.700 54.870 188.080 ;
        RECT 54.670 186.380 54.930 186.700 ;
        RECT 54.200 185.165 54.480 185.535 ;
        RECT 53.750 184.680 54.010 185.000 ;
        RECT 53.750 182.980 54.010 183.300 ;
        RECT 53.810 182.815 53.950 182.980 ;
        RECT 53.740 182.445 54.020 182.815 ;
        RECT 53.750 181.960 54.010 182.280 ;
        RECT 53.810 181.455 53.950 181.960 ;
        RECT 53.740 181.085 54.020 181.455 ;
        RECT 53.740 180.405 54.020 180.775 ;
        RECT 53.810 177.860 53.950 180.405 ;
        RECT 54.270 177.860 54.410 185.165 ;
        RECT 54.670 183.320 54.930 183.640 ;
        RECT 54.730 180.240 54.870 183.320 ;
        RECT 54.670 179.920 54.930 180.240 ;
        RECT 55.190 178.620 55.330 188.420 ;
        RECT 54.730 178.480 55.330 178.620 ;
        RECT 53.750 177.540 54.010 177.860 ;
        RECT 54.210 177.540 54.470 177.860 ;
        RECT 52.890 177.180 53.490 177.260 ;
        RECT 52.830 177.120 53.490 177.180 ;
        RECT 53.810 177.260 53.950 177.540 ;
        RECT 53.810 177.120 54.410 177.260 ;
        RECT 52.830 176.860 53.090 177.120 ;
        RECT 53.750 176.520 54.010 176.840 ;
        RECT 53.290 175.500 53.550 175.820 ;
        RECT 52.830 175.160 53.090 175.480 ;
        RECT 50.130 173.890 50.730 174.030 ;
        RECT 48.680 172.925 48.960 173.295 ;
        RECT 48.750 170.040 48.890 172.925 ;
        RECT 48.690 169.720 48.950 170.040 ;
        RECT 48.230 169.040 48.490 169.360 ;
        RECT 47.770 162.920 48.030 163.240 ;
        RECT 47.770 161.735 48.030 161.880 ;
        RECT 47.760 161.365 48.040 161.735 ;
        RECT 47.770 160.880 48.030 161.200 ;
        RECT 47.310 160.200 47.570 160.520 ;
        RECT 46.850 158.160 47.110 158.480 ;
        RECT 46.910 156.100 47.050 158.160 ;
        RECT 47.370 156.100 47.510 160.200 ;
        RECT 47.830 159.695 47.970 160.880 ;
        RECT 47.760 159.325 48.040 159.695 ;
        RECT 47.830 156.100 47.970 159.325 ;
        RECT 46.850 155.780 47.110 156.100 ;
        RECT 47.310 155.780 47.570 156.100 ;
        RECT 47.770 155.780 48.030 156.100 ;
        RECT 45.010 153.740 45.270 154.060 ;
        RECT 46.390 153.740 46.650 154.060 ;
        RECT 43.170 152.720 43.430 153.040 ;
        RECT 44.550 152.720 44.810 153.040 ;
        RECT 43.230 147.600 43.370 152.720 ;
        RECT 44.610 147.600 44.750 152.720 ;
        RECT 43.170 147.280 43.430 147.600 ;
        RECT 44.550 147.280 44.810 147.600 ;
        RECT 43.230 145.900 43.370 147.280 ;
        RECT 43.170 145.580 43.430 145.900 ;
        RECT 42.710 144.900 42.970 145.220 ;
        RECT 42.770 143.180 42.910 144.900 ;
        RECT 43.230 143.180 43.370 145.580 ;
        RECT 44.610 145.560 44.750 147.280 ;
        RECT 44.550 145.240 44.810 145.560 ;
        RECT 47.370 145.220 47.510 155.780 ;
        RECT 47.830 151.340 47.970 155.780 ;
        RECT 47.770 151.020 48.030 151.340 ;
        RECT 48.290 149.980 48.430 169.040 ;
        RECT 48.690 165.640 48.950 165.960 ;
        RECT 48.750 160.520 48.890 165.640 ;
        RECT 48.690 160.200 48.950 160.520 ;
        RECT 48.750 158.480 48.890 160.200 ;
        RECT 48.690 158.160 48.950 158.480 ;
        RECT 49.210 153.720 49.350 173.605 ;
        RECT 49.670 173.295 49.810 173.800 ;
        RECT 49.600 172.925 49.880 173.295 ;
        RECT 49.600 172.245 49.880 172.615 ;
        RECT 49.670 167.060 49.810 172.245 ;
        RECT 50.130 171.740 50.270 173.890 ;
        RECT 50.530 172.440 50.790 172.760 ;
        RECT 50.070 171.420 50.330 171.740 ;
        RECT 50.590 167.660 50.730 172.440 ;
        RECT 51.050 170.040 51.190 174.480 ;
        RECT 51.440 174.285 51.720 174.655 ;
        RECT 52.370 174.140 52.630 174.460 ;
        RECT 51.450 173.800 51.710 174.120 ;
        RECT 51.910 173.800 52.170 174.120 ;
        RECT 51.510 173.295 51.650 173.800 ;
        RECT 51.440 172.925 51.720 173.295 ;
        RECT 51.970 172.760 52.110 173.800 ;
        RECT 52.430 172.760 52.570 174.140 ;
        RECT 51.910 172.440 52.170 172.760 ;
        RECT 52.370 172.440 52.630 172.760 ;
        RECT 51.450 172.100 51.710 172.420 ;
        RECT 50.990 169.720 51.250 170.040 ;
        RECT 51.510 169.020 51.650 172.100 ;
        RECT 51.450 168.700 51.710 169.020 ;
        RECT 50.990 168.360 51.250 168.680 ;
        RECT 50.530 167.340 50.790 167.660 ;
        RECT 49.670 166.920 50.730 167.060 ;
        RECT 49.610 163.600 49.870 163.920 ;
        RECT 49.670 162.220 49.810 163.600 ;
        RECT 50.070 162.920 50.330 163.240 ;
        RECT 49.610 161.900 49.870 162.220 ;
        RECT 50.130 158.480 50.270 162.920 ;
        RECT 50.070 158.160 50.330 158.480 ;
        RECT 50.590 156.440 50.730 166.920 ;
        RECT 51.050 161.880 51.190 168.360 ;
        RECT 52.430 167.320 52.570 172.440 ;
        RECT 52.890 171.255 53.030 175.160 ;
        RECT 53.350 175.140 53.490 175.500 ;
        RECT 53.290 174.820 53.550 175.140 ;
        RECT 53.810 174.800 53.950 176.520 ;
        RECT 53.750 174.480 54.010 174.800 ;
        RECT 54.270 174.460 54.410 177.120 ;
        RECT 54.210 174.140 54.470 174.460 ;
        RECT 53.290 173.800 53.550 174.120 ;
        RECT 52.820 170.885 53.100 171.255 ;
        RECT 52.830 168.360 53.090 168.680 ;
        RECT 52.370 167.060 52.630 167.320 ;
        RECT 51.510 167.000 52.630 167.060 ;
        RECT 51.510 166.920 52.570 167.000 ;
        RECT 52.890 166.980 53.030 168.360 ;
        RECT 53.350 167.660 53.490 173.800 ;
        RECT 54.200 173.605 54.480 173.975 ;
        RECT 53.750 172.100 54.010 172.420 ;
        RECT 53.290 167.340 53.550 167.660 ;
        RECT 53.810 166.980 53.950 172.100 ;
        RECT 51.510 166.640 51.650 166.920 ;
        RECT 52.830 166.660 53.090 166.980 ;
        RECT 53.750 166.660 54.010 166.980 ;
        RECT 51.450 166.320 51.710 166.640 ;
        RECT 53.810 164.940 53.950 166.660 ;
        RECT 53.750 164.620 54.010 164.940 ;
        RECT 51.910 163.600 52.170 163.920 ;
        RECT 51.450 162.920 51.710 163.240 ;
        RECT 51.510 161.880 51.650 162.920 ;
        RECT 50.990 161.560 51.250 161.880 ;
        RECT 51.450 161.560 51.710 161.880 ;
        RECT 51.050 160.860 51.190 161.560 ;
        RECT 50.990 160.540 51.250 160.860 ;
        RECT 51.970 160.520 52.110 163.600 ;
        RECT 52.830 163.260 53.090 163.580 ;
        RECT 52.890 162.220 53.030 163.260 ;
        RECT 54.270 162.220 54.410 173.605 ;
        RECT 54.730 173.100 54.870 178.480 ;
        RECT 55.120 174.285 55.400 174.655 ;
        RECT 54.670 172.780 54.930 173.100 ;
        RECT 55.190 167.740 55.330 174.285 ;
        RECT 55.650 173.100 55.790 191.400 ;
        RECT 56.110 188.400 56.250 193.520 ;
        RECT 56.050 188.080 56.310 188.400 ;
        RECT 56.040 183.805 56.320 184.175 ;
        RECT 56.110 181.260 56.250 183.805 ;
        RECT 56.050 180.940 56.310 181.260 ;
        RECT 56.570 180.660 56.710 198.280 ;
        RECT 57.030 191.120 57.170 202.360 ;
        RECT 57.490 201.855 57.630 212.900 ;
        RECT 58.410 207.780 58.550 213.160 ;
        RECT 59.270 212.560 59.530 212.880 ;
        RECT 58.810 210.180 59.070 210.500 ;
        RECT 58.350 207.460 58.610 207.780 ;
        RECT 58.870 207.100 59.010 210.180 ;
        RECT 59.330 207.440 59.470 212.560 ;
        RECT 60.650 210.860 60.910 211.180 ;
        RECT 65.250 210.860 65.510 211.180 ;
        RECT 59.270 207.120 59.530 207.440 ;
        RECT 58.810 206.780 59.070 207.100 ;
        RECT 59.330 205.650 59.470 207.120 ;
        RECT 57.950 205.510 59.470 205.650 ;
        RECT 57.950 202.000 58.090 205.510 ;
        RECT 58.810 204.740 59.070 205.060 ;
        RECT 58.350 204.400 58.610 204.720 ;
        RECT 57.420 201.485 57.700 201.855 ;
        RECT 57.890 201.680 58.150 202.000 ;
        RECT 57.950 197.580 58.090 201.680 ;
        RECT 58.410 201.660 58.550 204.400 ;
        RECT 58.350 201.340 58.610 201.660 ;
        RECT 58.350 198.960 58.610 199.280 ;
        RECT 58.410 198.455 58.550 198.960 ;
        RECT 58.340 198.085 58.620 198.455 ;
        RECT 57.890 197.260 58.150 197.580 ;
        RECT 57.890 194.200 58.150 194.520 ;
        RECT 57.430 193.860 57.690 194.180 ;
        RECT 56.970 190.800 57.230 191.120 ;
        RECT 56.970 188.760 57.230 189.080 ;
        RECT 57.030 185.000 57.170 188.760 ;
        RECT 57.490 186.360 57.630 193.860 ;
        RECT 57.950 189.080 58.090 194.200 ;
        RECT 58.870 193.160 59.010 204.740 ;
        RECT 59.270 204.400 59.530 204.720 ;
        RECT 59.330 201.320 59.470 204.400 ;
        RECT 59.730 204.060 59.990 204.380 ;
        RECT 59.270 201.000 59.530 201.320 ;
        RECT 58.810 192.840 59.070 193.160 ;
        RECT 58.800 191.965 59.080 192.335 ;
        RECT 58.870 191.800 59.010 191.965 ;
        RECT 58.810 191.480 59.070 191.800 ;
        RECT 57.890 188.760 58.150 189.080 ;
        RECT 57.890 188.080 58.150 188.400 ;
        RECT 57.430 186.040 57.690 186.360 ;
        RECT 56.970 184.680 57.230 185.000 ;
        RECT 57.950 183.980 58.090 188.080 ;
        RECT 58.870 185.680 59.010 191.480 ;
        RECT 59.330 191.120 59.470 201.000 ;
        RECT 59.790 199.620 59.930 204.060 ;
        RECT 60.190 201.000 60.450 201.320 ;
        RECT 59.730 199.300 59.990 199.620 ;
        RECT 60.250 199.280 60.390 201.000 ;
        RECT 60.710 199.620 60.850 210.860 ;
        RECT 63.870 210.520 64.130 210.840 ;
        RECT 61.570 206.780 61.830 207.100 ;
        RECT 61.110 201.680 61.370 202.000 ;
        RECT 60.650 199.300 60.910 199.620 ;
        RECT 60.190 198.960 60.450 199.280 ;
        RECT 60.650 198.620 60.910 198.940 ;
        RECT 60.710 196.900 60.850 198.620 ;
        RECT 60.650 196.580 60.910 196.900 ;
        RECT 59.730 196.240 59.990 196.560 ;
        RECT 59.790 193.160 59.930 196.240 ;
        RECT 59.730 192.840 59.990 193.160 ;
        RECT 61.170 193.015 61.310 201.680 ;
        RECT 61.630 201.320 61.770 206.780 ;
        RECT 62.950 204.740 63.210 205.060 ;
        RECT 62.030 204.400 62.290 204.720 ;
        RECT 61.570 201.000 61.830 201.320 ;
        RECT 61.630 199.620 61.770 201.000 ;
        RECT 61.570 199.300 61.830 199.620 ;
        RECT 61.570 198.620 61.830 198.940 ;
        RECT 61.100 192.645 61.380 193.015 ;
        RECT 59.720 191.965 60.000 192.335 ;
        RECT 59.790 191.120 59.930 191.965 ;
        RECT 61.630 191.540 61.770 198.620 ;
        RECT 62.090 198.340 62.230 204.400 ;
        RECT 62.090 198.200 62.690 198.340 ;
        RECT 62.030 195.560 62.290 195.880 ;
        RECT 61.170 191.400 61.770 191.540 ;
        RECT 59.270 190.800 59.530 191.120 ;
        RECT 59.730 190.800 59.990 191.120 ;
        RECT 59.330 187.720 59.470 190.800 ;
        RECT 59.270 187.400 59.530 187.720 ;
        RECT 59.260 186.525 59.540 186.895 ;
        RECT 58.810 185.360 59.070 185.680 ;
        RECT 59.330 183.980 59.470 186.525 ;
        RECT 57.890 183.660 58.150 183.980 ;
        RECT 58.810 183.660 59.070 183.980 ;
        RECT 59.270 183.660 59.530 183.980 ;
        RECT 57.430 182.640 57.690 182.960 ;
        RECT 57.490 180.920 57.630 182.640 ;
        RECT 58.870 182.280 59.010 183.660 ;
        RECT 59.260 183.125 59.540 183.495 ;
        RECT 59.270 182.980 59.530 183.125 ;
        RECT 59.790 182.960 59.930 190.800 ;
        RECT 61.170 188.935 61.310 191.400 ;
        RECT 62.090 191.120 62.230 195.560 ;
        RECT 61.570 190.800 61.830 191.120 ;
        RECT 62.030 190.800 62.290 191.120 ;
        RECT 61.100 188.565 61.380 188.935 ;
        RECT 60.180 187.205 60.460 187.575 ;
        RECT 60.650 187.400 60.910 187.720 ;
        RECT 60.250 183.980 60.390 187.205 ;
        RECT 60.190 183.660 60.450 183.980 ;
        RECT 59.730 182.640 59.990 182.960 ;
        RECT 58.810 181.960 59.070 182.280 ;
        RECT 59.730 181.960 59.990 182.280 ;
        RECT 56.110 180.520 56.710 180.660 ;
        RECT 57.430 180.600 57.690 180.920 ;
        RECT 58.350 180.600 58.610 180.920 ;
        RECT 58.870 180.775 59.010 181.960 ;
        RECT 59.260 181.085 59.540 181.455 ;
        RECT 56.110 176.840 56.250 180.520 ;
        RECT 56.500 179.725 56.780 180.095 ;
        RECT 57.430 179.920 57.690 180.240 ;
        RECT 56.510 179.580 56.770 179.725 ;
        RECT 56.570 178.735 56.710 179.580 ;
        RECT 56.500 178.365 56.780 178.735 ;
        RECT 57.490 178.110 57.630 179.920 ;
        RECT 58.410 178.735 58.550 180.600 ;
        RECT 58.800 180.405 59.080 180.775 ;
        RECT 59.330 180.240 59.470 181.085 ;
        RECT 59.790 180.240 59.930 181.960 ;
        RECT 59.270 180.150 59.530 180.240 ;
        RECT 58.870 180.010 59.530 180.150 ;
        RECT 58.340 178.365 58.620 178.735 ;
        RECT 57.890 178.110 58.150 178.200 ;
        RECT 56.500 177.685 56.780 178.055 ;
        RECT 57.490 177.970 58.150 178.110 ;
        RECT 57.890 177.880 58.150 177.970 ;
        RECT 56.050 176.520 56.310 176.840 ;
        RECT 56.050 175.160 56.310 175.480 ;
        RECT 56.110 174.655 56.250 175.160 ;
        RECT 56.040 174.285 56.320 174.655 ;
        RECT 56.050 173.800 56.310 174.120 ;
        RECT 56.110 173.100 56.250 173.800 ;
        RECT 55.590 172.780 55.850 173.100 ;
        RECT 56.050 172.780 56.310 173.100 ;
        RECT 56.570 172.420 56.710 177.685 ;
        RECT 56.970 177.200 57.230 177.520 ;
        RECT 57.030 176.840 57.170 177.200 ;
        RECT 57.420 177.005 57.700 177.375 ;
        RECT 56.970 176.520 57.230 176.840 ;
        RECT 56.510 172.100 56.770 172.420 ;
        RECT 57.030 171.820 57.170 176.520 ;
        RECT 57.490 174.120 57.630 177.005 ;
        RECT 57.950 174.800 58.090 177.880 ;
        RECT 58.340 177.685 58.620 178.055 ;
        RECT 58.870 177.860 59.010 180.010 ;
        RECT 59.270 179.920 59.530 180.010 ;
        RECT 59.730 179.920 59.990 180.240 ;
        RECT 57.890 174.480 58.150 174.800 ;
        RECT 57.430 173.800 57.690 174.120 ;
        RECT 57.890 173.975 58.150 174.120 ;
        RECT 57.880 173.605 58.160 173.975 ;
        RECT 57.890 172.330 58.150 172.420 ;
        RECT 58.410 172.330 58.550 177.685 ;
        RECT 58.810 177.540 59.070 177.860 ;
        RECT 59.270 177.770 59.530 177.860 ;
        RECT 59.790 177.770 59.930 179.920 ;
        RECT 60.190 179.580 60.450 179.900 ;
        RECT 60.250 177.860 60.390 179.580 ;
        RECT 59.270 177.630 59.930 177.770 ;
        RECT 59.270 177.540 59.530 177.630 ;
        RECT 60.190 177.540 60.450 177.860 ;
        RECT 59.270 176.520 59.530 176.840 ;
        RECT 58.810 173.800 59.070 174.120 ;
        RECT 58.870 172.420 59.010 173.800 ;
        RECT 57.890 172.190 58.550 172.330 ;
        RECT 57.890 172.100 58.150 172.190 ;
        RECT 58.810 172.100 59.070 172.420 ;
        RECT 57.030 171.680 58.550 171.820 ;
        RECT 56.050 170.060 56.310 170.380 ;
        RECT 55.190 167.600 55.790 167.740 ;
        RECT 55.130 166.660 55.390 166.980 ;
        RECT 54.670 166.320 54.930 166.640 ;
        RECT 52.830 161.900 53.090 162.220 ;
        RECT 54.210 161.900 54.470 162.220 ;
        RECT 54.270 161.540 54.410 161.900 ;
        RECT 54.210 161.220 54.470 161.540 ;
        RECT 53.290 160.540 53.550 160.860 ;
        RECT 51.910 160.200 52.170 160.520 ;
        RECT 51.450 159.070 51.710 159.160 ;
        RECT 51.450 158.930 53.030 159.070 ;
        RECT 51.450 158.840 51.710 158.930 ;
        RECT 50.530 156.120 50.790 156.440 ;
        RECT 51.910 155.780 52.170 156.100 ;
        RECT 51.450 155.440 51.710 155.760 ;
        RECT 51.510 155.080 51.650 155.440 ;
        RECT 50.990 154.760 51.250 155.080 ;
        RECT 51.450 154.760 51.710 155.080 ;
        RECT 49.150 153.400 49.410 153.720 ;
        RECT 50.070 153.060 50.330 153.380 ;
        RECT 50.130 152.700 50.270 153.060 ;
        RECT 51.050 153.040 51.190 154.760 ;
        RECT 50.990 152.720 51.250 153.040 ;
        RECT 49.610 152.380 49.870 152.700 ;
        RECT 50.070 152.380 50.330 152.700 ;
        RECT 49.670 151.000 49.810 152.380 ;
        RECT 49.610 150.680 49.870 151.000 ;
        RECT 50.130 150.660 50.270 152.380 ;
        RECT 51.970 150.660 52.110 155.780 ;
        RECT 52.890 155.420 53.030 158.930 ;
        RECT 53.350 158.820 53.490 160.540 ;
        RECT 53.290 158.500 53.550 158.820 ;
        RECT 52.830 155.100 53.090 155.420 ;
        RECT 53.290 155.100 53.550 155.420 ;
        RECT 52.370 153.400 52.630 153.720 ;
        RECT 52.890 153.460 53.030 155.100 ;
        RECT 53.350 154.060 53.490 155.100 ;
        RECT 53.290 153.740 53.550 154.060 ;
        RECT 53.750 153.460 54.010 153.720 ;
        RECT 52.890 153.400 54.010 153.460 ;
        RECT 52.430 152.950 52.570 153.400 ;
        RECT 52.890 153.320 53.950 153.400 ;
        RECT 52.830 152.950 53.090 153.040 ;
        RECT 52.430 152.810 53.090 152.950 ;
        RECT 52.830 152.720 53.090 152.810 ;
        RECT 50.070 150.340 50.330 150.660 ;
        RECT 51.910 150.340 52.170 150.660 ;
        RECT 52.830 150.340 53.090 150.660 ;
        RECT 48.230 149.660 48.490 149.980 ;
        RECT 52.890 149.640 53.030 150.340 ;
        RECT 52.830 149.320 53.090 149.640 ;
        RECT 53.350 147.600 53.490 153.320 ;
        RECT 53.750 152.040 54.010 152.360 ;
        RECT 53.810 150.660 53.950 152.040 ;
        RECT 54.730 151.000 54.870 166.320 ;
        RECT 55.190 154.060 55.330 166.660 ;
        RECT 55.130 153.740 55.390 154.060 ;
        RECT 55.130 152.380 55.390 152.700 ;
        RECT 54.670 150.680 54.930 151.000 ;
        RECT 55.190 150.660 55.330 152.380 ;
        RECT 53.750 150.340 54.010 150.660 ;
        RECT 55.130 150.340 55.390 150.660 ;
        RECT 55.190 148.620 55.330 150.340 ;
        RECT 55.130 148.300 55.390 148.620 ;
        RECT 55.650 147.940 55.790 167.600 ;
        RECT 56.110 166.980 56.250 170.060 ;
        RECT 56.510 169.040 56.770 169.360 ;
        RECT 57.890 169.040 58.150 169.360 ;
        RECT 56.050 166.660 56.310 166.980 ;
        RECT 56.570 164.260 56.710 169.040 ;
        RECT 56.970 166.660 57.230 166.980 ;
        RECT 56.510 163.940 56.770 164.260 ;
        RECT 56.050 160.880 56.310 161.200 ;
        RECT 56.110 158.480 56.250 160.880 ;
        RECT 56.510 160.540 56.770 160.860 ;
        RECT 56.050 158.160 56.310 158.480 ;
        RECT 56.570 157.800 56.710 160.540 ;
        RECT 57.030 157.800 57.170 166.660 ;
        RECT 57.950 163.920 58.090 169.040 ;
        RECT 58.410 166.980 58.550 171.680 ;
        RECT 58.870 167.320 59.010 172.100 ;
        RECT 59.330 172.080 59.470 176.520 ;
        RECT 59.720 175.645 60.000 176.015 ;
        RECT 59.790 174.120 59.930 175.645 ;
        RECT 60.190 174.480 60.450 174.800 ;
        RECT 59.730 173.800 59.990 174.120 ;
        RECT 60.250 172.615 60.390 174.480 ;
        RECT 60.180 172.245 60.460 172.615 ;
        RECT 59.270 171.760 59.530 172.080 ;
        RECT 58.810 167.000 59.070 167.320 ;
        RECT 58.350 166.660 58.610 166.980 ;
        RECT 58.410 164.940 58.550 166.660 ;
        RECT 58.350 164.620 58.610 164.940 ;
        RECT 57.890 163.600 58.150 163.920 ;
        RECT 56.510 157.480 56.770 157.800 ;
        RECT 56.970 157.480 57.230 157.800 ;
        RECT 57.950 156.780 58.090 163.600 ;
        RECT 58.350 161.560 58.610 161.880 ;
        RECT 58.410 160.520 58.550 161.560 ;
        RECT 58.350 160.200 58.610 160.520 ;
        RECT 57.890 156.460 58.150 156.780 ;
        RECT 57.890 155.100 58.150 155.420 ;
        RECT 56.510 153.740 56.770 154.060 ;
        RECT 56.050 152.720 56.310 153.040 ;
        RECT 56.110 150.660 56.250 152.720 ;
        RECT 56.050 150.340 56.310 150.660 ;
        RECT 56.570 149.640 56.710 153.740 ;
        RECT 57.950 153.040 58.090 155.100 ;
        RECT 58.810 154.760 59.070 155.080 ;
        RECT 58.870 153.040 59.010 154.760 ;
        RECT 56.970 152.950 57.230 153.040 ;
        RECT 56.970 152.810 57.630 152.950 ;
        RECT 56.970 152.720 57.230 152.810 ;
        RECT 57.490 150.660 57.630 152.810 ;
        RECT 57.890 152.720 58.150 153.040 ;
        RECT 58.810 152.720 59.070 153.040 ;
        RECT 57.950 151.000 58.090 152.720 ;
        RECT 57.890 150.680 58.150 151.000 ;
        RECT 57.430 150.340 57.690 150.660 ;
        RECT 57.890 150.000 58.150 150.320 ;
        RECT 56.510 149.320 56.770 149.640 ;
        RECT 55.590 147.620 55.850 147.940 ;
        RECT 53.290 147.280 53.550 147.600 ;
        RECT 47.310 144.900 47.570 145.220 ;
        RECT 55.650 144.540 55.790 147.620 ;
        RECT 57.950 145.560 58.090 150.000 ;
        RECT 58.870 148.620 59.010 152.720 ;
        RECT 58.810 148.300 59.070 148.620 ;
        RECT 58.870 147.260 59.010 148.300 ;
        RECT 59.330 147.600 59.470 171.760 ;
        RECT 59.730 171.650 59.990 171.740 ;
        RECT 60.250 171.650 60.390 172.245 ;
        RECT 59.730 171.510 60.390 171.650 ;
        RECT 59.730 171.420 59.990 171.510 ;
        RECT 60.710 170.575 60.850 187.400 ;
        RECT 61.630 183.980 61.770 190.800 ;
        RECT 62.550 187.720 62.690 198.200 ;
        RECT 63.010 189.420 63.150 204.740 ;
        RECT 63.410 204.400 63.670 204.720 ;
        RECT 63.470 192.335 63.610 204.400 ;
        RECT 63.930 203.215 64.070 210.520 ;
        RECT 65.310 208.460 65.450 210.860 ;
        RECT 66.170 209.160 66.430 209.480 ;
        RECT 65.250 208.140 65.510 208.460 ;
        RECT 65.710 207.295 65.970 207.440 ;
        RECT 65.700 206.925 65.980 207.295 ;
        RECT 65.250 205.080 65.510 205.400 ;
        RECT 64.790 204.400 65.050 204.720 ;
        RECT 64.330 203.720 64.590 204.040 ;
        RECT 63.860 202.845 64.140 203.215 ;
        RECT 64.390 195.880 64.530 203.720 ;
        RECT 64.850 199.135 64.990 204.400 ;
        RECT 64.780 198.765 65.060 199.135 ;
        RECT 65.310 198.340 65.450 205.080 ;
        RECT 65.710 204.740 65.970 205.060 ;
        RECT 64.850 198.200 65.450 198.340 ;
        RECT 64.330 195.560 64.590 195.880 ;
        RECT 63.400 191.965 63.680 192.335 ;
        RECT 62.950 189.100 63.210 189.420 ;
        RECT 63.410 188.080 63.670 188.400 ;
        RECT 62.490 187.400 62.750 187.720 ;
        RECT 63.470 186.700 63.610 188.080 ;
        RECT 63.410 186.380 63.670 186.700 ;
        RECT 62.030 184.680 62.290 185.000 ;
        RECT 61.570 183.660 61.830 183.980 ;
        RECT 61.570 183.210 61.830 183.300 ;
        RECT 62.090 183.210 62.230 184.680 ;
        RECT 61.570 183.070 62.230 183.210 ;
        RECT 62.480 183.125 62.760 183.495 ;
        RECT 63.470 183.300 63.610 186.380 ;
        RECT 63.870 185.700 64.130 186.020 ;
        RECT 61.570 182.980 61.830 183.070 ;
        RECT 62.090 181.260 62.230 183.070 ;
        RECT 62.490 182.980 62.750 183.125 ;
        RECT 63.410 182.980 63.670 183.300 ;
        RECT 62.490 182.300 62.750 182.620 ;
        RECT 62.950 182.300 63.210 182.620 ;
        RECT 62.030 180.940 62.290 181.260 ;
        RECT 61.570 180.260 61.830 180.580 ;
        RECT 61.110 179.920 61.370 180.240 ;
        RECT 61.170 178.540 61.310 179.920 ;
        RECT 61.110 178.220 61.370 178.540 ;
        RECT 61.110 177.540 61.370 177.860 ;
        RECT 61.170 175.820 61.310 177.540 ;
        RECT 61.630 176.840 61.770 180.260 ;
        RECT 61.570 176.520 61.830 176.840 ;
        RECT 61.110 175.500 61.370 175.820 ;
        RECT 61.170 175.140 61.310 175.500 ;
        RECT 61.110 174.820 61.370 175.140 ;
        RECT 61.570 174.820 61.830 175.140 ;
        RECT 61.100 174.285 61.380 174.655 ;
        RECT 61.110 174.140 61.370 174.285 ;
        RECT 60.640 170.205 60.920 170.575 ;
        RECT 61.170 169.700 61.310 174.140 ;
        RECT 61.630 172.420 61.770 174.820 ;
        RECT 62.090 174.800 62.230 180.940 ;
        RECT 62.550 178.200 62.690 182.300 ;
        RECT 62.490 177.880 62.750 178.200 ;
        RECT 62.490 177.200 62.750 177.520 ;
        RECT 62.550 176.840 62.690 177.200 ;
        RECT 62.490 176.520 62.750 176.840 ;
        RECT 62.490 175.500 62.750 175.820 ;
        RECT 62.550 175.335 62.690 175.500 ;
        RECT 62.480 174.965 62.760 175.335 ;
        RECT 62.030 174.480 62.290 174.800 ;
        RECT 62.490 174.480 62.750 174.800 ;
        RECT 61.570 172.100 61.830 172.420 ;
        RECT 62.550 171.740 62.690 174.480 ;
        RECT 63.010 172.615 63.150 182.300 ;
        RECT 63.470 180.240 63.610 182.980 ;
        RECT 63.930 181.260 64.070 185.700 ;
        RECT 64.850 182.280 64.990 198.200 ;
        RECT 65.250 195.560 65.510 195.880 ;
        RECT 65.310 194.260 65.450 195.560 ;
        RECT 65.770 194.860 65.910 204.740 ;
        RECT 66.230 196.220 66.370 209.160 ;
        RECT 66.690 198.455 66.830 215.085 ;
        RECT 69.390 212.220 69.650 212.540 ;
        RECT 69.450 210.840 69.590 212.220 ;
        RECT 69.840 211.005 70.120 211.375 ;
        RECT 69.390 210.520 69.650 210.840 ;
        RECT 67.090 210.180 67.350 210.500 ;
        RECT 67.550 210.180 67.810 210.500 ;
        RECT 68.470 210.180 68.730 210.500 ;
        RECT 67.150 206.615 67.290 210.180 ;
        RECT 67.080 206.245 67.360 206.615 ;
        RECT 67.090 205.420 67.350 205.740 ;
        RECT 67.150 204.720 67.290 205.420 ;
        RECT 67.090 204.400 67.350 204.720 ;
        RECT 67.150 200.300 67.290 204.400 ;
        RECT 67.090 199.980 67.350 200.300 ;
        RECT 67.610 199.620 67.750 210.180 ;
        RECT 68.010 207.460 68.270 207.780 ;
        RECT 68.070 205.740 68.210 207.460 ;
        RECT 68.010 205.420 68.270 205.740 ;
        RECT 68.530 204.720 68.670 210.180 ;
        RECT 69.910 207.295 70.050 211.005 ;
        RECT 68.930 206.780 69.190 207.100 ;
        RECT 69.840 206.925 70.120 207.295 ;
        RECT 68.990 204.720 69.130 206.780 ;
        RECT 69.390 206.440 69.650 206.760 ;
        RECT 69.450 205.740 69.590 206.440 ;
        RECT 69.390 205.420 69.650 205.740 ;
        RECT 69.840 204.885 70.120 205.255 ;
        RECT 68.470 204.400 68.730 204.720 ;
        RECT 68.930 204.400 69.190 204.720 ;
        RECT 69.390 204.400 69.650 204.720 ;
        RECT 69.450 201.175 69.590 204.400 ;
        RECT 69.380 200.805 69.660 201.175 ;
        RECT 68.010 199.980 68.270 200.300 ;
        RECT 67.550 199.300 67.810 199.620 ;
        RECT 66.620 198.085 66.900 198.455 ;
        RECT 67.080 196.725 67.360 197.095 ;
        RECT 66.170 195.900 66.430 196.220 ;
        RECT 66.630 195.560 66.890 195.880 ;
        RECT 65.710 194.540 65.970 194.860 ;
        RECT 65.310 194.120 65.910 194.260 ;
        RECT 65.770 193.840 65.910 194.120 ;
        RECT 65.710 193.520 65.970 193.840 ;
        RECT 65.250 186.380 65.510 186.700 ;
        RECT 65.310 184.910 65.450 186.380 ;
        RECT 65.770 185.680 65.910 193.520 ;
        RECT 66.170 191.140 66.430 191.460 ;
        RECT 65.710 185.360 65.970 185.680 ;
        RECT 65.310 184.770 65.910 184.910 ;
        RECT 64.790 181.960 65.050 182.280 ;
        RECT 63.870 180.940 64.130 181.260 ;
        RECT 64.790 180.260 65.050 180.580 ;
        RECT 63.410 179.920 63.670 180.240 ;
        RECT 63.860 179.725 64.140 180.095 ;
        RECT 63.930 179.300 64.070 179.725 ;
        RECT 63.470 179.160 64.070 179.300 ;
        RECT 63.470 177.520 63.610 179.160 ;
        RECT 64.850 177.520 64.990 180.260 ;
        RECT 65.770 178.620 65.910 184.770 ;
        RECT 66.230 183.980 66.370 191.140 ;
        RECT 66.170 183.660 66.430 183.980 ;
        RECT 65.310 178.480 65.910 178.620 ;
        RECT 65.310 177.860 65.450 178.480 ;
        RECT 66.160 178.365 66.440 178.735 ;
        RECT 65.250 177.540 65.510 177.860 ;
        RECT 65.700 177.685 65.980 178.055 ;
        RECT 63.410 177.200 63.670 177.520 ;
        RECT 64.790 177.200 65.050 177.520 ;
        RECT 64.850 176.840 64.990 177.200 ;
        RECT 63.410 176.520 63.670 176.840 ;
        RECT 64.790 176.520 65.050 176.840 ;
        RECT 62.940 172.245 63.220 172.615 ;
        RECT 62.490 171.420 62.750 171.740 ;
        RECT 63.470 171.255 63.610 176.520 ;
        RECT 64.330 174.655 64.590 174.800 ;
        RECT 64.320 174.285 64.600 174.655 ;
        RECT 64.790 174.480 65.050 174.800 ;
        RECT 64.850 174.120 64.990 174.480 ;
        RECT 64.790 173.800 65.050 174.120 ;
        RECT 64.780 172.925 65.060 173.295 ;
        RECT 64.850 171.740 64.990 172.925 ;
        RECT 65.310 171.820 65.450 177.540 ;
        RECT 65.770 174.800 65.910 177.685 ;
        RECT 65.710 174.480 65.970 174.800 ;
        RECT 65.700 173.605 65.980 173.975 ;
        RECT 65.770 172.420 65.910 173.605 ;
        RECT 66.230 173.100 66.370 178.365 ;
        RECT 66.170 172.780 66.430 173.100 ;
        RECT 66.690 172.760 66.830 195.560 ;
        RECT 67.150 183.495 67.290 196.725 ;
        RECT 68.070 193.840 68.210 199.980 ;
        RECT 69.910 199.960 70.050 204.885 ;
        RECT 69.850 199.640 70.110 199.960 ;
        RECT 68.470 199.300 68.730 199.620 ;
        RECT 68.530 196.900 68.670 199.300 ;
        RECT 68.470 196.580 68.730 196.900 ;
        RECT 69.850 196.580 70.110 196.900 ;
        RECT 69.390 196.240 69.650 196.560 ;
        RECT 68.930 193.860 69.190 194.180 ;
        RECT 68.010 193.520 68.270 193.840 ;
        RECT 68.000 191.965 68.280 192.335 ;
        RECT 67.550 190.120 67.810 190.440 ;
        RECT 67.080 183.125 67.360 183.495 ;
        RECT 67.090 182.300 67.350 182.620 ;
        RECT 67.150 180.240 67.290 182.300 ;
        RECT 67.610 180.240 67.750 190.120 ;
        RECT 67.090 179.920 67.350 180.240 ;
        RECT 67.550 179.920 67.810 180.240 ;
        RECT 67.090 179.240 67.350 179.560 ;
        RECT 67.150 178.200 67.290 179.240 ;
        RECT 67.090 177.880 67.350 178.200 ;
        RECT 66.630 172.440 66.890 172.760 ;
        RECT 65.710 172.100 65.970 172.420 ;
        RECT 67.150 171.990 67.290 177.880 ;
        RECT 67.540 177.685 67.820 178.055 ;
        RECT 67.610 175.140 67.750 177.685 ;
        RECT 68.070 175.820 68.210 191.965 ;
        RECT 68.990 190.440 69.130 193.860 ;
        RECT 69.450 192.140 69.590 196.240 ;
        RECT 69.390 191.820 69.650 192.140 ;
        RECT 69.450 191.120 69.590 191.820 ;
        RECT 69.390 190.800 69.650 191.120 ;
        RECT 68.930 190.120 69.190 190.440 ;
        RECT 68.470 184.680 68.730 185.000 ;
        RECT 68.530 179.560 68.670 184.680 ;
        RECT 68.990 180.240 69.130 190.120 ;
        RECT 69.390 189.100 69.650 189.420 ;
        RECT 69.450 181.260 69.590 189.100 ;
        RECT 69.390 180.940 69.650 181.260 ;
        RECT 69.380 180.405 69.660 180.775 ;
        RECT 68.930 179.920 69.190 180.240 ;
        RECT 68.470 179.240 68.730 179.560 ;
        RECT 68.010 175.500 68.270 175.820 ;
        RECT 67.550 174.820 67.810 175.140 ;
        RECT 68.530 174.540 68.670 179.240 ;
        RECT 68.930 178.450 69.190 178.540 ;
        RECT 69.450 178.450 69.590 180.405 ;
        RECT 68.930 178.310 69.590 178.450 ;
        RECT 68.930 178.220 69.190 178.310 ;
        RECT 68.930 177.540 69.190 177.860 ;
        RECT 68.990 176.840 69.130 177.540 ;
        RECT 69.390 176.860 69.650 177.180 ;
        RECT 68.930 176.520 69.190 176.840 ;
        RECT 67.610 174.400 68.670 174.540 ;
        RECT 67.610 172.420 67.750 174.400 ;
        RECT 68.010 173.975 68.270 174.120 ;
        RECT 68.000 173.605 68.280 173.975 ;
        RECT 67.550 172.100 67.810 172.420 ;
        RECT 66.230 171.850 67.290 171.990 ;
        RECT 63.870 171.420 64.130 171.740 ;
        RECT 64.790 171.420 65.050 171.740 ;
        RECT 65.310 171.680 65.910 171.820 ;
        RECT 63.400 170.885 63.680 171.255 ;
        RECT 62.950 170.060 63.210 170.380 ;
        RECT 59.730 169.380 59.990 169.700 ;
        RECT 61.110 169.380 61.370 169.700 ;
        RECT 59.790 158.480 59.930 169.380 ;
        RECT 63.010 169.360 63.150 170.060 ;
        RECT 62.950 169.040 63.210 169.360 ;
        RECT 63.410 169.040 63.670 169.360 ;
        RECT 63.930 169.270 64.070 171.420 ;
        RECT 64.790 169.895 65.050 170.040 ;
        RECT 64.780 169.525 65.060 169.895 ;
        RECT 65.250 169.270 65.510 169.360 ;
        RECT 63.930 169.130 65.510 169.270 ;
        RECT 63.470 166.300 63.610 169.040 ;
        RECT 63.410 165.980 63.670 166.300 ;
        RECT 63.930 164.260 64.070 169.130 ;
        RECT 65.250 169.040 65.510 169.130 ;
        RECT 64.790 168.360 65.050 168.680 ;
        RECT 64.850 167.320 64.990 168.360 ;
        RECT 64.790 167.000 65.050 167.320 ;
        RECT 65.770 167.060 65.910 171.680 ;
        RECT 66.230 167.660 66.370 171.850 ;
        RECT 67.080 170.885 67.360 171.255 ;
        RECT 66.630 169.040 66.890 169.360 ;
        RECT 66.170 167.340 66.430 167.660 ;
        RECT 63.870 163.940 64.130 164.260 ;
        RECT 61.110 162.920 61.370 163.240 ;
        RECT 61.570 162.920 61.830 163.240 ;
        RECT 61.170 162.220 61.310 162.920 ;
        RECT 61.110 161.900 61.370 162.220 ;
        RECT 61.170 161.540 61.310 161.900 ;
        RECT 61.110 161.220 61.370 161.540 ;
        RECT 60.190 160.880 60.450 161.200 ;
        RECT 60.250 158.480 60.390 160.880 ;
        RECT 61.170 158.480 61.310 161.220 ;
        RECT 61.630 158.820 61.770 162.920 ;
        RECT 62.490 161.560 62.750 161.880 ;
        RECT 61.570 158.500 61.830 158.820 ;
        RECT 59.730 158.160 59.990 158.480 ;
        RECT 60.190 158.160 60.450 158.480 ;
        RECT 61.110 158.160 61.370 158.480 ;
        RECT 61.170 153.040 61.310 158.160 ;
        RECT 62.550 158.140 62.690 161.560 ;
        RECT 62.950 160.880 63.210 161.200 ;
        RECT 63.010 158.480 63.150 160.880 ;
        RECT 64.850 159.500 64.990 167.000 ;
        RECT 65.770 166.920 66.370 167.060 ;
        RECT 65.710 166.320 65.970 166.640 ;
        RECT 65.770 162.220 65.910 166.320 ;
        RECT 65.710 161.900 65.970 162.220 ;
        RECT 63.410 159.180 63.670 159.500 ;
        RECT 64.790 159.180 65.050 159.500 ;
        RECT 62.950 158.160 63.210 158.480 ;
        RECT 62.490 157.820 62.750 158.140 ;
        RECT 62.950 157.480 63.210 157.800 ;
        RECT 61.110 152.720 61.370 153.040 ;
        RECT 59.730 150.340 59.990 150.660 ;
        RECT 59.790 148.620 59.930 150.340 ;
        RECT 61.170 148.620 61.310 152.720 ;
        RECT 62.490 152.610 62.750 152.700 ;
        RECT 63.010 152.610 63.150 157.480 ;
        RECT 63.470 153.720 63.610 159.180 ;
        RECT 63.870 158.500 64.130 158.820 ;
        RECT 63.930 154.060 64.070 158.500 ;
        RECT 66.230 155.420 66.370 166.920 ;
        RECT 66.690 160.520 66.830 169.040 ;
        RECT 66.630 160.200 66.890 160.520 ;
        RECT 66.170 155.100 66.430 155.420 ;
        RECT 63.870 153.740 64.130 154.060 ;
        RECT 63.410 153.400 63.670 153.720 ;
        RECT 62.490 152.470 63.150 152.610 ;
        RECT 62.490 152.380 62.750 152.470 ;
        RECT 62.550 149.980 62.690 152.380 ;
        RECT 63.470 151.340 63.610 153.400 ;
        RECT 63.410 151.020 63.670 151.340 ;
        RECT 62.490 149.660 62.750 149.980 ;
        RECT 59.730 148.300 59.990 148.620 ;
        RECT 61.110 148.300 61.370 148.620 ;
        RECT 63.930 147.600 64.070 153.740 ;
        RECT 67.150 153.040 67.290 170.885 ;
        RECT 67.550 169.090 67.810 169.410 ;
        RECT 67.610 166.300 67.750 169.090 ;
        RECT 68.070 167.320 68.210 173.605 ;
        RECT 68.470 172.100 68.730 172.420 ;
        RECT 68.530 169.700 68.670 172.100 ;
        RECT 68.470 169.380 68.730 169.700 ;
        RECT 68.990 169.020 69.130 176.520 ;
        RECT 69.450 174.800 69.590 176.860 ;
        RECT 69.910 175.480 70.050 196.580 ;
        RECT 69.850 175.160 70.110 175.480 ;
        RECT 69.390 174.480 69.650 174.800 ;
        RECT 69.850 172.615 70.110 172.760 ;
        RECT 69.840 172.245 70.120 172.615 ;
        RECT 69.850 169.270 70.110 169.360 ;
        RECT 69.450 169.130 70.110 169.270 ;
        RECT 68.930 168.700 69.190 169.020 ;
        RECT 68.010 167.000 68.270 167.320 ;
        RECT 68.920 166.805 69.200 167.175 ;
        RECT 67.550 165.980 67.810 166.300 ;
        RECT 68.470 161.220 68.730 161.540 ;
        RECT 68.530 159.160 68.670 161.220 ;
        RECT 68.470 158.840 68.730 159.160 ;
        RECT 68.010 158.160 68.270 158.480 ;
        RECT 67.550 155.780 67.810 156.100 ;
        RECT 67.610 153.040 67.750 155.780 ;
        RECT 68.070 154.060 68.210 158.160 ;
        RECT 68.530 157.800 68.670 158.840 ;
        RECT 68.470 157.480 68.730 157.800 ;
        RECT 68.990 156.780 69.130 166.805 ;
        RECT 69.450 160.520 69.590 169.130 ;
        RECT 69.850 169.040 70.110 169.130 ;
        RECT 69.850 166.890 70.110 166.980 ;
        RECT 70.370 166.890 70.510 219.280 ;
        RECT 71.680 219.000 71.960 223.000 ;
        RECT 74.900 219.000 75.180 223.000 ;
        RECT 76.350 219.280 77.870 219.420 ;
        RECT 71.750 213.415 71.890 219.000 ;
        RECT 74.970 218.175 75.110 219.000 ;
        RECT 74.900 217.805 75.180 218.175 ;
        RECT 71.680 213.045 71.960 213.415 ;
        RECT 71.230 210.520 71.490 210.840 ;
        RECT 70.770 208.140 71.030 208.460 ;
        RECT 70.830 203.895 70.970 208.140 ;
        RECT 70.760 203.525 71.040 203.895 ;
        RECT 70.770 202.020 71.030 202.340 ;
        RECT 70.830 196.560 70.970 202.020 ;
        RECT 70.770 196.240 71.030 196.560 ;
        RECT 71.290 193.160 71.430 210.520 ;
        RECT 73.070 210.180 73.330 210.500 ;
        RECT 73.130 209.820 73.270 210.180 ;
        RECT 73.070 209.500 73.330 209.820 ;
        RECT 71.690 204.740 71.950 205.060 ;
        RECT 72.140 204.885 72.420 205.255 ;
        RECT 72.150 204.740 72.410 204.885 ;
        RECT 71.750 204.040 71.890 204.740 ;
        RECT 71.690 203.720 71.950 204.040 ;
        RECT 72.610 193.520 72.870 193.840 ;
        RECT 71.230 192.840 71.490 193.160 ;
        RECT 72.150 192.840 72.410 193.160 ;
        RECT 71.290 188.400 71.430 192.840 ;
        RECT 72.210 188.740 72.350 192.840 ;
        RECT 72.150 188.420 72.410 188.740 ;
        RECT 71.230 188.080 71.490 188.400 ;
        RECT 72.670 188.140 72.810 193.520 ;
        RECT 73.130 189.080 73.270 209.500 ;
        RECT 75.370 207.800 75.630 208.120 ;
        RECT 75.430 207.440 75.570 207.800 ;
        RECT 73.530 207.120 73.790 207.440 ;
        RECT 75.370 207.120 75.630 207.440 ;
        RECT 73.590 203.215 73.730 207.120 ;
        RECT 74.450 203.720 74.710 204.040 ;
        RECT 73.520 202.845 73.800 203.215 ;
        RECT 73.990 202.700 74.250 203.020 ;
        RECT 73.520 194.685 73.800 195.055 ;
        RECT 73.070 188.760 73.330 189.080 ;
        RECT 70.770 186.380 71.030 186.700 ;
        RECT 70.830 180.920 70.970 186.380 ;
        RECT 70.770 180.600 71.030 180.920 ;
        RECT 70.770 179.580 71.030 179.900 ;
        RECT 69.850 166.750 70.510 166.890 ;
        RECT 69.850 166.660 70.110 166.750 ;
        RECT 69.840 166.125 70.120 166.495 ;
        RECT 69.850 165.980 70.110 166.125 ;
        RECT 70.370 164.940 70.510 166.750 ;
        RECT 70.830 166.300 70.970 179.580 ;
        RECT 71.290 177.180 71.430 188.080 ;
        RECT 72.670 188.000 73.270 188.140 ;
        RECT 72.610 187.400 72.870 187.720 ;
        RECT 72.670 185.680 72.810 187.400 ;
        RECT 73.130 186.360 73.270 188.000 ;
        RECT 73.070 186.040 73.330 186.360 ;
        RECT 72.610 185.360 72.870 185.680 ;
        RECT 71.690 183.660 71.950 183.980 ;
        RECT 71.750 180.240 71.890 183.660 ;
        RECT 72.610 183.320 72.870 183.640 ;
        RECT 71.690 179.920 71.950 180.240 ;
        RECT 72.150 179.920 72.410 180.240 ;
        RECT 71.230 176.860 71.490 177.180 ;
        RECT 72.210 176.580 72.350 179.920 ;
        RECT 72.670 177.520 72.810 183.320 ;
        RECT 73.070 177.540 73.330 177.860 ;
        RECT 72.610 177.200 72.870 177.520 ;
        RECT 71.290 176.440 72.350 176.580 ;
        RECT 71.290 175.820 71.430 176.440 ;
        RECT 72.670 175.820 72.810 177.200 ;
        RECT 71.230 175.500 71.490 175.820 ;
        RECT 72.150 175.500 72.410 175.820 ;
        RECT 72.610 175.500 72.870 175.820 ;
        RECT 71.230 172.100 71.490 172.420 ;
        RECT 71.690 172.100 71.950 172.420 ;
        RECT 71.290 170.040 71.430 172.100 ;
        RECT 71.230 169.720 71.490 170.040 ;
        RECT 71.750 169.360 71.890 172.100 ;
        RECT 71.690 169.040 71.950 169.360 ;
        RECT 71.230 167.230 71.490 167.320 ;
        RECT 71.750 167.230 71.890 169.040 ;
        RECT 71.230 167.090 71.890 167.230 ;
        RECT 71.230 167.000 71.490 167.090 ;
        RECT 70.770 165.980 71.030 166.300 ;
        RECT 70.310 164.620 70.570 164.940 ;
        RECT 70.770 164.620 71.030 164.940 ;
        RECT 69.850 163.260 70.110 163.580 ;
        RECT 69.910 161.880 70.050 163.260 ;
        RECT 69.850 161.560 70.110 161.880 ;
        RECT 70.310 161.220 70.570 161.540 ;
        RECT 69.850 160.540 70.110 160.860 ;
        RECT 69.390 160.200 69.650 160.520 ;
        RECT 68.930 156.460 69.190 156.780 ;
        RECT 68.930 155.780 69.190 156.100 ;
        RECT 68.010 153.740 68.270 154.060 ;
        RECT 68.990 153.040 69.130 155.780 ;
        RECT 69.450 155.420 69.590 160.200 ;
        RECT 69.910 159.500 70.050 160.540 ;
        RECT 70.370 160.430 70.510 161.220 ;
        RECT 70.830 160.520 70.970 164.620 ;
        RECT 71.230 161.560 71.490 161.880 ;
        RECT 70.770 160.430 71.030 160.520 ;
        RECT 70.370 160.290 71.030 160.430 ;
        RECT 69.850 159.180 70.110 159.500 ;
        RECT 70.370 156.780 70.510 160.290 ;
        RECT 70.770 160.200 71.030 160.290 ;
        RECT 71.290 158.480 71.430 161.560 ;
        RECT 71.750 159.500 71.890 167.090 ;
        RECT 72.210 166.980 72.350 175.500 ;
        RECT 72.610 174.820 72.870 175.140 ;
        RECT 72.670 169.360 72.810 174.820 ;
        RECT 72.610 169.040 72.870 169.360 ;
        RECT 72.150 166.660 72.410 166.980 ;
        RECT 72.670 166.300 72.810 169.040 ;
        RECT 73.130 167.175 73.270 177.540 ;
        RECT 73.590 171.740 73.730 194.685 ;
        RECT 74.050 188.740 74.190 202.700 ;
        RECT 74.510 194.180 74.650 203.720 ;
        RECT 74.450 193.860 74.710 194.180 ;
        RECT 75.370 193.860 75.630 194.180 ;
        RECT 74.440 192.645 74.720 193.015 ;
        RECT 73.990 188.420 74.250 188.740 ;
        RECT 74.510 185.535 74.650 192.645 ;
        RECT 75.430 191.460 75.570 193.860 ;
        RECT 75.370 191.140 75.630 191.460 ;
        RECT 75.370 190.460 75.630 190.780 ;
        RECT 74.910 189.100 75.170 189.420 ;
        RECT 74.970 186.895 75.110 189.100 ;
        RECT 74.900 186.525 75.180 186.895 ;
        RECT 75.430 186.020 75.570 190.460 ;
        RECT 75.830 188.420 76.090 188.740 ;
        RECT 75.370 185.700 75.630 186.020 ;
        RECT 74.440 185.165 74.720 185.535 ;
        RECT 73.990 184.680 74.250 185.000 ;
        RECT 74.050 183.300 74.190 184.680 ;
        RECT 73.990 182.980 74.250 183.300 ;
        RECT 74.910 182.980 75.170 183.300 ;
        RECT 74.970 177.860 75.110 182.980 ;
        RECT 75.430 180.920 75.570 185.700 ;
        RECT 75.370 180.600 75.630 180.920 ;
        RECT 75.890 180.240 76.030 188.420 ;
        RECT 75.830 179.920 76.090 180.240 ;
        RECT 76.350 179.300 76.490 219.280 ;
        RECT 77.730 218.740 77.870 219.280 ;
        RECT 78.120 219.000 78.400 223.000 ;
        RECT 81.340 219.000 81.620 223.000 ;
        RECT 84.560 219.000 84.840 223.000 ;
        RECT 87.780 219.000 88.060 223.000 ;
        RECT 91.000 219.000 91.280 223.000 ;
        RECT 78.190 218.740 78.330 219.000 ;
        RECT 77.730 218.600 78.330 218.740 ;
        RECT 77.660 215.765 77.940 216.135 ;
        RECT 77.200 208.965 77.480 209.335 ;
        RECT 77.270 207.780 77.410 208.965 ;
        RECT 77.210 207.460 77.470 207.780 ;
        RECT 77.730 202.680 77.870 215.765 ;
        RECT 78.130 214.600 78.390 214.920 ;
        RECT 78.190 203.950 78.330 214.600 ;
        RECT 79.510 214.260 79.770 214.580 ;
        RECT 79.570 211.180 79.710 214.260 ;
        RECT 81.410 214.095 81.550 219.000 ;
        RECT 81.340 213.725 81.620 214.095 ;
        RECT 80.430 212.900 80.690 213.220 ;
        RECT 79.510 210.860 79.770 211.180 ;
        RECT 79.050 210.180 79.310 210.500 ;
        RECT 79.960 210.325 80.240 210.695 ;
        RECT 78.590 209.840 78.850 210.160 ;
        RECT 78.650 204.720 78.790 209.840 ;
        RECT 79.110 207.295 79.250 210.180 ;
        RECT 80.030 209.820 80.170 210.325 ;
        RECT 79.970 209.500 80.230 209.820 ;
        RECT 80.030 207.440 80.170 209.500 ;
        RECT 79.040 206.925 79.320 207.295 ;
        RECT 79.970 207.120 80.230 207.440 ;
        RECT 79.510 206.440 79.770 206.760 ;
        RECT 78.590 204.400 78.850 204.720 ;
        RECT 78.190 203.810 79.250 203.950 ;
        RECT 77.670 202.360 77.930 202.680 ;
        RECT 79.110 201.060 79.250 203.810 ;
        RECT 79.570 202.000 79.710 206.440 ;
        RECT 80.490 202.000 80.630 212.900 ;
        RECT 80.890 210.015 81.150 210.160 ;
        RECT 80.880 209.645 81.160 210.015 ;
        RECT 84.100 209.645 84.380 210.015 ;
        RECT 82.270 209.160 82.530 209.480 ;
        RECT 83.190 209.160 83.450 209.480 ;
        RECT 81.810 204.740 82.070 205.060 ;
        RECT 82.330 204.970 82.470 209.160 ;
        RECT 83.250 207.780 83.390 209.160 ;
        RECT 83.190 207.460 83.450 207.780 ;
        RECT 82.730 207.120 82.990 207.440 ;
        RECT 82.790 206.615 82.930 207.120 ;
        RECT 83.650 206.780 83.910 207.100 ;
        RECT 82.720 206.245 83.000 206.615 ;
        RECT 83.710 205.820 83.850 206.780 ;
        RECT 84.170 206.760 84.310 209.645 ;
        RECT 84.110 206.440 84.370 206.760 ;
        RECT 83.710 205.740 84.310 205.820 ;
        RECT 83.710 205.680 84.370 205.740 ;
        RECT 84.110 205.420 84.370 205.680 ;
        RECT 83.650 204.970 83.910 205.060 ;
        RECT 82.330 204.830 83.910 204.970 ;
        RECT 83.650 204.740 83.910 204.830 ;
        RECT 79.510 201.680 79.770 202.000 ;
        RECT 80.430 201.680 80.690 202.000 ;
        RECT 81.350 201.680 81.610 202.000 ;
        RECT 78.190 200.920 79.250 201.060 ;
        RECT 76.750 198.960 77.010 199.280 ;
        RECT 76.810 196.900 76.950 198.960 ;
        RECT 78.190 198.600 78.330 200.920 ;
        RECT 78.580 200.125 78.860 200.495 ;
        RECT 78.590 199.980 78.850 200.125 ;
        RECT 78.650 199.620 78.790 199.980 ;
        RECT 79.110 199.620 79.250 200.920 ;
        RECT 78.590 199.300 78.850 199.620 ;
        RECT 79.050 199.300 79.310 199.620 ;
        RECT 79.500 199.445 79.780 199.815 ;
        RECT 79.050 198.620 79.310 198.940 ;
        RECT 78.130 198.280 78.390 198.600 ;
        RECT 78.590 197.260 78.850 197.580 ;
        RECT 76.750 196.580 77.010 196.900 ;
        RECT 77.670 193.180 77.930 193.500 ;
        RECT 77.730 192.100 77.870 193.180 ;
        RECT 77.270 191.960 77.870 192.100 ;
        RECT 76.750 191.480 77.010 191.800 ;
        RECT 75.890 179.160 76.490 179.300 ;
        RECT 74.910 177.540 75.170 177.860 ;
        RECT 73.990 177.200 74.250 177.520 ;
        RECT 75.890 177.375 76.030 179.160 ;
        RECT 76.290 178.220 76.550 178.540 ;
        RECT 74.050 176.840 74.190 177.200 ;
        RECT 75.820 177.005 76.100 177.375 ;
        RECT 73.990 176.520 74.250 176.840 ;
        RECT 75.370 175.500 75.630 175.820 ;
        RECT 73.990 174.480 74.250 174.800 ;
        RECT 74.450 174.480 74.710 174.800 ;
        RECT 74.050 171.740 74.190 174.480 ;
        RECT 74.510 173.180 74.650 174.480 ;
        RECT 74.510 173.040 75.110 173.180 ;
        RECT 74.450 172.100 74.710 172.420 ;
        RECT 73.530 171.420 73.790 171.740 ;
        RECT 73.990 171.420 74.250 171.740 ;
        RECT 74.510 171.400 74.650 172.100 ;
        RECT 74.970 171.935 75.110 173.040 ;
        RECT 74.900 171.565 75.180 171.935 ;
        RECT 75.430 171.400 75.570 175.500 ;
        RECT 76.350 175.335 76.490 178.220 ;
        RECT 76.810 176.695 76.950 191.480 ;
        RECT 77.270 185.420 77.410 191.960 ;
        RECT 77.670 186.100 77.930 186.360 ;
        RECT 77.670 186.040 78.330 186.100 ;
        RECT 77.730 185.960 78.330 186.040 ;
        RECT 78.190 185.680 78.330 185.960 ;
        RECT 77.670 185.420 77.930 185.680 ;
        RECT 77.270 185.360 77.930 185.420 ;
        RECT 78.130 185.360 78.390 185.680 ;
        RECT 77.270 185.280 77.870 185.360 ;
        RECT 77.270 177.520 77.410 185.280 ;
        RECT 78.130 184.680 78.390 185.000 ;
        RECT 78.190 182.280 78.330 184.680 ;
        RECT 78.130 181.960 78.390 182.280 ;
        RECT 77.210 177.200 77.470 177.520 ;
        RECT 76.740 176.325 77.020 176.695 ;
        RECT 76.280 174.965 76.560 175.335 ;
        RECT 76.750 175.160 77.010 175.480 ;
        RECT 77.210 175.160 77.470 175.480 ;
        RECT 75.830 174.480 76.090 174.800 ;
        RECT 75.890 172.760 76.030 174.480 ;
        RECT 75.830 172.440 76.090 172.760 ;
        RECT 76.290 172.100 76.550 172.420 ;
        RECT 75.830 171.420 76.090 171.740 ;
        RECT 74.510 171.260 75.570 171.400 ;
        RECT 74.440 170.205 74.720 170.575 ;
        RECT 75.430 170.460 75.570 171.260 ;
        RECT 75.890 171.255 76.030 171.420 ;
        RECT 75.820 170.885 76.100 171.255 ;
        RECT 75.430 170.320 76.030 170.460 ;
        RECT 74.510 169.360 74.650 170.205 ;
        RECT 75.370 169.720 75.630 170.040 ;
        RECT 74.450 169.040 74.710 169.360 ;
        RECT 73.530 168.360 73.790 168.680 ;
        RECT 73.060 166.805 73.340 167.175 ;
        RECT 73.070 166.660 73.330 166.805 ;
        RECT 72.610 165.980 72.870 166.300 ;
        RECT 72.670 164.940 72.810 165.980 ;
        RECT 73.070 165.640 73.330 165.960 ;
        RECT 72.610 164.620 72.870 164.940 ;
        RECT 72.610 163.600 72.870 163.920 ;
        RECT 72.670 160.860 72.810 163.600 ;
        RECT 73.130 162.220 73.270 165.640 ;
        RECT 73.590 164.600 73.730 168.360 ;
        RECT 73.990 166.660 74.250 166.980 ;
        RECT 74.450 166.660 74.710 166.980 ;
        RECT 74.050 164.940 74.190 166.660 ;
        RECT 73.990 164.620 74.250 164.940 ;
        RECT 73.530 164.280 73.790 164.600 ;
        RECT 73.980 164.085 74.260 164.455 ;
        RECT 74.510 164.260 74.650 166.660 ;
        RECT 75.430 165.960 75.570 169.720 ;
        RECT 75.890 169.020 76.030 170.320 ;
        RECT 76.350 170.040 76.490 172.100 ;
        RECT 76.290 169.720 76.550 170.040 ;
        RECT 75.830 168.700 76.090 169.020 ;
        RECT 75.890 167.320 76.030 168.700 ;
        RECT 75.830 167.000 76.090 167.320 ;
        RECT 76.290 166.660 76.550 166.980 ;
        RECT 76.350 166.300 76.490 166.660 ;
        RECT 76.290 165.980 76.550 166.300 ;
        RECT 75.370 165.640 75.630 165.960 ;
        RECT 75.370 164.620 75.630 164.940 ;
        RECT 74.050 163.920 74.190 164.085 ;
        RECT 74.450 163.940 74.710 164.260 ;
        RECT 73.990 163.600 74.250 163.920 ;
        RECT 74.900 163.405 75.180 163.775 ;
        RECT 74.970 163.240 75.110 163.405 ;
        RECT 74.910 162.920 75.170 163.240 ;
        RECT 75.430 162.220 75.570 164.620 ;
        RECT 76.810 163.920 76.950 175.160 ;
        RECT 77.270 172.615 77.410 175.160 ;
        RECT 77.200 172.245 77.480 172.615 ;
        RECT 77.200 169.525 77.480 169.895 ;
        RECT 77.270 166.300 77.410 169.525 ;
        RECT 78.190 169.020 78.330 181.960 ;
        RECT 78.650 180.920 78.790 197.260 ;
        RECT 79.110 192.335 79.250 198.620 ;
        RECT 79.570 193.500 79.710 199.445 ;
        RECT 80.430 196.415 80.690 196.560 ;
        RECT 79.970 195.900 80.230 196.220 ;
        RECT 80.420 196.045 80.700 196.415 ;
        RECT 80.890 196.240 81.150 196.560 ;
        RECT 80.030 193.500 80.170 195.900 ;
        RECT 80.430 195.560 80.690 195.880 ;
        RECT 80.950 195.735 81.090 196.240 ;
        RECT 79.510 193.180 79.770 193.500 ;
        RECT 79.970 193.180 80.230 193.500 ;
        RECT 79.040 191.965 79.320 192.335 ;
        RECT 79.050 191.140 79.310 191.460 ;
        RECT 79.110 185.000 79.250 191.140 ;
        RECT 79.050 184.680 79.310 185.000 ;
        RECT 79.050 182.300 79.310 182.620 ;
        RECT 78.590 180.600 78.850 180.920 ;
        RECT 79.110 180.240 79.250 182.300 ;
        RECT 79.050 179.920 79.310 180.240 ;
        RECT 79.050 178.220 79.310 178.540 ;
        RECT 79.110 177.430 79.250 178.220 ;
        RECT 79.570 178.200 79.710 193.180 ;
        RECT 80.490 191.120 80.630 195.560 ;
        RECT 80.880 195.365 81.160 195.735 ;
        RECT 81.410 193.695 81.550 201.680 ;
        RECT 81.340 193.325 81.620 193.695 ;
        RECT 81.350 191.820 81.610 192.140 ;
        RECT 80.890 191.140 81.150 191.460 ;
        RECT 80.430 190.800 80.690 191.120 ;
        RECT 79.970 190.460 80.230 190.780 ;
        RECT 79.510 177.880 79.770 178.200 ;
        RECT 79.110 177.290 79.710 177.430 ;
        RECT 78.130 168.700 78.390 169.020 ;
        RECT 78.130 166.320 78.390 166.640 ;
        RECT 78.590 166.320 78.850 166.640 ;
        RECT 77.210 165.980 77.470 166.300 ;
        RECT 78.190 164.260 78.330 166.320 ;
        RECT 78.130 163.940 78.390 164.260 ;
        RECT 76.750 163.600 77.010 163.920 ;
        RECT 73.070 161.900 73.330 162.220 ;
        RECT 75.370 161.900 75.630 162.220 ;
        RECT 73.530 161.560 73.790 161.880 ;
        RECT 74.450 161.560 74.710 161.880 ;
        RECT 72.610 160.540 72.870 160.860 ;
        RECT 71.690 159.180 71.950 159.500 ;
        RECT 71.230 158.160 71.490 158.480 ;
        RECT 70.310 156.460 70.570 156.780 ;
        RECT 69.850 155.440 70.110 155.760 ;
        RECT 69.390 155.100 69.650 155.420 ;
        RECT 69.910 153.040 70.050 155.440 ;
        RECT 73.590 153.720 73.730 161.560 ;
        RECT 74.510 158.480 74.650 161.560 ;
        RECT 76.810 159.500 76.950 163.600 ;
        RECT 78.650 163.580 78.790 166.320 ;
        RECT 79.570 165.960 79.710 177.290 ;
        RECT 80.030 175.820 80.170 190.460 ;
        RECT 80.950 190.295 81.090 191.140 ;
        RECT 80.880 189.925 81.160 190.295 ;
        RECT 80.420 187.885 80.700 188.255 ;
        RECT 79.970 175.500 80.230 175.820 ;
        RECT 79.960 174.965 80.240 175.335 ;
        RECT 80.030 167.230 80.170 174.965 ;
        RECT 80.490 173.100 80.630 187.885 ;
        RECT 80.890 185.360 81.150 185.680 ;
        RECT 80.950 176.840 81.090 185.360 ;
        RECT 80.890 176.520 81.150 176.840 ;
        RECT 80.880 175.645 81.160 176.015 ;
        RECT 80.430 172.780 80.690 173.100 ;
        RECT 80.030 167.090 80.630 167.230 ;
        RECT 79.970 166.320 80.230 166.640 ;
        RECT 79.510 165.640 79.770 165.960 ;
        RECT 78.590 163.260 78.850 163.580 ;
        RECT 78.120 160.685 78.400 161.055 ;
        RECT 78.190 159.500 78.330 160.685 ;
        RECT 76.750 159.180 77.010 159.500 ;
        RECT 78.130 159.180 78.390 159.500 ;
        RECT 74.450 158.160 74.710 158.480 ;
        RECT 78.650 157.540 78.790 163.260 ;
        RECT 79.050 162.920 79.310 163.240 ;
        RECT 79.110 158.480 79.250 162.920 ;
        RECT 79.050 158.160 79.310 158.480 ;
        RECT 80.030 158.140 80.170 166.320 ;
        RECT 80.490 163.920 80.630 167.090 ;
        RECT 80.950 166.640 81.090 175.645 ;
        RECT 81.410 173.100 81.550 191.820 ;
        RECT 81.870 191.540 82.010 204.740 ;
        RECT 84.630 204.460 84.770 219.000 ;
        RECT 85.480 211.685 85.760 212.055 ;
        RECT 85.550 210.500 85.690 211.685 ;
        RECT 85.490 210.180 85.750 210.500 ;
        RECT 85.030 209.840 85.290 210.160 ;
        RECT 84.170 204.320 84.770 204.460 ;
        RECT 82.270 201.340 82.530 201.660 ;
        RECT 82.330 201.175 82.470 201.340 ;
        RECT 82.260 200.805 82.540 201.175 ;
        RECT 82.270 199.980 82.530 200.300 ;
        RECT 82.330 199.620 82.470 199.980 ;
        RECT 82.270 199.300 82.530 199.620 ;
        RECT 83.650 199.300 83.910 199.620 ;
        RECT 82.730 196.920 82.990 197.240 ;
        RECT 82.270 193.180 82.530 193.500 ;
        RECT 82.330 192.140 82.470 193.180 ;
        RECT 82.270 191.820 82.530 192.140 ;
        RECT 81.870 191.400 82.470 191.540 ;
        RECT 82.330 187.720 82.470 191.400 ;
        RECT 82.270 187.400 82.530 187.720 ;
        RECT 81.810 184.680 82.070 185.000 ;
        RECT 81.870 180.920 82.010 184.680 ;
        RECT 82.330 183.640 82.470 187.400 ;
        RECT 82.270 183.320 82.530 183.640 ;
        RECT 81.810 180.600 82.070 180.920 ;
        RECT 82.270 179.920 82.530 180.240 ;
        RECT 82.330 178.540 82.470 179.920 ;
        RECT 82.270 178.220 82.530 178.540 ;
        RECT 81.810 176.860 82.070 177.180 ;
        RECT 81.870 175.820 82.010 176.860 ;
        RECT 82.270 176.520 82.530 176.840 ;
        RECT 81.810 175.500 82.070 175.820 ;
        RECT 81.350 172.780 81.610 173.100 ;
        RECT 80.890 166.320 81.150 166.640 ;
        RECT 80.890 165.640 81.150 165.960 ;
        RECT 80.430 163.600 80.690 163.920 ;
        RECT 80.950 160.940 81.090 165.640 ;
        RECT 81.410 161.880 81.550 172.780 ;
        RECT 81.870 169.270 82.010 175.500 ;
        RECT 82.330 175.140 82.470 176.520 ;
        RECT 82.270 174.820 82.530 175.140 ;
        RECT 82.790 169.700 82.930 196.920 ;
        RECT 83.190 196.240 83.450 196.560 ;
        RECT 83.250 192.140 83.390 196.240 ;
        RECT 83.190 191.820 83.450 192.140 ;
        RECT 83.190 190.460 83.450 190.780 ;
        RECT 83.250 189.420 83.390 190.460 ;
        RECT 83.190 189.100 83.450 189.420 ;
        RECT 83.190 188.420 83.450 188.740 ;
        RECT 83.250 186.700 83.390 188.420 ;
        RECT 83.190 186.380 83.450 186.700 ;
        RECT 83.190 185.020 83.450 185.340 ;
        RECT 83.250 180.920 83.390 185.020 ;
        RECT 83.710 183.380 83.850 199.300 ;
        RECT 84.170 189.080 84.310 204.320 ;
        RECT 85.090 197.580 85.230 209.840 ;
        RECT 85.480 207.605 85.760 207.975 ;
        RECT 85.550 207.440 85.690 207.605 ;
        RECT 85.490 207.120 85.750 207.440 ;
        RECT 87.330 199.980 87.590 200.300 ;
        RECT 85.950 199.300 86.210 199.620 ;
        RECT 85.030 197.260 85.290 197.580 ;
        RECT 84.570 196.240 84.830 196.560 ;
        RECT 84.630 194.860 84.770 196.240 ;
        RECT 85.030 195.560 85.290 195.880 ;
        RECT 84.570 194.540 84.830 194.860 ;
        RECT 85.090 194.520 85.230 195.560 ;
        RECT 85.030 194.200 85.290 194.520 ;
        RECT 85.490 193.860 85.750 194.180 ;
        RECT 85.030 190.800 85.290 191.120 ;
        RECT 84.570 190.120 84.830 190.440 ;
        RECT 84.110 188.760 84.370 189.080 ;
        RECT 83.710 183.240 84.310 183.380 ;
        RECT 84.170 182.960 84.310 183.240 ;
        RECT 84.110 182.640 84.370 182.960 ;
        RECT 83.190 180.600 83.450 180.920 ;
        RECT 83.650 175.500 83.910 175.820 ;
        RECT 83.710 175.140 83.850 175.500 ;
        RECT 83.650 174.820 83.910 175.140 ;
        RECT 83.190 174.480 83.450 174.800 ;
        RECT 83.250 173.295 83.390 174.480 ;
        RECT 83.180 172.925 83.460 173.295 ;
        RECT 82.730 169.380 82.990 169.700 ;
        RECT 82.270 169.270 82.530 169.360 ;
        RECT 81.870 169.130 82.530 169.270 ;
        RECT 82.270 169.040 82.530 169.130 ;
        RECT 81.800 167.485 82.080 167.855 ;
        RECT 81.810 167.340 82.070 167.485 ;
        RECT 82.270 166.320 82.530 166.640 ;
        RECT 82.330 165.960 82.470 166.320 ;
        RECT 81.810 165.640 82.070 165.960 ;
        RECT 82.270 165.640 82.530 165.960 ;
        RECT 81.350 161.560 81.610 161.880 ;
        RECT 80.950 160.800 81.550 160.940 ;
        RECT 79.970 157.820 80.230 158.140 ;
        RECT 79.050 157.540 79.310 157.800 ;
        RECT 78.650 157.480 79.310 157.540 ;
        RECT 78.650 157.400 79.250 157.480 ;
        RECT 79.110 156.440 79.250 157.400 ;
        RECT 79.050 156.120 79.310 156.440 ;
        RECT 79.510 154.760 79.770 155.080 ;
        RECT 73.530 153.400 73.790 153.720 ;
        RECT 65.710 152.720 65.970 153.040 ;
        RECT 67.090 152.720 67.350 153.040 ;
        RECT 67.550 152.720 67.810 153.040 ;
        RECT 68.930 152.720 69.190 153.040 ;
        RECT 69.850 152.720 70.110 153.040 ;
        RECT 79.570 152.895 79.710 154.760 ;
        RECT 64.790 152.380 65.050 152.700 ;
        RECT 64.850 149.640 64.990 152.380 ;
        RECT 65.770 150.660 65.910 152.720 ;
        RECT 66.170 152.040 66.430 152.360 ;
        RECT 66.230 151.000 66.370 152.040 ;
        RECT 67.150 151.000 67.290 152.720 ;
        RECT 79.500 152.525 79.780 152.895 ;
        RECT 79.510 152.380 79.770 152.525 ;
        RECT 66.170 150.680 66.430 151.000 ;
        RECT 67.090 150.680 67.350 151.000 ;
        RECT 65.710 150.340 65.970 150.660 ;
        RECT 80.030 149.980 80.170 157.820 ;
        RECT 80.430 155.780 80.690 156.100 ;
        RECT 80.490 154.255 80.630 155.780 ;
        RECT 81.410 155.760 81.550 160.800 ;
        RECT 81.870 156.100 82.010 165.640 ;
        RECT 82.260 164.085 82.540 164.455 ;
        RECT 82.330 156.780 82.470 164.085 ;
        RECT 82.790 163.920 82.930 169.380 ;
        RECT 83.250 166.300 83.390 172.925 ;
        RECT 84.170 167.660 84.310 182.640 ;
        RECT 84.630 174.120 84.770 190.120 ;
        RECT 85.090 186.215 85.230 190.800 ;
        RECT 85.020 185.845 85.300 186.215 ;
        RECT 85.030 185.360 85.290 185.680 ;
        RECT 85.090 183.980 85.230 185.360 ;
        RECT 85.030 183.660 85.290 183.980 ;
        RECT 85.550 181.455 85.690 193.860 ;
        RECT 86.010 184.855 86.150 199.300 ;
        RECT 86.860 193.325 87.140 193.695 ;
        RECT 86.410 185.020 86.670 185.340 ;
        RECT 85.940 184.485 86.220 184.855 ;
        RECT 85.480 181.085 85.760 181.455 ;
        RECT 85.030 179.240 85.290 179.560 ;
        RECT 85.090 178.055 85.230 179.240 ;
        RECT 85.020 177.685 85.300 178.055 ;
        RECT 85.020 174.285 85.300 174.655 ;
        RECT 86.470 174.460 86.610 185.020 ;
        RECT 86.930 175.820 87.070 193.325 ;
        RECT 87.390 185.340 87.530 199.980 ;
        RECT 87.330 185.020 87.590 185.340 ;
        RECT 87.850 180.095 87.990 219.000 ;
        RECT 91.070 213.415 91.210 219.000 ;
        RECT 91.000 213.045 91.280 213.415 ;
        RECT 87.780 179.725 88.060 180.095 ;
        RECT 86.870 175.500 87.130 175.820 ;
        RECT 85.090 174.120 85.230 174.285 ;
        RECT 86.410 174.140 86.670 174.460 ;
        RECT 84.570 173.800 84.830 174.120 ;
        RECT 85.030 173.800 85.290 174.120 ;
        RECT 84.110 167.340 84.370 167.660 ;
        RECT 83.190 165.980 83.450 166.300 ;
        RECT 82.730 163.600 82.990 163.920 ;
        RECT 83.190 163.600 83.450 163.920 ;
        RECT 83.250 162.220 83.390 163.600 ;
        RECT 83.190 161.900 83.450 162.220 ;
        RECT 84.170 158.480 84.310 167.340 ;
        RECT 85.490 167.000 85.750 167.320 ;
        RECT 84.570 165.870 84.830 165.960 ;
        RECT 84.570 165.730 85.230 165.870 ;
        RECT 84.570 165.640 84.830 165.730 ;
        RECT 84.570 163.600 84.830 163.920 ;
        RECT 84.630 158.480 84.770 163.600 ;
        RECT 84.110 158.160 84.370 158.480 ;
        RECT 84.570 158.160 84.830 158.480 ;
        RECT 82.730 157.480 82.990 157.800 ;
        RECT 82.270 156.460 82.530 156.780 ;
        RECT 81.810 155.780 82.070 156.100 ;
        RECT 81.350 155.440 81.610 155.760 ;
        RECT 80.420 153.885 80.700 154.255 ;
        RECT 82.790 153.040 82.930 157.480 ;
        RECT 83.640 157.285 83.920 157.655 ;
        RECT 83.710 154.060 83.850 157.285 ;
        RECT 85.090 156.780 85.230 165.730 ;
        RECT 85.550 157.800 85.690 167.000 ;
        RECT 85.490 157.480 85.750 157.800 ;
        RECT 85.030 156.460 85.290 156.780 ;
        RECT 84.570 156.120 84.830 156.440 ;
        RECT 83.650 153.740 83.910 154.060 ;
        RECT 82.730 152.720 82.990 153.040 ;
        RECT 79.970 149.660 80.230 149.980 ;
        RECT 64.790 149.320 65.050 149.640 ;
        RECT 64.850 148.280 64.990 149.320 ;
        RECT 84.630 148.620 84.770 156.120 ;
        RECT 85.550 155.420 85.690 157.480 ;
        RECT 86.930 156.440 87.070 175.500 ;
        RECT 86.870 156.120 87.130 156.440 ;
        RECT 85.490 155.100 85.750 155.420 ;
        RECT 85.550 153.720 85.690 155.100 ;
        RECT 85.490 153.400 85.750 153.720 ;
        RECT 85.480 150.485 85.760 150.855 ;
        RECT 85.490 150.340 85.750 150.485 ;
        RECT 84.570 148.300 84.830 148.620 ;
        RECT 64.790 147.960 65.050 148.280 ;
        RECT 59.270 147.280 59.530 147.600 ;
        RECT 62.950 147.280 63.210 147.600 ;
        RECT 63.870 147.280 64.130 147.600 ;
        RECT 58.810 146.940 59.070 147.260 ;
        RECT 57.890 145.240 58.150 145.560 ;
        RECT 58.870 144.880 59.010 146.940 ;
        RECT 63.010 145.220 63.150 147.280 ;
        RECT 63.930 145.220 64.070 147.280 ;
        RECT 85.020 147.085 85.300 147.455 ;
        RECT 85.030 146.940 85.290 147.085 ;
        RECT 62.950 144.900 63.210 145.220 ;
        RECT 63.870 144.900 64.130 145.220 ;
        RECT 58.810 144.560 59.070 144.880 ;
        RECT 85.490 144.560 85.750 144.880 ;
        RECT 55.590 144.220 55.850 144.540 ;
        RECT 46.390 143.880 46.650 144.200 ;
        RECT 85.550 144.055 85.690 144.560 ;
        RECT 42.710 142.860 42.970 143.180 ;
        RECT 43.170 142.860 43.430 143.180 ;
        RECT 41.790 142.520 42.050 142.840 ;
        RECT 40.410 142.180 40.670 142.500 ;
        RECT 43.230 142.160 43.370 142.860 ;
        RECT 46.450 142.160 46.590 143.880 ;
        RECT 85.480 143.685 85.760 144.055 ;
        RECT 23.390 141.840 23.650 142.160 ;
        RECT 33.050 141.840 33.310 142.160 ;
        RECT 36.730 141.840 36.990 142.160 ;
        RECT 39.950 142.070 40.210 142.160 ;
        RECT 39.550 141.930 40.210 142.070 ;
        RECT 23.450 133.930 23.590 141.840 ;
        RECT 33.110 133.930 33.250 141.840 ;
        RECT 34.780 140.625 36.320 140.995 ;
        RECT 36.790 136.460 36.930 141.840 ;
        RECT 36.330 136.320 36.930 136.460 ;
        RECT 36.330 133.930 36.470 136.320 ;
        RECT 39.550 133.930 39.690 141.930 ;
        RECT 39.950 141.840 40.210 141.930 ;
        RECT 43.170 141.840 43.430 142.160 ;
        RECT 46.390 141.840 46.650 142.160 ;
        RECT 42.710 141.500 42.970 141.820 ;
        RECT 42.770 133.930 42.910 141.500 ;
        RECT 45.930 141.160 46.190 141.480 ;
        RECT 45.990 133.930 46.130 141.160 ;
        RECT 23.380 129.930 23.660 133.930 ;
        RECT 33.040 129.930 33.320 133.930 ;
        RECT 36.260 129.930 36.540 133.930 ;
        RECT 39.480 129.930 39.760 133.930 ;
        RECT 42.700 129.930 42.980 133.930 ;
        RECT 45.920 129.930 46.200 133.930 ;
      LAYER met3 ;
        RECT 29.080 222.220 29.460 222.230 ;
        RECT 88.760 222.220 92.760 222.370 ;
        RECT 29.080 221.920 92.760 222.220 ;
        RECT 29.080 221.910 29.460 221.920 ;
        RECT 88.760 221.770 92.760 221.920 ;
        RECT 20.595 218.820 20.925 218.835 ;
        RECT 88.760 218.820 92.760 218.970 ;
        RECT 20.595 218.520 92.760 218.820 ;
        RECT 20.595 218.505 20.925 218.520 ;
        RECT 88.760 218.370 92.760 218.520 ;
        RECT 16.200 218.140 16.580 218.150 ;
        RECT 74.875 218.140 75.205 218.155 ;
        RECT 16.200 217.840 75.205 218.140 ;
        RECT 16.200 217.830 16.580 217.840 ;
        RECT 74.875 217.825 75.205 217.840 ;
        RECT 10.475 216.100 10.805 216.115 ;
        RECT 24.480 216.100 24.860 216.110 ;
        RECT 10.475 215.800 24.860 216.100 ;
        RECT 10.475 215.785 10.805 215.800 ;
        RECT 24.480 215.790 24.860 215.800 ;
        RECT 61.995 216.100 62.325 216.115 ;
        RECT 77.635 216.100 77.965 216.115 ;
        RECT 61.995 215.800 77.965 216.100 ;
        RECT 61.995 215.785 62.325 215.800 ;
        RECT 77.635 215.785 77.965 215.800 ;
        RECT 40.120 215.420 40.500 215.430 ;
        RECT 65.215 215.420 65.545 215.435 ;
        RECT 40.120 215.120 65.545 215.420 ;
        RECT 40.120 215.110 40.500 215.120 ;
        RECT 65.215 215.105 65.545 215.120 ;
        RECT 66.595 215.420 66.925 215.435 ;
        RECT 88.760 215.420 92.760 215.570 ;
        RECT 66.595 215.120 92.760 215.420 ;
        RECT 66.595 215.105 66.925 215.120 ;
        RECT 88.760 214.970 92.760 215.120 ;
        RECT 29.335 214.060 29.665 214.075 ;
        RECT 49.115 214.060 49.445 214.075 ;
        RECT 29.335 213.760 49.445 214.060 ;
        RECT 29.335 213.745 29.665 213.760 ;
        RECT 49.115 213.745 49.445 213.760 ;
        RECT 56.680 214.060 57.060 214.070 ;
        RECT 81.315 214.060 81.645 214.075 ;
        RECT 56.680 213.760 81.645 214.060 ;
        RECT 56.680 213.750 57.060 213.760 ;
        RECT 81.315 213.745 81.645 213.760 ;
        RECT 20.800 213.380 21.180 213.390 ;
        RECT 23.355 213.380 23.685 213.395 ;
        RECT 20.800 213.080 23.685 213.380 ;
        RECT 20.800 213.070 21.180 213.080 ;
        RECT 23.355 213.065 23.685 213.080 ;
        RECT 27.955 213.380 28.285 213.395 ;
        RECT 42.880 213.380 43.260 213.390 ;
        RECT 27.955 213.080 43.260 213.380 ;
        RECT 27.955 213.065 28.285 213.080 ;
        RECT 42.880 213.070 43.260 213.080 ;
        RECT 53.920 213.380 54.300 213.390 ;
        RECT 71.655 213.380 71.985 213.395 ;
        RECT 90.975 213.380 91.305 213.395 ;
        RECT 53.920 213.080 71.985 213.380 ;
        RECT 53.920 213.070 54.300 213.080 ;
        RECT 71.655 213.065 71.985 213.080 ;
        RECT 72.360 213.080 91.305 213.380 ;
        RECT 18.755 212.700 19.085 212.715 ;
        RECT 37.615 212.700 37.945 212.715 ;
        RECT 18.755 212.400 37.945 212.700 ;
        RECT 18.755 212.385 19.085 212.400 ;
        RECT 37.615 212.385 37.945 212.400 ;
        RECT 54.175 212.700 54.505 212.715 ;
        RECT 72.360 212.700 72.660 213.080 ;
        RECT 90.975 213.065 91.305 213.080 ;
        RECT 54.175 212.400 72.660 212.700 ;
        RECT 54.175 212.385 54.505 212.400 ;
        RECT 10.410 212.020 14.410 212.170 ;
        RECT 15.535 212.020 15.865 212.035 ;
        RECT 10.410 211.720 15.865 212.020 ;
        RECT 10.410 211.570 14.410 211.720 ;
        RECT 15.535 211.705 15.865 211.720 ;
        RECT 55.555 212.020 55.885 212.035 ;
        RECT 85.455 212.020 85.785 212.035 ;
        RECT 88.760 212.020 92.760 212.170 ;
        RECT 55.555 211.720 85.785 212.020 ;
        RECT 55.555 211.705 55.885 211.720 ;
        RECT 85.455 211.705 85.785 211.720 ;
        RECT 86.160 211.720 92.760 212.020 ;
        RECT 34.760 211.365 36.340 211.695 ;
        RECT 21.055 211.340 21.385 211.355 ;
        RECT 33.015 211.340 33.345 211.355 ;
        RECT 21.055 211.040 33.345 211.340 ;
        RECT 21.055 211.025 21.385 211.040 ;
        RECT 33.015 211.025 33.345 211.040 ;
        RECT 36.695 211.340 37.025 211.355 ;
        RECT 69.815 211.340 70.145 211.355 ;
        RECT 36.695 211.040 70.145 211.340 ;
        RECT 36.695 211.025 37.025 211.040 ;
        RECT 69.815 211.025 70.145 211.040 ;
        RECT 76.920 211.340 77.300 211.350 ;
        RECT 86.160 211.340 86.460 211.720 ;
        RECT 88.760 211.570 92.760 211.720 ;
        RECT 76.920 211.040 86.460 211.340 ;
        RECT 76.920 211.030 77.300 211.040 ;
        RECT 28.415 210.660 28.745 210.675 ;
        RECT 79.935 210.660 80.265 210.675 ;
        RECT 28.415 210.360 80.265 210.660 ;
        RECT 28.415 210.345 28.745 210.360 ;
        RECT 79.935 210.345 80.265 210.360 ;
        RECT 22.640 209.980 23.020 209.990 ;
        RECT 23.815 209.980 24.145 209.995 ;
        RECT 31.635 209.980 31.965 209.995 ;
        RECT 35.315 209.980 35.645 209.995 ;
        RECT 22.640 209.680 24.145 209.980 ;
        RECT 22.640 209.670 23.020 209.680 ;
        RECT 23.815 209.665 24.145 209.680 ;
        RECT 25.440 209.680 35.645 209.980 ;
        RECT 10.410 208.620 14.410 208.770 ;
        RECT 16.915 208.620 17.245 208.635 ;
        RECT 10.410 208.320 17.245 208.620 ;
        RECT 10.410 208.170 14.410 208.320 ;
        RECT 16.915 208.305 17.245 208.320 ;
        RECT 19.215 207.260 19.545 207.275 ;
        RECT 25.440 207.270 25.740 209.680 ;
        RECT 31.635 209.665 31.965 209.680 ;
        RECT 35.315 209.665 35.645 209.680 ;
        RECT 36.235 209.980 36.565 209.995 ;
        RECT 41.755 209.980 42.085 209.995 ;
        RECT 80.855 209.980 81.185 209.995 ;
        RECT 36.235 209.680 81.185 209.980 ;
        RECT 36.235 209.665 36.565 209.680 ;
        RECT 41.755 209.665 42.085 209.680 ;
        RECT 80.855 209.665 81.185 209.680 ;
        RECT 83.360 209.980 83.740 209.990 ;
        RECT 84.075 209.980 84.405 209.995 ;
        RECT 83.360 209.680 84.405 209.980 ;
        RECT 83.360 209.670 83.740 209.680 ;
        RECT 84.075 209.665 84.405 209.680 ;
        RECT 35.775 209.300 36.105 209.315 ;
        RECT 40.835 209.300 41.165 209.315 ;
        RECT 35.775 209.000 41.165 209.300 ;
        RECT 35.775 208.985 36.105 209.000 ;
        RECT 40.835 208.985 41.165 209.000 ;
        RECT 54.840 209.300 55.220 209.310 ;
        RECT 56.015 209.300 56.345 209.315 ;
        RECT 77.175 209.300 77.505 209.315 ;
        RECT 54.840 209.000 77.505 209.300 ;
        RECT 54.840 208.990 55.220 209.000 ;
        RECT 56.015 208.985 56.345 209.000 ;
        RECT 77.175 208.985 77.505 209.000 ;
        RECT 31.460 208.645 33.040 208.975 ;
        RECT 44.055 208.620 44.385 208.635 ;
        RECT 75.080 208.620 75.460 208.630 ;
        RECT 88.760 208.620 92.760 208.770 ;
        RECT 33.720 208.320 58.860 208.620 ;
        RECT 26.115 207.940 26.445 207.955 ;
        RECT 33.720 207.940 34.020 208.320 ;
        RECT 44.055 208.305 44.385 208.320 ;
        RECT 26.115 207.640 34.020 207.940 ;
        RECT 35.315 207.940 35.645 207.955 ;
        RECT 44.720 207.940 45.100 207.950 ;
        RECT 35.315 207.640 45.100 207.940 ;
        RECT 58.560 207.940 58.860 208.320 ;
        RECT 75.080 208.320 92.760 208.620 ;
        RECT 75.080 208.310 75.460 208.320 ;
        RECT 88.760 208.170 92.760 208.320 ;
        RECT 85.455 207.940 85.785 207.955 ;
        RECT 58.560 207.640 85.785 207.940 ;
        RECT 26.115 207.625 26.445 207.640 ;
        RECT 35.315 207.625 35.645 207.640 ;
        RECT 44.720 207.630 45.100 207.640 ;
        RECT 85.455 207.625 85.785 207.640 ;
        RECT 25.400 207.260 25.780 207.270 ;
        RECT 19.215 206.960 25.780 207.260 ;
        RECT 19.215 206.945 19.545 206.960 ;
        RECT 25.400 206.950 25.780 206.960 ;
        RECT 27.035 207.260 27.365 207.275 ;
        RECT 65.675 207.260 66.005 207.275 ;
        RECT 27.035 206.960 66.005 207.260 ;
        RECT 27.035 206.945 27.365 206.960 ;
        RECT 65.675 206.945 66.005 206.960 ;
        RECT 69.815 207.260 70.145 207.275 ;
        RECT 79.015 207.260 79.345 207.275 ;
        RECT 69.815 206.960 79.345 207.260 ;
        RECT 69.815 206.945 70.145 206.960 ;
        RECT 79.015 206.945 79.345 206.960 ;
        RECT 23.815 206.580 24.145 206.595 ;
        RECT 27.050 206.580 27.350 206.945 ;
        RECT 23.815 206.280 27.350 206.580 ;
        RECT 27.955 206.580 28.285 206.595 ;
        RECT 37.155 206.590 37.485 206.595 ;
        RECT 33.680 206.580 34.060 206.590 ;
        RECT 27.955 206.280 34.060 206.580 ;
        RECT 23.815 206.265 24.145 206.280 ;
        RECT 27.955 206.265 28.285 206.280 ;
        RECT 33.680 206.270 34.060 206.280 ;
        RECT 37.155 206.580 37.740 206.590 ;
        RECT 52.080 206.580 52.460 206.590 ;
        RECT 53.255 206.580 53.585 206.595 ;
        RECT 37.155 206.280 37.940 206.580 ;
        RECT 52.080 206.280 53.585 206.580 ;
        RECT 37.155 206.270 37.740 206.280 ;
        RECT 52.080 206.270 52.460 206.280 ;
        RECT 37.155 206.265 37.485 206.270 ;
        RECT 53.255 206.265 53.585 206.280 ;
        RECT 67.055 206.580 67.385 206.595 ;
        RECT 67.720 206.580 68.100 206.590 ;
        RECT 67.055 206.280 68.100 206.580 ;
        RECT 67.055 206.265 67.385 206.280 ;
        RECT 67.720 206.270 68.100 206.280 ;
        RECT 69.560 206.580 69.940 206.590 ;
        RECT 82.695 206.580 83.025 206.595 ;
        RECT 69.560 206.280 83.025 206.580 ;
        RECT 69.560 206.270 69.940 206.280 ;
        RECT 82.695 206.265 83.025 206.280 ;
        RECT 34.760 205.925 36.340 206.255 ;
        RECT 23.355 205.900 23.685 205.915 ;
        RECT 33.935 205.900 34.265 205.915 ;
        RECT 23.355 205.600 34.265 205.900 ;
        RECT 23.355 205.585 23.685 205.600 ;
        RECT 33.935 205.585 34.265 205.600 ;
        RECT 36.695 205.900 37.025 205.915 ;
        RECT 55.095 205.900 55.425 205.915 ;
        RECT 36.695 205.600 71.740 205.900 ;
        RECT 36.695 205.585 37.025 205.600 ;
        RECT 55.095 205.585 55.425 205.600 ;
        RECT 10.410 205.220 14.410 205.370 ;
        RECT 16.455 205.220 16.785 205.235 ;
        RECT 10.410 204.920 16.785 205.220 ;
        RECT 10.410 204.770 14.410 204.920 ;
        RECT 16.455 204.905 16.785 204.920 ;
        RECT 25.655 205.220 25.985 205.235 ;
        RECT 28.415 205.220 28.745 205.235 ;
        RECT 66.800 205.220 67.180 205.230 ;
        RECT 69.815 205.220 70.145 205.235 ;
        RECT 25.655 204.920 28.745 205.220 ;
        RECT 25.655 204.905 25.985 204.920 ;
        RECT 28.415 204.905 28.745 204.920 ;
        RECT 30.040 204.920 70.145 205.220 ;
        RECT 71.440 205.220 71.740 205.600 ;
        RECT 72.115 205.220 72.445 205.235 ;
        RECT 71.440 204.920 72.445 205.220 ;
        RECT 25.195 203.860 25.525 203.875 ;
        RECT 30.040 203.860 30.340 204.920 ;
        RECT 66.800 204.910 67.180 204.920 ;
        RECT 69.815 204.905 70.145 204.920 ;
        RECT 72.115 204.905 72.445 204.920 ;
        RECT 76.000 205.220 76.380 205.230 ;
        RECT 88.760 205.220 92.760 205.370 ;
        RECT 76.000 204.920 92.760 205.220 ;
        RECT 76.000 204.910 76.380 204.920 ;
        RECT 88.760 204.770 92.760 204.920 ;
        RECT 31.635 204.540 31.965 204.555 ;
        RECT 39.200 204.540 39.580 204.550 ;
        RECT 31.635 204.240 39.580 204.540 ;
        RECT 31.635 204.225 31.965 204.240 ;
        RECT 39.200 204.230 39.580 204.240 ;
        RECT 40.375 204.540 40.705 204.555 ;
        RECT 54.840 204.540 55.220 204.550 ;
        RECT 40.375 204.240 55.220 204.540 ;
        RECT 40.375 204.225 40.705 204.240 ;
        RECT 54.840 204.230 55.220 204.240 ;
        RECT 56.935 204.540 57.265 204.555 ;
        RECT 57.600 204.540 57.980 204.550 ;
        RECT 56.935 204.240 57.980 204.540 ;
        RECT 56.935 204.225 57.265 204.240 ;
        RECT 57.600 204.230 57.980 204.240 ;
        RECT 25.195 203.560 30.340 203.860 ;
        RECT 34.395 203.860 34.725 203.875 ;
        RECT 41.960 203.860 42.340 203.870 ;
        RECT 34.395 203.560 42.340 203.860 ;
        RECT 25.195 203.545 25.525 203.560 ;
        RECT 34.395 203.545 34.725 203.560 ;
        RECT 41.960 203.550 42.340 203.560 ;
        RECT 44.515 203.860 44.845 203.875 ;
        RECT 50.240 203.860 50.620 203.870 ;
        RECT 70.735 203.860 71.065 203.875 ;
        RECT 44.515 203.560 71.065 203.860 ;
        RECT 44.515 203.545 44.845 203.560 ;
        RECT 50.240 203.550 50.620 203.560 ;
        RECT 70.735 203.545 71.065 203.560 ;
        RECT 31.460 203.205 33.040 203.535 ;
        RECT 21.515 203.180 21.845 203.195 ;
        RECT 22.640 203.180 23.020 203.190 ;
        RECT 21.515 202.880 23.020 203.180 ;
        RECT 21.515 202.865 21.845 202.880 ;
        RECT 22.640 202.870 23.020 202.880 ;
        RECT 24.275 203.180 24.605 203.195 ;
        RECT 29.795 203.180 30.125 203.195 ;
        RECT 24.275 202.880 30.125 203.180 ;
        RECT 24.275 202.865 24.605 202.880 ;
        RECT 29.795 202.865 30.125 202.880 ;
        RECT 33.935 203.180 34.265 203.195 ;
        RECT 36.235 203.180 36.565 203.195 ;
        RECT 38.280 203.180 38.660 203.190 ;
        RECT 33.935 202.880 38.660 203.180 ;
        RECT 33.935 202.865 34.265 202.880 ;
        RECT 36.235 202.865 36.565 202.880 ;
        RECT 38.280 202.870 38.660 202.880 ;
        RECT 40.375 203.180 40.705 203.195 ;
        RECT 63.120 203.180 63.500 203.190 ;
        RECT 63.835 203.180 64.165 203.195 ;
        RECT 40.375 202.880 64.165 203.180 ;
        RECT 40.375 202.865 40.705 202.880 ;
        RECT 63.120 202.870 63.500 202.880 ;
        RECT 63.835 202.865 64.165 202.880 ;
        RECT 71.400 203.180 71.780 203.190 ;
        RECT 73.495 203.180 73.825 203.195 ;
        RECT 71.400 202.880 73.825 203.180 ;
        RECT 71.400 202.870 71.780 202.880 ;
        RECT 73.495 202.865 73.825 202.880 ;
        RECT 26.320 202.500 26.700 202.510 ;
        RECT 30.715 202.500 31.045 202.515 ;
        RECT 26.320 202.200 31.045 202.500 ;
        RECT 26.320 202.190 26.700 202.200 ;
        RECT 30.715 202.185 31.045 202.200 ;
        RECT 31.635 202.500 31.965 202.515 ;
        RECT 50.035 202.500 50.365 202.515 ;
        RECT 31.635 202.200 50.365 202.500 ;
        RECT 31.635 202.185 31.965 202.200 ;
        RECT 50.035 202.185 50.365 202.200 ;
        RECT 10.410 201.820 14.410 201.970 ;
        RECT 15.535 201.820 15.865 201.835 ;
        RECT 10.410 201.520 15.865 201.820 ;
        RECT 10.410 201.370 14.410 201.520 ;
        RECT 15.535 201.505 15.865 201.520 ;
        RECT 22.895 201.820 23.225 201.835 ;
        RECT 33.475 201.820 33.805 201.835 ;
        RECT 43.800 201.820 44.180 201.830 ;
        RECT 22.895 201.520 29.650 201.820 ;
        RECT 22.895 201.505 23.225 201.520 ;
        RECT 24.275 201.140 24.605 201.155 ;
        RECT 28.160 201.140 28.540 201.150 ;
        RECT 24.275 200.840 28.540 201.140 ;
        RECT 29.350 201.140 29.650 201.520 ;
        RECT 33.475 201.520 44.180 201.820 ;
        RECT 33.475 201.505 33.805 201.520 ;
        RECT 43.800 201.510 44.180 201.520 ;
        RECT 53.000 201.820 53.380 201.830 ;
        RECT 57.395 201.820 57.725 201.835 ;
        RECT 53.000 201.520 57.725 201.820 ;
        RECT 53.000 201.510 53.380 201.520 ;
        RECT 57.395 201.505 57.725 201.520 ;
        RECT 73.240 201.820 73.620 201.830 ;
        RECT 88.760 201.820 92.760 201.970 ;
        RECT 73.240 201.520 92.760 201.820 ;
        RECT 73.240 201.510 73.620 201.520 ;
        RECT 88.760 201.370 92.760 201.520 ;
        RECT 33.935 201.140 34.265 201.155 ;
        RECT 29.350 200.840 34.265 201.140 ;
        RECT 24.275 200.825 24.605 200.840 ;
        RECT 28.160 200.830 28.540 200.840 ;
        RECT 33.935 200.825 34.265 200.840 ;
        RECT 37.615 201.140 37.945 201.155 ;
        RECT 58.520 201.140 58.900 201.150 ;
        RECT 69.355 201.140 69.685 201.155 ;
        RECT 37.615 200.840 69.685 201.140 ;
        RECT 37.615 200.825 37.945 200.840 ;
        RECT 58.520 200.830 58.900 200.840 ;
        RECT 69.355 200.825 69.685 200.840 ;
        RECT 80.600 201.140 80.980 201.150 ;
        RECT 82.235 201.140 82.565 201.155 ;
        RECT 80.600 200.840 82.565 201.140 ;
        RECT 80.600 200.830 80.980 200.840 ;
        RECT 82.235 200.825 82.565 200.840 ;
        RECT 34.760 200.485 36.340 200.815 ;
        RECT 22.640 200.460 23.020 200.470 ;
        RECT 25.655 200.460 25.985 200.475 ;
        RECT 22.640 200.160 25.985 200.460 ;
        RECT 22.640 200.150 23.020 200.160 ;
        RECT 25.655 200.145 25.985 200.160 ;
        RECT 30.000 200.460 30.380 200.470 ;
        RECT 32.095 200.460 32.425 200.475 ;
        RECT 30.000 200.160 32.425 200.460 ;
        RECT 30.000 200.150 30.380 200.160 ;
        RECT 32.095 200.145 32.425 200.160 ;
        RECT 36.695 200.460 37.025 200.475 ;
        RECT 49.575 200.460 49.905 200.475 ;
        RECT 36.695 200.160 49.905 200.460 ;
        RECT 36.695 200.145 37.025 200.160 ;
        RECT 49.575 200.145 49.905 200.160 ;
        RECT 55.555 200.460 55.885 200.475 ;
        RECT 78.555 200.460 78.885 200.475 ;
        RECT 55.555 200.160 78.885 200.460 ;
        RECT 55.555 200.145 55.885 200.160 ;
        RECT 78.555 200.145 78.885 200.160 ;
        RECT 29.335 199.780 29.665 199.795 ;
        RECT 31.175 199.780 31.505 199.795 ;
        RECT 36.710 199.780 37.010 200.145 ;
        RECT 29.335 199.480 37.010 199.780 ;
        RECT 44.975 199.780 45.305 199.795 ;
        RECT 79.475 199.780 79.805 199.795 ;
        RECT 44.975 199.480 79.805 199.780 ;
        RECT 29.335 199.465 29.665 199.480 ;
        RECT 31.175 199.465 31.505 199.480 ;
        RECT 44.975 199.465 45.305 199.480 ;
        RECT 79.475 199.465 79.805 199.480 ;
        RECT 38.280 199.100 38.660 199.110 ;
        RECT 39.455 199.100 39.785 199.115 ;
        RECT 30.040 198.800 34.020 199.100 ;
        RECT 10.410 198.420 14.410 198.570 ;
        RECT 17.835 198.420 18.165 198.435 ;
        RECT 10.410 198.120 18.165 198.420 ;
        RECT 10.410 197.970 14.410 198.120 ;
        RECT 17.835 198.105 18.165 198.120 ;
        RECT 24.735 197.740 25.065 197.755 ;
        RECT 25.655 197.740 25.985 197.755 ;
        RECT 30.040 197.740 30.340 198.800 ;
        RECT 33.720 198.420 34.020 198.800 ;
        RECT 38.280 198.800 39.785 199.100 ;
        RECT 38.280 198.790 38.660 198.800 ;
        RECT 39.455 198.785 39.785 198.800 ;
        RECT 40.835 199.110 41.165 199.115 ;
        RECT 40.835 199.100 41.420 199.110 ;
        RECT 42.215 199.100 42.545 199.115 ;
        RECT 56.475 199.100 56.805 199.115 ;
        RECT 40.835 198.800 41.620 199.100 ;
        RECT 42.215 198.800 56.805 199.100 ;
        RECT 40.835 198.790 41.420 198.800 ;
        RECT 40.835 198.785 41.165 198.790 ;
        RECT 42.215 198.785 42.545 198.800 ;
        RECT 56.475 198.785 56.805 198.800 ;
        RECT 64.755 199.110 65.085 199.115 ;
        RECT 64.755 199.100 65.340 199.110 ;
        RECT 64.755 198.800 65.540 199.100 ;
        RECT 64.755 198.790 65.340 198.800 ;
        RECT 64.755 198.785 65.085 198.790 ;
        RECT 46.815 198.420 47.145 198.435 ;
        RECT 58.315 198.420 58.645 198.435 ;
        RECT 33.720 198.120 41.380 198.420 ;
        RECT 31.460 197.765 33.040 198.095 ;
        RECT 24.735 197.440 30.340 197.740 ;
        RECT 33.935 197.740 34.265 197.755 ;
        RECT 37.155 197.740 37.485 197.755 ;
        RECT 38.535 197.750 38.865 197.755 ;
        RECT 38.280 197.740 38.865 197.750 ;
        RECT 33.935 197.440 37.485 197.740 ;
        RECT 38.080 197.440 38.865 197.740 ;
        RECT 24.735 197.425 25.065 197.440 ;
        RECT 25.655 197.425 25.985 197.440 ;
        RECT 33.935 197.425 34.265 197.440 ;
        RECT 37.155 197.425 37.485 197.440 ;
        RECT 38.280 197.430 38.865 197.440 ;
        RECT 38.535 197.425 38.865 197.430 ;
        RECT 28.415 197.060 28.745 197.075 ;
        RECT 40.120 197.060 40.500 197.070 ;
        RECT 28.415 196.760 40.500 197.060 ;
        RECT 41.080 197.060 41.380 198.120 ;
        RECT 46.815 198.120 58.645 198.420 ;
        RECT 46.815 198.105 47.145 198.120 ;
        RECT 58.315 198.105 58.645 198.120 ;
        RECT 64.040 198.420 64.420 198.430 ;
        RECT 66.595 198.420 66.925 198.435 ;
        RECT 88.760 198.420 92.760 198.570 ;
        RECT 64.040 198.120 66.925 198.420 ;
        RECT 64.040 198.110 64.420 198.120 ;
        RECT 66.595 198.105 66.925 198.120 ;
        RECT 72.360 198.120 92.760 198.420 ;
        RECT 50.955 197.740 51.285 197.755 ;
        RECT 72.360 197.740 72.660 198.120 ;
        RECT 88.760 197.970 92.760 198.120 ;
        RECT 50.955 197.440 72.660 197.740 ;
        RECT 50.955 197.425 51.285 197.440 ;
        RECT 67.055 197.060 67.385 197.075 ;
        RECT 41.080 196.760 67.385 197.060 ;
        RECT 28.415 196.745 28.745 196.760 ;
        RECT 40.120 196.750 40.500 196.760 ;
        RECT 67.055 196.745 67.385 196.760 ;
        RECT 23.560 196.380 23.940 196.390 ;
        RECT 26.575 196.380 26.905 196.395 ;
        RECT 29.335 196.390 29.665 196.395 ;
        RECT 29.080 196.380 29.665 196.390 ;
        RECT 37.615 196.380 37.945 196.395 ;
        RECT 23.560 196.080 26.905 196.380 ;
        RECT 28.880 196.080 29.665 196.380 ;
        RECT 23.560 196.070 23.940 196.080 ;
        RECT 26.575 196.065 26.905 196.080 ;
        RECT 29.080 196.070 29.665 196.080 ;
        RECT 29.335 196.065 29.665 196.070 ;
        RECT 33.950 196.080 37.945 196.380 ;
        RECT 22.435 195.700 22.765 195.715 ;
        RECT 33.950 195.700 34.250 196.080 ;
        RECT 37.615 196.065 37.945 196.080 ;
        RECT 40.120 196.380 40.500 196.390 ;
        RECT 41.755 196.380 42.085 196.395 ;
        RECT 40.120 196.080 42.085 196.380 ;
        RECT 40.120 196.070 40.500 196.080 ;
        RECT 41.755 196.065 42.085 196.080 ;
        RECT 44.055 196.380 44.385 196.395 ;
        RECT 48.195 196.380 48.525 196.395 ;
        RECT 44.055 196.080 48.525 196.380 ;
        RECT 44.055 196.065 44.385 196.080 ;
        RECT 48.195 196.065 48.525 196.080 ;
        RECT 57.600 196.380 57.980 196.390 ;
        RECT 80.395 196.380 80.725 196.395 ;
        RECT 57.600 196.080 80.725 196.380 ;
        RECT 57.600 196.070 57.980 196.080 ;
        RECT 80.395 196.065 80.725 196.080 ;
        RECT 22.435 195.400 34.250 195.700 ;
        RECT 40.835 195.700 41.165 195.715 ;
        RECT 45.640 195.700 46.020 195.710 ;
        RECT 80.855 195.700 81.185 195.715 ;
        RECT 40.835 195.400 81.185 195.700 ;
        RECT 22.435 195.385 22.765 195.400 ;
        RECT 40.835 195.385 41.165 195.400 ;
        RECT 45.640 195.390 46.020 195.400 ;
        RECT 80.855 195.385 81.185 195.400 ;
        RECT 10.410 195.020 14.410 195.170 ;
        RECT 34.760 195.045 36.340 195.375 ;
        RECT 15.075 195.020 15.405 195.035 ;
        RECT 10.410 194.720 15.405 195.020 ;
        RECT 10.410 194.570 14.410 194.720 ;
        RECT 15.075 194.705 15.405 194.720 ;
        RECT 23.355 195.020 23.685 195.035 ;
        RECT 31.635 195.020 31.965 195.035 ;
        RECT 23.355 194.720 31.965 195.020 ;
        RECT 23.355 194.705 23.685 194.720 ;
        RECT 31.635 194.705 31.965 194.720 ;
        RECT 44.975 195.020 45.305 195.035 ;
        RECT 53.255 195.020 53.585 195.035 ;
        RECT 44.975 194.720 53.585 195.020 ;
        RECT 44.975 194.705 45.305 194.720 ;
        RECT 53.255 194.705 53.585 194.720 ;
        RECT 73.495 195.020 73.825 195.035 ;
        RECT 88.760 195.020 92.760 195.170 ;
        RECT 73.495 194.720 92.760 195.020 ;
        RECT 73.495 194.705 73.825 194.720 ;
        RECT 88.760 194.570 92.760 194.720 ;
        RECT 31.175 194.340 31.505 194.355 ;
        RECT 47.275 194.340 47.605 194.355 ;
        RECT 31.175 194.040 47.605 194.340 ;
        RECT 31.175 194.025 31.505 194.040 ;
        RECT 47.275 194.025 47.605 194.040 ;
        RECT 29.335 193.660 29.665 193.675 ;
        RECT 33.015 193.660 33.345 193.675 ;
        RECT 29.335 193.360 33.345 193.660 ;
        RECT 29.335 193.345 29.665 193.360 ;
        RECT 33.015 193.345 33.345 193.360 ;
        RECT 37.155 193.660 37.485 193.675 ;
        RECT 81.315 193.660 81.645 193.675 ;
        RECT 86.835 193.660 87.165 193.675 ;
        RECT 37.155 193.360 87.165 193.660 ;
        RECT 37.155 193.345 37.485 193.360 ;
        RECT 81.315 193.345 81.645 193.360 ;
        RECT 86.835 193.345 87.165 193.360 ;
        RECT 26.320 192.980 26.700 192.990 ;
        RECT 30.715 192.980 31.045 192.995 ;
        RECT 35.315 192.980 35.645 192.995 ;
        RECT 26.320 192.680 31.045 192.980 ;
        RECT 26.320 192.670 26.700 192.680 ;
        RECT 30.715 192.665 31.045 192.680 ;
        RECT 33.490 192.680 35.645 192.980 ;
        RECT 31.460 192.325 33.040 192.655 ;
        RECT 14.615 192.300 14.945 192.315 ;
        RECT 14.400 191.985 14.945 192.300 ;
        RECT 27.955 192.300 28.285 192.315 ;
        RECT 30.255 192.300 30.585 192.315 ;
        RECT 27.955 192.000 30.585 192.300 ;
        RECT 27.955 191.985 28.285 192.000 ;
        RECT 30.255 191.985 30.585 192.000 ;
        RECT 14.400 191.770 14.700 191.985 ;
        RECT 10.410 191.320 14.700 191.770 ;
        RECT 26.575 191.630 26.905 191.635 ;
        RECT 26.320 191.620 26.905 191.630 ;
        RECT 26.120 191.320 26.905 191.620 ;
        RECT 10.410 191.170 14.410 191.320 ;
        RECT 26.320 191.310 26.905 191.320 ;
        RECT 27.240 191.620 27.620 191.630 ;
        RECT 33.490 191.620 33.790 192.680 ;
        RECT 35.315 192.665 35.645 192.680 ;
        RECT 38.280 192.980 38.660 192.990 ;
        RECT 51.875 192.980 52.205 192.995 ;
        RECT 61.075 192.980 61.405 192.995 ;
        RECT 38.280 192.680 52.205 192.980 ;
        RECT 38.280 192.670 38.660 192.680 ;
        RECT 51.875 192.665 52.205 192.680 ;
        RECT 58.790 192.680 61.405 192.980 ;
        RECT 58.790 192.315 59.090 192.680 ;
        RECT 61.075 192.665 61.405 192.680 ;
        RECT 74.415 192.980 74.745 192.995 ;
        RECT 76.920 192.980 77.300 192.990 ;
        RECT 74.415 192.680 77.300 192.980 ;
        RECT 74.415 192.665 74.745 192.680 ;
        RECT 76.920 192.670 77.300 192.680 ;
        RECT 35.315 192.300 35.645 192.315 ;
        RECT 45.435 192.300 45.765 192.315 ;
        RECT 35.315 192.000 45.765 192.300 ;
        RECT 50.955 192.130 51.285 192.145 ;
        RECT 35.315 191.985 35.645 192.000 ;
        RECT 45.435 191.985 45.765 192.000 ;
        RECT 50.280 191.830 51.285 192.130 ;
        RECT 58.775 191.985 59.105 192.315 ;
        RECT 59.695 192.300 60.025 192.315 ;
        RECT 63.375 192.300 63.705 192.315 ;
        RECT 59.695 192.000 63.705 192.300 ;
        RECT 59.695 191.985 60.025 192.000 ;
        RECT 63.375 191.985 63.705 192.000 ;
        RECT 67.975 192.300 68.305 192.315 ;
        RECT 79.015 192.300 79.345 192.315 ;
        RECT 67.975 192.000 79.345 192.300 ;
        RECT 67.975 191.985 68.305 192.000 ;
        RECT 79.015 191.985 79.345 192.000 ;
        RECT 27.240 191.320 33.790 191.620 ;
        RECT 34.855 191.620 35.185 191.635 ;
        RECT 50.280 191.620 50.580 191.830 ;
        RECT 50.955 191.815 51.285 191.830 ;
        RECT 34.855 191.320 50.580 191.620 ;
        RECT 51.875 191.620 52.205 191.635 ;
        RECT 88.760 191.620 92.760 191.770 ;
        RECT 51.875 191.320 92.760 191.620 ;
        RECT 27.240 191.310 27.620 191.320 ;
        RECT 26.575 191.305 26.905 191.310 ;
        RECT 34.855 191.305 35.185 191.320 ;
        RECT 51.875 191.305 52.205 191.320 ;
        RECT 88.760 191.170 92.760 191.320 ;
        RECT 22.895 190.940 23.225 190.955 ;
        RECT 31.635 190.940 31.965 190.955 ;
        RECT 22.895 190.640 31.965 190.940 ;
        RECT 22.895 190.625 23.225 190.640 ;
        RECT 31.635 190.625 31.965 190.640 ;
        RECT 35.775 190.940 36.105 190.955 ;
        RECT 53.000 190.940 53.380 190.950 ;
        RECT 73.240 190.940 73.620 190.950 ;
        RECT 35.775 190.640 53.380 190.940 ;
        RECT 35.775 190.625 36.105 190.640 ;
        RECT 53.000 190.630 53.380 190.640 ;
        RECT 61.320 190.640 73.620 190.940 ;
        RECT 29.080 190.260 29.460 190.270 ;
        RECT 32.095 190.260 32.425 190.275 ;
        RECT 41.755 190.270 42.085 190.275 ;
        RECT 41.755 190.260 42.340 190.270 ;
        RECT 50.495 190.260 50.825 190.275 ;
        RECT 29.080 189.960 32.425 190.260 ;
        RECT 41.530 189.960 42.340 190.260 ;
        RECT 29.080 189.950 29.460 189.960 ;
        RECT 32.095 189.945 32.425 189.960 ;
        RECT 41.755 189.950 42.340 189.960 ;
        RECT 43.150 189.960 50.825 190.260 ;
        RECT 41.755 189.945 42.085 189.950 ;
        RECT 34.760 189.605 36.340 189.935 ;
        RECT 14.615 189.590 14.945 189.595 ;
        RECT 14.360 189.580 14.945 189.590 ;
        RECT 14.160 189.280 14.945 189.580 ;
        RECT 14.360 189.270 14.945 189.280 ;
        RECT 14.615 189.265 14.945 189.270 ;
        RECT 20.595 189.580 20.925 189.595 ;
        RECT 24.275 189.580 24.605 189.595 ;
        RECT 20.595 189.280 24.605 189.580 ;
        RECT 20.595 189.265 20.925 189.280 ;
        RECT 24.275 189.265 24.605 189.280 ;
        RECT 29.795 189.265 30.125 189.595 ;
        RECT 33.015 189.580 33.345 189.595 ;
        RECT 33.935 189.580 34.265 189.595 ;
        RECT 33.015 189.280 34.265 189.580 ;
        RECT 33.015 189.265 33.345 189.280 ;
        RECT 33.935 189.265 34.265 189.280 ;
        RECT 40.835 189.580 41.165 189.595 ;
        RECT 43.150 189.580 43.450 189.960 ;
        RECT 50.495 189.945 50.825 189.960 ;
        RECT 55.760 190.260 56.140 190.270 ;
        RECT 61.320 190.260 61.620 190.640 ;
        RECT 73.240 190.630 73.620 190.640 ;
        RECT 80.855 190.260 81.185 190.275 ;
        RECT 55.760 189.960 61.620 190.260 ;
        RECT 72.360 189.960 81.185 190.260 ;
        RECT 55.760 189.950 56.140 189.960 ;
        RECT 40.835 189.280 43.450 189.580 ;
        RECT 44.720 189.580 45.100 189.590 ;
        RECT 46.815 189.580 47.145 189.595 ;
        RECT 44.720 189.280 47.145 189.580 ;
        RECT 40.835 189.265 41.165 189.280 ;
        RECT 44.720 189.270 45.100 189.280 ;
        RECT 46.815 189.265 47.145 189.280 ;
        RECT 49.575 189.580 49.905 189.595 ;
        RECT 51.160 189.580 51.540 189.590 ;
        RECT 72.360 189.580 72.660 189.960 ;
        RECT 80.855 189.945 81.185 189.960 ;
        RECT 49.575 189.280 72.660 189.580 ;
        RECT 49.575 189.265 49.905 189.280 ;
        RECT 51.160 189.270 51.540 189.280 ;
        RECT 29.810 188.900 30.110 189.265 ;
        RECT 37.615 188.900 37.945 188.915 ;
        RECT 29.810 188.600 37.945 188.900 ;
        RECT 37.615 188.585 37.945 188.600 ;
        RECT 44.515 188.900 44.845 188.915 ;
        RECT 47.275 188.900 47.605 188.915 ;
        RECT 61.075 188.900 61.405 188.915 ;
        RECT 44.515 188.600 46.900 188.900 ;
        RECT 44.515 188.585 44.845 188.600 ;
        RECT 10.410 188.230 14.410 188.370 ;
        RECT 10.410 187.910 14.740 188.230 ;
        RECT 29.795 188.220 30.125 188.235 ;
        RECT 39.915 188.220 40.245 188.235 ;
        RECT 29.795 187.920 40.245 188.220 ;
        RECT 10.410 187.770 14.410 187.910 ;
        RECT 29.795 187.905 30.125 187.920 ;
        RECT 39.915 187.905 40.245 187.920 ;
        RECT 46.600 187.550 46.900 188.600 ;
        RECT 47.275 188.600 61.405 188.900 ;
        RECT 47.275 188.585 47.605 188.600 ;
        RECT 61.075 188.585 61.405 188.600 ;
        RECT 49.320 188.220 49.700 188.230 ;
        RECT 50.955 188.220 51.285 188.235 ;
        RECT 49.320 187.920 51.285 188.220 ;
        RECT 49.320 187.910 49.700 187.920 ;
        RECT 50.955 187.905 51.285 187.920 ;
        RECT 53.255 188.220 53.585 188.235 ;
        RECT 54.840 188.220 55.220 188.230 ;
        RECT 53.255 187.920 55.220 188.220 ;
        RECT 53.255 187.905 53.585 187.920 ;
        RECT 54.840 187.910 55.220 187.920 ;
        RECT 80.395 188.220 80.725 188.235 ;
        RECT 88.760 188.220 92.760 188.370 ;
        RECT 80.395 187.920 92.760 188.220 ;
        RECT 80.395 187.905 80.725 187.920 ;
        RECT 88.760 187.770 92.760 187.920 ;
        RECT 46.560 187.540 46.940 187.550 ;
        RECT 54.175 187.540 54.505 187.555 ;
        RECT 60.155 187.540 60.485 187.555 ;
        RECT 46.560 187.240 60.485 187.540 ;
        RECT 46.560 187.230 46.940 187.240 ;
        RECT 54.175 187.225 54.505 187.240 ;
        RECT 60.155 187.225 60.485 187.240 ;
        RECT 31.460 186.885 33.040 187.215 ;
        RECT 23.560 186.860 23.940 186.870 ;
        RECT 29.795 186.860 30.125 186.875 ;
        RECT 38.995 186.860 39.325 186.875 ;
        RECT 23.560 186.560 30.125 186.860 ;
        RECT 23.560 186.550 23.940 186.560 ;
        RECT 29.795 186.545 30.125 186.560 ;
        RECT 35.790 186.560 39.325 186.860 ;
        RECT 35.790 186.195 36.090 186.560 ;
        RECT 38.995 186.545 39.325 186.560 ;
        RECT 40.120 186.860 40.500 186.870 ;
        RECT 43.595 186.860 43.925 186.875 ;
        RECT 40.120 186.560 43.925 186.860 ;
        RECT 40.120 186.550 40.500 186.560 ;
        RECT 43.595 186.545 43.925 186.560 ;
        RECT 59.235 186.860 59.565 186.875 ;
        RECT 74.875 186.860 75.205 186.875 ;
        RECT 59.235 186.560 75.205 186.860 ;
        RECT 59.235 186.545 59.565 186.560 ;
        RECT 74.875 186.545 75.205 186.560 ;
        RECT 25.195 186.180 25.525 186.195 ;
        RECT 27.955 186.180 28.285 186.195 ;
        RECT 31.175 186.180 31.505 186.195 ;
        RECT 25.195 185.880 27.580 186.180 ;
        RECT 25.195 185.865 25.525 185.880 ;
        RECT 24.480 185.500 24.860 185.510 ;
        RECT 25.655 185.500 25.985 185.515 ;
        RECT 24.480 185.200 25.985 185.500 ;
        RECT 27.280 185.500 27.580 185.880 ;
        RECT 27.955 185.880 31.505 186.180 ;
        RECT 27.955 185.865 28.285 185.880 ;
        RECT 31.175 185.865 31.505 185.880 ;
        RECT 32.095 186.180 32.425 186.195 ;
        RECT 33.680 186.180 34.060 186.190 ;
        RECT 32.095 185.880 34.060 186.180 ;
        RECT 32.095 185.865 32.425 185.880 ;
        RECT 33.680 185.870 34.060 185.880 ;
        RECT 35.775 185.865 36.105 186.195 ;
        RECT 45.435 186.180 45.765 186.195 ;
        RECT 84.995 186.180 85.325 186.195 ;
        RECT 45.435 185.880 85.325 186.180 ;
        RECT 45.435 185.865 45.765 185.880 ;
        RECT 84.995 185.865 85.325 185.880 ;
        RECT 31.635 185.500 31.965 185.515 ;
        RECT 27.280 185.200 31.965 185.500 ;
        RECT 24.480 185.190 24.860 185.200 ;
        RECT 25.655 185.185 25.985 185.200 ;
        RECT 31.635 185.185 31.965 185.200 ;
        RECT 41.295 185.500 41.625 185.515 ;
        RECT 47.275 185.500 47.605 185.515 ;
        RECT 52.795 185.500 53.125 185.515 ;
        RECT 54.175 185.510 54.505 185.515 ;
        RECT 53.920 185.500 54.505 185.510 ;
        RECT 74.415 185.500 74.745 185.515 ;
        RECT 41.295 185.200 53.125 185.500 ;
        RECT 53.720 185.200 54.505 185.500 ;
        RECT 41.295 185.185 41.625 185.200 ;
        RECT 47.275 185.185 47.605 185.200 ;
        RECT 52.795 185.185 53.125 185.200 ;
        RECT 53.920 185.190 54.505 185.200 ;
        RECT 54.175 185.185 54.505 185.190 ;
        RECT 61.320 185.200 74.745 185.500 ;
        RECT 10.410 184.820 14.410 184.970 ;
        RECT 17.375 184.820 17.705 184.835 ;
        RECT 10.410 184.520 17.705 184.820 ;
        RECT 10.410 184.370 14.410 184.520 ;
        RECT 17.375 184.505 17.705 184.520 ;
        RECT 20.800 184.820 21.180 184.830 ;
        RECT 27.035 184.820 27.365 184.835 ;
        RECT 20.800 184.520 27.365 184.820 ;
        RECT 20.800 184.510 21.180 184.520 ;
        RECT 27.035 184.505 27.365 184.520 ;
        RECT 29.080 184.820 29.460 184.830 ;
        RECT 33.475 184.820 33.805 184.835 ;
        RECT 29.080 184.520 33.805 184.820 ;
        RECT 29.080 184.510 29.460 184.520 ;
        RECT 33.475 184.505 33.805 184.520 ;
        RECT 41.755 184.820 42.085 184.835 ;
        RECT 42.880 184.820 43.260 184.830 ;
        RECT 41.755 184.520 43.260 184.820 ;
        RECT 41.755 184.505 42.085 184.520 ;
        RECT 42.880 184.510 43.260 184.520 ;
        RECT 43.800 184.820 44.180 184.830 ;
        RECT 47.275 184.820 47.605 184.835 ;
        RECT 43.800 184.520 47.605 184.820 ;
        RECT 43.800 184.510 44.180 184.520 ;
        RECT 47.275 184.505 47.605 184.520 ;
        RECT 50.955 184.820 51.285 184.835 ;
        RECT 61.320 184.820 61.620 185.200 ;
        RECT 74.415 185.185 74.745 185.200 ;
        RECT 50.955 184.520 61.620 184.820 ;
        RECT 85.915 184.820 86.245 184.835 ;
        RECT 88.760 184.820 92.760 184.970 ;
        RECT 85.915 184.520 92.760 184.820 ;
        RECT 50.955 184.505 51.285 184.520 ;
        RECT 85.915 184.505 86.245 184.520 ;
        RECT 34.760 184.165 36.340 184.495 ;
        RECT 88.760 184.370 92.760 184.520 ;
        RECT 22.640 184.140 23.020 184.150 ;
        RECT 23.815 184.140 24.145 184.155 ;
        RECT 22.640 183.840 24.145 184.140 ;
        RECT 22.640 183.830 23.020 183.840 ;
        RECT 23.815 183.825 24.145 183.840 ;
        RECT 25.400 184.140 25.780 184.150 ;
        RECT 27.955 184.140 28.285 184.155 ;
        RECT 25.400 183.840 28.285 184.140 ;
        RECT 25.400 183.830 25.780 183.840 ;
        RECT 27.955 183.825 28.285 183.840 ;
        RECT 30.255 184.140 30.585 184.155 ;
        RECT 33.680 184.140 34.060 184.150 ;
        RECT 30.255 183.840 34.060 184.140 ;
        RECT 30.255 183.825 30.585 183.840 ;
        RECT 33.680 183.830 34.060 183.840 ;
        RECT 42.675 184.140 43.005 184.155 ;
        RECT 56.015 184.140 56.345 184.155 ;
        RECT 42.675 183.840 56.345 184.140 ;
        RECT 42.675 183.825 43.005 183.840 ;
        RECT 56.015 183.825 56.345 183.840 ;
        RECT 64.960 184.140 65.340 184.150 ;
        RECT 73.240 184.140 73.620 184.150 ;
        RECT 64.960 183.840 73.620 184.140 ;
        RECT 64.960 183.830 65.340 183.840 ;
        RECT 73.240 183.830 73.620 183.840 ;
        RECT 20.595 183.460 20.925 183.475 ;
        RECT 52.080 183.460 52.460 183.470 ;
        RECT 20.595 183.160 52.460 183.460 ;
        RECT 20.595 183.145 20.925 183.160 ;
        RECT 52.080 183.150 52.460 183.160 ;
        RECT 59.235 183.460 59.565 183.475 ;
        RECT 61.280 183.460 61.660 183.470 ;
        RECT 62.455 183.460 62.785 183.475 ;
        RECT 59.235 183.160 62.785 183.460 ;
        RECT 59.235 183.145 59.565 183.160 ;
        RECT 61.280 183.150 61.660 183.160 ;
        RECT 62.455 183.145 62.785 183.160 ;
        RECT 67.055 183.460 67.385 183.475 ;
        RECT 69.560 183.460 69.940 183.470 ;
        RECT 67.055 183.160 69.940 183.460 ;
        RECT 67.055 183.145 67.385 183.160 ;
        RECT 69.560 183.150 69.940 183.160 ;
        RECT 13.695 182.780 14.025 182.795 ;
        RECT 25.655 182.780 25.985 182.795 ;
        RECT 13.695 182.480 25.985 182.780 ;
        RECT 13.695 182.465 14.025 182.480 ;
        RECT 25.655 182.465 25.985 182.480 ;
        RECT 26.320 182.780 26.700 182.790 ;
        RECT 29.795 182.780 30.125 182.795 ;
        RECT 26.320 182.480 30.125 182.780 ;
        RECT 26.320 182.470 26.700 182.480 ;
        RECT 29.795 182.465 30.125 182.480 ;
        RECT 30.715 182.780 31.045 182.795 ;
        RECT 40.375 182.780 40.705 182.795 ;
        RECT 30.715 182.480 40.705 182.780 ;
        RECT 30.715 182.465 31.045 182.480 ;
        RECT 40.375 182.465 40.705 182.480 ;
        RECT 42.215 182.780 42.545 182.795 ;
        RECT 47.275 182.780 47.605 182.795 ;
        RECT 42.215 182.480 47.605 182.780 ;
        RECT 42.215 182.465 42.545 182.480 ;
        RECT 47.275 182.465 47.605 182.480 ;
        RECT 52.795 182.780 53.125 182.795 ;
        RECT 53.715 182.780 54.045 182.795 ;
        RECT 52.795 182.480 54.045 182.780 ;
        RECT 52.795 182.465 53.125 182.480 ;
        RECT 53.715 182.465 54.045 182.480 ;
        RECT 25.655 182.100 25.985 182.115 ;
        RECT 27.240 182.100 27.620 182.110 ;
        RECT 25.655 181.800 27.620 182.100 ;
        RECT 25.655 181.785 25.985 181.800 ;
        RECT 27.240 181.790 27.620 181.800 ;
        RECT 33.680 182.100 34.060 182.110 ;
        RECT 47.735 182.100 48.065 182.115 ;
        RECT 50.495 182.110 50.825 182.115 ;
        RECT 33.680 181.800 48.065 182.100 ;
        RECT 33.680 181.790 34.060 181.800 ;
        RECT 47.735 181.785 48.065 181.800 ;
        RECT 50.240 182.100 50.825 182.110 ;
        RECT 50.240 181.800 51.050 182.100 ;
        RECT 50.240 181.790 50.825 181.800 ;
        RECT 50.495 181.785 50.825 181.790 ;
        RECT 31.460 181.445 33.040 181.775 ;
        RECT 35.315 181.420 35.645 181.435 ;
        RECT 36.695 181.420 37.025 181.435 ;
        RECT 38.995 181.420 39.325 181.435 ;
        RECT 47.735 181.420 48.065 181.435 ;
        RECT 35.315 181.120 48.065 181.420 ;
        RECT 35.315 181.105 35.645 181.120 ;
        RECT 36.695 181.105 37.025 181.120 ;
        RECT 38.995 181.105 39.325 181.120 ;
        RECT 47.735 181.105 48.065 181.120 ;
        RECT 53.715 181.420 54.045 181.435 ;
        RECT 59.235 181.420 59.565 181.435 ;
        RECT 53.715 181.120 59.565 181.420 ;
        RECT 53.715 181.105 54.045 181.120 ;
        RECT 59.235 181.105 59.565 181.120 ;
        RECT 85.455 181.420 85.785 181.435 ;
        RECT 88.760 181.420 92.760 181.570 ;
        RECT 85.455 181.120 92.760 181.420 ;
        RECT 85.455 181.105 85.785 181.120 ;
        RECT 88.760 180.970 92.760 181.120 ;
        RECT 38.280 180.740 38.660 180.750 ;
        RECT 39.915 180.740 40.245 180.755 ;
        RECT 46.355 180.740 46.685 180.755 ;
        RECT 38.280 180.440 46.685 180.740 ;
        RECT 38.280 180.430 38.660 180.440 ;
        RECT 39.915 180.425 40.245 180.440 ;
        RECT 46.355 180.425 46.685 180.440 ;
        RECT 53.715 180.740 54.045 180.755 ;
        RECT 57.600 180.740 57.980 180.750 ;
        RECT 53.715 180.440 57.980 180.740 ;
        RECT 53.715 180.425 54.045 180.440 ;
        RECT 57.600 180.430 57.980 180.440 ;
        RECT 58.775 180.740 59.105 180.755 ;
        RECT 69.355 180.740 69.685 180.755 ;
        RECT 58.775 180.440 69.685 180.740 ;
        RECT 58.775 180.425 59.105 180.440 ;
        RECT 69.355 180.425 69.685 180.440 ;
        RECT 26.115 180.060 26.445 180.075 ;
        RECT 39.200 180.060 39.580 180.070 ;
        RECT 26.115 179.760 39.580 180.060 ;
        RECT 26.115 179.745 26.445 179.760 ;
        RECT 39.200 179.750 39.580 179.760 ;
        RECT 40.835 180.060 41.165 180.075 ;
        RECT 50.955 180.060 51.285 180.075 ;
        RECT 40.835 179.760 51.285 180.060 ;
        RECT 40.835 179.745 41.165 179.760 ;
        RECT 50.955 179.745 51.285 179.760 ;
        RECT 56.475 180.060 56.805 180.075 ;
        RECT 63.835 180.060 64.165 180.075 ;
        RECT 56.475 179.760 64.165 180.060 ;
        RECT 56.475 179.745 56.805 179.760 ;
        RECT 63.835 179.745 64.165 179.760 ;
        RECT 64.960 180.060 65.340 180.070 ;
        RECT 87.755 180.060 88.085 180.075 ;
        RECT 64.960 179.760 88.085 180.060 ;
        RECT 64.960 179.750 65.340 179.760 ;
        RECT 87.755 179.745 88.085 179.760 ;
        RECT 46.815 179.380 47.145 179.395 ;
        RECT 53.000 179.380 53.380 179.390 ;
        RECT 54.840 179.380 55.220 179.390 ;
        RECT 68.640 179.380 69.020 179.390 ;
        RECT 46.815 179.080 69.020 179.380 ;
        RECT 46.815 179.065 47.145 179.080 ;
        RECT 53.000 179.070 53.380 179.080 ;
        RECT 54.840 179.070 55.220 179.080 ;
        RECT 68.640 179.070 69.020 179.080 ;
        RECT 34.760 178.725 36.340 179.055 ;
        RECT 36.695 178.700 37.025 178.715 ;
        RECT 46.355 178.700 46.685 178.715 ;
        RECT 48.655 178.710 48.985 178.715 ;
        RECT 48.400 178.700 48.985 178.710 ;
        RECT 50.955 178.710 51.285 178.715 ;
        RECT 50.955 178.700 51.540 178.710 ;
        RECT 36.695 178.400 46.685 178.700 ;
        RECT 48.200 178.400 48.985 178.700 ;
        RECT 50.730 178.400 51.540 178.700 ;
        RECT 36.695 178.385 37.025 178.400 ;
        RECT 46.355 178.385 46.685 178.400 ;
        RECT 48.400 178.390 48.985 178.400 ;
        RECT 48.655 178.385 48.985 178.390 ;
        RECT 50.955 178.390 51.540 178.400 ;
        RECT 51.875 178.700 52.205 178.715 ;
        RECT 53.920 178.700 54.300 178.710 ;
        RECT 56.475 178.700 56.805 178.715 ;
        RECT 51.875 178.400 56.805 178.700 ;
        RECT 50.955 178.385 51.285 178.390 ;
        RECT 51.875 178.385 52.205 178.400 ;
        RECT 53.920 178.390 54.300 178.400 ;
        RECT 56.475 178.385 56.805 178.400 ;
        RECT 58.315 178.385 58.645 178.715 ;
        RECT 66.135 178.700 66.465 178.715 ;
        RECT 76.000 178.700 76.380 178.710 ;
        RECT 66.135 178.400 76.380 178.700 ;
        RECT 66.135 178.385 66.465 178.400 ;
        RECT 76.000 178.390 76.380 178.400 ;
        RECT 10.410 178.020 14.410 178.170 ;
        RECT 58.330 178.035 58.630 178.385 ;
        RECT 17.375 178.020 17.705 178.035 ;
        RECT 10.410 177.720 17.705 178.020 ;
        RECT 10.410 177.570 14.410 177.720 ;
        RECT 17.375 177.705 17.705 177.720 ;
        RECT 38.535 178.020 38.865 178.035 ;
        RECT 44.975 178.020 45.305 178.035 ;
        RECT 38.535 177.720 45.305 178.020 ;
        RECT 38.535 177.705 38.865 177.720 ;
        RECT 44.975 177.705 45.305 177.720 ;
        RECT 45.640 178.020 46.020 178.030 ;
        RECT 51.875 178.020 52.205 178.035 ;
        RECT 45.640 177.720 52.205 178.020 ;
        RECT 45.640 177.710 46.020 177.720 ;
        RECT 51.875 177.705 52.205 177.720 ;
        RECT 56.475 178.030 56.805 178.035 ;
        RECT 56.475 178.020 57.060 178.030 ;
        RECT 56.475 177.720 57.260 178.020 ;
        RECT 56.475 177.710 57.060 177.720 ;
        RECT 56.475 177.705 56.805 177.710 ;
        RECT 58.315 177.705 58.645 178.035 ;
        RECT 65.675 178.020 66.005 178.035 ;
        RECT 67.515 178.030 67.845 178.035 ;
        RECT 66.800 178.020 67.180 178.030 ;
        RECT 65.675 177.720 67.180 178.020 ;
        RECT 65.675 177.705 66.005 177.720 ;
        RECT 66.800 177.710 67.180 177.720 ;
        RECT 67.515 178.020 68.100 178.030 ;
        RECT 84.995 178.020 85.325 178.035 ;
        RECT 88.760 178.020 92.760 178.170 ;
        RECT 67.515 177.720 68.300 178.020 ;
        RECT 84.995 177.720 92.760 178.020 ;
        RECT 67.515 177.710 68.100 177.720 ;
        RECT 67.515 177.705 67.845 177.710 ;
        RECT 84.995 177.705 85.325 177.720 ;
        RECT 88.760 177.570 92.760 177.720 ;
        RECT 30.000 177.340 30.380 177.350 ;
        RECT 41.040 177.340 41.420 177.350 ;
        RECT 48.195 177.340 48.525 177.355 ;
        RECT 30.000 177.040 40.690 177.340 ;
        RECT 30.000 177.030 30.380 177.040 ;
        RECT 40.390 176.660 40.690 177.040 ;
        RECT 41.040 177.040 48.525 177.340 ;
        RECT 41.040 177.030 41.420 177.040 ;
        RECT 48.195 177.025 48.525 177.040 ;
        RECT 50.955 177.340 51.285 177.355 ;
        RECT 55.760 177.340 56.140 177.350 ;
        RECT 50.955 177.040 56.140 177.340 ;
        RECT 50.955 177.025 51.285 177.040 ;
        RECT 55.760 177.030 56.140 177.040 ;
        RECT 57.395 177.340 57.725 177.355 ;
        RECT 75.795 177.340 76.125 177.355 ;
        RECT 57.395 177.040 76.125 177.340 ;
        RECT 57.395 177.025 57.725 177.040 ;
        RECT 75.795 177.025 76.125 177.040 ;
        RECT 48.655 176.660 48.985 176.675 ;
        RECT 76.715 176.660 77.045 176.675 ;
        RECT 40.390 176.360 48.985 176.660 ;
        RECT 48.655 176.345 48.985 176.360 ;
        RECT 63.160 176.360 77.045 176.660 ;
        RECT 31.460 176.005 33.040 176.335 ;
        RECT 37.360 175.980 37.740 175.990 ;
        RECT 59.695 175.980 60.025 175.995 ;
        RECT 37.360 175.680 60.025 175.980 ;
        RECT 37.360 175.670 37.740 175.680 ;
        RECT 59.695 175.665 60.025 175.680 ;
        RECT 28.160 175.300 28.540 175.310 ;
        RECT 47.275 175.300 47.605 175.315 ;
        RECT 62.455 175.300 62.785 175.315 ;
        RECT 28.160 175.000 62.785 175.300 ;
        RECT 28.160 174.990 28.540 175.000 ;
        RECT 47.275 174.985 47.605 175.000 ;
        RECT 62.455 174.985 62.785 175.000 ;
        RECT 16.200 174.620 16.580 174.630 ;
        RECT 51.415 174.620 51.745 174.635 ;
        RECT 55.095 174.630 55.425 174.635 ;
        RECT 16.200 174.320 51.745 174.620 ;
        RECT 16.200 174.310 16.580 174.320 ;
        RECT 51.415 174.305 51.745 174.320 ;
        RECT 54.840 174.620 55.425 174.630 ;
        RECT 56.015 174.620 56.345 174.635 ;
        RECT 61.075 174.630 61.405 174.635 ;
        RECT 58.520 174.620 58.900 174.630 ;
        RECT 54.840 174.320 55.650 174.620 ;
        RECT 56.015 174.320 58.900 174.620 ;
        RECT 54.840 174.310 55.425 174.320 ;
        RECT 55.095 174.305 55.425 174.310 ;
        RECT 56.015 174.305 56.345 174.320 ;
        RECT 58.520 174.310 58.900 174.320 ;
        RECT 61.075 174.620 61.660 174.630 ;
        RECT 61.075 174.320 61.860 174.620 ;
        RECT 61.075 174.310 61.660 174.320 ;
        RECT 61.075 174.305 61.405 174.310 ;
        RECT 46.355 173.950 46.685 173.955 ;
        RECT 49.115 173.950 49.445 173.955 ;
        RECT 54.175 173.950 54.505 173.955 ;
        RECT 46.355 173.940 46.940 173.950 ;
        RECT 49.115 173.940 49.700 173.950 ;
        RECT 53.920 173.940 54.505 173.950 ;
        RECT 46.130 173.640 46.940 173.940 ;
        RECT 48.890 173.640 49.700 173.940 ;
        RECT 53.720 173.640 54.505 173.940 ;
        RECT 46.355 173.630 46.940 173.640 ;
        RECT 49.115 173.630 49.700 173.640 ;
        RECT 53.920 173.630 54.505 173.640 ;
        RECT 46.355 173.625 46.685 173.630 ;
        RECT 49.115 173.625 49.445 173.630 ;
        RECT 54.175 173.625 54.505 173.630 ;
        RECT 57.855 173.940 58.185 173.955 ;
        RECT 63.160 173.940 63.460 176.360 ;
        RECT 76.715 176.345 77.045 176.360 ;
        RECT 80.855 175.980 81.185 175.995 ;
        RECT 72.360 175.680 81.185 175.980 ;
        RECT 64.295 174.620 64.625 174.635 ;
        RECT 64.960 174.620 65.340 174.630 ;
        RECT 72.360 174.620 72.660 175.680 ;
        RECT 80.855 175.665 81.185 175.680 ;
        RECT 76.255 175.300 76.585 175.315 ;
        RECT 79.935 175.300 80.265 175.315 ;
        RECT 80.600 175.300 80.980 175.310 ;
        RECT 76.255 175.000 80.980 175.300 ;
        RECT 76.255 174.985 76.585 175.000 ;
        RECT 79.935 174.985 80.265 175.000 ;
        RECT 80.600 174.990 80.980 175.000 ;
        RECT 64.295 174.320 65.340 174.620 ;
        RECT 64.295 174.305 64.625 174.320 ;
        RECT 64.960 174.310 65.340 174.320 ;
        RECT 66.840 174.320 72.660 174.620 ;
        RECT 84.995 174.620 85.325 174.635 ;
        RECT 88.760 174.620 92.760 174.770 ;
        RECT 84.995 174.320 92.760 174.620 ;
        RECT 57.855 173.640 63.460 173.940 ;
        RECT 64.040 173.940 64.420 173.950 ;
        RECT 65.675 173.940 66.005 173.955 ;
        RECT 64.040 173.640 66.005 173.940 ;
        RECT 57.855 173.625 58.185 173.640 ;
        RECT 64.040 173.630 64.420 173.640 ;
        RECT 65.675 173.625 66.005 173.640 ;
        RECT 34.760 173.285 36.340 173.615 ;
        RECT 42.880 173.260 43.260 173.270 ;
        RECT 44.975 173.260 45.305 173.275 ;
        RECT 48.655 173.270 48.985 173.275 ;
        RECT 42.880 172.960 45.305 173.260 ;
        RECT 42.880 172.950 43.260 172.960 ;
        RECT 44.975 172.945 45.305 172.960 ;
        RECT 48.400 173.260 48.985 173.270 ;
        RECT 49.575 173.260 49.905 173.275 ;
        RECT 51.415 173.260 51.745 173.275 ;
        RECT 48.400 172.960 49.210 173.260 ;
        RECT 49.575 172.960 51.745 173.260 ;
        RECT 48.400 172.950 48.985 172.960 ;
        RECT 48.655 172.945 48.985 172.950 ;
        RECT 49.575 172.945 49.905 172.960 ;
        RECT 51.415 172.945 51.745 172.960 ;
        RECT 63.120 173.260 63.500 173.270 ;
        RECT 64.755 173.260 65.085 173.275 ;
        RECT 63.120 172.960 65.085 173.260 ;
        RECT 63.120 172.950 63.500 172.960 ;
        RECT 64.755 172.945 65.085 172.960 ;
        RECT 30.255 172.580 30.585 172.595 ;
        RECT 37.155 172.580 37.485 172.595 ;
        RECT 30.255 172.280 37.485 172.580 ;
        RECT 30.255 172.265 30.585 172.280 ;
        RECT 37.155 172.265 37.485 172.280 ;
        RECT 44.515 172.580 44.845 172.595 ;
        RECT 49.575 172.580 49.905 172.595 ;
        RECT 44.515 172.280 49.905 172.580 ;
        RECT 44.515 172.265 44.845 172.280 ;
        RECT 49.575 172.265 49.905 172.280 ;
        RECT 60.155 172.580 60.485 172.595 ;
        RECT 62.915 172.580 63.245 172.595 ;
        RECT 66.840 172.580 67.140 174.320 ;
        RECT 84.995 174.305 85.325 174.320 ;
        RECT 88.760 174.170 92.760 174.320 ;
        RECT 67.975 173.940 68.305 173.955 ;
        RECT 69.560 173.940 69.940 173.950 ;
        RECT 67.975 173.640 69.940 173.940 ;
        RECT 67.975 173.625 68.305 173.640 ;
        RECT 69.560 173.630 69.940 173.640 ;
        RECT 68.640 173.260 69.020 173.270 ;
        RECT 83.155 173.260 83.485 173.275 ;
        RECT 68.640 172.960 83.485 173.260 ;
        RECT 68.640 172.950 69.020 172.960 ;
        RECT 83.155 172.945 83.485 172.960 ;
        RECT 60.155 172.280 67.140 172.580 ;
        RECT 69.815 172.580 70.145 172.595 ;
        RECT 77.175 172.580 77.505 172.595 ;
        RECT 69.815 172.280 77.505 172.580 ;
        RECT 60.155 172.265 60.485 172.280 ;
        RECT 62.915 172.265 63.245 172.280 ;
        RECT 69.815 172.265 70.145 172.280 ;
        RECT 77.175 172.265 77.505 172.280 ;
        RECT 18.295 171.900 18.625 171.915 ;
        RECT 74.875 171.900 75.205 171.915 ;
        RECT 18.295 171.600 75.205 171.900 ;
        RECT 18.295 171.585 18.625 171.600 ;
        RECT 74.875 171.585 75.205 171.600 ;
        RECT 44.975 171.220 45.305 171.235 ;
        RECT 52.795 171.220 53.125 171.235 ;
        RECT 44.975 170.920 53.125 171.220 ;
        RECT 44.975 170.905 45.305 170.920 ;
        RECT 52.795 170.905 53.125 170.920 ;
        RECT 63.375 171.220 63.705 171.235 ;
        RECT 67.055 171.220 67.385 171.235 ;
        RECT 63.375 170.920 67.385 171.220 ;
        RECT 63.375 170.905 63.705 170.920 ;
        RECT 67.055 170.905 67.385 170.920 ;
        RECT 75.795 171.220 76.125 171.235 ;
        RECT 88.760 171.220 92.760 171.370 ;
        RECT 75.795 170.920 92.760 171.220 ;
        RECT 75.795 170.905 76.125 170.920 ;
        RECT 31.460 170.565 33.040 170.895 ;
        RECT 88.760 170.770 92.760 170.920 ;
        RECT 60.615 170.540 60.945 170.555 ;
        RECT 74.415 170.540 74.745 170.555 ;
        RECT 60.615 170.240 74.745 170.540 ;
        RECT 60.615 170.225 60.945 170.240 ;
        RECT 74.415 170.225 74.745 170.240 ;
        RECT 28.875 169.860 29.205 169.875 ;
        RECT 40.375 169.860 40.705 169.875 ;
        RECT 28.875 169.560 40.705 169.860 ;
        RECT 28.875 169.545 29.205 169.560 ;
        RECT 40.375 169.545 40.705 169.560 ;
        RECT 64.755 169.860 65.085 169.875 ;
        RECT 77.175 169.860 77.505 169.875 ;
        RECT 64.755 169.560 77.505 169.860 ;
        RECT 64.755 169.545 65.085 169.560 ;
        RECT 77.175 169.545 77.505 169.560 ;
        RECT 35.315 169.180 35.645 169.195 ;
        RECT 36.695 169.180 37.025 169.195 ;
        RECT 44.975 169.180 45.305 169.195 ;
        RECT 35.315 168.880 45.305 169.180 ;
        RECT 35.315 168.865 35.645 168.880 ;
        RECT 36.695 168.865 37.025 168.880 ;
        RECT 44.975 168.865 45.305 168.880 ;
        RECT 34.760 167.845 36.340 168.175 ;
        RECT 81.775 167.820 82.105 167.835 ;
        RECT 88.760 167.820 92.760 167.970 ;
        RECT 81.775 167.520 92.760 167.820 ;
        RECT 81.775 167.505 82.105 167.520 ;
        RECT 88.760 167.370 92.760 167.520 ;
        RECT 25.195 167.140 25.525 167.155 ;
        RECT 30.255 167.140 30.585 167.155 ;
        RECT 68.895 167.140 69.225 167.155 ;
        RECT 73.035 167.140 73.365 167.155 ;
        RECT 25.195 166.840 73.365 167.140 ;
        RECT 25.195 166.825 25.525 166.840 ;
        RECT 30.255 166.825 30.585 166.840 ;
        RECT 68.895 166.825 69.225 166.840 ;
        RECT 73.035 166.825 73.365 166.840 ;
        RECT 69.815 166.460 70.145 166.475 ;
        RECT 71.400 166.460 71.780 166.470 ;
        RECT 69.815 166.160 71.780 166.460 ;
        RECT 69.815 166.145 70.145 166.160 ;
        RECT 71.400 166.150 71.780 166.160 ;
        RECT 31.460 165.125 33.040 165.455 ;
        RECT 73.240 164.420 73.620 164.430 ;
        RECT 73.955 164.420 74.285 164.435 ;
        RECT 73.240 164.120 74.285 164.420 ;
        RECT 73.240 164.110 73.620 164.120 ;
        RECT 73.955 164.105 74.285 164.120 ;
        RECT 82.235 164.420 82.565 164.435 ;
        RECT 88.760 164.420 92.760 164.570 ;
        RECT 82.235 164.120 92.760 164.420 ;
        RECT 82.235 164.105 82.565 164.120 ;
        RECT 88.760 163.970 92.760 164.120 ;
        RECT 74.875 163.750 75.205 163.755 ;
        RECT 74.875 163.740 75.460 163.750 ;
        RECT 74.650 163.440 75.460 163.740 ;
        RECT 74.875 163.430 75.460 163.440 ;
        RECT 74.875 163.425 75.205 163.430 ;
        RECT 34.760 162.405 36.340 162.735 ;
        RECT 45.895 161.700 46.225 161.715 ;
        RECT 47.735 161.700 48.065 161.715 ;
        RECT 45.895 161.400 48.065 161.700 ;
        RECT 45.895 161.385 46.225 161.400 ;
        RECT 47.735 161.385 48.065 161.400 ;
        RECT 10.410 161.020 14.410 161.170 ;
        RECT 17.835 161.020 18.165 161.035 ;
        RECT 10.410 160.720 18.165 161.020 ;
        RECT 10.410 160.570 14.410 160.720 ;
        RECT 17.835 160.705 18.165 160.720 ;
        RECT 41.295 161.020 41.625 161.035 ;
        RECT 45.895 161.020 46.225 161.035 ;
        RECT 41.295 160.720 46.225 161.020 ;
        RECT 41.295 160.705 41.625 160.720 ;
        RECT 45.895 160.705 46.225 160.720 ;
        RECT 78.095 161.020 78.425 161.035 ;
        RECT 88.760 161.020 92.760 161.170 ;
        RECT 78.095 160.720 92.760 161.020 ;
        RECT 78.095 160.705 78.425 160.720 ;
        RECT 88.760 160.570 92.760 160.720 ;
        RECT 31.460 159.685 33.040 160.015 ;
        RECT 44.975 159.660 45.305 159.675 ;
        RECT 47.735 159.660 48.065 159.675 ;
        RECT 44.975 159.360 48.065 159.660 ;
        RECT 44.975 159.345 45.305 159.360 ;
        RECT 47.735 159.345 48.065 159.360 ;
        RECT 10.410 157.620 14.410 157.770 ;
        RECT 19.675 157.620 20.005 157.635 ;
        RECT 10.410 157.320 20.005 157.620 ;
        RECT 10.410 157.170 14.410 157.320 ;
        RECT 19.675 157.305 20.005 157.320 ;
        RECT 83.615 157.620 83.945 157.635 ;
        RECT 88.760 157.620 92.760 157.770 ;
        RECT 83.615 157.320 92.760 157.620 ;
        RECT 83.615 157.305 83.945 157.320 ;
        RECT 34.760 156.965 36.340 157.295 ;
        RECT 88.760 157.170 92.760 157.320 ;
        RECT 17.375 154.900 17.705 154.915 ;
        RECT 14.400 154.600 17.705 154.900 ;
        RECT 14.400 154.370 14.700 154.600 ;
        RECT 17.375 154.585 17.705 154.600 ;
        RECT 10.410 153.920 14.700 154.370 ;
        RECT 31.460 154.245 33.040 154.575 ;
        RECT 80.395 154.220 80.725 154.235 ;
        RECT 88.760 154.220 92.760 154.370 ;
        RECT 80.395 153.920 92.760 154.220 ;
        RECT 10.410 153.770 14.410 153.920 ;
        RECT 80.395 153.905 80.725 153.920 ;
        RECT 88.760 153.770 92.760 153.920 ;
        RECT 38.535 152.860 38.865 152.875 ;
        RECT 79.475 152.860 79.805 152.875 ;
        RECT 38.535 152.560 79.805 152.860 ;
        RECT 38.535 152.545 38.865 152.560 ;
        RECT 79.475 152.545 79.805 152.560 ;
        RECT 34.760 151.525 36.340 151.855 ;
        RECT 10.410 150.820 14.410 150.970 ;
        RECT 85.455 150.820 85.785 150.835 ;
        RECT 88.760 150.820 92.760 150.970 ;
        RECT 10.410 150.370 14.700 150.820 ;
        RECT 85.455 150.520 92.760 150.820 ;
        RECT 85.455 150.505 85.785 150.520 ;
        RECT 88.760 150.370 92.760 150.520 ;
        RECT 14.400 150.140 14.700 150.370 ;
        RECT 17.835 150.140 18.165 150.155 ;
        RECT 14.400 149.840 18.165 150.140 ;
        RECT 17.835 149.825 18.165 149.840 ;
        RECT 31.460 148.805 33.040 149.135 ;
        RECT 84.995 147.420 85.325 147.435 ;
        RECT 88.760 147.420 92.760 147.570 ;
        RECT 84.995 147.120 92.760 147.420 ;
        RECT 84.995 147.105 85.325 147.120 ;
        RECT 88.760 146.970 92.760 147.120 ;
        RECT 34.760 146.085 36.340 146.415 ;
        RECT 85.455 144.020 85.785 144.035 ;
        RECT 88.760 144.020 92.760 144.170 ;
        RECT 85.455 143.720 92.760 144.020 ;
        RECT 85.455 143.705 85.785 143.720 ;
        RECT 31.460 143.365 33.040 143.695 ;
        RECT 88.760 143.570 92.760 143.720 ;
        RECT 34.760 140.645 36.340 140.975 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 29.105 221.905 29.435 222.235 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 16.225 217.825 16.555 218.155 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 14.385 189.265 14.715 189.595 ;
        RECT 14.400 188.235 14.700 189.265 ;
        RECT 14.385 187.905 14.715 188.235 ;
        RECT 16.240 174.635 16.540 217.825 ;
        RECT 24.505 215.785 24.835 216.115 ;
        RECT 20.825 213.065 21.155 213.395 ;
        RECT 20.840 184.835 21.140 213.065 ;
        RECT 22.240 209.240 23.420 210.420 ;
        RECT 22.240 202.440 23.420 203.620 ;
        RECT 22.665 200.145 22.995 200.475 ;
        RECT 20.825 184.505 21.155 184.835 ;
        RECT 22.680 184.155 22.980 200.145 ;
        RECT 23.585 196.065 23.915 196.395 ;
        RECT 23.600 186.875 23.900 196.065 ;
        RECT 23.585 186.545 23.915 186.875 ;
        RECT 24.520 185.515 24.820 215.785 ;
        RECT 25.425 206.945 25.755 207.275 ;
        RECT 24.505 185.185 24.835 185.515 ;
        RECT 25.440 184.155 25.740 206.945 ;
        RECT 26.345 202.185 26.675 202.515 ;
        RECT 26.360 192.995 26.660 202.185 ;
        RECT 28.185 200.825 28.515 201.155 ;
        RECT 28.200 193.420 28.500 200.825 ;
        RECT 29.120 196.395 29.420 221.905 ;
        RECT 40.145 215.105 40.475 215.435 ;
        RECT 30.025 200.145 30.355 200.475 ;
        RECT 29.105 196.065 29.435 196.395 ;
        RECT 26.345 192.665 26.675 192.995 ;
        RECT 27.760 192.240 28.940 193.420 ;
        RECT 26.345 191.305 26.675 191.635 ;
        RECT 27.265 191.305 27.595 191.635 ;
        RECT 22.665 183.825 22.995 184.155 ;
        RECT 25.425 183.825 25.755 184.155 ;
        RECT 26.360 182.795 26.660 191.305 ;
        RECT 26.345 182.465 26.675 182.795 ;
        RECT 27.280 182.115 27.580 191.305 ;
        RECT 27.265 181.785 27.595 182.115 ;
        RECT 28.200 175.315 28.500 192.240 ;
        RECT 29.105 189.945 29.435 190.275 ;
        RECT 29.120 184.835 29.420 189.945 ;
        RECT 29.105 184.505 29.435 184.835 ;
        RECT 30.040 177.355 30.340 200.145 ;
        RECT 30.025 177.025 30.355 177.355 ;
        RECT 28.185 174.985 28.515 175.315 ;
        RECT 16.225 174.305 16.555 174.635 ;
        RECT 31.450 140.570 33.050 211.770 ;
        RECT 33.705 206.265 34.035 206.595 ;
        RECT 33.720 186.195 34.020 206.265 ;
        RECT 33.705 185.865 34.035 186.195 ;
        RECT 33.705 183.825 34.035 184.155 ;
        RECT 33.720 182.115 34.020 183.825 ;
        RECT 33.705 181.785 34.035 182.115 ;
        RECT 34.750 140.570 36.350 211.770 ;
        RECT 37.385 206.265 37.715 206.595 ;
        RECT 37.400 175.995 37.700 206.265 ;
        RECT 39.225 204.225 39.555 204.555 ;
        RECT 38.305 202.865 38.635 203.195 ;
        RECT 38.320 199.115 38.620 202.865 ;
        RECT 38.305 198.785 38.635 199.115 ;
        RECT 38.305 197.425 38.635 197.755 ;
        RECT 38.320 192.995 38.620 197.425 ;
        RECT 38.305 192.665 38.635 192.995 ;
        RECT 38.320 180.755 38.620 192.665 ;
        RECT 38.305 180.425 38.635 180.755 ;
        RECT 39.240 180.075 39.540 204.225 ;
        RECT 40.160 197.075 40.460 215.105 ;
        RECT 56.705 213.745 57.035 214.075 ;
        RECT 42.905 213.065 43.235 213.395 ;
        RECT 53.945 213.065 54.275 213.395 ;
        RECT 41.985 203.545 42.315 203.875 ;
        RECT 41.065 198.785 41.395 199.115 ;
        RECT 40.145 196.745 40.475 197.075 ;
        RECT 40.145 196.065 40.475 196.395 ;
        RECT 40.160 186.875 40.460 196.065 ;
        RECT 40.145 186.545 40.475 186.875 ;
        RECT 39.225 179.745 39.555 180.075 ;
        RECT 41.080 177.355 41.380 198.785 ;
        RECT 42.000 190.275 42.300 203.545 ;
        RECT 41.985 189.945 42.315 190.275 ;
        RECT 42.920 184.835 43.220 213.065 ;
        RECT 44.745 207.625 45.075 207.955 ;
        RECT 43.825 201.505 44.155 201.835 ;
        RECT 43.840 184.835 44.140 201.505 ;
        RECT 44.760 189.595 45.060 207.625 ;
        RECT 52.105 206.265 52.435 206.595 ;
        RECT 50.265 203.545 50.595 203.875 ;
        RECT 45.665 195.385 45.995 195.715 ;
        RECT 44.745 189.265 45.075 189.595 ;
        RECT 42.905 184.505 43.235 184.835 ;
        RECT 43.825 184.505 44.155 184.835 ;
        RECT 41.065 177.025 41.395 177.355 ;
        RECT 37.385 175.665 37.715 175.995 ;
        RECT 42.920 173.275 43.220 184.505 ;
        RECT 45.680 178.035 45.980 195.385 ;
        RECT 49.345 187.905 49.675 188.235 ;
        RECT 46.585 187.225 46.915 187.555 ;
        RECT 45.665 177.705 45.995 178.035 ;
        RECT 46.600 173.955 46.900 187.225 ;
        RECT 48.425 178.385 48.755 178.715 ;
        RECT 46.585 173.625 46.915 173.955 ;
        RECT 48.440 173.275 48.740 178.385 ;
        RECT 49.360 173.955 49.660 187.905 ;
        RECT 50.280 182.115 50.580 203.545 ;
        RECT 51.185 189.265 51.515 189.595 ;
        RECT 50.265 181.785 50.595 182.115 ;
        RECT 51.200 178.715 51.500 189.265 ;
        RECT 52.120 183.475 52.420 206.265 ;
        RECT 53.025 201.505 53.355 201.835 ;
        RECT 53.040 190.955 53.340 201.505 ;
        RECT 53.025 190.625 53.355 190.955 ;
        RECT 52.105 183.145 52.435 183.475 ;
        RECT 53.040 179.395 53.340 190.625 ;
        RECT 53.960 185.515 54.260 213.065 ;
        RECT 54.865 208.985 55.195 209.315 ;
        RECT 54.880 204.555 55.180 208.985 ;
        RECT 54.865 204.225 55.195 204.555 ;
        RECT 54.880 188.235 55.180 204.225 ;
        RECT 55.785 189.945 56.115 190.275 ;
        RECT 54.865 187.905 55.195 188.235 ;
        RECT 53.945 185.185 54.275 185.515 ;
        RECT 53.025 179.065 53.355 179.395 ;
        RECT 54.865 179.065 55.195 179.395 ;
        RECT 51.185 178.385 51.515 178.715 ;
        RECT 53.945 178.385 54.275 178.715 ;
        RECT 53.960 173.955 54.260 178.385 ;
        RECT 54.880 174.635 55.180 179.065 ;
        RECT 55.800 177.355 56.100 189.945 ;
        RECT 56.720 178.035 57.020 213.745 ;
        RECT 76.945 211.025 77.275 211.355 ;
        RECT 75.105 208.305 75.435 208.635 ;
        RECT 67.745 206.265 68.075 206.595 ;
        RECT 69.585 206.265 69.915 206.595 ;
        RECT 66.825 204.905 67.155 205.235 ;
        RECT 57.625 204.225 57.955 204.555 ;
        RECT 57.640 196.395 57.940 204.225 ;
        RECT 63.145 202.865 63.475 203.195 ;
        RECT 58.545 200.825 58.875 201.155 ;
        RECT 57.625 196.065 57.955 196.395 ;
        RECT 57.640 180.755 57.940 196.065 ;
        RECT 57.625 180.425 57.955 180.755 ;
        RECT 56.705 177.705 57.035 178.035 ;
        RECT 55.785 177.025 56.115 177.355 ;
        RECT 58.560 174.635 58.860 200.825 ;
        RECT 61.305 183.145 61.635 183.475 ;
        RECT 61.320 174.635 61.620 183.145 ;
        RECT 54.865 174.305 55.195 174.635 ;
        RECT 58.545 174.305 58.875 174.635 ;
        RECT 61.305 174.305 61.635 174.635 ;
        RECT 49.345 173.625 49.675 173.955 ;
        RECT 53.945 173.625 54.275 173.955 ;
        RECT 63.160 173.275 63.460 202.865 ;
        RECT 64.985 198.785 65.315 199.115 ;
        RECT 64.065 198.105 64.395 198.435 ;
        RECT 64.080 173.955 64.380 198.105 ;
        RECT 65.000 184.155 65.300 198.785 ;
        RECT 64.985 183.825 65.315 184.155 ;
        RECT 64.985 179.745 65.315 180.075 ;
        RECT 65.000 174.635 65.300 179.745 ;
        RECT 66.840 178.035 67.140 204.905 ;
        RECT 67.760 178.035 68.060 206.265 ;
        RECT 69.600 193.420 69.900 206.265 ;
        RECT 71.000 202.440 72.180 203.620 ;
        RECT 69.160 192.240 70.340 193.420 ;
        RECT 69.585 183.145 69.915 183.475 ;
        RECT 68.665 179.065 68.995 179.395 ;
        RECT 66.825 177.705 67.155 178.035 ;
        RECT 67.745 177.705 68.075 178.035 ;
        RECT 64.985 174.305 65.315 174.635 ;
        RECT 64.065 173.625 64.395 173.955 ;
        RECT 68.680 173.275 68.980 179.065 ;
        RECT 69.600 173.955 69.900 183.145 ;
        RECT 69.585 173.625 69.915 173.955 ;
        RECT 42.905 172.945 43.235 173.275 ;
        RECT 48.425 172.945 48.755 173.275 ;
        RECT 63.145 172.945 63.475 173.275 ;
        RECT 68.665 172.945 68.995 173.275 ;
        RECT 71.440 166.475 71.740 202.440 ;
        RECT 73.265 201.505 73.595 201.835 ;
        RECT 73.280 190.955 73.580 201.505 ;
        RECT 73.265 190.625 73.595 190.955 ;
        RECT 73.265 183.825 73.595 184.155 ;
        RECT 71.425 166.145 71.755 166.475 ;
        RECT 73.280 164.435 73.580 183.825 ;
        RECT 73.265 164.105 73.595 164.435 ;
        RECT 75.120 163.755 75.420 208.305 ;
        RECT 76.025 204.905 76.355 205.235 ;
        RECT 76.040 178.715 76.340 204.905 ;
        RECT 76.960 192.995 77.260 211.025 ;
        RECT 82.960 209.240 84.140 210.420 ;
        RECT 80.625 200.825 80.955 201.155 ;
        RECT 76.945 192.665 77.275 192.995 ;
        RECT 76.025 178.385 76.355 178.715 ;
        RECT 80.640 175.315 80.940 200.825 ;
        RECT 80.625 174.985 80.955 175.315 ;
        RECT 75.105 163.425 75.435 163.755 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
      LAYER met5 ;
        RECT 22.030 209.030 84.350 210.630 ;
        RECT 22.030 202.230 72.390 203.830 ;
        RECT 27.550 192.030 70.550 193.630 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

