magic
tech sky130A
magscale 1 2
timestamp 1757965599
<< locali >>
rect 29958 10332 30413 10462
<< metal1 >>
rect 2293 44822 2299 44874
rect 2351 44868 2357 44874
rect 17724 44868 17730 44874
rect 2351 44828 17730 44868
rect 2351 44822 2357 44828
rect 17724 44822 17730 44828
rect 17782 44822 17788 44874
rect 2376 44724 2382 44776
rect 2434 44774 2440 44776
rect 16072 44774 16078 44776
rect 2434 44726 16078 44774
rect 2434 44724 2440 44726
rect 16072 44724 16078 44726
rect 16130 44724 16136 44776
rect 15516 44604 15522 44656
rect 15574 44604 15580 44656
rect 7728 44564 7816 44578
rect 7728 44512 7748 44564
rect 7800 44552 7816 44564
rect 14968 44552 14974 44564
rect 7800 44524 14974 44552
rect 7800 44512 7816 44524
rect 14968 44512 14974 44524
rect 15026 44512 15032 44564
rect 7728 44498 7816 44512
rect 2496 44368 2502 44420
rect 2554 44418 2560 44420
rect 17174 44418 17180 44421
rect 2554 44371 17180 44418
rect 2554 44368 2560 44371
rect 17174 44369 17180 44371
rect 17232 44369 17238 44421
rect 21587 44084 21593 44139
rect 21648 44084 25457 44139
rect 25512 44084 25518 44139
rect 23784 43743 23790 43816
rect 23863 43743 26457 43816
rect 26530 43743 26536 43816
rect 24314 43695 24396 43710
rect 24314 43641 24327 43695
rect 24381 43641 26589 43695
rect 26643 43641 26649 43695
rect 24314 43624 24396 43641
rect 24889 43536 26713 43575
rect 24874 43519 26713 43536
rect 24874 43457 24889 43519
rect 24951 43513 26713 43519
rect 26775 43513 26781 43575
rect 24951 43457 24968 43513
rect 24874 43436 24968 43457
rect 23229 43403 23307 43409
rect 26790 43394 26850 43400
rect 23307 43334 26790 43394
rect 26790 43328 26850 43334
rect 23229 43319 23307 43325
rect 22690 43230 22696 43290
rect 22756 43230 26910 43290
rect 26970 43230 26976 43290
rect 17401 33662 17407 33717
rect 17462 33662 25570 33717
rect 25625 33662 25631 33717
rect 2495 33466 2501 33518
rect 2553 33515 2559 33518
rect 10963 33515 10969 33517
rect 2553 33468 10969 33515
rect 2553 33466 2559 33468
rect 10963 33465 10969 33468
rect 11021 33465 11027 33517
rect 15468 33496 15474 33552
rect 15530 33496 26232 33552
rect 26288 33496 26294 33552
rect 2376 33374 2382 33426
rect 2434 33424 2440 33426
rect 6178 33424 6184 33426
rect 2434 33376 6184 33424
rect 2434 33374 2440 33376
rect 6178 33374 6184 33376
rect 6236 33374 6242 33426
rect 14172 33340 14178 33413
rect 14251 33340 26333 33413
rect 26406 33340 26412 33413
rect 2293 33271 2299 33323
rect 2351 33321 2357 33323
rect 5811 33321 5817 33322
rect 2351 33272 5817 33321
rect 2351 33271 2357 33272
rect 5811 33270 5817 33272
rect 5869 33270 5875 33322
rect 26471 33291 26525 33297
rect 13537 33237 13543 33291
rect 13597 33237 26471 33291
rect 26471 33231 26525 33237
rect 2147 33175 2153 33227
rect 2205 33223 2211 33227
rect 5167 33223 5173 33226
rect 2205 33178 5173 33223
rect 2205 33175 2211 33178
rect 5167 33174 5173 33178
rect 5225 33174 5231 33226
rect 12251 33191 12313 33197
rect 12313 33129 26565 33191
rect 26627 33129 26633 33191
rect 12251 33123 12313 33129
rect 200 26788 4666 27116
rect 194 26388 200 26788
rect 600 26716 4666 26788
rect 600 26388 606 26716
rect 24684 16644 26414 16724
rect 1860 14724 1866 14776
rect 1918 14724 1924 14776
rect 1873 14088 1911 14724
rect 3448 14420 3666 14472
rect 3718 14420 3724 14472
rect 2156 14088 2229 14094
rect 1868 14015 2156 14088
rect 2156 14009 2229 14015
rect 3448 13580 3500 14420
rect 3540 14268 3546 14328
rect 3606 14268 3612 14328
rect 3546 13694 3606 14268
rect 24684 13705 24764 16644
rect 3546 13628 3606 13634
rect 3440 13524 3446 13580
rect 3502 13524 3508 13580
rect 23500 13512 24924 13705
rect 24731 13284 24924 13512
rect 29235 13302 30479 13397
rect 29235 13211 29330 13302
rect 23863 12033 23869 12233
rect 24000 12033 24006 12233
rect 25828 12199 25959 12205
rect 25828 12062 25959 12068
rect 26490 12019 26670 12025
rect 16676 11844 16772 11850
rect 11700 11815 11820 11838
rect 11700 11742 11724 11815
rect 11797 11742 11820 11815
rect 11700 11726 11820 11742
rect 21700 11846 21772 11852
rect 16676 11742 16772 11748
rect 18491 11743 18563 11817
rect 20133 11769 20221 11843
rect 21772 11774 21852 11846
rect 21700 11768 21772 11774
rect 23331 11749 23403 11839
rect 26490 11833 26670 11839
rect 30384 11627 30479 13302
rect 30036 11334 30096 11340
rect 30036 11268 30096 11274
rect 30350 11010 30410 11016
rect 30410 10950 30464 11010
rect 30350 10944 30410 10950
rect 3238 10822 3244 10874
rect 3296 10862 3302 10874
rect 10554 10862 10560 10874
rect 3296 10834 10560 10862
rect 3296 10822 3302 10834
rect 10554 10822 10560 10834
rect 10612 10822 10618 10874
rect 24335 10785 24831 10911
rect 31983 10882 31989 11082
rect 32073 10882 32079 11082
rect 3125 10715 3131 10781
rect 3197 10715 16861 10781
rect 16927 10715 16933 10781
rect 30183 10659 30333 10665
rect 17170 10625 17176 10626
rect 3004 10573 3010 10625
rect 3062 10574 17176 10625
rect 17228 10574 17234 10626
rect 3062 10573 3068 10574
rect 17564 10514 17628 10520
rect 2854 10450 2860 10514
rect 2924 10450 17564 10514
rect 17564 10444 17628 10450
rect 30183 10403 30333 10509
rect 29951 10253 30403 10403
rect 587 9933 683 9990
rect 497 9837 503 9933
rect 768 9837 774 9933
rect 948 7045 1101 7051
rect 1486 7017 1584 7159
rect 1101 6919 1584 7017
rect 948 6886 1101 6892
rect 199 6653 205 6806
rect 595 6653 806 6806
rect 935 3839 1073 3845
rect 1486 3819 1584 3953
rect 1073 3721 1584 3819
rect 935 3695 1073 3701
rect 200 3458 206 3594
rect 594 3458 754 3594
rect 318 616 417 803
rect 912 616 918 637
rect 318 517 918 616
rect 912 497 918 517
rect 1058 497 1064 637
<< via1 >>
rect 2299 44822 2351 44874
rect 17730 44822 17782 44874
rect 2382 44724 2434 44776
rect 16078 44724 16130 44776
rect 15522 44604 15574 44656
rect 7748 44512 7800 44564
rect 14974 44512 15026 44564
rect 2502 44368 2554 44420
rect 17180 44369 17232 44421
rect 21593 44084 21648 44139
rect 25457 44084 25512 44139
rect 23790 43743 23863 43816
rect 26457 43743 26530 43816
rect 24327 43641 24381 43695
rect 26589 43641 26643 43695
rect 24889 43457 24951 43519
rect 26713 43513 26775 43575
rect 23229 43325 23307 43403
rect 26790 43334 26850 43394
rect 22696 43230 22756 43290
rect 26910 43230 26970 43290
rect 17407 33662 17462 33717
rect 25570 33662 25625 33717
rect 2501 33466 2553 33518
rect 10969 33465 11021 33517
rect 15474 33496 15530 33552
rect 26232 33496 26288 33552
rect 2382 33374 2434 33426
rect 6184 33374 6236 33426
rect 14178 33340 14251 33413
rect 26333 33340 26406 33413
rect 2299 33271 2351 33323
rect 5817 33270 5869 33322
rect 13543 33237 13597 33291
rect 26471 33237 26525 33291
rect 2153 33175 2205 33227
rect 5173 33174 5225 33226
rect 12251 33129 12313 33191
rect 26565 33129 26627 33191
rect 200 26388 600 26788
rect 1866 14724 1918 14776
rect 3666 14420 3718 14472
rect 2156 14015 2229 14088
rect 3546 14268 3606 14328
rect 3546 13634 3606 13694
rect 3446 13524 3502 13580
rect 23869 12033 24000 12233
rect 25828 12068 25959 12199
rect 11724 11742 11797 11815
rect 13382 11750 13442 11810
rect 15087 11739 15149 11801
rect 16676 11748 16772 11844
rect 18417 11743 18491 11817
rect 20059 11769 20133 11843
rect 21700 11774 21772 11846
rect 26490 11839 26670 12019
rect 23403 11749 23493 11839
rect 30036 11274 30096 11334
rect 30350 10950 30410 11010
rect 3244 10822 3296 10874
rect 10560 10822 10612 10874
rect 31989 10882 32073 11082
rect 3131 10715 3197 10781
rect 16861 10715 16927 10781
rect 3010 10573 3062 10625
rect 17176 10574 17228 10626
rect 2860 10450 2924 10514
rect 17564 10450 17628 10514
rect 30183 10509 30333 10659
rect 503 9837 768 9933
rect 948 6892 1101 7045
rect 205 6653 595 6806
rect 935 3701 1073 3839
rect 206 3458 594 3594
rect 918 497 1058 637
<< metal2 >>
rect 14970 45068 15030 45077
rect 14970 44999 15030 45008
rect 15518 45076 15578 45085
rect 15518 45007 15578 45016
rect 16074 45054 16134 45063
rect 2299 44874 2351 44880
rect 2149 44830 2209 44839
rect 2299 44816 2351 44822
rect 2149 44761 2209 44770
rect 1281 38587 1371 38588
rect 1273 38579 1379 38587
rect 1273 38489 1281 38579
rect 1371 38489 1379 38579
rect 1273 38407 1379 38489
rect 200 26788 600 26794
rect 196 26393 200 26783
rect 600 26393 604 26783
rect 200 26382 600 26388
rect 1294 11770 1358 38407
rect 1423 37904 1513 37908
rect 1418 37899 1518 37904
rect 1418 37809 1423 37899
rect 1513 37809 1518 37899
rect 1418 37684 1518 37809
rect 1443 11882 1494 37684
rect 1559 37225 1649 37228
rect 1554 37219 1655 37225
rect 1554 37129 1559 37219
rect 1649 37129 1655 37219
rect 1554 37062 1655 37129
rect 1571 12029 1637 37062
rect 1744 35793 1844 35798
rect 1740 35703 1749 35793
rect 1839 35703 1848 35793
rect 1744 35632 1844 35703
rect 1750 34690 1839 35632
rect 1750 34218 1814 34690
rect 1864 34418 1920 34425
rect 1862 34416 1922 34418
rect 1862 34360 1864 34416
rect 1920 34360 1922 34416
rect 1862 34262 1922 34360
rect 1750 14846 1839 34218
rect 1750 14668 1822 14846
rect 1873 14782 1911 34262
rect 1866 14776 1918 14782
rect 1866 14718 1918 14724
rect 1750 13851 1839 14668
rect 1964 14532 1992 31566
rect 1750 13753 1839 13762
rect 1930 14406 1992 14532
rect 1930 13450 1990 14406
rect 1930 13394 1932 13450
rect 1988 13394 1990 13450
rect 1930 13392 1990 13394
rect 1932 13385 1988 13392
rect 2056 12104 2084 36786
rect 2156 36386 2202 44761
rect 2305 36407 2345 44816
rect 2382 44776 2434 44782
rect 2382 44718 2434 44724
rect 2164 36164 2195 36386
rect 2157 33233 2202 36164
rect 2310 36156 2341 36407
rect 2301 33329 2350 36156
rect 2384 33432 2432 44718
rect 7728 44564 7816 44578
rect 14986 44570 15014 44999
rect 15534 44662 15562 45007
rect 16074 44985 16134 44994
rect 17726 45046 17786 45055
rect 16080 44782 16128 44985
rect 17726 44977 17786 44986
rect 17736 44880 17776 44977
rect 17730 44874 17782 44880
rect 17730 44816 17782 44822
rect 26326 44834 26422 44843
rect 22545 44785 22627 44794
rect 16078 44776 16130 44782
rect 16078 44718 16130 44724
rect 18683 44679 18761 44731
rect 15522 44656 15574 44662
rect 15522 44598 15574 44604
rect 18683 44592 18761 44601
rect 7728 44512 7748 44564
rect 7800 44512 7816 44564
rect 7728 44498 7816 44512
rect 14974 44564 15026 44570
rect 14974 44506 15026 44512
rect 19329 44530 19404 44742
rect 20608 44655 20617 44729
rect 20691 44655 20700 44729
rect 17170 44488 17243 44497
rect 2502 44420 2554 44426
rect 2502 44362 2554 44368
rect 19329 44446 19404 44455
rect 21261 44457 21335 44715
rect 21905 44625 21979 44709
rect 22545 44651 22627 44703
rect 26326 44650 26422 44738
rect 21905 44542 21979 44551
rect 17170 44369 17180 44415
rect 17232 44369 17243 44415
rect 21261 44374 21335 44383
rect 2504 33524 2551 44362
rect 17170 44359 17243 44369
rect 21580 44310 21661 44319
rect 10964 44212 11046 44272
rect 11106 44212 11115 44272
rect 21580 44175 21661 44229
rect 25861 44283 25936 44292
rect 26037 44211 26101 44301
rect 26191 44211 26200 44301
rect 21593 44139 21648 44175
rect 25861 44157 25936 44208
rect 21593 44078 21648 44084
rect 25457 44139 25512 44145
rect 4810 44046 4870 44055
rect 4810 43977 4870 43986
rect 2592 43858 2652 43867
rect 2592 43789 2652 43798
rect 2595 43755 2649 43789
rect 2608 35284 2636 43755
rect 2714 43700 2774 43709
rect 2714 43631 2774 43640
rect 2716 33680 2772 43631
rect 4810 42627 4869 43977
rect 25457 43873 25512 44084
rect 25572 44100 25644 44110
rect 25572 43940 25644 44028
rect 23770 43816 23882 43836
rect 25457 43818 25548 43873
rect 23770 43743 23790 43816
rect 23863 43743 23882 43816
rect 23770 43724 23882 43743
rect 24314 43698 24396 43710
rect 24314 43638 24324 43698
rect 24384 43638 24396 43698
rect 24314 43624 24396 43638
rect 24874 43519 24968 43536
rect 24874 43457 24889 43519
rect 24951 43457 24968 43519
rect 22664 43442 22789 43451
rect 24874 43436 24968 43457
rect 22664 43290 22789 43317
rect 23207 43426 23330 43435
rect 23207 43294 23330 43303
rect 22664 43230 22696 43290
rect 22756 43230 22789 43290
rect 22664 43198 22789 43230
rect 6440 42700 6532 42722
rect 6440 42640 6456 42700
rect 6516 42640 6532 42700
rect 6440 42624 6532 42640
rect 25493 38479 25548 43818
rect 25582 38722 25634 43940
rect 25884 39792 25912 44157
rect 25582 38670 25740 38722
rect 25493 38424 25625 38479
rect 25688 38458 25740 38670
rect 2716 33624 3294 33680
rect 2501 33518 2553 33524
rect 2501 33460 2553 33466
rect 2382 33426 2434 33432
rect 2382 33368 2434 33374
rect 2299 33323 2351 33329
rect 2299 33265 2351 33271
rect 2153 33227 2205 33233
rect 2153 33169 2205 33175
rect 2240 14241 2268 31886
rect 3238 31396 3294 33624
rect 3424 33622 3484 33624
rect 3417 33566 3426 33622
rect 3482 33566 3491 33622
rect 3424 14672 3484 33566
rect 10971 33523 11018 33704
rect 10969 33517 11021 33523
rect 10969 33459 11021 33465
rect 6184 33426 6236 33432
rect 6184 33368 6236 33374
rect 5817 33322 5869 33328
rect 5817 33264 5869 33270
rect 5176 33232 5221 33251
rect 5173 33226 5225 33232
rect 5173 33168 5225 33174
rect 3548 33134 3604 33141
rect 3402 14590 3484 14672
rect 3546 33132 3606 33134
rect 3546 33076 3548 33132
rect 3604 33076 3606 33132
rect 2224 14232 2284 14241
rect 2224 14163 2284 14172
rect 3402 14201 3463 14590
rect 3546 14328 3606 33076
rect 5176 33004 5221 33168
rect 5818 33006 5867 33264
rect 6186 33256 6234 33368
rect 12251 33191 12313 33659
rect 13543 33291 13597 33649
rect 14178 33413 14251 33693
rect 15474 33552 15530 33736
rect 17407 33717 17462 33723
rect 17407 33611 17462 33662
rect 25570 33717 25625 38424
rect 26056 37070 26108 44211
rect 26346 37390 26402 44650
rect 26232 37334 26402 37390
rect 26457 43816 26530 43822
rect 25570 33656 25625 33662
rect 15474 33490 15530 33496
rect 26232 33552 26288 37334
rect 26457 37264 26530 43743
rect 26232 33490 26288 33496
rect 26333 37191 26530 37264
rect 26589 43695 26643 43701
rect 14178 33334 14251 33340
rect 26333 33413 26406 37191
rect 26589 37135 26643 43641
rect 26713 43575 26775 43581
rect 26713 43487 26775 43513
rect 26333 33334 26406 33340
rect 26471 37081 26643 37135
rect 26675 43425 26775 43487
rect 26471 33291 26525 37081
rect 26675 37027 26737 43425
rect 26784 43334 26790 43394
rect 26850 43334 26856 43394
rect 26565 36965 26737 37027
rect 26465 33237 26471 33291
rect 26525 33237 26531 33291
rect 13543 33231 13597 33237
rect 26565 33191 26627 36965
rect 26790 36886 26850 43334
rect 12245 33129 12251 33191
rect 12313 33129 12319 33191
rect 26565 33123 26627 33129
rect 26706 36826 26850 36886
rect 26910 43290 26970 43296
rect 26706 32860 26766 36826
rect 26910 36774 26970 43230
rect 26706 32804 26708 32860
rect 26764 32804 26766 32860
rect 26706 32802 26766 32804
rect 26810 36714 26970 36774
rect 26708 32795 26764 32802
rect 26810 32724 26870 36714
rect 26810 32668 26812 32724
rect 26868 32668 26870 32724
rect 26810 32666 26870 32668
rect 26812 32659 26868 32666
rect 3662 32456 3722 32465
rect 3662 32387 3722 32396
rect 3666 14472 3718 32387
rect 3666 14414 3718 14420
rect 4274 14324 4330 14331
rect 3546 14262 3606 14268
rect 4272 14322 17886 14324
rect 4272 14266 4274 14322
rect 4330 14266 17886 14322
rect 4272 14264 17886 14266
rect 17946 14264 17955 14324
rect 4274 14257 4330 14264
rect 3402 14198 17504 14201
rect 3402 14142 17445 14198
rect 17501 14142 17510 14198
rect 3402 14140 17504 14142
rect 2150 14015 2156 14088
rect 2229 14083 17096 14088
rect 2229 14020 17028 14083
rect 17091 14020 17100 14083
rect 2229 14015 17096 14020
rect 2464 13957 2596 13964
rect 2464 13952 17373 13957
rect 2464 13938 17312 13952
rect 2464 13882 2522 13938
rect 2578 13896 17312 13938
rect 17368 13896 17377 13952
rect 2578 13892 17373 13896
rect 2578 13882 2596 13892
rect 2522 13873 2578 13882
rect 2162 13763 2171 13833
rect 2241 13828 17783 13833
rect 2241 13768 17718 13828
rect 17778 13768 17787 13828
rect 2241 13763 17783 13768
rect 3540 13634 3546 13694
rect 3606 13634 3612 13694
rect 3446 13580 3502 13586
rect 2143 13392 2152 13452
rect 2212 13449 2221 13452
rect 2212 13395 3405 13449
rect 2212 13392 2221 13395
rect 2056 12076 3284 12104
rect 1571 11963 3197 12029
rect 1443 11831 3061 11882
rect 1294 11706 2924 11770
rect 2860 10514 2924 11706
rect 3010 10631 3061 11831
rect 3131 10781 3197 11963
rect 3256 10880 3284 12076
rect 3244 10874 3296 10880
rect 3244 10816 3296 10822
rect 3351 10785 3405 13395
rect 3446 10870 3502 13524
rect 3546 10963 3606 13634
rect 23869 12233 24000 12239
rect 24000 12068 25828 12199
rect 25959 12068 25965 12199
rect 23869 12027 24000 12033
rect 26458 12019 26716 12044
rect 11700 11815 11820 11838
rect 11700 11742 11724 11815
rect 11797 11742 11820 11815
rect 11700 11726 11820 11742
rect 13364 11810 13484 11846
rect 16716 11844 16844 11872
rect 13364 11750 13382 11810
rect 13442 11750 13484 11810
rect 13364 11734 13484 11750
rect 15064 11801 15184 11834
rect 15064 11739 15087 11801
rect 15149 11739 15184 11801
rect 16670 11748 16676 11844
rect 16772 11839 16844 11844
rect 16825 11753 16844 11839
rect 16772 11748 16844 11753
rect 15064 11722 15184 11739
rect 16716 11736 16844 11748
rect 18402 11817 18530 11866
rect 18402 11743 18417 11817
rect 18491 11743 18530 11817
rect 20042 11843 20170 11888
rect 20042 11769 20059 11843
rect 20133 11769 20170 11843
rect 20042 11752 20170 11769
rect 21688 11846 21816 11892
rect 21688 11774 21700 11846
rect 21772 11774 21816 11846
rect 21688 11756 21816 11774
rect 23388 11839 23516 11874
rect 18402 11730 18530 11743
rect 23388 11749 23403 11839
rect 23493 11749 23516 11839
rect 26458 11839 26490 12019
rect 26670 11839 26716 12019
rect 26458 11806 26716 11839
rect 23388 11738 23516 11749
rect 30096 11334 30152 11341
rect 30030 11274 30036 11334
rect 30096 11332 30154 11334
rect 30152 11276 30154 11332
rect 30096 11274 30154 11276
rect 30096 11267 30152 11274
rect 30220 11209 30303 14036
rect 30145 11126 30303 11209
rect 16687 10972 16777 10976
rect 16682 10967 16782 10972
rect 3546 10921 11458 10963
rect 3546 10916 3606 10921
rect 10560 10874 10612 10880
rect 3446 10814 5986 10870
rect 10612 10834 11320 10862
rect 10560 10816 10612 10822
rect 3351 10731 5804 10785
rect 3131 10709 3197 10715
rect 3010 10625 3062 10631
rect 3010 10567 3062 10573
rect 5546 10621 5646 10682
rect 5750 10628 5804 10731
rect 5930 10628 5986 10814
rect 11114 10778 11170 10782
rect 11110 10773 11175 10778
rect 11110 10717 11114 10773
rect 11170 10717 11175 10773
rect 5546 10531 5551 10621
rect 5641 10531 5646 10621
rect 11110 10618 11175 10717
rect 11292 10598 11320 10834
rect 11416 10654 11458 10921
rect 16682 10877 16687 10967
rect 16777 10877 16782 10967
rect 16682 10594 16782 10877
rect 30145 10871 30228 11126
rect 31989 11082 32073 11088
rect 30292 11010 30348 11017
rect 30290 11008 30350 11010
rect 30290 10952 30292 11008
rect 30348 10952 30350 11008
rect 30290 10950 30350 10952
rect 30410 10950 30416 11010
rect 30292 10943 30348 10950
rect 31980 10882 31989 11082
rect 32073 10882 32082 11082
rect 31989 10876 32073 10882
rect 30145 10797 30300 10871
rect 30145 10788 30333 10797
rect 16861 10781 16927 10787
rect 16861 10587 16927 10715
rect 17023 10774 17096 10783
rect 17442 10728 17503 10737
rect 17023 10598 17096 10701
rect 17307 10714 17372 10723
rect 17176 10626 17228 10632
rect 17307 10601 17372 10649
rect 17442 10585 17503 10667
rect 17864 10691 17942 10700
rect 30183 10659 30333 10788
rect 17176 10568 17228 10574
rect 17864 10561 17942 10613
rect 5546 10526 5646 10531
rect 5551 10522 5641 10526
rect 17558 10450 17564 10514
rect 17628 10450 17634 10514
rect 30177 10509 30183 10659
rect 30333 10509 30339 10659
rect 2860 10444 2924 10450
rect 503 9933 768 9939
rect 494 9842 503 9928
rect 768 9842 777 9928
rect 503 9831 768 9837
rect 870 7045 1130 7080
rect 196 6653 205 7043
rect 595 6653 604 7043
rect 870 6892 948 7045
rect 1101 6892 1130 7045
rect 870 6688 1130 6892
rect 205 6647 595 6653
rect 904 3839 1130 3878
rect 904 3701 935 3839
rect 1073 3701 1130 3839
rect 197 3458 206 3680
rect 594 3458 603 3680
rect 904 3650 1130 3701
rect 206 3452 594 3458
rect 918 637 1058 643
rect 909 497 918 637
rect 1058 497 1067 637
rect 918 491 1058 497
<< via2 >>
rect 14970 45008 15030 45068
rect 15518 45016 15578 45076
rect 2149 44770 2209 44830
rect 1281 38489 1371 38579
rect 205 26393 595 26783
rect 1423 37809 1513 37899
rect 1559 37129 1649 37219
rect 1749 35703 1839 35793
rect 1864 34360 1920 34416
rect 1750 13762 1839 13851
rect 1932 13394 1988 13450
rect 16074 44994 16134 45054
rect 17726 44986 17786 45046
rect 18683 44601 18761 44679
rect 20617 44655 20691 44729
rect 17170 44421 17243 44488
rect 19329 44455 19404 44530
rect 22545 44703 22627 44785
rect 26326 44738 26422 44834
rect 21905 44551 21979 44625
rect 17170 44415 17180 44421
rect 17180 44415 17232 44421
rect 17232 44415 17243 44421
rect 21261 44383 21335 44457
rect 11046 44212 11106 44272
rect 21580 44229 21661 44310
rect 25861 44208 25936 44283
rect 26101 44211 26191 44301
rect 4810 43986 4870 44046
rect 2592 43798 2652 43858
rect 2714 43640 2774 43700
rect 25572 44028 25644 44100
rect 23790 43743 23863 43816
rect 24324 43695 24384 43698
rect 24324 43641 24327 43695
rect 24327 43641 24381 43695
rect 24381 43641 24384 43695
rect 24324 43638 24384 43641
rect 24889 43457 24951 43519
rect 22664 43317 22789 43442
rect 23207 43403 23330 43426
rect 23207 43325 23229 43403
rect 23229 43325 23307 43403
rect 23307 43325 23330 43403
rect 23207 43303 23330 43325
rect 6456 42640 6516 42700
rect 3426 33566 3482 33622
rect 3548 33076 3604 33132
rect 2224 14172 2284 14232
rect 26708 32804 26764 32860
rect 26812 32668 26868 32724
rect 3662 32396 3722 32456
rect 4274 14266 4330 14322
rect 17886 14264 17946 14324
rect 17445 14142 17501 14198
rect 17028 14020 17091 14083
rect 2522 13882 2578 13938
rect 17312 13896 17368 13952
rect 2171 13763 2241 13833
rect 17718 13768 17778 13828
rect 2152 13392 2212 13452
rect 11729 11747 11792 11810
rect 13384 11752 13440 11808
rect 15090 11742 15146 11798
rect 16739 11753 16772 11839
rect 16772 11753 16825 11839
rect 18422 11748 18486 11812
rect 20064 11774 20128 11838
rect 21705 11779 21767 11841
rect 23408 11754 23488 11834
rect 26490 11839 26670 12019
rect 30096 11276 30152 11332
rect 11114 10717 11170 10773
rect 5551 10531 5641 10621
rect 16687 10877 16777 10967
rect 30292 10952 30348 11008
rect 31989 10882 32073 11082
rect 17023 10701 17096 10774
rect 17307 10649 17372 10714
rect 17442 10667 17503 10728
rect 17713 10581 17783 10651
rect 17864 10613 17942 10691
rect 503 9842 768 9928
rect 205 6806 595 7043
rect 205 6653 595 6806
rect 948 6892 1101 7045
rect 935 3701 1073 3839
rect 206 3594 594 3680
rect 206 3458 594 3594
rect 918 497 1058 637
<< metal3 >>
rect 14950 45073 15062 45090
rect 14950 45003 14965 45073
rect 15035 45003 15062 45073
rect 14950 44976 15062 45003
rect 15494 45081 15596 45100
rect 15494 45011 15513 45081
rect 15583 45011 15596 45081
rect 15494 44992 15596 45011
rect 16056 45059 16154 45076
rect 16056 44989 16069 45059
rect 16139 44989 16154 45059
rect 16056 44972 16154 44989
rect 17170 45054 17243 45120
rect 2144 44830 2214 44835
rect 16596 44830 16602 44832
rect 2144 44770 2149 44830
rect 2209 44770 16602 44830
rect 2144 44765 2214 44770
rect 16596 44768 16602 44770
rect 16666 44768 16672 44832
rect 17170 44493 17243 44981
rect 17702 45051 17800 45142
rect 17702 44981 17721 45051
rect 17791 44981 17800 45051
rect 17702 44954 17800 44981
rect 26321 44834 26427 44839
rect 22540 44785 22632 44790
rect 20612 44729 20696 44734
rect 18678 44679 18766 44684
rect 18678 44601 18683 44679
rect 18761 44601 19371 44679
rect 19449 44601 19455 44679
rect 20479 44655 20485 44729
rect 20559 44655 20617 44729
rect 20691 44655 20696 44729
rect 21025 44703 21031 44785
rect 21113 44703 22545 44785
rect 22627 44703 22632 44785
rect 25436 44738 25442 44834
rect 25538 44738 26326 44834
rect 26422 44738 26427 44834
rect 26321 44733 26427 44738
rect 22540 44698 22632 44703
rect 20612 44650 20696 44655
rect 21900 44625 21984 44630
rect 18678 44596 18766 44601
rect 21900 44551 21905 44625
rect 21979 44551 26541 44625
rect 26615 44551 26621 44625
rect 21900 44546 21984 44551
rect 19324 44530 19409 44535
rect 17165 44488 17248 44493
rect 17165 44415 17170 44488
rect 17243 44415 17248 44488
rect 19324 44455 19329 44530
rect 19404 44455 19928 44530
rect 20003 44455 20009 44530
rect 21256 44457 21340 44462
rect 19324 44450 19409 44455
rect 17165 44410 17248 44415
rect 21256 44383 21261 44457
rect 21335 44383 25995 44457
rect 26069 44383 26075 44457
rect 21256 44378 21340 44383
rect 21566 44315 21674 44322
rect 11041 44272 11111 44277
rect 17960 44274 18024 44280
rect 11376 44272 11382 44274
rect 11041 44212 11046 44272
rect 11106 44212 11382 44272
rect 11041 44207 11111 44212
rect 11376 44210 11382 44212
rect 11446 44210 11452 44274
rect 19026 44272 19032 44274
rect 18024 44212 19032 44272
rect 19026 44210 19032 44212
rect 19096 44210 19102 44274
rect 21566 44224 21575 44315
rect 21666 44224 21674 44315
rect 26096 44301 26196 44306
rect 25856 44283 25941 44288
rect 21566 44216 21674 44224
rect 17960 44204 18024 44210
rect 22141 44208 22147 44283
rect 22222 44208 25861 44283
rect 25936 44208 25941 44283
rect 25856 44203 25941 44208
rect 26096 44211 26101 44301
rect 26191 44211 27645 44301
rect 27735 44211 27741 44301
rect 26096 44206 26196 44211
rect 25567 44100 25649 44105
rect 4805 44046 4875 44051
rect 4805 43986 4810 44046
rect 4870 43986 25284 44046
rect 25567 44028 25572 44100
rect 25644 44028 27104 44100
rect 27176 44028 27182 44100
rect 25567 44023 25649 44028
rect 4805 43981 4875 43986
rect 25224 43922 25284 43986
rect 28766 43924 28830 43930
rect 2587 43858 2657 43863
rect 25224 43862 28766 43922
rect 18272 43858 18278 43860
rect 1413 43820 1731 43825
rect 248 43500 254 43820
rect 574 43819 1732 43820
rect 574 43501 1413 43819
rect 1731 43501 1732 43819
rect 2587 43798 2592 43858
rect 2652 43798 18278 43858
rect 2587 43793 2657 43798
rect 18272 43796 18278 43798
rect 18342 43796 18348 43860
rect 28766 43854 28830 43860
rect 23770 43821 23882 43836
rect 23770 43738 23785 43821
rect 23868 43738 23882 43821
rect 23770 43724 23882 43738
rect 2709 43700 2779 43705
rect 18824 43700 18830 43702
rect 2709 43640 2714 43700
rect 2774 43640 18830 43700
rect 2709 43635 2779 43640
rect 18824 43638 18830 43640
rect 18894 43638 18900 43702
rect 24294 43698 24422 43712
rect 24294 43697 24324 43698
rect 24384 43697 24422 43698
rect 24294 43633 24319 43697
rect 24389 43633 24422 43697
rect 24294 43610 24422 43633
rect 574 43500 1732 43501
rect 24856 43524 24992 43570
rect 1413 43495 1731 43500
rect 22659 43447 22794 43453
rect 24856 43452 24884 43524
rect 24956 43452 24992 43524
rect 690 43248 1844 43348
rect 22659 43317 22664 43322
rect 22789 43317 22794 43322
rect 22659 43312 22794 43317
rect 23186 43431 23356 43444
rect 23186 43298 23202 43431
rect 23335 43298 23356 43431
rect 24856 43426 24992 43452
rect 23186 43284 23356 43298
rect 200 26787 600 26788
rect 195 26389 201 26787
rect 599 26389 605 26787
rect 200 26388 600 26389
rect 690 10626 790 43248
rect 6440 42700 6532 42722
rect 21166 42700 21772 42712
rect 28198 42700 28204 42702
rect 6440 42640 6456 42700
rect 6516 42650 28204 42700
rect 6516 42640 21238 42650
rect 21690 42640 28204 42650
rect 6440 42624 6532 42640
rect 28198 42638 28204 42640
rect 28268 42638 28274 42702
rect 931 41895 1833 41973
rect 931 10783 1009 41895
rect 1106 40524 1844 40624
rect 1106 10972 1206 40524
rect 1988 39582 2048 39934
rect 1986 39576 2050 39582
rect 1986 39506 2050 39512
rect 1276 38579 1844 38584
rect 1276 38489 1281 38579
rect 1371 38489 1844 38579
rect 1276 38484 1844 38489
rect 1418 37899 1844 37904
rect 1418 37809 1423 37899
rect 1513 37809 1844 37899
rect 1418 37804 1844 37809
rect 1554 37219 1844 37224
rect 1554 37129 1559 37219
rect 1649 37129 1844 37219
rect 1554 37124 1844 37129
rect 1744 35793 1844 35864
rect 1744 35703 1749 35793
rect 1839 35703 1844 35793
rect 1744 35698 1844 35703
rect 1266 35114 1906 35174
rect 1266 13978 1326 35114
rect 1876 34464 1936 34494
rect 1784 34416 1936 34464
rect 1784 34360 1864 34416
rect 1920 34360 1936 34416
rect 1784 34352 1936 34360
rect 1876 34292 1936 34352
rect 3334 33754 3484 33814
rect 3424 33627 3484 33754
rect 3421 33622 3487 33627
rect 3421 33566 3426 33622
rect 3482 33566 3487 33622
rect 3421 33561 3487 33566
rect 3543 33134 3609 33137
rect 3543 33132 3784 33134
rect 3543 33076 3548 33132
rect 3604 33076 3784 33132
rect 3543 33074 3784 33076
rect 3543 33071 3609 33074
rect 26703 32862 26769 32865
rect 8284 32860 26769 32862
rect 8284 32804 26708 32860
rect 26764 32804 26769 32860
rect 8284 32802 26769 32804
rect 26703 32799 26769 32802
rect 26807 32726 26873 32729
rect 7644 32724 26873 32726
rect 7644 32668 26812 32724
rect 26868 32668 26873 32724
rect 7644 32666 26873 32668
rect 26807 32663 26873 32666
rect 3657 32456 3727 32461
rect 3657 32396 3662 32456
rect 3722 32396 3822 32456
rect 3657 32391 3727 32396
rect 26072 21110 26078 21174
rect 26142 21110 26148 21174
rect 11246 19168 11310 19174
rect 11310 19106 25598 19166
rect 11246 19098 11310 19104
rect 4269 14324 4335 14327
rect 3994 14322 4335 14324
rect 3994 14266 4274 14322
rect 4330 14266 4335 14322
rect 17881 14324 17951 14329
rect 17881 14293 17886 14324
rect 3994 14264 4335 14266
rect 2219 14232 2289 14237
rect 3994 14232 4054 14264
rect 4269 14261 4335 14264
rect 17864 14264 17886 14293
rect 17946 14264 17951 14324
rect 2219 14172 2224 14232
rect 2284 14172 4054 14232
rect 17864 14259 17951 14264
rect 17440 14198 17506 14203
rect 2219 14167 2289 14172
rect 17440 14142 17445 14198
rect 17501 14142 17506 14198
rect 17440 14137 17506 14142
rect 17023 14083 17096 14088
rect 17023 14020 17028 14083
rect 17091 14020 17096 14083
rect 1266 13964 2540 13978
rect 1266 13941 2596 13964
rect 1266 13938 2781 13941
rect 1266 13918 2522 13938
rect 2464 13882 2522 13918
rect 2578 13882 2781 13938
rect 2517 13879 2781 13882
rect 2517 13877 2583 13879
rect 1745 13851 1844 13856
rect 1745 13762 1750 13851
rect 1839 13833 2272 13851
rect 1839 13763 2171 13833
rect 2241 13763 2272 13833
rect 1839 13762 2272 13763
rect 1745 13757 1844 13762
rect 2166 13758 2246 13762
rect 1927 13452 1993 13455
rect 2147 13452 2217 13457
rect 1927 13450 2152 13452
rect 1927 13394 1932 13450
rect 1988 13394 2152 13450
rect 1927 13392 2152 13394
rect 2212 13392 2217 13452
rect 1927 13389 1993 13392
rect 2147 13387 2217 13392
rect 11700 11814 11820 11838
rect 11700 11743 11725 11814
rect 11796 11743 11820 11814
rect 11700 11726 11820 11743
rect 13364 11812 13484 11846
rect 16716 11844 16844 11872
rect 13364 11748 13380 11812
rect 13444 11748 13484 11812
rect 13364 11734 13484 11748
rect 15064 11802 15184 11834
rect 15064 11738 15086 11802
rect 15150 11738 15184 11802
rect 15064 11722 15184 11738
rect 16716 11748 16734 11844
rect 16830 11748 16844 11844
rect 16716 11736 16844 11748
rect 1106 10967 16782 10972
rect 1106 10877 16687 10967
rect 16777 10877 16782 10967
rect 1106 10872 16782 10877
rect 931 10777 3253 10783
rect 17023 10779 17096 14020
rect 17307 13952 17373 13957
rect 17307 13896 17312 13952
rect 17368 13896 17373 13952
rect 17307 13891 17373 13896
rect 11109 10777 11175 10778
rect 931 10773 11175 10777
rect 931 10717 11114 10773
rect 11170 10717 11175 10773
rect 931 10712 11175 10717
rect 17018 10774 17101 10779
rect 931 10705 3253 10712
rect 17018 10701 17023 10774
rect 17096 10701 17101 10774
rect 17307 10719 17372 13891
rect 17442 10733 17503 14137
rect 17864 14128 17946 14259
rect 17713 13828 17783 13833
rect 17713 13768 17718 13828
rect 17778 13768 17783 13828
rect 17437 10728 17508 10733
rect 17018 10696 17101 10701
rect 17302 10714 17377 10719
rect 17302 10649 17307 10714
rect 17372 10649 17377 10714
rect 17437 10667 17442 10728
rect 17503 10667 17508 10728
rect 17437 10662 17508 10667
rect 17713 10656 17783 13768
rect 17864 10696 17942 14128
rect 25538 13592 25598 19106
rect 26080 13758 26140 21110
rect 26080 13698 30480 13758
rect 25538 13532 30154 13592
rect 26485 12019 26675 12024
rect 18402 11816 18530 11866
rect 18402 11744 18418 11816
rect 18490 11744 18530 11816
rect 20042 11842 20170 11888
rect 20042 11770 20060 11842
rect 20132 11770 20170 11842
rect 20042 11752 20170 11770
rect 21688 11845 21816 11892
rect 21688 11775 21701 11845
rect 21771 11775 21816 11845
rect 21688 11756 21816 11775
rect 23388 11838 23516 11874
rect 18402 11730 18530 11744
rect 23388 11750 23404 11838
rect 23492 11750 23516 11838
rect 26485 11839 26490 12019
rect 26670 11839 26675 12019
rect 26485 11834 26675 11839
rect 23388 11738 23516 11750
rect 17859 10691 17947 10696
rect 17302 10644 17377 10649
rect 17708 10651 17788 10656
rect 690 10621 5646 10626
rect 690 10531 5551 10621
rect 5641 10531 5646 10621
rect 17708 10581 17713 10651
rect 17783 10581 17788 10651
rect 17859 10613 17864 10691
rect 17942 10613 17947 10691
rect 17859 10608 17947 10613
rect 17708 10576 17788 10581
rect 690 10526 5646 10531
rect 26490 10220 26670 11834
rect 30094 11337 30154 13532
rect 30091 11332 30157 11337
rect 30091 11276 30096 11332
rect 30152 11276 30157 11332
rect 30091 11271 30157 11276
rect 30287 11010 30353 11013
rect 30420 11010 30480 13698
rect 30287 11008 30480 11010
rect 30287 10952 30292 11008
rect 30348 10952 30480 11008
rect 30287 10950 30480 10952
rect 31984 11082 31994 11087
rect 30287 10947 30353 10950
rect 31984 10882 31989 11082
rect 31984 10877 31994 10882
rect 32078 10877 32084 11087
rect 326 10173 599 10179
rect 325 9837 326 10112
rect 599 9928 773 10112
rect 26490 10040 31816 10220
rect 31996 10040 32002 10220
rect 768 9842 773 9928
rect 599 9837 773 9842
rect 326 9769 599 9775
rect 900 7080 1148 7092
rect 200 7047 600 7048
rect 195 6649 201 7047
rect 599 6649 605 7047
rect 870 7045 1148 7080
rect 870 6966 948 7045
rect 1101 6966 1148 7045
rect 870 6718 900 6966
rect 870 6712 1148 6718
rect 870 6688 1130 6712
rect 200 6648 600 6649
rect 195 3453 201 3851
rect 599 3453 605 3851
rect 904 3844 1130 3878
rect 904 3696 930 3844
rect 1078 3696 1130 3844
rect 904 3650 1130 3696
rect 896 659 1080 665
rect 896 469 1080 475
rect 28235 207 28301 1489
rect 28235 135 28301 141
<< via3 >>
rect 14965 45068 15035 45073
rect 14965 45008 14970 45068
rect 14970 45008 15030 45068
rect 15030 45008 15035 45068
rect 14965 45003 15035 45008
rect 15513 45076 15583 45081
rect 15513 45016 15518 45076
rect 15518 45016 15578 45076
rect 15578 45016 15583 45076
rect 15513 45011 15583 45016
rect 16069 45054 16139 45059
rect 16069 44994 16074 45054
rect 16074 44994 16134 45054
rect 16134 44994 16139 45054
rect 16069 44989 16139 44994
rect 17170 44981 17243 45054
rect 16602 44768 16666 44832
rect 17721 45046 17791 45051
rect 17721 44986 17726 45046
rect 17726 44986 17786 45046
rect 17786 44986 17791 45046
rect 17721 44981 17791 44986
rect 19371 44601 19449 44679
rect 20485 44655 20559 44729
rect 21031 44703 21113 44785
rect 25442 44738 25538 44834
rect 26541 44551 26615 44625
rect 19928 44455 20003 44530
rect 25995 44383 26069 44457
rect 11382 44210 11446 44274
rect 17960 44210 18024 44274
rect 19032 44210 19096 44274
rect 21575 44310 21666 44315
rect 21575 44229 21580 44310
rect 21580 44229 21661 44310
rect 21661 44229 21666 44310
rect 21575 44224 21666 44229
rect 22147 44208 22222 44283
rect 27645 44211 27735 44301
rect 27104 44028 27176 44100
rect 28766 43860 28830 43924
rect 254 43500 574 43820
rect 1413 43501 1731 43819
rect 18278 43796 18342 43860
rect 23785 43816 23868 43821
rect 23785 43743 23790 43816
rect 23790 43743 23863 43816
rect 23863 43743 23868 43816
rect 23785 43738 23868 43743
rect 18830 43638 18894 43702
rect 24319 43638 24324 43697
rect 24324 43638 24384 43697
rect 24384 43638 24389 43697
rect 24319 43633 24389 43638
rect 22659 43442 22794 43447
rect 24884 43519 24956 43524
rect 24884 43457 24889 43519
rect 24889 43457 24951 43519
rect 24951 43457 24956 43519
rect 24884 43452 24956 43457
rect 22659 43322 22664 43442
rect 22664 43322 22789 43442
rect 22789 43322 22794 43442
rect 23202 43426 23335 43431
rect 23202 43303 23207 43426
rect 23207 43303 23330 43426
rect 23330 43303 23335 43426
rect 23202 43298 23335 43303
rect 201 26783 599 26787
rect 201 26393 205 26783
rect 205 26393 595 26783
rect 595 26393 599 26783
rect 201 26389 599 26393
rect 28204 42638 28268 42702
rect 1986 39512 2050 39576
rect 26078 21110 26142 21174
rect 11246 19104 11310 19168
rect 11725 11810 11796 11814
rect 11725 11747 11729 11810
rect 11729 11747 11792 11810
rect 11792 11747 11796 11810
rect 11725 11743 11796 11747
rect 13380 11808 13444 11812
rect 13380 11752 13384 11808
rect 13384 11752 13440 11808
rect 13440 11752 13444 11808
rect 13380 11748 13444 11752
rect 15086 11798 15150 11802
rect 15086 11742 15090 11798
rect 15090 11742 15146 11798
rect 15146 11742 15150 11798
rect 15086 11738 15150 11742
rect 16734 11839 16830 11844
rect 16734 11753 16739 11839
rect 16739 11753 16825 11839
rect 16825 11753 16830 11839
rect 16734 11748 16830 11753
rect 18418 11812 18490 11816
rect 18418 11748 18422 11812
rect 18422 11748 18486 11812
rect 18486 11748 18490 11812
rect 18418 11744 18490 11748
rect 20060 11838 20132 11842
rect 20060 11774 20064 11838
rect 20064 11774 20128 11838
rect 20128 11774 20132 11838
rect 20060 11770 20132 11774
rect 21701 11841 21771 11845
rect 21701 11779 21705 11841
rect 21705 11779 21767 11841
rect 21767 11779 21771 11841
rect 21701 11775 21771 11779
rect 23404 11834 23492 11838
rect 23404 11754 23408 11834
rect 23408 11754 23488 11834
rect 23488 11754 23492 11834
rect 23404 11750 23492 11754
rect 31994 11082 32078 11087
rect 31994 10882 32073 11082
rect 32073 10882 32078 11082
rect 31994 10877 32078 10882
rect 326 9928 599 10173
rect 31816 10040 31996 10220
rect 326 9842 503 9928
rect 503 9842 599 9928
rect 326 9775 599 9842
rect 201 7043 599 7047
rect 201 6653 205 7043
rect 205 6653 595 7043
rect 595 6653 599 7043
rect 201 6649 599 6653
rect 900 6892 948 6966
rect 948 6892 1101 6966
rect 1101 6892 1148 6966
rect 900 6718 1148 6892
rect 201 3680 599 3851
rect 201 3458 206 3680
rect 206 3458 594 3680
rect 594 3458 599 3680
rect 201 3453 599 3458
rect 930 3839 1078 3844
rect 930 3701 935 3839
rect 935 3701 1073 3839
rect 1073 3701 1078 3839
rect 930 3696 1078 3701
rect 896 637 1080 659
rect 896 497 918 637
rect 918 497 1058 637
rect 1058 497 1080 637
rect 896 475 1080 497
rect 28235 141 28301 207
<< metal4 >>
rect 6134 45106 6194 45152
rect 6686 45106 6746 45152
rect 7238 45106 7298 45152
rect 7790 45106 7850 45152
rect 6128 45099 7850 45106
rect 988 45098 7850 45099
rect 8342 45098 8402 45152
rect 988 45096 8444 45098
rect 8894 45096 8954 45152
rect 9446 45096 9506 45152
rect 9998 45096 10058 45152
rect 988 45094 10058 45096
rect 10550 45110 10610 45152
rect 11102 45110 11162 45152
rect 11654 45110 11714 45152
rect 12206 45110 12266 45152
rect 12758 45110 12818 45152
rect 13310 45110 13370 45152
rect 13862 45110 13922 45152
rect 14414 45110 14474 45152
rect 10550 45094 14474 45110
rect 988 45002 14474 45094
rect 14966 45090 15026 45152
rect 15518 45100 15578 45152
rect 330 44152 442 44154
rect 988 44152 1085 45002
rect 6128 44996 14474 45002
rect 6128 44994 12266 44996
rect 6134 44952 6194 44994
rect 6686 44952 6746 44994
rect 7238 44952 7298 44994
rect 7734 44990 12266 44994
rect 7790 44952 7850 44990
rect 8342 44984 12266 44990
rect 8342 44952 8402 44984
rect 8894 44952 8954 44984
rect 9122 44982 9234 44984
rect 9446 44952 9506 44984
rect 9998 44952 10058 44984
rect 10550 44968 12266 44984
rect 10550 44912 10610 44968
rect 11102 44952 11162 44968
rect 11654 44952 11714 44968
rect 12206 44952 12266 44968
rect 12758 44952 12818 44996
rect 13310 44952 13370 44996
rect 13862 44952 13922 44996
rect 14414 44952 14474 44996
rect 14950 45073 15062 45090
rect 14950 45003 14965 45073
rect 15035 45003 15062 45073
rect 14950 44976 15062 45003
rect 15494 45081 15596 45100
rect 15494 45011 15513 45081
rect 15583 45011 15596 45081
rect 16070 45076 16130 45152
rect 16622 45128 16682 45152
rect 15494 44992 15596 45011
rect 16056 45059 16154 45076
rect 14966 44952 15026 44976
rect 15518 44952 15578 44992
rect 16056 44989 16069 45059
rect 16139 44989 16154 45059
rect 16056 44972 16154 44989
rect 16070 44952 16130 44972
rect 16604 44952 16682 45128
rect 17174 45100 17234 45152
rect 17726 45142 17786 45152
rect 17170 45055 17243 45100
rect 17169 45054 17244 45055
rect 17169 44981 17170 45054
rect 17243 44981 17244 45054
rect 17169 44980 17244 44981
rect 17702 45051 17800 45142
rect 17702 44981 17721 45051
rect 17791 44981 17800 45051
rect 17174 44952 17234 44980
rect 17702 44954 17800 44981
rect 18278 45060 18338 45152
rect 17726 44952 17786 44954
rect 18278 44952 18340 45060
rect 18830 45029 18890 45152
rect 19382 45101 19442 45152
rect 19934 45130 19994 45152
rect 18830 45012 18891 45029
rect 18830 44952 18892 45012
rect 16604 44833 16664 44952
rect 16601 44832 16667 44833
rect 16601 44768 16602 44832
rect 16666 44768 16667 44832
rect 16601 44767 16667 44768
rect 11381 44274 11447 44275
rect 11381 44210 11382 44274
rect 11446 44272 11447 44274
rect 17959 44274 18025 44275
rect 17959 44272 17960 44274
rect 11446 44212 17960 44272
rect 11446 44210 11447 44212
rect 11381 44209 11447 44210
rect 17959 44210 17960 44212
rect 18024 44210 18025 44274
rect 17959 44209 18025 44210
rect 200 43820 600 44152
rect 200 43500 254 43820
rect 574 43500 600 43820
rect 200 26787 600 43500
rect 200 26389 201 26787
rect 599 26389 600 26787
rect 200 10173 600 26389
rect 200 9775 326 10173
rect 599 9775 600 10173
rect 200 7047 600 9775
rect 200 6649 201 7047
rect 599 6649 600 7047
rect 200 4620 600 6649
rect 800 44148 1200 44152
rect 800 44088 1204 44148
rect 800 43022 1200 44088
rect 18280 43861 18340 44952
rect 18277 43860 18343 43861
rect 1412 43819 1948 43820
rect 1412 43501 1413 43819
rect 1731 43540 1948 43819
rect 18277 43796 18278 43860
rect 18342 43796 18343 43860
rect 18277 43795 18343 43796
rect 18832 43703 18892 44952
rect 19371 44680 19449 45101
rect 19930 44985 19994 45130
rect 20486 45064 20546 45152
rect 21038 45089 21098 45152
rect 20486 45055 20550 45064
rect 19370 44679 19450 44680
rect 19370 44601 19371 44679
rect 19449 44601 19450 44679
rect 19370 44600 19450 44601
rect 19928 44531 20003 44985
rect 20485 44730 20559 45055
rect 21031 44786 21113 45089
rect 21590 45038 21650 45152
rect 22142 45079 22202 45152
rect 22694 45142 22754 45152
rect 22142 45054 22222 45079
rect 21590 45016 21652 45038
rect 21030 44785 21114 44786
rect 20484 44729 20560 44730
rect 20484 44655 20485 44729
rect 20559 44655 20560 44729
rect 21030 44703 21031 44785
rect 21113 44703 21114 44785
rect 21030 44702 21114 44703
rect 20484 44654 20560 44655
rect 19927 44530 20004 44531
rect 19927 44455 19928 44530
rect 20003 44455 20004 44530
rect 19927 44454 20004 44455
rect 21580 44322 21661 45016
rect 22140 44880 22222 45054
rect 21566 44315 21674 44322
rect 19031 44274 19097 44275
rect 19031 44210 19032 44274
rect 19096 44272 19097 44274
rect 19096 44212 21282 44272
rect 21566 44224 21575 44315
rect 21666 44224 21674 44315
rect 22147 44284 22222 44880
rect 21566 44216 21674 44224
rect 22146 44283 22223 44284
rect 19096 44210 19097 44212
rect 19031 44209 19097 44210
rect 21222 43814 21282 44212
rect 22146 44208 22147 44283
rect 22222 44208 22223 44283
rect 22146 44207 22223 44208
rect 21222 43754 22476 43814
rect 18829 43702 18895 43703
rect 18829 43638 18830 43702
rect 18894 43638 18895 43702
rect 18829 43637 18895 43638
rect 1731 43501 22288 43540
rect 1412 43500 22288 43501
rect 1628 43220 22288 43500
rect 800 42988 1482 43022
rect 800 42668 21628 42988
rect 800 42622 1482 42668
rect 800 42412 1202 42622
rect 800 22076 1200 42412
rect 21308 41508 21628 42668
rect 21968 41100 22288 43220
rect 22416 42888 22476 43754
rect 22664 43448 22789 45142
rect 23246 45054 23306 45152
rect 22658 43447 22795 43448
rect 22658 43322 22659 43447
rect 22794 43322 22795 43447
rect 23230 43444 23306 45054
rect 23798 45040 23858 45152
rect 24350 45108 24410 45152
rect 23790 43836 23863 45040
rect 24324 44952 24410 45108
rect 24902 45021 24962 45152
rect 25454 45070 25514 45152
rect 24889 44952 24962 45021
rect 23770 43821 23882 43836
rect 23770 43738 23785 43821
rect 23868 43738 23882 43821
rect 23770 43724 23882 43738
rect 22658 43321 22795 43322
rect 23186 43431 23356 43444
rect 23186 43298 23202 43431
rect 23335 43298 23356 43431
rect 23186 43284 23356 43298
rect 23790 43045 23863 43724
rect 24324 43710 24384 44952
rect 24314 43697 24396 43710
rect 24314 43633 24319 43697
rect 24389 43633 24396 43697
rect 24314 43624 24396 43633
rect 24324 43186 24384 43624
rect 24889 43536 24951 44952
rect 25442 44835 25538 45070
rect 26006 45053 26066 45152
rect 26558 45123 26618 45152
rect 25441 44834 25539 44835
rect 25441 44738 25442 44834
rect 25538 44738 25539 44834
rect 25441 44737 25539 44738
rect 25442 43578 25538 44737
rect 25995 44458 26069 45053
rect 26541 44952 26618 45123
rect 27110 45050 27170 45152
rect 27662 45137 27722 45152
rect 26541 44626 26615 44952
rect 26540 44625 26616 44626
rect 26540 44551 26541 44625
rect 26615 44551 26616 44625
rect 26540 44550 26616 44551
rect 25994 44457 26070 44458
rect 25994 44383 25995 44457
rect 26069 44383 26070 44457
rect 25994 44382 26070 44383
rect 25995 43733 26069 44382
rect 26541 43897 26615 44550
rect 27104 44101 27176 45050
rect 27645 44302 27735 45137
rect 28214 45120 28274 45152
rect 28206 44952 28274 45120
rect 28766 45076 28826 45152
rect 28766 44952 28828 45076
rect 29318 44952 29378 45152
rect 27644 44301 27736 44302
rect 27644 44211 27645 44301
rect 27735 44211 27736 44301
rect 27644 44210 27736 44211
rect 27103 44100 27177 44101
rect 27103 44028 27104 44100
rect 27176 44044 27177 44100
rect 27176 44028 27512 44044
rect 27103 44027 27512 44028
rect 27104 43972 27512 44027
rect 26541 43823 27335 43897
rect 25995 43659 27141 43733
rect 24874 43524 24968 43536
rect 24874 43452 24884 43524
rect 24956 43452 24968 43524
rect 25442 43482 26952 43578
rect 24874 43436 24968 43452
rect 24889 43361 24951 43436
rect 24889 43299 26725 43361
rect 24324 43126 26494 43186
rect 23790 42972 26328 43045
rect 22416 42828 26140 42888
rect 1985 39576 2051 39577
rect 1985 39512 1986 39576
rect 2050 39512 2051 39576
rect 1985 39511 2051 39512
rect 1988 22076 2048 39511
rect 800 21676 4666 22076
rect 800 6966 1200 21676
rect 1988 19166 2048 21676
rect 26080 21175 26140 42828
rect 26077 21174 26143 21175
rect 26077 21110 26078 21174
rect 26142 21110 26143 21174
rect 26077 21109 26143 21110
rect 26255 20843 26328 42972
rect 11724 20770 26328 20843
rect 11245 19168 11311 19169
rect 11245 19166 11246 19168
rect 1988 19106 11246 19166
rect 11245 19104 11246 19106
rect 11310 19104 11311 19168
rect 11245 19103 11311 19104
rect 11724 11814 11797 20770
rect 26434 20636 26494 43126
rect 11724 11743 11725 11814
rect 11796 11743 11797 11814
rect 13382 20576 26494 20636
rect 13382 11813 13442 20576
rect 26663 20419 26725 43299
rect 15087 20357 26725 20419
rect 13379 11812 13445 11813
rect 13379 11748 13380 11812
rect 13444 11748 13445 11812
rect 15087 11803 15149 20357
rect 26856 20192 26952 43482
rect 16734 20096 26952 20192
rect 16734 11845 16830 20096
rect 27067 19927 27141 43659
rect 18417 19853 27141 19927
rect 16733 11844 16831 11845
rect 13379 11747 13445 11748
rect 15085 11802 15151 11803
rect 11724 11742 11797 11743
rect 15085 11738 15086 11802
rect 15150 11738 15151 11802
rect 16733 11748 16734 11844
rect 16830 11748 16831 11844
rect 16733 11747 16831 11748
rect 18417 11816 18491 19853
rect 27261 19737 27335 43823
rect 18417 11744 18418 11816
rect 18490 11744 18491 11816
rect 20059 19663 27335 19737
rect 20059 11842 20133 19663
rect 27440 19522 27512 43972
rect 20059 11770 20060 11842
rect 20132 11770 20133 11842
rect 21700 19450 27512 19522
rect 21700 11845 21772 19450
rect 27645 19339 27735 44210
rect 28206 42703 28266 44952
rect 28768 43925 28828 44952
rect 28765 43924 28831 43925
rect 28765 43860 28766 43924
rect 28830 43860 28831 43924
rect 28765 43859 28831 43860
rect 28203 42702 28269 42703
rect 28203 42638 28204 42702
rect 28268 42638 28269 42702
rect 28203 42637 28269 42638
rect 21700 11775 21701 11845
rect 21771 11775 21772 11845
rect 21700 11774 21772 11775
rect 23403 19249 27735 19339
rect 23403 11838 23493 19249
rect 31857 13836 31930 14036
rect 20059 11769 20133 11770
rect 23403 11750 23404 11838
rect 23492 11750 23493 11838
rect 23403 11749 23493 11750
rect 18417 11743 18491 11744
rect 15085 11737 15151 11738
rect 31802 11088 32054 13836
rect 31802 11087 32079 11088
rect 31802 10877 31994 11087
rect 32078 10877 32079 11087
rect 31802 10876 32079 10877
rect 31802 10220 32054 10876
rect 31802 10040 31816 10220
rect 31996 10040 32054 10220
rect 31802 7464 32054 10040
rect 800 6718 900 6966
rect 1148 6718 1200 6966
rect 200 3866 602 4620
rect 200 3851 600 3866
rect 200 3453 201 3851
rect 599 3453 600 3851
rect 200 1000 600 3453
rect 800 3844 1200 6718
rect 800 3696 930 3844
rect 1078 3696 1200 3844
rect 800 1000 1200 3696
rect 30306 7212 32054 7464
rect 896 660 1080 1000
rect 895 659 1081 660
rect 895 475 896 659
rect 1080 475 1081 659
rect 895 474 1081 475
rect 30306 348 30558 7212
rect 28234 207 28302 208
rect 30298 207 30586 348
rect 3314 0 3494 204
rect 7178 0 7358 204
rect 11042 0 11222 204
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 28234 141 28235 207
rect 28301 141 30586 207
rect 28234 140 28302 141
rect 30298 96 30586 141
rect 30362 0 30542 96
use anl_switch  anl_switch_0
timestamp 1757923025
transform 1 0 28556 0 1 12962
box 1756 -3202 3533 463
use compr  compr_0
timestamp 1757923025
transform 1 0 24174 0 1 11715
box 510 -1403 5975 1713
use digital  digital_0
timestamp 1757921826
transform -1 0 26496 0 -1 44732
box 0 0 24752 13370
use flash_adc  flash_adc_0
timestamp 1757923025
transform 1 0 18258 0 1 6076
box -18000 -5600 12898 5562
use r2r_dac  r2r_dac_0
timestamp 1757914993
transform 1 0 7799 0 1 33431
box 2901 -22615 16695 -19768
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
