magic
tech sky130A
magscale 1 2
timestamp 1757923025
<< locali >>
rect 1826 -1247 2224 -1205
rect 1826 -1293 1862 -1247
rect 1788 -1370 1862 -1293
rect 2196 -1370 2224 -1247
rect 1788 -1404 2224 -1370
rect 1788 -1414 1838 -1404
rect 2114 -1938 2215 -1404
rect 1801 -2540 1847 -2536
rect 1801 -2566 1911 -2540
rect 2118 -2566 2219 -2027
rect 1801 -2604 1849 -2566
rect 1816 -2631 1849 -2604
rect 1828 -2651 1849 -2631
rect 2175 -2568 2219 -2566
rect 2175 -2651 2224 -2568
rect 1828 -2679 2224 -2651
<< viali >>
rect 1862 -1370 2196 -1247
rect 1849 -2651 2175 -2566
<< metal1 >>
rect 2346 294 2407 346
rect 2664 339 2725 348
rect 2657 296 2725 339
rect 2979 296 3040 348
rect 2657 287 2718 296
rect 3292 294 3353 346
rect 1983 -1205 2183 -1199
rect 1820 -1247 2222 -1205
rect 1820 -1311 1862 -1247
rect 1792 -1370 1862 -1311
rect 2196 -1370 2222 -1247
rect 1792 -1408 2222 -1370
rect 1792 -1565 1859 -1408
rect 1933 -1510 2000 -1457
rect 1792 -1646 1937 -1565
rect 1813 -1737 1937 -1646
rect 1995 -1736 2124 -1568
rect 2071 -1796 2124 -1736
rect 2275 -1626 2344 234
rect 2406 -1358 2475 237
rect 2586 -1355 2655 234
rect 2406 -1379 2476 -1358
rect 2406 -1389 2492 -1379
rect 2406 -1501 2410 -1389
rect 2477 -1501 2492 -1389
rect 2406 -1508 2492 -1501
rect 2406 -1561 2476 -1508
rect 2586 -1558 2656 -1355
rect 2719 -1387 2789 238
rect 2719 -1499 2721 -1387
rect 2788 -1499 2789 -1387
rect 2903 -1335 2972 236
rect 2903 -1388 2974 -1335
rect 3034 -1336 3103 243
rect 3221 -1333 3290 229
rect 3034 -1380 3107 -1336
rect 3034 -1388 3115 -1380
rect 3221 -1388 3292 -1333
rect 3354 -1335 3423 236
rect 2275 -1738 2281 -1626
rect 2275 -1743 2344 -1738
rect 2406 -1740 2475 -1561
rect 2586 -1624 2655 -1558
rect 2586 -1736 2592 -1624
rect 2586 -1743 2655 -1736
rect 2719 -1748 2789 -1499
rect 2904 -1511 2974 -1388
rect 3037 -1500 3041 -1388
rect 3108 -1500 3115 -1388
rect 3037 -1509 3115 -1500
rect 3037 -1511 3107 -1509
rect 3222 -1511 3292 -1388
rect 2903 -1538 2974 -1511
rect 2903 -1623 2972 -1538
rect 3034 -1539 3107 -1511
rect 3221 -1536 3292 -1511
rect 3353 -1390 3423 -1335
rect 3420 -1502 3423 -1390
rect 2903 -1735 2907 -1623
rect 3034 -1734 3103 -1539
rect 3221 -1624 3290 -1536
rect 3353 -1538 3423 -1502
rect 2903 -1741 2972 -1735
rect 3221 -1736 3226 -1624
rect 3354 -1651 3423 -1538
rect 3221 -1748 3290 -1736
rect 3354 -1741 3481 -1651
rect 1936 -1876 1994 -1799
rect 2071 -1848 3359 -1796
rect 2071 -1855 2752 -1848
rect 3035 -1852 3359 -1848
rect 3035 -1855 3273 -1852
rect 1833 -1941 2033 -1876
rect 1833 -2021 1966 -1941
rect 2025 -2021 2033 -1941
rect 1833 -2076 2033 -2021
rect 1936 -2161 1994 -2076
rect 1822 -2313 1931 -2212
rect 2071 -2215 2124 -1855
rect 3387 -1880 3481 -1741
rect 2787 -1885 2987 -1881
rect 2787 -1896 3137 -1885
rect 2154 -1950 2246 -1940
rect 2154 -2010 2166 -1950
rect 2238 -2010 2246 -1950
rect 2154 -2021 2246 -2010
rect 2162 -2107 2217 -2021
rect 2787 -2058 3037 -1896
rect 3103 -2058 3137 -1896
rect 2787 -2081 3137 -2058
rect 3317 -2080 3517 -1880
rect 2162 -2109 2380 -2107
rect 2162 -2159 3356 -2109
rect 2192 -2163 3356 -2159
rect 2346 -2164 3356 -2163
rect 1805 -2383 1931 -2313
rect 1995 -2383 2124 -2215
rect 2264 -2229 2338 -2214
rect 2264 -2341 2268 -2229
rect 2335 -2341 2338 -2229
rect 1805 -2547 1865 -2383
rect 1923 -2481 1990 -2428
rect 1996 -2547 2196 -2536
rect 1805 -2566 2196 -2547
rect 1805 -2651 1849 -2566
rect 2175 -2651 2196 -2566
rect 1805 -2685 2196 -2651
rect 1836 -2689 2196 -2685
rect 1996 -2736 2196 -2689
rect 2264 -2988 2338 -2341
rect 2411 -2431 2485 -2209
rect 2477 -2543 2485 -2431
rect 2411 -2983 2485 -2543
rect 2586 -2229 2660 -2214
rect 2586 -2341 2592 -2229
rect 2659 -2341 2660 -2229
rect 2586 -2988 2660 -2341
rect 2724 -2430 2798 -2214
rect 2724 -2542 2725 -2430
rect 2792 -2542 2798 -2430
rect 2724 -2988 2798 -2542
rect 2896 -2229 2970 -2211
rect 3387 -2214 3481 -2080
rect 2896 -2341 2903 -2229
rect 2896 -2985 2970 -2341
rect 3041 -2432 3115 -2214
rect 3103 -2544 3115 -2432
rect 3041 -2988 3115 -2544
rect 3205 -2230 3279 -2220
rect 3205 -2342 3212 -2230
rect 3205 -2994 3279 -2342
rect 3361 -2375 3481 -2214
rect 3361 -2428 3435 -2375
rect 3422 -2540 3435 -2428
rect 3361 -2988 3435 -2540
rect 2340 -3087 2407 -3034
rect 2655 -3087 2722 -3034
rect 2970 -3087 3037 -3034
rect 3285 -3084 3352 -3031
<< via1 >>
rect 2410 -1501 2477 -1389
rect 2721 -1499 2788 -1387
rect 2281 -1738 2348 -1626
rect 2592 -1736 2659 -1624
rect 3041 -1500 3108 -1388
rect 3353 -1502 3420 -1390
rect 2907 -1735 2974 -1623
rect 3226 -1736 3293 -1624
rect 1966 -2021 2025 -1941
rect 2166 -2010 2238 -1950
rect 3037 -2058 3103 -1896
rect 2268 -2341 2335 -2229
rect 2410 -2543 2477 -2431
rect 2592 -2341 2659 -2229
rect 2725 -2542 2792 -2430
rect 2903 -2341 2970 -2229
rect 3036 -2544 3103 -2432
rect 3212 -2342 3279 -2230
rect 3355 -2540 3422 -2428
<< metal2 >>
rect 2407 -1381 3414 -1374
rect 2407 -1387 3432 -1381
rect 2407 -1389 2721 -1387
rect 2407 -1501 2410 -1389
rect 2477 -1499 2721 -1389
rect 2788 -1388 3432 -1387
rect 2788 -1499 3041 -1388
rect 2477 -1500 3041 -1499
rect 3108 -1390 3432 -1388
rect 3108 -1500 3353 -1390
rect 2477 -1501 3353 -1500
rect 2407 -1502 3353 -1501
rect 3420 -1502 3432 -1390
rect 2407 -1509 3432 -1502
rect 3404 -1510 3432 -1509
rect 3276 -1618 3304 -1617
rect 2277 -1623 3304 -1618
rect 2277 -1624 2907 -1623
rect 2277 -1626 2592 -1624
rect 2277 -1637 2281 -1626
rect 2267 -1738 2281 -1637
rect 2348 -1736 2592 -1626
rect 2659 -1735 2907 -1624
rect 2974 -1624 3304 -1623
rect 2974 -1735 3226 -1624
rect 2659 -1736 3226 -1735
rect 3293 -1736 3304 -1624
rect 2348 -1738 3304 -1736
rect 2267 -1741 3304 -1738
rect 2267 -1748 2299 -1741
rect 3018 -1896 3124 -1741
rect 3276 -1746 3304 -1741
rect 1955 -1941 2252 -1932
rect 1955 -2021 1966 -1941
rect 2025 -1950 2252 -1941
rect 2025 -2010 2166 -1950
rect 2238 -2010 2252 -1950
rect 2025 -2021 2252 -2010
rect 1955 -2030 2252 -2021
rect 3018 -2058 3037 -1896
rect 3103 -2058 3124 -1896
rect 3018 -2223 3124 -2058
rect 3269 -2223 3297 -2221
rect 2260 -2229 3297 -2223
rect 2260 -2341 2268 -2229
rect 2335 -2341 2592 -2229
rect 2659 -2341 2903 -2229
rect 2970 -2230 3297 -2229
rect 2970 -2341 3212 -2230
rect 2260 -2342 3212 -2341
rect 3279 -2342 3297 -2230
rect 2260 -2346 3297 -2342
rect 2260 -2348 2310 -2346
rect 3269 -2350 3297 -2346
rect 3407 -2425 3435 -2419
rect 2397 -2428 3435 -2425
rect 2397 -2430 3355 -2428
rect 2397 -2431 2725 -2430
rect 2397 -2543 2410 -2431
rect 2477 -2542 2725 -2431
rect 2792 -2432 3355 -2430
rect 2792 -2542 3036 -2432
rect 2477 -2543 3036 -2542
rect 2397 -2544 3036 -2543
rect 3103 -2540 3355 -2432
rect 3422 -2540 3435 -2428
rect 3103 -2544 3435 -2540
rect 2397 -2548 3435 -2544
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 1757903622
transform 1 0 1967 0 1 -2293
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM4
timestamp 1757903622
transform 1 0 1967 0 1 -1640
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_PWNS5P  XM5
timestamp 1757903622
transform 1 0 2374 0 1 -2592
box -211 -610 211 610
use sky130_fd_pr__nfet_01v8_PWNS5P  XM6
timestamp 1757903622
transform 1 0 2690 0 1 -2592
box -211 -610 211 610
use sky130_fd_pr__nfet_01v8_PWNS5P  XM7
timestamp 1757903622
transform 1 0 3006 0 1 -2592
box -211 -610 211 610
use sky130_fd_pr__nfet_01v8_PWNS5P  XM8
timestamp 1757903622
transform 1 0 3322 0 1 -2592
box -211 -610 211 610
use sky130_fd_pr__pfet_01v8_XGA8MR  XM9
timestamp 1757903622
transform 1 0 2374 0 1 -756
box -211 -1219 211 1219
use sky130_fd_pr__pfet_01v8_XGA8MR  XM10
timestamp 1757903622
transform 1 0 2690 0 1 -756
box -211 -1219 211 1219
use sky130_fd_pr__pfet_01v8_XGA8MR  XM11
timestamp 1757903622
transform 1 0 3006 0 1 -756
box -211 -1219 211 1219
use sky130_fd_pr__pfet_01v8_XGA8MR  XM12
timestamp 1757903622
transform 1 0 3322 0 1 -756
box -211 -1219 211 1219
<< labels >>
flabel metal1 1833 -2076 2033 -1876 0 FreeSans 256 0 0 0 EN
port 1 nsew
flabel metal1 2787 -2081 2987 -1881 0 FreeSans 256 0 0 0 IN
port 2 nsew
flabel metal1 3317 -2080 3517 -1880 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel metal1 1996 -2736 2196 -2536 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 1983 -1399 2183 -1199 0 FreeSans 256 0 0 0 VDD
port 0 nsew
<< end >>
