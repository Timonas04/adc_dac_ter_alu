VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 27.305 209.005 27.475 209.195 ;
        RECT 30.065 209.005 30.235 209.195 ;
        RECT 31.445 209.025 31.615 209.195 ;
        RECT 31.905 209.005 32.075 209.195 ;
        RECT 37.425 209.005 37.595 209.195 ;
        RECT 40.645 209.005 40.815 209.195 ;
        RECT 46.165 209.005 46.335 209.195 ;
        RECT 51.685 209.005 51.855 209.195 ;
        RECT 53.525 209.005 53.695 209.195 ;
        RECT 55.180 209.005 55.350 209.195 ;
        RECT 59.045 209.005 59.215 209.195 ;
        RECT 64.565 209.005 64.735 209.195 ;
        RECT 66.415 209.050 66.575 209.160 ;
        RECT 67.325 209.005 67.495 209.195 ;
        RECT 68.705 209.005 68.875 209.195 ;
        RECT 74.220 209.055 74.340 209.165 ;
        RECT 74.690 209.005 74.860 209.195 ;
        RECT 78.360 209.055 78.480 209.165 ;
        RECT 79.285 209.005 79.455 209.195 ;
        RECT 81.120 209.055 81.240 209.165 ;
        RECT 81.595 209.005 81.765 209.195 ;
        RECT 83.425 209.045 83.595 209.195 ;
        RECT 27.165 208.195 28.535 209.005 ;
        RECT 28.545 208.325 30.375 209.005 ;
        RECT 28.545 208.095 29.890 208.325 ;
        RECT 31.765 208.195 37.275 209.005 ;
        RECT 37.285 208.195 40.035 209.005 ;
        RECT 40.055 208.135 40.485 208.920 ;
        RECT 40.505 208.195 46.015 209.005 ;
        RECT 46.025 208.195 51.535 209.005 ;
        RECT 51.545 208.195 52.915 209.005 ;
        RECT 52.935 208.135 53.365 208.920 ;
        RECT 53.385 208.195 54.755 209.005 ;
        RECT 54.765 208.325 58.665 209.005 ;
        RECT 54.765 208.095 55.695 208.325 ;
        RECT 58.905 208.195 64.415 209.005 ;
        RECT 64.425 208.195 65.795 209.005 ;
        RECT 65.815 208.135 66.245 208.920 ;
        RECT 67.185 208.225 68.555 209.005 ;
        RECT 68.565 208.195 74.075 209.005 ;
        RECT 74.545 208.325 78.215 209.005 ;
        RECT 74.545 208.095 75.470 208.325 ;
        RECT 78.695 208.135 79.125 208.920 ;
        RECT 79.145 208.195 80.975 209.005 ;
        RECT 81.445 208.225 82.815 209.005 ;
        RECT 82.825 208.095 83.715 209.045 ;
        RECT 84.795 209.005 84.965 209.195 ;
        RECT 85.265 209.005 85.435 209.195 ;
        RECT 87.105 209.045 87.275 209.195 ;
        RECT 87.575 209.050 87.735 209.160 ;
        RECT 83.745 208.225 85.115 209.005 ;
        RECT 85.125 208.225 86.495 209.005 ;
        RECT 86.505 208.095 87.395 209.045 ;
        RECT 88.495 209.005 88.665 209.195 ;
        RECT 91.245 209.005 91.415 209.195 ;
        RECT 92.160 209.055 92.280 209.165 ;
        RECT 92.635 209.005 92.805 209.195 ;
        RECT 94.015 209.050 94.175 209.160 ;
        RECT 96.765 209.025 96.935 209.195 ;
        RECT 96.765 209.005 96.930 209.025 ;
        RECT 97.225 209.005 97.395 209.195 ;
        RECT 99.060 209.055 99.180 209.165 ;
        RECT 99.500 209.025 99.670 209.195 ;
        RECT 104.120 209.055 104.240 209.165 ;
        RECT 105.055 209.050 105.215 209.160 ;
        RECT 99.560 209.005 99.670 209.025 ;
        RECT 107.345 209.005 107.515 209.195 ;
        RECT 107.805 209.005 107.975 209.195 ;
        RECT 110.095 209.005 110.265 209.195 ;
        RECT 111.485 209.005 111.655 209.195 ;
        RECT 111.940 209.055 112.060 209.165 ;
        RECT 113.785 209.005 113.955 209.195 ;
        RECT 115.160 209.005 115.330 209.195 ;
        RECT 117.005 209.005 117.175 209.195 ;
        RECT 117.935 209.050 118.095 209.160 ;
        RECT 120.225 209.005 120.395 209.195 ;
        RECT 121.605 209.005 121.775 209.195 ;
        RECT 122.065 209.005 122.235 209.195 ;
        RECT 125.755 209.005 125.925 209.195 ;
        RECT 127.125 209.005 127.295 209.195 ;
        RECT 128.505 209.005 128.675 209.195 ;
        RECT 130.800 209.055 130.920 209.165 ;
        RECT 131.270 209.005 131.440 209.195 ;
        RECT 137.695 209.005 137.865 209.195 ;
        RECT 138.160 209.055 138.280 209.165 ;
        RECT 139.545 209.005 139.715 209.195 ;
        RECT 88.345 208.225 89.715 209.005 ;
        RECT 89.725 208.325 91.555 209.005 ;
        RECT 89.725 208.095 91.070 208.325 ;
        RECT 91.575 208.135 92.005 208.920 ;
        RECT 92.485 208.225 93.855 209.005 ;
        RECT 95.095 208.325 96.930 209.005 ;
        RECT 97.085 208.325 98.915 209.005 ;
        RECT 99.560 208.325 103.975 209.005 ;
        RECT 95.095 208.095 96.025 208.325 ;
        RECT 97.570 208.095 98.915 208.325 ;
        RECT 100.045 208.095 103.975 208.325 ;
        RECT 104.455 208.135 104.885 208.920 ;
        RECT 105.825 208.325 107.655 209.005 ;
        RECT 105.825 208.095 107.170 208.325 ;
        RECT 107.675 208.095 109.025 209.005 ;
        RECT 109.045 208.225 110.415 209.005 ;
        RECT 110.425 208.225 111.795 209.005 ;
        RECT 112.265 208.325 114.095 209.005 ;
        RECT 112.265 208.095 113.610 208.325 ;
        RECT 114.125 208.095 115.475 209.005 ;
        RECT 115.485 208.325 117.315 209.005 ;
        RECT 115.485 208.095 116.830 208.325 ;
        RECT 117.335 208.135 117.765 208.920 ;
        RECT 118.705 208.325 120.535 209.005 ;
        RECT 118.705 208.095 120.050 208.325 ;
        RECT 120.545 208.225 121.915 209.005 ;
        RECT 121.925 208.195 125.595 209.005 ;
        RECT 125.605 208.225 126.975 209.005 ;
        RECT 126.985 208.225 128.355 209.005 ;
        RECT 128.365 208.325 130.195 209.005 ;
        RECT 128.850 208.095 130.195 208.325 ;
        RECT 130.215 208.135 130.645 208.920 ;
        RECT 131.125 208.095 136.255 209.005 ;
        RECT 136.645 208.225 138.015 209.005 ;
        RECT 138.485 208.195 139.855 209.005 ;
      LAYER nwell ;
        RECT 26.970 204.975 140.050 207.805 ;
      LAYER pwell ;
        RECT 27.165 203.775 28.535 204.585 ;
        RECT 28.545 204.455 29.890 204.685 ;
        RECT 28.545 203.775 30.375 204.455 ;
        RECT 30.385 203.775 34.055 204.585 ;
        RECT 34.065 203.775 35.435 204.585 ;
        RECT 35.445 203.775 36.815 204.555 ;
        RECT 36.825 203.775 40.035 204.685 ;
        RECT 40.055 203.860 40.485 204.645 ;
        RECT 40.505 204.455 41.435 204.685 ;
        RECT 40.505 203.775 44.405 204.455 ;
        RECT 44.645 203.775 50.155 204.585 ;
        RECT 50.180 203.775 51.995 204.685 ;
        RECT 52.005 203.775 55.215 204.685 ;
        RECT 55.225 204.455 56.155 204.685 ;
        RECT 55.225 203.775 59.125 204.455 ;
        RECT 59.365 203.775 63.035 204.585 ;
        RECT 63.980 203.775 65.795 204.685 ;
        RECT 65.815 203.860 66.245 204.645 ;
        RECT 66.735 203.775 69.465 204.685 ;
        RECT 69.485 203.775 72.235 204.585 ;
        RECT 73.295 204.455 74.225 204.685 ;
        RECT 72.390 203.775 74.225 204.455 ;
        RECT 74.545 204.455 75.470 204.685 ;
        RECT 74.545 203.775 78.215 204.455 ;
        RECT 78.225 203.775 80.055 204.585 ;
        RECT 80.065 204.455 80.995 204.685 ;
        RECT 80.065 203.775 83.965 204.455 ;
        RECT 84.665 203.775 86.015 204.685 ;
        RECT 27.305 203.565 27.475 203.775 ;
        RECT 28.685 203.565 28.855 203.755 ;
        RECT 30.065 203.585 30.235 203.775 ;
        RECT 30.525 203.585 30.695 203.775 ;
        RECT 32.365 203.565 32.535 203.755 ;
        RECT 32.825 203.565 32.995 203.755 ;
        RECT 34.205 203.585 34.375 203.775 ;
        RECT 36.505 203.585 36.675 203.775 ;
        RECT 36.965 203.585 37.135 203.775 ;
        RECT 38.345 203.565 38.515 203.755 ;
        RECT 40.460 203.565 40.630 203.755 ;
        RECT 40.920 203.585 41.090 203.775 ;
        RECT 44.785 203.585 44.955 203.775 ;
        RECT 46.165 203.585 46.335 203.755 ;
        RECT 46.635 203.610 46.795 203.720 ;
        RECT 47.545 203.585 47.715 203.755 ;
        RECT 50.305 203.585 50.475 203.775 ;
        RECT 52.145 203.585 52.315 203.775 ;
        RECT 46.165 203.565 46.330 203.585 ;
        RECT 27.165 202.755 28.535 203.565 ;
        RECT 28.545 202.755 31.295 203.565 ;
        RECT 31.305 202.785 32.675 203.565 ;
        RECT 32.685 202.755 38.195 203.565 ;
        RECT 38.205 202.755 40.035 203.565 ;
        RECT 40.045 202.885 43.945 203.565 ;
        RECT 44.495 202.885 46.330 203.565 ;
        RECT 47.550 203.565 47.715 203.585 ;
        RECT 52.605 203.565 52.775 203.755 ;
        RECT 53.525 203.565 53.695 203.755 ;
        RECT 55.360 203.615 55.480 203.725 ;
        RECT 55.640 203.585 55.810 203.775 ;
        RECT 56.100 203.565 56.270 203.755 ;
        RECT 59.505 203.585 59.675 203.775 ;
        RECT 62.265 203.565 62.435 203.755 ;
        RECT 62.735 203.610 62.895 203.720 ;
        RECT 63.195 203.620 63.355 203.730 ;
        RECT 64.105 203.585 64.275 203.775 ;
        RECT 64.570 203.565 64.740 203.755 ;
        RECT 65.020 203.615 65.140 203.725 ;
        RECT 65.490 203.565 65.660 203.755 ;
        RECT 66.400 203.615 66.520 203.725 ;
        RECT 68.710 203.565 68.880 203.755 ;
        RECT 69.165 203.585 69.335 203.775 ;
        RECT 69.625 203.585 69.795 203.775 ;
        RECT 72.390 203.755 72.555 203.775 ;
        RECT 72.385 203.585 72.555 203.755 ;
        RECT 74.690 203.585 74.860 203.775 ;
        RECT 77.010 203.565 77.180 203.755 ;
        RECT 77.440 203.565 77.610 203.755 ;
        RECT 78.365 203.585 78.535 203.775 ;
        RECT 79.285 203.565 79.455 203.755 ;
        RECT 80.480 203.585 80.650 203.775 ;
        RECT 81.120 203.615 81.240 203.725 ;
        RECT 84.340 203.615 84.460 203.725 ;
        RECT 84.990 203.565 85.160 203.755 ;
        RECT 85.730 203.585 85.900 203.775 ;
        RECT 86.045 203.755 86.935 204.685 ;
        RECT 86.965 203.775 88.335 204.555 ;
        RECT 86.000 203.735 86.935 203.755 ;
        RECT 86.000 203.565 86.170 203.735 ;
        RECT 86.645 203.585 86.815 203.735 ;
        RECT 88.015 203.585 88.185 203.775 ;
        RECT 89.265 203.735 90.155 204.685 ;
        RECT 90.185 203.775 91.555 204.555 ;
        RECT 91.575 203.860 92.005 204.645 ;
        RECT 92.025 203.775 93.395 204.555 ;
        RECT 93.865 203.775 96.615 204.685 ;
        RECT 96.825 204.595 97.775 204.685 ;
        RECT 96.825 203.775 98.755 204.595 ;
        RECT 101.210 204.485 102.595 204.685 ;
        RECT 98.925 203.805 102.595 204.485 ;
        RECT 90.335 203.755 90.505 203.775 ;
        RECT 88.495 203.620 88.655 203.730 ;
        RECT 89.865 203.605 90.035 203.735 ;
        RECT 90.325 203.605 90.505 203.755 ;
        RECT 47.550 202.885 49.385 203.565 ;
        RECT 40.045 202.655 40.975 202.885 ;
        RECT 44.495 202.655 45.425 202.885 ;
        RECT 48.455 202.655 49.385 202.885 ;
        RECT 49.705 202.655 52.915 203.565 ;
        RECT 52.935 202.695 53.365 203.480 ;
        RECT 53.385 202.755 55.215 203.565 ;
        RECT 55.685 202.885 59.585 203.565 ;
        RECT 55.685 202.655 56.615 202.885 ;
        RECT 59.835 202.655 62.565 203.565 ;
        RECT 63.505 202.655 64.855 203.565 ;
        RECT 65.345 202.655 68.265 203.565 ;
        RECT 68.565 202.655 72.865 203.565 ;
        RECT 73.165 202.655 77.240 203.565 ;
        RECT 77.325 202.655 78.675 203.565 ;
        RECT 78.695 202.695 79.125 203.480 ;
        RECT 79.145 202.755 80.975 203.565 ;
        RECT 81.675 202.885 85.575 203.565 ;
        RECT 84.645 202.655 85.575 202.885 ;
        RECT 85.585 202.885 89.485 203.565 ;
        RECT 85.585 202.655 86.515 202.885 ;
        RECT 89.725 202.655 90.615 203.605 ;
        RECT 90.785 203.565 90.955 203.755 ;
        RECT 92.170 203.565 92.340 203.755 ;
        RECT 93.085 203.585 93.255 203.775 ;
        RECT 93.540 203.615 93.660 203.725 ;
        RECT 95.850 203.565 96.020 203.755 ;
        RECT 96.305 203.585 96.475 203.775 ;
        RECT 98.605 203.755 98.755 203.775 ;
        RECT 98.605 203.585 98.775 203.755 ;
        RECT 99.065 203.585 99.235 203.805 ;
        RECT 101.225 203.775 102.595 203.805 ;
        RECT 102.605 203.775 103.975 204.555 ;
        RECT 104.005 203.775 105.355 204.685 ;
        RECT 105.375 203.775 106.725 204.685 ;
        RECT 107.305 203.775 109.495 204.685 ;
        RECT 110.845 204.485 112.255 204.685 ;
        RECT 109.520 203.805 112.255 204.485 ;
        RECT 101.360 203.565 101.530 203.755 ;
        RECT 101.820 203.615 101.940 203.725 ;
        RECT 102.285 203.585 102.455 203.755 ;
        RECT 102.755 203.585 102.925 203.775 ;
        RECT 105.040 203.755 105.210 203.775 ;
        RECT 105.040 203.585 105.215 203.755 ;
        RECT 105.505 203.585 105.675 203.775 ;
        RECT 106.880 203.615 107.000 203.725 ;
        RECT 109.180 203.585 109.350 203.775 ;
        RECT 109.645 203.585 109.815 203.805 ;
        RECT 110.860 203.775 112.255 203.805 ;
        RECT 112.265 203.775 115.935 204.685 ;
        RECT 115.945 203.775 117.295 204.685 ;
        RECT 117.335 203.860 117.765 204.645 ;
        RECT 117.785 204.005 119.620 204.685 ;
        RECT 117.930 203.775 119.620 204.005 ;
        RECT 120.545 203.775 124.645 204.685 ;
        RECT 125.145 203.775 134.250 204.455 ;
        RECT 134.345 203.775 135.715 204.555 ;
        RECT 135.725 203.775 137.095 204.555 ;
        RECT 137.520 203.775 138.475 204.455 ;
        RECT 138.485 203.775 139.855 204.585 ;
        RECT 102.305 203.565 102.455 203.585 ;
        RECT 105.045 203.565 105.215 203.585 ;
        RECT 110.100 203.565 110.270 203.755 ;
        RECT 110.565 203.585 110.735 203.755 ;
        RECT 115.620 203.585 115.790 203.775 ;
        RECT 117.010 203.585 117.180 203.775 ;
        RECT 117.930 203.585 118.100 203.775 ;
        RECT 120.220 203.615 120.340 203.725 ;
        RECT 120.690 203.585 120.860 203.775 ;
        RECT 110.570 203.565 110.735 203.585 ;
        RECT 121.605 203.565 121.775 203.755 ;
        RECT 90.645 202.785 92.015 203.565 ;
        RECT 92.025 202.655 95.695 203.565 ;
        RECT 95.705 202.655 99.375 203.565 ;
        RECT 99.485 202.655 101.675 203.565 ;
        RECT 102.305 202.745 104.235 203.565 ;
        RECT 103.285 202.655 104.235 202.745 ;
        RECT 104.455 202.695 104.885 203.480 ;
        RECT 104.905 202.885 106.735 203.565 ;
        RECT 105.390 202.655 106.735 202.885 ;
        RECT 106.745 202.655 110.415 203.565 ;
        RECT 110.570 202.885 112.405 203.565 ;
        RECT 112.810 202.885 121.915 203.565 ;
        RECT 122.065 203.335 122.235 203.755 ;
        RECT 124.820 203.615 124.940 203.725 ;
        RECT 125.285 203.585 125.455 203.775 ;
        RECT 129.885 203.565 130.055 203.755 ;
        RECT 130.805 203.565 130.975 203.755 ;
        RECT 134.485 203.565 134.655 203.755 ;
        RECT 134.940 203.615 135.060 203.725 ;
        RECT 135.405 203.585 135.575 203.775 ;
        RECT 136.325 203.565 136.495 203.755 ;
        RECT 136.785 203.565 136.955 203.775 ;
        RECT 137.245 203.585 137.415 203.755 ;
        RECT 139.545 203.565 139.715 203.775 ;
        RECT 123.345 203.335 127.435 203.565 ;
        RECT 111.475 202.655 112.405 202.885 ;
        RECT 121.960 202.655 127.435 203.335 ;
        RECT 127.455 202.885 130.195 203.565 ;
        RECT 130.215 202.695 130.645 203.480 ;
        RECT 130.665 202.885 133.405 203.565 ;
        RECT 133.435 202.655 134.785 203.565 ;
        RECT 135.265 202.785 136.635 203.565 ;
        RECT 136.645 202.885 138.475 203.565 ;
        RECT 137.130 202.655 138.475 202.885 ;
        RECT 138.485 202.755 139.855 203.565 ;
      LAYER nwell ;
        RECT 26.970 199.535 140.050 202.365 ;
      LAYER pwell ;
        RECT 27.165 198.335 28.535 199.145 ;
        RECT 28.545 198.335 34.055 199.145 ;
        RECT 34.065 198.335 37.735 199.145 ;
        RECT 38.685 198.335 40.035 199.245 ;
        RECT 40.055 198.420 40.485 199.205 ;
        RECT 42.575 199.155 44.165 199.245 ;
        RECT 41.595 198.335 44.165 199.155 ;
        RECT 44.195 198.335 45.545 199.245 ;
        RECT 46.505 198.335 47.855 199.245 ;
        RECT 47.865 198.335 49.680 199.245 ;
        RECT 49.705 198.335 52.455 199.145 ;
        RECT 52.775 199.015 53.705 199.245 ;
        RECT 54.765 199.015 55.695 199.245 ;
        RECT 52.775 198.335 54.610 199.015 ;
        RECT 54.765 198.335 58.665 199.015 ;
        RECT 58.905 198.335 62.575 199.145 ;
        RECT 62.585 198.335 63.935 199.245 ;
        RECT 63.965 198.335 65.795 199.145 ;
        RECT 65.815 198.420 66.245 199.205 ;
        RECT 66.265 198.335 68.095 199.145 ;
        RECT 68.565 198.335 71.775 199.245 ;
        RECT 71.785 198.335 77.295 199.145 ;
        RECT 77.305 198.335 78.675 199.145 ;
        RECT 78.705 198.335 80.055 199.245 ;
        RECT 80.065 199.015 80.995 199.245 ;
        RECT 80.065 198.335 83.965 199.015 ;
        RECT 84.285 198.335 87.285 199.245 ;
        RECT 87.425 198.335 88.775 199.245 ;
        RECT 88.805 198.335 91.555 199.145 ;
        RECT 91.575 198.420 92.005 199.205 ;
        RECT 92.035 198.335 94.765 199.245 ;
        RECT 95.260 198.335 97.075 199.245 ;
        RECT 97.085 198.335 100.295 199.245 ;
        RECT 100.305 198.335 104.175 199.245 ;
        RECT 104.445 198.335 107.655 199.245 ;
        RECT 107.665 199.015 109.010 199.245 ;
        RECT 109.505 199.015 111.095 199.245 ;
        RECT 107.665 198.335 109.495 199.015 ;
        RECT 109.505 198.335 113.175 199.015 ;
        RECT 113.185 198.335 117.315 199.245 ;
        RECT 117.335 198.420 117.765 199.205 ;
        RECT 117.785 198.335 121.455 199.145 ;
        RECT 121.935 198.335 123.285 199.245 ;
        RECT 123.315 198.335 124.665 199.245 ;
        RECT 124.685 198.335 126.055 199.115 ;
        RECT 126.525 198.335 135.630 199.015 ;
        RECT 27.305 198.125 27.475 198.335 ;
        RECT 28.685 198.125 28.855 198.335 ;
        RECT 34.205 198.145 34.375 198.335 ;
        RECT 37.895 198.180 38.055 198.290 ;
        RECT 38.530 198.125 38.700 198.315 ;
        RECT 38.800 198.145 38.970 198.335 ;
        RECT 41.595 198.315 41.735 198.335 ;
        RECT 40.655 198.180 40.815 198.290 ;
        RECT 41.565 198.145 41.735 198.315 ;
        RECT 42.670 198.125 42.840 198.315 ;
        RECT 43.405 198.125 43.575 198.315 ;
        RECT 45.245 198.145 45.415 198.335 ;
        RECT 45.715 198.180 45.875 198.290 ;
        RECT 46.620 198.145 46.790 198.335 ;
        RECT 49.385 198.145 49.555 198.335 ;
        RECT 49.845 198.125 50.015 198.335 ;
        RECT 54.445 198.315 54.610 198.335 ;
        RECT 50.315 198.170 50.475 198.280 ;
        RECT 52.605 198.125 52.775 198.315 ;
        RECT 53.525 198.125 53.695 198.315 ;
        RECT 54.445 198.145 54.615 198.315 ;
        RECT 55.180 198.145 55.350 198.335 ;
        RECT 59.045 198.125 59.215 198.335 ;
        RECT 63.650 198.145 63.820 198.335 ;
        RECT 64.105 198.145 64.275 198.335 ;
        RECT 64.560 198.175 64.680 198.285 ;
        RECT 65.025 198.125 65.195 198.315 ;
        RECT 66.405 198.145 66.575 198.335 ;
        RECT 67.790 198.125 67.960 198.315 ;
        RECT 68.240 198.175 68.360 198.285 ;
        RECT 71.460 198.145 71.630 198.335 ;
        RECT 71.925 198.145 72.095 198.335 ;
        RECT 72.845 198.125 73.015 198.315 ;
        RECT 73.305 198.125 73.475 198.315 ;
        RECT 77.445 198.145 77.615 198.335 ;
        RECT 78.820 198.145 78.990 198.335 ;
        RECT 79.280 198.175 79.400 198.285 ;
        RECT 79.750 198.125 79.920 198.315 ;
        RECT 80.480 198.145 80.650 198.335 ;
        RECT 81.595 198.170 81.755 198.280 ;
        RECT 82.505 198.125 82.675 198.315 ;
        RECT 84.345 198.145 84.515 198.335 ;
        RECT 85.725 198.125 85.895 198.315 ;
        RECT 88.490 198.145 88.660 198.335 ;
        RECT 88.945 198.145 89.115 198.335 ;
        RECT 89.405 198.125 89.575 198.315 ;
        RECT 91.245 198.165 91.415 198.315 ;
        RECT 27.165 197.315 28.535 198.125 ;
        RECT 28.545 197.315 34.055 198.125 ;
        RECT 35.215 197.445 39.115 198.125 ;
        RECT 39.355 197.445 43.255 198.125 ;
        RECT 38.185 197.215 39.115 197.445 ;
        RECT 42.325 197.215 43.255 197.445 ;
        RECT 43.265 197.315 48.775 198.125 ;
        RECT 48.795 197.215 50.145 198.125 ;
        RECT 51.085 197.215 52.900 198.125 ;
        RECT 52.935 197.255 53.365 198.040 ;
        RECT 53.385 197.315 58.895 198.125 ;
        RECT 58.905 197.315 64.415 198.125 ;
        RECT 64.885 197.215 67.605 198.125 ;
        RECT 67.645 197.215 71.315 198.125 ;
        RECT 71.325 197.445 73.155 198.125 ;
        RECT 73.165 197.315 78.675 198.125 ;
        RECT 78.695 197.255 79.125 198.040 ;
        RECT 79.605 197.215 81.435 198.125 ;
        RECT 82.445 197.215 85.445 198.125 ;
        RECT 85.585 197.315 89.255 198.125 ;
        RECT 89.265 197.315 90.635 198.125 ;
        RECT 90.645 197.215 91.535 198.165 ;
        RECT 91.715 198.125 91.885 198.315 ;
        RECT 92.165 198.145 92.335 198.335 ;
        RECT 93.085 198.125 93.255 198.315 ;
        RECT 94.920 198.175 95.040 198.285 ;
        RECT 95.385 198.145 95.555 198.335 ;
        RECT 96.765 198.145 96.935 198.315 ;
        RECT 97.235 198.170 97.395 198.280 ;
        RECT 99.985 198.145 100.155 198.335 ;
        RECT 100.450 198.145 100.620 198.335 ;
        RECT 101.825 198.145 101.995 198.315 ;
        RECT 104.125 198.145 104.295 198.315 ;
        RECT 96.765 198.125 96.930 198.145 ;
        RECT 101.825 198.125 101.985 198.145 ;
        RECT 104.125 198.125 104.275 198.145 ;
        RECT 105.045 198.125 105.215 198.315 ;
        RECT 106.430 198.125 106.600 198.315 ;
        RECT 107.345 198.145 107.515 198.335 ;
        RECT 109.185 198.145 109.355 198.335 ;
        RECT 109.650 198.125 109.820 198.315 ;
        RECT 112.860 198.145 113.030 198.335 ;
        RECT 113.330 198.145 113.500 198.335 ;
        RECT 113.785 198.125 113.955 198.315 ;
        RECT 117.925 198.145 118.095 198.335 ;
        RECT 121.600 198.175 121.720 198.285 ;
        RECT 122.985 198.145 123.155 198.335 ;
        RECT 123.445 198.145 123.615 198.335 ;
        RECT 125.735 198.145 125.905 198.335 ;
        RECT 126.665 198.315 126.835 198.335 ;
        RECT 126.200 198.175 126.320 198.285 ;
        RECT 126.665 198.145 126.860 198.315 ;
        RECT 126.690 198.125 126.860 198.145 ;
        RECT 129.885 198.125 130.055 198.315 ;
        RECT 130.810 198.125 130.980 198.315 ;
        RECT 134.485 198.125 134.655 198.315 ;
        RECT 135.745 198.295 136.635 199.245 ;
        RECT 136.645 198.335 138.475 199.245 ;
        RECT 138.485 198.335 139.855 199.145 ;
        RECT 135.865 198.145 136.035 198.295 ;
        RECT 137.715 198.170 137.875 198.280 ;
        RECT 138.160 198.145 138.330 198.335 ;
        RECT 139.545 198.125 139.715 198.335 ;
        RECT 91.565 197.345 92.935 198.125 ;
        RECT 92.960 197.215 94.775 198.125 ;
        RECT 95.095 197.445 96.930 198.125 ;
        RECT 95.095 197.215 96.025 197.445 ;
        RECT 98.330 197.215 101.985 198.125 ;
        RECT 102.345 197.305 104.275 198.125 ;
        RECT 102.345 197.215 103.295 197.305 ;
        RECT 104.455 197.255 104.885 198.040 ;
        RECT 104.915 197.215 106.265 198.125 ;
        RECT 106.285 197.215 109.400 198.125 ;
        RECT 109.505 197.215 113.635 198.125 ;
        RECT 113.645 197.445 122.750 198.125 ;
        RECT 122.845 197.215 126.920 198.125 ;
        RECT 126.985 197.215 130.195 198.125 ;
        RECT 130.215 197.255 130.645 198.040 ;
        RECT 130.665 197.215 134.335 198.125 ;
        RECT 134.345 198.095 136.185 198.125 ;
        RECT 134.345 197.445 137.510 198.095 ;
        RECT 134.830 197.415 137.510 197.445 ;
        RECT 134.830 197.215 136.185 197.415 ;
        RECT 138.485 197.315 139.855 198.125 ;
      LAYER nwell ;
        RECT 26.970 194.095 140.050 196.925 ;
      LAYER pwell ;
        RECT 27.165 192.895 28.535 193.705 ;
        RECT 28.545 193.575 29.890 193.805 ;
        RECT 28.545 192.895 30.375 193.575 ;
        RECT 30.385 192.895 35.895 193.705 ;
        RECT 35.905 192.895 39.575 193.705 ;
        RECT 40.055 192.980 40.485 193.765 ;
        RECT 40.505 192.895 43.715 193.805 ;
        RECT 44.180 193.125 46.015 193.805 ;
        RECT 44.180 192.895 45.870 193.125 ;
        RECT 46.025 192.895 47.395 193.705 ;
        RECT 47.405 192.895 49.220 193.805 ;
        RECT 49.245 192.895 52.915 193.705 ;
        RECT 53.095 192.895 56.595 193.805 ;
        RECT 56.605 192.895 57.975 193.705 ;
        RECT 57.985 192.895 59.815 193.805 ;
        RECT 59.825 192.895 61.655 193.705 ;
        RECT 62.140 193.575 63.510 193.805 ;
        RECT 62.140 192.895 64.415 193.575 ;
        RECT 64.425 192.895 65.795 193.705 ;
        RECT 65.815 192.980 66.245 193.765 ;
        RECT 66.265 193.575 67.185 193.805 ;
        RECT 66.265 192.895 69.850 193.575 ;
        RECT 69.960 192.895 73.615 193.805 ;
        RECT 73.640 192.895 75.455 193.805 ;
        RECT 75.465 192.895 79.135 193.705 ;
        RECT 79.605 192.895 81.435 193.805 ;
        RECT 82.420 192.895 86.495 193.805 ;
        RECT 86.505 192.895 90.160 193.805 ;
        RECT 90.185 192.895 91.555 193.705 ;
        RECT 91.575 192.980 92.005 193.765 ;
        RECT 92.110 192.895 101.215 193.575 ;
        RECT 102.155 192.895 104.895 193.575 ;
        RECT 104.905 192.895 108.115 193.805 ;
        RECT 108.125 192.895 117.230 193.575 ;
        RECT 117.335 192.980 117.765 193.765 ;
        RECT 137.130 193.575 138.475 193.805 ;
        RECT 117.785 192.895 126.890 193.575 ;
        RECT 126.985 192.895 136.090 193.575 ;
        RECT 136.645 192.895 138.475 193.575 ;
        RECT 138.485 192.895 139.855 193.705 ;
        RECT 27.305 192.685 27.475 192.895 ;
        RECT 28.685 192.685 28.855 192.875 ;
        RECT 30.065 192.705 30.235 192.895 ;
        RECT 30.525 192.705 30.695 192.895 ;
        RECT 32.365 192.685 32.535 192.875 ;
        RECT 32.825 192.685 32.995 192.875 ;
        RECT 36.045 192.705 36.215 192.895 ;
        RECT 38.345 192.685 38.515 192.875 ;
        RECT 39.720 192.735 39.840 192.845 ;
        RECT 41.100 192.685 41.270 192.875 ;
        RECT 41.565 192.685 41.735 192.875 ;
        RECT 42.945 192.685 43.115 192.875 ;
        RECT 43.405 192.705 43.575 192.895 ;
        RECT 44.325 192.685 44.495 192.875 ;
        RECT 45.700 192.705 45.870 192.895 ;
        RECT 46.165 192.705 46.335 192.895 ;
        RECT 48.005 192.685 48.175 192.875 ;
        RECT 48.925 192.705 49.095 192.895 ;
        RECT 49.385 192.705 49.555 192.895 ;
        RECT 53.095 192.875 53.230 192.895 ;
        RECT 50.765 192.685 50.935 192.875 ;
        RECT 51.225 192.685 51.395 192.875 ;
        RECT 53.060 192.705 53.230 192.875 ;
        RECT 53.510 192.685 53.680 192.875 ;
        RECT 56.745 192.705 56.915 192.895 ;
        RECT 58.130 192.705 58.300 192.895 ;
        RECT 59.045 192.705 59.215 192.875 ;
        RECT 59.965 192.705 60.135 192.895 ;
        RECT 59.045 192.685 59.195 192.705 ;
        RECT 60.430 192.685 60.600 192.875 ;
        RECT 60.885 192.685 61.055 192.875 ;
        RECT 61.800 192.735 61.920 192.845 ;
        RECT 64.100 192.705 64.270 192.895 ;
        RECT 64.565 192.705 64.735 192.895 ;
        RECT 66.410 192.705 66.580 192.895 ;
        RECT 69.165 192.685 69.335 192.875 ;
        RECT 69.625 192.685 69.795 192.875 ;
        RECT 72.385 192.685 72.555 192.875 ;
        RECT 73.300 192.705 73.470 192.895 ;
        RECT 73.765 192.705 73.935 192.895 ;
        RECT 75.605 192.705 75.775 192.895 ;
        RECT 79.285 192.845 79.455 192.875 ;
        RECT 77.915 192.730 78.075 192.840 ;
        RECT 79.280 192.735 79.455 192.845 ;
        RECT 79.285 192.685 79.455 192.735 ;
        RECT 79.750 192.705 79.920 192.895 ;
        RECT 81.595 192.740 81.755 192.850 ;
        RECT 82.040 192.685 82.210 192.875 ;
        RECT 82.480 192.705 82.650 192.895 ;
        RECT 86.650 192.705 86.820 192.895 ;
        RECT 88.025 192.685 88.195 192.875 ;
        RECT 88.485 192.685 88.655 192.875 ;
        RECT 90.325 192.705 90.495 192.895 ;
        RECT 91.245 192.685 91.415 192.875 ;
        RECT 93.545 192.685 93.715 192.875 ;
        RECT 94.000 192.685 94.170 192.875 ;
        RECT 98.145 192.685 98.315 192.875 ;
        RECT 99.530 192.685 99.700 192.875 ;
        RECT 99.985 192.685 100.155 192.875 ;
        RECT 100.905 192.705 101.075 192.895 ;
        RECT 101.375 192.740 101.535 192.850 ;
        RECT 104.125 192.685 104.295 192.875 ;
        RECT 104.585 192.705 104.755 192.895 ;
        RECT 105.050 192.705 105.220 192.895 ;
        RECT 105.965 192.685 106.135 192.875 ;
        RECT 108.265 192.705 108.435 192.895 ;
        RECT 115.165 192.685 115.335 192.875 ;
        RECT 117.925 192.705 118.095 192.895 ;
        RECT 124.365 192.685 124.535 192.875 ;
        RECT 124.830 192.685 125.000 192.875 ;
        RECT 127.125 192.705 127.295 192.895 ;
        RECT 129.890 192.685 130.060 192.875 ;
        RECT 130.810 192.685 130.980 192.875 ;
        RECT 134.485 192.705 134.655 192.875 ;
        RECT 136.320 192.735 136.440 192.845 ;
        RECT 136.785 192.705 136.955 192.895 ;
        RECT 138.160 192.735 138.280 192.845 ;
        RECT 134.485 192.685 134.685 192.705 ;
        RECT 139.545 192.685 139.715 192.895 ;
        RECT 27.165 191.875 28.535 192.685 ;
        RECT 28.545 192.005 30.375 192.685 ;
        RECT 31.305 191.905 32.675 192.685 ;
        RECT 32.685 191.875 38.195 192.685 ;
        RECT 38.205 191.875 40.035 192.685 ;
        RECT 40.065 191.775 41.415 192.685 ;
        RECT 41.425 191.875 42.795 192.685 ;
        RECT 42.815 191.775 44.165 192.685 ;
        RECT 44.185 191.875 47.855 192.685 ;
        RECT 47.865 191.875 49.235 192.685 ;
        RECT 49.245 191.775 51.060 192.685 ;
        RECT 51.100 191.775 52.915 192.685 ;
        RECT 52.935 191.815 53.365 192.600 ;
        RECT 53.395 191.775 57.055 192.685 ;
        RECT 57.265 191.865 59.195 192.685 ;
        RECT 57.265 191.775 58.215 191.865 ;
        RECT 59.365 191.775 60.715 192.685 ;
        RECT 60.745 191.875 66.255 192.685 ;
        RECT 66.265 192.005 69.475 192.685 ;
        RECT 69.485 192.005 72.235 192.685 ;
        RECT 66.265 191.775 67.400 192.005 ;
        RECT 71.305 191.775 72.235 192.005 ;
        RECT 72.245 191.875 77.755 192.685 ;
        RECT 78.695 191.815 79.125 192.600 ;
        RECT 79.145 191.875 81.895 192.685 ;
        RECT 81.915 191.775 85.115 192.685 ;
        RECT 85.125 191.775 88.335 192.685 ;
        RECT 88.345 191.875 91.095 192.685 ;
        RECT 91.105 191.905 92.475 192.685 ;
        RECT 92.485 191.905 93.855 192.685 ;
        RECT 93.885 191.775 95.235 192.685 ;
        RECT 95.245 191.775 98.455 192.685 ;
        RECT 98.465 191.775 99.815 192.685 ;
        RECT 99.845 192.005 102.595 192.685 ;
        RECT 101.665 191.775 102.595 192.005 ;
        RECT 102.605 191.775 104.420 192.685 ;
        RECT 104.455 191.815 104.885 192.600 ;
        RECT 104.915 191.775 106.265 192.685 ;
        RECT 106.370 192.005 115.475 192.685 ;
        RECT 115.570 192.005 124.675 192.685 ;
        RECT 124.685 191.775 128.815 192.685 ;
        RECT 128.825 191.775 130.175 192.685 ;
        RECT 130.215 191.815 130.645 192.600 ;
        RECT 130.665 191.775 134.320 192.685 ;
        RECT 134.485 192.005 138.015 192.685 ;
        RECT 135.190 191.775 138.015 192.005 ;
        RECT 138.485 191.875 139.855 192.685 ;
      LAYER nwell ;
        RECT 26.970 188.655 140.050 191.485 ;
      LAYER pwell ;
        RECT 27.165 187.455 28.535 188.265 ;
        RECT 28.545 187.455 31.295 188.265 ;
        RECT 31.315 187.455 32.665 188.365 ;
        RECT 32.685 187.455 36.355 188.265 ;
        RECT 36.365 187.455 38.195 188.365 ;
        RECT 38.205 187.455 40.035 188.365 ;
        RECT 40.055 187.540 40.485 188.325 ;
        RECT 40.505 188.165 41.435 188.365 ;
        RECT 42.765 188.165 43.715 188.365 ;
        RECT 40.505 187.685 43.715 188.165 ;
        RECT 40.650 187.485 43.715 187.685 ;
        RECT 27.305 187.245 27.475 187.455 ;
        RECT 28.685 187.435 28.855 187.455 ;
        RECT 28.660 187.265 28.855 187.435 ;
        RECT 31.445 187.265 31.615 187.455 ;
        RECT 32.825 187.265 32.995 187.455 ;
        RECT 28.720 187.245 28.830 187.265 ;
        RECT 33.285 187.245 33.455 187.435 ;
        RECT 35.120 187.295 35.240 187.405 ;
        RECT 35.590 187.245 35.760 187.435 ;
        RECT 36.510 187.265 36.680 187.455 ;
        RECT 38.350 187.265 38.520 187.455 ;
        RECT 38.805 187.245 38.975 187.435 ;
        RECT 40.650 187.265 40.820 187.485 ;
        RECT 42.780 187.455 43.715 187.485 ;
        RECT 43.725 187.455 49.235 188.265 ;
        RECT 49.245 187.455 51.075 188.265 ;
        RECT 51.555 187.455 55.675 188.365 ;
        RECT 55.685 187.455 57.035 188.365 ;
        RECT 57.065 187.455 58.415 188.365 ;
        RECT 58.445 187.455 62.115 188.265 ;
        RECT 63.055 187.455 64.405 188.365 ;
        RECT 64.425 187.455 65.795 188.265 ;
        RECT 65.815 187.540 66.245 188.325 ;
        RECT 68.545 188.135 69.475 188.365 ;
        RECT 66.725 187.455 69.475 188.135 ;
        RECT 69.495 187.455 72.225 188.365 ;
        RECT 72.245 188.165 73.190 188.365 ;
        RECT 74.525 188.165 75.455 188.365 ;
        RECT 72.245 187.685 75.455 188.165 ;
        RECT 72.245 187.485 75.315 187.685 ;
        RECT 72.245 187.455 73.190 187.485 ;
        RECT 27.165 186.435 28.535 187.245 ;
        RECT 28.720 186.565 33.135 187.245 ;
        RECT 29.205 186.335 33.135 186.565 ;
        RECT 33.145 186.435 34.975 187.245 ;
        RECT 35.445 186.565 38.655 187.245 ;
        RECT 38.665 186.565 42.335 187.245 ;
        RECT 42.490 187.215 42.660 187.435 ;
        RECT 43.865 187.265 44.035 187.455 ;
        RECT 45.705 187.245 45.875 187.435 ;
        RECT 48.475 187.290 48.635 187.400 ;
        RECT 49.385 187.265 49.555 187.455 ;
        RECT 51.225 187.405 51.395 187.435 ;
        RECT 51.220 187.295 51.395 187.405 ;
        RECT 51.225 187.265 51.395 187.295 ;
        RECT 51.225 187.245 51.375 187.265 ;
        RECT 51.685 187.245 51.855 187.435 ;
        RECT 53.525 187.265 53.695 187.455 ;
        RECT 55.365 187.265 55.535 187.455 ;
        RECT 56.750 187.435 56.920 187.455 ;
        RECT 57.210 187.435 57.380 187.455 ;
        RECT 56.745 187.265 56.920 187.435 ;
        RECT 57.205 187.265 57.380 187.435 ;
        RECT 58.585 187.265 58.755 187.455 ;
        RECT 62.275 187.300 62.435 187.410 ;
        RECT 56.745 187.245 56.915 187.265 ;
        RECT 57.205 187.245 57.375 187.265 ;
        RECT 62.725 187.245 62.895 187.435 ;
        RECT 63.185 187.265 63.355 187.455 ;
        RECT 64.565 187.265 64.735 187.455 ;
        RECT 65.480 187.245 65.650 187.435 ;
        RECT 66.400 187.295 66.520 187.405 ;
        RECT 66.865 187.245 67.035 187.455 ;
        RECT 71.925 187.435 72.095 187.455 ;
        RECT 71.920 187.265 72.095 187.435 ;
        RECT 71.920 187.245 72.090 187.265 ;
        RECT 72.390 187.245 72.560 187.435 ;
        RECT 75.145 187.265 75.315 187.485 ;
        RECT 75.465 187.455 80.975 188.265 ;
        RECT 80.985 187.455 84.655 188.265 ;
        RECT 84.665 187.455 86.035 188.265 ;
        RECT 86.060 187.455 87.875 188.365 ;
        RECT 88.805 187.455 90.155 188.365 ;
        RECT 90.205 187.455 91.555 188.365 ;
        RECT 91.575 187.540 92.005 188.325 ;
        RECT 92.025 187.455 95.235 188.365 ;
        RECT 95.705 187.455 97.055 188.365 ;
        RECT 97.170 187.455 106.275 188.135 ;
        RECT 106.285 187.455 108.115 188.365 ;
        RECT 108.210 187.455 117.315 188.135 ;
        RECT 117.335 187.540 117.765 188.325 ;
        RECT 117.870 187.455 126.975 188.135 ;
        RECT 126.985 187.455 136.090 188.135 ;
        RECT 136.285 187.455 138.475 188.365 ;
        RECT 138.485 187.455 139.855 188.265 ;
        RECT 75.605 187.265 75.775 187.455 ;
        RECT 77.905 187.265 78.075 187.435 ;
        RECT 78.360 187.295 78.480 187.405 ;
        RECT 77.905 187.245 78.070 187.265 ;
        RECT 80.210 187.245 80.380 187.435 ;
        RECT 80.665 187.245 80.835 187.435 ;
        RECT 81.125 187.265 81.295 187.455 ;
        RECT 82.505 187.245 82.675 187.435 ;
        RECT 84.345 187.245 84.515 187.435 ;
        RECT 84.805 187.265 84.975 187.455 ;
        RECT 86.185 187.265 86.355 187.455 ;
        RECT 88.035 187.300 88.195 187.410 ;
        RECT 89.870 187.265 90.040 187.455 ;
        RECT 90.320 187.265 90.490 187.455 ;
        RECT 86.185 187.245 86.385 187.265 ;
        RECT 91.710 187.245 91.880 187.435 ;
        RECT 92.170 187.245 92.340 187.435 ;
        RECT 94.925 187.265 95.095 187.455 ;
        RECT 95.380 187.295 95.500 187.405 ;
        RECT 95.850 187.265 96.020 187.455 ;
        RECT 105.965 187.435 106.135 187.455 ;
        RECT 97.685 187.245 97.855 187.435 ;
        RECT 98.145 187.265 98.315 187.435 ;
        RECT 102.280 187.295 102.400 187.405 ;
        RECT 98.155 187.245 98.315 187.265 ;
        RECT 104.125 187.245 104.295 187.435 ;
        RECT 105.965 187.265 106.140 187.435 ;
        RECT 106.430 187.265 106.600 187.455 ;
        RECT 109.645 187.265 109.815 187.435 ;
        RECT 110.100 187.295 110.220 187.405 ;
        RECT 105.970 187.245 106.140 187.265 ;
        RECT 109.615 187.245 109.815 187.265 ;
        RECT 110.565 187.245 110.735 187.435 ;
        RECT 117.005 187.265 117.175 187.455 ;
        RECT 119.765 187.245 119.935 187.435 ;
        RECT 126.665 187.265 126.835 187.455 ;
        RECT 127.125 187.265 127.295 187.455 ;
        RECT 128.970 187.245 129.140 187.435 ;
        RECT 130.810 187.245 130.980 187.435 ;
        RECT 134.485 187.265 134.655 187.435 ;
        RECT 138.160 187.265 138.330 187.455 ;
        RECT 134.485 187.245 134.685 187.265 ;
        RECT 139.545 187.245 139.715 187.455 ;
        RECT 44.620 187.215 45.555 187.245 ;
        RECT 42.490 187.015 45.555 187.215 ;
        RECT 37.290 186.335 38.655 186.565 ;
        RECT 41.405 186.335 42.335 186.565 ;
        RECT 42.345 186.535 45.555 187.015 ;
        RECT 45.565 186.565 48.315 187.245 ;
        RECT 42.345 186.335 43.275 186.535 ;
        RECT 44.605 186.335 45.555 186.535 ;
        RECT 47.385 186.335 48.315 186.565 ;
        RECT 49.445 186.425 51.375 187.245 ;
        RECT 51.545 186.435 52.915 187.245 ;
        RECT 49.445 186.335 50.395 186.425 ;
        RECT 52.935 186.375 53.365 187.160 ;
        RECT 53.525 186.335 56.975 187.245 ;
        RECT 57.065 186.435 62.575 187.245 ;
        RECT 62.585 186.435 65.335 187.245 ;
        RECT 65.365 186.335 66.715 187.245 ;
        RECT 66.725 186.435 68.555 187.245 ;
        RECT 68.565 186.565 72.235 187.245 ;
        RECT 71.310 186.335 72.235 186.565 ;
        RECT 72.245 186.335 75.720 187.245 ;
        RECT 76.235 186.565 78.070 187.245 ;
        RECT 76.235 186.335 77.165 186.565 ;
        RECT 78.695 186.375 79.125 187.160 ;
        RECT 79.145 186.335 80.495 187.245 ;
        RECT 80.540 186.335 82.355 187.245 ;
        RECT 82.380 186.335 84.195 187.245 ;
        RECT 84.220 186.335 86.035 187.245 ;
        RECT 86.185 186.565 89.715 187.245 ;
        RECT 86.890 186.335 89.715 186.565 ;
        RECT 90.645 186.335 91.995 187.245 ;
        RECT 92.025 186.335 94.775 187.245 ;
        RECT 94.785 186.335 97.995 187.245 ;
        RECT 98.155 186.335 101.810 187.245 ;
        RECT 102.605 186.335 104.420 187.245 ;
        RECT 104.455 186.375 104.885 187.160 ;
        RECT 104.905 186.335 106.255 187.245 ;
        RECT 106.285 186.565 109.815 187.245 ;
        RECT 110.425 186.565 119.530 187.245 ;
        RECT 119.625 186.565 128.730 187.245 ;
        RECT 106.285 186.335 109.110 186.565 ;
        RECT 128.825 186.335 130.175 187.245 ;
        RECT 130.215 186.375 130.645 187.160 ;
        RECT 130.665 186.335 134.265 187.245 ;
        RECT 134.485 186.565 138.015 187.245 ;
        RECT 135.190 186.335 138.015 186.565 ;
        RECT 138.485 186.435 139.855 187.245 ;
      LAYER nwell ;
        RECT 26.970 183.215 140.050 186.045 ;
      LAYER pwell ;
        RECT 31.995 182.835 33.585 182.925 ;
        RECT 27.165 182.015 28.535 182.825 ;
        RECT 28.545 182.015 30.375 182.695 ;
        RECT 31.015 182.015 33.585 182.835 ;
        RECT 33.605 182.015 39.115 182.825 ;
        RECT 40.055 182.100 40.485 182.885 ;
        RECT 43.270 182.695 44.610 182.925 ;
        RECT 45.305 182.835 46.255 182.925 ;
        RECT 40.505 182.015 45.095 182.695 ;
        RECT 45.305 182.015 47.235 182.835 ;
        RECT 47.715 182.695 48.645 182.925 ;
        RECT 47.715 182.015 49.550 182.695 ;
        RECT 27.305 181.805 27.475 182.015 ;
        RECT 28.685 181.825 28.855 182.015 ;
        RECT 31.015 181.995 31.155 182.015 ;
        RECT 30.065 181.805 30.235 181.995 ;
        RECT 30.520 181.960 30.640 181.965 ;
        RECT 30.520 181.855 30.695 181.960 ;
        RECT 30.535 181.850 30.695 181.855 ;
        RECT 30.985 181.825 31.155 181.995 ;
        RECT 32.365 181.805 32.535 181.995 ;
        RECT 32.825 181.805 32.995 181.995 ;
        RECT 33.745 181.825 33.915 182.015 ;
        RECT 38.345 181.805 38.515 181.995 ;
        RECT 39.275 181.860 39.435 181.970 ;
        RECT 42.020 181.855 42.140 181.965 ;
        RECT 43.865 181.805 44.035 181.995 ;
        RECT 44.780 181.825 44.950 182.015 ;
        RECT 47.085 181.995 47.235 182.015 ;
        RECT 49.385 181.995 49.550 182.015 ;
        RECT 49.855 182.015 53.510 182.925 ;
        RECT 53.845 182.015 57.055 182.925 ;
        RECT 57.065 182.015 59.815 182.825 ;
        RECT 61.670 182.695 63.035 182.925 ;
        RECT 59.825 182.015 63.035 182.695 ;
        RECT 63.045 182.015 65.795 182.825 ;
        RECT 65.815 182.100 66.245 182.885 ;
        RECT 66.265 182.015 69.935 182.825 ;
        RECT 70.405 182.015 73.325 182.925 ;
        RECT 74.545 182.725 75.475 182.925 ;
        RECT 76.810 182.725 77.755 182.925 ;
        RECT 74.545 182.245 77.755 182.725 ;
        RECT 74.685 182.045 77.755 182.245 ;
        RECT 49.855 181.995 50.015 182.015 ;
        RECT 47.085 181.825 47.265 181.995 ;
        RECT 47.095 181.805 47.265 181.825 ;
        RECT 47.545 181.805 47.715 181.995 ;
        RECT 49.385 181.825 49.555 181.995 ;
        RECT 49.845 181.825 50.015 181.995 ;
        RECT 50.305 181.805 50.475 181.995 ;
        RECT 52.155 181.850 52.315 181.960 ;
        RECT 53.975 181.825 54.145 182.015 ;
        RECT 57.205 181.995 57.375 182.015 ;
        RECT 56.740 181.805 56.910 181.995 ;
        RECT 57.205 181.825 57.380 181.995 ;
        RECT 59.970 181.825 60.140 182.015 ;
        RECT 57.210 181.805 57.380 181.825 ;
        RECT 63.185 181.805 63.355 182.015 ;
        RECT 63.645 181.805 63.815 181.995 ;
        RECT 65.025 181.805 65.195 181.995 ;
        RECT 66.405 181.825 66.575 182.015 ;
        RECT 66.865 181.805 67.035 181.995 ;
        RECT 70.085 181.965 70.255 181.995 ;
        RECT 69.620 181.855 69.740 181.965 ;
        RECT 70.080 181.855 70.255 181.965 ;
        RECT 70.085 181.805 70.255 181.855 ;
        RECT 70.550 181.825 70.720 182.015 ;
        RECT 71.465 181.805 71.635 181.995 ;
        RECT 73.300 181.855 73.420 181.965 ;
        RECT 73.775 181.860 73.935 181.970 ;
        RECT 74.685 181.805 74.855 182.045 ;
        RECT 76.810 182.015 77.755 182.045 ;
        RECT 77.765 182.015 80.545 182.925 ;
        RECT 80.985 182.015 82.815 182.695 ;
        RECT 82.825 182.015 84.195 182.795 ;
        RECT 84.205 182.695 87.030 182.925 ;
        RECT 84.205 182.015 87.735 182.695 ;
        RECT 76.055 181.805 76.225 181.995 ;
        RECT 76.985 181.845 77.155 181.995 ;
        RECT 27.165 180.995 28.535 181.805 ;
        RECT 28.545 181.125 30.375 181.805 ;
        RECT 28.545 180.895 29.890 181.125 ;
        RECT 31.305 181.025 32.675 181.805 ;
        RECT 32.685 180.995 38.195 181.805 ;
        RECT 38.205 180.995 41.875 181.805 ;
        RECT 42.345 181.125 44.175 181.805 ;
        RECT 42.345 180.895 43.690 181.125 ;
        RECT 44.185 180.895 47.395 181.805 ;
        RECT 47.415 180.895 50.145 181.805 ;
        RECT 50.165 181.125 51.995 181.805 ;
        RECT 50.650 180.895 51.995 181.125 ;
        RECT 52.935 180.935 53.365 181.720 ;
        RECT 53.385 180.895 57.055 181.805 ;
        RECT 57.210 181.575 60.265 181.805 ;
        RECT 57.065 180.895 60.265 181.575 ;
        RECT 60.285 180.895 63.495 181.805 ;
        RECT 63.505 180.995 64.875 181.805 ;
        RECT 64.885 181.125 66.715 181.805 ;
        RECT 65.370 180.895 66.715 181.125 ;
        RECT 66.725 180.995 69.475 181.805 ;
        RECT 69.955 180.895 71.305 181.805 ;
        RECT 71.325 180.995 73.155 181.805 ;
        RECT 73.635 180.895 74.985 181.805 ;
        RECT 75.005 181.025 76.375 181.805 ;
        RECT 76.385 180.895 77.275 181.845 ;
        RECT 77.455 181.805 77.625 181.995 ;
        RECT 77.905 181.825 78.075 182.015 ;
        RECT 79.290 181.805 79.460 181.995 ;
        RECT 81.125 181.825 81.295 182.015 ;
        RECT 82.975 181.825 83.145 182.015 ;
        RECT 87.535 181.995 87.735 182.015 ;
        RECT 83.895 181.850 84.055 181.960 ;
        RECT 85.725 181.805 85.895 181.995 ;
        RECT 86.185 181.805 86.355 181.995 ;
        RECT 87.565 181.825 87.745 181.995 ;
        RECT 87.885 181.975 88.775 182.925 ;
        RECT 88.805 182.015 90.175 182.795 ;
        RECT 90.185 182.015 91.535 182.925 ;
        RECT 91.575 182.100 92.005 182.885 ;
        RECT 92.485 182.015 95.695 182.925 ;
        RECT 96.625 182.695 97.545 182.925 ;
        RECT 96.625 182.015 100.210 182.695 ;
        RECT 101.225 182.015 104.700 182.925 ;
        RECT 104.905 182.015 114.010 182.695 ;
        RECT 114.105 182.015 117.145 182.925 ;
        RECT 117.335 182.100 117.765 182.885 ;
        RECT 118.705 182.015 121.915 182.925 ;
        RECT 122.010 182.015 131.115 182.695 ;
        RECT 131.125 182.015 138.035 182.925 ;
        RECT 138.485 182.015 139.855 182.825 ;
        RECT 88.485 181.825 88.655 181.975 ;
        RECT 88.955 181.825 89.125 182.015 ;
        RECT 91.250 181.995 91.420 182.015 ;
        RECT 87.575 181.805 87.745 181.825 ;
        RECT 89.860 181.805 90.030 181.995 ;
        RECT 91.245 181.825 91.420 181.995 ;
        RECT 92.160 181.855 92.280 181.965 ;
        RECT 91.245 181.805 91.415 181.825 ;
        RECT 92.625 181.805 92.795 181.995 ;
        RECT 93.090 181.805 93.260 181.995 ;
        RECT 95.385 181.825 95.555 182.015 ;
        RECT 95.855 181.850 96.015 181.970 ;
        RECT 96.770 181.825 96.940 182.015 ;
        RECT 99.065 181.805 99.235 181.995 ;
        RECT 100.455 181.860 100.615 181.970 ;
        RECT 101.370 181.825 101.540 182.015 ;
        RECT 102.285 181.805 102.455 181.995 ;
        RECT 102.745 181.805 102.915 181.995 ;
        RECT 105.045 181.965 105.215 182.015 ;
        RECT 117.000 181.995 117.145 182.015 ;
        RECT 105.040 181.855 105.215 181.965 ;
        RECT 105.045 181.825 105.215 181.855 ;
        RECT 114.245 181.805 114.415 181.995 ;
        RECT 117.000 181.825 117.170 181.995 ;
        RECT 117.935 181.860 118.095 181.970 ;
        RECT 121.600 181.825 121.770 182.015 ;
        RECT 123.445 181.805 123.615 181.995 ;
        RECT 127.580 181.805 127.750 181.995 ;
        RECT 129.880 181.805 130.050 181.995 ;
        RECT 130.805 181.965 130.975 182.015 ;
        RECT 130.800 181.855 130.975 181.965 ;
        RECT 130.805 181.825 130.975 181.855 ;
        RECT 131.265 181.995 131.435 182.015 ;
        RECT 131.265 181.825 131.440 181.995 ;
        RECT 131.270 181.805 131.440 181.825 ;
        RECT 138.160 181.805 138.330 181.995 ;
        RECT 139.545 181.805 139.715 182.015 ;
        RECT 77.305 181.025 78.675 181.805 ;
        RECT 78.695 180.935 79.125 181.720 ;
        RECT 79.145 180.895 83.535 181.805 ;
        RECT 84.675 180.895 86.025 181.805 ;
        RECT 86.045 181.025 87.415 181.805 ;
        RECT 87.425 181.025 88.795 181.805 ;
        RECT 88.825 180.895 90.175 181.805 ;
        RECT 90.195 180.895 91.545 181.805 ;
        RECT 91.575 180.895 92.925 181.805 ;
        RECT 92.945 180.895 95.695 181.805 ;
        RECT 96.635 181.125 99.375 181.805 ;
        RECT 99.385 180.895 102.595 181.805 ;
        RECT 102.605 181.125 104.435 181.805 ;
        RECT 103.090 180.895 104.435 181.125 ;
        RECT 104.455 180.935 104.885 181.720 ;
        RECT 105.450 181.125 114.555 181.805 ;
        RECT 114.650 181.125 123.755 181.805 ;
        RECT 123.765 180.895 127.895 181.805 ;
        RECT 127.985 180.895 130.195 181.805 ;
        RECT 130.215 180.935 130.645 181.720 ;
        RECT 131.125 180.895 134.670 181.805 ;
        RECT 134.930 180.895 138.475 181.805 ;
        RECT 138.485 180.995 139.855 181.805 ;
      LAYER nwell ;
        RECT 26.970 177.775 140.050 180.605 ;
      LAYER pwell ;
        RECT 27.165 176.575 28.535 177.385 ;
        RECT 28.545 176.575 34.055 177.385 ;
        RECT 34.065 176.575 39.575 177.385 ;
        RECT 40.055 176.660 40.485 177.445 ;
        RECT 42.810 177.255 44.175 177.485 ;
        RECT 40.965 176.575 44.175 177.255 ;
        RECT 44.645 176.575 47.395 177.485 ;
        RECT 47.405 176.575 52.915 177.385 ;
        RECT 52.925 176.575 54.755 177.385 ;
        RECT 55.225 176.805 57.060 177.485 ;
        RECT 55.370 176.575 57.060 176.805 ;
        RECT 57.525 176.575 60.275 177.385 ;
        RECT 60.765 176.575 62.115 177.485 ;
        RECT 62.125 176.575 65.795 177.485 ;
        RECT 65.815 176.660 66.245 177.445 ;
        RECT 66.265 176.575 69.935 177.485 ;
        RECT 69.965 176.575 71.315 177.485 ;
        RECT 27.305 176.365 27.475 176.575 ;
        RECT 28.685 176.365 28.855 176.575 ;
        RECT 34.205 176.365 34.375 176.575 ;
        RECT 39.725 176.525 39.895 176.555 ;
        RECT 39.720 176.415 39.895 176.525 ;
        RECT 40.640 176.415 40.760 176.525 ;
        RECT 39.725 176.365 39.895 176.415 ;
        RECT 41.110 176.385 41.280 176.575 ;
        RECT 41.565 176.365 41.735 176.555 ;
        RECT 44.320 176.415 44.440 176.525 ;
        RECT 44.785 176.385 44.955 176.575 ;
        RECT 45.705 176.365 45.875 176.555 ;
        RECT 46.165 176.365 46.335 176.555 ;
        RECT 47.545 176.385 47.715 176.575 ;
        RECT 49.385 176.385 49.555 176.555 ;
        RECT 49.385 176.365 49.535 176.385 ;
        RECT 51.225 176.365 51.395 176.555 ;
        RECT 51.685 176.365 51.855 176.555 ;
        RECT 53.065 176.385 53.235 176.575 ;
        RECT 53.525 176.365 53.695 176.555 ;
        RECT 54.900 176.415 55.020 176.525 ;
        RECT 55.370 176.385 55.540 176.575 ;
        RECT 57.665 176.385 57.835 176.575 ;
        RECT 59.040 176.365 59.210 176.555 ;
        RECT 60.420 176.365 60.590 176.555 ;
        RECT 61.800 176.385 61.970 176.575 ;
        RECT 62.720 176.365 62.890 176.555 ;
        RECT 65.025 176.385 65.195 176.555 ;
        RECT 65.485 176.525 65.655 176.575 ;
        RECT 65.480 176.415 65.655 176.525 ;
        RECT 65.485 176.385 65.655 176.415 ;
        RECT 65.025 176.365 65.190 176.385 ;
        RECT 65.955 176.365 66.125 176.555 ;
        RECT 69.625 176.365 69.795 176.575 ;
        RECT 71.000 176.555 71.170 176.575 ;
        RECT 70.080 176.415 70.200 176.525 ;
        RECT 71.000 176.405 71.175 176.555 ;
        RECT 27.165 175.555 28.535 176.365 ;
        RECT 28.545 175.555 34.055 176.365 ;
        RECT 34.065 175.555 39.575 176.365 ;
        RECT 39.585 175.555 41.415 176.365 ;
        RECT 41.425 175.685 44.175 176.365 ;
        RECT 44.185 175.685 46.015 176.365 ;
        RECT 43.245 175.455 44.175 175.685 ;
        RECT 46.025 175.555 47.395 176.365 ;
        RECT 47.605 175.545 49.535 176.365 ;
        RECT 49.705 175.685 51.535 176.365 ;
        RECT 51.545 175.555 52.915 176.365 ;
        RECT 47.605 175.455 48.555 175.545 ;
        RECT 52.935 175.495 53.365 176.280 ;
        RECT 53.385 175.555 58.895 176.365 ;
        RECT 58.925 175.455 60.275 176.365 ;
        RECT 60.305 175.455 61.655 176.365 ;
        RECT 61.685 175.455 63.035 176.365 ;
        RECT 63.355 175.685 65.190 176.365 ;
        RECT 63.355 175.455 64.285 175.685 ;
        RECT 65.805 175.585 67.175 176.365 ;
        RECT 67.195 175.455 69.925 176.365 ;
        RECT 70.405 175.455 71.295 176.405 ;
        RECT 71.475 176.365 71.645 176.555 ;
        RECT 72.385 176.385 72.555 176.555 ;
        RECT 72.705 176.535 73.595 177.485 ;
        RECT 73.625 176.575 74.995 177.355 ;
        RECT 75.015 176.575 77.745 177.485 ;
        RECT 77.780 176.575 79.595 177.485 ;
        RECT 80.525 176.575 81.895 177.355 ;
        RECT 81.925 176.575 83.275 177.485 ;
        RECT 83.285 176.575 86.495 177.485 ;
        RECT 86.965 176.575 88.335 177.355 ;
        RECT 88.345 176.575 89.715 177.355 ;
        RECT 89.725 176.575 91.540 177.485 ;
        RECT 91.575 176.660 92.005 177.445 ;
        RECT 92.945 176.805 94.780 177.485 ;
        RECT 93.090 176.575 94.780 176.805 ;
        RECT 95.255 177.395 96.845 177.485 ;
        RECT 95.255 176.575 97.825 177.395 ;
        RECT 98.295 176.575 101.215 177.485 ;
        RECT 101.240 176.575 104.895 177.485 ;
        RECT 104.990 176.575 114.095 177.255 ;
        RECT 114.105 176.575 117.315 177.485 ;
        RECT 117.335 176.660 117.765 177.445 ;
        RECT 117.840 176.575 121.915 177.485 ;
        RECT 122.385 176.575 131.490 177.255 ;
        RECT 131.595 176.805 134.795 177.485 ;
        RECT 135.650 177.255 138.475 177.485 ;
        RECT 131.595 176.575 134.650 176.805 ;
        RECT 72.845 176.365 73.015 176.535 ;
        RECT 73.305 176.385 73.475 176.535 ;
        RECT 73.765 176.385 73.935 176.575 ;
        RECT 74.225 176.405 74.395 176.555 ;
        RECT 75.145 176.525 75.315 176.575 ;
        RECT 75.140 176.415 75.315 176.525 ;
        RECT 71.325 175.585 72.695 176.365 ;
        RECT 72.705 175.585 74.075 176.365 ;
        RECT 74.105 175.455 74.995 176.405 ;
        RECT 75.145 176.385 75.315 176.415 ;
        RECT 75.610 176.335 75.780 176.555 ;
        RECT 77.905 176.385 78.075 176.575 ;
        RECT 81.585 176.555 81.755 176.575 ;
        RECT 78.360 176.415 78.480 176.525 ;
        RECT 79.285 176.365 79.455 176.555 ;
        RECT 79.755 176.420 79.915 176.530 ;
        RECT 81.585 176.385 81.765 176.555 ;
        RECT 82.040 176.385 82.210 176.575 ;
        RECT 83.415 176.555 83.585 176.575 ;
        RECT 82.960 176.415 83.080 176.525 ;
        RECT 83.415 176.385 83.605 176.555 ;
        RECT 81.595 176.365 81.765 176.385 ;
        RECT 83.435 176.365 83.605 176.385 ;
        RECT 84.810 176.365 84.980 176.555 ;
        RECT 86.640 176.415 86.760 176.525 ;
        RECT 88.025 176.385 88.195 176.575 ;
        RECT 88.485 176.385 88.655 176.575 ;
        RECT 89.865 176.365 90.035 176.555 ;
        RECT 91.245 176.385 91.415 176.575 ;
        RECT 92.160 176.530 92.330 176.555 ;
        RECT 92.160 176.420 92.335 176.530 ;
        RECT 92.160 176.365 92.330 176.420 ;
        RECT 93.090 176.385 93.260 176.575 ;
        RECT 97.685 176.555 97.825 176.575 ;
        RECT 94.460 176.365 94.630 176.555 ;
        RECT 96.760 176.365 96.930 176.555 ;
        RECT 97.230 176.365 97.400 176.555 ;
        RECT 97.685 176.385 97.855 176.555 ;
        RECT 100.455 176.410 100.615 176.520 ;
        RECT 100.900 176.385 101.070 176.575 ;
        RECT 101.370 176.365 101.540 176.555 ;
        RECT 104.580 176.385 104.750 176.575 ;
        RECT 105.045 176.365 105.215 176.555 ;
        RECT 107.810 176.365 107.980 176.555 ;
        RECT 111.485 176.365 111.655 176.555 ;
        RECT 113.785 176.385 113.955 176.575 ;
        RECT 117.000 176.385 117.170 176.575 ;
        RECT 117.900 176.385 118.070 176.575 ;
        RECT 122.060 176.415 122.180 176.525 ;
        RECT 122.525 176.385 122.695 176.575 ;
        RECT 129.425 176.365 129.595 176.555 ;
        RECT 129.880 176.415 130.000 176.525 ;
        RECT 130.810 176.365 130.980 176.555 ;
        RECT 134.480 176.385 134.650 176.575 ;
        RECT 134.945 176.575 138.475 177.255 ;
        RECT 138.485 176.575 139.855 177.385 ;
        RECT 134.945 176.555 135.145 176.575 ;
        RECT 134.945 176.385 135.115 176.555 ;
        RECT 135.860 176.415 135.980 176.525 ;
        RECT 136.330 176.365 136.500 176.555 ;
        RECT 139.545 176.365 139.715 176.575 ;
        RECT 77.270 176.335 78.215 176.365 ;
        RECT 75.465 175.655 78.215 176.335 ;
        RECT 77.270 175.455 78.215 175.655 ;
        RECT 78.695 175.495 79.125 176.280 ;
        RECT 79.145 175.685 81.435 176.365 ;
        RECT 80.515 175.455 81.435 175.685 ;
        RECT 81.445 175.585 82.815 176.365 ;
        RECT 83.285 175.585 84.655 176.365 ;
        RECT 84.665 175.455 88.320 176.365 ;
        RECT 88.345 175.455 90.160 176.365 ;
        RECT 90.200 175.685 92.475 176.365 ;
        RECT 90.200 175.455 91.570 175.685 ;
        RECT 92.565 175.455 94.775 176.365 ;
        RECT 94.865 175.455 97.075 176.365 ;
        RECT 97.230 176.135 100.285 176.365 ;
        RECT 97.085 175.455 100.285 176.135 ;
        RECT 101.225 175.455 104.145 176.365 ;
        RECT 104.455 175.495 104.885 176.280 ;
        RECT 104.905 175.685 107.645 176.365 ;
        RECT 107.665 175.455 111.335 176.365 ;
        RECT 111.345 175.685 120.450 176.365 ;
        RECT 120.630 175.685 129.735 176.365 ;
        RECT 130.215 175.495 130.645 176.280 ;
        RECT 130.665 175.455 135.620 176.365 ;
        RECT 136.185 175.455 138.475 176.365 ;
        RECT 138.485 175.555 139.855 176.365 ;
      LAYER nwell ;
        RECT 26.970 172.335 140.050 175.165 ;
      LAYER pwell ;
        RECT 27.165 171.135 28.535 171.945 ;
        RECT 28.545 171.135 34.055 171.945 ;
        RECT 34.065 171.135 39.575 171.945 ;
        RECT 40.055 171.220 40.485 172.005 ;
        RECT 40.505 171.135 46.015 171.945 ;
        RECT 46.025 171.135 51.535 171.945 ;
        RECT 51.545 171.135 57.055 171.945 ;
        RECT 57.065 171.135 58.435 171.945 ;
        RECT 58.455 171.135 61.185 172.045 ;
        RECT 61.205 171.135 63.020 172.045 ;
        RECT 63.965 171.135 65.780 172.045 ;
        RECT 65.815 171.220 66.245 172.005 ;
        RECT 66.265 171.135 69.475 172.045 ;
        RECT 69.485 171.135 72.695 172.045 ;
        RECT 74.535 171.815 75.455 172.045 ;
        RECT 73.165 171.135 75.455 171.815 ;
        RECT 75.465 171.135 78.675 172.045 ;
        RECT 80.020 171.845 80.975 172.045 ;
        RECT 78.695 171.165 80.975 171.845 ;
        RECT 27.305 170.925 27.475 171.135 ;
        RECT 28.685 170.945 28.855 171.135 ;
        RECT 29.605 170.945 29.775 171.115 ;
        RECT 30.065 170.925 30.235 171.115 ;
        RECT 34.205 170.945 34.375 171.135 ;
        RECT 35.585 170.925 35.755 171.115 ;
        RECT 39.720 170.975 39.840 171.085 ;
        RECT 40.645 170.945 40.815 171.135 ;
        RECT 41.105 170.925 41.275 171.115 ;
        RECT 46.165 170.945 46.335 171.135 ;
        RECT 46.625 170.925 46.795 171.115 ;
        RECT 51.685 170.945 51.855 171.135 ;
        RECT 52.155 170.970 52.315 171.080 ;
        RECT 53.525 170.925 53.695 171.115 ;
        RECT 56.285 170.925 56.455 171.115 ;
        RECT 56.750 170.925 56.920 171.115 ;
        RECT 57.205 170.945 57.375 171.135 ;
        RECT 60.885 171.085 61.055 171.135 ;
        RECT 60.880 170.975 61.055 171.085 ;
        RECT 60.885 170.945 61.055 170.975 ;
        RECT 61.345 170.925 61.515 171.115 ;
        RECT 62.725 170.945 62.895 171.135 ;
        RECT 63.195 170.980 63.355 171.090 ;
        RECT 65.485 170.945 65.655 171.135 ;
        RECT 27.165 170.115 28.535 170.925 ;
        RECT 29.925 170.115 35.435 170.925 ;
        RECT 35.445 170.115 40.955 170.925 ;
        RECT 40.965 170.115 46.475 170.925 ;
        RECT 46.485 170.115 51.995 170.925 ;
        RECT 52.935 170.055 53.365 170.840 ;
        RECT 53.385 170.115 54.755 170.925 ;
        RECT 54.765 170.245 56.595 170.925 ;
        RECT 56.605 170.245 60.700 170.925 ;
        RECT 61.205 170.245 63.035 170.925 ;
        RECT 54.765 170.015 56.110 170.245 ;
        RECT 57.090 170.015 60.700 170.245 ;
        RECT 61.690 170.015 63.035 170.245 ;
        RECT 63.050 170.695 66.210 170.925 ;
        RECT 67.320 170.695 67.490 171.115 ;
        RECT 69.165 170.945 69.335 171.135 ;
        RECT 71.460 170.925 71.630 171.115 ;
        RECT 71.935 170.970 72.095 171.080 ;
        RECT 72.385 170.945 72.555 171.135 ;
        RECT 72.845 171.085 73.015 171.115 ;
        RECT 72.840 170.975 73.015 171.085 ;
        RECT 72.845 170.925 73.015 170.975 ;
        RECT 73.305 170.945 73.475 171.135 ;
        RECT 74.225 170.925 74.395 171.115 ;
        RECT 76.525 170.925 76.695 171.115 ;
        RECT 78.365 170.945 78.535 171.135 ;
        RECT 78.820 170.945 78.990 171.165 ;
        RECT 80.020 171.135 80.975 171.165 ;
        RECT 81.115 171.135 84.115 172.045 ;
        RECT 84.345 171.135 87.795 172.045 ;
        RECT 89.220 171.845 90.175 172.045 ;
        RECT 87.895 171.165 90.175 171.845 ;
        RECT 82.505 170.925 82.675 171.115 ;
        RECT 82.965 170.925 83.135 171.115 ;
        RECT 83.885 170.945 84.055 171.135 ;
        RECT 84.805 170.925 84.975 171.115 ;
        RECT 87.565 170.945 87.735 171.135 ;
        RECT 88.020 170.945 88.190 171.165 ;
        RECT 89.220 171.135 90.175 171.165 ;
        RECT 90.195 171.135 91.545 172.045 ;
        RECT 91.575 171.220 92.005 172.005 ;
        RECT 92.035 171.135 94.970 172.045 ;
        RECT 95.705 171.815 96.635 172.045 ;
        RECT 98.465 171.815 99.600 172.045 ;
        RECT 95.705 171.135 98.455 171.815 ;
        RECT 98.465 171.135 101.675 171.815 ;
        RECT 101.685 171.135 110.790 171.815 ;
        RECT 110.885 171.135 116.955 172.045 ;
        RECT 117.335 171.220 117.765 172.005 ;
        RECT 137.235 171.815 138.165 172.045 ;
        RECT 117.785 171.135 126.890 171.815 ;
        RECT 126.985 171.135 136.090 171.815 ;
        RECT 136.330 171.135 138.165 171.815 ;
        RECT 138.485 171.135 139.855 171.945 ;
        RECT 88.485 170.945 88.655 171.115 ;
        RECT 88.485 170.925 88.635 170.945 ;
        RECT 88.950 170.925 89.120 171.115 ;
        RECT 91.245 170.945 91.415 171.135 ;
        RECT 94.925 171.115 94.970 171.135 ;
        RECT 94.925 170.945 95.095 171.115 ;
        RECT 95.380 170.975 95.500 171.085 ;
        RECT 96.305 170.945 96.475 171.115 ;
        RECT 96.765 170.945 96.935 171.115 ;
        RECT 98.145 170.945 98.315 171.135 ;
        RECT 101.365 170.945 101.535 171.135 ;
        RECT 101.825 170.945 101.995 171.135 ;
        RECT 111.030 171.115 111.200 171.135 ;
        RECT 96.305 170.925 96.350 170.945 ;
        RECT 63.050 170.245 67.595 170.695 ;
        RECT 63.050 170.015 64.430 170.245 ;
        RECT 66.220 170.015 67.595 170.245 ;
        RECT 67.680 170.245 71.775 170.925 ;
        RECT 67.680 170.015 71.290 170.245 ;
        RECT 72.705 170.145 74.075 170.925 ;
        RECT 74.085 170.245 76.375 170.925 ;
        RECT 76.385 170.245 78.675 170.925 ;
        RECT 75.455 170.015 76.375 170.245 ;
        RECT 77.755 170.015 78.675 170.245 ;
        RECT 78.695 170.055 79.125 170.840 ;
        RECT 79.285 170.015 82.735 170.925 ;
        RECT 82.825 170.245 84.655 170.925 ;
        RECT 84.665 170.245 86.495 170.925 ;
        RECT 86.705 170.105 88.635 170.925 ;
        RECT 88.805 170.245 93.395 170.925 ;
        RECT 86.705 170.015 87.655 170.105 ;
        RECT 89.290 170.015 90.630 170.245 ;
        RECT 93.415 170.015 96.350 170.925 ;
        RECT 96.795 170.925 96.935 170.945 ;
        RECT 102.740 170.925 102.910 171.115 ;
        RECT 103.205 170.925 103.375 171.115 ;
        RECT 107.800 170.925 107.970 171.115 ;
        RECT 108.265 170.925 108.435 171.115 ;
        RECT 111.025 170.945 111.200 171.115 ;
        RECT 117.925 170.945 118.095 171.135 ;
        RECT 127.125 170.945 127.295 171.135 ;
        RECT 136.330 171.115 136.495 171.135 ;
        RECT 111.025 170.925 111.195 170.945 ;
        RECT 128.965 170.925 129.135 171.115 ;
        RECT 129.435 170.970 129.595 171.080 ;
        RECT 130.805 170.945 130.975 171.115 ;
        RECT 134.485 170.945 134.655 171.115 ;
        RECT 136.325 170.945 136.495 171.115 ;
        RECT 138.160 170.975 138.280 171.085 ;
        RECT 130.805 170.925 131.005 170.945 ;
        RECT 134.485 170.925 134.685 170.945 ;
        RECT 139.545 170.925 139.715 171.135 ;
        RECT 96.795 170.105 99.365 170.925 ;
        RECT 97.775 170.015 99.365 170.105 ;
        RECT 99.465 170.015 103.050 170.925 ;
        RECT 103.065 170.145 104.435 170.925 ;
        RECT 104.455 170.055 104.885 170.840 ;
        RECT 104.915 170.695 107.970 170.925 ;
        RECT 104.915 170.015 108.115 170.695 ;
        RECT 108.125 170.245 110.865 170.925 ;
        RECT 110.885 170.245 119.990 170.925 ;
        RECT 120.170 170.245 129.275 170.925 ;
        RECT 130.215 170.055 130.645 170.840 ;
        RECT 130.805 170.245 134.335 170.925 ;
        RECT 134.485 170.245 138.015 170.925 ;
        RECT 131.510 170.015 134.335 170.245 ;
        RECT 135.190 170.015 138.015 170.245 ;
        RECT 138.485 170.115 139.855 170.925 ;
      LAYER nwell ;
        RECT 26.970 166.895 140.050 169.725 ;
      LAYER pwell ;
        RECT 27.165 165.695 28.535 166.505 ;
        RECT 28.545 165.695 34.055 166.505 ;
        RECT 34.065 165.695 39.575 166.505 ;
        RECT 40.055 165.780 40.485 166.565 ;
        RECT 41.425 165.695 42.795 166.475 ;
        RECT 42.805 165.695 44.635 166.505 ;
        RECT 44.645 165.695 46.015 166.475 ;
        RECT 46.025 165.695 47.855 166.505 ;
        RECT 48.350 166.375 49.695 166.605 ;
        RECT 47.865 165.695 49.695 166.375 ;
        RECT 50.165 165.695 51.535 166.475 ;
        RECT 51.545 165.695 52.915 166.475 ;
        RECT 52.935 165.780 53.365 166.565 ;
        RECT 54.305 165.695 55.675 166.475 ;
        RECT 55.720 166.375 57.095 166.605 ;
        RECT 58.865 166.375 59.815 166.605 ;
        RECT 55.720 165.925 59.815 166.375 ;
        RECT 27.305 165.505 27.475 165.695 ;
        RECT 28.685 165.505 28.855 165.695 ;
        RECT 34.205 165.505 34.375 165.695 ;
        RECT 39.720 165.535 39.840 165.645 ;
        RECT 40.655 165.540 40.815 165.650 ;
        RECT 41.575 165.505 41.745 165.695 ;
        RECT 42.945 165.505 43.115 165.695 ;
        RECT 44.785 165.505 44.955 165.695 ;
        RECT 46.165 165.505 46.335 165.695 ;
        RECT 48.005 165.505 48.175 165.695 ;
        RECT 49.840 165.535 49.960 165.645 ;
        RECT 50.315 165.505 50.485 165.695 ;
        RECT 51.695 165.505 51.865 165.695 ;
        RECT 53.535 165.540 53.695 165.650 ;
        RECT 54.455 165.505 54.625 165.695 ;
        RECT 55.825 165.505 55.995 165.925 ;
        RECT 57.105 165.695 59.815 165.925 ;
        RECT 59.825 166.375 61.170 166.605 ;
        RECT 59.825 165.695 61.655 166.375 ;
        RECT 61.665 165.695 63.495 166.375 ;
        RECT 64.425 165.695 65.795 166.475 ;
        RECT 65.815 165.780 66.245 166.565 ;
        RECT 66.265 166.375 67.610 166.605 ;
        RECT 66.265 165.695 68.095 166.375 ;
        RECT 69.025 165.695 70.395 166.475 ;
        RECT 70.405 165.695 71.775 166.475 ;
        RECT 71.805 165.695 73.155 166.605 ;
        RECT 73.165 165.695 74.535 166.475 ;
        RECT 74.545 165.695 75.915 166.475 ;
        RECT 75.925 165.695 77.295 166.475 ;
        RECT 77.305 165.695 78.675 166.475 ;
        RECT 78.695 165.780 79.125 166.565 ;
        RECT 80.550 166.375 81.895 166.605 ;
        RECT 80.065 165.695 81.895 166.375 ;
        RECT 81.905 166.375 83.250 166.605 ;
        RECT 81.905 165.695 83.735 166.375 ;
        RECT 83.745 165.925 85.580 166.605 ;
        RECT 83.890 165.695 85.580 165.925 ;
        RECT 86.055 165.695 88.785 166.605 ;
        RECT 88.805 166.405 90.215 166.605 ;
        RECT 88.805 165.725 91.540 166.405 ;
        RECT 91.575 165.780 92.005 166.565 ;
        RECT 101.695 166.515 103.285 166.605 ;
        RECT 88.805 165.695 90.200 165.725 ;
        RECT 61.345 165.505 61.515 165.695 ;
        RECT 61.805 165.505 61.975 165.695 ;
        RECT 63.655 165.540 63.815 165.650 ;
        RECT 64.575 165.505 64.745 165.695 ;
        RECT 67.785 165.505 67.955 165.695 ;
        RECT 68.255 165.540 68.415 165.650 ;
        RECT 69.165 165.505 69.335 165.695 ;
        RECT 70.555 165.505 70.725 165.695 ;
        RECT 72.840 165.505 73.010 165.695 ;
        RECT 73.315 165.505 73.485 165.695 ;
        RECT 74.695 165.505 74.865 165.695 ;
        RECT 76.075 165.505 76.245 165.695 ;
        RECT 77.455 165.505 77.625 165.695 ;
        RECT 79.295 165.540 79.455 165.650 ;
        RECT 80.205 165.505 80.375 165.695 ;
        RECT 83.425 165.505 83.595 165.695 ;
        RECT 83.890 165.505 84.060 165.695 ;
        RECT 88.485 165.505 88.655 165.695 ;
        RECT 91.245 165.505 91.415 165.725 ;
        RECT 92.570 165.695 101.675 166.375 ;
        RECT 101.695 165.695 104.265 166.515 ;
        RECT 104.455 165.780 104.885 166.565 ;
        RECT 104.905 165.695 107.945 166.605 ;
        RECT 108.125 165.695 111.335 166.605 ;
        RECT 111.345 165.695 114.555 166.605 ;
        RECT 114.575 165.695 117.315 166.375 ;
        RECT 117.335 165.780 117.765 166.565 ;
        RECT 118.270 166.375 119.615 166.605 ;
        RECT 117.785 165.695 119.615 166.375 ;
        RECT 119.625 165.695 128.730 166.375 ;
        RECT 128.825 165.695 130.195 166.475 ;
        RECT 130.215 165.780 130.645 166.565 ;
        RECT 130.865 166.515 131.815 166.605 ;
        RECT 130.865 165.695 132.795 166.515 ;
        RECT 133.810 166.375 136.635 166.605 ;
        RECT 137.130 166.375 138.475 166.605 ;
        RECT 92.160 165.535 92.280 165.645 ;
        RECT 101.365 165.505 101.535 165.695 ;
        RECT 104.125 165.675 104.265 165.695 ;
        RECT 107.800 165.675 107.945 165.695 ;
        RECT 104.125 165.505 104.295 165.675 ;
        RECT 107.800 165.505 107.970 165.675 ;
        RECT 108.265 165.505 108.435 165.695 ;
        RECT 111.485 165.505 111.655 165.695 ;
        RECT 117.005 165.505 117.175 165.695 ;
        RECT 117.925 165.505 118.095 165.695 ;
        RECT 119.765 165.505 119.935 165.695 ;
        RECT 129.875 165.505 130.045 165.695 ;
        RECT 132.645 165.675 132.795 165.695 ;
        RECT 133.105 165.695 136.635 166.375 ;
        RECT 136.645 165.695 138.475 166.375 ;
        RECT 138.485 165.695 139.855 166.505 ;
        RECT 133.105 165.675 133.305 165.695 ;
        RECT 132.645 165.505 132.815 165.675 ;
        RECT 133.105 165.505 133.275 165.675 ;
        RECT 136.785 165.505 136.955 165.695 ;
        RECT 139.545 165.505 139.715 165.695 ;
      LAYER li1 ;
        RECT 27.160 209.025 139.860 209.195 ;
        RECT 27.245 208.275 28.455 209.025 ;
        RECT 27.245 207.735 27.765 208.275 ;
        RECT 28.630 208.185 28.890 209.025 ;
        RECT 29.065 208.280 29.320 208.855 ;
        RECT 29.490 208.645 29.820 209.025 ;
        RECT 30.035 208.475 30.205 208.855 ;
        RECT 29.490 208.305 30.205 208.475 ;
        RECT 30.645 208.365 30.985 209.025 ;
        RECT 27.935 207.565 28.455 208.105 ;
        RECT 27.245 206.475 28.455 207.565 ;
        RECT 28.630 206.475 28.890 207.625 ;
        RECT 29.065 207.550 29.235 208.280 ;
        RECT 29.490 208.115 29.660 208.305 ;
        RECT 29.405 207.785 29.660 208.115 ;
        RECT 29.490 207.575 29.660 207.785 ;
        RECT 29.940 207.755 30.295 208.125 ;
        RECT 29.065 206.645 29.320 207.550 ;
        RECT 29.490 207.405 30.205 207.575 ;
        RECT 29.490 206.475 29.820 207.235 ;
        RECT 30.035 206.645 30.205 207.405 ;
        RECT 30.465 206.645 30.985 208.195 ;
        RECT 31.155 207.370 31.675 208.855 ;
        RECT 31.845 208.480 37.190 209.025 ;
        RECT 33.430 207.650 33.770 208.480 ;
        RECT 37.365 208.255 39.955 209.025 ;
        RECT 40.125 208.300 40.415 209.025 ;
        RECT 40.585 208.480 45.930 209.025 ;
        RECT 46.105 208.480 51.450 209.025 ;
        RECT 31.155 206.475 31.485 207.200 ;
        RECT 35.250 206.910 35.600 208.160 ;
        RECT 37.365 207.735 38.575 208.255 ;
        RECT 38.745 207.565 39.955 208.085 ;
        RECT 42.170 207.650 42.510 208.480 ;
        RECT 31.845 206.475 37.190 206.910 ;
        RECT 37.365 206.475 39.955 207.565 ;
        RECT 40.125 206.475 40.415 207.640 ;
        RECT 43.990 206.910 44.340 208.160 ;
        RECT 47.690 207.650 48.030 208.480 ;
        RECT 51.625 208.275 52.835 209.025 ;
        RECT 53.005 208.300 53.295 209.025 ;
        RECT 53.465 208.275 54.675 209.025 ;
        RECT 54.850 208.285 55.105 208.855 ;
        RECT 55.275 208.625 55.605 209.025 ;
        RECT 56.030 208.490 56.560 208.855 ;
        RECT 56.030 208.455 56.205 208.490 ;
        RECT 55.275 208.285 56.205 208.455 ;
        RECT 49.510 206.910 49.860 208.160 ;
        RECT 51.625 207.735 52.145 208.275 ;
        RECT 52.315 207.565 52.835 208.105 ;
        RECT 53.465 207.735 53.985 208.275 ;
        RECT 40.585 206.475 45.930 206.910 ;
        RECT 46.105 206.475 51.450 206.910 ;
        RECT 51.625 206.475 52.835 207.565 ;
        RECT 53.005 206.475 53.295 207.640 ;
        RECT 54.155 207.565 54.675 208.105 ;
        RECT 53.465 206.475 54.675 207.565 ;
        RECT 54.850 207.615 55.020 208.285 ;
        RECT 55.275 208.115 55.445 208.285 ;
        RECT 55.190 207.785 55.445 208.115 ;
        RECT 55.670 207.785 55.865 208.115 ;
        RECT 54.850 206.645 55.185 207.615 ;
        RECT 55.355 206.475 55.525 207.615 ;
        RECT 55.695 206.815 55.865 207.785 ;
        RECT 56.035 207.155 56.205 208.285 ;
        RECT 56.375 207.495 56.545 208.295 ;
        RECT 56.750 208.005 57.025 208.855 ;
        RECT 56.745 207.835 57.025 208.005 ;
        RECT 56.750 207.695 57.025 207.835 ;
        RECT 57.195 207.495 57.385 208.855 ;
        RECT 57.565 208.490 58.075 209.025 ;
        RECT 58.295 208.215 58.540 208.820 ;
        RECT 58.985 208.480 64.330 209.025 ;
        RECT 57.585 208.045 58.815 208.215 ;
        RECT 56.375 207.325 57.385 207.495 ;
        RECT 57.555 207.480 58.305 207.670 ;
        RECT 56.035 206.985 57.160 207.155 ;
        RECT 57.555 206.815 57.725 207.480 ;
        RECT 58.475 207.235 58.815 208.045 ;
        RECT 60.570 207.650 60.910 208.480 ;
        RECT 64.505 208.275 65.715 209.025 ;
        RECT 65.885 208.300 66.175 209.025 ;
        RECT 67.355 208.475 67.525 208.855 ;
        RECT 67.705 208.645 68.035 209.025 ;
        RECT 67.355 208.305 68.020 208.475 ;
        RECT 68.215 208.350 68.475 208.855 ;
        RECT 68.645 208.480 73.990 209.025 ;
        RECT 55.695 206.645 57.725 206.815 ;
        RECT 57.895 206.475 58.065 207.235 ;
        RECT 58.300 206.825 58.815 207.235 ;
        RECT 62.390 206.910 62.740 208.160 ;
        RECT 64.505 207.735 65.025 208.275 ;
        RECT 65.195 207.565 65.715 208.105 ;
        RECT 67.285 207.755 67.615 208.125 ;
        RECT 67.850 208.050 68.020 208.305 ;
        RECT 67.850 207.720 68.135 208.050 ;
        RECT 58.985 206.475 64.330 206.910 ;
        RECT 64.505 206.475 65.715 207.565 ;
        RECT 65.885 206.475 66.175 207.640 ;
        RECT 67.850 207.575 68.020 207.720 ;
        RECT 67.355 207.405 68.020 207.575 ;
        RECT 68.305 207.550 68.475 208.350 ;
        RECT 70.230 207.650 70.570 208.480 ;
        RECT 74.625 208.285 74.965 208.855 ;
        RECT 75.160 208.360 75.330 209.025 ;
        RECT 75.610 208.685 75.830 208.730 ;
        RECT 75.605 208.515 75.830 208.685 ;
        RECT 76.000 208.545 76.445 208.715 ;
        RECT 75.610 208.375 75.830 208.515 ;
        RECT 67.355 206.645 67.525 207.405 ;
        RECT 67.705 206.475 68.035 207.235 ;
        RECT 68.205 206.645 68.475 207.550 ;
        RECT 72.050 206.910 72.400 208.160 ;
        RECT 74.625 207.315 74.800 208.285 ;
        RECT 75.610 208.205 76.105 208.375 ;
        RECT 74.970 207.665 75.140 208.115 ;
        RECT 75.310 207.835 75.760 208.035 ;
        RECT 75.930 208.010 76.105 208.205 ;
        RECT 76.275 207.755 76.445 208.545 ;
        RECT 76.615 208.420 76.865 208.790 ;
        RECT 76.695 208.035 76.865 208.420 ;
        RECT 77.035 208.385 77.285 208.790 ;
        RECT 77.455 208.555 77.625 209.025 ;
        RECT 77.795 208.385 78.135 208.790 ;
        RECT 77.035 208.205 78.135 208.385 ;
        RECT 78.765 208.300 79.055 209.025 ;
        RECT 79.225 208.255 80.895 209.025 ;
        RECT 81.615 208.475 81.785 208.855 ;
        RECT 81.965 208.645 82.295 209.025 ;
        RECT 81.615 208.305 82.280 208.475 ;
        RECT 82.475 208.350 82.735 208.855 ;
        RECT 76.695 207.865 76.890 208.035 ;
        RECT 74.970 207.495 75.365 207.665 ;
        RECT 76.275 207.615 76.550 207.755 ;
        RECT 68.645 206.475 73.990 206.910 ;
        RECT 74.625 206.645 74.885 207.315 ;
        RECT 75.195 207.225 75.365 207.495 ;
        RECT 75.535 207.395 76.550 207.615 ;
        RECT 76.720 207.615 76.890 207.865 ;
        RECT 77.060 207.785 77.620 208.035 ;
        RECT 76.720 207.225 77.275 207.615 ;
        RECT 75.195 207.055 77.275 207.225 ;
        RECT 75.055 206.475 75.385 206.875 ;
        RECT 76.255 206.475 76.655 206.875 ;
        RECT 76.945 206.820 77.275 207.055 ;
        RECT 77.445 206.685 77.620 207.785 ;
        RECT 77.790 207.465 78.135 208.035 ;
        RECT 79.225 207.735 79.975 208.255 ;
        RECT 77.790 206.475 78.135 207.295 ;
        RECT 78.765 206.475 79.055 207.640 ;
        RECT 80.145 207.565 80.895 208.085 ;
        RECT 81.545 207.755 81.885 208.125 ;
        RECT 82.110 208.050 82.280 208.305 ;
        RECT 82.110 207.720 82.385 208.050 ;
        RECT 82.110 207.575 82.280 207.720 ;
        RECT 79.225 206.475 80.895 207.565 ;
        RECT 81.605 207.405 82.280 207.575 ;
        RECT 82.555 207.550 82.735 208.350 ;
        RECT 81.605 206.645 81.785 207.405 ;
        RECT 81.965 206.475 82.295 207.235 ;
        RECT 82.465 206.645 82.735 207.550 ;
        RECT 82.905 206.645 83.655 208.855 ;
        RECT 83.825 208.350 84.085 208.855 ;
        RECT 84.265 208.645 84.595 209.025 ;
        RECT 84.775 208.475 84.945 208.855 ;
        RECT 83.825 207.550 84.005 208.350 ;
        RECT 84.280 208.305 84.945 208.475 ;
        RECT 85.295 208.475 85.465 208.855 ;
        RECT 85.645 208.645 85.975 209.025 ;
        RECT 85.295 208.305 85.960 208.475 ;
        RECT 86.155 208.350 86.415 208.855 ;
        RECT 84.280 208.050 84.450 208.305 ;
        RECT 84.175 207.720 84.450 208.050 ;
        RECT 84.675 207.755 85.015 208.125 ;
        RECT 85.225 207.755 85.555 208.125 ;
        RECT 85.790 208.050 85.960 208.305 ;
        RECT 84.280 207.575 84.450 207.720 ;
        RECT 85.790 207.720 86.075 208.050 ;
        RECT 85.790 207.575 85.960 207.720 ;
        RECT 83.825 206.645 84.095 207.550 ;
        RECT 84.280 207.405 84.955 207.575 ;
        RECT 84.265 206.475 84.595 207.235 ;
        RECT 84.775 206.645 84.955 207.405 ;
        RECT 85.295 207.405 85.960 207.575 ;
        RECT 86.245 207.550 86.415 208.350 ;
        RECT 85.295 206.645 85.465 207.405 ;
        RECT 85.645 206.475 85.975 207.235 ;
        RECT 86.145 206.645 86.415 207.550 ;
        RECT 86.585 206.645 87.335 208.855 ;
        RECT 88.515 208.475 88.685 208.855 ;
        RECT 88.865 208.645 89.195 209.025 ;
        RECT 88.515 208.305 89.180 208.475 ;
        RECT 89.375 208.350 89.635 208.855 ;
        RECT 88.445 207.755 88.785 208.125 ;
        RECT 89.010 208.050 89.180 208.305 ;
        RECT 89.010 207.720 89.285 208.050 ;
        RECT 89.010 207.575 89.180 207.720 ;
        RECT 88.505 207.405 89.180 207.575 ;
        RECT 89.455 207.550 89.635 208.350 ;
        RECT 89.810 208.185 90.070 209.025 ;
        RECT 90.245 208.280 90.500 208.855 ;
        RECT 90.670 208.645 91.000 209.025 ;
        RECT 91.215 208.475 91.385 208.855 ;
        RECT 90.670 208.305 91.385 208.475 ;
        RECT 88.505 206.645 88.685 207.405 ;
        RECT 88.865 206.475 89.195 207.235 ;
        RECT 89.365 206.645 89.635 207.550 ;
        RECT 89.810 206.475 90.070 207.625 ;
        RECT 90.245 207.550 90.415 208.280 ;
        RECT 90.670 208.115 90.840 208.305 ;
        RECT 91.645 208.300 91.935 209.025 ;
        RECT 92.655 208.475 92.825 208.855 ;
        RECT 93.005 208.645 93.335 209.025 ;
        RECT 92.655 208.305 93.320 208.475 ;
        RECT 93.515 208.350 93.775 208.855 ;
        RECT 90.585 207.785 90.840 208.115 ;
        RECT 90.670 207.575 90.840 207.785 ;
        RECT 91.120 207.755 91.475 208.125 ;
        RECT 92.585 207.755 92.925 208.125 ;
        RECT 93.150 208.050 93.320 208.305 ;
        RECT 93.150 207.720 93.425 208.050 ;
        RECT 90.245 206.645 90.500 207.550 ;
        RECT 90.670 207.405 91.385 207.575 ;
        RECT 90.670 206.475 91.000 207.235 ;
        RECT 91.215 206.645 91.385 207.405 ;
        RECT 91.645 206.475 91.935 207.640 ;
        RECT 93.150 207.575 93.320 207.720 ;
        RECT 92.645 207.405 93.320 207.575 ;
        RECT 93.595 207.550 93.775 208.350 ;
        RECT 92.645 206.645 92.825 207.405 ;
        RECT 93.005 206.475 93.335 207.235 ;
        RECT 93.505 206.645 93.775 207.550 ;
        RECT 94.900 208.285 95.515 208.855 ;
        RECT 95.685 208.515 95.900 209.025 ;
        RECT 96.130 208.515 96.410 208.845 ;
        RECT 96.590 208.515 96.830 209.025 ;
        RECT 94.900 207.265 95.215 208.285 ;
        RECT 95.385 207.615 95.555 208.115 ;
        RECT 95.805 207.785 96.070 208.345 ;
        RECT 96.240 207.615 96.410 208.515 ;
        RECT 97.255 208.475 97.425 208.855 ;
        RECT 97.640 208.645 97.970 209.025 ;
        RECT 96.580 207.785 96.935 208.345 ;
        RECT 97.255 208.305 97.970 208.475 ;
        RECT 97.165 207.755 97.520 208.125 ;
        RECT 97.800 208.115 97.970 208.305 ;
        RECT 98.140 208.280 98.395 208.855 ;
        RECT 97.800 207.785 98.055 208.115 ;
        RECT 95.385 207.445 96.810 207.615 ;
        RECT 97.800 207.575 97.970 207.785 ;
        RECT 94.900 206.645 95.435 207.265 ;
        RECT 95.605 206.475 95.935 207.275 ;
        RECT 96.420 207.270 96.810 207.445 ;
        RECT 97.255 207.405 97.970 207.575 ;
        RECT 98.225 207.550 98.395 208.280 ;
        RECT 98.570 208.185 98.830 209.025 ;
        RECT 99.465 208.455 99.900 208.855 ;
        RECT 100.070 208.625 100.455 209.025 ;
        RECT 99.465 208.285 100.455 208.455 ;
        RECT 100.625 208.285 101.050 208.855 ;
        RECT 101.240 208.455 101.495 208.855 ;
        RECT 101.665 208.625 102.050 209.025 ;
        RECT 101.240 208.285 102.050 208.455 ;
        RECT 102.220 208.285 102.465 208.855 ;
        RECT 102.655 208.455 102.910 208.855 ;
        RECT 103.080 208.625 103.465 209.025 ;
        RECT 102.655 208.285 103.465 208.455 ;
        RECT 103.635 208.285 103.895 208.855 ;
        RECT 104.525 208.300 104.815 209.025 ;
        RECT 100.120 208.115 100.455 208.285 ;
        RECT 100.700 208.115 101.050 208.285 ;
        RECT 101.700 208.115 102.050 208.285 ;
        RECT 102.295 208.115 102.465 208.285 ;
        RECT 103.115 208.115 103.465 208.285 ;
        RECT 97.255 206.645 97.425 207.405 ;
        RECT 97.640 206.475 97.970 207.235 ;
        RECT 98.140 206.645 98.395 207.550 ;
        RECT 98.570 206.475 98.830 207.625 ;
        RECT 99.465 207.410 99.950 208.115 ;
        RECT 100.120 207.785 100.530 208.115 ;
        RECT 100.120 207.240 100.455 207.785 ;
        RECT 100.700 207.615 101.530 208.115 ;
        RECT 99.465 207.070 100.455 207.240 ;
        RECT 100.625 207.435 101.530 207.615 ;
        RECT 101.700 207.785 102.125 208.115 ;
        RECT 99.465 206.645 99.900 207.070 ;
        RECT 100.070 206.475 100.455 206.900 ;
        RECT 100.625 206.645 101.050 207.435 ;
        RECT 101.700 207.265 102.050 207.785 ;
        RECT 102.295 207.615 102.945 208.115 ;
        RECT 101.220 207.070 102.050 207.265 ;
        RECT 102.220 207.435 102.945 207.615 ;
        RECT 103.115 207.785 103.540 208.115 ;
        RECT 101.220 206.645 101.495 207.070 ;
        RECT 101.665 206.475 102.050 206.900 ;
        RECT 102.220 206.645 102.465 207.435 ;
        RECT 103.115 207.265 103.465 207.785 ;
        RECT 103.710 207.615 103.895 208.285 ;
        RECT 105.910 208.185 106.170 209.025 ;
        RECT 106.345 208.280 106.600 208.855 ;
        RECT 106.770 208.645 107.100 209.025 ;
        RECT 107.315 208.475 107.485 208.855 ;
        RECT 106.770 208.305 107.485 208.475 ;
        RECT 102.655 207.070 103.465 207.265 ;
        RECT 102.655 206.645 102.910 207.070 ;
        RECT 103.080 206.475 103.465 206.900 ;
        RECT 103.635 206.645 103.895 207.615 ;
        RECT 104.525 206.475 104.815 207.640 ;
        RECT 105.910 206.475 106.170 207.625 ;
        RECT 106.345 207.550 106.515 208.280 ;
        RECT 106.770 208.115 106.940 208.305 ;
        RECT 107.785 208.205 108.015 209.025 ;
        RECT 108.185 208.225 108.515 208.855 ;
        RECT 106.685 207.785 106.940 208.115 ;
        RECT 106.770 207.575 106.940 207.785 ;
        RECT 107.220 207.755 107.575 208.125 ;
        RECT 107.765 207.785 108.095 208.035 ;
        RECT 108.265 207.625 108.515 208.225 ;
        RECT 108.685 208.205 108.895 209.025 ;
        RECT 109.125 208.350 109.385 208.855 ;
        RECT 109.565 208.645 109.895 209.025 ;
        RECT 110.075 208.475 110.245 208.855 ;
        RECT 106.345 206.645 106.600 207.550 ;
        RECT 106.770 207.405 107.485 207.575 ;
        RECT 106.770 206.475 107.100 207.235 ;
        RECT 107.315 206.645 107.485 207.405 ;
        RECT 107.785 206.475 108.015 207.615 ;
        RECT 108.185 206.645 108.515 207.625 ;
        RECT 108.685 206.475 108.895 207.615 ;
        RECT 109.125 207.550 109.305 208.350 ;
        RECT 109.580 208.305 110.245 208.475 ;
        RECT 110.505 208.350 110.765 208.855 ;
        RECT 110.945 208.645 111.275 209.025 ;
        RECT 111.455 208.475 111.625 208.855 ;
        RECT 109.580 208.050 109.750 208.305 ;
        RECT 109.475 207.720 109.750 208.050 ;
        RECT 109.975 207.755 110.315 208.125 ;
        RECT 109.580 207.575 109.750 207.720 ;
        RECT 109.125 206.645 109.395 207.550 ;
        RECT 109.580 207.405 110.255 207.575 ;
        RECT 109.565 206.475 109.895 207.235 ;
        RECT 110.075 206.645 110.255 207.405 ;
        RECT 110.505 207.550 110.675 208.350 ;
        RECT 110.960 208.305 111.625 208.475 ;
        RECT 110.960 208.050 111.130 208.305 ;
        RECT 112.350 208.185 112.610 209.025 ;
        RECT 112.785 208.280 113.040 208.855 ;
        RECT 113.210 208.645 113.540 209.025 ;
        RECT 113.755 208.475 113.925 208.855 ;
        RECT 113.210 208.305 113.925 208.475 ;
        RECT 110.845 207.720 111.130 208.050 ;
        RECT 111.365 207.755 111.695 208.125 ;
        RECT 110.960 207.575 111.130 207.720 ;
        RECT 110.505 206.645 110.775 207.550 ;
        RECT 110.960 207.405 111.625 207.575 ;
        RECT 110.945 206.475 111.275 207.235 ;
        RECT 111.455 206.645 111.625 207.405 ;
        RECT 112.350 206.475 112.610 207.625 ;
        RECT 112.785 207.550 112.955 208.280 ;
        RECT 113.210 208.115 113.380 208.305 ;
        RECT 114.195 208.215 114.465 209.025 ;
        RECT 114.635 208.215 114.965 208.855 ;
        RECT 115.135 208.215 115.375 209.025 ;
        RECT 113.125 207.785 113.380 208.115 ;
        RECT 113.210 207.575 113.380 207.785 ;
        RECT 113.660 207.755 114.015 208.125 ;
        RECT 114.185 207.785 114.535 208.035 ;
        RECT 114.705 207.615 114.875 208.215 ;
        RECT 115.570 208.185 115.830 209.025 ;
        RECT 116.005 208.280 116.260 208.855 ;
        RECT 116.430 208.645 116.760 209.025 ;
        RECT 116.975 208.475 117.145 208.855 ;
        RECT 116.430 208.305 117.145 208.475 ;
        RECT 115.045 207.785 115.395 208.035 ;
        RECT 112.785 206.645 113.040 207.550 ;
        RECT 113.210 207.405 113.925 207.575 ;
        RECT 113.210 206.475 113.540 207.235 ;
        RECT 113.755 206.645 113.925 207.405 ;
        RECT 114.195 206.475 114.525 207.615 ;
        RECT 114.705 207.445 115.385 207.615 ;
        RECT 115.055 206.660 115.385 207.445 ;
        RECT 115.570 206.475 115.830 207.625 ;
        RECT 116.005 207.550 116.175 208.280 ;
        RECT 116.430 208.115 116.600 208.305 ;
        RECT 117.405 208.300 117.695 209.025 ;
        RECT 118.790 208.185 119.050 209.025 ;
        RECT 119.225 208.280 119.480 208.855 ;
        RECT 119.650 208.645 119.980 209.025 ;
        RECT 120.195 208.475 120.365 208.855 ;
        RECT 119.650 208.305 120.365 208.475 ;
        RECT 120.625 208.350 120.885 208.855 ;
        RECT 121.065 208.645 121.395 209.025 ;
        RECT 121.575 208.475 121.745 208.855 ;
        RECT 116.345 207.785 116.600 208.115 ;
        RECT 116.430 207.575 116.600 207.785 ;
        RECT 116.880 207.755 117.235 208.125 ;
        RECT 116.005 206.645 116.260 207.550 ;
        RECT 116.430 207.405 117.145 207.575 ;
        RECT 116.430 206.475 116.760 207.235 ;
        RECT 116.975 206.645 117.145 207.405 ;
        RECT 117.405 206.475 117.695 207.640 ;
        RECT 118.790 206.475 119.050 207.625 ;
        RECT 119.225 207.550 119.395 208.280 ;
        RECT 119.650 208.115 119.820 208.305 ;
        RECT 119.565 207.785 119.820 208.115 ;
        RECT 119.650 207.575 119.820 207.785 ;
        RECT 120.100 207.755 120.455 208.125 ;
        RECT 119.225 206.645 119.480 207.550 ;
        RECT 119.650 207.405 120.365 207.575 ;
        RECT 119.650 206.475 119.980 207.235 ;
        RECT 120.195 206.645 120.365 207.405 ;
        RECT 120.625 207.550 120.795 208.350 ;
        RECT 121.080 208.305 121.745 208.475 ;
        RECT 121.080 208.050 121.250 208.305 ;
        RECT 122.005 208.255 125.515 209.025 ;
        RECT 125.775 208.475 125.945 208.855 ;
        RECT 126.125 208.645 126.455 209.025 ;
        RECT 125.775 208.305 126.440 208.475 ;
        RECT 126.635 208.350 126.895 208.855 ;
        RECT 120.965 207.720 121.250 208.050 ;
        RECT 121.485 207.755 121.815 208.125 ;
        RECT 122.005 207.735 123.655 208.255 ;
        RECT 121.080 207.575 121.250 207.720 ;
        RECT 120.625 206.645 120.895 207.550 ;
        RECT 121.080 207.405 121.745 207.575 ;
        RECT 123.825 207.565 125.515 208.085 ;
        RECT 125.705 207.755 126.045 208.125 ;
        RECT 126.270 208.050 126.440 208.305 ;
        RECT 126.270 207.720 126.545 208.050 ;
        RECT 126.270 207.575 126.440 207.720 ;
        RECT 121.065 206.475 121.395 207.235 ;
        RECT 121.575 206.645 121.745 207.405 ;
        RECT 122.005 206.475 125.515 207.565 ;
        RECT 125.765 207.405 126.440 207.575 ;
        RECT 126.715 207.550 126.895 208.350 ;
        RECT 127.155 208.475 127.325 208.855 ;
        RECT 127.505 208.645 127.835 209.025 ;
        RECT 127.155 208.305 127.820 208.475 ;
        RECT 128.015 208.350 128.275 208.855 ;
        RECT 127.085 207.755 127.415 208.125 ;
        RECT 127.650 208.050 127.820 208.305 ;
        RECT 127.650 207.720 127.935 208.050 ;
        RECT 127.650 207.575 127.820 207.720 ;
        RECT 125.765 206.645 125.945 207.405 ;
        RECT 126.125 206.475 126.455 207.235 ;
        RECT 126.625 206.645 126.895 207.550 ;
        RECT 127.155 207.405 127.820 207.575 ;
        RECT 128.105 207.550 128.275 208.350 ;
        RECT 128.535 208.475 128.705 208.855 ;
        RECT 128.920 208.645 129.250 209.025 ;
        RECT 128.535 208.305 129.250 208.475 ;
        RECT 128.445 207.755 128.800 208.125 ;
        RECT 129.080 208.115 129.250 208.305 ;
        RECT 129.420 208.280 129.675 208.855 ;
        RECT 129.080 207.785 129.335 208.115 ;
        RECT 129.080 207.575 129.250 207.785 ;
        RECT 127.155 206.645 127.325 207.405 ;
        RECT 127.505 206.475 127.835 207.235 ;
        RECT 128.005 206.645 128.275 207.550 ;
        RECT 128.535 207.405 129.250 207.575 ;
        RECT 129.505 207.550 129.675 208.280 ;
        RECT 129.850 208.185 130.110 209.025 ;
        RECT 130.285 208.300 130.575 209.025 ;
        RECT 131.295 208.375 131.465 208.855 ;
        RECT 131.635 208.545 131.965 209.025 ;
        RECT 132.135 208.375 132.305 208.850 ;
        RECT 132.475 208.545 132.805 209.025 ;
        RECT 132.975 208.375 133.145 208.855 ;
        RECT 133.315 208.545 133.645 209.025 ;
        RECT 133.815 208.375 133.985 208.855 ;
        RECT 134.155 208.545 134.485 209.025 ;
        RECT 134.655 208.375 134.825 208.855 ;
        RECT 134.995 208.545 135.325 209.025 ;
        RECT 135.495 208.375 135.665 208.855 ;
        RECT 131.295 208.205 132.715 208.375 ;
        RECT 132.975 208.205 135.665 208.375 ;
        RECT 135.835 208.225 136.165 209.025 ;
        RECT 136.725 208.350 136.985 208.855 ;
        RECT 137.165 208.645 137.495 209.025 ;
        RECT 137.675 208.475 137.845 208.855 ;
        RECT 132.540 208.035 132.715 208.205 ;
        RECT 131.260 207.835 132.360 208.035 ;
        RECT 132.540 207.865 135.165 208.035 ;
        RECT 132.540 207.665 132.715 207.865 ;
        RECT 135.410 207.665 135.665 208.205 ;
        RECT 128.535 206.645 128.705 207.405 ;
        RECT 128.920 206.475 129.250 207.235 ;
        RECT 129.420 206.645 129.675 207.550 ;
        RECT 129.850 206.475 130.110 207.625 ;
        RECT 130.285 206.475 130.575 207.640 ;
        RECT 131.215 207.495 132.715 207.665 ;
        RECT 132.975 207.495 135.665 207.665 ;
        RECT 131.215 206.645 131.545 207.495 ;
        RECT 131.715 206.475 131.885 207.275 ;
        RECT 132.055 206.645 132.385 207.495 ;
        RECT 132.555 206.475 132.725 207.275 ;
        RECT 132.975 206.645 133.145 207.495 ;
        RECT 133.315 206.475 133.645 207.275 ;
        RECT 133.815 206.645 133.985 207.495 ;
        RECT 134.155 206.475 134.485 207.275 ;
        RECT 134.655 206.645 134.825 207.495 ;
        RECT 134.995 206.475 135.325 207.275 ;
        RECT 135.495 206.645 135.665 207.495 ;
        RECT 135.835 206.475 136.165 207.625 ;
        RECT 136.725 207.550 136.905 208.350 ;
        RECT 137.180 208.305 137.845 208.475 ;
        RECT 137.180 208.050 137.350 208.305 ;
        RECT 138.565 208.275 139.775 209.025 ;
        RECT 137.075 207.720 137.350 208.050 ;
        RECT 137.575 207.755 137.915 208.125 ;
        RECT 137.180 207.575 137.350 207.720 ;
        RECT 136.725 206.645 136.995 207.550 ;
        RECT 137.180 207.405 137.855 207.575 ;
        RECT 137.165 206.475 137.495 207.235 ;
        RECT 137.675 206.645 137.855 207.405 ;
        RECT 138.565 207.565 139.085 208.105 ;
        RECT 139.255 207.735 139.775 208.275 ;
        RECT 138.565 206.475 139.775 207.565 ;
        RECT 27.160 206.305 139.860 206.475 ;
        RECT 27.245 205.215 28.455 206.305 ;
        RECT 27.245 204.505 27.765 205.045 ;
        RECT 27.935 204.675 28.455 205.215 ;
        RECT 28.630 205.155 28.890 206.305 ;
        RECT 29.065 205.230 29.320 206.135 ;
        RECT 29.490 205.545 29.820 206.305 ;
        RECT 30.035 205.375 30.205 206.135 ;
        RECT 27.245 203.755 28.455 204.505 ;
        RECT 28.630 203.755 28.890 204.595 ;
        RECT 29.065 204.500 29.235 205.230 ;
        RECT 29.490 205.205 30.205 205.375 ;
        RECT 30.465 205.215 33.975 206.305 ;
        RECT 34.145 205.215 35.355 206.305 ;
        RECT 29.490 204.995 29.660 205.205 ;
        RECT 29.405 204.665 29.660 204.995 ;
        RECT 29.065 203.925 29.320 204.500 ;
        RECT 29.490 204.475 29.660 204.665 ;
        RECT 29.940 204.655 30.295 205.025 ;
        RECT 30.465 204.525 32.115 205.045 ;
        RECT 32.285 204.695 33.975 205.215 ;
        RECT 29.490 204.305 30.205 204.475 ;
        RECT 29.490 203.755 29.820 204.135 ;
        RECT 30.035 203.925 30.205 204.305 ;
        RECT 30.465 203.755 33.975 204.525 ;
        RECT 34.145 204.505 34.665 205.045 ;
        RECT 34.835 204.675 35.355 205.215 ;
        RECT 35.525 205.230 35.795 206.135 ;
        RECT 35.965 205.545 36.295 206.305 ;
        RECT 36.475 205.375 36.645 206.135 ;
        RECT 34.145 203.755 35.355 204.505 ;
        RECT 35.525 204.430 35.695 205.230 ;
        RECT 35.980 205.205 36.645 205.375 ;
        RECT 35.980 205.060 36.150 205.205 ;
        RECT 35.865 204.730 36.150 205.060 ;
        RECT 35.980 204.475 36.150 204.730 ;
        RECT 36.385 204.655 36.715 205.025 ;
        RECT 35.525 203.925 35.785 204.430 ;
        RECT 35.980 204.305 36.645 204.475 ;
        RECT 35.965 203.755 36.295 204.135 ;
        RECT 36.475 203.925 36.645 204.305 ;
        RECT 36.905 204.035 37.185 206.135 ;
        RECT 37.375 205.545 38.160 206.305 ;
        RECT 38.555 205.475 38.940 206.135 ;
        RECT 38.555 205.375 38.965 205.475 ;
        RECT 37.355 205.165 38.965 205.375 ;
        RECT 39.265 205.285 39.465 206.075 ;
        RECT 37.355 204.565 37.630 205.165 ;
        RECT 39.135 205.115 39.465 205.285 ;
        RECT 39.635 205.125 39.955 206.305 ;
        RECT 40.125 205.140 40.415 206.305 ;
        RECT 40.590 205.165 40.925 206.135 ;
        RECT 41.095 205.165 41.265 206.305 ;
        RECT 41.435 205.965 43.465 206.135 ;
        RECT 39.135 204.995 39.315 205.115 ;
        RECT 37.800 204.745 38.155 204.995 ;
        RECT 38.350 204.945 38.815 204.995 ;
        RECT 38.345 204.775 38.815 204.945 ;
        RECT 38.350 204.745 38.815 204.775 ;
        RECT 38.985 204.745 39.315 204.995 ;
        RECT 39.490 204.745 39.955 204.945 ;
        RECT 37.355 204.385 38.605 204.565 ;
        RECT 38.240 204.315 38.605 204.385 ;
        RECT 38.775 204.365 39.955 204.535 ;
        RECT 40.590 204.495 40.760 205.165 ;
        RECT 41.435 204.995 41.605 205.965 ;
        RECT 40.930 204.665 41.185 204.995 ;
        RECT 41.410 204.665 41.605 204.995 ;
        RECT 41.775 205.625 42.900 205.795 ;
        RECT 41.015 204.495 41.185 204.665 ;
        RECT 41.775 204.495 41.945 205.625 ;
        RECT 37.415 203.755 37.585 204.215 ;
        RECT 38.775 204.145 39.105 204.365 ;
        RECT 37.855 203.965 39.105 204.145 ;
        RECT 39.275 203.755 39.445 204.195 ;
        RECT 39.615 203.950 39.955 204.365 ;
        RECT 40.125 203.755 40.415 204.480 ;
        RECT 40.590 203.925 40.845 204.495 ;
        RECT 41.015 204.325 41.945 204.495 ;
        RECT 42.115 205.285 43.125 205.455 ;
        RECT 42.115 204.485 42.285 205.285 ;
        RECT 41.770 204.290 41.945 204.325 ;
        RECT 41.015 203.755 41.345 204.155 ;
        RECT 41.770 203.925 42.300 204.290 ;
        RECT 42.490 204.265 42.765 205.085 ;
        RECT 42.485 204.095 42.765 204.265 ;
        RECT 42.490 203.925 42.765 204.095 ;
        RECT 42.935 203.925 43.125 205.285 ;
        RECT 43.295 205.300 43.465 205.965 ;
        RECT 43.635 205.545 43.805 206.305 ;
        RECT 44.040 205.545 44.555 205.955 ;
        RECT 44.725 205.870 50.070 206.305 ;
        RECT 43.295 205.110 44.045 205.300 ;
        RECT 44.215 204.735 44.555 205.545 ;
        RECT 43.325 204.565 44.555 204.735 ;
        RECT 43.305 203.755 43.815 204.290 ;
        RECT 44.035 203.960 44.280 204.565 ;
        RECT 46.310 204.300 46.650 205.130 ;
        RECT 48.130 204.620 48.480 205.870 ;
        RECT 50.255 205.355 50.530 206.125 ;
        RECT 50.700 205.695 51.030 206.125 ;
        RECT 51.200 205.865 51.395 206.305 ;
        RECT 51.575 205.695 51.905 206.125 ;
        RECT 50.700 205.525 51.905 205.695 ;
        RECT 50.255 205.165 50.840 205.355 ;
        RECT 51.010 205.195 51.905 205.525 ;
        RECT 50.255 204.345 50.495 204.995 ;
        RECT 50.665 204.495 50.840 205.165 ;
        RECT 51.010 204.665 51.425 204.995 ;
        RECT 51.605 204.665 51.900 204.995 ;
        RECT 50.665 204.315 50.995 204.495 ;
        RECT 44.725 203.755 50.070 204.300 ;
        RECT 50.270 203.755 50.600 204.145 ;
        RECT 50.770 203.935 50.995 204.315 ;
        RECT 51.195 204.045 51.425 204.665 ;
        RECT 51.605 203.755 51.905 204.485 ;
        RECT 52.085 204.035 52.365 206.135 ;
        RECT 52.555 205.545 53.340 206.305 ;
        RECT 53.735 205.475 54.120 206.135 ;
        RECT 53.735 205.375 54.145 205.475 ;
        RECT 52.535 205.165 54.145 205.375 ;
        RECT 54.445 205.285 54.645 206.075 ;
        RECT 52.535 204.565 52.810 205.165 ;
        RECT 54.315 205.115 54.645 205.285 ;
        RECT 54.815 205.125 55.135 206.305 ;
        RECT 55.310 205.165 55.645 206.135 ;
        RECT 55.815 205.165 55.985 206.305 ;
        RECT 56.155 205.965 58.185 206.135 ;
        RECT 54.315 204.995 54.495 205.115 ;
        RECT 52.980 204.745 53.335 204.995 ;
        RECT 53.530 204.945 53.995 204.995 ;
        RECT 53.525 204.775 53.995 204.945 ;
        RECT 53.530 204.745 53.995 204.775 ;
        RECT 54.165 204.745 54.495 204.995 ;
        RECT 54.670 204.745 55.135 204.945 ;
        RECT 52.535 204.385 53.785 204.565 ;
        RECT 53.420 204.315 53.785 204.385 ;
        RECT 53.955 204.365 55.135 204.535 ;
        RECT 52.595 203.755 52.765 204.215 ;
        RECT 53.955 204.145 54.285 204.365 ;
        RECT 53.035 203.965 54.285 204.145 ;
        RECT 54.455 203.755 54.625 204.195 ;
        RECT 54.795 203.950 55.135 204.365 ;
        RECT 55.310 204.495 55.480 205.165 ;
        RECT 56.155 204.995 56.325 205.965 ;
        RECT 55.650 204.665 55.905 204.995 ;
        RECT 56.130 204.665 56.325 204.995 ;
        RECT 56.495 205.625 57.620 205.795 ;
        RECT 55.735 204.495 55.905 204.665 ;
        RECT 56.495 204.495 56.665 205.625 ;
        RECT 55.310 203.925 55.565 204.495 ;
        RECT 55.735 204.325 56.665 204.495 ;
        RECT 56.835 205.285 57.845 205.455 ;
        RECT 56.835 204.485 57.005 205.285 ;
        RECT 57.210 204.605 57.485 205.085 ;
        RECT 57.205 204.435 57.485 204.605 ;
        RECT 56.490 204.290 56.665 204.325 ;
        RECT 55.735 203.755 56.065 204.155 ;
        RECT 56.490 203.925 57.020 204.290 ;
        RECT 57.210 203.925 57.485 204.435 ;
        RECT 57.655 203.925 57.845 205.285 ;
        RECT 58.015 205.300 58.185 205.965 ;
        RECT 58.355 205.545 58.525 206.305 ;
        RECT 58.760 205.545 59.275 205.955 ;
        RECT 58.015 205.110 58.765 205.300 ;
        RECT 58.935 204.735 59.275 205.545 ;
        RECT 59.445 205.215 62.955 206.305 ;
        RECT 58.045 204.565 59.275 204.735 ;
        RECT 58.025 203.755 58.535 204.290 ;
        RECT 58.755 203.960 59.000 204.565 ;
        RECT 59.445 204.525 61.095 205.045 ;
        RECT 61.265 204.695 62.955 205.215 ;
        RECT 64.055 205.355 64.330 206.125 ;
        RECT 64.500 205.695 64.830 206.125 ;
        RECT 65.000 205.865 65.195 206.305 ;
        RECT 65.375 205.695 65.705 206.125 ;
        RECT 64.500 205.525 65.705 205.695 ;
        RECT 64.055 205.165 64.640 205.355 ;
        RECT 64.810 205.195 65.705 205.525 ;
        RECT 59.445 203.755 62.955 204.525 ;
        RECT 64.055 204.345 64.295 204.995 ;
        RECT 64.465 204.495 64.640 205.165 ;
        RECT 65.885 205.140 66.175 206.305 ;
        RECT 66.825 205.415 67.085 206.125 ;
        RECT 67.255 205.595 67.585 206.305 ;
        RECT 67.755 205.415 67.985 206.125 ;
        RECT 66.825 205.175 67.985 205.415 ;
        RECT 68.165 205.395 68.435 206.125 ;
        RECT 68.615 205.575 68.955 206.305 ;
        RECT 68.165 205.175 68.935 205.395 ;
        RECT 64.810 204.665 65.225 204.995 ;
        RECT 65.405 204.665 65.700 204.995 ;
        RECT 66.815 204.665 67.115 204.995 ;
        RECT 67.295 204.685 67.820 204.995 ;
        RECT 68.000 204.685 68.465 204.995 ;
        RECT 64.465 204.315 64.795 204.495 ;
        RECT 64.070 203.755 64.400 204.145 ;
        RECT 64.570 203.935 64.795 204.315 ;
        RECT 64.995 204.045 65.225 204.665 ;
        RECT 65.405 203.755 65.705 204.485 ;
        RECT 65.885 203.755 66.175 204.480 ;
        RECT 66.825 203.755 67.115 204.485 ;
        RECT 67.295 204.045 67.525 204.685 ;
        RECT 68.645 204.505 68.935 205.175 ;
        RECT 67.705 204.305 68.935 204.505 ;
        RECT 67.705 203.935 68.015 204.305 ;
        RECT 68.195 203.755 68.865 204.125 ;
        RECT 69.125 203.935 69.385 206.125 ;
        RECT 69.565 205.215 72.155 206.305 ;
        RECT 69.565 204.525 70.775 205.045 ;
        RECT 70.945 204.695 72.155 205.215 ;
        RECT 72.510 205.335 72.900 205.510 ;
        RECT 73.385 205.505 73.715 206.305 ;
        RECT 73.885 205.515 74.420 206.135 ;
        RECT 72.510 205.165 73.935 205.335 ;
        RECT 69.565 203.755 72.155 204.525 ;
        RECT 72.385 204.435 72.740 204.995 ;
        RECT 72.910 204.265 73.080 205.165 ;
        RECT 73.250 204.435 73.515 204.995 ;
        RECT 73.765 204.665 73.935 205.165 ;
        RECT 74.105 204.495 74.420 205.515 ;
        RECT 72.490 203.755 72.730 204.265 ;
        RECT 72.910 203.935 73.190 204.265 ;
        RECT 73.420 203.755 73.635 204.265 ;
        RECT 73.805 203.925 74.420 204.495 ;
        RECT 74.625 205.465 74.885 206.135 ;
        RECT 75.055 205.905 75.385 206.305 ;
        RECT 76.255 205.905 76.655 206.305 ;
        RECT 76.945 205.725 77.275 205.960 ;
        RECT 75.195 205.555 77.275 205.725 ;
        RECT 74.625 204.495 74.800 205.465 ;
        RECT 75.195 205.285 75.365 205.555 ;
        RECT 74.970 205.115 75.365 205.285 ;
        RECT 75.535 205.165 76.550 205.385 ;
        RECT 74.970 204.665 75.140 205.115 ;
        RECT 76.275 205.025 76.550 205.165 ;
        RECT 76.720 205.165 77.275 205.555 ;
        RECT 75.310 204.745 75.760 204.945 ;
        RECT 75.930 204.575 76.105 204.770 ;
        RECT 74.625 203.925 74.965 204.495 ;
        RECT 75.160 203.755 75.330 204.420 ;
        RECT 75.610 204.405 76.105 204.575 ;
        RECT 75.610 204.265 75.830 204.405 ;
        RECT 75.605 204.095 75.830 204.265 ;
        RECT 76.275 204.235 76.445 205.025 ;
        RECT 76.720 204.915 76.890 205.165 ;
        RECT 77.445 204.995 77.620 206.095 ;
        RECT 77.790 205.485 78.135 206.305 ;
        RECT 76.695 204.745 76.890 204.915 ;
        RECT 77.060 204.745 77.620 204.995 ;
        RECT 77.790 204.745 78.135 205.315 ;
        RECT 78.305 205.215 79.975 206.305 ;
        RECT 76.695 204.360 76.865 204.745 ;
        RECT 75.610 204.050 75.830 204.095 ;
        RECT 76.000 204.065 76.445 204.235 ;
        RECT 76.615 203.990 76.865 204.360 ;
        RECT 77.035 204.395 78.135 204.575 ;
        RECT 77.035 203.990 77.285 204.395 ;
        RECT 77.455 203.755 77.625 204.225 ;
        RECT 77.795 203.990 78.135 204.395 ;
        RECT 78.305 204.525 79.055 205.045 ;
        RECT 79.225 204.695 79.975 205.215 ;
        RECT 80.150 205.165 80.485 206.135 ;
        RECT 80.655 205.165 80.825 206.305 ;
        RECT 80.995 205.965 83.025 206.135 ;
        RECT 78.305 203.755 79.975 204.525 ;
        RECT 80.150 204.495 80.320 205.165 ;
        RECT 80.995 204.995 81.165 205.965 ;
        RECT 80.490 204.665 80.745 204.995 ;
        RECT 80.970 204.665 81.165 204.995 ;
        RECT 81.335 205.625 82.460 205.795 ;
        RECT 80.575 204.495 80.745 204.665 ;
        RECT 81.335 204.495 81.505 205.625 ;
        RECT 80.150 203.925 80.405 204.495 ;
        RECT 80.575 204.325 81.505 204.495 ;
        RECT 81.675 205.285 82.685 205.455 ;
        RECT 81.675 204.485 81.845 205.285 ;
        RECT 81.330 204.290 81.505 204.325 ;
        RECT 80.575 203.755 80.905 204.155 ;
        RECT 81.330 203.925 81.860 204.290 ;
        RECT 82.050 204.265 82.325 205.085 ;
        RECT 82.045 204.095 82.325 204.265 ;
        RECT 82.050 203.925 82.325 204.095 ;
        RECT 82.495 203.925 82.685 205.285 ;
        RECT 82.855 205.300 83.025 205.965 ;
        RECT 83.195 205.545 83.365 206.305 ;
        RECT 83.600 205.545 84.115 205.955 ;
        RECT 82.855 205.110 83.605 205.300 ;
        RECT 83.775 204.735 84.115 205.545 ;
        RECT 84.745 205.165 85.005 206.305 ;
        RECT 85.175 205.155 85.505 206.135 ;
        RECT 85.675 205.165 85.955 206.305 ;
        RECT 84.765 204.745 85.100 204.995 ;
        RECT 82.885 204.565 84.115 204.735 ;
        RECT 82.865 203.755 83.375 204.290 ;
        RECT 83.595 203.960 83.840 204.565 ;
        RECT 85.270 204.555 85.440 205.155 ;
        RECT 85.610 204.725 85.945 204.995 ;
        RECT 84.745 203.925 85.440 204.555 ;
        RECT 85.645 203.755 85.955 204.555 ;
        RECT 86.125 203.925 86.875 206.135 ;
        RECT 87.045 205.230 87.315 206.135 ;
        RECT 87.485 205.545 87.815 206.305 ;
        RECT 87.995 205.375 88.175 206.135 ;
        RECT 87.045 204.430 87.225 205.230 ;
        RECT 87.500 205.205 88.175 205.375 ;
        RECT 87.500 205.060 87.670 205.205 ;
        RECT 87.395 204.730 87.670 205.060 ;
        RECT 87.500 204.475 87.670 204.730 ;
        RECT 87.895 204.655 88.235 205.025 ;
        RECT 87.045 203.925 87.305 204.430 ;
        RECT 87.500 204.305 88.165 204.475 ;
        RECT 87.485 203.755 87.815 204.135 ;
        RECT 87.995 203.925 88.165 204.305 ;
        RECT 89.345 203.925 90.095 206.135 ;
        RECT 90.345 205.375 90.525 206.135 ;
        RECT 90.705 205.545 91.035 206.305 ;
        RECT 90.345 205.205 91.020 205.375 ;
        RECT 91.205 205.230 91.475 206.135 ;
        RECT 90.850 205.060 91.020 205.205 ;
        RECT 90.285 204.655 90.625 205.025 ;
        RECT 90.850 204.730 91.125 205.060 ;
        RECT 90.850 204.475 91.020 204.730 ;
        RECT 90.355 204.305 91.020 204.475 ;
        RECT 91.295 204.430 91.475 205.230 ;
        RECT 91.645 205.140 91.935 206.305 ;
        RECT 92.105 205.230 92.375 206.135 ;
        RECT 92.545 205.545 92.875 206.305 ;
        RECT 93.055 205.375 93.225 206.135 ;
        RECT 93.955 205.585 94.285 206.305 ;
        RECT 90.355 203.925 90.525 204.305 ;
        RECT 90.705 203.755 91.035 204.135 ;
        RECT 91.215 203.925 91.475 204.430 ;
        RECT 91.645 203.755 91.935 204.480 ;
        RECT 92.105 204.430 92.275 205.230 ;
        RECT 92.560 205.205 93.225 205.375 ;
        RECT 92.560 205.060 92.730 205.205 ;
        RECT 92.445 204.730 92.730 205.060 ;
        RECT 92.560 204.475 92.730 204.730 ;
        RECT 92.965 204.655 93.295 205.025 ;
        RECT 93.945 204.945 94.175 205.285 ;
        RECT 94.465 204.945 94.680 206.060 ;
        RECT 94.875 205.360 95.205 206.135 ;
        RECT 95.375 205.530 96.085 206.305 ;
        RECT 94.875 205.145 96.025 205.360 ;
        RECT 93.945 204.745 94.275 204.945 ;
        RECT 94.465 204.765 94.915 204.945 ;
        RECT 94.585 204.745 94.915 204.765 ;
        RECT 95.085 204.745 95.555 204.975 ;
        RECT 95.740 204.575 96.025 205.145 ;
        RECT 96.255 204.700 96.535 206.135 ;
        RECT 92.105 203.925 92.365 204.430 ;
        RECT 92.560 204.305 93.225 204.475 ;
        RECT 92.545 203.755 92.875 204.135 ;
        RECT 93.055 203.925 93.225 204.305 ;
        RECT 93.945 204.385 95.125 204.575 ;
        RECT 93.945 203.925 94.285 204.385 ;
        RECT 94.795 204.305 95.125 204.385 ;
        RECT 95.315 204.385 96.025 204.575 ;
        RECT 95.315 204.245 95.615 204.385 ;
        RECT 95.300 204.235 95.615 204.245 ;
        RECT 95.290 204.225 95.615 204.235 ;
        RECT 95.280 204.220 95.615 204.225 ;
        RECT 94.455 203.755 94.625 204.215 ;
        RECT 95.275 204.210 95.615 204.220 ;
        RECT 95.270 204.205 95.615 204.210 ;
        RECT 95.265 204.195 95.615 204.205 ;
        RECT 95.260 204.190 95.615 204.195 ;
        RECT 95.255 203.925 95.615 204.190 ;
        RECT 95.855 203.755 96.025 204.215 ;
        RECT 96.195 203.925 96.535 204.700 ;
        RECT 96.705 205.585 97.165 206.135 ;
        RECT 97.355 205.585 97.685 206.305 ;
        RECT 96.705 204.215 96.955 205.585 ;
        RECT 97.885 205.415 98.185 205.965 ;
        RECT 98.355 205.635 98.635 206.305 ;
        RECT 97.245 205.245 98.185 205.415 ;
        RECT 97.245 204.995 97.415 205.245 ;
        RECT 98.555 204.995 98.820 205.355 ;
        RECT 99.005 205.245 99.320 206.305 ;
        RECT 99.950 205.800 100.565 206.305 ;
        RECT 97.125 204.665 97.415 204.995 ;
        RECT 97.585 204.745 97.925 204.995 ;
        RECT 98.145 204.745 98.820 204.995 ;
        RECT 97.245 204.575 97.415 204.665 ;
        RECT 97.245 204.385 98.635 204.575 ;
        RECT 99.065 204.415 99.330 204.995 ;
        RECT 99.500 204.915 99.775 205.575 ;
        RECT 99.970 205.265 100.205 205.630 ;
        RECT 100.375 205.625 100.565 205.800 ;
        RECT 100.735 205.795 101.210 206.135 ;
        RECT 100.375 205.435 100.705 205.625 ;
        RECT 100.930 205.265 101.120 205.560 ;
        RECT 101.380 205.460 101.595 206.305 ;
        RECT 101.795 205.465 102.080 206.135 ;
        RECT 99.970 205.095 101.740 205.265 ;
        RECT 99.500 204.685 100.335 204.915 ;
        RECT 96.705 203.925 97.265 204.215 ;
        RECT 97.435 203.755 97.685 204.215 ;
        RECT 98.305 204.025 98.635 204.385 ;
        RECT 99.005 203.755 99.275 204.245 ;
        RECT 99.500 203.975 99.775 204.685 ;
        RECT 100.505 204.240 100.760 205.095 ;
        RECT 99.975 203.975 100.760 204.240 ;
        RECT 100.930 204.435 101.340 204.915 ;
        RECT 101.510 204.665 101.740 205.095 ;
        RECT 101.910 205.115 102.080 205.465 ;
        RECT 102.250 205.295 102.515 206.305 ;
        RECT 102.765 205.375 102.945 206.135 ;
        RECT 103.125 205.545 103.455 206.305 ;
        RECT 102.765 205.205 103.440 205.375 ;
        RECT 103.625 205.230 103.895 206.135 ;
        RECT 101.910 204.595 102.515 205.115 ;
        RECT 103.270 205.060 103.440 205.205 ;
        RECT 102.705 204.655 103.045 205.025 ;
        RECT 103.270 204.730 103.545 205.060 ;
        RECT 100.930 203.975 101.140 204.435 ;
        RECT 101.910 204.385 102.080 204.595 ;
        RECT 103.270 204.475 103.440 204.730 ;
        RECT 101.330 203.755 101.660 204.250 ;
        RECT 101.835 203.925 102.080 204.385 ;
        RECT 102.250 203.755 102.515 204.415 ;
        RECT 102.775 204.305 103.440 204.475 ;
        RECT 103.715 204.430 103.895 205.230 ;
        RECT 104.075 205.165 104.405 206.305 ;
        RECT 104.935 205.335 105.265 206.120 ;
        RECT 104.585 205.165 105.265 205.335 ;
        RECT 105.485 205.165 105.715 206.305 ;
        RECT 104.065 204.745 104.415 204.995 ;
        RECT 104.585 204.565 104.755 205.165 ;
        RECT 105.885 205.155 106.215 206.135 ;
        RECT 106.385 205.165 106.595 206.305 ;
        RECT 107.390 205.505 107.645 206.305 ;
        RECT 107.815 205.335 108.145 206.135 ;
        RECT 108.315 205.505 108.485 206.305 ;
        RECT 108.655 205.335 108.985 206.135 ;
        RECT 107.285 205.165 108.985 205.335 ;
        RECT 109.155 205.165 109.415 206.305 ;
        RECT 109.585 205.800 110.215 206.305 ;
        RECT 109.600 205.265 109.855 205.630 ;
        RECT 110.025 205.625 110.215 205.800 ;
        RECT 110.395 205.795 110.870 206.135 ;
        RECT 110.025 205.435 110.355 205.625 ;
        RECT 110.580 205.265 110.830 205.560 ;
        RECT 111.055 205.460 111.270 206.305 ;
        RECT 111.470 205.465 111.745 206.135 ;
        RECT 111.485 205.455 111.745 205.465 ;
        RECT 104.925 204.745 105.275 204.995 ;
        RECT 105.465 204.745 105.795 204.995 ;
        RECT 102.775 203.925 102.945 204.305 ;
        RECT 103.125 203.755 103.455 204.135 ;
        RECT 103.635 203.925 103.895 204.430 ;
        RECT 104.075 203.755 104.345 204.565 ;
        RECT 104.515 203.925 104.845 204.565 ;
        RECT 105.015 203.755 105.255 204.565 ;
        RECT 105.485 203.755 105.715 204.575 ;
        RECT 105.965 204.555 106.215 205.155 ;
        RECT 107.285 204.575 107.565 205.165 ;
        RECT 109.600 205.095 111.390 205.265 ;
        RECT 111.575 205.115 111.745 205.455 ;
        RECT 111.915 205.295 112.175 206.305 ;
        RECT 112.355 205.330 112.685 205.995 ;
        RECT 113.145 205.690 113.475 206.135 ;
        RECT 113.710 205.860 113.985 206.305 ;
        RECT 114.155 205.690 114.485 206.135 ;
        RECT 113.145 205.510 114.485 205.690 ;
        RECT 114.685 205.500 114.940 206.305 ;
        RECT 112.355 205.160 114.940 205.330 ;
        RECT 107.735 204.745 108.485 204.995 ;
        RECT 108.655 204.745 109.415 204.995 ;
        RECT 105.885 203.925 106.215 204.555 ;
        RECT 106.385 203.755 106.595 204.575 ;
        RECT 107.285 204.325 108.145 204.575 ;
        RECT 108.315 204.385 109.415 204.555 ;
        RECT 109.585 204.435 109.970 204.915 ;
        RECT 107.395 204.135 107.725 204.155 ;
        RECT 108.315 204.135 108.565 204.385 ;
        RECT 107.395 203.925 108.565 204.135 ;
        RECT 108.735 203.755 108.905 204.215 ;
        RECT 109.075 203.925 109.415 204.385 ;
        RECT 110.140 204.240 110.395 205.095 ;
        RECT 109.605 203.975 110.395 204.240 ;
        RECT 110.565 204.420 110.975 204.915 ;
        RECT 111.160 204.665 111.390 205.095 ;
        RECT 111.560 204.595 112.175 205.115 ;
        RECT 112.345 204.715 112.680 204.945 ;
        RECT 112.865 204.775 113.320 204.945 ;
        RECT 112.870 204.715 113.320 204.775 ;
        RECT 113.490 204.715 113.960 204.945 ;
        RECT 114.130 204.715 114.460 204.945 ;
        RECT 110.565 203.975 110.795 204.420 ;
        RECT 111.560 204.385 111.730 204.595 ;
        RECT 114.630 204.545 114.940 205.160 ;
        RECT 110.975 203.755 111.305 204.250 ;
        RECT 111.480 203.925 111.730 204.385 ;
        RECT 111.900 203.755 112.175 204.415 ;
        RECT 112.355 204.365 114.940 204.545 ;
        RECT 112.355 203.945 112.685 204.365 ;
        RECT 112.855 203.755 113.130 204.195 ;
        RECT 113.335 203.945 113.665 204.365 ;
        RECT 115.155 204.305 115.385 206.005 ;
        RECT 115.555 205.160 115.850 206.305 ;
        RECT 116.025 205.165 116.285 206.305 ;
        RECT 116.455 205.155 116.785 206.135 ;
        RECT 116.955 205.165 117.235 206.305 ;
        RECT 116.045 204.745 116.380 204.995 ;
        RECT 114.145 203.755 114.995 204.115 ;
        RECT 115.165 203.925 115.385 204.305 ;
        RECT 115.555 203.755 115.850 204.575 ;
        RECT 116.550 204.555 116.720 205.155 ;
        RECT 117.405 205.140 117.695 206.305 ;
        RECT 118.360 205.505 118.610 206.305 ;
        RECT 118.780 205.675 119.110 206.135 ;
        RECT 119.280 205.845 119.495 206.305 ;
        RECT 118.780 205.505 119.950 205.675 ;
        RECT 117.870 205.335 118.150 205.495 ;
        RECT 117.870 205.165 119.205 205.335 ;
        RECT 119.035 204.995 119.205 205.165 ;
        RECT 116.890 204.725 117.225 204.995 ;
        RECT 117.870 204.745 118.220 204.985 ;
        RECT 118.390 204.745 118.865 204.985 ;
        RECT 119.035 204.745 119.410 204.995 ;
        RECT 119.035 204.575 119.205 204.745 ;
        RECT 116.025 203.925 116.720 204.555 ;
        RECT 116.925 203.755 117.235 204.555 ;
        RECT 117.405 203.755 117.695 204.480 ;
        RECT 117.870 204.405 119.205 204.575 ;
        RECT 117.870 204.195 118.140 204.405 ;
        RECT 119.580 204.215 119.950 205.505 ;
        RECT 120.715 205.295 120.885 206.135 ;
        RECT 121.055 205.965 122.225 206.135 ;
        RECT 121.055 205.465 121.385 205.965 ;
        RECT 121.895 205.925 122.225 205.965 ;
        RECT 122.415 205.885 122.770 206.305 ;
        RECT 121.555 205.705 121.785 205.795 ;
        RECT 122.940 205.705 123.190 206.135 ;
        RECT 121.555 205.465 123.190 205.705 ;
        RECT 123.360 205.545 123.690 206.305 ;
        RECT 123.860 205.465 124.115 206.135 ;
        RECT 120.715 205.125 123.775 205.295 ;
        RECT 120.625 204.745 120.980 204.955 ;
        RECT 121.150 204.745 121.595 204.945 ;
        RECT 121.765 204.745 122.240 204.945 ;
        RECT 118.360 203.755 118.690 204.215 ;
        RECT 119.200 203.925 119.950 204.215 ;
        RECT 120.715 204.405 121.780 204.575 ;
        RECT 120.715 203.925 120.885 204.405 ;
        RECT 121.055 203.755 121.385 204.235 ;
        RECT 121.610 204.175 121.780 204.405 ;
        RECT 121.960 204.345 122.240 204.745 ;
        RECT 122.510 204.745 122.840 204.945 ;
        RECT 123.010 204.745 123.375 204.945 ;
        RECT 122.510 204.345 122.795 204.745 ;
        RECT 123.605 204.575 123.775 205.125 ;
        RECT 122.975 204.405 123.775 204.575 ;
        RECT 122.975 204.175 123.145 204.405 ;
        RECT 123.945 204.335 124.115 205.465 ;
        RECT 124.285 205.115 124.455 206.305 ;
        RECT 125.235 205.495 125.530 206.305 ;
        RECT 125.710 204.995 125.955 206.135 ;
        RECT 126.130 205.495 126.390 206.305 ;
        RECT 126.990 206.300 133.265 206.305 ;
        RECT 126.570 204.995 126.820 206.130 ;
        RECT 126.990 205.505 127.250 206.300 ;
        RECT 127.420 205.405 127.680 206.130 ;
        RECT 127.850 205.575 128.110 206.300 ;
        RECT 128.280 205.405 128.540 206.130 ;
        RECT 128.710 205.575 128.970 206.300 ;
        RECT 129.140 205.405 129.400 206.130 ;
        RECT 129.570 205.575 129.830 206.300 ;
        RECT 130.000 205.405 130.260 206.130 ;
        RECT 130.430 205.575 130.675 206.300 ;
        RECT 130.845 205.405 131.105 206.130 ;
        RECT 131.290 205.575 131.535 206.300 ;
        RECT 131.705 205.405 131.965 206.130 ;
        RECT 132.150 205.575 132.395 206.300 ;
        RECT 132.565 205.405 132.825 206.130 ;
        RECT 133.010 205.575 133.265 206.300 ;
        RECT 127.420 205.390 132.825 205.405 ;
        RECT 133.435 205.390 133.725 206.130 ;
        RECT 133.895 205.560 134.165 206.305 ;
        RECT 127.420 205.165 134.165 205.390 ;
        RECT 123.930 204.255 124.115 204.335 ;
        RECT 121.610 203.925 123.145 204.175 ;
        RECT 123.315 203.755 123.645 204.235 ;
        RECT 123.860 203.925 124.115 204.255 ;
        RECT 124.285 203.755 124.455 204.650 ;
        RECT 125.225 204.435 125.540 204.995 ;
        RECT 125.710 204.745 132.830 204.995 ;
        RECT 125.225 203.755 125.530 204.265 ;
        RECT 125.710 203.935 125.960 204.745 ;
        RECT 126.130 203.755 126.390 204.280 ;
        RECT 126.570 203.935 126.820 204.745 ;
        RECT 133.000 204.575 134.165 205.165 ;
        RECT 127.420 204.405 134.165 204.575 ;
        RECT 134.425 205.230 134.695 206.135 ;
        RECT 134.865 205.545 135.195 206.305 ;
        RECT 135.375 205.375 135.545 206.135 ;
        RECT 134.425 204.430 134.595 205.230 ;
        RECT 134.880 205.205 135.545 205.375 ;
        RECT 135.805 205.230 136.075 206.135 ;
        RECT 136.245 205.545 136.575 206.305 ;
        RECT 136.755 205.375 136.925 206.135 ;
        RECT 134.880 205.060 135.050 205.205 ;
        RECT 134.765 204.730 135.050 205.060 ;
        RECT 134.880 204.475 135.050 204.730 ;
        RECT 135.285 204.655 135.615 205.025 ;
        RECT 126.990 203.755 127.250 204.315 ;
        RECT 127.420 203.950 127.680 204.405 ;
        RECT 127.850 203.755 128.110 204.235 ;
        RECT 128.280 203.950 128.540 204.405 ;
        RECT 128.710 203.755 128.970 204.235 ;
        RECT 129.140 203.950 129.400 204.405 ;
        RECT 129.570 203.755 129.815 204.235 ;
        RECT 129.985 203.950 130.260 204.405 ;
        RECT 130.430 203.755 130.675 204.235 ;
        RECT 130.845 203.950 131.105 204.405 ;
        RECT 131.285 203.755 131.535 204.235 ;
        RECT 131.705 203.950 131.965 204.405 ;
        RECT 132.145 203.755 132.395 204.235 ;
        RECT 132.565 203.950 132.825 204.405 ;
        RECT 133.005 203.755 133.265 204.235 ;
        RECT 133.435 203.950 133.695 204.405 ;
        RECT 133.865 203.755 134.165 204.235 ;
        RECT 134.425 203.925 134.685 204.430 ;
        RECT 134.880 204.305 135.545 204.475 ;
        RECT 134.865 203.755 135.195 204.135 ;
        RECT 135.375 203.925 135.545 204.305 ;
        RECT 135.805 204.430 135.975 205.230 ;
        RECT 136.260 205.205 136.925 205.375 ;
        RECT 137.185 205.335 137.445 206.305 ;
        RECT 136.260 205.060 136.430 205.205 ;
        RECT 136.145 204.730 136.430 205.060 ;
        RECT 136.260 204.475 136.430 204.730 ;
        RECT 136.665 204.655 136.995 205.025 ;
        RECT 135.805 203.925 136.065 204.430 ;
        RECT 136.260 204.305 136.925 204.475 ;
        RECT 136.245 203.755 136.575 204.135 ;
        RECT 136.755 203.925 136.925 204.305 ;
        RECT 137.185 204.045 137.425 204.995 ;
        RECT 137.615 204.960 137.945 206.135 ;
        RECT 138.115 205.335 138.395 206.305 ;
        RECT 138.565 205.215 139.775 206.305 ;
        RECT 137.615 204.430 138.395 204.960 ;
        RECT 138.565 204.675 139.085 205.215 ;
        RECT 139.255 204.505 139.775 205.045 ;
        RECT 137.615 203.925 137.940 204.430 ;
        RECT 138.110 203.755 138.395 204.260 ;
        RECT 138.565 203.755 139.775 204.505 ;
        RECT 27.160 203.585 139.860 203.755 ;
        RECT 27.245 202.835 28.455 203.585 ;
        RECT 27.245 202.295 27.765 202.835 ;
        RECT 28.625 202.815 31.215 203.585 ;
        RECT 31.385 202.910 31.645 203.415 ;
        RECT 31.825 203.205 32.155 203.585 ;
        RECT 32.335 203.035 32.505 203.415 ;
        RECT 32.765 203.040 38.110 203.585 ;
        RECT 27.935 202.125 28.455 202.665 ;
        RECT 28.625 202.295 29.835 202.815 ;
        RECT 30.005 202.125 31.215 202.645 ;
        RECT 27.245 201.035 28.455 202.125 ;
        RECT 28.625 201.035 31.215 202.125 ;
        RECT 31.385 202.110 31.555 202.910 ;
        RECT 31.840 202.865 32.505 203.035 ;
        RECT 31.840 202.610 32.010 202.865 ;
        RECT 31.725 202.280 32.010 202.610 ;
        RECT 32.245 202.315 32.575 202.685 ;
        RECT 31.840 202.135 32.010 202.280 ;
        RECT 34.350 202.210 34.690 203.040 ;
        RECT 38.285 202.815 39.955 203.585 ;
        RECT 40.130 202.845 40.385 203.415 ;
        RECT 40.555 203.185 40.885 203.585 ;
        RECT 41.310 203.050 41.840 203.415 ;
        RECT 41.310 203.015 41.485 203.050 ;
        RECT 40.555 202.845 41.485 203.015 ;
        RECT 42.030 202.905 42.305 203.415 ;
        RECT 31.385 201.205 31.655 202.110 ;
        RECT 31.840 201.965 32.505 202.135 ;
        RECT 31.825 201.035 32.155 201.795 ;
        RECT 32.335 201.205 32.505 201.965 ;
        RECT 36.170 201.470 36.520 202.720 ;
        RECT 38.285 202.295 39.035 202.815 ;
        RECT 39.205 202.125 39.955 202.645 ;
        RECT 32.765 201.035 38.110 201.470 ;
        RECT 38.285 201.035 39.955 202.125 ;
        RECT 40.130 202.175 40.300 202.845 ;
        RECT 40.555 202.675 40.725 202.845 ;
        RECT 40.470 202.345 40.725 202.675 ;
        RECT 40.950 202.345 41.145 202.675 ;
        RECT 40.130 201.205 40.465 202.175 ;
        RECT 40.635 201.035 40.805 202.175 ;
        RECT 40.975 201.375 41.145 202.345 ;
        RECT 41.315 201.715 41.485 202.845 ;
        RECT 41.655 202.055 41.825 202.855 ;
        RECT 42.025 202.735 42.305 202.905 ;
        RECT 42.030 202.255 42.305 202.735 ;
        RECT 42.475 202.055 42.665 203.415 ;
        RECT 42.845 203.050 43.355 203.585 ;
        RECT 43.575 202.775 43.820 203.380 ;
        RECT 44.300 202.845 44.915 203.415 ;
        RECT 45.085 203.075 45.300 203.585 ;
        RECT 45.530 203.075 45.810 203.405 ;
        RECT 45.990 203.075 46.230 203.585 ;
        RECT 47.650 203.075 47.890 203.585 ;
        RECT 48.070 203.075 48.350 203.405 ;
        RECT 48.580 203.075 48.795 203.585 ;
        RECT 42.865 202.605 44.095 202.775 ;
        RECT 41.655 201.885 42.665 202.055 ;
        RECT 42.835 202.040 43.585 202.230 ;
        RECT 41.315 201.545 42.440 201.715 ;
        RECT 42.835 201.375 43.005 202.040 ;
        RECT 43.755 201.795 44.095 202.605 ;
        RECT 40.975 201.205 43.005 201.375 ;
        RECT 43.175 201.035 43.345 201.795 ;
        RECT 43.580 201.385 44.095 201.795 ;
        RECT 44.300 201.825 44.615 202.845 ;
        RECT 44.785 202.175 44.955 202.675 ;
        RECT 45.205 202.345 45.470 202.905 ;
        RECT 45.640 202.175 45.810 203.075 ;
        RECT 45.980 202.345 46.335 202.905 ;
        RECT 47.545 202.345 47.900 202.905 ;
        RECT 48.070 202.175 48.240 203.075 ;
        RECT 48.410 202.345 48.675 202.905 ;
        RECT 48.965 202.845 49.580 203.415 ;
        RECT 48.925 202.175 49.095 202.675 ;
        RECT 44.785 202.005 46.210 202.175 ;
        RECT 44.300 201.205 44.835 201.825 ;
        RECT 45.005 201.035 45.335 201.835 ;
        RECT 45.820 201.830 46.210 202.005 ;
        RECT 47.670 202.005 49.095 202.175 ;
        RECT 47.670 201.830 48.060 202.005 ;
        RECT 48.545 201.035 48.875 201.835 ;
        RECT 49.265 201.825 49.580 202.845 ;
        RECT 49.785 202.975 50.125 203.390 ;
        RECT 50.295 203.145 50.465 203.585 ;
        RECT 50.635 203.195 51.885 203.375 ;
        RECT 50.635 202.975 50.965 203.195 ;
        RECT 52.155 203.125 52.325 203.585 ;
        RECT 49.785 202.805 50.965 202.975 ;
        RECT 51.135 202.955 51.500 203.025 ;
        RECT 51.135 202.775 52.385 202.955 ;
        RECT 49.785 202.395 50.250 202.595 ;
        RECT 50.425 202.345 50.755 202.595 ;
        RECT 50.925 202.565 51.390 202.595 ;
        RECT 50.925 202.395 51.395 202.565 ;
        RECT 50.925 202.345 51.390 202.395 ;
        RECT 51.585 202.345 51.940 202.595 ;
        RECT 50.425 202.225 50.605 202.345 ;
        RECT 49.045 201.205 49.580 201.825 ;
        RECT 49.785 201.035 50.105 202.215 ;
        RECT 50.275 202.055 50.605 202.225 ;
        RECT 52.110 202.175 52.385 202.775 ;
        RECT 50.275 201.265 50.475 202.055 ;
        RECT 50.775 201.965 52.385 202.175 ;
        RECT 50.775 201.865 51.185 201.965 ;
        RECT 50.800 201.205 51.185 201.865 ;
        RECT 51.580 201.035 52.365 201.795 ;
        RECT 52.555 201.205 52.835 203.305 ;
        RECT 53.005 202.860 53.295 203.585 ;
        RECT 53.465 202.815 55.135 203.585 ;
        RECT 55.770 202.845 56.025 203.415 ;
        RECT 56.195 203.185 56.525 203.585 ;
        RECT 56.950 203.050 57.480 203.415 ;
        RECT 57.670 203.245 57.945 203.415 ;
        RECT 57.665 203.075 57.945 203.245 ;
        RECT 56.950 203.015 57.125 203.050 ;
        RECT 56.195 202.845 57.125 203.015 ;
        RECT 53.465 202.295 54.215 202.815 ;
        RECT 53.005 201.035 53.295 202.200 ;
        RECT 54.385 202.125 55.135 202.645 ;
        RECT 53.465 201.035 55.135 202.125 ;
        RECT 55.770 202.175 55.940 202.845 ;
        RECT 56.195 202.675 56.365 202.845 ;
        RECT 56.110 202.345 56.365 202.675 ;
        RECT 56.590 202.345 56.785 202.675 ;
        RECT 55.770 201.205 56.105 202.175 ;
        RECT 56.275 201.035 56.445 202.175 ;
        RECT 56.615 201.375 56.785 202.345 ;
        RECT 56.955 201.715 57.125 202.845 ;
        RECT 57.295 202.055 57.465 202.855 ;
        RECT 57.670 202.255 57.945 203.075 ;
        RECT 58.115 202.055 58.305 203.415 ;
        RECT 58.485 203.050 58.995 203.585 ;
        RECT 59.215 202.775 59.460 203.380 ;
        RECT 59.925 202.855 60.215 203.585 ;
        RECT 58.505 202.605 59.735 202.775 ;
        RECT 57.295 201.885 58.305 202.055 ;
        RECT 58.475 202.040 59.225 202.230 ;
        RECT 56.955 201.545 58.080 201.715 ;
        RECT 58.475 201.375 58.645 202.040 ;
        RECT 59.395 201.795 59.735 202.605 ;
        RECT 59.915 202.345 60.215 202.675 ;
        RECT 60.395 202.655 60.625 203.295 ;
        RECT 60.805 203.035 61.115 203.405 ;
        RECT 61.295 203.215 61.965 203.585 ;
        RECT 60.805 202.835 62.035 203.035 ;
        RECT 60.395 202.345 60.920 202.655 ;
        RECT 61.100 202.345 61.565 202.655 ;
        RECT 61.745 202.165 62.035 202.835 ;
        RECT 56.615 201.205 58.645 201.375 ;
        RECT 58.815 201.035 58.985 201.795 ;
        RECT 59.220 201.385 59.735 201.795 ;
        RECT 59.925 201.925 61.085 202.165 ;
        RECT 59.925 201.215 60.185 201.925 ;
        RECT 60.355 201.035 60.685 201.745 ;
        RECT 60.855 201.215 61.085 201.925 ;
        RECT 61.265 201.945 62.035 202.165 ;
        RECT 61.265 201.215 61.535 201.945 ;
        RECT 61.715 201.035 62.055 201.765 ;
        RECT 62.225 201.215 62.485 203.405 ;
        RECT 63.585 202.785 64.280 203.415 ;
        RECT 64.485 202.785 64.795 203.585 ;
        RECT 65.435 202.860 65.765 203.370 ;
        RECT 65.935 203.185 66.265 203.585 ;
        RECT 67.315 203.015 67.645 203.355 ;
        RECT 67.815 203.185 68.145 203.585 ;
        RECT 63.605 202.345 63.940 202.595 ;
        RECT 64.110 202.185 64.280 202.785 ;
        RECT 64.450 202.345 64.785 202.615 ;
        RECT 63.585 201.035 63.845 202.175 ;
        RECT 64.015 201.205 64.345 202.185 ;
        RECT 64.515 201.035 64.795 202.175 ;
        RECT 65.435 202.095 65.625 202.860 ;
        RECT 65.935 202.845 68.300 203.015 ;
        RECT 65.935 202.675 66.105 202.845 ;
        RECT 65.795 202.345 66.105 202.675 ;
        RECT 66.275 202.345 66.580 202.675 ;
        RECT 65.435 201.245 65.765 202.095 ;
        RECT 65.935 201.035 66.185 202.175 ;
        RECT 66.365 202.015 66.580 202.345 ;
        RECT 66.755 202.015 67.040 202.675 ;
        RECT 67.235 202.015 67.500 202.675 ;
        RECT 67.715 202.015 67.960 202.675 ;
        RECT 68.130 201.845 68.300 202.845 ;
        RECT 68.695 202.785 68.905 203.585 ;
        RECT 66.375 201.675 67.665 201.845 ;
        RECT 66.375 201.255 66.625 201.675 ;
        RECT 66.855 201.035 67.185 201.505 ;
        RECT 67.415 201.255 67.665 201.675 ;
        RECT 67.845 201.675 68.300 201.845 ;
        RECT 67.845 201.245 68.175 201.675 ;
        RECT 68.695 201.035 68.905 202.175 ;
        RECT 69.075 201.205 69.415 203.415 ;
        RECT 69.595 203.125 69.845 203.585 ;
        RECT 70.035 202.955 70.365 203.415 ;
        RECT 69.590 202.785 70.365 202.955 ;
        RECT 70.565 202.905 70.950 203.415 ;
        RECT 69.590 201.885 69.865 202.785 ;
        RECT 70.545 202.735 70.950 202.905 ;
        RECT 71.425 203.045 71.755 203.415 ;
        RECT 71.945 203.215 72.275 203.585 ;
        RECT 72.445 203.045 72.775 203.415 ;
        RECT 73.335 203.105 73.505 203.585 ;
        RECT 71.425 202.845 72.775 203.045 ;
        RECT 73.675 202.935 74.005 203.405 ;
        RECT 70.065 202.055 70.395 202.595 ;
        RECT 70.565 202.055 70.950 202.735 ;
        RECT 73.245 202.765 74.005 202.935 ;
        RECT 74.175 202.765 74.345 203.585 ;
        RECT 74.515 202.935 74.845 203.400 ;
        RECT 75.015 203.115 75.185 203.585 ;
        RECT 75.445 203.205 76.630 203.375 ;
        RECT 76.800 203.035 77.130 203.415 ;
        RECT 75.830 202.935 76.215 203.025 ;
        RECT 74.515 202.765 76.215 202.935 ;
        RECT 76.585 202.865 77.130 203.035 ;
        RECT 71.240 202.055 71.660 202.595 ;
        RECT 71.860 202.345 72.220 202.675 ;
        RECT 72.390 202.355 73.075 202.665 ;
        RECT 69.590 201.645 71.755 201.885 ;
        RECT 69.595 201.035 70.215 201.475 ;
        RECT 70.420 201.205 70.700 201.645 ;
        RECT 70.885 201.035 71.215 201.415 ;
        RECT 71.425 201.205 71.755 201.645 ;
        RECT 71.930 201.545 72.220 202.345 ;
        RECT 71.925 201.375 72.220 201.545 ;
        RECT 71.930 201.300 72.220 201.375 ;
        RECT 72.445 201.035 72.700 202.175 ;
        RECT 72.870 201.315 73.075 202.355 ;
        RECT 73.245 201.795 73.555 202.765 ;
        RECT 73.725 202.385 74.055 202.595 ;
        RECT 74.225 202.385 74.665 202.595 ;
        RECT 74.835 202.385 75.320 202.595 ;
        RECT 73.885 202.215 74.055 202.385 ;
        RECT 73.885 202.045 74.845 202.215 ;
        RECT 73.245 201.625 74.005 201.795 ;
        RECT 73.245 201.035 73.585 201.455 ;
        RECT 73.755 201.205 74.005 201.625 ;
        RECT 74.175 201.035 74.505 201.875 ;
        RECT 74.675 201.795 74.845 202.045 ;
        RECT 75.015 201.965 75.320 202.385 ;
        RECT 75.510 202.395 75.900 202.595 ;
        RECT 76.070 202.395 76.415 202.595 ;
        RECT 75.510 201.965 75.800 202.395 ;
        RECT 76.585 202.225 76.755 202.865 ;
        RECT 77.385 202.785 77.695 203.585 ;
        RECT 77.900 202.785 78.595 203.415 ;
        RECT 78.765 202.860 79.055 203.585 ;
        RECT 79.225 202.815 80.895 203.585 ;
        RECT 76.955 202.345 77.215 202.695 ;
        RECT 77.395 202.345 77.730 202.615 ;
        RECT 75.970 202.175 76.755 202.225 ;
        RECT 77.900 202.185 78.070 202.785 ;
        RECT 78.240 202.345 78.575 202.595 ;
        RECT 79.225 202.295 79.975 202.815 ;
        RECT 81.800 202.775 82.045 203.380 ;
        RECT 82.265 203.050 82.775 203.585 ;
        RECT 75.970 202.000 77.050 202.175 ;
        RECT 75.970 201.795 76.140 202.000 ;
        RECT 74.675 201.625 76.140 201.795 ;
        RECT 74.995 201.205 75.750 201.625 ;
        RECT 76.310 201.035 76.550 201.820 ;
        RECT 76.720 201.205 77.050 202.000 ;
        RECT 77.385 201.035 77.665 202.175 ;
        RECT 77.835 201.205 78.165 202.185 ;
        RECT 78.335 201.035 78.595 202.175 ;
        RECT 78.765 201.035 79.055 202.200 ;
        RECT 80.145 202.125 80.895 202.645 ;
        RECT 79.225 201.035 80.895 202.125 ;
        RECT 81.525 202.605 82.755 202.775 ;
        RECT 81.525 201.795 81.865 202.605 ;
        RECT 82.035 202.040 82.785 202.230 ;
        RECT 81.525 201.385 82.040 201.795 ;
        RECT 82.275 201.035 82.445 201.795 ;
        RECT 82.615 201.375 82.785 202.040 ;
        RECT 82.955 202.055 83.145 203.415 ;
        RECT 83.315 202.565 83.590 203.415 ;
        RECT 83.780 203.050 84.310 203.415 ;
        RECT 84.735 203.185 85.065 203.585 ;
        RECT 84.135 203.015 84.310 203.050 ;
        RECT 83.315 202.395 83.595 202.565 ;
        RECT 83.315 202.255 83.590 202.395 ;
        RECT 83.795 202.055 83.965 202.855 ;
        RECT 82.955 201.885 83.965 202.055 ;
        RECT 84.135 202.845 85.065 203.015 ;
        RECT 85.235 202.845 85.490 203.415 ;
        RECT 84.135 201.715 84.305 202.845 ;
        RECT 84.895 202.675 85.065 202.845 ;
        RECT 83.180 201.545 84.305 201.715 ;
        RECT 84.475 202.345 84.670 202.675 ;
        RECT 84.895 202.345 85.150 202.675 ;
        RECT 84.475 201.375 84.645 202.345 ;
        RECT 85.320 202.175 85.490 202.845 ;
        RECT 82.615 201.205 84.645 201.375 ;
        RECT 84.815 201.035 84.985 202.175 ;
        RECT 85.155 201.205 85.490 202.175 ;
        RECT 85.670 202.845 85.925 203.415 ;
        RECT 86.095 203.185 86.425 203.585 ;
        RECT 86.850 203.050 87.380 203.415 ;
        RECT 86.850 203.015 87.025 203.050 ;
        RECT 86.095 202.845 87.025 203.015 ;
        RECT 85.670 202.175 85.840 202.845 ;
        RECT 86.095 202.675 86.265 202.845 ;
        RECT 86.010 202.345 86.265 202.675 ;
        RECT 86.490 202.345 86.685 202.675 ;
        RECT 85.670 201.205 86.005 202.175 ;
        RECT 86.175 201.035 86.345 202.175 ;
        RECT 86.515 201.375 86.685 202.345 ;
        RECT 86.855 201.715 87.025 202.845 ;
        RECT 87.195 202.055 87.365 202.855 ;
        RECT 87.570 202.565 87.845 203.415 ;
        RECT 87.565 202.395 87.845 202.565 ;
        RECT 87.570 202.255 87.845 202.395 ;
        RECT 88.015 202.055 88.205 203.415 ;
        RECT 88.385 203.050 88.895 203.585 ;
        RECT 89.115 202.775 89.360 203.380 ;
        RECT 88.405 202.605 89.635 202.775 ;
        RECT 87.195 201.885 88.205 202.055 ;
        RECT 88.375 202.040 89.125 202.230 ;
        RECT 86.855 201.545 87.980 201.715 ;
        RECT 88.375 201.375 88.545 202.040 ;
        RECT 89.295 201.795 89.635 202.605 ;
        RECT 86.515 201.205 88.545 201.375 ;
        RECT 88.715 201.035 88.885 201.795 ;
        RECT 89.120 201.385 89.635 201.795 ;
        RECT 89.805 201.205 90.555 203.415 ;
        RECT 90.815 203.035 90.985 203.415 ;
        RECT 91.165 203.205 91.495 203.585 ;
        RECT 90.815 202.865 91.480 203.035 ;
        RECT 91.675 202.910 91.935 203.415 ;
        RECT 90.745 202.315 91.075 202.685 ;
        RECT 91.310 202.610 91.480 202.865 ;
        RECT 91.310 202.280 91.595 202.610 ;
        RECT 91.310 202.135 91.480 202.280 ;
        RECT 90.815 201.965 91.480 202.135 ;
        RECT 91.765 202.110 91.935 202.910 ;
        RECT 90.815 201.205 90.985 201.965 ;
        RECT 91.165 201.035 91.495 201.795 ;
        RECT 91.665 201.205 91.935 202.110 ;
        RECT 92.110 203.110 92.445 203.370 ;
        RECT 92.615 203.185 92.945 203.585 ;
        RECT 93.115 203.185 94.730 203.355 ;
        RECT 92.110 201.755 92.365 203.110 ;
        RECT 93.115 203.015 93.285 203.185 ;
        RECT 92.725 202.845 93.285 203.015 ;
        RECT 92.725 202.675 92.895 202.845 ;
        RECT 92.590 202.345 92.895 202.675 ;
        RECT 93.090 202.565 93.340 202.675 ;
        RECT 93.550 202.565 93.820 203.005 ;
        RECT 94.010 202.905 94.300 203.005 ;
        RECT 94.005 202.735 94.300 202.905 ;
        RECT 93.085 202.395 93.340 202.565 ;
        RECT 93.545 202.395 93.820 202.565 ;
        RECT 93.090 202.345 93.340 202.395 ;
        RECT 93.550 202.345 93.820 202.395 ;
        RECT 94.010 202.345 94.300 202.735 ;
        RECT 94.470 202.345 94.890 203.010 ;
        RECT 95.275 202.865 95.605 203.585 ;
        RECT 95.790 203.110 96.125 203.370 ;
        RECT 96.295 203.185 96.625 203.585 ;
        RECT 96.795 203.185 98.410 203.355 ;
        RECT 95.200 202.345 95.550 202.675 ;
        RECT 92.725 202.175 92.895 202.345 ;
        RECT 95.345 202.225 95.550 202.345 ;
        RECT 92.725 202.005 95.095 202.175 ;
        RECT 95.345 202.055 95.555 202.225 ;
        RECT 92.110 201.245 92.445 201.755 ;
        RECT 92.695 201.035 93.025 201.835 ;
        RECT 93.270 201.625 94.695 201.795 ;
        RECT 93.270 201.205 93.555 201.625 ;
        RECT 93.810 201.035 94.140 201.455 ;
        RECT 94.365 201.375 94.695 201.625 ;
        RECT 94.925 201.545 95.095 202.005 ;
        RECT 95.355 201.375 95.525 201.875 ;
        RECT 94.365 201.205 95.525 201.375 ;
        RECT 95.790 201.755 96.045 203.110 ;
        RECT 96.795 203.015 96.965 203.185 ;
        RECT 96.405 202.845 96.965 203.015 ;
        RECT 96.405 202.675 96.575 202.845 ;
        RECT 96.270 202.345 96.575 202.675 ;
        RECT 96.770 202.565 97.020 202.675 ;
        RECT 97.230 202.565 97.500 203.005 ;
        RECT 97.690 202.905 97.980 203.005 ;
        RECT 97.685 202.735 97.980 202.905 ;
        RECT 96.765 202.395 97.020 202.565 ;
        RECT 97.225 202.395 97.500 202.565 ;
        RECT 96.770 202.345 97.020 202.395 ;
        RECT 97.230 202.345 97.500 202.395 ;
        RECT 97.690 202.345 97.980 202.735 ;
        RECT 98.150 202.345 98.570 203.010 ;
        RECT 98.955 202.865 99.285 203.585 ;
        RECT 99.575 203.205 100.745 203.415 ;
        RECT 99.575 203.185 99.905 203.205 ;
        RECT 99.465 202.765 100.325 203.015 ;
        RECT 100.495 202.955 100.745 203.205 ;
        RECT 100.915 203.125 101.085 203.585 ;
        RECT 101.255 202.955 101.595 203.415 ;
        RECT 100.495 202.785 101.595 202.955 ;
        RECT 102.425 202.955 102.755 203.315 ;
        RECT 103.375 203.125 103.625 203.585 ;
        RECT 103.795 203.125 104.355 203.415 ;
        RECT 102.425 202.765 103.815 202.955 ;
        RECT 98.880 202.345 99.230 202.675 ;
        RECT 96.405 202.175 96.575 202.345 ;
        RECT 99.025 202.225 99.230 202.345 ;
        RECT 96.405 202.005 98.775 202.175 ;
        RECT 99.025 202.055 99.235 202.225 ;
        RECT 99.465 202.175 99.745 202.765 ;
        RECT 103.645 202.675 103.815 202.765 ;
        RECT 99.915 202.345 100.665 202.595 ;
        RECT 100.835 202.345 101.595 202.595 ;
        RECT 102.240 202.345 102.915 202.595 ;
        RECT 103.135 202.345 103.475 202.595 ;
        RECT 103.645 202.345 103.935 202.675 ;
        RECT 99.465 202.005 101.165 202.175 ;
        RECT 95.790 201.245 96.125 201.755 ;
        RECT 96.375 201.035 96.705 201.835 ;
        RECT 96.950 201.625 98.375 201.795 ;
        RECT 96.950 201.205 97.235 201.625 ;
        RECT 97.490 201.035 97.820 201.455 ;
        RECT 98.045 201.375 98.375 201.625 ;
        RECT 98.605 201.545 98.775 202.005 ;
        RECT 99.035 201.375 99.205 201.875 ;
        RECT 98.045 201.205 99.205 201.375 ;
        RECT 99.570 201.035 99.825 201.835 ;
        RECT 99.995 201.205 100.325 202.005 ;
        RECT 100.495 201.035 100.665 201.835 ;
        RECT 100.835 201.205 101.165 202.005 ;
        RECT 101.335 201.035 101.595 202.175 ;
        RECT 102.240 201.985 102.505 202.345 ;
        RECT 103.645 202.095 103.815 202.345 ;
        RECT 102.875 201.925 103.815 202.095 ;
        RECT 102.425 201.035 102.705 201.705 ;
        RECT 102.875 201.375 103.175 201.925 ;
        RECT 104.105 201.755 104.355 203.125 ;
        RECT 104.525 202.860 104.815 203.585 ;
        RECT 105.075 203.035 105.245 203.415 ;
        RECT 105.460 203.205 105.790 203.585 ;
        RECT 105.075 202.865 105.790 203.035 ;
        RECT 104.985 202.315 105.340 202.685 ;
        RECT 105.620 202.675 105.790 202.865 ;
        RECT 105.960 202.840 106.215 203.415 ;
        RECT 105.620 202.345 105.875 202.675 ;
        RECT 103.375 201.035 103.705 201.755 ;
        RECT 103.895 201.205 104.355 201.755 ;
        RECT 104.525 201.035 104.815 202.200 ;
        RECT 105.620 202.135 105.790 202.345 ;
        RECT 105.075 201.965 105.790 202.135 ;
        RECT 106.045 202.110 106.215 202.840 ;
        RECT 106.390 202.745 106.650 203.585 ;
        RECT 106.835 202.865 107.165 203.585 ;
        RECT 107.710 203.185 109.325 203.355 ;
        RECT 109.495 203.185 109.825 203.585 ;
        RECT 109.155 203.015 109.325 203.185 ;
        RECT 109.995 203.110 110.330 203.370 ;
        RECT 106.890 202.565 107.240 202.675 ;
        RECT 106.885 202.395 107.240 202.565 ;
        RECT 106.890 202.345 107.240 202.395 ;
        RECT 107.550 202.345 107.970 203.010 ;
        RECT 108.140 202.905 108.430 203.005 ;
        RECT 108.620 202.905 108.890 203.005 ;
        RECT 108.140 202.735 108.435 202.905 ;
        RECT 108.620 202.735 108.895 202.905 ;
        RECT 109.155 202.845 109.715 203.015 ;
        RECT 108.140 202.345 108.430 202.735 ;
        RECT 108.620 202.345 108.890 202.735 ;
        RECT 109.545 202.675 109.715 202.845 ;
        RECT 109.100 202.565 109.350 202.675 ;
        RECT 109.100 202.395 109.355 202.565 ;
        RECT 109.100 202.345 109.350 202.395 ;
        RECT 109.545 202.345 109.850 202.675 ;
        RECT 105.075 201.205 105.245 201.965 ;
        RECT 105.460 201.035 105.790 201.795 ;
        RECT 105.960 201.205 106.215 202.110 ;
        RECT 106.390 201.035 106.650 202.185 ;
        RECT 106.890 202.055 107.095 202.345 ;
        RECT 109.545 202.175 109.715 202.345 ;
        RECT 107.345 202.005 109.715 202.175 ;
        RECT 106.915 201.375 107.085 201.875 ;
        RECT 107.345 201.545 107.515 202.005 ;
        RECT 107.745 201.625 109.170 201.795 ;
        RECT 107.745 201.375 108.075 201.625 ;
        RECT 106.915 201.205 108.075 201.375 ;
        RECT 108.300 201.035 108.630 201.455 ;
        RECT 108.885 201.205 109.170 201.625 ;
        RECT 109.415 201.035 109.745 201.835 ;
        RECT 110.075 201.755 110.330 203.110 ;
        RECT 110.670 203.075 110.910 203.585 ;
        RECT 111.090 203.075 111.370 203.405 ;
        RECT 111.600 203.075 111.815 203.585 ;
        RECT 110.565 202.345 110.920 202.905 ;
        RECT 111.090 202.175 111.260 203.075 ;
        RECT 111.430 202.345 111.695 202.905 ;
        RECT 111.985 202.845 112.600 203.415 ;
        RECT 112.895 203.105 113.195 203.585 ;
        RECT 113.365 202.935 113.625 203.390 ;
        RECT 113.795 203.105 114.055 203.585 ;
        RECT 114.235 202.935 114.495 203.390 ;
        RECT 114.665 203.105 114.915 203.585 ;
        RECT 115.095 202.935 115.355 203.390 ;
        RECT 115.525 203.105 115.775 203.585 ;
        RECT 115.955 202.935 116.215 203.390 ;
        RECT 116.385 203.105 116.630 203.585 ;
        RECT 116.800 202.935 117.075 203.390 ;
        RECT 117.245 203.105 117.490 203.585 ;
        RECT 117.660 202.935 117.920 203.390 ;
        RECT 118.090 203.105 118.350 203.585 ;
        RECT 118.520 202.935 118.780 203.390 ;
        RECT 118.950 203.105 119.210 203.585 ;
        RECT 119.380 202.935 119.640 203.390 ;
        RECT 119.810 203.025 120.070 203.585 ;
        RECT 111.945 202.175 112.115 202.675 ;
        RECT 110.690 202.005 112.115 202.175 ;
        RECT 110.690 201.830 111.080 202.005 ;
        RECT 109.995 201.245 110.330 201.755 ;
        RECT 111.565 201.035 111.895 201.835 ;
        RECT 112.285 201.825 112.600 202.845 ;
        RECT 112.895 202.765 119.640 202.935 ;
        RECT 112.895 202.225 114.060 202.765 ;
        RECT 120.240 202.595 120.490 203.405 ;
        RECT 120.670 203.060 120.930 203.585 ;
        RECT 121.100 202.595 121.350 203.405 ;
        RECT 121.530 203.075 121.835 203.585 ;
        RECT 114.230 202.345 121.350 202.595 ;
        RECT 121.520 202.345 121.835 202.905 ;
        RECT 122.005 202.845 122.320 203.220 ;
        RECT 122.575 202.845 122.745 203.585 ;
        RECT 122.995 203.015 123.165 203.220 ;
        RECT 123.435 203.190 123.765 203.585 ;
        RECT 124.015 203.015 124.185 203.365 ;
        RECT 124.385 203.185 124.715 203.585 ;
        RECT 124.885 203.015 125.055 203.365 ;
        RECT 125.275 203.185 125.655 203.585 ;
        RECT 122.995 202.845 123.515 203.015 ;
        RECT 112.865 202.175 114.060 202.225 ;
        RECT 112.865 202.055 119.640 202.175 ;
        RECT 112.895 201.950 119.640 202.055 ;
        RECT 112.065 201.205 112.600 201.825 ;
        RECT 112.895 201.035 113.165 201.780 ;
        RECT 113.335 201.210 113.625 201.950 ;
        RECT 114.235 201.935 119.640 201.950 ;
        RECT 113.795 201.040 114.050 201.765 ;
        RECT 114.235 201.210 114.495 201.935 ;
        RECT 114.665 201.040 114.910 201.765 ;
        RECT 115.095 201.210 115.355 201.935 ;
        RECT 115.525 201.040 115.770 201.765 ;
        RECT 115.955 201.210 116.215 201.935 ;
        RECT 116.385 201.040 116.630 201.765 ;
        RECT 116.800 201.210 117.060 201.935 ;
        RECT 117.230 201.040 117.490 201.765 ;
        RECT 117.660 201.210 117.920 201.935 ;
        RECT 118.090 201.040 118.350 201.765 ;
        RECT 118.520 201.210 118.780 201.935 ;
        RECT 118.950 201.040 119.210 201.765 ;
        RECT 119.380 201.210 119.640 201.935 ;
        RECT 119.810 201.040 120.070 201.835 ;
        RECT 120.240 201.210 120.490 202.345 ;
        RECT 113.795 201.035 120.070 201.040 ;
        RECT 120.670 201.035 120.930 201.845 ;
        RECT 121.105 201.205 121.350 202.345 ;
        RECT 121.530 201.035 121.825 201.845 ;
        RECT 122.005 201.805 122.175 202.845 ;
        RECT 123.325 202.675 123.515 202.845 ;
        RECT 123.855 202.845 125.665 203.015 ;
        RECT 122.345 201.975 122.695 202.675 ;
        RECT 122.865 202.345 123.155 202.675 ;
        RECT 123.325 202.345 123.615 202.675 ;
        RECT 123.325 202.145 123.515 202.345 ;
        RECT 122.910 201.975 123.515 202.145 ;
        RECT 122.005 201.635 123.215 201.805 ;
        RECT 123.855 201.715 124.025 202.845 ;
        RECT 122.005 201.215 122.265 201.635 ;
        RECT 122.435 201.035 122.765 201.465 ;
        RECT 123.045 201.375 123.215 201.635 ;
        RECT 123.430 201.545 124.025 201.715 ;
        RECT 124.195 201.375 124.365 202.675 ;
        RECT 124.595 202.220 124.925 202.675 ;
        RECT 123.045 201.205 124.365 201.375 ;
        RECT 124.715 201.885 124.925 202.220 ;
        RECT 125.155 202.225 125.325 202.675 ;
        RECT 125.495 202.595 125.665 202.845 ;
        RECT 125.835 202.945 126.085 203.415 ;
        RECT 126.255 203.115 126.425 203.585 ;
        RECT 126.595 202.945 126.925 203.415 ;
        RECT 127.095 203.115 127.265 203.585 ;
        RECT 127.585 203.105 127.865 203.585 ;
        RECT 125.835 202.765 127.355 202.945 ;
        RECT 128.035 202.935 128.295 203.325 ;
        RECT 128.470 203.105 128.725 203.585 ;
        RECT 128.895 202.935 129.190 203.325 ;
        RECT 129.370 203.105 129.645 203.585 ;
        RECT 129.815 203.085 130.115 203.415 ;
        RECT 125.495 202.425 126.955 202.595 ;
        RECT 125.155 202.055 125.590 202.225 ;
        RECT 127.125 202.215 127.355 202.765 ;
        RECT 125.795 202.045 127.355 202.215 ;
        RECT 127.540 202.765 129.190 202.935 ;
        RECT 127.540 202.255 127.945 202.765 ;
        RECT 128.115 202.425 129.255 202.595 ;
        RECT 127.540 202.085 128.295 202.255 ;
        RECT 124.715 201.295 125.035 201.885 ;
        RECT 125.320 201.035 125.570 201.875 ;
        RECT 125.795 201.205 126.045 202.045 ;
        RECT 126.215 201.035 126.465 201.875 ;
        RECT 126.635 201.205 126.885 202.045 ;
        RECT 127.055 201.035 127.305 201.875 ;
        RECT 127.580 201.035 127.865 201.905 ;
        RECT 128.035 201.835 128.295 202.085 ;
        RECT 129.085 202.175 129.255 202.425 ;
        RECT 129.425 202.345 129.775 202.915 ;
        RECT 129.945 202.175 130.115 203.085 ;
        RECT 130.285 202.860 130.575 203.585 ;
        RECT 130.745 203.085 131.045 203.415 ;
        RECT 131.215 203.105 131.490 203.585 ;
        RECT 129.085 202.005 130.115 202.175 ;
        RECT 128.035 201.665 129.155 201.835 ;
        RECT 128.035 201.205 128.295 201.665 ;
        RECT 128.470 201.035 128.725 201.495 ;
        RECT 128.895 201.205 129.155 201.665 ;
        RECT 129.325 201.035 129.635 201.835 ;
        RECT 129.805 201.205 130.115 202.005 ;
        RECT 130.285 201.035 130.575 202.200 ;
        RECT 130.745 202.175 130.915 203.085 ;
        RECT 131.670 202.935 131.965 203.325 ;
        RECT 132.135 203.105 132.390 203.585 ;
        RECT 132.565 202.935 132.825 203.325 ;
        RECT 132.995 203.105 133.275 203.585 ;
        RECT 131.085 202.345 131.435 202.915 ;
        RECT 131.670 202.765 133.320 202.935 ;
        RECT 133.565 202.765 133.775 203.585 ;
        RECT 133.945 202.785 134.275 203.415 ;
        RECT 131.605 202.425 132.745 202.595 ;
        RECT 131.605 202.175 131.775 202.425 ;
        RECT 132.915 202.255 133.320 202.765 ;
        RECT 130.745 202.005 131.775 202.175 ;
        RECT 132.565 202.085 133.320 202.255 ;
        RECT 133.945 202.185 134.195 202.785 ;
        RECT 134.445 202.765 134.675 203.585 ;
        RECT 135.345 202.910 135.605 203.415 ;
        RECT 135.785 203.205 136.115 203.585 ;
        RECT 136.295 203.035 136.465 203.415 ;
        RECT 134.365 202.345 134.695 202.595 ;
        RECT 130.745 201.205 131.055 202.005 ;
        RECT 132.565 201.835 132.825 202.085 ;
        RECT 131.225 201.035 131.535 201.835 ;
        RECT 131.705 201.665 132.825 201.835 ;
        RECT 131.705 201.205 131.965 201.665 ;
        RECT 132.135 201.035 132.390 201.495 ;
        RECT 132.565 201.205 132.825 201.665 ;
        RECT 132.995 201.035 133.280 201.905 ;
        RECT 133.565 201.035 133.775 202.175 ;
        RECT 133.945 201.205 134.275 202.185 ;
        RECT 134.445 201.035 134.675 202.175 ;
        RECT 135.345 202.110 135.515 202.910 ;
        RECT 135.800 202.865 136.465 203.035 ;
        RECT 136.815 203.035 136.985 203.415 ;
        RECT 137.200 203.205 137.530 203.585 ;
        RECT 136.815 202.865 137.530 203.035 ;
        RECT 135.800 202.610 135.970 202.865 ;
        RECT 135.685 202.280 135.970 202.610 ;
        RECT 136.205 202.315 136.535 202.685 ;
        RECT 136.725 202.315 137.080 202.685 ;
        RECT 137.360 202.675 137.530 202.865 ;
        RECT 137.700 202.840 137.955 203.415 ;
        RECT 137.360 202.345 137.615 202.675 ;
        RECT 135.800 202.135 135.970 202.280 ;
        RECT 137.360 202.135 137.530 202.345 ;
        RECT 135.345 201.205 135.615 202.110 ;
        RECT 135.800 201.965 136.465 202.135 ;
        RECT 135.785 201.035 136.115 201.795 ;
        RECT 136.295 201.205 136.465 201.965 ;
        RECT 136.815 201.965 137.530 202.135 ;
        RECT 137.785 202.110 137.955 202.840 ;
        RECT 138.130 202.745 138.390 203.585 ;
        RECT 138.565 202.835 139.775 203.585 ;
        RECT 136.815 201.205 136.985 201.965 ;
        RECT 137.200 201.035 137.530 201.795 ;
        RECT 137.700 201.205 137.955 202.110 ;
        RECT 138.130 201.035 138.390 202.185 ;
        RECT 138.565 202.125 139.085 202.665 ;
        RECT 139.255 202.295 139.775 202.835 ;
        RECT 138.565 201.035 139.775 202.125 ;
        RECT 27.160 200.865 139.860 201.035 ;
        RECT 27.245 199.775 28.455 200.865 ;
        RECT 28.625 200.430 33.970 200.865 ;
        RECT 27.245 199.065 27.765 199.605 ;
        RECT 27.935 199.235 28.455 199.775 ;
        RECT 27.245 198.315 28.455 199.065 ;
        RECT 30.210 198.860 30.550 199.690 ;
        RECT 32.030 199.180 32.380 200.430 ;
        RECT 34.145 199.775 37.655 200.865 ;
        RECT 34.145 199.085 35.795 199.605 ;
        RECT 35.965 199.255 37.655 199.775 ;
        RECT 38.745 199.725 39.025 200.865 ;
        RECT 39.195 199.715 39.525 200.695 ;
        RECT 39.695 199.725 39.955 200.865 ;
        RECT 38.755 199.285 39.090 199.555 ;
        RECT 39.260 199.115 39.430 199.715 ;
        RECT 40.125 199.700 40.415 200.865 ;
        RECT 41.705 200.195 41.985 200.865 ;
        RECT 41.505 199.555 41.820 199.995 ;
        RECT 42.155 199.975 42.455 200.525 ;
        RECT 42.665 200.145 42.995 200.865 ;
        RECT 43.185 200.145 43.635 200.695 ;
        RECT 42.155 199.805 43.095 199.975 ;
        RECT 42.925 199.555 43.095 199.805 ;
        RECT 39.600 199.305 39.935 199.555 ;
        RECT 41.505 199.305 42.195 199.555 ;
        RECT 42.425 199.305 42.755 199.555 ;
        RECT 42.925 199.225 43.215 199.555 ;
        RECT 42.925 199.135 43.095 199.225 ;
        RECT 28.625 198.315 33.970 198.860 ;
        RECT 34.145 198.315 37.655 199.085 ;
        RECT 38.745 198.315 39.055 199.115 ;
        RECT 39.260 198.485 39.955 199.115 ;
        RECT 40.125 198.315 40.415 199.040 ;
        RECT 41.705 198.945 43.095 199.135 ;
        RECT 41.705 198.585 42.035 198.945 ;
        RECT 43.385 198.775 43.635 200.145 ;
        RECT 43.805 199.725 44.095 200.865 ;
        RECT 44.325 199.725 44.535 200.865 ;
        RECT 44.705 199.715 45.035 200.695 ;
        RECT 45.205 199.725 45.435 200.865 ;
        RECT 46.565 199.725 46.845 200.865 ;
        RECT 47.015 199.715 47.345 200.695 ;
        RECT 47.515 199.725 47.775 200.865 ;
        RECT 47.955 200.255 48.285 200.685 ;
        RECT 48.465 200.425 48.660 200.865 ;
        RECT 48.830 200.255 49.160 200.685 ;
        RECT 47.955 200.085 49.160 200.255 ;
        RECT 47.955 199.755 48.850 200.085 ;
        RECT 49.330 199.915 49.605 200.685 ;
        RECT 49.020 199.725 49.605 199.915 ;
        RECT 49.785 199.775 52.375 200.865 ;
        RECT 42.665 198.315 42.915 198.775 ;
        RECT 43.085 198.485 43.635 198.775 ;
        RECT 43.805 198.315 44.095 199.115 ;
        RECT 44.325 198.315 44.535 199.135 ;
        RECT 44.705 199.115 44.955 199.715 ;
        RECT 45.125 199.305 45.455 199.555 ;
        RECT 46.575 199.285 46.910 199.555 ;
        RECT 44.705 198.485 45.035 199.115 ;
        RECT 45.205 198.315 45.435 199.135 ;
        RECT 47.080 199.115 47.250 199.715 ;
        RECT 47.420 199.305 47.755 199.555 ;
        RECT 47.960 199.225 48.255 199.555 ;
        RECT 48.435 199.225 48.850 199.555 ;
        RECT 46.565 198.315 46.875 199.115 ;
        RECT 47.080 198.485 47.775 199.115 ;
        RECT 47.955 198.315 48.255 199.045 ;
        RECT 48.435 198.605 48.665 199.225 ;
        RECT 49.020 199.055 49.195 199.725 ;
        RECT 48.865 198.875 49.195 199.055 ;
        RECT 49.365 198.905 49.605 199.555 ;
        RECT 49.785 199.085 50.995 199.605 ;
        RECT 51.165 199.255 52.375 199.775 ;
        RECT 52.580 200.075 53.115 200.695 ;
        RECT 48.865 198.495 49.090 198.875 ;
        RECT 49.260 198.315 49.590 198.705 ;
        RECT 49.785 198.315 52.375 199.085 ;
        RECT 52.580 199.055 52.895 200.075 ;
        RECT 53.285 200.065 53.615 200.865 ;
        RECT 54.100 199.895 54.490 200.070 ;
        RECT 53.065 199.725 54.490 199.895 ;
        RECT 54.850 199.725 55.185 200.695 ;
        RECT 55.355 199.725 55.525 200.865 ;
        RECT 55.695 200.525 57.725 200.695 ;
        RECT 53.065 199.225 53.235 199.725 ;
        RECT 52.580 198.485 53.195 199.055 ;
        RECT 53.485 198.995 53.750 199.555 ;
        RECT 53.920 198.825 54.090 199.725 ;
        RECT 54.260 198.995 54.615 199.555 ;
        RECT 54.850 199.055 55.020 199.725 ;
        RECT 55.695 199.555 55.865 200.525 ;
        RECT 55.190 199.225 55.445 199.555 ;
        RECT 55.670 199.225 55.865 199.555 ;
        RECT 56.035 200.185 57.160 200.355 ;
        RECT 55.275 199.055 55.445 199.225 ;
        RECT 56.035 199.055 56.205 200.185 ;
        RECT 53.365 198.315 53.580 198.825 ;
        RECT 53.810 198.495 54.090 198.825 ;
        RECT 54.270 198.315 54.510 198.825 ;
        RECT 54.850 198.485 55.105 199.055 ;
        RECT 55.275 198.885 56.205 199.055 ;
        RECT 56.375 199.845 57.385 200.015 ;
        RECT 56.375 199.045 56.545 199.845 ;
        RECT 56.750 199.505 57.025 199.645 ;
        RECT 56.745 199.335 57.025 199.505 ;
        RECT 56.030 198.850 56.205 198.885 ;
        RECT 55.275 198.315 55.605 198.715 ;
        RECT 56.030 198.485 56.560 198.850 ;
        RECT 56.750 198.485 57.025 199.335 ;
        RECT 57.195 198.485 57.385 199.845 ;
        RECT 57.555 199.860 57.725 200.525 ;
        RECT 57.895 200.105 58.065 200.865 ;
        RECT 58.300 200.105 58.815 200.515 ;
        RECT 57.555 199.670 58.305 199.860 ;
        RECT 58.475 199.295 58.815 200.105 ;
        RECT 58.985 199.775 62.495 200.865 ;
        RECT 57.585 199.125 58.815 199.295 ;
        RECT 57.565 198.315 58.075 198.850 ;
        RECT 58.295 198.520 58.540 199.125 ;
        RECT 58.985 199.085 60.635 199.605 ;
        RECT 60.805 199.255 62.495 199.775 ;
        RECT 62.665 199.725 62.925 200.865 ;
        RECT 63.095 199.715 63.425 200.695 ;
        RECT 63.595 199.725 63.875 200.865 ;
        RECT 64.045 199.775 65.715 200.865 ;
        RECT 62.685 199.305 63.020 199.555 ;
        RECT 63.190 199.115 63.360 199.715 ;
        RECT 63.530 199.285 63.865 199.555 ;
        RECT 58.985 198.315 62.495 199.085 ;
        RECT 62.665 198.485 63.360 199.115 ;
        RECT 63.565 198.315 63.875 199.115 ;
        RECT 64.045 199.085 64.795 199.605 ;
        RECT 64.965 199.255 65.715 199.775 ;
        RECT 65.885 199.700 66.175 200.865 ;
        RECT 66.345 199.775 68.015 200.865 ;
        RECT 68.660 199.880 68.985 200.865 ;
        RECT 69.555 200.235 69.815 200.695 ;
        RECT 69.985 200.415 70.835 200.865 ;
        RECT 69.170 200.185 69.375 200.215 ;
        RECT 69.165 200.015 69.375 200.185 ;
        RECT 69.555 200.015 70.675 200.235 ;
        RECT 66.345 199.085 67.095 199.605 ;
        RECT 67.265 199.255 68.015 199.775 ;
        RECT 68.655 199.225 68.915 199.680 ;
        RECT 69.170 199.630 69.375 200.015 ;
        RECT 69.170 199.255 69.755 199.630 ;
        RECT 69.925 199.240 70.335 199.845 ;
        RECT 70.505 199.560 70.675 200.015 ;
        RECT 64.045 198.315 65.715 199.085 ;
        RECT 65.885 198.315 66.175 199.040 ;
        RECT 66.345 198.315 68.015 199.085 ;
        RECT 70.505 199.070 70.835 199.560 ;
        RECT 68.660 198.865 69.815 199.055 ;
        RECT 68.660 198.725 68.935 198.865 ;
        RECT 69.605 198.695 69.815 198.865 ;
        RECT 69.985 198.865 70.835 199.070 ;
        RECT 69.105 198.315 69.435 198.695 ;
        RECT 69.985 198.485 70.315 198.865 ;
        RECT 70.505 198.315 70.835 198.695 ;
        RECT 71.005 198.485 71.250 200.695 ;
        RECT 71.435 199.865 71.690 200.865 ;
        RECT 71.865 200.430 77.210 200.865 ;
        RECT 71.435 198.315 71.675 199.115 ;
        RECT 73.450 198.860 73.790 199.690 ;
        RECT 75.270 199.180 75.620 200.430 ;
        RECT 77.385 199.775 78.595 200.865 ;
        RECT 77.385 199.065 77.905 199.605 ;
        RECT 78.075 199.235 78.595 199.775 ;
        RECT 78.765 199.725 79.045 200.865 ;
        RECT 79.215 199.715 79.545 200.695 ;
        RECT 79.715 199.725 79.975 200.865 ;
        RECT 80.150 199.725 80.485 200.695 ;
        RECT 80.655 199.725 80.825 200.865 ;
        RECT 80.995 200.525 83.025 200.695 ;
        RECT 78.775 199.285 79.110 199.555 ;
        RECT 79.280 199.115 79.450 199.715 ;
        RECT 79.620 199.305 79.955 199.555 ;
        RECT 71.865 198.315 77.210 198.860 ;
        RECT 77.385 198.315 78.595 199.065 ;
        RECT 78.765 198.315 79.075 199.115 ;
        RECT 79.280 198.485 79.975 199.115 ;
        RECT 80.150 199.055 80.320 199.725 ;
        RECT 80.995 199.555 81.165 200.525 ;
        RECT 80.490 199.225 80.745 199.555 ;
        RECT 80.970 199.225 81.165 199.555 ;
        RECT 81.335 200.185 82.460 200.355 ;
        RECT 80.575 199.055 80.745 199.225 ;
        RECT 81.335 199.055 81.505 200.185 ;
        RECT 80.150 198.485 80.405 199.055 ;
        RECT 80.575 198.885 81.505 199.055 ;
        RECT 81.675 199.845 82.685 200.015 ;
        RECT 81.675 199.045 81.845 199.845 ;
        RECT 82.050 199.505 82.325 199.645 ;
        RECT 82.045 199.335 82.325 199.505 ;
        RECT 81.330 198.850 81.505 198.885 ;
        RECT 80.575 198.315 80.905 198.715 ;
        RECT 81.330 198.485 81.860 198.850 ;
        RECT 82.050 198.485 82.325 199.335 ;
        RECT 82.495 198.485 82.685 199.845 ;
        RECT 82.855 199.860 83.025 200.525 ;
        RECT 83.195 200.105 83.365 200.865 ;
        RECT 83.600 200.105 84.115 200.515 ;
        RECT 82.855 199.670 83.605 199.860 ;
        RECT 83.775 199.295 84.115 200.105 ;
        RECT 82.885 199.125 84.115 199.295 ;
        RECT 84.285 200.065 84.725 200.695 ;
        RECT 82.865 198.315 83.375 198.850 ;
        RECT 83.595 198.520 83.840 199.125 ;
        RECT 84.285 199.055 84.595 200.065 ;
        RECT 84.900 200.015 85.215 200.865 ;
        RECT 85.385 200.525 86.815 200.695 ;
        RECT 85.385 199.845 85.555 200.525 ;
        RECT 84.765 199.675 85.555 199.845 ;
        RECT 84.765 199.225 84.935 199.675 ;
        RECT 85.725 199.555 85.925 200.355 ;
        RECT 85.105 199.225 85.495 199.505 ;
        RECT 85.680 199.225 85.925 199.555 ;
        RECT 86.125 199.225 86.375 200.355 ;
        RECT 86.565 199.895 86.815 200.525 ;
        RECT 86.995 200.065 87.325 200.865 ;
        RECT 86.565 199.725 87.335 199.895 ;
        RECT 87.505 199.725 87.765 200.865 ;
        RECT 86.590 199.225 86.995 199.555 ;
        RECT 87.165 199.055 87.335 199.725 ;
        RECT 87.935 199.715 88.265 200.695 ;
        RECT 88.435 199.725 88.715 200.865 ;
        RECT 88.885 199.775 91.475 200.865 ;
        RECT 87.525 199.305 87.860 199.555 ;
        RECT 88.030 199.165 88.200 199.715 ;
        RECT 88.370 199.285 88.705 199.555 ;
        RECT 88.025 199.115 88.200 199.165 ;
        RECT 84.285 198.495 84.725 199.055 ;
        RECT 84.895 198.315 85.345 199.055 ;
        RECT 85.515 198.885 86.675 199.055 ;
        RECT 85.515 198.485 85.685 198.885 ;
        RECT 85.855 198.315 86.275 198.715 ;
        RECT 86.445 198.485 86.675 198.885 ;
        RECT 86.845 198.485 87.335 199.055 ;
        RECT 87.505 198.485 88.200 199.115 ;
        RECT 88.405 198.315 88.715 199.115 ;
        RECT 88.885 199.085 90.095 199.605 ;
        RECT 90.265 199.255 91.475 199.775 ;
        RECT 91.645 199.700 91.935 200.865 ;
        RECT 88.885 198.315 91.475 199.085 ;
        RECT 91.645 198.315 91.935 199.040 ;
        RECT 92.115 198.495 92.375 200.685 ;
        RECT 92.545 200.135 92.885 200.865 ;
        RECT 93.065 199.955 93.335 200.685 ;
        RECT 92.565 199.735 93.335 199.955 ;
        RECT 93.515 199.975 93.745 200.685 ;
        RECT 93.915 200.155 94.245 200.865 ;
        RECT 94.415 199.975 94.675 200.685 ;
        RECT 93.515 199.735 94.675 199.975 ;
        RECT 95.335 199.915 95.610 200.685 ;
        RECT 95.780 200.255 96.110 200.685 ;
        RECT 96.280 200.425 96.475 200.865 ;
        RECT 96.655 200.255 96.985 200.685 ;
        RECT 95.780 200.085 96.985 200.255 ;
        RECT 92.565 199.065 92.855 199.735 ;
        RECT 95.335 199.725 95.920 199.915 ;
        RECT 96.090 199.755 96.985 200.085 ;
        RECT 97.165 200.015 97.425 200.695 ;
        RECT 97.595 200.085 97.845 200.865 ;
        RECT 98.095 200.315 98.345 200.695 ;
        RECT 98.515 200.485 98.870 200.865 ;
        RECT 99.875 200.475 100.210 200.695 ;
        RECT 99.475 200.315 99.705 200.355 ;
        RECT 98.095 200.115 99.705 200.315 ;
        RECT 98.095 200.105 98.930 200.115 ;
        RECT 99.520 200.025 99.705 200.115 ;
        RECT 93.035 199.245 93.500 199.555 ;
        RECT 93.680 199.245 94.205 199.555 ;
        RECT 92.565 198.865 93.795 199.065 ;
        RECT 92.635 198.315 93.305 198.685 ;
        RECT 93.485 198.495 93.795 198.865 ;
        RECT 93.975 198.605 94.205 199.245 ;
        RECT 94.385 199.225 94.685 199.555 ;
        RECT 94.385 198.315 94.675 199.045 ;
        RECT 95.335 198.905 95.575 199.555 ;
        RECT 95.745 199.055 95.920 199.725 ;
        RECT 96.090 199.225 96.505 199.555 ;
        RECT 96.685 199.225 96.980 199.555 ;
        RECT 95.745 198.875 96.075 199.055 ;
        RECT 95.350 198.315 95.680 198.705 ;
        RECT 95.850 198.495 96.075 198.875 ;
        RECT 96.275 198.605 96.505 199.225 ;
        RECT 96.685 198.315 96.985 199.045 ;
        RECT 97.165 198.825 97.335 200.015 ;
        RECT 99.035 199.915 99.365 199.945 ;
        RECT 97.565 199.855 99.365 199.915 ;
        RECT 99.955 199.855 100.210 200.475 ;
        RECT 97.505 199.745 100.210 199.855 ;
        RECT 97.505 199.710 97.705 199.745 ;
        RECT 97.505 199.135 97.675 199.710 ;
        RECT 99.035 199.685 100.210 199.745 ;
        RECT 100.390 199.725 100.645 200.865 ;
        RECT 100.815 199.895 101.145 200.695 ;
        RECT 101.315 200.065 101.485 200.865 ;
        RECT 101.655 199.895 101.985 200.695 ;
        RECT 102.155 200.065 102.325 200.865 ;
        RECT 102.495 199.895 102.825 200.695 ;
        RECT 102.995 200.065 103.165 200.865 ;
        RECT 103.335 199.895 103.665 200.695 ;
        RECT 103.835 200.065 104.085 200.865 ;
        RECT 100.815 199.725 103.665 199.895 ;
        RECT 104.525 200.015 104.785 200.695 ;
        RECT 104.955 200.085 105.205 200.865 ;
        RECT 105.455 200.315 105.705 200.695 ;
        RECT 105.875 200.485 106.230 200.865 ;
        RECT 107.235 200.475 107.570 200.695 ;
        RECT 106.835 200.315 107.065 200.355 ;
        RECT 105.455 200.115 107.065 200.315 ;
        RECT 105.455 200.105 106.290 200.115 ;
        RECT 106.880 200.025 107.065 200.115 ;
        RECT 97.905 199.270 98.315 199.575 ;
        RECT 98.485 199.305 98.815 199.515 ;
        RECT 97.505 199.015 97.775 199.135 ;
        RECT 97.505 198.970 98.350 199.015 ;
        RECT 97.595 198.845 98.350 198.970 ;
        RECT 98.605 198.905 98.815 199.305 ;
        RECT 99.060 199.305 99.535 199.515 ;
        RECT 99.725 199.305 100.215 199.505 ;
        RECT 100.410 199.305 102.030 199.555 ;
        RECT 102.210 199.305 102.745 199.725 ;
        RECT 102.915 199.305 104.355 199.555 ;
        RECT 99.060 198.905 99.280 199.305 ;
        RECT 97.165 198.815 97.395 198.825 ;
        RECT 97.165 198.485 97.425 198.815 ;
        RECT 98.180 198.695 98.350 198.845 ;
        RECT 97.595 198.315 97.925 198.675 ;
        RECT 98.180 198.485 99.480 198.695 ;
        RECT 99.755 198.315 100.210 199.080 ;
        RECT 100.390 198.945 102.325 199.135 ;
        RECT 100.390 198.485 100.725 198.945 ;
        RECT 100.895 198.315 101.065 198.775 ;
        RECT 101.235 198.485 101.565 198.945 ;
        RECT 101.735 198.315 101.905 198.775 ;
        RECT 102.075 198.695 102.325 198.945 ;
        RECT 102.495 199.035 102.745 199.305 ;
        RECT 102.495 198.865 103.665 199.035 ;
        RECT 103.835 198.695 104.085 199.115 ;
        RECT 102.075 198.485 104.085 198.695 ;
        RECT 104.525 198.825 104.695 200.015 ;
        RECT 106.395 199.915 106.725 199.945 ;
        RECT 104.925 199.855 106.725 199.915 ;
        RECT 107.315 199.855 107.570 200.475 ;
        RECT 104.865 199.745 107.570 199.855 ;
        RECT 104.865 199.710 105.065 199.745 ;
        RECT 104.865 199.135 105.035 199.710 ;
        RECT 106.395 199.685 107.570 199.745 ;
        RECT 107.750 199.715 108.010 200.865 ;
        RECT 108.185 199.790 108.440 200.695 ;
        RECT 108.610 200.105 108.940 200.865 ;
        RECT 109.155 199.935 109.325 200.695 ;
        RECT 109.605 200.065 109.935 200.865 ;
        RECT 105.265 199.270 105.675 199.575 ;
        RECT 105.845 199.305 106.175 199.515 ;
        RECT 104.865 199.015 105.135 199.135 ;
        RECT 104.865 198.970 105.710 199.015 ;
        RECT 104.955 198.845 105.710 198.970 ;
        RECT 105.965 198.905 106.175 199.305 ;
        RECT 106.420 199.305 106.895 199.515 ;
        RECT 107.085 199.305 107.575 199.505 ;
        RECT 106.420 198.905 106.640 199.305 ;
        RECT 104.525 198.815 104.755 198.825 ;
        RECT 104.525 198.485 104.785 198.815 ;
        RECT 105.540 198.695 105.710 198.845 ;
        RECT 104.955 198.315 105.285 198.675 ;
        RECT 105.540 198.485 106.840 198.695 ;
        RECT 107.115 198.315 107.570 199.080 ;
        RECT 107.750 198.315 108.010 199.155 ;
        RECT 108.185 199.060 108.355 199.790 ;
        RECT 108.610 199.765 109.325 199.935 ;
        RECT 108.610 199.555 108.780 199.765 ;
        RECT 110.110 199.725 110.445 200.695 ;
        RECT 110.615 200.065 110.945 200.865 ;
        RECT 111.345 199.895 111.595 200.695 ;
        RECT 111.780 200.145 112.110 200.865 ;
        RECT 112.330 199.895 112.580 200.695 ;
        RECT 112.755 200.485 113.085 200.865 ;
        RECT 110.625 199.725 112.680 199.895 ;
        RECT 108.525 199.225 108.780 199.555 ;
        RECT 108.185 198.485 108.440 199.060 ;
        RECT 108.610 199.035 108.780 199.225 ;
        RECT 109.060 199.215 109.415 199.585 ;
        RECT 110.110 199.505 110.285 199.725 ;
        RECT 110.625 199.545 110.850 199.725 ;
        RECT 110.105 199.335 110.285 199.505 ;
        RECT 108.610 198.865 109.325 199.035 ;
        RECT 108.610 198.315 108.940 198.695 ;
        RECT 109.155 198.485 109.325 198.865 ;
        RECT 109.595 198.315 109.925 199.040 ;
        RECT 110.110 199.035 110.285 199.335 ;
        RECT 110.455 199.305 110.850 199.545 ;
        RECT 110.110 198.570 110.445 199.035 ;
        RECT 110.115 198.525 110.445 198.570 ;
        RECT 110.615 198.315 110.850 199.120 ;
        RECT 111.020 198.645 111.280 199.555 ;
        RECT 111.590 199.535 111.760 199.555 ;
        RECT 111.460 198.645 111.760 199.535 ;
        RECT 111.935 198.650 112.290 199.555 ;
        RECT 112.510 198.815 112.680 199.725 ;
        RECT 112.850 198.985 113.055 200.305 ;
        RECT 113.265 199.725 113.525 200.865 ;
        RECT 112.510 198.485 113.005 198.815 ;
        RECT 113.265 198.315 113.525 199.115 ;
        RECT 113.695 198.485 114.025 200.695 ;
        RECT 114.195 200.355 114.705 200.865 ;
        RECT 115.875 200.185 116.205 200.695 ;
        RECT 114.195 200.015 116.705 200.185 ;
        RECT 114.195 199.225 114.505 200.015 ;
        RECT 114.675 199.225 114.895 199.845 ;
        RECT 115.165 199.225 115.340 199.845 ;
        RECT 115.595 199.225 115.815 199.845 ;
        RECT 116.090 199.505 116.335 199.845 ;
        RECT 116.085 199.335 116.335 199.505 ;
        RECT 116.090 199.225 116.335 199.335 ;
        RECT 116.505 199.055 116.705 200.015 ;
        RECT 116.875 199.725 117.235 200.865 ;
        RECT 117.405 199.700 117.695 200.865 ;
        RECT 117.865 199.775 121.375 200.865 ;
        RECT 116.905 199.475 117.235 199.555 ;
        RECT 116.875 199.305 117.235 199.475 ;
        RECT 114.275 198.315 114.605 199.055 ;
        RECT 114.875 198.885 116.205 199.055 ;
        RECT 114.875 198.485 115.205 198.885 ;
        RECT 115.375 198.315 115.705 198.715 ;
        RECT 115.875 198.655 116.205 198.885 ;
        RECT 116.375 198.825 116.705 199.055 ;
        RECT 116.875 198.655 117.235 199.135 ;
        RECT 117.865 199.085 119.515 199.605 ;
        RECT 119.685 199.255 121.375 199.775 ;
        RECT 122.065 199.725 122.275 200.865 ;
        RECT 122.445 199.715 122.775 200.695 ;
        RECT 122.945 199.725 123.175 200.865 ;
        RECT 123.425 199.725 123.655 200.865 ;
        RECT 123.825 199.715 124.155 200.695 ;
        RECT 124.325 199.725 124.535 200.865 ;
        RECT 124.765 199.790 125.035 200.695 ;
        RECT 125.205 200.105 125.535 200.865 ;
        RECT 125.715 199.935 125.895 200.695 ;
        RECT 126.615 200.055 126.910 200.865 ;
        RECT 115.875 198.485 117.235 198.655 ;
        RECT 117.405 198.315 117.695 199.040 ;
        RECT 117.865 198.315 121.375 199.085 ;
        RECT 122.065 198.315 122.275 199.135 ;
        RECT 122.445 199.115 122.695 199.715 ;
        RECT 122.865 199.305 123.195 199.555 ;
        RECT 123.405 199.305 123.735 199.555 ;
        RECT 122.445 198.485 122.775 199.115 ;
        RECT 122.945 198.315 123.175 199.135 ;
        RECT 123.425 198.315 123.655 199.135 ;
        RECT 123.905 199.115 124.155 199.715 ;
        RECT 123.825 198.485 124.155 199.115 ;
        RECT 124.325 198.315 124.535 199.135 ;
        RECT 124.765 198.990 124.945 199.790 ;
        RECT 125.220 199.765 125.895 199.935 ;
        RECT 125.220 199.620 125.390 199.765 ;
        RECT 125.115 199.290 125.390 199.620 ;
        RECT 125.220 199.035 125.390 199.290 ;
        RECT 125.615 199.215 125.955 199.585 ;
        RECT 127.090 199.555 127.335 200.695 ;
        RECT 127.510 200.055 127.770 200.865 ;
        RECT 128.370 200.860 134.645 200.865 ;
        RECT 127.950 199.555 128.200 200.690 ;
        RECT 128.370 200.065 128.630 200.860 ;
        RECT 128.800 199.965 129.060 200.690 ;
        RECT 129.230 200.135 129.490 200.860 ;
        RECT 129.660 199.965 129.920 200.690 ;
        RECT 130.090 200.135 130.350 200.860 ;
        RECT 130.520 199.965 130.780 200.690 ;
        RECT 130.950 200.135 131.210 200.860 ;
        RECT 131.380 199.965 131.640 200.690 ;
        RECT 131.810 200.135 132.055 200.860 ;
        RECT 132.225 199.965 132.485 200.690 ;
        RECT 132.670 200.135 132.915 200.860 ;
        RECT 133.085 199.965 133.345 200.690 ;
        RECT 133.530 200.135 133.775 200.860 ;
        RECT 133.945 199.965 134.205 200.690 ;
        RECT 134.390 200.135 134.645 200.860 ;
        RECT 128.800 199.950 134.205 199.965 ;
        RECT 134.815 199.950 135.105 200.690 ;
        RECT 135.275 200.120 135.545 200.865 ;
        RECT 128.800 199.725 135.545 199.950 ;
        RECT 124.765 198.485 125.025 198.990 ;
        RECT 125.220 198.865 125.885 199.035 ;
        RECT 126.605 198.995 126.920 199.555 ;
        RECT 127.090 199.305 134.210 199.555 ;
        RECT 125.205 198.315 125.535 198.695 ;
        RECT 125.715 198.485 125.885 198.865 ;
        RECT 126.605 198.315 126.910 198.825 ;
        RECT 127.090 198.495 127.340 199.305 ;
        RECT 127.510 198.315 127.770 198.840 ;
        RECT 127.950 198.495 128.200 199.305 ;
        RECT 134.380 199.135 135.545 199.725 ;
        RECT 128.800 198.965 135.545 199.135 ;
        RECT 128.370 198.315 128.630 198.875 ;
        RECT 128.800 198.510 129.060 198.965 ;
        RECT 129.230 198.315 129.490 198.795 ;
        RECT 129.660 198.510 129.920 198.965 ;
        RECT 130.090 198.315 130.350 198.795 ;
        RECT 130.520 198.510 130.780 198.965 ;
        RECT 130.950 198.315 131.195 198.795 ;
        RECT 131.365 198.510 131.640 198.965 ;
        RECT 131.810 198.315 132.055 198.795 ;
        RECT 132.225 198.510 132.485 198.965 ;
        RECT 132.665 198.315 132.915 198.795 ;
        RECT 133.085 198.510 133.345 198.965 ;
        RECT 133.525 198.315 133.775 198.795 ;
        RECT 133.945 198.510 134.205 198.965 ;
        RECT 134.385 198.315 134.645 198.795 ;
        RECT 134.815 198.510 135.075 198.965 ;
        RECT 135.245 198.315 135.545 198.795 ;
        RECT 135.805 198.485 136.555 200.695 ;
        RECT 136.730 200.065 136.985 200.865 ;
        RECT 137.185 200.015 137.515 200.695 ;
        RECT 136.730 199.525 136.975 199.885 ;
        RECT 137.165 199.735 137.515 200.015 ;
        RECT 137.165 199.355 137.335 199.735 ;
        RECT 137.695 199.555 137.890 200.605 ;
        RECT 138.070 199.725 138.390 200.865 ;
        RECT 138.565 199.775 139.775 200.865 ;
        RECT 136.815 199.185 137.335 199.355 ;
        RECT 137.505 199.225 137.890 199.555 ;
        RECT 138.070 199.505 138.330 199.555 ;
        RECT 138.070 199.335 138.335 199.505 ;
        RECT 138.070 199.225 138.330 199.335 ;
        RECT 138.565 199.235 139.085 199.775 ;
        RECT 136.815 199.165 136.985 199.185 ;
        RECT 136.785 198.995 136.985 199.165 ;
        RECT 139.255 199.065 139.775 199.605 ;
        RECT 136.815 198.620 136.985 198.995 ;
        RECT 137.175 198.845 138.390 199.015 ;
        RECT 137.175 198.540 137.405 198.845 ;
        RECT 137.575 198.315 137.905 198.675 ;
        RECT 138.100 198.495 138.390 198.845 ;
        RECT 138.565 198.315 139.775 199.065 ;
        RECT 27.160 198.145 139.860 198.315 ;
        RECT 27.245 197.395 28.455 198.145 ;
        RECT 28.625 197.600 33.970 198.145 ;
        RECT 27.245 196.855 27.765 197.395 ;
        RECT 27.935 196.685 28.455 197.225 ;
        RECT 30.210 196.770 30.550 197.600 ;
        RECT 35.340 197.335 35.585 197.940 ;
        RECT 35.805 197.610 36.315 198.145 ;
        RECT 27.245 195.595 28.455 196.685 ;
        RECT 32.030 196.030 32.380 197.280 ;
        RECT 35.065 197.165 36.295 197.335 ;
        RECT 35.065 196.355 35.405 197.165 ;
        RECT 35.575 196.600 36.325 196.790 ;
        RECT 28.625 195.595 33.970 196.030 ;
        RECT 35.065 195.945 35.580 196.355 ;
        RECT 35.815 195.595 35.985 196.355 ;
        RECT 36.155 195.935 36.325 196.600 ;
        RECT 36.495 196.615 36.685 197.975 ;
        RECT 36.855 197.125 37.130 197.975 ;
        RECT 37.320 197.610 37.850 197.975 ;
        RECT 38.275 197.745 38.605 198.145 ;
        RECT 37.675 197.575 37.850 197.610 ;
        RECT 36.855 196.955 37.135 197.125 ;
        RECT 36.855 196.815 37.130 196.955 ;
        RECT 37.335 196.615 37.505 197.415 ;
        RECT 36.495 196.445 37.505 196.615 ;
        RECT 37.675 197.405 38.605 197.575 ;
        RECT 38.775 197.405 39.030 197.975 ;
        RECT 37.675 196.275 37.845 197.405 ;
        RECT 38.435 197.235 38.605 197.405 ;
        RECT 36.720 196.105 37.845 196.275 ;
        RECT 38.015 196.905 38.210 197.235 ;
        RECT 38.435 196.905 38.690 197.235 ;
        RECT 38.015 195.935 38.185 196.905 ;
        RECT 38.860 196.735 39.030 197.405 ;
        RECT 39.480 197.335 39.725 197.940 ;
        RECT 39.945 197.610 40.455 198.145 ;
        RECT 36.155 195.765 38.185 195.935 ;
        RECT 38.355 195.595 38.525 196.735 ;
        RECT 38.695 195.765 39.030 196.735 ;
        RECT 39.205 197.165 40.435 197.335 ;
        RECT 39.205 196.355 39.545 197.165 ;
        RECT 39.715 196.600 40.465 196.790 ;
        RECT 39.205 195.945 39.720 196.355 ;
        RECT 39.955 195.595 40.125 196.355 ;
        RECT 40.295 195.935 40.465 196.600 ;
        RECT 40.635 196.615 40.825 197.975 ;
        RECT 40.995 197.465 41.270 197.975 ;
        RECT 41.460 197.610 41.990 197.975 ;
        RECT 42.415 197.745 42.745 198.145 ;
        RECT 41.815 197.575 41.990 197.610 ;
        RECT 40.995 197.295 41.275 197.465 ;
        RECT 40.995 196.815 41.270 197.295 ;
        RECT 41.475 196.615 41.645 197.415 ;
        RECT 40.635 196.445 41.645 196.615 ;
        RECT 41.815 197.405 42.745 197.575 ;
        RECT 42.915 197.405 43.170 197.975 ;
        RECT 43.345 197.600 48.690 198.145 ;
        RECT 41.815 196.275 41.985 197.405 ;
        RECT 42.575 197.235 42.745 197.405 ;
        RECT 40.860 196.105 41.985 196.275 ;
        RECT 42.155 196.905 42.350 197.235 ;
        RECT 42.575 196.905 42.830 197.235 ;
        RECT 42.155 195.935 42.325 196.905 ;
        RECT 43.000 196.735 43.170 197.405 ;
        RECT 44.930 196.770 45.270 197.600 ;
        RECT 48.925 197.325 49.135 198.145 ;
        RECT 49.305 197.345 49.635 197.975 ;
        RECT 40.295 195.765 42.325 195.935 ;
        RECT 42.495 195.595 42.665 196.735 ;
        RECT 42.835 195.765 43.170 196.735 ;
        RECT 46.750 196.030 47.100 197.280 ;
        RECT 49.305 196.745 49.555 197.345 ;
        RECT 49.805 197.325 50.035 198.145 ;
        RECT 51.175 197.415 51.475 198.145 ;
        RECT 51.655 197.235 51.885 197.855 ;
        RECT 52.085 197.585 52.310 197.965 ;
        RECT 52.480 197.755 52.810 198.145 ;
        RECT 52.085 197.405 52.415 197.585 ;
        RECT 49.725 196.905 50.055 197.155 ;
        RECT 51.180 196.905 51.475 197.235 ;
        RECT 51.655 196.905 52.070 197.235 ;
        RECT 43.345 195.595 48.690 196.030 ;
        RECT 48.925 195.595 49.135 196.735 ;
        RECT 49.305 195.765 49.635 196.745 ;
        RECT 52.240 196.735 52.415 197.405 ;
        RECT 52.585 196.905 52.825 197.555 ;
        RECT 53.005 197.420 53.295 198.145 ;
        RECT 53.465 197.600 58.810 198.145 ;
        RECT 58.985 197.600 64.330 198.145 ;
        RECT 64.975 197.615 65.305 197.975 ;
        RECT 65.475 197.785 65.805 198.145 ;
        RECT 66.005 197.615 66.335 197.975 ;
        RECT 55.050 196.770 55.390 197.600 ;
        RECT 49.805 195.595 50.035 196.735 ;
        RECT 51.175 196.375 52.070 196.705 ;
        RECT 52.240 196.545 52.825 196.735 ;
        RECT 51.175 196.205 52.380 196.375 ;
        RECT 51.175 195.775 51.505 196.205 ;
        RECT 51.685 195.595 51.880 196.035 ;
        RECT 52.050 195.775 52.380 196.205 ;
        RECT 52.550 195.775 52.825 196.545 ;
        RECT 53.005 195.595 53.295 196.760 ;
        RECT 56.870 196.030 57.220 197.280 ;
        RECT 60.570 196.770 60.910 197.600 ;
        RECT 64.975 197.405 66.335 197.615 ;
        RECT 66.845 197.385 67.555 197.975 ;
        RECT 62.390 196.030 62.740 197.280 ;
        RECT 64.965 196.905 65.275 197.235 ;
        RECT 65.485 196.905 65.860 197.235 ;
        RECT 66.180 196.905 66.675 197.235 ;
        RECT 53.465 195.595 58.810 196.030 ;
        RECT 58.985 195.595 64.330 196.030 ;
        RECT 64.975 195.595 65.305 196.655 ;
        RECT 65.485 195.935 65.655 196.905 ;
        RECT 65.825 196.415 66.155 196.635 ;
        RECT 66.350 196.615 66.675 196.905 ;
        RECT 66.850 196.615 67.180 197.155 ;
        RECT 67.350 196.415 67.555 197.385 ;
        RECT 65.825 196.185 67.555 196.415 ;
        RECT 65.825 195.785 66.155 196.185 ;
        RECT 66.325 195.595 66.655 195.955 ;
        RECT 66.855 195.765 67.555 196.185 ;
        RECT 67.730 197.670 68.065 197.930 ;
        RECT 68.235 197.745 68.565 198.145 ;
        RECT 68.735 197.745 70.350 197.915 ;
        RECT 67.730 196.315 67.985 197.670 ;
        RECT 68.735 197.575 68.905 197.745 ;
        RECT 68.345 197.405 68.905 197.575 ;
        RECT 68.345 197.235 68.515 197.405 ;
        RECT 68.210 196.905 68.515 197.235 ;
        RECT 68.710 196.905 68.960 197.235 ;
        RECT 69.170 197.125 69.440 197.565 ;
        RECT 69.630 197.125 69.920 197.565 ;
        RECT 69.165 196.955 69.440 197.125 ;
        RECT 69.625 196.955 69.920 197.125 ;
        RECT 69.170 196.905 69.440 196.955 ;
        RECT 69.630 196.905 69.920 196.955 ;
        RECT 70.090 196.905 70.510 197.570 ;
        RECT 70.895 197.425 71.225 198.145 ;
        RECT 71.410 197.745 71.745 198.145 ;
        RECT 71.915 197.575 72.120 197.975 ;
        RECT 72.330 197.665 72.605 198.145 ;
        RECT 72.815 197.645 73.075 197.975 ;
        RECT 71.435 197.405 72.120 197.575 ;
        RECT 70.820 196.905 71.170 197.235 ;
        RECT 68.345 196.735 68.515 196.905 ;
        RECT 70.965 196.785 71.170 196.905 ;
        RECT 68.345 196.565 70.715 196.735 ;
        RECT 70.965 196.615 71.175 196.785 ;
        RECT 67.730 195.805 68.065 196.315 ;
        RECT 68.315 195.595 68.645 196.395 ;
        RECT 68.890 196.185 70.315 196.355 ;
        RECT 68.890 195.765 69.175 196.185 ;
        RECT 69.430 195.595 69.760 196.015 ;
        RECT 69.985 195.935 70.315 196.185 ;
        RECT 70.545 196.105 70.715 196.565 ;
        RECT 70.975 195.935 71.145 196.435 ;
        RECT 71.435 196.375 71.775 197.405 ;
        RECT 71.945 196.735 72.195 197.235 ;
        RECT 72.375 196.905 72.735 197.485 ;
        RECT 72.905 196.735 73.075 197.645 ;
        RECT 73.245 197.600 78.590 198.145 ;
        RECT 74.830 196.770 75.170 197.600 ;
        RECT 78.765 197.420 79.055 198.145 ;
        RECT 79.690 197.615 79.980 197.965 ;
        RECT 80.175 197.785 80.505 198.145 ;
        RECT 80.675 197.615 80.905 197.920 ;
        RECT 79.690 197.445 80.905 197.615 ;
        RECT 81.095 197.805 81.265 197.840 ;
        RECT 81.095 197.635 81.295 197.805 ;
        RECT 71.945 196.565 73.075 196.735 ;
        RECT 71.435 196.200 72.100 196.375 ;
        RECT 69.985 195.765 71.145 195.935 ;
        RECT 71.410 195.595 71.745 196.020 ;
        RECT 71.915 195.795 72.100 196.200 ;
        RECT 72.305 195.595 72.635 196.375 ;
        RECT 72.805 195.795 73.075 196.565 ;
        RECT 76.650 196.030 77.000 197.280 ;
        RECT 81.095 197.275 81.265 197.635 ;
        RECT 79.750 197.125 80.010 197.235 ;
        RECT 79.745 196.955 80.010 197.125 ;
        RECT 79.750 196.905 80.010 196.955 ;
        RECT 80.190 196.905 80.575 197.235 ;
        RECT 80.745 197.105 81.265 197.275 ;
        RECT 82.445 197.405 82.885 197.965 ;
        RECT 83.055 197.405 83.505 198.145 ;
        RECT 83.675 197.575 83.845 197.975 ;
        RECT 84.015 197.745 84.435 198.145 ;
        RECT 84.605 197.575 84.835 197.975 ;
        RECT 83.675 197.405 84.835 197.575 ;
        RECT 85.005 197.405 85.495 197.975 ;
        RECT 73.245 195.595 78.590 196.030 ;
        RECT 78.765 195.595 79.055 196.760 ;
        RECT 79.690 195.595 80.010 196.735 ;
        RECT 80.190 195.855 80.385 196.905 ;
        RECT 80.745 196.725 80.915 197.105 ;
        RECT 80.565 196.445 80.915 196.725 ;
        RECT 81.105 196.575 81.350 196.935 ;
        RECT 80.565 195.765 80.895 196.445 ;
        RECT 82.445 196.395 82.755 197.405 ;
        RECT 82.925 196.785 83.095 197.235 ;
        RECT 83.265 196.955 83.655 197.235 ;
        RECT 83.840 196.905 84.085 197.235 ;
        RECT 82.925 196.615 83.715 196.785 ;
        RECT 81.095 195.595 81.350 196.395 ;
        RECT 82.445 195.765 82.885 196.395 ;
        RECT 83.060 195.595 83.375 196.445 ;
        RECT 83.545 195.935 83.715 196.615 ;
        RECT 83.885 196.105 84.085 196.905 ;
        RECT 84.285 196.105 84.535 197.235 ;
        RECT 84.750 196.905 85.155 197.235 ;
        RECT 85.325 196.735 85.495 197.405 ;
        RECT 85.665 197.375 89.175 198.145 ;
        RECT 89.345 197.395 90.555 198.145 ;
        RECT 85.665 196.855 87.315 197.375 ;
        RECT 84.725 196.565 85.495 196.735 ;
        RECT 87.485 196.685 89.175 197.205 ;
        RECT 89.345 196.855 89.865 197.395 ;
        RECT 90.035 196.685 90.555 197.225 ;
        RECT 84.725 195.935 84.975 196.565 ;
        RECT 83.545 195.765 84.975 195.935 ;
        RECT 85.155 195.595 85.485 196.395 ;
        RECT 85.665 195.595 89.175 196.685 ;
        RECT 89.345 195.595 90.555 196.685 ;
        RECT 90.725 195.765 91.475 197.975 ;
        RECT 91.735 197.595 91.905 197.975 ;
        RECT 92.085 197.765 92.415 198.145 ;
        RECT 91.735 197.425 92.400 197.595 ;
        RECT 92.595 197.470 92.855 197.975 ;
        RECT 93.050 197.755 93.380 198.145 ;
        RECT 93.550 197.585 93.775 197.965 ;
        RECT 91.665 196.875 92.005 197.245 ;
        RECT 92.230 197.170 92.400 197.425 ;
        RECT 92.230 196.840 92.505 197.170 ;
        RECT 92.230 196.695 92.400 196.840 ;
        RECT 91.725 196.525 92.400 196.695 ;
        RECT 92.675 196.670 92.855 197.470 ;
        RECT 93.035 196.905 93.275 197.555 ;
        RECT 93.445 197.405 93.775 197.585 ;
        RECT 93.445 196.735 93.620 197.405 ;
        RECT 93.975 197.235 94.205 197.855 ;
        RECT 94.385 197.415 94.685 198.145 ;
        RECT 94.900 197.405 95.515 197.975 ;
        RECT 95.685 197.635 95.900 198.145 ;
        RECT 96.130 197.635 96.410 197.965 ;
        RECT 96.590 197.635 96.830 198.145 ;
        RECT 93.790 196.905 94.205 197.235 ;
        RECT 94.385 196.905 94.680 197.235 ;
        RECT 91.725 195.765 91.905 196.525 ;
        RECT 92.085 195.595 92.415 196.355 ;
        RECT 92.585 195.765 92.855 196.670 ;
        RECT 93.035 196.545 93.620 196.735 ;
        RECT 93.035 195.775 93.310 196.545 ;
        RECT 93.790 196.375 94.685 196.705 ;
        RECT 93.480 196.205 94.685 196.375 ;
        RECT 93.480 195.775 93.810 196.205 ;
        RECT 93.980 195.595 94.175 196.035 ;
        RECT 94.355 195.775 94.685 196.205 ;
        RECT 94.900 196.385 95.215 197.405 ;
        RECT 95.385 196.735 95.555 197.235 ;
        RECT 95.805 196.905 96.070 197.465 ;
        RECT 96.240 196.735 96.410 197.635 ;
        RECT 96.580 196.905 96.935 197.465 ;
        RECT 98.085 197.325 98.770 197.965 ;
        RECT 98.940 197.325 99.110 198.145 ;
        RECT 99.280 197.495 99.610 197.960 ;
        RECT 99.780 197.675 99.950 198.145 ;
        RECT 100.210 197.755 101.395 197.925 ;
        RECT 101.565 197.585 101.895 197.975 ;
        RECT 100.595 197.495 100.980 197.585 ;
        RECT 99.280 197.325 100.980 197.495 ;
        RECT 101.385 197.405 101.895 197.585 ;
        RECT 102.225 197.685 102.785 197.975 ;
        RECT 102.955 197.685 103.205 198.145 ;
        RECT 95.385 196.565 96.810 196.735 ;
        RECT 94.900 195.765 95.435 196.385 ;
        RECT 95.605 195.595 95.935 196.395 ;
        RECT 96.420 196.390 96.810 196.565 ;
        RECT 98.085 196.355 98.335 197.325 ;
        RECT 98.505 196.945 98.840 197.155 ;
        RECT 99.010 196.945 99.460 197.155 ;
        RECT 99.650 196.945 100.135 197.155 ;
        RECT 98.670 196.775 98.840 196.945 ;
        RECT 99.760 196.785 100.135 196.945 ;
        RECT 100.325 196.905 100.705 197.155 ;
        RECT 100.885 196.945 101.215 197.155 ;
        RECT 98.670 196.605 99.590 196.775 ;
        RECT 98.085 195.765 98.750 196.355 ;
        RECT 98.920 195.595 99.250 196.435 ;
        RECT 99.420 196.355 99.590 196.605 ;
        RECT 99.760 196.615 100.155 196.785 ;
        RECT 99.760 196.525 100.135 196.615 ;
        RECT 100.325 196.525 100.645 196.905 ;
        RECT 101.385 196.775 101.555 197.405 ;
        RECT 101.725 196.945 102.055 197.235 ;
        RECT 100.815 196.605 101.900 196.775 ;
        RECT 100.815 196.355 100.985 196.605 ;
        RECT 99.420 196.185 100.985 196.355 ;
        RECT 99.760 195.765 100.565 196.185 ;
        RECT 101.155 195.595 101.405 196.435 ;
        RECT 101.600 195.765 101.900 196.605 ;
        RECT 102.225 196.315 102.475 197.685 ;
        RECT 103.825 197.515 104.155 197.875 ;
        RECT 102.765 197.325 104.155 197.515 ;
        RECT 104.525 197.420 104.815 198.145 ;
        RECT 105.025 197.325 105.255 198.145 ;
        RECT 105.425 197.345 105.755 197.975 ;
        RECT 102.765 197.235 102.935 197.325 ;
        RECT 102.645 196.905 102.935 197.235 ;
        RECT 103.105 196.905 103.445 197.155 ;
        RECT 103.665 196.905 104.340 197.155 ;
        RECT 105.005 196.905 105.335 197.155 ;
        RECT 102.765 196.655 102.935 196.905 ;
        RECT 102.765 196.485 103.705 196.655 ;
        RECT 104.075 196.545 104.340 196.905 ;
        RECT 102.225 195.765 102.685 196.315 ;
        RECT 102.875 195.595 103.205 196.315 ;
        RECT 103.405 195.935 103.705 196.485 ;
        RECT 103.875 195.595 104.155 196.265 ;
        RECT 104.525 195.595 104.815 196.760 ;
        RECT 105.505 196.745 105.755 197.345 ;
        RECT 105.925 197.325 106.135 198.145 ;
        RECT 106.385 197.635 106.625 198.145 ;
        RECT 106.370 196.905 106.625 197.465 ;
        RECT 106.795 197.405 107.125 197.940 ;
        RECT 107.340 197.405 107.510 198.145 ;
        RECT 107.720 197.495 108.050 197.965 ;
        RECT 108.220 197.665 108.390 198.145 ;
        RECT 108.560 197.495 108.890 197.965 ;
        RECT 109.060 197.665 109.230 198.145 ;
        RECT 105.025 195.595 105.255 196.735 ;
        RECT 105.425 195.765 105.755 196.745 ;
        RECT 106.795 196.735 106.975 197.405 ;
        RECT 107.720 197.325 109.415 197.495 ;
        RECT 109.585 197.345 109.845 198.145 ;
        RECT 107.145 196.905 107.520 197.235 ;
        RECT 107.690 196.985 108.900 197.155 ;
        RECT 107.690 196.735 107.895 196.985 ;
        RECT 109.070 196.735 109.415 197.325 ;
        RECT 105.925 195.595 106.135 196.735 ;
        RECT 106.435 196.565 107.895 196.735 ;
        RECT 108.560 196.565 109.415 196.735 ;
        RECT 106.435 195.765 106.795 196.565 ;
        RECT 108.560 196.395 108.890 196.565 ;
        RECT 107.340 195.595 107.510 196.395 ;
        RECT 107.720 196.225 108.890 196.395 ;
        RECT 107.720 195.765 108.050 196.225 ;
        RECT 108.220 195.595 108.390 196.055 ;
        RECT 108.560 195.765 108.890 196.225 ;
        RECT 109.060 195.595 109.230 196.395 ;
        RECT 109.585 195.595 109.845 196.735 ;
        RECT 110.015 195.765 110.345 197.975 ;
        RECT 110.595 197.405 110.925 198.145 ;
        RECT 111.195 197.575 111.525 197.975 ;
        RECT 111.695 197.745 112.025 198.145 ;
        RECT 112.195 197.805 113.555 197.975 ;
        RECT 112.195 197.575 112.525 197.805 ;
        RECT 111.195 197.405 112.525 197.575 ;
        RECT 112.695 197.405 113.025 197.635 ;
        RECT 110.515 196.445 110.825 197.235 ;
        RECT 110.995 196.615 111.215 197.235 ;
        RECT 111.485 196.615 111.660 197.235 ;
        RECT 111.915 196.615 112.135 197.235 ;
        RECT 112.410 196.785 112.655 197.235 ;
        RECT 112.405 196.615 112.655 196.785 ;
        RECT 112.825 196.445 113.025 197.405 ;
        RECT 113.195 197.325 113.555 197.805 ;
        RECT 113.725 197.635 114.030 198.145 ;
        RECT 113.195 196.985 113.555 197.155 ;
        RECT 113.225 196.905 113.555 196.985 ;
        RECT 113.725 196.905 114.040 197.465 ;
        RECT 114.210 197.155 114.460 197.965 ;
        RECT 114.630 197.620 114.890 198.145 ;
        RECT 115.070 197.155 115.320 197.965 ;
        RECT 115.490 197.585 115.750 198.145 ;
        RECT 115.920 197.495 116.180 197.950 ;
        RECT 116.350 197.665 116.610 198.145 ;
        RECT 116.780 197.495 117.040 197.950 ;
        RECT 117.210 197.665 117.470 198.145 ;
        RECT 117.640 197.495 117.900 197.950 ;
        RECT 118.070 197.665 118.315 198.145 ;
        RECT 118.485 197.495 118.760 197.950 ;
        RECT 118.930 197.665 119.175 198.145 ;
        RECT 119.345 197.495 119.605 197.950 ;
        RECT 119.785 197.665 120.035 198.145 ;
        RECT 120.205 197.495 120.465 197.950 ;
        RECT 120.645 197.665 120.895 198.145 ;
        RECT 121.065 197.495 121.325 197.950 ;
        RECT 121.505 197.665 121.765 198.145 ;
        RECT 121.935 197.495 122.195 197.950 ;
        RECT 122.365 197.665 122.665 198.145 ;
        RECT 123.015 197.665 123.185 198.145 ;
        RECT 123.355 197.495 123.685 197.965 ;
        RECT 115.920 197.325 122.665 197.495 ;
        RECT 114.210 196.905 121.330 197.155 ;
        RECT 121.500 197.125 122.665 197.325 ;
        RECT 122.925 197.325 123.685 197.495 ;
        RECT 123.855 197.325 124.025 198.145 ;
        RECT 124.195 197.495 124.525 197.960 ;
        RECT 124.695 197.675 124.865 198.145 ;
        RECT 125.125 197.765 126.310 197.935 ;
        RECT 126.480 197.595 126.810 197.975 ;
        RECT 125.510 197.495 125.895 197.585 ;
        RECT 124.195 197.325 125.895 197.495 ;
        RECT 126.265 197.425 126.810 197.595 ;
        RECT 127.065 197.645 127.325 197.975 ;
        RECT 127.495 197.785 127.825 198.145 ;
        RECT 128.080 197.765 129.380 197.975 ;
        RECT 121.500 196.955 122.695 197.125 ;
        RECT 110.515 196.275 113.025 196.445 ;
        RECT 110.515 195.595 111.025 196.105 ;
        RECT 112.195 195.765 112.525 196.275 ;
        RECT 113.195 195.595 113.555 196.735 ;
        RECT 113.735 195.595 114.030 196.405 ;
        RECT 114.210 195.765 114.455 196.905 ;
        RECT 114.630 195.595 114.890 196.405 ;
        RECT 115.070 195.770 115.320 196.905 ;
        RECT 121.500 196.735 122.665 196.955 ;
        RECT 115.920 196.510 122.665 196.735 ;
        RECT 115.920 196.495 121.325 196.510 ;
        RECT 115.490 195.600 115.750 196.395 ;
        RECT 115.920 195.770 116.180 196.495 ;
        RECT 116.350 195.600 116.610 196.325 ;
        RECT 116.780 195.770 117.040 196.495 ;
        RECT 117.210 195.600 117.470 196.325 ;
        RECT 117.640 195.770 117.900 196.495 ;
        RECT 118.070 195.600 118.330 196.325 ;
        RECT 118.500 195.770 118.760 196.495 ;
        RECT 118.930 195.600 119.175 196.325 ;
        RECT 119.345 195.770 119.605 196.495 ;
        RECT 119.790 195.600 120.035 196.325 ;
        RECT 120.205 195.770 120.465 196.495 ;
        RECT 120.650 195.600 120.895 196.325 ;
        RECT 121.065 195.770 121.325 196.495 ;
        RECT 121.510 195.600 121.765 196.325 ;
        RECT 121.935 195.770 122.225 196.510 ;
        RECT 122.925 196.355 123.235 197.325 ;
        RECT 123.405 196.945 123.735 197.155 ;
        RECT 123.905 196.945 124.345 197.155 ;
        RECT 124.515 196.945 125.000 197.155 ;
        RECT 123.565 196.775 123.735 196.945 ;
        RECT 123.565 196.605 124.525 196.775 ;
        RECT 115.490 195.595 121.765 195.600 ;
        RECT 122.395 195.595 122.665 196.340 ;
        RECT 122.925 196.185 123.685 196.355 ;
        RECT 122.925 195.595 123.265 196.015 ;
        RECT 123.435 195.765 123.685 196.185 ;
        RECT 123.855 195.595 124.185 196.435 ;
        RECT 124.355 196.355 124.525 196.605 ;
        RECT 124.695 196.525 125.000 196.945 ;
        RECT 125.190 196.955 125.580 197.155 ;
        RECT 125.750 196.955 126.095 197.155 ;
        RECT 125.190 196.525 125.480 196.955 ;
        RECT 126.265 196.785 126.435 197.425 ;
        RECT 126.635 196.905 126.895 197.255 ;
        RECT 125.650 196.735 126.435 196.785 ;
        RECT 125.650 196.560 126.730 196.735 ;
        RECT 125.650 196.355 125.820 196.560 ;
        RECT 124.355 196.185 125.820 196.355 ;
        RECT 124.675 195.765 125.430 196.185 ;
        RECT 125.990 195.595 126.230 196.380 ;
        RECT 126.400 195.765 126.730 196.560 ;
        RECT 127.065 196.445 127.235 197.645 ;
        RECT 128.080 197.615 128.250 197.765 ;
        RECT 127.495 197.490 128.250 197.615 ;
        RECT 127.405 197.445 128.250 197.490 ;
        RECT 127.405 197.325 127.675 197.445 ;
        RECT 127.405 196.750 127.575 197.325 ;
        RECT 127.805 196.885 128.215 197.190 ;
        RECT 128.505 197.155 128.715 197.555 ;
        RECT 128.385 196.945 128.715 197.155 ;
        RECT 128.960 197.155 129.180 197.555 ;
        RECT 129.655 197.380 130.110 198.145 ;
        RECT 130.285 197.420 130.575 198.145 ;
        RECT 130.750 197.325 131.045 198.145 ;
        RECT 131.215 197.595 131.435 197.975 ;
        RECT 131.605 197.785 132.455 198.145 ;
        RECT 128.960 196.945 129.435 197.155 ;
        RECT 129.625 196.955 130.115 197.155 ;
        RECT 127.405 196.715 127.605 196.750 ;
        RECT 128.935 196.715 130.110 196.775 ;
        RECT 127.405 196.605 130.110 196.715 ;
        RECT 127.465 196.545 129.265 196.605 ;
        RECT 128.935 196.515 129.265 196.545 ;
        RECT 127.065 195.765 127.325 196.445 ;
        RECT 127.495 195.595 127.745 196.375 ;
        RECT 127.995 196.345 128.830 196.355 ;
        RECT 129.420 196.345 129.605 196.435 ;
        RECT 127.995 196.145 129.605 196.345 ;
        RECT 127.995 195.765 128.245 196.145 ;
        RECT 129.375 196.105 129.605 196.145 ;
        RECT 129.855 195.985 130.110 196.605 ;
        RECT 128.415 195.595 128.770 195.975 ;
        RECT 129.775 195.765 130.110 195.985 ;
        RECT 130.285 195.595 130.575 196.760 ;
        RECT 130.750 195.595 131.045 196.740 ;
        RECT 131.215 195.895 131.445 197.595 ;
        RECT 132.935 197.535 133.265 197.955 ;
        RECT 133.470 197.705 133.745 198.145 ;
        RECT 133.915 197.535 134.245 197.955 ;
        RECT 131.660 197.355 134.245 197.535 ;
        RECT 134.425 197.495 134.685 197.940 ;
        RECT 134.935 197.665 135.105 198.145 ;
        RECT 135.275 197.635 135.625 197.965 ;
        RECT 135.860 197.665 136.030 198.145 ;
        RECT 131.660 196.740 131.970 197.355 ;
        RECT 134.425 197.325 135.105 197.495 ;
        RECT 132.140 196.955 132.470 197.185 ;
        RECT 132.640 196.955 133.110 197.185 ;
        RECT 133.280 197.125 133.730 197.185 ;
        RECT 133.280 196.955 133.735 197.125 ;
        RECT 133.920 196.955 134.255 197.185 ;
        RECT 131.660 196.570 134.245 196.740 ;
        RECT 134.425 196.590 134.765 197.155 ;
        RECT 131.660 195.595 131.915 196.400 ;
        RECT 132.115 196.210 133.455 196.390 ;
        RECT 132.115 195.765 132.445 196.210 ;
        RECT 132.615 195.595 132.890 196.040 ;
        RECT 133.125 195.765 133.455 196.210 ;
        RECT 133.915 195.905 134.245 196.570 ;
        RECT 134.935 196.420 135.105 197.325 ;
        RECT 135.275 196.735 135.445 197.635 ;
        RECT 136.330 197.575 136.500 197.925 ;
        RECT 136.670 197.745 137.000 198.145 ;
        RECT 137.170 197.625 137.425 197.925 ;
        RECT 137.170 197.575 137.475 197.625 ;
        RECT 136.330 197.495 137.475 197.575 ;
        RECT 135.765 197.465 137.475 197.495 ;
        RECT 135.615 197.405 137.475 197.465 ;
        RECT 135.615 197.325 136.500 197.405 ;
        RECT 135.615 197.295 135.935 197.325 ;
        RECT 135.615 196.905 135.785 197.295 ;
        RECT 135.275 196.530 135.670 196.735 ;
        RECT 136.035 196.615 136.570 197.155 ;
        RECT 136.830 196.905 137.130 197.235 ;
        RECT 136.830 196.445 137.000 196.905 ;
        RECT 137.305 196.735 137.475 197.405 ;
        RECT 138.565 197.395 139.775 198.145 ;
        RECT 134.425 196.360 135.105 196.420 ;
        RECT 135.890 196.360 137.000 196.445 ;
        RECT 134.425 196.275 137.000 196.360 ;
        RECT 137.170 196.305 137.475 196.735 ;
        RECT 138.565 196.685 139.085 197.225 ;
        RECT 139.255 196.855 139.775 197.395 ;
        RECT 134.425 196.190 136.060 196.275 ;
        RECT 134.425 196.010 134.685 196.190 ;
        RECT 134.890 195.595 135.250 196.020 ;
        RECT 135.765 195.595 136.095 196.020 ;
        RECT 136.275 195.865 137.475 196.105 ;
        RECT 138.565 195.595 139.775 196.685 ;
        RECT 27.160 195.425 139.860 195.595 ;
        RECT 27.245 194.335 28.455 195.425 ;
        RECT 27.245 193.625 27.765 194.165 ;
        RECT 27.935 193.795 28.455 194.335 ;
        RECT 28.630 194.275 28.890 195.425 ;
        RECT 29.065 194.350 29.320 195.255 ;
        RECT 29.490 194.665 29.820 195.425 ;
        RECT 30.035 194.495 30.205 195.255 ;
        RECT 30.465 194.990 35.810 195.425 ;
        RECT 27.245 192.875 28.455 193.625 ;
        RECT 28.630 192.875 28.890 193.715 ;
        RECT 29.065 193.620 29.235 194.350 ;
        RECT 29.490 194.325 30.205 194.495 ;
        RECT 29.490 194.115 29.660 194.325 ;
        RECT 29.405 193.785 29.660 194.115 ;
        RECT 29.065 193.045 29.320 193.620 ;
        RECT 29.490 193.595 29.660 193.785 ;
        RECT 29.940 193.775 30.295 194.145 ;
        RECT 29.490 193.425 30.205 193.595 ;
        RECT 29.490 192.875 29.820 193.255 ;
        RECT 30.035 193.045 30.205 193.425 ;
        RECT 32.050 193.420 32.390 194.250 ;
        RECT 33.870 193.740 34.220 194.990 ;
        RECT 35.985 194.335 39.495 195.425 ;
        RECT 35.985 193.645 37.635 194.165 ;
        RECT 37.805 193.815 39.495 194.335 ;
        RECT 40.125 194.260 40.415 195.425 ;
        RECT 40.585 194.245 40.905 195.425 ;
        RECT 41.075 194.405 41.275 195.195 ;
        RECT 41.600 194.595 41.985 195.255 ;
        RECT 42.380 194.665 43.165 195.425 ;
        RECT 41.575 194.495 41.985 194.595 ;
        RECT 41.075 194.235 41.405 194.405 ;
        RECT 41.575 194.285 43.185 194.495 ;
        RECT 41.225 194.115 41.405 194.235 ;
        RECT 40.585 193.865 41.050 194.065 ;
        RECT 41.225 193.865 41.555 194.115 ;
        RECT 41.725 194.065 42.190 194.115 ;
        RECT 41.725 193.895 42.195 194.065 ;
        RECT 41.725 193.865 42.190 193.895 ;
        RECT 42.385 193.865 42.740 194.115 ;
        RECT 42.910 193.685 43.185 194.285 ;
        RECT 30.465 192.875 35.810 193.420 ;
        RECT 35.985 192.875 39.495 193.645 ;
        RECT 40.125 192.875 40.415 193.600 ;
        RECT 40.585 193.485 41.765 193.655 ;
        RECT 40.585 193.070 40.925 193.485 ;
        RECT 41.095 192.875 41.265 193.315 ;
        RECT 41.435 193.265 41.765 193.485 ;
        RECT 41.935 193.505 43.185 193.685 ;
        RECT 41.935 193.435 42.300 193.505 ;
        RECT 41.435 193.085 42.685 193.265 ;
        RECT 42.955 192.875 43.125 193.335 ;
        RECT 43.355 193.155 43.635 195.255 ;
        RECT 44.305 194.965 44.520 195.425 ;
        RECT 44.690 194.795 45.020 195.255 ;
        RECT 43.850 194.625 45.020 194.795 ;
        RECT 45.190 194.625 45.440 195.425 ;
        RECT 43.850 193.335 44.220 194.625 ;
        RECT 45.650 194.455 45.930 194.615 ;
        RECT 44.595 194.285 45.930 194.455 ;
        RECT 46.105 194.335 47.315 195.425 ;
        RECT 44.595 194.115 44.765 194.285 ;
        RECT 44.390 193.865 44.765 194.115 ;
        RECT 44.935 193.865 45.410 194.105 ;
        RECT 45.580 193.865 45.930 194.105 ;
        RECT 44.595 193.695 44.765 193.865 ;
        RECT 44.595 193.525 45.930 193.695 ;
        RECT 43.850 193.045 44.600 193.335 ;
        RECT 45.110 192.875 45.440 193.335 ;
        RECT 45.660 193.315 45.930 193.525 ;
        RECT 46.105 193.625 46.625 194.165 ;
        RECT 46.795 193.795 47.315 194.335 ;
        RECT 47.495 194.815 47.825 195.245 ;
        RECT 48.005 194.985 48.200 195.425 ;
        RECT 48.370 194.815 48.700 195.245 ;
        RECT 47.495 194.645 48.700 194.815 ;
        RECT 47.495 194.315 48.390 194.645 ;
        RECT 48.870 194.475 49.145 195.245 ;
        RECT 48.560 194.285 49.145 194.475 ;
        RECT 49.325 194.335 52.835 195.425 ;
        RECT 47.500 193.785 47.795 194.115 ;
        RECT 47.975 193.785 48.390 194.115 ;
        RECT 46.105 192.875 47.315 193.625 ;
        RECT 47.495 192.875 47.795 193.605 ;
        RECT 47.975 193.165 48.205 193.785 ;
        RECT 48.560 193.615 48.735 194.285 ;
        RECT 48.405 193.435 48.735 193.615 ;
        RECT 48.905 193.465 49.145 194.115 ;
        RECT 49.325 193.645 50.975 194.165 ;
        RECT 51.145 193.815 52.835 194.335 ;
        RECT 53.005 194.285 53.390 195.245 ;
        RECT 53.605 194.625 53.895 195.425 ;
        RECT 54.065 195.085 55.430 195.255 ;
        RECT 54.065 194.455 54.235 195.085 ;
        RECT 53.560 194.285 54.235 194.455 ;
        RECT 48.405 193.055 48.630 193.435 ;
        RECT 48.800 192.875 49.130 193.265 ;
        RECT 49.325 192.875 52.835 193.645 ;
        RECT 53.005 193.615 53.180 194.285 ;
        RECT 53.560 194.115 53.730 194.285 ;
        RECT 54.405 194.115 54.730 194.915 ;
        RECT 55.100 194.875 55.430 195.085 ;
        RECT 55.100 194.625 56.055 194.875 ;
        RECT 53.365 193.865 53.730 194.115 ;
        RECT 53.925 193.865 54.175 194.115 ;
        RECT 53.365 193.785 53.555 193.865 ;
        RECT 53.925 193.785 54.095 193.865 ;
        RECT 54.385 193.785 54.730 194.115 ;
        RECT 54.900 193.785 55.175 194.450 ;
        RECT 55.360 193.785 55.715 194.450 ;
        RECT 55.885 193.615 56.055 194.625 ;
        RECT 56.225 194.285 56.515 195.425 ;
        RECT 56.685 194.335 57.895 195.425 ;
        RECT 56.240 193.785 56.515 194.115 ;
        RECT 53.005 193.045 53.515 193.615 ;
        RECT 54.060 193.445 55.460 193.615 ;
        RECT 53.685 192.875 53.855 193.435 ;
        RECT 54.060 193.045 54.390 193.445 ;
        RECT 54.565 192.875 54.895 193.275 ;
        RECT 55.130 193.255 55.460 193.445 ;
        RECT 55.630 193.425 56.055 193.615 ;
        RECT 56.685 193.625 57.205 194.165 ;
        RECT 57.375 193.795 57.895 194.335 ;
        RECT 58.070 194.285 58.390 195.425 ;
        RECT 58.570 194.115 58.765 195.165 ;
        RECT 58.945 194.575 59.275 195.255 ;
        RECT 59.475 194.625 59.730 195.425 ;
        RECT 58.945 194.295 59.295 194.575 ;
        RECT 58.130 194.065 58.390 194.115 ;
        RECT 58.125 193.895 58.390 194.065 ;
        RECT 58.130 193.785 58.390 193.895 ;
        RECT 58.570 193.785 58.955 194.115 ;
        RECT 59.125 193.915 59.295 194.295 ;
        RECT 59.485 194.085 59.730 194.445 ;
        RECT 59.905 194.335 61.575 195.425 ;
        RECT 62.310 194.965 62.480 195.425 ;
        RECT 62.650 194.795 62.980 195.255 ;
        RECT 59.125 193.745 59.645 193.915 ;
        RECT 59.475 193.725 59.645 193.745 ;
        RECT 56.225 193.255 56.515 193.525 ;
        RECT 55.130 193.045 56.515 193.255 ;
        RECT 56.685 192.875 57.895 193.625 ;
        RECT 58.070 193.405 59.285 193.575 ;
        RECT 58.070 193.055 58.360 193.405 ;
        RECT 58.555 192.875 58.885 193.235 ;
        RECT 59.055 193.100 59.285 193.405 ;
        RECT 59.475 193.555 59.675 193.725 ;
        RECT 59.905 193.645 60.655 194.165 ;
        RECT 60.825 193.815 61.575 194.335 ;
        RECT 62.205 194.625 62.980 194.795 ;
        RECT 63.150 194.625 63.320 195.425 ;
        RECT 59.475 193.180 59.645 193.555 ;
        RECT 59.905 192.875 61.575 193.645 ;
        RECT 62.205 193.615 62.635 194.625 ;
        RECT 63.905 194.455 64.265 194.630 ;
        RECT 62.805 194.285 64.265 194.455 ;
        RECT 64.505 194.335 65.715 195.425 ;
        RECT 62.805 193.785 62.975 194.285 ;
        RECT 62.205 193.445 62.900 193.615 ;
        RECT 63.145 193.555 63.555 194.115 ;
        RECT 62.230 192.875 62.560 193.275 ;
        RECT 62.730 193.175 62.900 193.445 ;
        RECT 63.725 193.385 63.905 194.285 ;
        RECT 64.075 193.725 64.270 194.115 ;
        RECT 64.075 193.555 64.275 193.725 ;
        RECT 64.505 193.625 65.025 194.165 ;
        RECT 65.195 193.795 65.715 194.335 ;
        RECT 65.885 194.260 66.175 195.425 ;
        RECT 66.345 194.315 66.605 195.255 ;
        RECT 66.775 195.025 67.105 195.425 ;
        RECT 68.250 195.160 68.505 195.255 ;
        RECT 67.365 194.990 68.505 195.160 ;
        RECT 68.675 195.045 69.005 195.215 ;
        RECT 67.365 194.765 67.535 194.990 ;
        RECT 66.775 194.595 67.535 194.765 ;
        RECT 68.250 194.855 68.505 194.990 ;
        RECT 63.070 192.875 63.385 193.385 ;
        RECT 63.615 193.045 63.905 193.385 ;
        RECT 64.075 192.875 64.315 193.385 ;
        RECT 64.505 192.875 65.715 193.625 ;
        RECT 66.345 193.600 66.520 194.315 ;
        RECT 66.775 194.115 66.945 194.595 ;
        RECT 67.800 194.505 67.970 194.695 ;
        RECT 68.250 194.685 68.660 194.855 ;
        RECT 66.690 193.785 66.945 194.115 ;
        RECT 67.170 193.785 67.500 194.405 ;
        RECT 67.800 194.335 68.320 194.505 ;
        RECT 67.670 193.785 67.960 194.165 ;
        RECT 68.150 193.615 68.320 194.335 ;
        RECT 65.885 192.875 66.175 193.600 ;
        RECT 66.345 193.045 66.605 193.600 ;
        RECT 67.440 193.445 68.320 193.615 ;
        RECT 68.490 193.660 68.660 194.685 ;
        RECT 68.835 194.795 69.005 195.045 ;
        RECT 69.175 194.965 69.425 195.425 ;
        RECT 69.595 194.795 69.775 195.255 ;
        RECT 68.835 194.625 69.775 194.795 ;
        RECT 70.045 194.585 70.300 195.255 ;
        RECT 70.470 194.665 70.800 195.425 ;
        RECT 70.970 194.825 71.220 195.255 ;
        RECT 71.390 195.005 71.745 195.425 ;
        RECT 71.935 195.085 73.105 195.255 ;
        RECT 71.935 195.045 72.265 195.085 ;
        RECT 72.375 194.825 72.605 194.915 ;
        RECT 70.970 194.585 72.605 194.825 ;
        RECT 72.775 194.585 73.105 195.085 ;
        RECT 68.860 194.145 69.340 194.445 ;
        RECT 68.490 193.490 68.840 193.660 ;
        RECT 69.080 193.555 69.340 194.145 ;
        RECT 69.540 193.555 69.800 194.445 ;
        RECT 66.775 192.875 67.205 193.320 ;
        RECT 67.440 193.045 67.610 193.445 ;
        RECT 67.780 192.875 68.500 193.275 ;
        RECT 68.670 193.045 68.840 193.490 ;
        RECT 70.045 193.455 70.215 194.585 ;
        RECT 73.275 194.415 73.445 195.255 ;
        RECT 70.385 194.245 73.445 194.415 ;
        RECT 73.715 194.475 73.990 195.245 ;
        RECT 74.160 194.815 74.490 195.245 ;
        RECT 74.660 194.985 74.855 195.425 ;
        RECT 75.035 194.815 75.365 195.245 ;
        RECT 74.160 194.645 75.365 194.815 ;
        RECT 73.715 194.285 74.300 194.475 ;
        RECT 74.470 194.315 75.365 194.645 ;
        RECT 75.545 194.335 79.055 195.425 ;
        RECT 70.385 193.695 70.555 194.245 ;
        RECT 70.785 193.865 71.150 194.065 ;
        RECT 71.320 193.865 71.650 194.065 ;
        RECT 70.385 193.525 71.185 193.695 ;
        RECT 69.415 192.875 69.815 193.385 ;
        RECT 70.045 193.375 70.230 193.455 ;
        RECT 70.045 193.045 70.300 193.375 ;
        RECT 70.515 192.875 70.845 193.355 ;
        RECT 71.015 193.295 71.185 193.525 ;
        RECT 71.365 193.465 71.650 193.865 ;
        RECT 71.920 193.865 72.395 194.065 ;
        RECT 72.565 193.865 73.010 194.065 ;
        RECT 73.180 193.865 73.530 194.075 ;
        RECT 71.920 193.465 72.200 193.865 ;
        RECT 72.380 193.525 73.445 193.695 ;
        RECT 72.380 193.295 72.550 193.525 ;
        RECT 71.015 193.045 72.550 193.295 ;
        RECT 72.775 192.875 73.105 193.355 ;
        RECT 73.275 193.045 73.445 193.525 ;
        RECT 73.715 193.465 73.955 194.115 ;
        RECT 74.125 193.615 74.300 194.285 ;
        RECT 74.470 193.785 74.885 194.115 ;
        RECT 75.065 193.785 75.360 194.115 ;
        RECT 74.125 193.435 74.455 193.615 ;
        RECT 73.730 192.875 74.060 193.265 ;
        RECT 74.230 193.055 74.455 193.435 ;
        RECT 74.655 193.165 74.885 193.785 ;
        RECT 75.545 193.645 77.195 194.165 ;
        RECT 77.365 193.815 79.055 194.335 ;
        RECT 79.690 194.285 80.010 195.425 ;
        RECT 80.190 194.115 80.385 195.165 ;
        RECT 80.565 194.575 80.895 195.255 ;
        RECT 81.095 194.625 81.350 195.425 ;
        RECT 80.565 194.295 80.915 194.575 ;
        RECT 82.610 194.460 82.940 195.255 ;
        RECT 83.110 194.640 83.350 195.425 ;
        RECT 83.910 194.835 84.665 195.255 ;
        RECT 83.520 194.665 84.985 194.835 ;
        RECT 83.520 194.460 83.690 194.665 ;
        RECT 79.750 194.065 80.010 194.115 ;
        RECT 79.745 193.895 80.010 194.065 ;
        RECT 79.750 193.785 80.010 193.895 ;
        RECT 80.190 193.785 80.575 194.115 ;
        RECT 80.745 193.915 80.915 194.295 ;
        RECT 81.105 194.085 81.350 194.445 ;
        RECT 82.610 194.285 83.690 194.460 ;
        RECT 82.905 194.235 83.690 194.285 ;
        RECT 80.745 193.745 81.265 193.915 ;
        RECT 82.445 193.765 82.705 194.115 ;
        RECT 75.065 192.875 75.365 193.605 ;
        RECT 75.545 192.875 79.055 193.645 ;
        RECT 79.690 193.405 80.905 193.575 ;
        RECT 79.690 193.055 79.980 193.405 ;
        RECT 80.175 192.875 80.505 193.235 ;
        RECT 80.675 193.100 80.905 193.405 ;
        RECT 81.095 193.180 81.265 193.745 ;
        RECT 82.905 193.595 83.075 194.235 ;
        RECT 83.860 194.065 84.150 194.495 ;
        RECT 83.245 193.865 83.590 194.065 ;
        RECT 83.760 193.865 84.150 194.065 ;
        RECT 84.340 194.075 84.645 194.495 ;
        RECT 84.815 194.415 84.985 194.665 ;
        RECT 85.155 194.585 85.485 195.425 ;
        RECT 85.655 194.835 85.905 195.255 ;
        RECT 86.075 195.005 86.415 195.425 ;
        RECT 85.655 194.665 86.415 194.835 ;
        RECT 84.815 194.245 85.775 194.415 ;
        RECT 85.605 194.075 85.775 194.245 ;
        RECT 84.340 193.865 84.825 194.075 ;
        RECT 84.995 193.865 85.435 194.075 ;
        RECT 85.605 193.865 85.935 194.075 ;
        RECT 86.105 193.695 86.415 194.665 ;
        RECT 86.590 194.555 86.855 195.255 ;
        RECT 87.025 194.725 87.355 195.425 ;
        RECT 87.525 194.555 88.195 195.255 ;
        RECT 88.700 194.725 89.130 195.425 ;
        RECT 89.310 194.865 89.500 195.255 ;
        RECT 89.670 195.045 90.000 195.425 ;
        RECT 89.310 194.695 90.040 194.865 ;
        RECT 86.590 194.300 89.165 194.555 ;
        RECT 86.585 193.785 86.860 194.115 ;
        RECT 82.530 193.425 83.075 193.595 ;
        RECT 83.445 193.525 85.145 193.695 ;
        RECT 83.445 193.435 83.830 193.525 ;
        RECT 82.530 193.045 82.860 193.425 ;
        RECT 83.030 193.085 84.215 193.255 ;
        RECT 84.475 192.875 84.645 193.345 ;
        RECT 84.815 193.060 85.145 193.525 ;
        RECT 85.315 192.875 85.485 193.695 ;
        RECT 85.655 193.525 86.415 193.695 ;
        RECT 87.030 193.615 87.210 194.300 ;
        RECT 88.995 194.115 89.165 194.300 ;
        RECT 87.380 193.785 87.740 194.115 ;
        RECT 88.030 194.065 88.320 194.115 ;
        RECT 88.025 193.895 88.320 194.065 ;
        RECT 88.030 193.785 88.320 193.895 ;
        RECT 88.490 193.785 88.825 194.115 ;
        RECT 88.995 193.785 89.675 194.115 ;
        RECT 85.655 193.055 85.985 193.525 ;
        RECT 86.155 192.875 86.325 193.355 ;
        RECT 86.595 193.215 87.210 193.615 ;
        RECT 87.380 193.425 88.650 193.615 ;
        RECT 89.845 193.575 90.040 194.695 ;
        RECT 90.265 194.335 91.475 195.425 ;
        RECT 89.220 193.405 90.040 193.575 ;
        RECT 90.265 193.625 90.785 194.165 ;
        RECT 90.955 193.795 91.475 194.335 ;
        RECT 91.645 194.260 91.935 195.425 ;
        RECT 92.195 194.680 92.465 195.425 ;
        RECT 93.095 195.420 99.370 195.425 ;
        RECT 92.635 194.510 92.925 195.250 ;
        RECT 93.095 194.695 93.350 195.420 ;
        RECT 93.535 194.525 93.795 195.250 ;
        RECT 93.965 194.695 94.210 195.420 ;
        RECT 94.395 194.525 94.655 195.250 ;
        RECT 94.825 194.695 95.070 195.420 ;
        RECT 95.255 194.525 95.515 195.250 ;
        RECT 95.685 194.695 95.930 195.420 ;
        RECT 96.100 194.525 96.360 195.250 ;
        RECT 96.530 194.695 96.790 195.420 ;
        RECT 96.960 194.525 97.220 195.250 ;
        RECT 97.390 194.695 97.650 195.420 ;
        RECT 97.820 194.525 98.080 195.250 ;
        RECT 98.250 194.695 98.510 195.420 ;
        RECT 98.680 194.525 98.940 195.250 ;
        RECT 99.110 194.625 99.370 195.420 ;
        RECT 93.535 194.510 98.940 194.525 ;
        RECT 92.195 194.405 98.940 194.510 ;
        RECT 92.165 194.285 98.940 194.405 ;
        RECT 92.165 194.235 93.360 194.285 ;
        RECT 92.195 193.695 93.360 194.235 ;
        RECT 99.540 194.115 99.790 195.250 ;
        RECT 99.970 194.615 100.230 195.425 ;
        RECT 100.405 194.115 100.650 195.255 ;
        RECT 100.830 194.615 101.125 195.425 ;
        RECT 102.280 194.555 102.565 195.425 ;
        RECT 102.735 194.795 102.995 195.255 ;
        RECT 103.170 194.965 103.425 195.425 ;
        RECT 103.595 194.795 103.855 195.255 ;
        RECT 102.735 194.625 103.855 194.795 ;
        RECT 104.025 194.625 104.335 195.425 ;
        RECT 102.735 194.375 102.995 194.625 ;
        RECT 104.505 194.455 104.815 195.255 ;
        RECT 105.035 194.965 105.285 195.425 ;
        RECT 105.495 194.795 105.665 195.255 ;
        RECT 102.240 194.205 102.995 194.375 ;
        RECT 103.785 194.285 104.815 194.455 ;
        RECT 93.530 193.865 100.650 194.115 ;
        RECT 86.595 193.045 86.930 193.215 ;
        RECT 87.890 192.875 88.225 193.255 ;
        RECT 88.815 192.875 89.050 193.315 ;
        RECT 89.220 193.045 89.550 193.405 ;
        RECT 89.720 192.875 90.050 193.235 ;
        RECT 90.265 192.875 91.475 193.625 ;
        RECT 91.645 192.875 91.935 193.600 ;
        RECT 92.195 193.525 98.940 193.695 ;
        RECT 92.195 192.875 92.495 193.355 ;
        RECT 92.665 193.070 92.925 193.525 ;
        RECT 93.095 192.875 93.355 193.355 ;
        RECT 93.535 193.070 93.795 193.525 ;
        RECT 93.965 192.875 94.215 193.355 ;
        RECT 94.395 193.070 94.655 193.525 ;
        RECT 94.825 192.875 95.075 193.355 ;
        RECT 95.255 193.070 95.515 193.525 ;
        RECT 95.685 192.875 95.930 193.355 ;
        RECT 96.100 193.070 96.375 193.525 ;
        RECT 96.545 192.875 96.790 193.355 ;
        RECT 96.960 193.070 97.220 193.525 ;
        RECT 97.390 192.875 97.650 193.355 ;
        RECT 97.820 193.070 98.080 193.525 ;
        RECT 98.250 192.875 98.510 193.355 ;
        RECT 98.680 193.070 98.940 193.525 ;
        RECT 99.110 192.875 99.370 193.435 ;
        RECT 99.540 193.055 99.790 193.865 ;
        RECT 99.970 192.875 100.230 193.400 ;
        RECT 100.400 193.055 100.650 193.865 ;
        RECT 100.820 193.555 101.135 194.115 ;
        RECT 102.240 193.695 102.645 194.205 ;
        RECT 103.785 194.035 103.955 194.285 ;
        RECT 102.815 193.865 103.955 194.035 ;
        RECT 102.240 193.525 103.890 193.695 ;
        RECT 104.125 193.545 104.475 194.115 ;
        RECT 100.830 192.875 101.135 193.385 ;
        RECT 102.285 192.875 102.565 193.355 ;
        RECT 102.735 193.135 102.995 193.525 ;
        RECT 103.170 192.875 103.425 193.355 ;
        RECT 103.595 193.135 103.890 193.525 ;
        RECT 104.645 193.375 104.815 194.285 ;
        RECT 104.990 194.625 105.665 194.795 ;
        RECT 105.835 194.625 106.085 195.425 ;
        RECT 106.255 194.795 106.505 195.215 ;
        RECT 106.715 194.965 107.045 195.425 ;
        RECT 107.235 194.795 107.485 195.215 ;
        RECT 106.255 194.625 107.545 194.795 ;
        RECT 104.990 193.675 105.245 194.625 ;
        RECT 107.775 194.455 107.945 195.255 ;
        RECT 108.215 194.615 108.510 195.425 ;
        RECT 105.455 194.285 107.945 194.455 ;
        RECT 105.455 194.035 105.625 194.285 ;
        RECT 105.455 193.865 105.785 194.035 ;
        RECT 105.965 193.785 106.295 194.115 ;
        RECT 106.525 194.035 106.695 194.050 ;
        RECT 106.525 193.865 106.855 194.035 ;
        RECT 104.990 193.505 105.665 193.675 ;
        RECT 105.965 193.550 106.170 193.785 ;
        RECT 106.525 193.655 106.695 193.865 ;
        RECT 107.085 193.660 107.255 194.115 ;
        RECT 104.070 192.875 104.345 193.355 ;
        RECT 104.515 193.045 104.815 193.375 ;
        RECT 105.495 193.385 105.665 193.505 ;
        RECT 106.430 193.485 106.695 193.655 ;
        RECT 106.865 193.490 107.255 193.660 ;
        RECT 106.430 193.385 106.600 193.485 ;
        RECT 104.990 192.875 105.245 193.335 ;
        RECT 105.495 193.215 105.675 193.385 ;
        RECT 105.915 193.255 106.085 193.335 ;
        RECT 105.495 193.045 105.665 193.215 ;
        RECT 105.855 192.875 106.185 193.255 ;
        RECT 106.425 193.215 106.600 193.385 ;
        RECT 106.430 193.190 106.600 193.215 ;
        RECT 106.865 193.205 107.075 193.490 ;
        RECT 107.435 193.295 107.605 194.285 ;
        RECT 108.690 194.115 108.935 195.255 ;
        RECT 109.110 194.615 109.370 195.425 ;
        RECT 109.970 195.420 116.245 195.425 ;
        RECT 109.550 194.115 109.800 195.250 ;
        RECT 109.970 194.625 110.230 195.420 ;
        RECT 110.400 194.525 110.660 195.250 ;
        RECT 110.830 194.695 111.090 195.420 ;
        RECT 111.260 194.525 111.520 195.250 ;
        RECT 111.690 194.695 111.950 195.420 ;
        RECT 112.120 194.525 112.380 195.250 ;
        RECT 112.550 194.695 112.810 195.420 ;
        RECT 112.980 194.525 113.240 195.250 ;
        RECT 113.410 194.695 113.655 195.420 ;
        RECT 113.825 194.525 114.085 195.250 ;
        RECT 114.270 194.695 114.515 195.420 ;
        RECT 114.685 194.525 114.945 195.250 ;
        RECT 115.130 194.695 115.375 195.420 ;
        RECT 115.545 194.525 115.805 195.250 ;
        RECT 115.990 194.695 116.245 195.420 ;
        RECT 110.400 194.510 115.805 194.525 ;
        RECT 116.415 194.510 116.705 195.250 ;
        RECT 116.875 194.680 117.145 195.425 ;
        RECT 110.400 194.285 117.145 194.510 ;
        RECT 107.795 193.545 107.990 194.115 ;
        RECT 108.205 193.555 108.520 194.115 ;
        RECT 108.690 193.865 115.810 194.115 ;
        RECT 115.980 194.065 117.145 194.285 ;
        RECT 117.405 194.260 117.695 195.425 ;
        RECT 117.875 194.615 118.170 195.425 ;
        RECT 118.350 194.115 118.595 195.255 ;
        RECT 118.770 194.615 119.030 195.425 ;
        RECT 119.630 195.420 125.905 195.425 ;
        RECT 119.210 194.115 119.460 195.250 ;
        RECT 119.630 194.625 119.890 195.420 ;
        RECT 120.060 194.525 120.320 195.250 ;
        RECT 120.490 194.695 120.750 195.420 ;
        RECT 120.920 194.525 121.180 195.250 ;
        RECT 121.350 194.695 121.610 195.420 ;
        RECT 121.780 194.525 122.040 195.250 ;
        RECT 122.210 194.695 122.470 195.420 ;
        RECT 122.640 194.525 122.900 195.250 ;
        RECT 123.070 194.695 123.315 195.420 ;
        RECT 123.485 194.525 123.745 195.250 ;
        RECT 123.930 194.695 124.175 195.420 ;
        RECT 124.345 194.525 124.605 195.250 ;
        RECT 124.790 194.695 125.035 195.420 ;
        RECT 125.205 194.525 125.465 195.250 ;
        RECT 125.650 194.695 125.905 195.420 ;
        RECT 120.060 194.510 125.465 194.525 ;
        RECT 126.075 194.510 126.365 195.250 ;
        RECT 126.535 194.680 126.805 195.425 ;
        RECT 127.075 194.615 127.370 195.425 ;
        RECT 120.060 194.285 126.805 194.510 ;
        RECT 115.980 193.895 117.175 194.065 ;
        RECT 107.275 193.125 107.605 193.295 ;
        RECT 107.360 193.045 107.605 193.125 ;
        RECT 107.775 192.875 108.035 193.355 ;
        RECT 108.205 192.875 108.510 193.385 ;
        RECT 108.690 193.055 108.940 193.865 ;
        RECT 109.110 192.875 109.370 193.400 ;
        RECT 109.550 193.055 109.800 193.865 ;
        RECT 115.980 193.695 117.145 193.895 ;
        RECT 110.400 193.525 117.145 193.695 ;
        RECT 109.970 192.875 110.230 193.435 ;
        RECT 110.400 193.070 110.660 193.525 ;
        RECT 110.830 192.875 111.090 193.355 ;
        RECT 111.260 193.070 111.520 193.525 ;
        RECT 111.690 192.875 111.950 193.355 ;
        RECT 112.120 193.070 112.380 193.525 ;
        RECT 112.550 192.875 112.795 193.355 ;
        RECT 112.965 193.070 113.240 193.525 ;
        RECT 113.410 192.875 113.655 193.355 ;
        RECT 113.825 193.070 114.085 193.525 ;
        RECT 114.265 192.875 114.515 193.355 ;
        RECT 114.685 193.070 114.945 193.525 ;
        RECT 115.125 192.875 115.375 193.355 ;
        RECT 115.545 193.070 115.805 193.525 ;
        RECT 115.985 192.875 116.245 193.355 ;
        RECT 116.415 193.070 116.675 193.525 ;
        RECT 116.845 192.875 117.145 193.355 ;
        RECT 117.405 192.875 117.695 193.600 ;
        RECT 117.865 193.555 118.180 194.115 ;
        RECT 118.350 193.865 125.470 194.115 ;
        RECT 117.865 192.875 118.170 193.385 ;
        RECT 118.350 193.055 118.600 193.865 ;
        RECT 118.770 192.875 119.030 193.400 ;
        RECT 119.210 193.055 119.460 193.865 ;
        RECT 125.640 193.695 126.805 194.285 ;
        RECT 127.550 194.115 127.795 195.255 ;
        RECT 127.970 194.615 128.230 195.425 ;
        RECT 128.830 195.420 135.105 195.425 ;
        RECT 128.410 194.115 128.660 195.250 ;
        RECT 128.830 194.625 129.090 195.420 ;
        RECT 129.260 194.525 129.520 195.250 ;
        RECT 129.690 194.695 129.950 195.420 ;
        RECT 130.120 194.525 130.380 195.250 ;
        RECT 130.550 194.695 130.810 195.420 ;
        RECT 130.980 194.525 131.240 195.250 ;
        RECT 131.410 194.695 131.670 195.420 ;
        RECT 131.840 194.525 132.100 195.250 ;
        RECT 132.270 194.695 132.515 195.420 ;
        RECT 132.685 194.525 132.945 195.250 ;
        RECT 133.130 194.695 133.375 195.420 ;
        RECT 133.545 194.525 133.805 195.250 ;
        RECT 133.990 194.695 134.235 195.420 ;
        RECT 134.405 194.525 134.665 195.250 ;
        RECT 134.850 194.695 135.105 195.420 ;
        RECT 129.260 194.510 134.665 194.525 ;
        RECT 135.275 194.510 135.565 195.250 ;
        RECT 135.735 194.680 136.005 195.425 ;
        RECT 129.260 194.285 136.005 194.510 ;
        RECT 136.815 194.495 136.985 195.255 ;
        RECT 137.200 194.665 137.530 195.425 ;
        RECT 136.815 194.325 137.530 194.495 ;
        RECT 137.700 194.350 137.955 195.255 ;
        RECT 120.060 193.525 126.805 193.695 ;
        RECT 127.065 193.555 127.380 194.115 ;
        RECT 127.550 193.865 134.670 194.115 ;
        RECT 119.630 192.875 119.890 193.435 ;
        RECT 120.060 193.070 120.320 193.525 ;
        RECT 120.490 192.875 120.750 193.355 ;
        RECT 120.920 193.070 121.180 193.525 ;
        RECT 121.350 192.875 121.610 193.355 ;
        RECT 121.780 193.070 122.040 193.525 ;
        RECT 122.210 192.875 122.455 193.355 ;
        RECT 122.625 193.070 122.900 193.525 ;
        RECT 123.070 192.875 123.315 193.355 ;
        RECT 123.485 193.070 123.745 193.525 ;
        RECT 123.925 192.875 124.175 193.355 ;
        RECT 124.345 193.070 124.605 193.525 ;
        RECT 124.785 192.875 125.035 193.355 ;
        RECT 125.205 193.070 125.465 193.525 ;
        RECT 125.645 192.875 125.905 193.355 ;
        RECT 126.075 193.070 126.335 193.525 ;
        RECT 126.505 192.875 126.805 193.355 ;
        RECT 127.065 192.875 127.370 193.385 ;
        RECT 127.550 193.055 127.800 193.865 ;
        RECT 127.970 192.875 128.230 193.400 ;
        RECT 128.410 193.055 128.660 193.865 ;
        RECT 134.840 193.695 136.005 194.285 ;
        RECT 136.725 193.775 137.080 194.145 ;
        RECT 137.360 194.115 137.530 194.325 ;
        RECT 137.360 193.785 137.615 194.115 ;
        RECT 129.260 193.525 136.005 193.695 ;
        RECT 137.360 193.595 137.530 193.785 ;
        RECT 137.785 193.620 137.955 194.350 ;
        RECT 138.130 194.275 138.390 195.425 ;
        RECT 138.565 194.335 139.775 195.425 ;
        RECT 138.565 193.795 139.085 194.335 ;
        RECT 128.830 192.875 129.090 193.435 ;
        RECT 129.260 193.070 129.520 193.525 ;
        RECT 129.690 192.875 129.950 193.355 ;
        RECT 130.120 193.070 130.380 193.525 ;
        RECT 130.550 192.875 130.810 193.355 ;
        RECT 130.980 193.070 131.240 193.525 ;
        RECT 131.410 192.875 131.655 193.355 ;
        RECT 131.825 193.070 132.100 193.525 ;
        RECT 132.270 192.875 132.515 193.355 ;
        RECT 132.685 193.070 132.945 193.525 ;
        RECT 133.125 192.875 133.375 193.355 ;
        RECT 133.545 193.070 133.805 193.525 ;
        RECT 133.985 192.875 134.235 193.355 ;
        RECT 134.405 193.070 134.665 193.525 ;
        RECT 134.845 192.875 135.105 193.355 ;
        RECT 135.275 193.070 135.535 193.525 ;
        RECT 136.815 193.425 137.530 193.595 ;
        RECT 135.705 192.875 136.005 193.355 ;
        RECT 136.815 193.045 136.985 193.425 ;
        RECT 137.200 192.875 137.530 193.255 ;
        RECT 137.700 193.045 137.955 193.620 ;
        RECT 138.130 192.875 138.390 193.715 ;
        RECT 139.255 193.625 139.775 194.165 ;
        RECT 138.565 192.875 139.775 193.625 ;
        RECT 27.160 192.705 139.860 192.875 ;
        RECT 27.245 191.955 28.455 192.705 ;
        RECT 28.625 192.205 28.885 192.535 ;
        RECT 29.095 192.225 29.370 192.705 ;
        RECT 27.245 191.415 27.765 191.955 ;
        RECT 27.935 191.245 28.455 191.785 ;
        RECT 27.245 190.155 28.455 191.245 ;
        RECT 28.625 191.295 28.795 192.205 ;
        RECT 29.580 192.135 29.785 192.535 ;
        RECT 29.955 192.305 30.290 192.705 ;
        RECT 28.965 191.465 29.325 192.045 ;
        RECT 29.580 191.965 30.265 192.135 ;
        RECT 29.505 191.295 29.755 191.795 ;
        RECT 28.625 191.125 29.755 191.295 ;
        RECT 28.625 190.355 28.895 191.125 ;
        RECT 29.925 190.935 30.265 191.965 ;
        RECT 29.065 190.155 29.395 190.935 ;
        RECT 29.600 190.760 30.265 190.935 ;
        RECT 31.385 192.030 31.645 192.535 ;
        RECT 31.825 192.325 32.155 192.705 ;
        RECT 32.335 192.155 32.505 192.535 ;
        RECT 32.765 192.160 38.110 192.705 ;
        RECT 31.385 191.230 31.555 192.030 ;
        RECT 31.840 191.985 32.505 192.155 ;
        RECT 31.840 191.730 32.010 191.985 ;
        RECT 31.725 191.400 32.010 191.730 ;
        RECT 32.245 191.435 32.575 191.805 ;
        RECT 31.840 191.255 32.010 191.400 ;
        RECT 34.350 191.330 34.690 192.160 ;
        RECT 38.285 191.935 39.955 192.705 ;
        RECT 29.600 190.355 29.785 190.760 ;
        RECT 29.955 190.155 30.290 190.580 ;
        RECT 31.385 190.325 31.655 191.230 ;
        RECT 31.840 191.085 32.505 191.255 ;
        RECT 31.825 190.155 32.155 190.915 ;
        RECT 32.335 190.325 32.505 191.085 ;
        RECT 36.170 190.590 36.520 191.840 ;
        RECT 38.285 191.415 39.035 191.935 ;
        RECT 40.135 191.895 40.405 192.705 ;
        RECT 40.575 191.895 40.905 192.535 ;
        RECT 41.075 191.895 41.315 192.705 ;
        RECT 41.505 191.955 42.715 192.705 ;
        RECT 39.205 191.245 39.955 191.765 ;
        RECT 40.125 191.465 40.475 191.715 ;
        RECT 40.645 191.295 40.815 191.895 ;
        RECT 40.985 191.465 41.335 191.715 ;
        RECT 41.505 191.415 42.025 191.955 ;
        RECT 42.925 191.885 43.155 192.705 ;
        RECT 43.325 191.905 43.655 192.535 ;
        RECT 32.765 190.155 38.110 190.590 ;
        RECT 38.285 190.155 39.955 191.245 ;
        RECT 40.135 190.155 40.465 191.295 ;
        RECT 40.645 191.125 41.325 191.295 ;
        RECT 42.195 191.245 42.715 191.785 ;
        RECT 42.905 191.465 43.235 191.715 ;
        RECT 43.405 191.305 43.655 191.905 ;
        RECT 43.825 191.885 44.035 192.705 ;
        RECT 44.265 191.935 47.775 192.705 ;
        RECT 47.945 191.955 49.155 192.705 ;
        RECT 49.335 191.975 49.635 192.705 ;
        RECT 44.265 191.415 45.915 191.935 ;
        RECT 40.995 190.340 41.325 191.125 ;
        RECT 41.505 190.155 42.715 191.245 ;
        RECT 42.925 190.155 43.155 191.295 ;
        RECT 43.325 190.325 43.655 191.305 ;
        RECT 43.825 190.155 44.035 191.295 ;
        RECT 46.085 191.245 47.775 191.765 ;
        RECT 47.945 191.415 48.465 191.955 ;
        RECT 49.815 191.795 50.045 192.415 ;
        RECT 50.245 192.145 50.470 192.525 ;
        RECT 50.640 192.315 50.970 192.705 ;
        RECT 51.190 192.315 51.520 192.705 ;
        RECT 51.690 192.145 51.915 192.525 ;
        RECT 50.245 191.965 50.575 192.145 ;
        RECT 48.635 191.245 49.155 191.785 ;
        RECT 49.340 191.465 49.635 191.795 ;
        RECT 49.815 191.465 50.230 191.795 ;
        RECT 50.400 191.295 50.575 191.965 ;
        RECT 50.745 191.465 50.985 192.115 ;
        RECT 51.175 191.465 51.415 192.115 ;
        RECT 51.585 191.965 51.915 192.145 ;
        RECT 51.585 191.295 51.760 191.965 ;
        RECT 52.115 191.795 52.345 192.415 ;
        RECT 52.525 191.975 52.825 192.705 ;
        RECT 53.005 191.980 53.295 192.705 ;
        RECT 53.565 191.905 53.735 192.705 ;
        RECT 51.930 191.465 52.345 191.795 ;
        RECT 52.525 191.465 52.820 191.795 ;
        RECT 44.265 190.155 47.775 191.245 ;
        RECT 47.945 190.155 49.155 191.245 ;
        RECT 49.335 190.935 50.230 191.265 ;
        RECT 50.400 191.105 50.985 191.295 ;
        RECT 49.335 190.765 50.540 190.935 ;
        RECT 49.335 190.335 49.665 190.765 ;
        RECT 49.845 190.155 50.040 190.595 ;
        RECT 50.210 190.335 50.540 190.765 ;
        RECT 50.710 190.335 50.985 191.105 ;
        RECT 51.175 191.105 51.760 191.295 ;
        RECT 51.175 190.335 51.450 191.105 ;
        RECT 51.930 190.935 52.825 191.265 ;
        RECT 51.620 190.765 52.825 190.935 ;
        RECT 51.620 190.335 51.950 190.765 ;
        RECT 52.120 190.155 52.315 190.595 ;
        RECT 52.495 190.335 52.825 190.765 ;
        RECT 53.005 190.155 53.295 191.320 ;
        RECT 53.495 190.155 53.745 191.345 ;
        RECT 53.970 190.325 54.185 192.425 ;
        RECT 54.405 192.245 54.585 192.705 ;
        RECT 54.845 192.315 56.110 192.495 ;
        RECT 55.230 192.075 55.595 192.145 ;
        RECT 54.355 191.895 55.595 192.075 ;
        RECT 55.770 192.095 56.110 192.315 ;
        RECT 56.295 192.265 56.465 192.705 ;
        RECT 56.635 192.095 56.970 192.510 ;
        RECT 55.770 191.965 56.970 192.095 ;
        RECT 55.940 191.925 56.970 191.965 ;
        RECT 57.145 192.245 57.705 192.535 ;
        RECT 57.875 192.245 58.125 192.705 ;
        RECT 54.355 191.295 54.635 191.895 ;
        RECT 54.815 191.465 55.170 191.715 ;
        RECT 55.340 191.465 55.805 191.715 ;
        RECT 55.975 191.465 56.305 191.715 ;
        RECT 56.475 191.515 56.970 191.715 ;
        RECT 56.125 191.345 56.305 191.465 ;
        RECT 54.355 191.085 55.955 191.295 ;
        RECT 56.125 191.175 56.480 191.345 ;
        RECT 56.650 191.175 56.970 191.515 ;
        RECT 54.375 190.155 55.175 190.915 ;
        RECT 55.570 190.325 55.955 191.085 ;
        RECT 56.280 190.385 56.480 191.175 ;
        RECT 56.650 190.155 56.970 190.995 ;
        RECT 57.145 190.875 57.395 192.245 ;
        RECT 58.745 192.075 59.075 192.435 ;
        RECT 57.685 191.885 59.075 192.075 ;
        RECT 59.445 191.905 60.140 192.535 ;
        RECT 60.345 191.905 60.655 192.705 ;
        RECT 60.825 192.160 66.170 192.705 ;
        RECT 57.685 191.795 57.855 191.885 ;
        RECT 57.565 191.465 57.855 191.795 ;
        RECT 58.025 191.465 58.365 191.715 ;
        RECT 58.585 191.465 59.260 191.715 ;
        RECT 59.465 191.465 59.800 191.715 ;
        RECT 57.685 191.215 57.855 191.465 ;
        RECT 57.685 191.045 58.625 191.215 ;
        RECT 58.995 191.105 59.260 191.465 ;
        RECT 59.970 191.305 60.140 191.905 ;
        RECT 60.310 191.465 60.645 191.735 ;
        RECT 62.410 191.330 62.750 192.160 ;
        RECT 66.345 191.985 66.685 192.495 ;
        RECT 57.145 190.325 57.605 190.875 ;
        RECT 57.795 190.155 58.125 190.875 ;
        RECT 58.325 190.495 58.625 191.045 ;
        RECT 58.795 190.155 59.075 190.825 ;
        RECT 59.445 190.155 59.705 191.295 ;
        RECT 59.875 190.325 60.205 191.305 ;
        RECT 60.375 190.155 60.655 191.295 ;
        RECT 64.230 190.590 64.580 191.840 ;
        RECT 60.825 190.155 66.170 190.590 ;
        RECT 66.345 190.585 66.605 191.985 ;
        RECT 66.855 191.905 67.125 192.705 ;
        RECT 66.780 191.465 67.110 191.715 ;
        RECT 67.305 191.465 67.585 192.435 ;
        RECT 67.765 191.465 68.065 192.435 ;
        RECT 68.245 191.465 68.595 192.430 ;
        RECT 68.815 192.205 69.310 192.535 ;
        RECT 66.795 191.295 67.110 191.465 ;
        RECT 68.815 191.295 68.985 192.205 ;
        RECT 69.570 192.200 69.905 192.705 ;
        RECT 70.075 192.135 70.315 192.510 ;
        RECT 70.595 192.375 70.765 192.520 ;
        RECT 70.595 192.180 70.970 192.375 ;
        RECT 71.330 192.210 71.725 192.705 ;
        RECT 66.795 191.125 68.985 191.295 ;
        RECT 66.345 190.325 66.685 190.585 ;
        RECT 66.855 190.155 67.185 190.955 ;
        RECT 67.650 190.325 67.900 191.125 ;
        RECT 68.085 190.155 68.415 190.875 ;
        RECT 68.635 190.325 68.885 191.125 ;
        RECT 69.155 190.715 69.395 192.025 ;
        RECT 69.625 191.175 69.925 192.025 ;
        RECT 70.095 191.985 70.315 192.135 ;
        RECT 70.095 191.655 70.630 191.985 ;
        RECT 70.800 191.845 70.970 192.180 ;
        RECT 71.895 192.015 72.135 192.535 ;
        RECT 72.325 192.160 77.670 192.705 ;
        RECT 70.095 191.005 70.330 191.655 ;
        RECT 70.800 191.485 71.785 191.845 ;
        RECT 69.655 190.775 70.330 191.005 ;
        RECT 70.500 191.465 71.785 191.485 ;
        RECT 70.500 191.315 71.360 191.465 ;
        RECT 69.055 190.155 69.390 190.535 ;
        RECT 69.655 190.345 69.825 190.775 ;
        RECT 69.995 190.155 70.325 190.605 ;
        RECT 70.500 190.370 70.785 191.315 ;
        RECT 71.960 191.210 72.135 192.015 ;
        RECT 73.910 191.330 74.250 192.160 ;
        RECT 78.765 191.980 79.055 192.705 ;
        RECT 79.225 191.935 81.815 192.705 ;
        RECT 82.005 192.075 82.335 192.535 ;
        RECT 82.515 192.245 82.685 192.705 ;
        RECT 82.865 192.075 83.195 192.535 ;
        RECT 83.425 192.245 83.595 192.705 ;
        RECT 83.835 192.365 85.025 192.535 ;
        RECT 83.835 192.075 84.165 192.365 ;
        RECT 84.715 192.195 85.025 192.365 ;
        RECT 70.960 190.835 71.655 191.145 ;
        RECT 70.965 190.155 71.650 190.625 ;
        RECT 71.830 190.425 72.135 191.210 ;
        RECT 75.730 190.590 76.080 191.840 ;
        RECT 79.225 191.415 80.435 191.935 ;
        RECT 82.005 191.905 84.165 192.075 ;
        RECT 72.325 190.155 77.670 190.590 ;
        RECT 78.765 190.155 79.055 191.320 ;
        RECT 80.605 191.245 81.815 191.765 ;
        RECT 79.225 190.155 81.815 191.245 ;
        RECT 82.020 191.345 82.350 191.735 ;
        RECT 82.520 191.515 83.320 191.715 ;
        RECT 83.500 191.345 83.995 191.715 ;
        RECT 82.020 191.175 83.995 191.345 ;
        RECT 84.335 191.005 84.545 192.195 ;
        RECT 85.205 192.095 85.545 192.510 ;
        RECT 85.715 192.265 85.885 192.705 ;
        RECT 86.055 192.315 87.305 192.495 ;
        RECT 86.055 192.095 86.385 192.315 ;
        RECT 87.575 192.245 87.745 192.705 ;
        RECT 84.715 191.390 85.030 192.025 ;
        RECT 85.205 191.925 86.385 192.095 ;
        RECT 86.555 192.075 86.920 192.145 ;
        RECT 86.555 191.895 87.805 192.075 ;
        RECT 85.205 191.515 85.670 191.715 ;
        RECT 85.845 191.465 86.175 191.715 ;
        RECT 86.345 191.685 86.810 191.715 ;
        RECT 86.345 191.515 86.815 191.685 ;
        RECT 86.345 191.465 86.810 191.515 ;
        RECT 87.005 191.465 87.360 191.715 ;
        RECT 85.845 191.345 86.025 191.465 ;
        RECT 82.005 190.155 82.335 191.005 ;
        RECT 82.505 190.495 82.725 191.005 ;
        RECT 82.895 190.825 84.545 191.005 ;
        RECT 82.895 190.665 83.195 190.825 ;
        RECT 83.425 190.495 83.615 190.655 ;
        RECT 82.505 190.325 83.615 190.495 ;
        RECT 83.810 190.155 84.140 190.615 ;
        RECT 84.310 190.325 84.545 190.825 ;
        RECT 84.715 190.155 85.025 191.220 ;
        RECT 85.205 190.155 85.525 191.335 ;
        RECT 85.695 191.175 86.025 191.345 ;
        RECT 87.530 191.295 87.805 191.895 ;
        RECT 85.695 190.385 85.895 191.175 ;
        RECT 86.195 191.085 87.805 191.295 ;
        RECT 86.195 190.985 86.605 191.085 ;
        RECT 86.220 190.325 86.605 190.985 ;
        RECT 87.000 190.155 87.785 190.915 ;
        RECT 87.975 190.325 88.255 192.425 ;
        RECT 88.425 191.935 91.015 192.705 ;
        RECT 91.275 192.155 91.445 192.535 ;
        RECT 91.625 192.325 91.955 192.705 ;
        RECT 91.275 191.985 91.940 192.155 ;
        RECT 92.135 192.030 92.395 192.535 ;
        RECT 88.425 191.415 89.635 191.935 ;
        RECT 89.805 191.245 91.015 191.765 ;
        RECT 91.205 191.435 91.535 191.805 ;
        RECT 91.770 191.730 91.940 191.985 ;
        RECT 91.770 191.400 92.055 191.730 ;
        RECT 91.770 191.255 91.940 191.400 ;
        RECT 88.425 190.155 91.015 191.245 ;
        RECT 91.275 191.085 91.940 191.255 ;
        RECT 92.225 191.230 92.395 192.030 ;
        RECT 91.275 190.325 91.445 191.085 ;
        RECT 91.625 190.155 91.955 190.915 ;
        RECT 92.125 190.325 92.395 191.230 ;
        RECT 92.565 192.030 92.825 192.535 ;
        RECT 93.005 192.325 93.335 192.705 ;
        RECT 93.515 192.155 93.685 192.535 ;
        RECT 92.565 191.230 92.735 192.030 ;
        RECT 93.020 191.985 93.685 192.155 ;
        RECT 93.020 191.730 93.190 191.985 ;
        RECT 93.945 191.905 94.255 192.705 ;
        RECT 94.460 191.905 95.155 192.535 ;
        RECT 95.325 192.205 95.585 192.535 ;
        RECT 95.755 192.345 96.085 192.705 ;
        RECT 96.340 192.325 97.640 192.535 ;
        RECT 92.905 191.400 93.190 191.730 ;
        RECT 93.425 191.435 93.755 191.805 ;
        RECT 93.955 191.465 94.290 191.735 ;
        RECT 93.020 191.255 93.190 191.400 ;
        RECT 94.460 191.305 94.630 191.905 ;
        RECT 94.800 191.465 95.135 191.715 ;
        RECT 92.565 190.325 92.835 191.230 ;
        RECT 93.020 191.085 93.685 191.255 ;
        RECT 93.005 190.155 93.335 190.915 ;
        RECT 93.515 190.325 93.685 191.085 ;
        RECT 93.945 190.155 94.225 191.295 ;
        RECT 94.395 190.325 94.725 191.305 ;
        RECT 94.895 190.155 95.155 191.295 ;
        RECT 95.325 191.005 95.495 192.205 ;
        RECT 96.340 192.175 96.510 192.325 ;
        RECT 95.755 192.050 96.510 192.175 ;
        RECT 95.665 192.005 96.510 192.050 ;
        RECT 95.665 191.885 95.935 192.005 ;
        RECT 95.665 191.310 95.835 191.885 ;
        RECT 96.065 191.445 96.475 191.750 ;
        RECT 96.765 191.715 96.975 192.115 ;
        RECT 96.645 191.505 96.975 191.715 ;
        RECT 97.220 191.715 97.440 192.115 ;
        RECT 97.915 191.940 98.370 192.705 ;
        RECT 98.545 191.905 99.240 192.535 ;
        RECT 99.445 191.905 99.755 192.705 ;
        RECT 99.930 192.200 100.265 192.705 ;
        RECT 100.435 192.135 100.675 192.510 ;
        RECT 100.955 192.375 101.125 192.520 ;
        RECT 100.955 192.180 101.330 192.375 ;
        RECT 101.690 192.210 102.085 192.705 ;
        RECT 99.065 191.855 99.240 191.905 ;
        RECT 97.220 191.505 97.695 191.715 ;
        RECT 97.885 191.515 98.375 191.715 ;
        RECT 98.565 191.465 98.900 191.715 ;
        RECT 95.665 191.275 95.865 191.310 ;
        RECT 97.195 191.275 98.370 191.335 ;
        RECT 99.070 191.305 99.240 191.855 ;
        RECT 99.410 191.465 99.745 191.735 ;
        RECT 95.665 191.165 98.370 191.275 ;
        RECT 95.725 191.105 97.525 191.165 ;
        RECT 97.195 191.075 97.525 191.105 ;
        RECT 95.325 190.325 95.585 191.005 ;
        RECT 95.755 190.155 96.005 190.935 ;
        RECT 96.255 190.905 97.090 190.915 ;
        RECT 97.680 190.905 97.865 190.995 ;
        RECT 96.255 190.705 97.865 190.905 ;
        RECT 96.255 190.325 96.505 190.705 ;
        RECT 97.635 190.665 97.865 190.705 ;
        RECT 98.115 190.545 98.370 191.165 ;
        RECT 96.675 190.155 97.030 190.535 ;
        RECT 98.035 190.325 98.370 190.545 ;
        RECT 98.545 190.155 98.805 191.295 ;
        RECT 98.975 190.325 99.305 191.305 ;
        RECT 99.475 190.155 99.755 191.295 ;
        RECT 99.985 191.175 100.285 192.025 ;
        RECT 100.455 191.985 100.675 192.135 ;
        RECT 100.455 191.655 100.990 191.985 ;
        RECT 101.160 191.845 101.330 192.180 ;
        RECT 102.255 192.015 102.495 192.535 ;
        RECT 100.455 191.005 100.690 191.655 ;
        RECT 101.160 191.485 102.145 191.845 ;
        RECT 100.015 190.775 100.690 191.005 ;
        RECT 100.860 191.465 102.145 191.485 ;
        RECT 100.860 191.315 101.720 191.465 ;
        RECT 100.015 190.345 100.185 190.775 ;
        RECT 100.355 190.155 100.685 190.605 ;
        RECT 100.860 190.370 101.145 191.315 ;
        RECT 102.320 191.210 102.495 192.015 ;
        RECT 102.695 191.975 102.995 192.705 ;
        RECT 103.175 191.795 103.405 192.415 ;
        RECT 103.605 192.145 103.830 192.525 ;
        RECT 104.000 192.315 104.330 192.705 ;
        RECT 103.605 191.965 103.935 192.145 ;
        RECT 102.700 191.465 102.995 191.795 ;
        RECT 103.175 191.465 103.590 191.795 ;
        RECT 103.760 191.295 103.935 191.965 ;
        RECT 104.105 191.465 104.345 192.115 ;
        RECT 104.525 191.980 104.815 192.705 ;
        RECT 105.045 191.885 105.255 192.705 ;
        RECT 105.425 191.905 105.755 192.535 ;
        RECT 101.320 190.835 102.015 191.145 ;
        RECT 101.325 190.155 102.010 190.625 ;
        RECT 102.190 190.425 102.495 191.210 ;
        RECT 102.695 190.935 103.590 191.265 ;
        RECT 103.760 191.105 104.345 191.295 ;
        RECT 102.695 190.765 103.900 190.935 ;
        RECT 102.695 190.335 103.025 190.765 ;
        RECT 103.205 190.155 103.400 190.595 ;
        RECT 103.570 190.335 103.900 190.765 ;
        RECT 104.070 190.335 104.345 191.105 ;
        RECT 104.525 190.155 104.815 191.320 ;
        RECT 105.425 191.305 105.675 191.905 ;
        RECT 105.925 191.885 106.155 192.705 ;
        RECT 106.455 192.225 106.755 192.705 ;
        RECT 106.925 192.055 107.185 192.510 ;
        RECT 107.355 192.225 107.615 192.705 ;
        RECT 107.795 192.055 108.055 192.510 ;
        RECT 108.225 192.225 108.475 192.705 ;
        RECT 108.655 192.055 108.915 192.510 ;
        RECT 109.085 192.225 109.335 192.705 ;
        RECT 109.515 192.055 109.775 192.510 ;
        RECT 109.945 192.225 110.190 192.705 ;
        RECT 110.360 192.055 110.635 192.510 ;
        RECT 110.805 192.225 111.050 192.705 ;
        RECT 111.220 192.055 111.480 192.510 ;
        RECT 111.650 192.225 111.910 192.705 ;
        RECT 112.080 192.055 112.340 192.510 ;
        RECT 112.510 192.225 112.770 192.705 ;
        RECT 112.940 192.055 113.200 192.510 ;
        RECT 113.370 192.145 113.630 192.705 ;
        RECT 106.455 191.885 113.200 192.055 ;
        RECT 105.845 191.465 106.175 191.715 ;
        RECT 105.045 190.155 105.255 191.295 ;
        RECT 105.425 190.325 105.755 191.305 ;
        RECT 106.455 191.295 107.620 191.885 ;
        RECT 113.800 191.715 114.050 192.525 ;
        RECT 114.230 192.180 114.490 192.705 ;
        RECT 114.660 191.715 114.910 192.525 ;
        RECT 115.090 192.195 115.395 192.705 ;
        RECT 115.655 192.225 115.955 192.705 ;
        RECT 116.125 192.055 116.385 192.510 ;
        RECT 116.555 192.225 116.815 192.705 ;
        RECT 116.995 192.055 117.255 192.510 ;
        RECT 117.425 192.225 117.675 192.705 ;
        RECT 117.855 192.055 118.115 192.510 ;
        RECT 118.285 192.225 118.535 192.705 ;
        RECT 118.715 192.055 118.975 192.510 ;
        RECT 119.145 192.225 119.390 192.705 ;
        RECT 119.560 192.055 119.835 192.510 ;
        RECT 120.005 192.225 120.250 192.705 ;
        RECT 120.420 192.055 120.680 192.510 ;
        RECT 120.850 192.225 121.110 192.705 ;
        RECT 121.280 192.055 121.540 192.510 ;
        RECT 121.710 192.225 121.970 192.705 ;
        RECT 122.140 192.055 122.400 192.510 ;
        RECT 122.570 192.145 122.830 192.705 ;
        RECT 115.655 192.025 122.400 192.055 ;
        RECT 107.790 191.465 114.910 191.715 ;
        RECT 115.080 191.465 115.395 192.025 ;
        RECT 115.625 191.885 122.400 192.025 ;
        RECT 115.625 191.855 116.820 191.885 ;
        RECT 105.925 190.155 106.155 191.295 ;
        RECT 106.455 191.070 113.200 191.295 ;
        RECT 106.455 190.155 106.725 190.900 ;
        RECT 106.895 190.330 107.185 191.070 ;
        RECT 107.795 191.055 113.200 191.070 ;
        RECT 107.355 190.160 107.610 190.885 ;
        RECT 107.795 190.330 108.055 191.055 ;
        RECT 108.225 190.160 108.470 190.885 ;
        RECT 108.655 190.330 108.915 191.055 ;
        RECT 109.085 190.160 109.330 190.885 ;
        RECT 109.515 190.330 109.775 191.055 ;
        RECT 109.945 190.160 110.190 190.885 ;
        RECT 110.360 190.330 110.620 191.055 ;
        RECT 110.790 190.160 111.050 190.885 ;
        RECT 111.220 190.330 111.480 191.055 ;
        RECT 111.650 190.160 111.910 190.885 ;
        RECT 112.080 190.330 112.340 191.055 ;
        RECT 112.510 190.160 112.770 190.885 ;
        RECT 112.940 190.330 113.200 191.055 ;
        RECT 113.370 190.160 113.630 190.955 ;
        RECT 113.800 190.330 114.050 191.465 ;
        RECT 107.355 190.155 113.630 190.160 ;
        RECT 114.230 190.155 114.490 190.965 ;
        RECT 114.665 190.325 114.910 191.465 ;
        RECT 115.655 191.295 116.820 191.855 ;
        RECT 123.000 191.715 123.250 192.525 ;
        RECT 123.430 192.180 123.690 192.705 ;
        RECT 123.860 191.715 124.110 192.525 ;
        RECT 124.290 192.195 124.595 192.705 ;
        RECT 116.990 191.465 124.110 191.715 ;
        RECT 124.280 191.465 124.595 192.025 ;
        RECT 124.765 191.905 125.060 192.705 ;
        RECT 125.230 191.795 125.505 192.535 ;
        RECT 125.675 191.965 126.345 192.705 ;
        RECT 126.515 192.135 126.800 192.480 ;
        RECT 126.980 192.305 127.355 192.705 ;
        RECT 127.570 192.135 127.900 192.480 ;
        RECT 126.515 191.965 127.900 192.135 ;
        RECT 128.150 191.965 128.735 192.535 ;
        RECT 125.230 191.735 125.585 191.795 ;
        RECT 124.765 191.475 125.585 191.735 ;
        RECT 115.655 191.070 122.400 191.295 ;
        RECT 115.090 190.155 115.385 190.965 ;
        RECT 115.655 190.155 115.925 190.900 ;
        RECT 116.095 190.330 116.385 191.070 ;
        RECT 116.995 191.055 122.400 191.070 ;
        RECT 116.555 190.160 116.810 190.885 ;
        RECT 116.995 190.330 117.255 191.055 ;
        RECT 117.425 190.160 117.670 190.885 ;
        RECT 117.855 190.330 118.115 191.055 ;
        RECT 118.285 190.160 118.530 190.885 ;
        RECT 118.715 190.330 118.975 191.055 ;
        RECT 119.145 190.160 119.390 190.885 ;
        RECT 119.560 190.330 119.820 191.055 ;
        RECT 119.990 190.160 120.250 190.885 ;
        RECT 120.420 190.330 120.680 191.055 ;
        RECT 120.850 190.160 121.110 190.885 ;
        RECT 121.280 190.330 121.540 191.055 ;
        RECT 121.710 190.160 121.970 190.885 ;
        RECT 122.140 190.330 122.400 191.055 ;
        RECT 122.570 190.160 122.830 190.955 ;
        RECT 123.000 190.330 123.250 191.465 ;
        RECT 116.555 190.155 122.830 190.160 ;
        RECT 123.430 190.155 123.690 190.965 ;
        RECT 123.865 190.325 124.110 191.465 ;
        RECT 124.290 190.155 124.585 190.965 ;
        RECT 124.765 190.155 125.060 191.305 ;
        RECT 125.230 190.325 125.585 191.475 ;
        RECT 125.755 191.295 125.925 191.795 ;
        RECT 126.095 191.465 126.430 191.795 ;
        RECT 126.600 191.465 126.930 191.795 ;
        RECT 125.755 191.125 126.490 191.295 ;
        RECT 125.755 190.155 126.150 190.955 ;
        RECT 126.320 190.495 126.490 191.125 ;
        RECT 126.660 190.720 126.930 191.465 ;
        RECT 127.120 191.465 127.410 191.795 ;
        RECT 127.580 191.465 127.980 191.795 ;
        RECT 127.120 190.720 127.355 191.465 ;
        RECT 128.150 191.295 128.320 191.965 ;
        RECT 128.905 191.905 129.600 192.535 ;
        RECT 129.805 191.905 130.115 192.705 ;
        RECT 130.285 191.980 130.575 192.705 ;
        RECT 130.755 192.365 131.090 192.535 ;
        RECT 130.755 191.965 131.370 192.365 ;
        RECT 132.050 192.325 132.385 192.705 ;
        RECT 132.975 192.265 133.210 192.705 ;
        RECT 133.380 192.175 133.710 192.535 ;
        RECT 133.880 192.345 134.210 192.705 ;
        RECT 131.540 191.965 132.810 192.155 ;
        RECT 133.380 192.005 134.200 192.175 ;
        RECT 129.425 191.855 129.600 191.905 ;
        RECT 128.490 191.465 128.735 191.795 ;
        RECT 128.925 191.465 129.260 191.715 ;
        RECT 129.430 191.305 129.600 191.855 ;
        RECT 129.770 191.465 130.105 191.735 ;
        RECT 130.745 191.465 131.020 191.795 ;
        RECT 127.525 191.125 128.735 191.295 ;
        RECT 127.525 190.495 127.855 191.125 ;
        RECT 126.320 190.325 127.855 190.495 ;
        RECT 128.040 190.155 128.275 190.955 ;
        RECT 128.445 190.325 128.735 191.125 ;
        RECT 128.905 190.155 129.165 191.295 ;
        RECT 129.335 190.325 129.665 191.305 ;
        RECT 129.835 190.155 130.115 191.295 ;
        RECT 130.285 190.155 130.575 191.320 ;
        RECT 131.190 191.280 131.370 191.965 ;
        RECT 131.540 191.465 131.900 191.795 ;
        RECT 132.190 191.685 132.480 191.795 ;
        RECT 132.185 191.515 132.480 191.685 ;
        RECT 132.190 191.465 132.480 191.515 ;
        RECT 132.650 191.465 132.985 191.795 ;
        RECT 133.155 191.465 133.835 191.795 ;
        RECT 133.155 191.280 133.325 191.465 ;
        RECT 130.750 191.025 133.325 191.280 ;
        RECT 130.750 190.325 131.015 191.025 ;
        RECT 131.185 190.155 131.515 190.855 ;
        RECT 131.685 190.325 132.355 191.025 ;
        RECT 134.005 190.885 134.200 192.005 ;
        RECT 134.445 191.125 134.675 192.465 ;
        RECT 134.855 191.625 135.085 192.525 ;
        RECT 135.285 191.925 135.530 192.705 ;
        RECT 135.700 192.165 136.130 192.525 ;
        RECT 136.710 192.335 137.440 192.705 ;
        RECT 135.700 191.975 137.440 192.165 ;
        RECT 135.700 191.745 135.920 191.975 ;
        RECT 134.855 190.945 135.195 191.625 ;
        RECT 132.860 190.155 133.290 190.855 ;
        RECT 133.470 190.715 134.200 190.885 ;
        RECT 134.445 190.745 135.195 190.945 ;
        RECT 135.375 191.445 135.920 191.745 ;
        RECT 133.470 190.325 133.660 190.715 ;
        RECT 133.830 190.155 134.160 190.535 ;
        RECT 134.445 190.355 134.685 190.745 ;
        RECT 134.855 190.155 135.205 190.565 ;
        RECT 135.375 190.335 135.705 191.445 ;
        RECT 136.090 191.175 136.515 191.795 ;
        RECT 136.710 191.175 136.970 191.795 ;
        RECT 137.180 191.465 137.440 191.975 ;
        RECT 135.875 190.805 136.900 191.005 ;
        RECT 135.875 190.335 136.055 190.805 ;
        RECT 136.225 190.155 136.555 190.635 ;
        RECT 136.730 190.335 136.900 190.805 ;
        RECT 137.165 190.155 137.450 191.295 ;
        RECT 137.640 190.335 137.920 192.525 ;
        RECT 138.565 191.955 139.775 192.705 ;
        RECT 138.565 191.245 139.085 191.785 ;
        RECT 139.255 191.415 139.775 191.955 ;
        RECT 138.565 190.155 139.775 191.245 ;
        RECT 27.160 189.985 139.860 190.155 ;
        RECT 27.245 188.895 28.455 189.985 ;
        RECT 28.625 188.895 31.215 189.985 ;
        RECT 27.245 188.185 27.765 188.725 ;
        RECT 27.935 188.355 28.455 188.895 ;
        RECT 28.625 188.205 29.835 188.725 ;
        RECT 30.005 188.375 31.215 188.895 ;
        RECT 31.425 188.845 31.655 189.985 ;
        RECT 31.825 188.835 32.155 189.815 ;
        RECT 32.325 188.845 32.535 189.985 ;
        RECT 32.765 188.895 36.275 189.985 ;
        RECT 31.405 188.425 31.735 188.675 ;
        RECT 27.245 187.435 28.455 188.185 ;
        RECT 28.625 187.435 31.215 188.205 ;
        RECT 31.425 187.435 31.655 188.255 ;
        RECT 31.905 188.235 32.155 188.835 ;
        RECT 31.825 187.605 32.155 188.235 ;
        RECT 32.325 187.435 32.535 188.255 ;
        RECT 32.765 188.205 34.415 188.725 ;
        RECT 34.585 188.375 36.275 188.895 ;
        RECT 36.450 188.845 36.770 189.985 ;
        RECT 36.950 188.675 37.145 189.725 ;
        RECT 37.325 189.135 37.655 189.815 ;
        RECT 37.855 189.185 38.110 189.985 ;
        RECT 37.325 188.855 37.675 189.135 ;
        RECT 36.510 188.625 36.770 188.675 ;
        RECT 36.505 188.455 36.770 188.625 ;
        RECT 36.510 188.345 36.770 188.455 ;
        RECT 36.950 188.345 37.335 188.675 ;
        RECT 37.505 188.475 37.675 188.855 ;
        RECT 37.865 188.645 38.110 189.005 ;
        RECT 38.290 188.845 38.610 189.985 ;
        RECT 38.790 188.675 38.985 189.725 ;
        RECT 39.165 189.135 39.495 189.815 ;
        RECT 39.695 189.185 39.950 189.985 ;
        RECT 39.165 188.855 39.515 189.135 ;
        RECT 38.350 188.625 38.610 188.675 ;
        RECT 37.505 188.305 38.025 188.475 ;
        RECT 38.345 188.455 38.610 188.625 ;
        RECT 38.350 188.345 38.610 188.455 ;
        RECT 38.790 188.345 39.175 188.675 ;
        RECT 39.345 188.475 39.515 188.855 ;
        RECT 39.705 188.645 39.950 189.005 ;
        RECT 40.125 188.820 40.415 189.985 ;
        RECT 40.585 189.475 40.845 189.985 ;
        RECT 39.345 188.305 39.865 188.475 ;
        RECT 40.585 188.425 40.925 189.305 ;
        RECT 41.095 188.595 41.265 189.815 ;
        RECT 41.505 189.480 42.120 189.985 ;
        RECT 41.505 188.945 41.755 189.310 ;
        RECT 41.925 189.305 42.120 189.480 ;
        RECT 42.290 189.475 42.765 189.815 ;
        RECT 42.935 189.440 43.150 189.985 ;
        RECT 41.925 189.115 42.255 189.305 ;
        RECT 42.475 188.945 43.190 189.240 ;
        RECT 43.360 189.115 43.635 189.815 ;
        RECT 43.805 189.550 49.150 189.985 ;
        RECT 41.505 188.775 43.295 188.945 ;
        RECT 32.765 187.435 36.275 188.205 ;
        RECT 36.450 187.965 37.665 188.135 ;
        RECT 36.450 187.615 36.740 187.965 ;
        RECT 36.935 187.435 37.265 187.795 ;
        RECT 37.435 187.660 37.665 187.965 ;
        RECT 37.855 187.740 38.025 188.305 ;
        RECT 38.290 187.965 39.505 188.135 ;
        RECT 38.290 187.615 38.580 187.965 ;
        RECT 38.775 187.435 39.105 187.795 ;
        RECT 39.275 187.660 39.505 187.965 ;
        RECT 39.695 187.945 39.865 188.305 ;
        RECT 41.095 188.345 41.890 188.595 ;
        RECT 41.095 188.255 41.345 188.345 ;
        RECT 39.695 187.775 39.895 187.945 ;
        RECT 39.695 187.740 39.865 187.775 ;
        RECT 40.125 187.435 40.415 188.160 ;
        RECT 40.585 187.435 40.845 188.255 ;
        RECT 41.015 187.835 41.345 188.255 ;
        RECT 42.060 187.920 42.315 188.775 ;
        RECT 41.525 187.655 42.315 187.920 ;
        RECT 42.485 188.075 42.895 188.595 ;
        RECT 43.065 188.345 43.295 188.775 ;
        RECT 43.465 188.085 43.635 189.115 ;
        RECT 42.485 187.655 42.685 188.075 ;
        RECT 42.875 187.435 43.205 187.895 ;
        RECT 43.375 187.605 43.635 188.085 ;
        RECT 45.390 187.980 45.730 188.810 ;
        RECT 47.210 188.300 47.560 189.550 ;
        RECT 49.325 188.895 50.995 189.985 ;
        RECT 49.325 188.205 50.075 188.725 ;
        RECT 50.245 188.375 50.995 188.895 ;
        RECT 51.690 189.015 51.960 189.810 ;
        RECT 52.140 189.185 52.355 189.985 ;
        RECT 52.535 189.015 52.820 189.810 ;
        RECT 51.690 188.845 52.820 189.015 ;
        RECT 51.670 188.375 52.170 188.640 ;
        RECT 52.390 188.345 52.775 188.675 ;
        RECT 53.000 188.345 53.280 189.815 ;
        RECT 53.460 188.400 53.790 189.815 ;
        RECT 53.960 188.640 54.165 189.815 ;
        RECT 54.335 188.995 54.545 189.810 ;
        RECT 54.785 189.165 55.115 189.985 ;
        RECT 54.335 188.815 54.985 188.995 ;
        RECT 55.290 188.970 55.545 189.810 ;
        RECT 53.960 188.400 54.390 188.640 ;
        RECT 43.805 187.435 49.150 187.980 ;
        RECT 49.325 187.435 50.995 188.205 ;
        RECT 52.390 188.195 52.695 188.345 ;
        RECT 51.725 187.435 51.965 188.110 ;
        RECT 52.140 187.635 52.695 188.195 ;
        RECT 54.765 188.175 54.985 188.815 ;
        RECT 52.875 188.005 54.985 188.175 ;
        RECT 52.875 187.610 53.080 188.005 ;
        RECT 53.765 188.000 54.985 188.005 ;
        RECT 53.250 187.435 53.595 187.835 ;
        RECT 53.765 187.610 54.095 188.000 ;
        RECT 54.370 187.435 55.045 187.820 ;
        RECT 55.215 187.605 55.545 188.970 ;
        RECT 55.765 188.845 56.025 189.985 ;
        RECT 56.195 188.835 56.525 189.815 ;
        RECT 56.695 188.845 56.975 189.985 ;
        RECT 57.155 189.015 57.485 189.800 ;
        RECT 57.155 188.845 57.835 189.015 ;
        RECT 58.015 188.845 58.345 189.985 ;
        RECT 58.525 188.895 62.035 189.985 ;
        RECT 55.785 188.425 56.120 188.675 ;
        RECT 56.290 188.235 56.460 188.835 ;
        RECT 56.630 188.405 56.965 188.675 ;
        RECT 57.145 188.425 57.495 188.675 ;
        RECT 57.665 188.245 57.835 188.845 ;
        RECT 58.005 188.425 58.355 188.675 ;
        RECT 55.765 187.605 56.460 188.235 ;
        RECT 56.665 187.435 56.975 188.235 ;
        RECT 57.165 187.435 57.405 188.245 ;
        RECT 57.575 187.605 57.905 188.245 ;
        RECT 58.075 187.435 58.345 188.245 ;
        RECT 58.525 188.205 60.175 188.725 ;
        RECT 60.345 188.375 62.035 188.895 ;
        RECT 63.165 188.845 63.395 189.985 ;
        RECT 63.565 188.835 63.895 189.815 ;
        RECT 64.065 188.845 64.275 189.985 ;
        RECT 64.505 188.895 65.715 189.985 ;
        RECT 63.145 188.425 63.475 188.675 ;
        RECT 58.525 187.435 62.035 188.205 ;
        RECT 63.165 187.435 63.395 188.255 ;
        RECT 63.645 188.235 63.895 188.835 ;
        RECT 63.565 187.605 63.895 188.235 ;
        RECT 64.065 187.435 64.275 188.255 ;
        RECT 64.505 188.185 65.025 188.725 ;
        RECT 65.195 188.355 65.715 188.895 ;
        RECT 65.885 188.820 66.175 189.985 ;
        RECT 66.895 189.365 67.065 189.795 ;
        RECT 67.235 189.535 67.565 189.985 ;
        RECT 66.895 189.135 67.570 189.365 ;
        RECT 64.505 187.435 65.715 188.185 ;
        RECT 65.885 187.435 66.175 188.160 ;
        RECT 66.865 188.115 67.165 188.965 ;
        RECT 67.335 188.485 67.570 189.135 ;
        RECT 67.740 188.825 68.025 189.770 ;
        RECT 68.205 189.515 68.890 189.985 ;
        RECT 68.200 188.995 68.895 189.305 ;
        RECT 69.070 188.930 69.375 189.715 ;
        RECT 67.740 188.675 68.600 188.825 ;
        RECT 69.165 188.795 69.375 188.930 ;
        RECT 69.585 189.095 69.845 189.805 ;
        RECT 70.015 189.275 70.345 189.985 ;
        RECT 70.515 189.095 70.745 189.805 ;
        RECT 69.585 188.855 70.745 189.095 ;
        RECT 70.925 189.075 71.195 189.805 ;
        RECT 71.375 189.255 71.715 189.985 ;
        RECT 70.925 188.855 71.695 189.075 ;
        RECT 67.740 188.655 69.025 188.675 ;
        RECT 67.335 188.155 67.870 188.485 ;
        RECT 68.040 188.295 69.025 188.655 ;
        RECT 67.335 188.005 67.555 188.155 ;
        RECT 66.810 187.435 67.145 187.940 ;
        RECT 67.315 187.630 67.555 188.005 ;
        RECT 68.040 187.960 68.210 188.295 ;
        RECT 69.200 188.125 69.375 188.795 ;
        RECT 69.575 188.345 69.875 188.675 ;
        RECT 70.055 188.365 70.580 188.675 ;
        RECT 70.760 188.365 71.225 188.675 ;
        RECT 67.835 187.765 68.210 187.960 ;
        RECT 67.835 187.620 68.005 187.765 ;
        RECT 68.570 187.435 68.965 187.930 ;
        RECT 69.135 187.605 69.375 188.125 ;
        RECT 69.585 187.435 69.875 188.165 ;
        RECT 70.055 187.725 70.285 188.365 ;
        RECT 71.405 188.185 71.695 188.855 ;
        RECT 70.465 187.985 71.695 188.185 ;
        RECT 70.465 187.615 70.775 187.985 ;
        RECT 70.955 187.435 71.625 187.805 ;
        RECT 71.885 187.615 72.145 189.805 ;
        RECT 72.325 188.845 72.600 189.815 ;
        RECT 72.810 189.185 73.090 189.985 ;
        RECT 73.260 189.475 74.875 189.805 ;
        RECT 73.260 189.135 74.435 189.305 ;
        RECT 73.260 189.015 73.430 189.135 ;
        RECT 72.770 188.845 73.430 189.015 ;
        RECT 72.325 188.110 72.495 188.845 ;
        RECT 72.770 188.675 72.940 188.845 ;
        RECT 73.690 188.675 73.935 188.965 ;
        RECT 74.105 188.845 74.435 189.135 ;
        RECT 74.695 188.675 74.865 189.235 ;
        RECT 75.115 188.845 75.375 189.985 ;
        RECT 75.545 189.550 80.890 189.985 ;
        RECT 72.665 188.345 72.940 188.675 ;
        RECT 73.110 188.345 73.935 188.675 ;
        RECT 74.150 188.345 74.865 188.675 ;
        RECT 75.035 188.425 75.370 188.675 ;
        RECT 72.770 188.175 72.940 188.345 ;
        RECT 74.615 188.255 74.865 188.345 ;
        RECT 72.325 187.765 72.600 188.110 ;
        RECT 72.770 188.005 74.435 188.175 ;
        RECT 72.790 187.435 73.165 187.835 ;
        RECT 73.335 187.655 73.505 188.005 ;
        RECT 73.675 187.435 74.005 187.835 ;
        RECT 74.175 187.605 74.435 188.005 ;
        RECT 74.615 187.835 74.945 188.255 ;
        RECT 75.115 187.435 75.375 188.255 ;
        RECT 77.130 187.980 77.470 188.810 ;
        RECT 78.950 188.300 79.300 189.550 ;
        RECT 81.065 188.895 84.575 189.985 ;
        RECT 84.745 188.895 85.955 189.985 ;
        RECT 81.065 188.205 82.715 188.725 ;
        RECT 82.885 188.375 84.575 188.895 ;
        RECT 75.545 187.435 80.890 187.980 ;
        RECT 81.065 187.435 84.575 188.205 ;
        RECT 84.745 188.185 85.265 188.725 ;
        RECT 85.435 188.355 85.955 188.895 ;
        RECT 86.135 189.035 86.410 189.805 ;
        RECT 86.580 189.375 86.910 189.805 ;
        RECT 87.080 189.545 87.275 189.985 ;
        RECT 87.455 189.375 87.785 189.805 ;
        RECT 86.580 189.205 87.785 189.375 ;
        RECT 86.135 188.845 86.720 189.035 ;
        RECT 86.890 188.875 87.785 189.205 ;
        RECT 88.885 188.845 89.145 189.985 ;
        RECT 84.745 187.435 85.955 188.185 ;
        RECT 86.135 188.025 86.375 188.675 ;
        RECT 86.545 188.175 86.720 188.845 ;
        RECT 89.315 188.835 89.645 189.815 ;
        RECT 89.815 188.845 90.095 189.985 ;
        RECT 90.265 188.845 90.545 189.985 ;
        RECT 90.715 188.835 91.045 189.815 ;
        RECT 91.215 188.845 91.475 189.985 ;
        RECT 86.890 188.345 87.305 188.675 ;
        RECT 87.485 188.345 87.780 188.675 ;
        RECT 88.905 188.425 89.240 188.675 ;
        RECT 86.545 187.995 86.875 188.175 ;
        RECT 86.150 187.435 86.480 187.825 ;
        RECT 86.650 187.615 86.875 187.995 ;
        RECT 87.075 187.725 87.305 188.345 ;
        RECT 89.410 188.235 89.580 188.835 ;
        RECT 89.750 188.405 90.085 188.675 ;
        RECT 90.275 188.405 90.610 188.675 ;
        RECT 90.780 188.235 90.950 188.835 ;
        RECT 91.645 188.820 91.935 189.985 ;
        RECT 92.105 189.135 92.365 189.815 ;
        RECT 92.535 189.205 92.785 189.985 ;
        RECT 93.035 189.435 93.285 189.815 ;
        RECT 93.455 189.605 93.810 189.985 ;
        RECT 94.815 189.595 95.150 189.815 ;
        RECT 94.415 189.435 94.645 189.475 ;
        RECT 93.035 189.235 94.645 189.435 ;
        RECT 93.035 189.225 93.870 189.235 ;
        RECT 94.460 189.145 94.645 189.235 ;
        RECT 91.120 188.425 91.455 188.675 ;
        RECT 87.485 187.435 87.785 188.165 ;
        RECT 88.885 187.605 89.580 188.235 ;
        RECT 89.785 187.435 90.095 188.235 ;
        RECT 90.265 187.435 90.575 188.235 ;
        RECT 90.780 187.605 91.475 188.235 ;
        RECT 91.645 187.435 91.935 188.160 ;
        RECT 92.105 187.945 92.275 189.135 ;
        RECT 93.975 189.035 94.305 189.065 ;
        RECT 92.505 188.975 94.305 189.035 ;
        RECT 94.895 188.975 95.150 189.595 ;
        RECT 92.445 188.865 95.150 188.975 ;
        RECT 92.445 188.830 92.645 188.865 ;
        RECT 92.445 188.255 92.615 188.830 ;
        RECT 93.975 188.805 95.150 188.865 ;
        RECT 95.795 189.015 96.125 189.800 ;
        RECT 95.795 188.845 96.475 189.015 ;
        RECT 96.655 188.845 96.985 189.985 ;
        RECT 97.255 189.240 97.525 189.985 ;
        RECT 98.155 189.980 104.430 189.985 ;
        RECT 97.695 189.070 97.985 189.810 ;
        RECT 98.155 189.255 98.410 189.980 ;
        RECT 98.595 189.085 98.855 189.810 ;
        RECT 99.025 189.255 99.270 189.980 ;
        RECT 99.455 189.085 99.715 189.810 ;
        RECT 99.885 189.255 100.130 189.980 ;
        RECT 100.315 189.085 100.575 189.810 ;
        RECT 100.745 189.255 100.990 189.980 ;
        RECT 101.160 189.085 101.420 189.810 ;
        RECT 101.590 189.255 101.850 189.980 ;
        RECT 102.020 189.085 102.280 189.810 ;
        RECT 102.450 189.255 102.710 189.980 ;
        RECT 102.880 189.085 103.140 189.810 ;
        RECT 103.310 189.255 103.570 189.980 ;
        RECT 103.740 189.085 104.000 189.810 ;
        RECT 104.170 189.185 104.430 189.980 ;
        RECT 98.595 189.070 104.000 189.085 ;
        RECT 97.255 188.845 104.000 189.070 ;
        RECT 92.845 188.390 93.255 188.695 ;
        RECT 93.425 188.425 93.755 188.635 ;
        RECT 92.445 188.135 92.715 188.255 ;
        RECT 92.445 188.090 93.290 188.135 ;
        RECT 92.535 187.965 93.290 188.090 ;
        RECT 93.545 188.025 93.755 188.425 ;
        RECT 94.000 188.425 94.475 188.635 ;
        RECT 94.665 188.425 95.155 188.625 ;
        RECT 95.785 188.425 96.135 188.675 ;
        RECT 94.000 188.025 94.220 188.425 ;
        RECT 96.305 188.245 96.475 188.845 ;
        RECT 96.645 188.425 96.995 188.675 ;
        RECT 97.255 188.255 98.420 188.845 ;
        RECT 104.600 188.675 104.850 189.810 ;
        RECT 105.030 189.175 105.290 189.985 ;
        RECT 105.465 188.675 105.710 189.815 ;
        RECT 105.890 189.175 106.185 189.985 ;
        RECT 106.370 188.845 106.690 189.985 ;
        RECT 106.870 188.675 107.065 189.725 ;
        RECT 107.245 189.135 107.575 189.815 ;
        RECT 107.775 189.185 108.030 189.985 ;
        RECT 108.295 189.240 108.565 189.985 ;
        RECT 109.195 189.980 115.470 189.985 ;
        RECT 107.245 188.855 107.595 189.135 ;
        RECT 108.735 189.070 109.025 189.810 ;
        RECT 109.195 189.255 109.450 189.980 ;
        RECT 109.635 189.085 109.895 189.810 ;
        RECT 110.065 189.255 110.310 189.980 ;
        RECT 110.495 189.085 110.755 189.810 ;
        RECT 110.925 189.255 111.170 189.980 ;
        RECT 111.355 189.085 111.615 189.810 ;
        RECT 111.785 189.255 112.030 189.980 ;
        RECT 112.200 189.085 112.460 189.810 ;
        RECT 112.630 189.255 112.890 189.980 ;
        RECT 113.060 189.085 113.320 189.810 ;
        RECT 113.490 189.255 113.750 189.980 ;
        RECT 113.920 189.085 114.180 189.810 ;
        RECT 114.350 189.255 114.610 189.980 ;
        RECT 114.780 189.085 115.040 189.810 ;
        RECT 115.210 189.185 115.470 189.980 ;
        RECT 109.635 189.070 115.040 189.085 ;
        RECT 98.590 188.425 105.710 188.675 ;
        RECT 92.105 187.935 92.335 187.945 ;
        RECT 92.105 187.605 92.365 187.935 ;
        RECT 93.120 187.815 93.290 187.965 ;
        RECT 92.535 187.435 92.865 187.795 ;
        RECT 93.120 187.605 94.420 187.815 ;
        RECT 94.695 187.435 95.150 188.200 ;
        RECT 95.805 187.435 96.045 188.245 ;
        RECT 96.215 187.605 96.545 188.245 ;
        RECT 96.715 187.435 96.985 188.245 ;
        RECT 97.255 188.085 104.000 188.255 ;
        RECT 97.255 187.435 97.555 187.915 ;
        RECT 97.725 187.630 97.985 188.085 ;
        RECT 98.155 187.435 98.415 187.915 ;
        RECT 98.595 187.630 98.855 188.085 ;
        RECT 99.025 187.435 99.275 187.915 ;
        RECT 99.455 187.630 99.715 188.085 ;
        RECT 99.885 187.435 100.135 187.915 ;
        RECT 100.315 187.630 100.575 188.085 ;
        RECT 100.745 187.435 100.990 187.915 ;
        RECT 101.160 187.630 101.435 188.085 ;
        RECT 101.605 187.435 101.850 187.915 ;
        RECT 102.020 187.630 102.280 188.085 ;
        RECT 102.450 187.435 102.710 187.915 ;
        RECT 102.880 187.630 103.140 188.085 ;
        RECT 103.310 187.435 103.570 187.915 ;
        RECT 103.740 187.630 104.000 188.085 ;
        RECT 104.170 187.435 104.430 187.995 ;
        RECT 104.600 187.615 104.850 188.425 ;
        RECT 105.030 187.435 105.290 187.960 ;
        RECT 105.460 187.615 105.710 188.425 ;
        RECT 105.880 188.115 106.195 188.675 ;
        RECT 106.430 188.625 106.690 188.675 ;
        RECT 106.425 188.455 106.690 188.625 ;
        RECT 106.430 188.345 106.690 188.455 ;
        RECT 106.870 188.345 107.255 188.675 ;
        RECT 107.425 188.475 107.595 188.855 ;
        RECT 107.785 188.645 108.030 189.005 ;
        RECT 108.295 188.845 115.040 189.070 ;
        RECT 107.425 188.305 107.945 188.475 ;
        RECT 106.370 187.965 107.585 188.135 ;
        RECT 105.890 187.435 106.195 187.945 ;
        RECT 106.370 187.615 106.660 187.965 ;
        RECT 106.855 187.435 107.185 187.795 ;
        RECT 107.355 187.660 107.585 187.965 ;
        RECT 107.775 187.945 107.945 188.305 ;
        RECT 108.295 188.255 109.460 188.845 ;
        RECT 115.640 188.675 115.890 189.810 ;
        RECT 116.070 189.175 116.330 189.985 ;
        RECT 116.505 188.675 116.750 189.815 ;
        RECT 116.930 189.175 117.225 189.985 ;
        RECT 117.405 188.820 117.695 189.985 ;
        RECT 117.955 189.240 118.225 189.985 ;
        RECT 118.855 189.980 125.130 189.985 ;
        RECT 118.395 189.070 118.685 189.810 ;
        RECT 118.855 189.255 119.110 189.980 ;
        RECT 119.295 189.085 119.555 189.810 ;
        RECT 119.725 189.255 119.970 189.980 ;
        RECT 120.155 189.085 120.415 189.810 ;
        RECT 120.585 189.255 120.830 189.980 ;
        RECT 121.015 189.085 121.275 189.810 ;
        RECT 121.445 189.255 121.690 189.980 ;
        RECT 121.860 189.085 122.120 189.810 ;
        RECT 122.290 189.255 122.550 189.980 ;
        RECT 122.720 189.085 122.980 189.810 ;
        RECT 123.150 189.255 123.410 189.980 ;
        RECT 123.580 189.085 123.840 189.810 ;
        RECT 124.010 189.255 124.270 189.980 ;
        RECT 124.440 189.085 124.700 189.810 ;
        RECT 124.870 189.185 125.130 189.980 ;
        RECT 119.295 189.070 124.700 189.085 ;
        RECT 117.955 188.845 124.700 189.070 ;
        RECT 109.630 188.425 116.750 188.675 ;
        RECT 108.295 188.085 115.040 188.255 ;
        RECT 107.775 187.775 107.975 187.945 ;
        RECT 107.775 187.740 107.945 187.775 ;
        RECT 108.295 187.435 108.595 187.915 ;
        RECT 108.765 187.630 109.025 188.085 ;
        RECT 109.195 187.435 109.455 187.915 ;
        RECT 109.635 187.630 109.895 188.085 ;
        RECT 110.065 187.435 110.315 187.915 ;
        RECT 110.495 187.630 110.755 188.085 ;
        RECT 110.925 187.435 111.175 187.915 ;
        RECT 111.355 187.630 111.615 188.085 ;
        RECT 111.785 187.435 112.030 187.915 ;
        RECT 112.200 187.630 112.475 188.085 ;
        RECT 112.645 187.435 112.890 187.915 ;
        RECT 113.060 187.630 113.320 188.085 ;
        RECT 113.490 187.435 113.750 187.915 ;
        RECT 113.920 187.630 114.180 188.085 ;
        RECT 114.350 187.435 114.610 187.915 ;
        RECT 114.780 187.630 115.040 188.085 ;
        RECT 115.210 187.435 115.470 187.995 ;
        RECT 115.640 187.615 115.890 188.425 ;
        RECT 116.070 187.435 116.330 187.960 ;
        RECT 116.500 187.615 116.750 188.425 ;
        RECT 116.920 188.115 117.235 188.675 ;
        RECT 117.955 188.255 119.120 188.845 ;
        RECT 125.300 188.675 125.550 189.810 ;
        RECT 125.730 189.175 125.990 189.985 ;
        RECT 126.165 188.675 126.410 189.815 ;
        RECT 126.590 189.175 126.885 189.985 ;
        RECT 127.075 189.175 127.370 189.985 ;
        RECT 127.550 188.675 127.795 189.815 ;
        RECT 127.970 189.175 128.230 189.985 ;
        RECT 128.830 189.980 135.105 189.985 ;
        RECT 128.410 188.675 128.660 189.810 ;
        RECT 128.830 189.185 129.090 189.980 ;
        RECT 129.260 189.085 129.520 189.810 ;
        RECT 129.690 189.255 129.950 189.980 ;
        RECT 130.120 189.085 130.380 189.810 ;
        RECT 130.550 189.255 130.810 189.980 ;
        RECT 130.980 189.085 131.240 189.810 ;
        RECT 131.410 189.255 131.670 189.980 ;
        RECT 131.840 189.085 132.100 189.810 ;
        RECT 132.270 189.255 132.515 189.980 ;
        RECT 132.685 189.085 132.945 189.810 ;
        RECT 133.130 189.255 133.375 189.980 ;
        RECT 133.545 189.085 133.805 189.810 ;
        RECT 133.990 189.255 134.235 189.980 ;
        RECT 134.405 189.085 134.665 189.810 ;
        RECT 134.850 189.255 135.105 189.980 ;
        RECT 129.260 189.070 134.665 189.085 ;
        RECT 135.275 189.070 135.565 189.810 ;
        RECT 135.735 189.240 136.005 189.985 ;
        RECT 136.370 189.185 136.625 189.985 ;
        RECT 129.260 188.845 136.005 189.070 ;
        RECT 136.795 189.015 137.125 189.815 ;
        RECT 137.295 189.185 137.465 189.985 ;
        RECT 137.635 189.015 137.965 189.815 ;
        RECT 119.290 188.425 126.410 188.675 ;
        RECT 116.930 187.435 117.235 187.945 ;
        RECT 117.405 187.435 117.695 188.160 ;
        RECT 117.955 188.085 124.700 188.255 ;
        RECT 117.955 187.435 118.255 187.915 ;
        RECT 118.425 187.630 118.685 188.085 ;
        RECT 118.855 187.435 119.115 187.915 ;
        RECT 119.295 187.630 119.555 188.085 ;
        RECT 119.725 187.435 119.975 187.915 ;
        RECT 120.155 187.630 120.415 188.085 ;
        RECT 120.585 187.435 120.835 187.915 ;
        RECT 121.015 187.630 121.275 188.085 ;
        RECT 121.445 187.435 121.690 187.915 ;
        RECT 121.860 187.630 122.135 188.085 ;
        RECT 122.305 187.435 122.550 187.915 ;
        RECT 122.720 187.630 122.980 188.085 ;
        RECT 123.150 187.435 123.410 187.915 ;
        RECT 123.580 187.630 123.840 188.085 ;
        RECT 124.010 187.435 124.270 187.915 ;
        RECT 124.440 187.630 124.700 188.085 ;
        RECT 124.870 187.435 125.130 187.995 ;
        RECT 125.300 187.615 125.550 188.425 ;
        RECT 125.730 187.435 125.990 187.960 ;
        RECT 126.160 187.615 126.410 188.425 ;
        RECT 126.580 188.115 126.895 188.675 ;
        RECT 127.065 188.115 127.380 188.675 ;
        RECT 127.550 188.425 134.670 188.675 ;
        RECT 126.590 187.435 126.895 187.945 ;
        RECT 127.065 187.435 127.370 187.945 ;
        RECT 127.550 187.615 127.800 188.425 ;
        RECT 127.970 187.435 128.230 187.960 ;
        RECT 128.410 187.615 128.660 188.425 ;
        RECT 134.840 188.255 136.005 188.845 ;
        RECT 129.260 188.085 136.005 188.255 ;
        RECT 136.265 188.845 137.965 189.015 ;
        RECT 138.135 188.845 138.395 189.985 ;
        RECT 138.565 188.895 139.775 189.985 ;
        RECT 136.265 188.255 136.545 188.845 ;
        RECT 136.715 188.425 137.465 188.675 ;
        RECT 137.635 188.425 138.395 188.675 ;
        RECT 138.565 188.355 139.085 188.895 ;
        RECT 128.830 187.435 129.090 187.995 ;
        RECT 129.260 187.630 129.520 188.085 ;
        RECT 129.690 187.435 129.950 187.915 ;
        RECT 130.120 187.630 130.380 188.085 ;
        RECT 130.550 187.435 130.810 187.915 ;
        RECT 130.980 187.630 131.240 188.085 ;
        RECT 131.410 187.435 131.655 187.915 ;
        RECT 131.825 187.630 132.100 188.085 ;
        RECT 132.270 187.435 132.515 187.915 ;
        RECT 132.685 187.630 132.945 188.085 ;
        RECT 133.125 187.435 133.375 187.915 ;
        RECT 133.545 187.630 133.805 188.085 ;
        RECT 133.985 187.435 134.235 187.915 ;
        RECT 134.405 187.630 134.665 188.085 ;
        RECT 134.845 187.435 135.105 187.915 ;
        RECT 135.275 187.630 135.535 188.085 ;
        RECT 136.265 188.005 137.125 188.255 ;
        RECT 137.295 188.065 138.395 188.235 ;
        RECT 139.255 188.185 139.775 188.725 ;
        RECT 135.705 187.435 136.005 187.915 ;
        RECT 136.375 187.815 136.705 187.835 ;
        RECT 137.295 187.815 137.545 188.065 ;
        RECT 136.375 187.605 137.545 187.815 ;
        RECT 137.715 187.435 137.885 187.895 ;
        RECT 138.055 187.605 138.395 188.065 ;
        RECT 138.565 187.435 139.775 188.185 ;
        RECT 27.160 187.265 139.860 187.435 ;
        RECT 27.245 186.515 28.455 187.265 ;
        RECT 28.625 186.695 29.060 187.095 ;
        RECT 29.230 186.865 29.615 187.265 ;
        RECT 28.625 186.525 29.615 186.695 ;
        RECT 29.785 186.525 30.210 187.095 ;
        RECT 30.400 186.695 30.655 187.095 ;
        RECT 30.825 186.865 31.210 187.265 ;
        RECT 30.400 186.525 31.210 186.695 ;
        RECT 31.380 186.525 31.625 187.095 ;
        RECT 31.815 186.695 32.070 187.095 ;
        RECT 32.240 186.865 32.625 187.265 ;
        RECT 31.815 186.525 32.625 186.695 ;
        RECT 32.795 186.525 33.055 187.095 ;
        RECT 27.245 185.975 27.765 186.515 ;
        RECT 29.280 186.355 29.615 186.525 ;
        RECT 29.860 186.355 30.210 186.525 ;
        RECT 30.860 186.355 31.210 186.525 ;
        RECT 31.455 186.355 31.625 186.525 ;
        RECT 32.275 186.355 32.625 186.525 ;
        RECT 27.935 185.805 28.455 186.345 ;
        RECT 27.245 184.715 28.455 185.805 ;
        RECT 28.625 185.650 29.110 186.355 ;
        RECT 29.280 186.025 29.690 186.355 ;
        RECT 29.280 185.480 29.615 186.025 ;
        RECT 29.860 185.855 30.690 186.355 ;
        RECT 28.625 185.310 29.615 185.480 ;
        RECT 29.785 185.675 30.690 185.855 ;
        RECT 30.860 186.025 31.285 186.355 ;
        RECT 28.625 184.885 29.060 185.310 ;
        RECT 29.230 184.715 29.615 185.140 ;
        RECT 29.785 184.885 30.210 185.675 ;
        RECT 30.860 185.505 31.210 186.025 ;
        RECT 31.455 185.855 32.105 186.355 ;
        RECT 30.380 185.310 31.210 185.505 ;
        RECT 31.380 185.675 32.105 185.855 ;
        RECT 32.275 186.025 32.700 186.355 ;
        RECT 30.380 184.885 30.655 185.310 ;
        RECT 30.825 184.715 31.210 185.140 ;
        RECT 31.380 184.885 31.625 185.675 ;
        RECT 32.275 185.505 32.625 186.025 ;
        RECT 32.870 185.855 33.055 186.525 ;
        RECT 33.225 186.495 34.895 187.265 ;
        RECT 35.535 186.760 35.865 187.265 ;
        RECT 36.035 186.695 36.275 187.070 ;
        RECT 36.555 186.935 36.725 187.080 ;
        RECT 36.555 186.740 36.955 186.935 ;
        RECT 37.315 186.770 37.715 187.265 ;
        RECT 33.225 185.975 33.975 186.495 ;
        RECT 31.815 185.310 32.625 185.505 ;
        RECT 31.815 184.885 32.070 185.310 ;
        RECT 32.240 184.715 32.625 185.140 ;
        RECT 32.795 184.885 33.055 185.855 ;
        RECT 34.145 185.805 34.895 186.325 ;
        RECT 35.590 185.905 35.890 186.585 ;
        RECT 33.225 184.715 34.895 185.805 ;
        RECT 35.585 185.735 35.890 185.905 ;
        RECT 36.060 186.545 36.275 186.695 ;
        RECT 36.060 186.215 36.615 186.545 ;
        RECT 36.785 186.405 36.955 186.740 ;
        RECT 37.885 186.575 38.120 187.095 ;
        RECT 38.305 186.630 38.575 187.265 ;
        RECT 38.830 186.695 39.005 187.095 ;
        RECT 39.175 186.885 39.505 187.265 ;
        RECT 39.750 186.765 39.980 187.095 ;
        RECT 36.060 185.565 36.295 186.215 ;
        RECT 36.785 186.045 37.775 186.405 ;
        RECT 35.615 185.335 36.295 185.565 ;
        RECT 36.485 186.025 37.775 186.045 ;
        RECT 36.485 185.875 37.345 186.025 ;
        RECT 35.615 184.905 35.785 185.335 ;
        RECT 35.955 184.715 36.285 185.165 ;
        RECT 36.485 184.930 36.770 185.875 ;
        RECT 37.945 185.770 38.120 186.575 ;
        RECT 38.830 186.525 39.460 186.695 ;
        RECT 39.290 186.355 39.460 186.525 ;
        RECT 36.945 185.395 37.640 185.705 ;
        RECT 36.950 184.715 37.635 185.185 ;
        RECT 37.815 184.985 38.120 185.770 ;
        RECT 38.745 185.675 39.110 186.355 ;
        RECT 39.290 186.025 39.640 186.355 ;
        RECT 38.305 184.715 38.575 185.670 ;
        RECT 39.290 185.505 39.460 186.025 ;
        RECT 38.830 185.335 39.460 185.505 ;
        RECT 39.810 185.475 39.980 186.765 ;
        RECT 40.180 185.655 40.460 186.930 ;
        RECT 40.685 185.905 40.955 186.930 ;
        RECT 41.415 186.885 41.745 187.265 ;
        RECT 41.915 187.010 42.250 187.055 ;
        RECT 40.645 185.735 40.955 185.905 ;
        RECT 40.685 185.655 40.955 185.735 ;
        RECT 41.145 185.655 41.485 186.685 ;
        RECT 41.915 186.545 42.255 187.010 ;
        RECT 41.655 186.025 41.915 186.355 ;
        RECT 41.655 185.475 41.825 186.025 ;
        RECT 42.085 185.855 42.255 186.545 ;
        RECT 42.425 186.445 42.685 187.265 ;
        RECT 42.855 186.445 43.185 186.865 ;
        RECT 43.365 186.780 44.155 187.045 ;
        RECT 42.935 186.355 43.185 186.445 ;
        RECT 38.830 184.885 39.005 185.335 ;
        RECT 39.810 185.305 41.825 185.475 ;
        RECT 39.175 184.715 39.505 185.155 ;
        RECT 39.810 184.885 39.980 185.305 ;
        RECT 40.215 184.715 40.885 185.125 ;
        RECT 41.100 184.885 41.270 185.305 ;
        RECT 41.470 184.715 41.800 185.125 ;
        RECT 41.995 184.885 42.255 185.855 ;
        RECT 42.425 185.395 42.765 186.275 ;
        RECT 42.935 186.105 43.730 186.355 ;
        RECT 42.425 184.715 42.685 185.225 ;
        RECT 42.935 184.885 43.105 186.105 ;
        RECT 43.900 185.925 44.155 186.780 ;
        RECT 44.325 186.625 44.525 187.045 ;
        RECT 44.715 186.805 45.045 187.265 ;
        RECT 44.325 186.105 44.735 186.625 ;
        RECT 45.215 186.615 45.475 187.095 ;
        RECT 45.650 186.760 45.985 187.265 ;
        RECT 46.155 186.695 46.395 187.070 ;
        RECT 46.675 186.935 46.845 187.080 ;
        RECT 46.675 186.740 47.050 186.935 ;
        RECT 47.410 186.770 47.805 187.265 ;
        RECT 44.905 185.925 45.135 186.355 ;
        RECT 43.345 185.755 45.135 185.925 ;
        RECT 43.345 185.390 43.595 185.755 ;
        RECT 43.765 185.395 44.095 185.585 ;
        RECT 44.315 185.460 45.030 185.755 ;
        RECT 45.305 185.585 45.475 186.615 ;
        RECT 45.705 185.735 46.005 186.585 ;
        RECT 46.175 186.545 46.395 186.695 ;
        RECT 46.175 186.215 46.710 186.545 ;
        RECT 46.880 186.405 47.050 186.740 ;
        RECT 47.975 186.575 48.215 187.095 ;
        RECT 43.765 185.220 43.960 185.395 ;
        RECT 43.345 184.715 43.960 185.220 ;
        RECT 44.130 184.885 44.605 185.225 ;
        RECT 44.775 184.715 44.990 185.260 ;
        RECT 45.200 184.885 45.475 185.585 ;
        RECT 46.175 185.565 46.410 186.215 ;
        RECT 46.880 186.045 47.865 186.405 ;
        RECT 45.735 185.335 46.410 185.565 ;
        RECT 46.580 186.025 47.865 186.045 ;
        RECT 46.580 185.875 47.440 186.025 ;
        RECT 45.735 184.905 45.905 185.335 ;
        RECT 46.075 184.715 46.405 185.165 ;
        RECT 46.580 184.930 46.865 185.875 ;
        RECT 48.040 185.770 48.215 186.575 ;
        RECT 47.040 185.395 47.735 185.705 ;
        RECT 47.045 184.715 47.730 185.185 ;
        RECT 47.910 184.985 48.215 185.770 ;
        RECT 49.325 186.805 49.885 187.095 ;
        RECT 50.055 186.805 50.305 187.265 ;
        RECT 49.325 185.435 49.575 186.805 ;
        RECT 50.925 186.635 51.255 186.995 ;
        RECT 49.865 186.445 51.255 186.635 ;
        RECT 51.625 186.515 52.835 187.265 ;
        RECT 53.005 186.540 53.295 187.265 ;
        RECT 53.620 186.615 53.950 187.080 ;
        RECT 54.120 186.795 54.290 187.265 ;
        RECT 54.460 186.615 54.790 187.095 ;
        RECT 49.865 186.355 50.035 186.445 ;
        RECT 49.745 186.025 50.035 186.355 ;
        RECT 50.205 186.025 50.545 186.275 ;
        RECT 50.765 186.025 51.440 186.275 ;
        RECT 49.865 185.775 50.035 186.025 ;
        RECT 49.865 185.605 50.805 185.775 ;
        RECT 51.175 185.665 51.440 186.025 ;
        RECT 51.625 185.975 52.145 186.515 ;
        RECT 53.620 186.445 54.790 186.615 ;
        RECT 52.315 185.805 52.835 186.345 ;
        RECT 53.465 186.065 54.110 186.275 ;
        RECT 54.280 186.065 54.850 186.275 ;
        RECT 55.020 185.895 55.190 187.095 ;
        RECT 55.730 186.695 55.900 186.900 ;
        RECT 49.325 184.885 49.785 185.435 ;
        RECT 49.975 184.715 50.305 185.435 ;
        RECT 50.505 185.055 50.805 185.605 ;
        RECT 50.975 184.715 51.255 185.385 ;
        RECT 51.625 184.715 52.835 185.805 ;
        RECT 53.005 184.715 53.295 185.880 ;
        RECT 53.680 184.715 54.010 185.815 ;
        RECT 54.485 185.485 55.190 185.895 ;
        RECT 55.360 186.525 55.900 186.695 ;
        RECT 56.180 186.525 56.350 187.265 ;
        RECT 56.615 186.525 56.975 186.900 ;
        RECT 57.145 186.720 62.490 187.265 ;
        RECT 55.360 185.825 55.530 186.525 ;
        RECT 55.700 186.025 56.030 186.355 ;
        RECT 56.200 186.025 56.550 186.355 ;
        RECT 55.360 185.655 55.985 185.825 ;
        RECT 56.200 185.485 56.465 186.025 ;
        RECT 56.720 185.870 56.975 186.525 ;
        RECT 58.730 185.890 59.070 186.720 ;
        RECT 62.665 186.495 65.255 187.265 ;
        RECT 54.485 185.315 56.465 185.485 ;
        RECT 54.485 184.885 54.810 185.315 ;
        RECT 54.980 184.715 55.310 185.135 ;
        RECT 56.055 184.715 56.465 185.145 ;
        RECT 56.635 184.885 56.975 185.870 ;
        RECT 60.550 185.150 60.900 186.400 ;
        RECT 62.665 185.975 63.875 186.495 ;
        RECT 65.425 186.465 65.735 187.265 ;
        RECT 65.940 186.465 66.635 187.095 ;
        RECT 66.805 186.495 68.475 187.265 ;
        RECT 68.645 186.625 68.985 187.030 ;
        RECT 69.155 186.795 69.325 187.265 ;
        RECT 69.495 186.625 69.745 187.030 ;
        RECT 64.045 185.805 65.255 186.325 ;
        RECT 65.435 186.025 65.770 186.295 ;
        RECT 65.940 185.865 66.110 186.465 ;
        RECT 66.280 186.025 66.615 186.275 ;
        RECT 66.805 185.975 67.555 186.495 ;
        RECT 68.645 186.445 69.745 186.625 ;
        RECT 69.915 186.660 70.165 187.030 ;
        RECT 70.335 186.785 70.780 186.955 ;
        RECT 70.950 186.925 71.170 186.970 ;
        RECT 57.145 184.715 62.490 185.150 ;
        RECT 62.665 184.715 65.255 185.805 ;
        RECT 65.425 184.715 65.705 185.855 ;
        RECT 65.875 184.885 66.205 185.865 ;
        RECT 66.375 184.715 66.635 185.855 ;
        RECT 67.725 185.805 68.475 186.325 ;
        RECT 69.915 186.275 70.085 186.660 ;
        RECT 66.805 184.715 68.475 185.805 ;
        RECT 68.645 185.705 68.990 186.275 ;
        RECT 69.160 186.025 69.720 186.275 ;
        RECT 69.890 186.105 70.085 186.275 ;
        RECT 68.645 184.715 68.990 185.535 ;
        RECT 69.160 184.925 69.335 186.025 ;
        RECT 69.890 185.855 70.060 186.105 ;
        RECT 70.335 185.995 70.505 186.785 ;
        RECT 70.950 186.755 71.175 186.925 ;
        RECT 70.950 186.615 71.170 186.755 ;
        RECT 70.675 186.445 71.170 186.615 ;
        RECT 71.450 186.600 71.620 187.265 ;
        RECT 71.815 186.525 72.155 187.095 ;
        RECT 70.675 186.250 70.850 186.445 ;
        RECT 71.020 186.075 71.470 186.275 ;
        RECT 69.505 185.465 70.060 185.855 ;
        RECT 70.230 185.855 70.505 185.995 ;
        RECT 71.640 185.905 71.810 186.355 ;
        RECT 70.230 185.635 71.245 185.855 ;
        RECT 71.415 185.735 71.810 185.905 ;
        RECT 71.415 185.465 71.585 185.735 ;
        RECT 71.980 185.555 72.155 186.525 ;
        RECT 69.505 185.295 71.585 185.465 ;
        RECT 69.505 185.060 69.835 185.295 ;
        RECT 70.125 184.715 70.525 185.115 ;
        RECT 71.395 184.715 71.725 185.115 ;
        RECT 71.895 184.885 72.155 185.555 ;
        RECT 72.325 186.465 72.665 187.095 ;
        RECT 72.835 186.465 73.085 187.265 ;
        RECT 73.275 186.615 73.605 187.095 ;
        RECT 73.775 186.805 74.000 187.265 ;
        RECT 74.170 186.615 74.500 187.095 ;
        RECT 72.325 185.855 72.500 186.465 ;
        RECT 73.275 186.445 74.500 186.615 ;
        RECT 75.130 186.485 75.630 187.095 ;
        RECT 76.040 186.525 76.655 187.095 ;
        RECT 76.825 186.755 77.040 187.265 ;
        RECT 77.270 186.755 77.550 187.085 ;
        RECT 77.730 186.755 77.970 187.265 ;
        RECT 72.670 186.105 73.365 186.275 ;
        RECT 73.195 185.855 73.365 186.105 ;
        RECT 73.540 186.075 73.960 186.275 ;
        RECT 74.130 186.075 74.460 186.275 ;
        RECT 74.630 186.075 74.960 186.275 ;
        RECT 75.130 185.855 75.300 186.485 ;
        RECT 75.485 186.025 75.835 186.275 ;
        RECT 72.325 184.885 72.665 185.855 ;
        RECT 72.835 184.715 73.005 185.855 ;
        RECT 73.195 185.685 75.630 185.855 ;
        RECT 73.275 184.715 73.525 185.515 ;
        RECT 74.170 184.885 74.500 185.685 ;
        RECT 74.800 184.715 75.130 185.515 ;
        RECT 75.300 184.885 75.630 185.685 ;
        RECT 76.040 185.505 76.355 186.525 ;
        RECT 76.525 185.855 76.695 186.355 ;
        RECT 76.945 186.025 77.210 186.585 ;
        RECT 77.380 185.855 77.550 186.755 ;
        RECT 77.720 186.025 78.075 186.585 ;
        RECT 78.765 186.540 79.055 187.265 ;
        RECT 79.225 186.465 79.920 187.095 ;
        RECT 80.125 186.465 80.435 187.265 ;
        RECT 80.630 186.875 80.960 187.265 ;
        RECT 81.130 186.705 81.355 187.085 ;
        RECT 79.245 186.025 79.580 186.275 ;
        RECT 76.525 185.685 77.950 185.855 ;
        RECT 76.040 184.885 76.575 185.505 ;
        RECT 76.745 184.715 77.075 185.515 ;
        RECT 77.560 185.510 77.950 185.685 ;
        RECT 78.765 184.715 79.055 185.880 ;
        RECT 79.750 185.865 79.920 186.465 ;
        RECT 80.090 186.025 80.425 186.295 ;
        RECT 80.615 186.025 80.855 186.675 ;
        RECT 81.025 186.525 81.355 186.705 ;
        RECT 79.225 184.715 79.485 185.855 ;
        RECT 79.655 184.885 79.985 185.865 ;
        RECT 81.025 185.855 81.200 186.525 ;
        RECT 81.555 186.355 81.785 186.975 ;
        RECT 81.965 186.535 82.265 187.265 ;
        RECT 82.470 186.875 82.800 187.265 ;
        RECT 82.970 186.705 83.195 187.085 ;
        RECT 81.370 186.025 81.785 186.355 ;
        RECT 81.965 186.025 82.260 186.355 ;
        RECT 82.455 186.025 82.695 186.675 ;
        RECT 82.865 186.525 83.195 186.705 ;
        RECT 82.865 185.855 83.040 186.525 ;
        RECT 83.395 186.355 83.625 186.975 ;
        RECT 83.805 186.535 84.105 187.265 ;
        RECT 84.310 186.875 84.640 187.265 ;
        RECT 84.810 186.705 85.035 187.085 ;
        RECT 83.210 186.025 83.625 186.355 ;
        RECT 83.805 186.025 84.100 186.355 ;
        RECT 84.295 186.025 84.535 186.675 ;
        RECT 84.705 186.525 85.035 186.705 ;
        RECT 84.705 185.855 84.880 186.525 ;
        RECT 85.235 186.355 85.465 186.975 ;
        RECT 85.645 186.535 85.945 187.265 ;
        RECT 85.050 186.025 85.465 186.355 ;
        RECT 85.645 186.025 85.940 186.355 ;
        RECT 80.155 184.715 80.435 185.855 ;
        RECT 80.615 185.665 81.200 185.855 ;
        RECT 80.615 184.895 80.890 185.665 ;
        RECT 81.370 185.495 82.265 185.825 ;
        RECT 81.060 185.325 82.265 185.495 ;
        RECT 81.060 184.895 81.390 185.325 ;
        RECT 81.560 184.715 81.755 185.155 ;
        RECT 81.935 184.895 82.265 185.325 ;
        RECT 82.455 185.665 83.040 185.855 ;
        RECT 82.455 184.895 82.730 185.665 ;
        RECT 83.210 185.495 84.105 185.825 ;
        RECT 82.900 185.325 84.105 185.495 ;
        RECT 82.900 184.895 83.230 185.325 ;
        RECT 83.400 184.715 83.595 185.155 ;
        RECT 83.775 184.895 84.105 185.325 ;
        RECT 84.295 185.665 84.880 185.855 ;
        RECT 84.295 184.895 84.570 185.665 ;
        RECT 85.050 185.495 85.945 185.825 ;
        RECT 86.145 185.685 86.375 187.025 ;
        RECT 86.555 186.185 86.785 187.085 ;
        RECT 86.985 186.485 87.230 187.265 ;
        RECT 87.400 186.725 87.830 187.085 ;
        RECT 88.410 186.895 89.140 187.265 ;
        RECT 87.400 186.535 89.140 186.725 ;
        RECT 87.400 186.305 87.620 186.535 ;
        RECT 86.555 185.505 86.895 186.185 ;
        RECT 84.740 185.325 85.945 185.495 ;
        RECT 84.740 184.895 85.070 185.325 ;
        RECT 85.240 184.715 85.435 185.155 ;
        RECT 85.615 184.895 85.945 185.325 ;
        RECT 86.145 185.305 86.895 185.505 ;
        RECT 87.075 186.005 87.620 186.305 ;
        RECT 86.145 184.915 86.385 185.305 ;
        RECT 86.555 184.715 86.905 185.125 ;
        RECT 87.075 184.895 87.405 186.005 ;
        RECT 87.790 185.735 88.215 186.355 ;
        RECT 88.410 185.735 88.670 186.355 ;
        RECT 88.880 186.025 89.140 186.535 ;
        RECT 87.575 185.365 88.600 185.565 ;
        RECT 87.575 184.895 87.755 185.365 ;
        RECT 87.925 184.715 88.255 185.195 ;
        RECT 88.430 184.895 88.600 185.365 ;
        RECT 88.865 184.715 89.150 185.855 ;
        RECT 89.340 184.895 89.620 187.085 ;
        RECT 90.725 186.465 91.420 187.095 ;
        RECT 91.625 186.465 91.935 187.265 ;
        RECT 92.115 186.755 92.565 187.265 ;
        RECT 92.840 186.845 94.145 187.095 ;
        RECT 94.325 186.865 94.655 187.265 ;
        RECT 93.965 186.695 94.145 186.845 ;
        RECT 94.865 186.765 95.125 187.095 ;
        RECT 95.295 186.905 95.625 187.265 ;
        RECT 95.880 186.885 97.180 187.095 ;
        RECT 94.865 186.755 95.095 186.765 ;
        RECT 90.745 186.025 91.080 186.275 ;
        RECT 91.250 185.865 91.420 186.465 ;
        RECT 91.590 186.025 91.925 186.295 ;
        RECT 92.145 186.075 92.595 186.585 ;
        RECT 93.010 186.275 93.260 186.675 ;
        RECT 92.785 186.075 93.260 186.275 ;
        RECT 93.510 186.275 93.720 186.675 ;
        RECT 93.965 186.525 94.695 186.695 ;
        RECT 93.510 186.075 93.860 186.275 ;
        RECT 94.030 186.025 94.355 186.355 ;
        RECT 90.725 184.715 90.985 185.855 ;
        RECT 91.155 184.885 91.485 185.865 ;
        RECT 92.115 185.855 93.860 185.905 ;
        RECT 94.525 185.855 94.695 186.525 ;
        RECT 91.655 184.715 91.935 185.855 ;
        RECT 92.115 185.725 94.695 185.855 ;
        RECT 92.115 185.055 92.445 185.725 ;
        RECT 93.635 185.685 94.695 185.725 ;
        RECT 94.865 185.565 95.035 186.755 ;
        RECT 95.880 186.735 96.050 186.885 ;
        RECT 95.295 186.610 96.050 186.735 ;
        RECT 95.205 186.565 96.050 186.610 ;
        RECT 95.205 186.445 95.475 186.565 ;
        RECT 95.205 185.870 95.375 186.445 ;
        RECT 95.605 186.005 96.015 186.310 ;
        RECT 96.305 186.275 96.515 186.675 ;
        RECT 96.185 186.065 96.515 186.275 ;
        RECT 96.760 186.275 96.980 186.675 ;
        RECT 97.455 186.500 97.910 187.265 ;
        RECT 98.245 186.705 98.575 187.095 ;
        RECT 98.745 186.875 99.930 187.045 ;
        RECT 100.190 186.795 100.360 187.265 ;
        RECT 98.245 186.525 98.755 186.705 ;
        RECT 96.760 186.065 97.235 186.275 ;
        RECT 97.425 186.075 97.915 186.275 ;
        RECT 98.085 186.065 98.415 186.355 ;
        RECT 98.585 185.895 98.755 186.525 ;
        RECT 99.160 186.615 99.545 186.705 ;
        RECT 100.530 186.615 100.860 187.080 ;
        RECT 99.160 186.445 100.860 186.615 ;
        RECT 101.030 186.445 101.200 187.265 ;
        RECT 101.370 186.445 102.055 187.085 ;
        RECT 102.695 186.535 102.995 187.265 ;
        RECT 98.925 186.065 99.255 186.275 ;
        RECT 99.435 186.025 99.815 186.275 ;
        RECT 95.205 185.835 95.405 185.870 ;
        RECT 96.735 185.835 97.910 185.895 ;
        RECT 95.205 185.725 97.910 185.835 ;
        RECT 95.265 185.665 97.065 185.725 ;
        RECT 96.735 185.635 97.065 185.665 ;
        RECT 92.615 185.515 93.495 185.555 ;
        RECT 92.615 185.315 94.145 185.515 ;
        RECT 92.615 185.265 93.230 185.315 ;
        RECT 92.615 185.225 92.845 185.265 ;
        RECT 93.975 185.185 94.145 185.315 ;
        RECT 92.955 185.055 93.285 185.095 ;
        RECT 92.115 184.885 93.285 185.055 ;
        RECT 93.455 184.715 93.830 185.095 ;
        RECT 94.380 184.715 94.645 185.495 ;
        RECT 94.865 184.885 95.125 185.565 ;
        RECT 95.295 184.715 95.545 185.495 ;
        RECT 95.795 185.465 96.630 185.475 ;
        RECT 97.220 185.465 97.405 185.555 ;
        RECT 95.795 185.265 97.405 185.465 ;
        RECT 95.795 184.885 96.045 185.265 ;
        RECT 97.175 185.225 97.405 185.265 ;
        RECT 97.655 185.105 97.910 185.725 ;
        RECT 96.215 184.715 96.570 185.095 ;
        RECT 97.575 184.885 97.910 185.105 ;
        RECT 98.240 185.725 99.325 185.895 ;
        RECT 98.240 184.885 98.540 185.725 ;
        RECT 98.735 184.715 98.985 185.555 ;
        RECT 99.155 185.475 99.325 185.725 ;
        RECT 99.495 185.645 99.815 186.025 ;
        RECT 100.005 186.065 100.490 186.275 ;
        RECT 100.680 186.065 101.130 186.275 ;
        RECT 101.300 186.065 101.635 186.275 ;
        RECT 100.005 185.905 100.380 186.065 ;
        RECT 99.985 185.735 100.380 185.905 ;
        RECT 101.300 185.895 101.470 186.065 ;
        RECT 100.005 185.645 100.380 185.735 ;
        RECT 100.550 185.725 101.470 185.895 ;
        RECT 100.550 185.475 100.720 185.725 ;
        RECT 99.155 185.305 100.720 185.475 ;
        RECT 99.575 184.885 100.380 185.305 ;
        RECT 100.890 184.715 101.220 185.555 ;
        RECT 101.805 185.475 102.055 186.445 ;
        RECT 103.175 186.355 103.405 186.975 ;
        RECT 103.605 186.705 103.830 187.085 ;
        RECT 104.000 186.875 104.330 187.265 ;
        RECT 103.605 186.525 103.935 186.705 ;
        RECT 102.700 186.025 102.995 186.355 ;
        RECT 103.175 186.025 103.590 186.355 ;
        RECT 103.760 185.855 103.935 186.525 ;
        RECT 104.105 186.025 104.345 186.675 ;
        RECT 104.525 186.540 104.815 187.265 ;
        RECT 104.985 186.465 105.680 187.095 ;
        RECT 105.885 186.465 106.195 187.265 ;
        RECT 105.005 186.025 105.340 186.275 ;
        RECT 101.390 184.885 102.055 185.475 ;
        RECT 102.695 185.495 103.590 185.825 ;
        RECT 103.760 185.665 104.345 185.855 ;
        RECT 102.695 185.325 103.900 185.495 ;
        RECT 102.695 184.895 103.025 185.325 ;
        RECT 103.205 184.715 103.400 185.155 ;
        RECT 103.570 184.895 103.900 185.325 ;
        RECT 104.070 184.895 104.345 185.665 ;
        RECT 104.525 184.715 104.815 185.880 ;
        RECT 105.510 185.865 105.680 186.465 ;
        RECT 105.850 186.025 106.185 186.295 ;
        RECT 104.985 184.715 105.245 185.855 ;
        RECT 105.415 184.885 105.745 185.865 ;
        RECT 105.915 184.715 106.195 185.855 ;
        RECT 106.380 184.895 106.660 187.085 ;
        RECT 106.860 186.895 107.590 187.265 ;
        RECT 108.170 186.725 108.600 187.085 ;
        RECT 106.860 186.535 108.600 186.725 ;
        RECT 106.860 186.025 107.120 186.535 ;
        RECT 106.850 184.715 107.135 185.855 ;
        RECT 107.330 185.735 107.590 186.355 ;
        RECT 107.785 185.735 108.210 186.355 ;
        RECT 108.380 186.305 108.600 186.535 ;
        RECT 108.770 186.485 109.015 187.265 ;
        RECT 108.380 186.005 108.925 186.305 ;
        RECT 109.215 186.185 109.445 187.085 ;
        RECT 107.400 185.365 108.425 185.565 ;
        RECT 107.400 184.895 107.570 185.365 ;
        RECT 107.745 184.715 108.075 185.195 ;
        RECT 108.245 184.895 108.425 185.365 ;
        RECT 108.595 184.895 108.925 186.005 ;
        RECT 109.105 185.505 109.445 186.185 ;
        RECT 109.625 185.685 109.855 187.025 ;
        RECT 110.505 186.755 110.810 187.265 ;
        RECT 110.505 186.025 110.820 186.585 ;
        RECT 110.990 186.275 111.240 187.085 ;
        RECT 111.410 186.740 111.670 187.265 ;
        RECT 111.850 186.275 112.100 187.085 ;
        RECT 112.270 186.705 112.530 187.265 ;
        RECT 112.700 186.615 112.960 187.070 ;
        RECT 113.130 186.785 113.390 187.265 ;
        RECT 113.560 186.615 113.820 187.070 ;
        RECT 113.990 186.785 114.250 187.265 ;
        RECT 114.420 186.615 114.680 187.070 ;
        RECT 114.850 186.785 115.095 187.265 ;
        RECT 115.265 186.615 115.540 187.070 ;
        RECT 115.710 186.785 115.955 187.265 ;
        RECT 116.125 186.615 116.385 187.070 ;
        RECT 116.565 186.785 116.815 187.265 ;
        RECT 116.985 186.615 117.245 187.070 ;
        RECT 117.425 186.785 117.675 187.265 ;
        RECT 117.845 186.615 118.105 187.070 ;
        RECT 118.285 186.785 118.545 187.265 ;
        RECT 118.715 186.615 118.975 187.070 ;
        RECT 119.145 186.785 119.445 187.265 ;
        RECT 119.705 186.755 120.010 187.265 ;
        RECT 112.700 186.445 119.445 186.615 ;
        RECT 110.990 186.025 118.110 186.275 ;
        RECT 109.105 185.305 109.855 185.505 ;
        RECT 109.095 184.715 109.445 185.125 ;
        RECT 109.615 184.915 109.855 185.305 ;
        RECT 110.515 184.715 110.810 185.525 ;
        RECT 110.990 184.885 111.235 186.025 ;
        RECT 111.410 184.715 111.670 185.525 ;
        RECT 111.850 184.890 112.100 186.025 ;
        RECT 118.280 185.855 119.445 186.445 ;
        RECT 119.705 186.025 120.020 186.585 ;
        RECT 120.190 186.275 120.440 187.085 ;
        RECT 120.610 186.740 120.870 187.265 ;
        RECT 121.050 186.275 121.300 187.085 ;
        RECT 121.470 186.705 121.730 187.265 ;
        RECT 121.900 186.615 122.160 187.070 ;
        RECT 122.330 186.785 122.590 187.265 ;
        RECT 122.760 186.615 123.020 187.070 ;
        RECT 123.190 186.785 123.450 187.265 ;
        RECT 123.620 186.615 123.880 187.070 ;
        RECT 124.050 186.785 124.295 187.265 ;
        RECT 124.465 186.615 124.740 187.070 ;
        RECT 124.910 186.785 125.155 187.265 ;
        RECT 125.325 186.615 125.585 187.070 ;
        RECT 125.765 186.785 126.015 187.265 ;
        RECT 126.185 186.615 126.445 187.070 ;
        RECT 126.625 186.785 126.875 187.265 ;
        RECT 127.045 186.615 127.305 187.070 ;
        RECT 127.485 186.785 127.745 187.265 ;
        RECT 127.915 186.615 128.175 187.070 ;
        RECT 128.345 186.785 128.645 187.265 ;
        RECT 121.900 186.585 128.645 186.615 ;
        RECT 121.900 186.445 128.675 186.585 ;
        RECT 128.925 186.455 129.165 187.265 ;
        RECT 129.335 186.455 129.665 187.095 ;
        RECT 129.835 186.455 130.105 187.265 ;
        RECT 130.285 186.540 130.575 187.265 ;
        RECT 130.750 186.885 132.765 187.055 ;
        RECT 132.955 186.885 133.285 187.265 ;
        RECT 130.750 186.565 131.005 186.885 ;
        RECT 127.480 186.415 128.675 186.445 ;
        RECT 120.190 186.025 127.310 186.275 ;
        RECT 112.700 185.630 119.445 185.855 ;
        RECT 112.700 185.615 118.105 185.630 ;
        RECT 112.270 184.720 112.530 185.515 ;
        RECT 112.700 184.890 112.960 185.615 ;
        RECT 113.130 184.720 113.390 185.445 ;
        RECT 113.560 184.890 113.820 185.615 ;
        RECT 113.990 184.720 114.250 185.445 ;
        RECT 114.420 184.890 114.680 185.615 ;
        RECT 114.850 184.720 115.110 185.445 ;
        RECT 115.280 184.890 115.540 185.615 ;
        RECT 115.710 184.720 115.955 185.445 ;
        RECT 116.125 184.890 116.385 185.615 ;
        RECT 116.570 184.720 116.815 185.445 ;
        RECT 116.985 184.890 117.245 185.615 ;
        RECT 117.430 184.720 117.675 185.445 ;
        RECT 117.845 184.890 118.105 185.615 ;
        RECT 118.290 184.720 118.545 185.445 ;
        RECT 118.715 184.890 119.005 185.630 ;
        RECT 112.270 184.715 118.545 184.720 ;
        RECT 119.175 184.715 119.445 185.460 ;
        RECT 119.715 184.715 120.010 185.525 ;
        RECT 120.190 184.885 120.435 186.025 ;
        RECT 120.610 184.715 120.870 185.525 ;
        RECT 121.050 184.890 121.300 186.025 ;
        RECT 127.480 185.855 128.645 186.415 ;
        RECT 128.905 186.025 129.255 186.275 ;
        RECT 129.425 185.855 129.595 186.455 ;
        RECT 129.765 186.025 130.115 186.275 ;
        RECT 130.750 186.025 130.990 186.355 ;
        RECT 131.175 185.905 131.505 186.715 ;
        RECT 132.015 186.445 133.705 186.715 ;
        RECT 133.875 186.465 134.255 187.265 ;
        RECT 131.730 186.075 132.820 186.275 ;
        RECT 133.130 186.245 134.255 186.275 ;
        RECT 133.105 186.075 134.255 186.245 ;
        RECT 121.900 185.630 128.645 185.855 ;
        RECT 128.915 185.685 129.595 185.855 ;
        RECT 121.900 185.615 127.305 185.630 ;
        RECT 121.470 184.720 121.730 185.515 ;
        RECT 121.900 184.890 122.160 185.615 ;
        RECT 122.330 184.720 122.590 185.445 ;
        RECT 122.760 184.890 123.020 185.615 ;
        RECT 123.190 184.720 123.450 185.445 ;
        RECT 123.620 184.890 123.880 185.615 ;
        RECT 124.050 184.720 124.310 185.445 ;
        RECT 124.480 184.890 124.740 185.615 ;
        RECT 124.910 184.720 125.155 185.445 ;
        RECT 125.325 184.890 125.585 185.615 ;
        RECT 125.770 184.720 126.015 185.445 ;
        RECT 126.185 184.890 126.445 185.615 ;
        RECT 126.630 184.720 126.875 185.445 ;
        RECT 127.045 184.890 127.305 185.615 ;
        RECT 127.490 184.720 127.745 185.445 ;
        RECT 127.915 184.890 128.205 185.630 ;
        RECT 121.470 184.715 127.745 184.720 ;
        RECT 128.375 184.715 128.645 185.460 ;
        RECT 128.915 184.900 129.245 185.685 ;
        RECT 129.775 184.715 130.105 185.855 ;
        RECT 130.285 184.715 130.575 185.880 ;
        RECT 130.750 184.715 131.005 185.855 ;
        RECT 131.175 185.685 133.705 185.905 ;
        RECT 131.175 184.885 131.505 185.685 ;
        RECT 131.675 184.715 131.845 185.515 ;
        RECT 132.015 184.885 132.345 185.685 ;
        RECT 132.515 184.715 133.205 185.515 ;
        RECT 133.375 184.885 133.705 185.685 ;
        RECT 133.875 184.715 134.255 185.905 ;
        RECT 134.445 185.685 134.675 187.025 ;
        RECT 134.855 186.185 135.085 187.085 ;
        RECT 135.285 186.485 135.530 187.265 ;
        RECT 135.700 186.725 136.130 187.085 ;
        RECT 136.710 186.895 137.440 187.265 ;
        RECT 135.700 186.535 137.440 186.725 ;
        RECT 135.700 186.305 135.920 186.535 ;
        RECT 134.855 185.505 135.195 186.185 ;
        RECT 134.445 185.305 135.195 185.505 ;
        RECT 135.375 186.005 135.920 186.305 ;
        RECT 134.445 184.915 134.685 185.305 ;
        RECT 134.855 184.715 135.205 185.125 ;
        RECT 135.375 184.895 135.705 186.005 ;
        RECT 136.090 185.735 136.515 186.355 ;
        RECT 136.710 185.735 136.970 186.355 ;
        RECT 137.180 186.025 137.440 186.535 ;
        RECT 135.875 185.365 136.900 185.565 ;
        RECT 135.875 184.895 136.055 185.365 ;
        RECT 136.225 184.715 136.555 185.195 ;
        RECT 136.730 184.895 136.900 185.365 ;
        RECT 137.165 184.715 137.450 185.855 ;
        RECT 137.640 184.895 137.920 187.085 ;
        RECT 138.565 186.515 139.775 187.265 ;
        RECT 138.565 185.805 139.085 186.345 ;
        RECT 139.255 185.975 139.775 186.515 ;
        RECT 138.565 184.715 139.775 185.805 ;
        RECT 27.160 184.545 139.860 184.715 ;
        RECT 27.245 183.455 28.455 184.545 ;
        RECT 27.245 182.745 27.765 183.285 ;
        RECT 27.935 182.915 28.455 183.455 ;
        RECT 28.625 183.575 28.895 184.345 ;
        RECT 29.065 183.765 29.395 184.545 ;
        RECT 29.600 183.940 29.785 184.345 ;
        RECT 29.955 184.120 30.290 184.545 ;
        RECT 29.600 183.765 30.265 183.940 ;
        RECT 31.125 183.875 31.405 184.545 ;
        RECT 28.625 183.405 29.755 183.575 ;
        RECT 27.245 181.995 28.455 182.745 ;
        RECT 28.625 182.495 28.795 183.405 ;
        RECT 28.965 182.655 29.325 183.235 ;
        RECT 29.505 182.905 29.755 183.405 ;
        RECT 29.925 182.735 30.265 183.765 ;
        RECT 30.925 183.235 31.240 183.675 ;
        RECT 31.575 183.655 31.875 184.205 ;
        RECT 32.085 183.825 32.415 184.545 ;
        RECT 32.605 183.825 33.055 184.375 ;
        RECT 31.575 183.485 32.515 183.655 ;
        RECT 32.345 183.235 32.515 183.485 ;
        RECT 30.925 182.985 31.615 183.235 ;
        RECT 31.845 182.985 32.175 183.235 ;
        RECT 32.345 182.905 32.635 183.235 ;
        RECT 32.345 182.815 32.515 182.905 ;
        RECT 29.580 182.565 30.265 182.735 ;
        RECT 31.125 182.625 32.515 182.815 ;
        RECT 28.625 182.165 28.885 182.495 ;
        RECT 29.095 181.995 29.370 182.475 ;
        RECT 29.580 182.165 29.785 182.565 ;
        RECT 29.955 181.995 30.290 182.395 ;
        RECT 31.125 182.265 31.455 182.625 ;
        RECT 32.805 182.455 33.055 183.825 ;
        RECT 33.225 183.405 33.515 184.545 ;
        RECT 33.685 184.110 39.030 184.545 ;
        RECT 32.085 181.995 32.335 182.455 ;
        RECT 32.505 182.165 33.055 182.455 ;
        RECT 33.225 181.995 33.515 182.795 ;
        RECT 35.270 182.540 35.610 183.370 ;
        RECT 37.090 182.860 37.440 184.110 ;
        RECT 40.125 183.380 40.415 184.545 ;
        RECT 40.585 183.995 40.845 184.375 ;
        RECT 41.015 184.165 41.345 184.545 ;
        RECT 41.685 183.995 41.855 184.375 ;
        RECT 42.025 184.165 42.365 184.545 ;
        RECT 42.535 183.995 42.705 184.375 ;
        RECT 42.940 184.165 43.610 184.545 ;
        RECT 44.255 184.165 44.585 184.545 ;
        RECT 40.585 183.825 41.515 183.995 ;
        RECT 41.685 183.825 42.865 183.995 ;
        RECT 44.755 183.965 44.925 184.375 ;
        RECT 33.685 181.995 39.030 182.540 ;
        RECT 40.125 181.995 40.415 182.720 ;
        RECT 40.585 182.495 40.755 183.825 ;
        RECT 41.345 183.655 41.515 183.825 ;
        RECT 41.345 183.485 42.525 183.655 ;
        RECT 40.925 182.675 41.275 183.215 ;
        RECT 40.585 182.165 40.845 182.495 ;
        RECT 41.015 181.995 41.265 182.495 ;
        RECT 41.445 182.335 41.750 183.315 ;
        RECT 42.355 183.310 42.525 183.485 ;
        RECT 41.925 182.845 42.190 183.185 ;
        RECT 41.925 182.675 42.195 182.845 ;
        RECT 42.695 182.715 42.865 183.825 ;
        RECT 43.175 183.795 44.925 183.965 ;
        RECT 45.185 183.825 45.645 184.375 ;
        RECT 45.835 183.825 46.165 184.545 ;
        RECT 43.175 183.235 43.345 183.795 ;
        RECT 43.780 183.455 44.110 183.625 ;
        RECT 43.035 182.905 43.345 183.235 ;
        RECT 43.515 182.715 43.685 183.235 ;
        RECT 41.925 182.330 42.190 182.675 ;
        RECT 42.695 182.545 43.685 182.715 ;
        RECT 42.920 182.165 43.090 182.545 ;
        RECT 43.360 181.995 43.690 182.375 ;
        RECT 43.860 182.165 44.085 183.455 ;
        RECT 44.430 182.715 44.600 183.795 ;
        RECT 44.770 183.525 44.950 183.545 ;
        RECT 44.770 183.355 44.955 183.525 ;
        RECT 44.770 182.905 44.950 183.355 ;
        RECT 44.430 182.545 44.925 182.715 ;
        RECT 44.255 181.995 44.585 182.375 ;
        RECT 44.755 182.165 44.925 182.545 ;
        RECT 45.185 182.455 45.435 183.825 ;
        RECT 46.365 183.655 46.665 184.205 ;
        RECT 46.835 183.875 47.115 184.545 ;
        RECT 45.725 183.485 46.665 183.655 ;
        RECT 47.520 183.755 48.055 184.375 ;
        RECT 45.725 183.235 45.895 183.485 ;
        RECT 47.035 183.235 47.300 183.595 ;
        RECT 45.605 182.905 45.895 183.235 ;
        RECT 46.065 182.985 46.405 183.235 ;
        RECT 46.625 182.985 47.300 183.235 ;
        RECT 45.725 182.815 45.895 182.905 ;
        RECT 45.725 182.625 47.115 182.815 ;
        RECT 45.185 182.165 45.745 182.455 ;
        RECT 45.915 181.995 46.165 182.455 ;
        RECT 46.785 182.265 47.115 182.625 ;
        RECT 47.520 182.735 47.835 183.755 ;
        RECT 48.225 183.745 48.555 184.545 ;
        RECT 49.040 183.575 49.430 183.750 ;
        RECT 48.005 183.405 49.430 183.575 ;
        RECT 49.940 183.535 50.240 184.375 ;
        RECT 50.435 183.705 50.685 184.545 ;
        RECT 51.275 183.955 52.080 184.375 ;
        RECT 50.855 183.785 52.420 183.955 ;
        RECT 50.855 183.535 51.025 183.785 ;
        RECT 48.005 182.905 48.175 183.405 ;
        RECT 47.520 182.165 48.135 182.735 ;
        RECT 48.425 182.675 48.690 183.235 ;
        RECT 48.860 182.505 49.030 183.405 ;
        RECT 49.940 183.365 51.025 183.535 ;
        RECT 49.200 182.675 49.555 183.235 ;
        RECT 49.785 182.905 50.115 183.195 ;
        RECT 50.285 182.735 50.455 183.365 ;
        RECT 51.195 183.235 51.515 183.615 ;
        RECT 51.705 183.525 52.080 183.615 ;
        RECT 51.685 183.355 52.080 183.525 ;
        RECT 52.250 183.535 52.420 183.785 ;
        RECT 52.590 183.705 52.920 184.545 ;
        RECT 53.090 183.785 53.755 184.375 ;
        RECT 52.250 183.365 53.170 183.535 ;
        RECT 50.625 182.985 50.955 183.195 ;
        RECT 51.135 182.985 51.515 183.235 ;
        RECT 51.705 183.195 52.080 183.355 ;
        RECT 53.000 183.195 53.170 183.365 ;
        RECT 51.705 182.985 52.190 183.195 ;
        RECT 52.380 182.985 52.830 183.195 ;
        RECT 53.000 182.985 53.335 183.195 ;
        RECT 53.505 182.815 53.755 183.785 ;
        RECT 49.945 182.555 50.455 182.735 ;
        RECT 50.860 182.645 52.560 182.815 ;
        RECT 50.860 182.555 51.245 182.645 ;
        RECT 48.305 181.995 48.520 182.505 ;
        RECT 48.750 182.175 49.030 182.505 ;
        RECT 49.210 181.995 49.450 182.505 ;
        RECT 49.945 182.165 50.275 182.555 ;
        RECT 50.445 182.215 51.630 182.385 ;
        RECT 51.890 181.995 52.060 182.465 ;
        RECT 52.230 182.180 52.560 182.645 ;
        RECT 52.730 181.995 52.900 182.815 ;
        RECT 53.070 182.175 53.755 182.815 ;
        RECT 53.930 183.595 54.195 184.365 ;
        RECT 54.365 183.825 54.695 184.545 ;
        RECT 54.885 184.005 55.145 184.365 ;
        RECT 55.315 184.175 55.645 184.545 ;
        RECT 55.815 184.005 56.075 184.365 ;
        RECT 54.885 183.775 56.075 184.005 ;
        RECT 56.645 183.595 56.935 184.365 ;
        RECT 53.930 182.175 54.265 183.595 ;
        RECT 54.440 183.415 56.935 183.595 ;
        RECT 57.145 183.455 59.735 184.545 ;
        RECT 59.995 183.925 60.165 184.355 ;
        RECT 60.335 184.095 60.665 184.545 ;
        RECT 59.995 183.695 60.675 183.925 ;
        RECT 54.440 182.725 54.665 183.415 ;
        RECT 54.865 182.905 55.145 183.235 ;
        RECT 55.325 182.905 55.900 183.235 ;
        RECT 56.080 182.905 56.515 183.235 ;
        RECT 56.695 182.905 56.965 183.235 ;
        RECT 57.145 182.765 58.355 183.285 ;
        RECT 58.525 182.935 59.735 183.455 ;
        RECT 59.965 183.355 60.270 183.525 ;
        RECT 54.440 182.535 56.925 182.725 ;
        RECT 54.445 181.995 55.190 182.365 ;
        RECT 55.755 182.175 56.010 182.535 ;
        RECT 56.190 181.995 56.520 182.365 ;
        RECT 56.700 182.175 56.925 182.535 ;
        RECT 57.145 181.995 59.735 182.765 ;
        RECT 59.970 182.675 60.270 183.355 ;
        RECT 60.440 183.045 60.675 183.695 ;
        RECT 60.865 183.385 61.150 184.330 ;
        RECT 61.330 184.075 62.015 184.545 ;
        RECT 61.325 183.555 62.020 183.865 ;
        RECT 62.195 183.490 62.500 184.275 ;
        RECT 62.685 183.590 62.955 184.545 ;
        RECT 60.865 183.235 61.725 183.385 ;
        RECT 60.865 183.215 62.155 183.235 ;
        RECT 60.440 182.715 60.995 183.045 ;
        RECT 61.165 182.855 62.155 183.215 ;
        RECT 60.440 182.565 60.655 182.715 ;
        RECT 59.915 181.995 60.245 182.500 ;
        RECT 60.415 182.190 60.655 182.565 ;
        RECT 61.165 182.520 61.335 182.855 ;
        RECT 62.325 182.685 62.500 183.490 ;
        RECT 63.125 183.455 65.715 184.545 ;
        RECT 60.935 182.325 61.335 182.520 ;
        RECT 60.935 182.180 61.105 182.325 ;
        RECT 61.695 181.995 62.095 182.490 ;
        RECT 62.265 182.165 62.500 182.685 ;
        RECT 63.125 182.765 64.335 183.285 ;
        RECT 64.505 182.935 65.715 183.455 ;
        RECT 65.885 183.380 66.175 184.545 ;
        RECT 66.345 183.455 69.855 184.545 ;
        RECT 66.345 182.765 67.995 183.285 ;
        RECT 68.165 182.935 69.855 183.455 ;
        RECT 70.495 183.485 70.825 184.335 ;
        RECT 62.685 181.995 62.955 182.630 ;
        RECT 63.125 181.995 65.715 182.765 ;
        RECT 65.885 181.995 66.175 182.720 ;
        RECT 66.345 181.995 69.855 182.765 ;
        RECT 70.495 182.720 70.685 183.485 ;
        RECT 70.995 183.405 71.245 184.545 ;
        RECT 71.435 183.905 71.685 184.325 ;
        RECT 71.915 184.075 72.245 184.545 ;
        RECT 72.475 183.905 72.725 184.325 ;
        RECT 71.435 183.735 72.725 183.905 ;
        RECT 72.905 183.905 73.235 184.335 ;
        RECT 72.905 183.735 73.360 183.905 ;
        RECT 71.425 183.235 71.640 183.565 ;
        RECT 70.855 182.905 71.165 183.235 ;
        RECT 71.335 182.905 71.640 183.235 ;
        RECT 71.815 182.905 72.100 183.565 ;
        RECT 72.295 182.905 72.560 183.565 ;
        RECT 72.775 182.905 73.020 183.565 ;
        RECT 70.995 182.735 71.165 182.905 ;
        RECT 73.190 182.735 73.360 183.735 ;
        RECT 74.625 183.405 74.885 184.545 ;
        RECT 75.125 184.035 76.740 184.365 ;
        RECT 75.135 183.235 75.305 183.795 ;
        RECT 75.565 183.695 76.740 183.865 ;
        RECT 76.910 183.745 77.190 184.545 ;
        RECT 75.565 183.405 75.895 183.695 ;
        RECT 76.570 183.575 76.740 183.695 ;
        RECT 76.065 183.235 76.310 183.525 ;
        RECT 76.570 183.405 77.230 183.575 ;
        RECT 77.400 183.405 77.675 184.375 ;
        RECT 77.845 184.165 79.105 184.375 ;
        RECT 77.845 183.745 78.105 184.165 ;
        RECT 77.060 183.235 77.230 183.405 ;
        RECT 74.630 182.985 74.965 183.235 ;
        RECT 75.135 182.905 75.850 183.235 ;
        RECT 76.065 182.905 76.890 183.235 ;
        RECT 77.060 182.905 77.335 183.235 ;
        RECT 75.135 182.815 75.385 182.905 ;
        RECT 70.495 182.210 70.825 182.720 ;
        RECT 70.995 182.565 73.360 182.735 ;
        RECT 70.995 181.995 71.325 182.395 ;
        RECT 72.375 182.225 72.705 182.565 ;
        RECT 72.875 181.995 73.205 182.395 ;
        RECT 74.625 181.995 74.885 182.815 ;
        RECT 75.055 182.395 75.385 182.815 ;
        RECT 77.060 182.735 77.230 182.905 ;
        RECT 75.565 182.565 77.230 182.735 ;
        RECT 77.505 182.670 77.675 183.405 ;
        RECT 78.275 183.695 78.625 183.995 ;
        RECT 78.855 183.865 79.105 184.165 ;
        RECT 79.315 184.045 79.565 184.545 ;
        RECT 79.775 183.865 79.945 184.375 ;
        RECT 78.855 183.695 79.945 183.865 ;
        RECT 77.845 182.905 78.105 183.235 ;
        RECT 75.565 182.165 75.825 182.565 ;
        RECT 75.995 181.995 76.325 182.395 ;
        RECT 76.495 182.215 76.665 182.565 ;
        RECT 76.835 181.995 77.210 182.395 ;
        RECT 77.400 182.325 77.675 182.670 ;
        RECT 78.275 182.715 78.445 183.695 ;
        RECT 79.775 183.655 79.945 183.695 ;
        RECT 78.615 183.335 79.015 183.525 ;
        RECT 80.115 183.405 80.455 184.545 ;
        RECT 81.065 183.575 81.335 184.345 ;
        RECT 81.505 183.765 81.835 184.545 ;
        RECT 82.040 183.940 82.225 184.345 ;
        RECT 82.395 184.120 82.730 184.545 ;
        RECT 82.040 183.765 82.705 183.940 ;
        RECT 81.065 183.405 82.195 183.575 ;
        RECT 78.615 182.905 78.785 183.335 ;
        RECT 78.990 182.985 79.355 183.165 ;
        RECT 78.275 182.545 78.925 182.715 ;
        RECT 77.855 181.995 78.185 182.375 ;
        RECT 78.675 182.205 78.925 182.545 ;
        RECT 79.165 182.675 79.355 182.985 ;
        RECT 79.565 182.905 79.925 183.235 ;
        RECT 80.095 182.925 80.510 183.235 ;
        RECT 79.165 182.255 79.465 182.675 ;
        RECT 79.725 182.325 79.925 182.905 ;
        RECT 80.115 181.995 80.455 182.715 ;
        RECT 81.065 182.495 81.235 183.405 ;
        RECT 81.405 182.655 81.765 183.235 ;
        RECT 81.945 182.905 82.195 183.405 ;
        RECT 82.365 182.735 82.705 183.765 ;
        RECT 82.985 183.615 83.165 184.375 ;
        RECT 83.345 183.785 83.675 184.545 ;
        RECT 82.985 183.445 83.660 183.615 ;
        RECT 83.845 183.470 84.115 184.375 ;
        RECT 83.490 183.300 83.660 183.445 ;
        RECT 82.925 182.895 83.265 183.265 ;
        RECT 83.490 182.970 83.765 183.300 ;
        RECT 82.020 182.565 82.705 182.735 ;
        RECT 83.490 182.715 83.660 182.970 ;
        RECT 81.065 182.165 81.325 182.495 ;
        RECT 81.535 181.995 81.810 182.475 ;
        RECT 82.020 182.165 82.225 182.565 ;
        RECT 82.995 182.545 83.660 182.715 ;
        RECT 83.935 182.670 84.115 183.470 ;
        RECT 82.395 181.995 82.730 182.395 ;
        RECT 82.995 182.165 83.165 182.545 ;
        RECT 83.345 181.995 83.675 182.375 ;
        RECT 83.855 182.165 84.115 182.670 ;
        RECT 84.300 182.175 84.580 184.365 ;
        RECT 84.770 183.405 85.055 184.545 ;
        RECT 85.320 183.895 85.490 184.365 ;
        RECT 85.665 184.065 85.995 184.545 ;
        RECT 86.165 183.895 86.345 184.365 ;
        RECT 85.320 183.695 86.345 183.895 ;
        RECT 84.780 182.725 85.040 183.235 ;
        RECT 85.250 182.905 85.510 183.525 ;
        RECT 85.705 182.905 86.130 183.525 ;
        RECT 86.515 183.255 86.845 184.365 ;
        RECT 87.015 184.135 87.365 184.545 ;
        RECT 87.535 183.955 87.775 184.345 ;
        RECT 86.300 182.955 86.845 183.255 ;
        RECT 87.025 183.755 87.775 183.955 ;
        RECT 87.025 183.075 87.365 183.755 ;
        RECT 86.300 182.725 86.520 182.955 ;
        RECT 84.780 182.535 86.520 182.725 ;
        RECT 84.780 181.995 85.510 182.365 ;
        RECT 86.090 182.175 86.520 182.535 ;
        RECT 86.690 181.995 86.935 182.775 ;
        RECT 87.135 182.175 87.365 183.075 ;
        RECT 87.545 182.235 87.775 183.575 ;
        RECT 87.965 182.165 88.715 184.375 ;
        RECT 88.965 183.615 89.145 184.375 ;
        RECT 89.325 183.785 89.655 184.545 ;
        RECT 88.965 183.445 89.640 183.615 ;
        RECT 89.825 183.470 90.095 184.375 ;
        RECT 89.470 183.300 89.640 183.445 ;
        RECT 88.905 182.895 89.245 183.265 ;
        RECT 89.470 182.970 89.745 183.300 ;
        RECT 89.470 182.715 89.640 182.970 ;
        RECT 88.975 182.545 89.640 182.715 ;
        RECT 89.915 182.670 90.095 183.470 ;
        RECT 90.265 183.405 90.525 184.545 ;
        RECT 90.695 183.395 91.025 184.375 ;
        RECT 91.195 183.405 91.475 184.545 ;
        RECT 90.285 182.985 90.620 183.235 ;
        RECT 90.790 182.795 90.960 183.395 ;
        RECT 91.645 183.380 91.935 184.545 ;
        RECT 92.565 183.695 92.825 184.375 ;
        RECT 92.995 183.765 93.245 184.545 ;
        RECT 93.495 183.995 93.745 184.375 ;
        RECT 93.915 184.165 94.270 184.545 ;
        RECT 95.275 184.155 95.610 184.375 ;
        RECT 94.875 183.995 95.105 184.035 ;
        RECT 93.495 183.795 95.105 183.995 ;
        RECT 93.495 183.785 94.330 183.795 ;
        RECT 94.920 183.705 95.105 183.795 ;
        RECT 91.130 182.965 91.465 183.235 ;
        RECT 88.975 182.165 89.145 182.545 ;
        RECT 89.325 181.995 89.655 182.375 ;
        RECT 89.835 182.165 90.095 182.670 ;
        RECT 90.265 182.165 90.960 182.795 ;
        RECT 91.165 181.995 91.475 182.795 ;
        RECT 91.645 181.995 91.935 182.720 ;
        RECT 92.565 182.505 92.735 183.695 ;
        RECT 94.435 183.595 94.765 183.625 ;
        RECT 92.965 183.535 94.765 183.595 ;
        RECT 95.355 183.535 95.610 184.155 ;
        RECT 92.905 183.425 95.610 183.535 ;
        RECT 92.905 183.390 93.105 183.425 ;
        RECT 92.905 182.815 93.075 183.390 ;
        RECT 94.435 183.365 95.610 183.425 ;
        RECT 96.705 183.435 96.965 184.375 ;
        RECT 97.135 184.145 97.465 184.545 ;
        RECT 98.610 184.280 98.865 184.375 ;
        RECT 97.725 184.110 98.865 184.280 ;
        RECT 99.035 184.165 99.365 184.335 ;
        RECT 97.725 183.885 97.895 184.110 ;
        RECT 97.135 183.715 97.895 183.885 ;
        RECT 98.610 183.975 98.865 184.110 ;
        RECT 93.305 182.950 93.715 183.255 ;
        RECT 93.885 182.985 94.215 183.195 ;
        RECT 92.905 182.695 93.175 182.815 ;
        RECT 92.905 182.650 93.750 182.695 ;
        RECT 92.995 182.525 93.750 182.650 ;
        RECT 94.005 182.585 94.215 182.985 ;
        RECT 94.460 182.985 94.935 183.195 ;
        RECT 95.125 182.985 95.615 183.185 ;
        RECT 94.460 182.585 94.680 182.985 ;
        RECT 92.565 182.495 92.795 182.505 ;
        RECT 92.565 182.165 92.825 182.495 ;
        RECT 93.580 182.375 93.750 182.525 ;
        RECT 92.995 181.995 93.325 182.355 ;
        RECT 93.580 182.165 94.880 182.375 ;
        RECT 95.155 181.995 95.610 182.760 ;
        RECT 96.705 182.720 96.880 183.435 ;
        RECT 97.135 183.235 97.305 183.715 ;
        RECT 98.160 183.625 98.330 183.815 ;
        RECT 98.610 183.805 99.020 183.975 ;
        RECT 97.050 182.905 97.305 183.235 ;
        RECT 97.530 182.905 97.860 183.525 ;
        RECT 98.160 183.455 98.680 183.625 ;
        RECT 98.030 182.905 98.320 183.285 ;
        RECT 98.510 182.735 98.680 183.455 ;
        RECT 96.705 182.165 96.965 182.720 ;
        RECT 97.800 182.565 98.680 182.735 ;
        RECT 98.850 182.780 99.020 183.805 ;
        RECT 99.195 183.915 99.365 184.165 ;
        RECT 99.535 184.085 99.785 184.545 ;
        RECT 99.955 183.915 100.135 184.375 ;
        RECT 99.195 183.745 100.135 183.915 ;
        RECT 99.220 183.265 99.700 183.565 ;
        RECT 98.850 182.610 99.200 182.780 ;
        RECT 99.440 182.675 99.700 183.265 ;
        RECT 99.900 182.675 100.160 183.565 ;
        RECT 101.305 183.405 101.645 184.375 ;
        RECT 101.815 183.405 101.985 184.545 ;
        RECT 102.255 183.745 102.505 184.545 ;
        RECT 103.150 183.575 103.480 184.375 ;
        RECT 103.780 183.745 104.110 184.545 ;
        RECT 104.280 183.575 104.610 184.375 ;
        RECT 104.995 183.735 105.290 184.545 ;
        RECT 102.175 183.405 104.610 183.575 ;
        RECT 101.305 182.795 101.480 183.405 ;
        RECT 102.175 183.155 102.345 183.405 ;
        RECT 101.650 182.985 102.345 183.155 ;
        RECT 102.520 182.985 102.940 183.185 ;
        RECT 103.110 182.985 103.440 183.185 ;
        RECT 103.610 182.985 103.940 183.185 ;
        RECT 97.135 181.995 97.565 182.440 ;
        RECT 97.800 182.165 97.970 182.565 ;
        RECT 98.140 181.995 98.860 182.395 ;
        RECT 99.030 182.165 99.200 182.610 ;
        RECT 99.775 181.995 100.175 182.505 ;
        RECT 101.305 182.165 101.645 182.795 ;
        RECT 101.815 181.995 102.065 182.795 ;
        RECT 102.255 182.645 103.480 182.815 ;
        RECT 102.255 182.165 102.585 182.645 ;
        RECT 102.755 181.995 102.980 182.455 ;
        RECT 103.150 182.165 103.480 182.645 ;
        RECT 104.110 182.775 104.280 183.405 ;
        RECT 105.470 183.235 105.715 184.375 ;
        RECT 105.890 183.735 106.150 184.545 ;
        RECT 106.750 184.540 113.025 184.545 ;
        RECT 106.330 183.235 106.580 184.370 ;
        RECT 106.750 183.745 107.010 184.540 ;
        RECT 107.180 183.645 107.440 184.370 ;
        RECT 107.610 183.815 107.870 184.540 ;
        RECT 108.040 183.645 108.300 184.370 ;
        RECT 108.470 183.815 108.730 184.540 ;
        RECT 108.900 183.645 109.160 184.370 ;
        RECT 109.330 183.815 109.590 184.540 ;
        RECT 109.760 183.645 110.020 184.370 ;
        RECT 110.190 183.815 110.435 184.540 ;
        RECT 110.605 183.645 110.865 184.370 ;
        RECT 111.050 183.815 111.295 184.540 ;
        RECT 111.465 183.645 111.725 184.370 ;
        RECT 111.910 183.815 112.155 184.540 ;
        RECT 112.325 183.645 112.585 184.370 ;
        RECT 112.770 183.815 113.025 184.540 ;
        RECT 107.180 183.630 112.585 183.645 ;
        RECT 113.195 183.630 113.485 184.370 ;
        RECT 113.655 183.800 113.925 184.545 ;
        RECT 114.245 183.845 114.465 184.375 ;
        RECT 114.635 184.035 114.965 184.545 ;
        RECT 115.135 183.845 115.360 184.375 ;
        RECT 107.180 183.405 113.925 183.630 ;
        RECT 114.245 183.580 115.360 183.845 ;
        RECT 115.530 183.830 115.845 184.375 ;
        RECT 116.035 184.130 116.365 184.545 ;
        RECT 115.530 183.600 116.365 183.830 ;
        RECT 104.465 182.985 104.815 183.235 ;
        RECT 104.110 182.165 104.610 182.775 ;
        RECT 104.985 182.675 105.300 183.235 ;
        RECT 105.470 182.985 112.590 183.235 ;
        RECT 104.985 181.995 105.290 182.505 ;
        RECT 105.470 182.175 105.720 182.985 ;
        RECT 105.890 181.995 106.150 182.520 ;
        RECT 106.330 182.175 106.580 182.985 ;
        RECT 112.760 182.815 113.925 183.405 ;
        RECT 107.180 182.645 113.925 182.815 ;
        RECT 114.195 182.660 114.510 183.235 ;
        RECT 106.750 181.995 107.010 182.555 ;
        RECT 107.180 182.190 107.440 182.645 ;
        RECT 107.610 181.995 107.870 182.475 ;
        RECT 108.040 182.190 108.300 182.645 ;
        RECT 108.470 181.995 108.730 182.475 ;
        RECT 108.900 182.190 109.160 182.645 ;
        RECT 109.330 181.995 109.575 182.475 ;
        RECT 109.745 182.190 110.020 182.645 ;
        RECT 110.190 181.995 110.435 182.475 ;
        RECT 110.605 182.190 110.865 182.645 ;
        RECT 111.045 181.995 111.295 182.475 ;
        RECT 111.465 182.190 111.725 182.645 ;
        RECT 111.905 181.995 112.155 182.475 ;
        RECT 112.325 182.190 112.585 182.645 ;
        RECT 112.765 181.995 113.025 182.475 ;
        RECT 113.195 182.190 113.455 182.645 ;
        RECT 113.625 181.995 113.925 182.475 ;
        RECT 114.185 181.995 114.515 182.475 ;
        RECT 114.700 182.275 115.080 183.235 ;
        RECT 115.530 182.905 115.855 183.320 ;
        RECT 116.025 182.905 116.365 183.600 ;
        RECT 116.025 182.735 116.195 182.905 ;
        RECT 116.535 182.735 116.765 184.375 ;
        RECT 116.935 183.575 117.225 184.545 ;
        RECT 117.405 183.380 117.695 184.545 ;
        RECT 118.875 183.575 119.045 184.375 ;
        RECT 119.335 183.915 119.585 184.335 ;
        RECT 119.775 184.085 120.105 184.545 ;
        RECT 120.315 183.915 120.565 184.335 ;
        RECT 119.275 183.745 120.565 183.915 ;
        RECT 120.735 183.745 120.985 184.545 ;
        RECT 121.155 183.915 121.325 184.375 ;
        RECT 121.535 184.085 121.785 184.545 ;
        RECT 121.155 183.745 121.830 183.915 ;
        RECT 122.095 183.800 122.365 184.545 ;
        RECT 122.995 184.540 129.270 184.545 ;
        RECT 118.875 183.405 121.365 183.575 ;
        RECT 115.455 182.565 116.195 182.735 ;
        RECT 115.455 182.165 115.645 182.565 ;
        RECT 116.365 182.545 116.765 182.735 ;
        RECT 115.865 181.995 116.195 182.355 ;
        RECT 116.365 182.165 116.555 182.545 ;
        RECT 116.725 181.995 117.055 182.375 ;
        RECT 117.405 181.995 117.695 182.720 ;
        RECT 118.830 182.665 119.025 183.235 ;
        RECT 118.785 181.995 119.045 182.475 ;
        RECT 119.215 182.415 119.385 183.405 ;
        RECT 119.565 182.780 119.735 183.235 ;
        RECT 120.125 183.155 120.295 183.170 ;
        RECT 119.965 182.985 120.295 183.155 ;
        RECT 119.565 182.610 119.955 182.780 ;
        RECT 119.215 182.245 119.545 182.415 ;
        RECT 119.745 182.325 119.955 182.610 ;
        RECT 120.125 182.775 120.295 182.985 ;
        RECT 120.525 182.905 120.855 183.235 ;
        RECT 121.195 183.155 121.365 183.405 ;
        RECT 121.035 182.985 121.365 183.155 ;
        RECT 120.125 182.605 120.390 182.775 ;
        RECT 120.650 182.670 120.855 182.905 ;
        RECT 121.575 182.795 121.830 183.745 ;
        RECT 122.535 183.630 122.825 184.370 ;
        RECT 122.995 183.815 123.250 184.540 ;
        RECT 123.435 183.645 123.695 184.370 ;
        RECT 123.865 183.815 124.110 184.540 ;
        RECT 124.295 183.645 124.555 184.370 ;
        RECT 124.725 183.815 124.970 184.540 ;
        RECT 125.155 183.645 125.415 184.370 ;
        RECT 125.585 183.815 125.830 184.540 ;
        RECT 126.000 183.645 126.260 184.370 ;
        RECT 126.430 183.815 126.690 184.540 ;
        RECT 126.860 183.645 127.120 184.370 ;
        RECT 127.290 183.815 127.550 184.540 ;
        RECT 127.720 183.645 127.980 184.370 ;
        RECT 128.150 183.815 128.410 184.540 ;
        RECT 128.580 183.645 128.840 184.370 ;
        RECT 129.010 183.745 129.270 184.540 ;
        RECT 123.435 183.630 128.840 183.645 ;
        RECT 120.220 182.505 120.390 182.605 ;
        RECT 121.155 182.625 121.830 182.795 ;
        RECT 122.095 183.405 128.840 183.630 ;
        RECT 122.095 182.815 123.260 183.405 ;
        RECT 129.440 183.235 129.690 184.370 ;
        RECT 129.870 183.735 130.130 184.545 ;
        RECT 130.305 183.235 130.550 184.375 ;
        RECT 130.730 183.735 131.025 184.545 ;
        RECT 131.260 183.705 131.465 184.545 ;
        RECT 131.675 184.205 132.765 184.375 ;
        RECT 131.675 183.695 131.925 184.205 ;
        RECT 132.515 184.035 132.765 184.205 ;
        RECT 132.935 184.035 133.185 184.545 ;
        RECT 132.095 183.865 132.345 184.035 ;
        RECT 133.355 183.875 133.645 184.375 ;
        RECT 133.815 184.045 134.545 184.545 ;
        RECT 135.135 184.045 135.385 184.545 ;
        RECT 134.715 183.875 134.965 184.035 ;
        RECT 135.555 183.875 135.805 184.375 ;
        RECT 133.355 183.865 133.735 183.875 ;
        RECT 132.095 183.695 133.735 183.865 ;
        RECT 131.205 183.355 133.015 183.525 ;
        RECT 123.430 182.985 130.550 183.235 ;
        RECT 122.095 182.645 128.840 182.815 ;
        RECT 120.220 182.335 120.395 182.505 ;
        RECT 120.735 182.375 120.905 182.455 ;
        RECT 120.220 182.310 120.390 182.335 ;
        RECT 119.215 182.165 119.460 182.245 ;
        RECT 120.635 181.995 120.965 182.375 ;
        RECT 121.155 182.165 121.325 182.625 ;
        RECT 121.575 181.995 121.830 182.455 ;
        RECT 122.095 181.995 122.395 182.475 ;
        RECT 122.565 182.190 122.825 182.645 ;
        RECT 122.995 181.995 123.255 182.475 ;
        RECT 123.435 182.190 123.695 182.645 ;
        RECT 123.865 181.995 124.115 182.475 ;
        RECT 124.295 182.190 124.555 182.645 ;
        RECT 124.725 181.995 124.975 182.475 ;
        RECT 125.155 182.190 125.415 182.645 ;
        RECT 125.585 181.995 125.830 182.475 ;
        RECT 126.000 182.190 126.275 182.645 ;
        RECT 126.445 181.995 126.690 182.475 ;
        RECT 126.860 182.190 127.120 182.645 ;
        RECT 127.290 181.995 127.550 182.475 ;
        RECT 127.720 182.190 127.980 182.645 ;
        RECT 128.150 181.995 128.410 182.475 ;
        RECT 128.580 182.190 128.840 182.645 ;
        RECT 129.010 181.995 129.270 182.555 ;
        RECT 129.440 182.175 129.690 182.985 ;
        RECT 129.870 181.995 130.130 182.520 ;
        RECT 130.300 182.175 130.550 182.985 ;
        RECT 130.720 182.675 131.035 183.235 ;
        RECT 131.205 182.985 131.695 183.355 ;
        RECT 132.685 183.185 133.015 183.355 ;
        RECT 131.925 182.985 132.465 183.185 ;
        RECT 132.645 183.015 133.015 183.185 ;
        RECT 132.685 182.985 133.015 183.015 ;
        RECT 133.185 183.325 133.735 183.695 ;
        RECT 134.075 183.695 135.805 183.875 ;
        RECT 135.975 183.705 136.225 184.545 ;
        RECT 136.395 183.865 136.645 184.375 ;
        RECT 136.815 184.075 137.065 184.545 ;
        RECT 137.235 183.865 137.485 184.375 ;
        RECT 136.395 183.695 137.485 183.865 ;
        RECT 137.655 183.735 137.905 184.545 ;
        RECT 133.185 182.985 133.565 183.325 ;
        RECT 134.075 183.155 134.265 183.695 ;
        RECT 137.235 183.565 137.485 183.695 ;
        RECT 133.735 182.985 134.265 183.155 ;
        RECT 134.435 183.355 136.085 183.525 ;
        RECT 134.435 182.985 134.765 183.355 ;
        RECT 134.935 182.985 135.555 183.185 ;
        RECT 135.725 182.985 136.085 183.355 ;
        RECT 136.285 183.155 136.575 183.525 ;
        RECT 137.235 183.325 138.030 183.565 ;
        RECT 136.285 182.985 137.555 183.155 ;
        RECT 131.215 182.645 133.145 182.815 ;
        RECT 131.215 182.635 132.385 182.645 ;
        RECT 130.730 181.995 131.035 182.505 ;
        RECT 131.215 182.165 131.545 182.635 ;
        RECT 131.715 181.995 131.885 182.465 ;
        RECT 132.055 182.165 132.385 182.635 ;
        RECT 132.555 181.995 132.725 182.465 ;
        RECT 132.895 182.385 133.145 182.645 ;
        RECT 133.315 182.725 133.565 182.985 ;
        RECT 134.075 182.815 134.265 182.985 ;
        RECT 137.725 182.815 138.030 183.325 ;
        RECT 138.565 183.455 139.775 184.545 ;
        RECT 138.565 182.915 139.085 183.455 ;
        RECT 133.315 182.555 133.645 182.725 ;
        RECT 134.075 182.635 135.425 182.815 ;
        RECT 135.095 182.555 135.425 182.635 ;
        RECT 132.895 182.165 134.065 182.385 ;
        RECT 134.335 181.995 134.505 182.465 ;
        RECT 135.595 182.385 135.845 182.805 ;
        RECT 134.675 182.215 135.845 182.385 ;
        RECT 136.015 181.995 136.185 182.805 ;
        RECT 136.355 182.635 138.030 182.815 ;
        RECT 139.255 182.745 139.775 183.285 ;
        RECT 136.355 182.185 136.685 182.635 ;
        RECT 136.855 181.995 137.025 182.465 ;
        RECT 137.195 182.185 137.525 182.635 ;
        RECT 137.695 181.995 137.865 182.465 ;
        RECT 138.565 181.995 139.775 182.745 ;
        RECT 27.160 181.825 139.860 181.995 ;
        RECT 27.245 181.075 28.455 181.825 ;
        RECT 27.245 180.535 27.765 181.075 ;
        RECT 28.630 180.985 28.890 181.825 ;
        RECT 29.065 181.080 29.320 181.655 ;
        RECT 29.490 181.445 29.820 181.825 ;
        RECT 30.035 181.275 30.205 181.655 ;
        RECT 29.490 181.105 30.205 181.275 ;
        RECT 31.385 181.150 31.645 181.655 ;
        RECT 31.825 181.445 32.155 181.825 ;
        RECT 32.335 181.275 32.505 181.655 ;
        RECT 32.765 181.280 38.110 181.825 ;
        RECT 27.935 180.365 28.455 180.905 ;
        RECT 27.245 179.275 28.455 180.365 ;
        RECT 28.630 179.275 28.890 180.425 ;
        RECT 29.065 180.350 29.235 181.080 ;
        RECT 29.490 180.915 29.660 181.105 ;
        RECT 29.405 180.585 29.660 180.915 ;
        RECT 29.490 180.375 29.660 180.585 ;
        RECT 29.940 180.555 30.295 180.925 ;
        RECT 29.065 179.445 29.320 180.350 ;
        RECT 29.490 180.205 30.205 180.375 ;
        RECT 29.490 179.275 29.820 180.035 ;
        RECT 30.035 179.445 30.205 180.205 ;
        RECT 31.385 180.350 31.555 181.150 ;
        RECT 31.840 181.105 32.505 181.275 ;
        RECT 31.840 180.850 32.010 181.105 ;
        RECT 31.725 180.520 32.010 180.850 ;
        RECT 32.245 180.555 32.575 180.925 ;
        RECT 31.840 180.375 32.010 180.520 ;
        RECT 34.350 180.450 34.690 181.280 ;
        RECT 38.285 181.055 41.795 181.825 ;
        RECT 31.385 179.445 31.655 180.350 ;
        RECT 31.840 180.205 32.505 180.375 ;
        RECT 31.825 179.275 32.155 180.035 ;
        RECT 32.335 179.445 32.505 180.205 ;
        RECT 36.170 179.710 36.520 180.960 ;
        RECT 38.285 180.535 39.935 181.055 ;
        RECT 42.430 180.985 42.690 181.825 ;
        RECT 42.865 181.080 43.120 181.655 ;
        RECT 43.290 181.445 43.620 181.825 ;
        RECT 43.835 181.275 44.005 181.655 ;
        RECT 43.290 181.105 44.005 181.275 ;
        RECT 44.315 181.285 44.540 181.645 ;
        RECT 44.720 181.455 45.050 181.825 ;
        RECT 45.230 181.285 45.485 181.645 ;
        RECT 46.050 181.455 46.795 181.825 ;
        RECT 40.105 180.365 41.795 180.885 ;
        RECT 32.765 179.275 38.110 179.710 ;
        RECT 38.285 179.275 41.795 180.365 ;
        RECT 42.430 179.275 42.690 180.425 ;
        RECT 42.865 180.350 43.035 181.080 ;
        RECT 43.290 180.915 43.460 181.105 ;
        RECT 44.315 181.095 46.800 181.285 ;
        RECT 43.205 180.585 43.460 180.915 ;
        RECT 43.290 180.375 43.460 180.585 ;
        RECT 43.740 180.555 44.095 180.925 ;
        RECT 44.275 180.585 44.545 180.915 ;
        RECT 44.725 180.585 45.160 180.915 ;
        RECT 45.340 180.585 45.915 180.915 ;
        RECT 46.095 180.585 46.375 180.915 ;
        RECT 46.575 180.405 46.800 181.095 ;
        RECT 42.865 179.445 43.120 180.350 ;
        RECT 43.290 180.205 44.005 180.375 ;
        RECT 43.290 179.275 43.620 180.035 ;
        RECT 43.835 179.445 44.005 180.205 ;
        RECT 44.305 180.225 46.800 180.405 ;
        RECT 46.975 180.225 47.310 181.645 ;
        RECT 44.305 179.455 44.595 180.225 ;
        RECT 45.165 179.815 46.355 180.045 ;
        RECT 45.165 179.455 45.425 179.815 ;
        RECT 45.595 179.275 45.925 179.645 ;
        RECT 46.095 179.455 46.355 179.815 ;
        RECT 46.545 179.275 46.875 179.995 ;
        RECT 47.045 179.455 47.310 180.225 ;
        RECT 47.495 179.455 47.755 181.645 ;
        RECT 48.015 181.455 48.685 181.825 ;
        RECT 48.865 181.275 49.175 181.645 ;
        RECT 47.945 181.075 49.175 181.275 ;
        RECT 47.945 180.405 48.235 181.075 ;
        RECT 49.355 180.895 49.585 181.535 ;
        RECT 49.765 181.095 50.055 181.825 ;
        RECT 50.335 181.275 50.505 181.655 ;
        RECT 50.720 181.445 51.050 181.825 ;
        RECT 50.335 181.105 51.050 181.275 ;
        RECT 48.415 180.585 48.880 180.895 ;
        RECT 49.060 180.585 49.585 180.895 ;
        RECT 49.765 180.585 50.065 180.915 ;
        RECT 50.245 180.555 50.600 180.925 ;
        RECT 50.880 180.915 51.050 181.105 ;
        RECT 51.220 181.080 51.475 181.655 ;
        RECT 50.880 180.585 51.135 180.915 ;
        RECT 47.945 180.185 48.715 180.405 ;
        RECT 47.925 179.275 48.265 180.005 ;
        RECT 48.445 179.455 48.715 180.185 ;
        RECT 48.895 180.165 50.055 180.405 ;
        RECT 50.880 180.375 51.050 180.585 ;
        RECT 48.895 179.455 49.125 180.165 ;
        RECT 49.295 179.275 49.625 179.985 ;
        RECT 49.795 179.455 50.055 180.165 ;
        RECT 50.335 180.205 51.050 180.375 ;
        RECT 51.305 180.350 51.475 181.080 ;
        RECT 51.650 180.985 51.910 181.825 ;
        RECT 53.005 181.100 53.295 181.825 ;
        RECT 53.475 181.105 53.805 181.825 ;
        RECT 54.350 181.425 55.965 181.595 ;
        RECT 56.135 181.425 56.465 181.825 ;
        RECT 55.795 181.255 55.965 181.425 ;
        RECT 56.635 181.350 56.970 181.610 ;
        RECT 53.530 180.585 53.880 180.915 ;
        RECT 54.190 180.585 54.610 181.250 ;
        RECT 54.780 180.805 55.070 181.245 ;
        RECT 55.260 180.805 55.530 181.245 ;
        RECT 55.795 181.085 56.355 181.255 ;
        RECT 56.185 180.915 56.355 181.085 ;
        RECT 55.740 180.805 55.990 180.915 ;
        RECT 54.780 180.635 55.075 180.805 ;
        RECT 55.260 180.635 55.535 180.805 ;
        RECT 55.740 180.635 55.995 180.805 ;
        RECT 54.780 180.585 55.070 180.635 ;
        RECT 55.260 180.585 55.530 180.635 ;
        RECT 55.740 180.585 55.990 180.635 ;
        RECT 56.185 180.585 56.490 180.915 ;
        RECT 53.530 180.465 53.735 180.585 ;
        RECT 50.335 179.445 50.505 180.205 ;
        RECT 50.720 179.275 51.050 180.035 ;
        RECT 51.220 179.445 51.475 180.350 ;
        RECT 51.650 179.275 51.910 180.425 ;
        RECT 53.005 179.275 53.295 180.440 ;
        RECT 53.525 180.295 53.735 180.465 ;
        RECT 56.185 180.415 56.355 180.585 ;
        RECT 53.985 180.245 56.355 180.415 ;
        RECT 53.555 179.615 53.725 180.115 ;
        RECT 53.985 179.785 54.155 180.245 ;
        RECT 54.385 179.865 55.810 180.035 ;
        RECT 54.385 179.615 54.715 179.865 ;
        RECT 53.555 179.445 54.715 179.615 ;
        RECT 54.940 179.275 55.270 179.695 ;
        RECT 55.525 179.445 55.810 179.865 ;
        RECT 56.055 179.275 56.385 180.075 ;
        RECT 56.715 179.995 56.970 181.350 ;
        RECT 57.170 181.070 57.405 181.400 ;
        RECT 57.575 181.085 57.905 181.825 ;
        RECT 58.140 181.445 59.335 181.655 ;
        RECT 57.170 180.415 57.340 181.070 ;
        RECT 58.140 181.005 58.415 181.445 ;
        RECT 58.585 181.105 58.915 181.275 ;
        RECT 58.590 181.005 58.915 181.105 ;
        RECT 59.085 181.215 59.335 181.445 ;
        RECT 59.505 181.385 59.675 181.825 ;
        RECT 59.845 181.215 60.195 181.655 ;
        RECT 59.085 181.005 60.195 181.215 ;
        RECT 60.365 181.325 60.625 181.655 ;
        RECT 60.795 181.465 61.125 181.825 ;
        RECT 61.380 181.445 62.680 181.655 ;
        RECT 60.365 181.315 60.595 181.325 ;
        RECT 57.515 180.585 57.860 180.915 ;
        RECT 58.090 180.415 58.420 180.835 ;
        RECT 57.170 180.245 58.420 180.415 ;
        RECT 57.170 180.050 57.470 180.245 ;
        RECT 58.590 180.075 58.870 181.005 ;
        RECT 59.050 180.635 60.195 180.835 ;
        RECT 59.050 180.255 59.240 180.635 ;
        RECT 59.505 180.415 59.675 180.465 ;
        RECT 59.420 180.075 59.695 180.415 ;
        RECT 56.635 179.485 56.970 179.995 ;
        RECT 57.640 179.275 57.895 180.075 ;
        RECT 58.095 179.905 59.695 180.075 ;
        RECT 58.095 179.445 58.425 179.905 ;
        RECT 58.595 179.275 59.170 179.735 ;
        RECT 59.340 179.445 59.695 179.905 ;
        RECT 59.865 179.275 60.195 180.415 ;
        RECT 60.365 180.125 60.535 181.315 ;
        RECT 61.380 181.295 61.550 181.445 ;
        RECT 60.795 181.170 61.550 181.295 ;
        RECT 60.705 181.125 61.550 181.170 ;
        RECT 60.705 181.005 60.975 181.125 ;
        RECT 60.705 180.430 60.875 181.005 ;
        RECT 61.105 180.565 61.515 180.870 ;
        RECT 61.805 180.835 62.015 181.235 ;
        RECT 61.685 180.625 62.015 180.835 ;
        RECT 62.260 180.835 62.480 181.235 ;
        RECT 62.955 181.060 63.410 181.825 ;
        RECT 63.585 181.075 64.795 181.825 ;
        RECT 65.055 181.275 65.225 181.655 ;
        RECT 65.440 181.445 65.770 181.825 ;
        RECT 65.055 181.105 65.770 181.275 ;
        RECT 62.260 180.625 62.735 180.835 ;
        RECT 62.925 180.635 63.415 180.835 ;
        RECT 63.585 180.535 64.105 181.075 ;
        RECT 60.705 180.395 60.905 180.430 ;
        RECT 62.235 180.395 63.410 180.455 ;
        RECT 60.705 180.285 63.410 180.395 ;
        RECT 64.275 180.365 64.795 180.905 ;
        RECT 64.965 180.555 65.320 180.925 ;
        RECT 65.600 180.915 65.770 181.105 ;
        RECT 65.940 181.080 66.195 181.655 ;
        RECT 65.600 180.585 65.855 180.915 ;
        RECT 65.600 180.375 65.770 180.585 ;
        RECT 60.765 180.225 62.565 180.285 ;
        RECT 62.235 180.195 62.565 180.225 ;
        RECT 60.365 179.445 60.625 180.125 ;
        RECT 60.795 179.275 61.045 180.055 ;
        RECT 61.295 180.025 62.130 180.035 ;
        RECT 62.720 180.025 62.905 180.115 ;
        RECT 61.295 179.825 62.905 180.025 ;
        RECT 61.295 179.445 61.545 179.825 ;
        RECT 62.675 179.785 62.905 179.825 ;
        RECT 63.155 179.665 63.410 180.285 ;
        RECT 61.715 179.275 62.070 179.655 ;
        RECT 63.075 179.445 63.410 179.665 ;
        RECT 63.585 179.275 64.795 180.365 ;
        RECT 65.055 180.205 65.770 180.375 ;
        RECT 66.025 180.350 66.195 181.080 ;
        RECT 66.370 180.985 66.630 181.825 ;
        RECT 66.805 181.055 69.395 181.825 ;
        RECT 66.805 180.535 68.015 181.055 ;
        RECT 70.065 181.005 70.295 181.825 ;
        RECT 70.465 181.025 70.795 181.655 ;
        RECT 65.055 179.445 65.225 180.205 ;
        RECT 65.440 179.275 65.770 180.035 ;
        RECT 65.940 179.445 66.195 180.350 ;
        RECT 66.370 179.275 66.630 180.425 ;
        RECT 68.185 180.365 69.395 180.885 ;
        RECT 70.045 180.585 70.375 180.835 ;
        RECT 70.545 180.425 70.795 181.025 ;
        RECT 70.965 181.005 71.175 181.825 ;
        RECT 71.405 181.055 73.075 181.825 ;
        RECT 71.405 180.535 72.155 181.055 ;
        RECT 73.765 181.005 73.975 181.825 ;
        RECT 74.145 181.025 74.475 181.655 ;
        RECT 66.805 179.275 69.395 180.365 ;
        RECT 70.065 179.275 70.295 180.415 ;
        RECT 70.465 179.445 70.795 180.425 ;
        RECT 70.965 179.275 71.175 180.415 ;
        RECT 72.325 180.365 73.075 180.885 ;
        RECT 74.145 180.425 74.395 181.025 ;
        RECT 74.645 181.005 74.875 181.825 ;
        RECT 75.085 181.150 75.345 181.655 ;
        RECT 75.525 181.445 75.855 181.825 ;
        RECT 76.035 181.275 76.205 181.655 ;
        RECT 74.565 180.585 74.895 180.835 ;
        RECT 71.405 179.275 73.075 180.365 ;
        RECT 73.765 179.275 73.975 180.415 ;
        RECT 74.145 179.445 74.475 180.425 ;
        RECT 74.645 179.275 74.875 180.415 ;
        RECT 75.085 180.350 75.265 181.150 ;
        RECT 75.540 181.105 76.205 181.275 ;
        RECT 75.540 180.850 75.710 181.105 ;
        RECT 75.435 180.520 75.710 180.850 ;
        RECT 75.935 180.555 76.275 180.925 ;
        RECT 75.540 180.375 75.710 180.520 ;
        RECT 75.085 179.445 75.355 180.350 ;
        RECT 75.540 180.205 76.215 180.375 ;
        RECT 75.525 179.275 75.855 180.035 ;
        RECT 76.035 179.445 76.215 180.205 ;
        RECT 76.465 179.445 77.215 181.655 ;
        RECT 77.475 181.275 77.645 181.655 ;
        RECT 77.825 181.445 78.155 181.825 ;
        RECT 77.475 181.105 78.140 181.275 ;
        RECT 78.335 181.150 78.595 181.655 ;
        RECT 77.405 180.555 77.745 180.925 ;
        RECT 77.970 180.850 78.140 181.105 ;
        RECT 77.970 180.520 78.245 180.850 ;
        RECT 77.970 180.375 78.140 180.520 ;
        RECT 77.465 180.205 78.140 180.375 ;
        RECT 78.415 180.350 78.595 181.150 ;
        RECT 78.765 181.100 79.055 181.825 ;
        RECT 79.235 181.230 79.485 181.655 ;
        RECT 79.655 181.400 79.985 181.825 ;
        RECT 80.155 181.405 81.245 181.655 ;
        RECT 81.435 181.405 82.525 181.655 ;
        RECT 80.155 181.230 80.325 181.405 ;
        RECT 79.235 181.060 80.325 181.230 ;
        RECT 80.495 181.065 82.185 181.235 ;
        RECT 82.355 181.230 82.525 181.405 ;
        RECT 82.695 181.400 83.025 181.825 ;
        RECT 83.195 181.230 83.515 181.655 ;
        RECT 79.290 180.635 79.920 180.835 ;
        RECT 80.210 180.805 80.840 180.835 ;
        RECT 80.205 180.635 80.840 180.805 ;
        RECT 77.465 179.445 77.645 180.205 ;
        RECT 77.825 179.275 78.155 180.035 ;
        RECT 78.325 179.445 78.595 180.350 ;
        RECT 78.765 179.275 79.055 180.440 ;
        RECT 79.285 180.425 79.455 180.465 ;
        RECT 81.010 180.425 81.300 181.065 ;
        RECT 82.355 181.060 83.515 181.230 ;
        RECT 84.805 181.005 85.015 181.825 ;
        RECT 85.185 181.025 85.515 181.655 ;
        RECT 81.585 180.635 82.240 180.835 ;
        RECT 82.530 180.805 83.640 180.835 ;
        RECT 82.505 180.635 83.640 180.805 ;
        RECT 85.185 180.425 85.435 181.025 ;
        RECT 85.685 181.005 85.915 181.825 ;
        RECT 86.215 181.275 86.385 181.655 ;
        RECT 86.565 181.445 86.895 181.825 ;
        RECT 86.215 181.105 86.880 181.275 ;
        RECT 87.075 181.150 87.335 181.655 ;
        RECT 85.605 180.585 85.935 180.835 ;
        RECT 86.145 180.555 86.475 180.925 ;
        RECT 86.710 180.850 86.880 181.105 ;
        RECT 86.710 180.520 86.995 180.850 ;
        RECT 79.235 180.255 81.300 180.425 ;
        RECT 79.235 179.445 79.485 180.255 ;
        RECT 79.655 179.615 79.905 180.085 ;
        RECT 80.075 179.785 80.405 180.255 ;
        RECT 80.575 179.615 80.745 180.085 ;
        RECT 80.915 179.785 81.300 180.255 ;
        RECT 81.515 180.255 83.445 180.425 ;
        RECT 81.515 179.615 81.765 180.255 ;
        RECT 79.655 179.445 81.765 179.615 ;
        RECT 81.935 179.275 82.105 180.085 ;
        RECT 82.275 179.445 82.605 180.255 ;
        RECT 82.775 179.275 82.945 180.085 ;
        RECT 83.115 179.445 83.445 180.255 ;
        RECT 84.805 179.275 85.015 180.415 ;
        RECT 85.185 179.445 85.515 180.425 ;
        RECT 85.685 179.275 85.915 180.415 ;
        RECT 86.710 180.375 86.880 180.520 ;
        RECT 86.215 180.205 86.880 180.375 ;
        RECT 87.165 180.350 87.335 181.150 ;
        RECT 87.595 181.275 87.765 181.655 ;
        RECT 87.945 181.445 88.275 181.825 ;
        RECT 87.595 181.105 88.260 181.275 ;
        RECT 88.455 181.150 88.715 181.655 ;
        RECT 87.525 180.555 87.865 180.925 ;
        RECT 88.090 180.850 88.260 181.105 ;
        RECT 88.090 180.520 88.365 180.850 ;
        RECT 88.090 180.375 88.260 180.520 ;
        RECT 86.215 179.445 86.385 180.205 ;
        RECT 86.565 179.275 86.895 180.035 ;
        RECT 87.065 179.445 87.335 180.350 ;
        RECT 87.585 180.205 88.260 180.375 ;
        RECT 88.535 180.350 88.715 181.150 ;
        RECT 88.895 181.015 89.165 181.825 ;
        RECT 89.335 181.015 89.665 181.655 ;
        RECT 89.835 181.015 90.075 181.825 ;
        RECT 88.885 180.585 89.235 180.835 ;
        RECT 89.405 180.415 89.575 181.015 ;
        RECT 90.325 181.005 90.535 181.825 ;
        RECT 90.705 181.025 91.035 181.655 ;
        RECT 89.745 180.585 90.095 180.835 ;
        RECT 90.705 180.425 90.955 181.025 ;
        RECT 91.205 181.005 91.435 181.825 ;
        RECT 91.705 181.005 91.915 181.825 ;
        RECT 92.085 181.025 92.415 181.655 ;
        RECT 91.125 180.585 91.455 180.835 ;
        RECT 92.085 180.425 92.335 181.025 ;
        RECT 92.585 181.005 92.815 181.825 ;
        RECT 93.035 181.315 93.485 181.825 ;
        RECT 93.760 181.405 95.065 181.655 ;
        RECT 95.245 181.425 95.575 181.825 ;
        RECT 94.885 181.255 95.065 181.405 ;
        RECT 96.765 181.345 97.045 181.825 ;
        RECT 92.505 180.585 92.835 180.835 ;
        RECT 93.065 180.635 93.515 181.145 ;
        RECT 93.930 180.835 94.180 181.235 ;
        RECT 93.705 180.635 94.180 180.835 ;
        RECT 94.430 180.835 94.640 181.235 ;
        RECT 94.885 181.085 95.615 181.255 ;
        RECT 97.215 181.175 97.475 181.565 ;
        RECT 97.650 181.345 97.905 181.825 ;
        RECT 98.075 181.175 98.370 181.565 ;
        RECT 98.550 181.345 98.825 181.825 ;
        RECT 98.995 181.325 99.295 181.655 ;
        RECT 94.430 180.635 94.780 180.835 ;
        RECT 94.950 180.585 95.275 180.915 ;
        RECT 87.585 179.445 87.765 180.205 ;
        RECT 87.945 179.275 88.275 180.035 ;
        RECT 88.445 179.445 88.715 180.350 ;
        RECT 88.895 179.275 89.225 180.415 ;
        RECT 89.405 180.245 90.085 180.415 ;
        RECT 89.755 179.460 90.085 180.245 ;
        RECT 90.325 179.275 90.535 180.415 ;
        RECT 90.705 179.445 91.035 180.425 ;
        RECT 91.205 179.275 91.435 180.415 ;
        RECT 91.705 179.275 91.915 180.415 ;
        RECT 92.085 179.445 92.415 180.425 ;
        RECT 93.035 180.415 94.780 180.465 ;
        RECT 95.445 180.415 95.615 181.085 ;
        RECT 92.585 179.275 92.815 180.415 ;
        RECT 93.035 180.285 95.615 180.415 ;
        RECT 96.720 181.005 98.370 181.175 ;
        RECT 96.720 180.495 97.125 181.005 ;
        RECT 97.295 180.665 98.435 180.835 ;
        RECT 96.720 180.325 97.475 180.495 ;
        RECT 93.035 179.615 93.365 180.285 ;
        RECT 94.555 180.245 95.615 180.285 ;
        RECT 93.535 180.075 94.415 180.115 ;
        RECT 93.535 179.875 95.065 180.075 ;
        RECT 93.535 179.825 94.150 179.875 ;
        RECT 93.535 179.785 93.765 179.825 ;
        RECT 94.895 179.745 95.065 179.875 ;
        RECT 93.875 179.615 94.205 179.655 ;
        RECT 93.035 179.445 94.205 179.615 ;
        RECT 94.375 179.275 94.750 179.655 ;
        RECT 95.300 179.275 95.565 180.055 ;
        RECT 96.760 179.275 97.045 180.145 ;
        RECT 97.215 180.075 97.475 180.325 ;
        RECT 98.265 180.415 98.435 180.665 ;
        RECT 98.605 180.585 98.955 181.155 ;
        RECT 99.125 180.415 99.295 181.325 ;
        RECT 98.265 180.245 99.295 180.415 ;
        RECT 97.215 179.905 98.335 180.075 ;
        RECT 97.215 179.445 97.475 179.905 ;
        RECT 97.650 179.275 97.905 179.735 ;
        RECT 98.075 179.445 98.335 179.905 ;
        RECT 98.505 179.275 98.815 180.075 ;
        RECT 98.985 179.445 99.295 180.245 ;
        RECT 99.465 181.325 99.725 181.655 ;
        RECT 99.895 181.465 100.225 181.825 ;
        RECT 100.480 181.445 101.780 181.655 ;
        RECT 99.465 180.125 99.635 181.325 ;
        RECT 100.480 181.295 100.650 181.445 ;
        RECT 99.895 181.170 100.650 181.295 ;
        RECT 99.805 181.125 100.650 181.170 ;
        RECT 99.805 181.005 100.075 181.125 ;
        RECT 99.805 180.430 99.975 181.005 ;
        RECT 100.205 180.565 100.615 180.870 ;
        RECT 100.905 180.835 101.115 181.235 ;
        RECT 100.785 180.625 101.115 180.835 ;
        RECT 101.360 180.835 101.580 181.235 ;
        RECT 102.055 181.060 102.510 181.825 ;
        RECT 102.775 181.275 102.945 181.655 ;
        RECT 103.160 181.445 103.490 181.825 ;
        RECT 102.775 181.105 103.490 181.275 ;
        RECT 101.360 180.625 101.835 180.835 ;
        RECT 102.025 180.635 102.515 180.835 ;
        RECT 102.685 180.555 103.040 180.925 ;
        RECT 103.320 180.915 103.490 181.105 ;
        RECT 103.660 181.080 103.915 181.655 ;
        RECT 103.320 180.585 103.575 180.915 ;
        RECT 99.805 180.395 100.005 180.430 ;
        RECT 101.335 180.395 102.510 180.455 ;
        RECT 99.805 180.285 102.510 180.395 ;
        RECT 103.320 180.375 103.490 180.585 ;
        RECT 99.865 180.225 101.665 180.285 ;
        RECT 101.335 180.195 101.665 180.225 ;
        RECT 99.465 179.445 99.725 180.125 ;
        RECT 99.895 179.275 100.145 180.055 ;
        RECT 100.395 180.025 101.230 180.035 ;
        RECT 101.820 180.025 102.005 180.115 ;
        RECT 100.395 179.825 102.005 180.025 ;
        RECT 100.395 179.445 100.645 179.825 ;
        RECT 101.775 179.785 102.005 179.825 ;
        RECT 102.255 179.665 102.510 180.285 ;
        RECT 100.815 179.275 101.170 179.655 ;
        RECT 102.175 179.445 102.510 179.665 ;
        RECT 102.775 180.205 103.490 180.375 ;
        RECT 103.745 180.350 103.915 181.080 ;
        RECT 104.090 180.985 104.350 181.825 ;
        RECT 104.525 181.100 104.815 181.825 ;
        RECT 105.535 181.345 105.835 181.825 ;
        RECT 106.005 181.175 106.265 181.630 ;
        RECT 106.435 181.345 106.695 181.825 ;
        RECT 106.875 181.175 107.135 181.630 ;
        RECT 107.305 181.345 107.555 181.825 ;
        RECT 107.735 181.175 107.995 181.630 ;
        RECT 108.165 181.345 108.415 181.825 ;
        RECT 108.595 181.175 108.855 181.630 ;
        RECT 109.025 181.345 109.270 181.825 ;
        RECT 109.440 181.175 109.715 181.630 ;
        RECT 109.885 181.345 110.130 181.825 ;
        RECT 110.300 181.175 110.560 181.630 ;
        RECT 110.730 181.345 110.990 181.825 ;
        RECT 111.160 181.175 111.420 181.630 ;
        RECT 111.590 181.345 111.850 181.825 ;
        RECT 112.020 181.175 112.280 181.630 ;
        RECT 112.450 181.265 112.710 181.825 ;
        RECT 105.535 181.005 112.280 181.175 ;
        RECT 102.775 179.445 102.945 180.205 ;
        RECT 103.160 179.275 103.490 180.035 ;
        RECT 103.660 179.445 103.915 180.350 ;
        RECT 104.090 179.275 104.350 180.425 ;
        RECT 104.525 179.275 104.815 180.440 ;
        RECT 105.535 180.415 106.700 181.005 ;
        RECT 112.880 180.835 113.130 181.645 ;
        RECT 113.310 181.300 113.570 181.825 ;
        RECT 113.740 180.835 113.990 181.645 ;
        RECT 114.170 181.315 114.475 181.825 ;
        RECT 114.735 181.345 115.035 181.825 ;
        RECT 115.205 181.175 115.465 181.630 ;
        RECT 115.635 181.345 115.895 181.825 ;
        RECT 116.075 181.175 116.335 181.630 ;
        RECT 116.505 181.345 116.755 181.825 ;
        RECT 116.935 181.175 117.195 181.630 ;
        RECT 117.365 181.345 117.615 181.825 ;
        RECT 117.795 181.175 118.055 181.630 ;
        RECT 118.225 181.345 118.470 181.825 ;
        RECT 118.640 181.175 118.915 181.630 ;
        RECT 119.085 181.345 119.330 181.825 ;
        RECT 119.500 181.175 119.760 181.630 ;
        RECT 119.930 181.345 120.190 181.825 ;
        RECT 120.360 181.175 120.620 181.630 ;
        RECT 120.790 181.345 121.050 181.825 ;
        RECT 121.220 181.175 121.480 181.630 ;
        RECT 121.650 181.265 121.910 181.825 ;
        RECT 106.870 180.585 113.990 180.835 ;
        RECT 114.160 180.585 114.475 181.145 ;
        RECT 114.735 181.005 121.480 181.175 ;
        RECT 105.535 180.190 112.280 180.415 ;
        RECT 105.535 179.275 105.805 180.020 ;
        RECT 105.975 179.450 106.265 180.190 ;
        RECT 106.875 180.175 112.280 180.190 ;
        RECT 106.435 179.280 106.690 180.005 ;
        RECT 106.875 179.450 107.135 180.175 ;
        RECT 107.305 179.280 107.550 180.005 ;
        RECT 107.735 179.450 107.995 180.175 ;
        RECT 108.165 179.280 108.410 180.005 ;
        RECT 108.595 179.450 108.855 180.175 ;
        RECT 109.025 179.280 109.270 180.005 ;
        RECT 109.440 179.450 109.700 180.175 ;
        RECT 109.870 179.280 110.130 180.005 ;
        RECT 110.300 179.450 110.560 180.175 ;
        RECT 110.730 179.280 110.990 180.005 ;
        RECT 111.160 179.450 111.420 180.175 ;
        RECT 111.590 179.280 111.850 180.005 ;
        RECT 112.020 179.450 112.280 180.175 ;
        RECT 112.450 179.280 112.710 180.075 ;
        RECT 112.880 179.450 113.130 180.585 ;
        RECT 106.435 179.275 112.710 179.280 ;
        RECT 113.310 179.275 113.570 180.085 ;
        RECT 113.745 179.445 113.990 180.585 ;
        RECT 114.735 180.415 115.900 181.005 ;
        RECT 122.080 180.835 122.330 181.645 ;
        RECT 122.510 181.300 122.770 181.825 ;
        RECT 122.940 180.835 123.190 181.645 ;
        RECT 123.370 181.315 123.675 181.825 ;
        RECT 123.845 181.485 125.205 181.655 ;
        RECT 116.070 180.585 123.190 180.835 ;
        RECT 123.360 180.585 123.675 181.145 ;
        RECT 123.845 181.005 124.205 181.485 ;
        RECT 124.375 181.085 124.705 181.315 ;
        RECT 124.875 181.255 125.205 181.485 ;
        RECT 125.375 181.425 125.705 181.825 ;
        RECT 125.875 181.255 126.205 181.655 ;
        RECT 124.875 181.085 126.205 181.255 ;
        RECT 126.475 181.085 126.805 181.825 ;
        RECT 123.845 180.665 124.205 180.835 ;
        RECT 123.845 180.585 124.175 180.665 ;
        RECT 114.735 180.190 121.480 180.415 ;
        RECT 114.170 179.275 114.465 180.085 ;
        RECT 114.735 179.275 115.005 180.020 ;
        RECT 115.175 179.450 115.465 180.190 ;
        RECT 116.075 180.175 121.480 180.190 ;
        RECT 115.635 179.280 115.890 180.005 ;
        RECT 116.075 179.450 116.335 180.175 ;
        RECT 116.505 179.280 116.750 180.005 ;
        RECT 116.935 179.450 117.195 180.175 ;
        RECT 117.365 179.280 117.610 180.005 ;
        RECT 117.795 179.450 118.055 180.175 ;
        RECT 118.225 179.280 118.470 180.005 ;
        RECT 118.640 179.450 118.900 180.175 ;
        RECT 119.070 179.280 119.330 180.005 ;
        RECT 119.500 179.450 119.760 180.175 ;
        RECT 119.930 179.280 120.190 180.005 ;
        RECT 120.360 179.450 120.620 180.175 ;
        RECT 120.790 179.280 121.050 180.005 ;
        RECT 121.220 179.450 121.480 180.175 ;
        RECT 121.650 179.280 121.910 180.075 ;
        RECT 122.080 179.450 122.330 180.585 ;
        RECT 115.635 179.275 121.910 179.280 ;
        RECT 122.510 179.275 122.770 180.085 ;
        RECT 122.945 179.445 123.190 180.585 ;
        RECT 123.370 179.275 123.665 180.085 ;
        RECT 123.845 179.275 124.205 180.415 ;
        RECT 124.375 180.125 124.575 181.085 ;
        RECT 124.745 180.465 124.990 180.915 ;
        RECT 124.745 180.295 124.995 180.465 ;
        RECT 125.265 180.295 125.485 180.915 ;
        RECT 125.740 180.295 125.915 180.915 ;
        RECT 126.185 180.295 126.405 180.915 ;
        RECT 126.575 180.125 126.885 180.915 ;
        RECT 124.375 179.955 126.885 180.125 ;
        RECT 124.875 179.445 125.205 179.955 ;
        RECT 126.375 179.275 126.885 179.785 ;
        RECT 127.055 179.445 127.385 181.655 ;
        RECT 127.555 181.025 127.815 181.825 ;
        RECT 128.035 181.355 128.325 181.825 ;
        RECT 128.495 181.185 128.825 181.655 ;
        RECT 128.995 181.355 129.165 181.825 ;
        RECT 129.335 181.185 129.665 181.655 ;
        RECT 128.495 181.175 129.665 181.185 ;
        RECT 128.065 181.145 129.665 181.175 ;
        RECT 128.045 181.005 129.665 181.145 ;
        RECT 129.835 181.005 130.110 181.825 ;
        RECT 130.285 181.100 130.575 181.825 ;
        RECT 131.205 181.005 131.500 181.825 ;
        RECT 131.670 181.085 132.110 181.645 ;
        RECT 132.280 181.085 132.730 181.825 ;
        RECT 132.900 181.255 133.070 181.655 ;
        RECT 133.240 181.425 133.660 181.825 ;
        RECT 133.830 181.255 134.060 181.655 ;
        RECT 132.900 181.085 134.060 181.255 ;
        RECT 134.230 181.085 134.715 181.655 ;
        RECT 128.045 180.975 128.280 181.005 ;
        RECT 128.065 180.465 128.280 180.975 ;
        RECT 131.670 180.835 131.980 181.085 ;
        RECT 128.450 180.635 129.220 180.835 ;
        RECT 129.390 180.635 130.110 180.835 ;
        RECT 131.205 180.615 131.980 180.835 ;
        RECT 127.555 179.275 127.815 180.415 ;
        RECT 128.065 180.245 128.825 180.465 ;
        RECT 128.025 179.615 128.325 180.075 ;
        RECT 128.495 179.785 128.825 180.245 ;
        RECT 128.995 180.245 130.110 180.455 ;
        RECT 128.995 179.615 129.165 180.245 ;
        RECT 128.025 179.445 129.165 179.615 ;
        RECT 129.335 179.275 129.665 180.075 ;
        RECT 129.835 179.445 130.110 180.245 ;
        RECT 130.285 179.275 130.575 180.440 ;
        RECT 131.205 179.275 131.500 180.445 ;
        RECT 131.670 180.075 131.980 180.615 ;
        RECT 132.150 180.465 132.320 180.915 ;
        RECT 132.490 180.635 132.880 180.915 ;
        RECT 133.065 180.585 133.310 180.915 ;
        RECT 132.150 180.295 132.940 180.465 ;
        RECT 131.670 179.445 132.110 180.075 ;
        RECT 132.285 179.275 132.600 180.125 ;
        RECT 132.770 179.615 132.940 180.295 ;
        RECT 133.110 179.785 133.310 180.585 ;
        RECT 133.510 179.785 133.760 180.915 ;
        RECT 133.975 180.585 134.375 180.915 ;
        RECT 134.545 180.415 134.715 181.085 ;
        RECT 133.950 180.245 134.715 180.415 ;
        RECT 134.885 181.085 135.370 181.655 ;
        RECT 135.540 181.255 135.770 181.655 ;
        RECT 135.940 181.425 136.360 181.825 ;
        RECT 136.530 181.255 136.700 181.655 ;
        RECT 135.540 181.085 136.700 181.255 ;
        RECT 136.870 181.085 137.320 181.825 ;
        RECT 137.490 181.085 137.930 181.645 ;
        RECT 134.885 180.415 135.055 181.085 ;
        RECT 135.225 180.585 135.625 180.915 ;
        RECT 134.885 180.245 135.650 180.415 ;
        RECT 133.950 179.615 134.200 180.245 ;
        RECT 132.770 179.445 134.200 179.615 ;
        RECT 134.375 179.275 134.710 180.075 ;
        RECT 134.890 179.275 135.225 180.075 ;
        RECT 135.400 179.615 135.650 180.245 ;
        RECT 135.840 179.785 136.090 180.915 ;
        RECT 136.290 180.585 136.535 180.915 ;
        RECT 136.720 180.635 137.110 180.915 ;
        RECT 136.290 179.785 136.490 180.585 ;
        RECT 137.280 180.465 137.450 180.915 ;
        RECT 136.660 180.295 137.450 180.465 ;
        RECT 137.620 180.835 137.930 181.085 ;
        RECT 138.100 181.005 138.395 181.825 ;
        RECT 138.565 181.075 139.775 181.825 ;
        RECT 137.620 180.615 138.395 180.835 ;
        RECT 136.660 179.615 136.830 180.295 ;
        RECT 135.400 179.445 136.830 179.615 ;
        RECT 137.000 179.275 137.315 180.125 ;
        RECT 137.620 180.075 137.930 180.615 ;
        RECT 137.490 179.445 137.930 180.075 ;
        RECT 138.100 179.275 138.395 180.445 ;
        RECT 138.565 180.365 139.085 180.905 ;
        RECT 139.255 180.535 139.775 181.075 ;
        RECT 138.565 179.275 139.775 180.365 ;
        RECT 27.160 179.105 139.860 179.275 ;
        RECT 27.245 178.015 28.455 179.105 ;
        RECT 28.625 178.670 33.970 179.105 ;
        RECT 34.145 178.670 39.490 179.105 ;
        RECT 27.245 177.305 27.765 177.845 ;
        RECT 27.935 177.475 28.455 178.015 ;
        RECT 27.245 176.555 28.455 177.305 ;
        RECT 30.210 177.100 30.550 177.930 ;
        RECT 32.030 177.420 32.380 178.670 ;
        RECT 35.730 177.100 36.070 177.930 ;
        RECT 37.550 177.420 37.900 178.670 ;
        RECT 40.125 177.940 40.415 179.105 ;
        RECT 41.135 178.485 41.305 178.915 ;
        RECT 41.475 178.655 41.805 179.105 ;
        RECT 41.135 178.255 41.815 178.485 ;
        RECT 41.110 177.405 41.410 178.085 ;
        RECT 28.625 176.555 33.970 177.100 ;
        RECT 34.145 176.555 39.490 177.100 ;
        RECT 40.125 176.555 40.415 177.280 ;
        RECT 41.105 177.235 41.410 177.405 ;
        RECT 41.580 177.605 41.815 178.255 ;
        RECT 42.005 177.945 42.290 178.890 ;
        RECT 42.470 178.635 43.155 179.105 ;
        RECT 42.465 178.115 43.160 178.425 ;
        RECT 43.335 178.050 43.640 178.835 ;
        RECT 43.825 178.150 44.095 179.105 ;
        RECT 42.005 177.795 42.865 177.945 ;
        RECT 42.005 177.775 43.295 177.795 ;
        RECT 41.580 177.275 42.135 177.605 ;
        RECT 42.305 177.415 43.295 177.775 ;
        RECT 41.580 177.125 41.795 177.275 ;
        RECT 41.055 176.555 41.385 177.060 ;
        RECT 41.555 176.750 41.795 177.125 ;
        RECT 42.305 177.080 42.475 177.415 ;
        RECT 43.465 177.245 43.640 178.050 ;
        RECT 42.075 176.885 42.475 177.080 ;
        RECT 42.075 176.740 42.245 176.885 ;
        RECT 42.835 176.555 43.235 177.050 ;
        RECT 43.405 176.725 43.640 177.245 ;
        RECT 44.725 177.500 45.005 178.935 ;
        RECT 45.175 178.330 45.885 179.105 ;
        RECT 46.055 178.160 46.385 178.935 ;
        RECT 45.235 177.945 46.385 178.160 ;
        RECT 43.825 176.555 44.095 177.190 ;
        RECT 44.725 176.725 45.065 177.500 ;
        RECT 45.235 177.375 45.520 177.945 ;
        RECT 45.705 177.545 46.175 177.775 ;
        RECT 46.580 177.745 46.795 178.860 ;
        RECT 46.975 178.385 47.305 179.105 ;
        RECT 47.485 178.670 52.830 179.105 ;
        RECT 47.085 177.745 47.315 178.085 ;
        RECT 46.345 177.565 46.795 177.745 ;
        RECT 46.345 177.545 46.675 177.565 ;
        RECT 46.985 177.545 47.315 177.745 ;
        RECT 45.235 177.185 45.945 177.375 ;
        RECT 45.645 177.045 45.945 177.185 ;
        RECT 46.135 177.185 47.315 177.375 ;
        RECT 46.135 177.105 46.465 177.185 ;
        RECT 45.645 177.035 45.960 177.045 ;
        RECT 45.645 177.025 45.970 177.035 ;
        RECT 45.645 177.020 45.980 177.025 ;
        RECT 45.235 176.555 45.405 177.015 ;
        RECT 45.645 177.010 45.985 177.020 ;
        RECT 45.645 177.005 45.990 177.010 ;
        RECT 45.645 176.995 45.995 177.005 ;
        RECT 45.645 176.990 46.000 176.995 ;
        RECT 45.645 176.725 46.005 176.990 ;
        RECT 46.635 176.555 46.805 177.015 ;
        RECT 46.975 176.725 47.315 177.185 ;
        RECT 49.070 177.100 49.410 177.930 ;
        RECT 50.890 177.420 51.240 178.670 ;
        RECT 53.005 178.015 54.675 179.105 ;
        RECT 55.800 178.305 56.050 179.105 ;
        RECT 56.220 178.475 56.550 178.935 ;
        RECT 56.720 178.645 56.935 179.105 ;
        RECT 56.220 178.305 57.390 178.475 ;
        RECT 53.005 177.325 53.755 177.845 ;
        RECT 53.925 177.495 54.675 178.015 ;
        RECT 55.310 178.135 55.590 178.295 ;
        RECT 55.310 177.965 56.645 178.135 ;
        RECT 56.475 177.795 56.645 177.965 ;
        RECT 55.310 177.545 55.660 177.785 ;
        RECT 55.830 177.545 56.305 177.785 ;
        RECT 56.475 177.545 56.850 177.795 ;
        RECT 56.475 177.375 56.645 177.545 ;
        RECT 47.485 176.555 52.830 177.100 ;
        RECT 53.005 176.555 54.675 177.325 ;
        RECT 55.310 177.205 56.645 177.375 ;
        RECT 55.310 176.995 55.580 177.205 ;
        RECT 57.020 177.015 57.390 178.305 ;
        RECT 57.605 178.015 60.195 179.105 ;
        RECT 55.800 176.555 56.130 177.015 ;
        RECT 56.640 176.725 57.390 177.015 ;
        RECT 57.605 177.325 58.815 177.845 ;
        RECT 58.985 177.495 60.195 178.015 ;
        RECT 60.835 177.965 61.165 179.105 ;
        RECT 61.695 178.135 62.025 178.920 ;
        RECT 61.345 177.965 62.025 178.135 ;
        RECT 62.295 178.135 62.465 178.935 ;
        RECT 63.225 178.475 63.475 178.935 ;
        RECT 63.675 178.725 64.345 179.105 ;
        RECT 64.535 178.475 64.785 178.935 ;
        RECT 64.960 178.645 65.205 179.105 ;
        RECT 63.225 178.305 64.785 178.475 ;
        RECT 65.375 178.255 65.715 178.895 ;
        RECT 62.295 177.965 65.235 178.135 ;
        RECT 60.825 177.545 61.175 177.795 ;
        RECT 61.345 177.365 61.515 177.965 ;
        RECT 65.065 177.795 65.235 177.965 ;
        RECT 61.685 177.545 62.035 177.795 ;
        RECT 62.265 177.465 62.450 177.795 ;
        RECT 62.705 177.465 63.180 177.795 ;
        RECT 63.490 177.465 63.835 177.795 ;
        RECT 57.605 176.555 60.195 177.325 ;
        RECT 60.835 176.555 61.105 177.365 ;
        RECT 61.275 176.725 61.605 177.365 ;
        RECT 61.775 176.555 62.015 177.365 ;
        RECT 62.295 177.125 63.475 177.295 ;
        RECT 63.645 177.235 63.835 177.465 ;
        RECT 64.095 177.220 64.290 177.795 ;
        RECT 64.560 177.465 64.895 177.795 ;
        RECT 65.065 177.465 65.375 177.795 ;
        RECT 65.065 177.295 65.235 177.465 ;
        RECT 62.295 176.725 62.465 177.125 ;
        RECT 62.705 176.555 63.035 176.955 ;
        RECT 63.305 176.895 63.475 177.125 ;
        RECT 64.540 177.125 65.235 177.295 ;
        RECT 65.545 177.140 65.715 178.255 ;
        RECT 65.885 177.940 66.175 179.105 ;
        RECT 66.435 178.135 66.605 178.935 ;
        RECT 67.365 178.475 67.615 178.935 ;
        RECT 67.815 178.725 68.485 179.105 ;
        RECT 68.675 178.475 68.925 178.935 ;
        RECT 69.100 178.645 69.345 179.105 ;
        RECT 67.365 178.305 68.925 178.475 ;
        RECT 69.515 178.255 69.855 178.895 ;
        RECT 66.435 177.965 69.375 178.135 ;
        RECT 69.205 177.795 69.375 177.965 ;
        RECT 66.405 177.465 66.590 177.795 ;
        RECT 66.845 177.465 67.320 177.795 ;
        RECT 67.630 177.465 67.975 177.795 ;
        RECT 64.540 176.895 64.710 177.125 ;
        RECT 63.305 176.725 64.710 176.895 ;
        RECT 64.880 176.555 65.210 176.935 ;
        RECT 65.405 176.725 65.715 177.140 ;
        RECT 65.885 176.555 66.175 177.280 ;
        RECT 66.435 177.125 67.615 177.295 ;
        RECT 67.785 177.235 67.975 177.465 ;
        RECT 68.235 177.220 68.430 177.795 ;
        RECT 68.700 177.465 69.035 177.795 ;
        RECT 69.205 177.465 69.515 177.795 ;
        RECT 69.205 177.295 69.375 177.465 ;
        RECT 66.435 176.725 66.605 177.125 ;
        RECT 66.845 176.555 67.175 176.955 ;
        RECT 67.445 176.895 67.615 177.125 ;
        RECT 68.680 177.125 69.375 177.295 ;
        RECT 69.685 177.140 69.855 178.255 ;
        RECT 70.035 177.965 70.365 179.105 ;
        RECT 70.895 178.135 71.225 178.920 ;
        RECT 70.545 177.965 71.225 178.135 ;
        RECT 70.025 177.545 70.375 177.795 ;
        RECT 70.545 177.365 70.715 177.965 ;
        RECT 70.885 177.545 71.235 177.795 ;
        RECT 71.405 177.385 71.925 178.935 ;
        RECT 72.095 178.380 72.425 179.105 ;
        RECT 68.680 176.895 68.850 177.125 ;
        RECT 67.445 176.725 68.850 176.895 ;
        RECT 69.020 176.555 69.350 176.935 ;
        RECT 69.545 176.725 69.855 177.140 ;
        RECT 70.035 176.555 70.305 177.365 ;
        RECT 70.475 176.725 70.805 177.365 ;
        RECT 70.975 176.555 71.215 177.365 ;
        RECT 71.585 176.555 71.925 177.215 ;
        RECT 72.095 176.725 72.615 178.210 ;
        RECT 72.785 176.725 73.535 178.935 ;
        RECT 73.795 178.175 73.965 178.935 ;
        RECT 74.145 178.345 74.475 179.105 ;
        RECT 73.795 178.005 74.460 178.175 ;
        RECT 74.645 178.030 74.915 178.935 ;
        RECT 74.290 177.860 74.460 178.005 ;
        RECT 73.725 177.455 74.055 177.825 ;
        RECT 74.290 177.530 74.575 177.860 ;
        RECT 74.290 177.275 74.460 177.530 ;
        RECT 73.795 177.105 74.460 177.275 ;
        RECT 74.745 177.230 74.915 178.030 ;
        RECT 73.795 176.725 73.965 177.105 ;
        RECT 74.145 176.555 74.475 176.935 ;
        RECT 74.655 176.725 74.915 177.230 ;
        RECT 75.095 176.735 75.355 178.925 ;
        RECT 75.525 178.375 75.865 179.105 ;
        RECT 76.045 178.195 76.315 178.925 ;
        RECT 75.545 177.975 76.315 178.195 ;
        RECT 76.495 178.215 76.725 178.925 ;
        RECT 76.895 178.395 77.225 179.105 ;
        RECT 77.395 178.215 77.655 178.925 ;
        RECT 76.495 177.975 77.655 178.215 ;
        RECT 77.855 178.155 78.130 178.925 ;
        RECT 78.300 178.495 78.630 178.925 ;
        RECT 78.800 178.665 78.995 179.105 ;
        RECT 79.175 178.495 79.505 178.925 ;
        RECT 78.300 178.325 79.505 178.495 ;
        RECT 75.545 177.305 75.835 177.975 ;
        RECT 77.855 177.965 78.440 178.155 ;
        RECT 78.610 177.995 79.505 178.325 ;
        RECT 80.605 178.030 80.875 178.935 ;
        RECT 81.045 178.345 81.375 179.105 ;
        RECT 81.555 178.175 81.725 178.935 ;
        RECT 76.015 177.485 76.480 177.795 ;
        RECT 76.660 177.485 77.185 177.795 ;
        RECT 75.545 177.105 76.775 177.305 ;
        RECT 75.615 176.555 76.285 176.925 ;
        RECT 76.465 176.735 76.775 177.105 ;
        RECT 76.955 176.845 77.185 177.485 ;
        RECT 77.365 177.465 77.665 177.795 ;
        RECT 77.365 176.555 77.655 177.285 ;
        RECT 77.855 177.145 78.095 177.795 ;
        RECT 78.265 177.295 78.440 177.965 ;
        RECT 78.610 177.465 79.025 177.795 ;
        RECT 79.205 177.465 79.500 177.795 ;
        RECT 78.265 177.115 78.595 177.295 ;
        RECT 77.870 176.555 78.200 176.945 ;
        RECT 78.370 176.735 78.595 177.115 ;
        RECT 78.795 176.845 79.025 177.465 ;
        RECT 79.205 176.555 79.505 177.285 ;
        RECT 80.605 177.230 80.775 178.030 ;
        RECT 81.060 178.005 81.725 178.175 ;
        RECT 81.060 177.860 81.230 178.005 ;
        RECT 81.985 177.965 82.265 179.105 ;
        RECT 82.435 177.955 82.765 178.935 ;
        RECT 82.935 177.965 83.195 179.105 ;
        RECT 83.370 178.155 83.635 178.925 ;
        RECT 83.805 178.385 84.135 179.105 ;
        RECT 84.325 178.565 84.585 178.925 ;
        RECT 84.755 178.735 85.085 179.105 ;
        RECT 85.255 178.565 85.515 178.925 ;
        RECT 84.325 178.335 85.515 178.565 ;
        RECT 86.085 178.155 86.375 178.925 ;
        RECT 80.945 177.530 81.230 177.860 ;
        RECT 81.060 177.275 81.230 177.530 ;
        RECT 81.465 177.455 81.795 177.825 ;
        RECT 81.995 177.525 82.330 177.795 ;
        RECT 82.500 177.355 82.670 177.955 ;
        RECT 82.840 177.545 83.175 177.795 ;
        RECT 80.605 176.725 80.865 177.230 ;
        RECT 81.060 177.105 81.725 177.275 ;
        RECT 81.045 176.555 81.375 176.935 ;
        RECT 81.555 176.725 81.725 177.105 ;
        RECT 81.985 176.555 82.295 177.355 ;
        RECT 82.500 176.725 83.195 177.355 ;
        RECT 83.370 176.735 83.705 178.155 ;
        RECT 83.880 177.975 86.375 178.155 ;
        RECT 87.045 178.030 87.315 178.935 ;
        RECT 87.485 178.345 87.815 179.105 ;
        RECT 87.995 178.175 88.165 178.935 ;
        RECT 83.880 177.285 84.105 177.975 ;
        RECT 84.305 177.465 84.585 177.795 ;
        RECT 84.765 177.465 85.340 177.795 ;
        RECT 85.520 177.465 85.955 177.795 ;
        RECT 86.135 177.465 86.405 177.795 ;
        RECT 83.880 177.095 86.365 177.285 ;
        RECT 83.885 176.555 84.630 176.925 ;
        RECT 85.195 176.735 85.450 177.095 ;
        RECT 85.630 176.555 85.960 176.925 ;
        RECT 86.140 176.735 86.365 177.095 ;
        RECT 87.045 177.230 87.215 178.030 ;
        RECT 87.500 178.005 88.165 178.175 ;
        RECT 88.515 178.175 88.685 178.935 ;
        RECT 88.865 178.345 89.195 179.105 ;
        RECT 88.515 178.005 89.180 178.175 ;
        RECT 89.365 178.030 89.635 178.935 ;
        RECT 87.500 177.860 87.670 178.005 ;
        RECT 87.385 177.530 87.670 177.860 ;
        RECT 89.010 177.860 89.180 178.005 ;
        RECT 87.500 177.275 87.670 177.530 ;
        RECT 87.905 177.455 88.235 177.825 ;
        RECT 88.445 177.455 88.775 177.825 ;
        RECT 89.010 177.530 89.295 177.860 ;
        RECT 89.010 177.275 89.180 177.530 ;
        RECT 87.045 176.725 87.305 177.230 ;
        RECT 87.500 177.105 88.165 177.275 ;
        RECT 87.485 176.555 87.815 176.935 ;
        RECT 87.995 176.725 88.165 177.105 ;
        RECT 88.515 177.105 89.180 177.275 ;
        RECT 89.465 177.230 89.635 178.030 ;
        RECT 89.815 178.495 90.145 178.925 ;
        RECT 90.325 178.665 90.520 179.105 ;
        RECT 90.690 178.495 91.020 178.925 ;
        RECT 89.815 178.325 91.020 178.495 ;
        RECT 89.815 177.995 90.710 178.325 ;
        RECT 91.190 178.155 91.465 178.925 ;
        RECT 90.880 177.965 91.465 178.155 ;
        RECT 89.820 177.465 90.115 177.795 ;
        RECT 90.295 177.465 90.710 177.795 ;
        RECT 88.515 176.725 88.685 177.105 ;
        RECT 88.865 176.555 89.195 176.935 ;
        RECT 89.375 176.725 89.635 177.230 ;
        RECT 89.815 176.555 90.115 177.285 ;
        RECT 90.295 176.845 90.525 177.465 ;
        RECT 90.880 177.295 91.055 177.965 ;
        RECT 91.645 177.940 91.935 179.105 ;
        RECT 93.520 178.305 93.770 179.105 ;
        RECT 93.940 178.475 94.270 178.935 ;
        RECT 94.440 178.645 94.655 179.105 ;
        RECT 93.940 178.305 95.110 178.475 ;
        RECT 93.030 178.135 93.310 178.295 ;
        RECT 93.030 177.965 94.365 178.135 ;
        RECT 94.195 177.795 94.365 177.965 ;
        RECT 90.725 177.115 91.055 177.295 ;
        RECT 91.225 177.145 91.465 177.795 ;
        RECT 93.030 177.545 93.380 177.785 ;
        RECT 93.550 177.545 94.025 177.785 ;
        RECT 94.195 177.545 94.570 177.795 ;
        RECT 94.195 177.375 94.365 177.545 ;
        RECT 90.725 176.735 90.950 177.115 ;
        RECT 91.120 176.555 91.450 176.945 ;
        RECT 91.645 176.555 91.935 177.280 ;
        RECT 93.030 177.205 94.365 177.375 ;
        RECT 93.030 176.995 93.300 177.205 ;
        RECT 94.740 177.015 95.110 178.305 ;
        RECT 95.325 177.965 95.615 179.105 ;
        RECT 95.785 178.385 96.235 178.935 ;
        RECT 96.425 178.385 96.755 179.105 ;
        RECT 93.520 176.555 93.850 177.015 ;
        RECT 94.360 176.725 95.110 177.015 ;
        RECT 95.325 176.555 95.615 177.355 ;
        RECT 95.785 177.015 96.035 178.385 ;
        RECT 96.965 178.215 97.265 178.765 ;
        RECT 97.435 178.435 97.715 179.105 ;
        RECT 98.385 178.465 98.715 178.895 ;
        RECT 98.260 178.295 98.715 178.465 ;
        RECT 98.895 178.465 99.145 178.885 ;
        RECT 99.375 178.635 99.705 179.105 ;
        RECT 99.935 178.465 100.185 178.885 ;
        RECT 98.895 178.295 100.185 178.465 ;
        RECT 96.325 178.045 97.265 178.215 ;
        RECT 96.325 177.795 96.495 178.045 ;
        RECT 97.600 177.795 97.915 178.235 ;
        RECT 96.205 177.465 96.495 177.795 ;
        RECT 96.665 177.545 96.995 177.795 ;
        RECT 97.225 177.545 97.915 177.795 ;
        RECT 96.325 177.375 96.495 177.465 ;
        RECT 96.325 177.185 97.715 177.375 ;
        RECT 95.785 176.725 96.335 177.015 ;
        RECT 96.505 176.555 96.755 177.015 ;
        RECT 97.385 176.825 97.715 177.185 ;
        RECT 98.260 177.295 98.430 178.295 ;
        RECT 98.600 177.465 98.845 178.125 ;
        RECT 99.060 177.465 99.325 178.125 ;
        RECT 99.520 177.465 99.805 178.125 ;
        RECT 99.980 177.795 100.195 178.125 ;
        RECT 100.375 177.965 100.625 179.105 ;
        RECT 100.795 178.045 101.125 178.895 ;
        RECT 101.400 178.725 101.730 179.105 ;
        RECT 101.900 178.545 102.090 178.935 ;
        RECT 99.980 177.465 100.285 177.795 ;
        RECT 100.455 177.465 100.765 177.795 ;
        RECT 100.455 177.295 100.625 177.465 ;
        RECT 98.260 177.125 100.625 177.295 ;
        RECT 100.935 177.280 101.125 178.045 ;
        RECT 98.415 176.555 98.745 176.955 ;
        RECT 98.915 176.785 99.245 177.125 ;
        RECT 100.295 176.555 100.625 176.955 ;
        RECT 100.795 176.770 101.125 177.280 ;
        RECT 101.360 178.375 102.090 178.545 ;
        RECT 102.270 178.405 102.700 179.105 ;
        RECT 101.360 177.255 101.555 178.375 ;
        RECT 103.205 178.235 103.875 178.935 ;
        RECT 104.045 178.405 104.375 179.105 ;
        RECT 104.545 178.235 104.810 178.935 ;
        RECT 105.075 178.360 105.345 179.105 ;
        RECT 105.975 179.100 112.250 179.105 ;
        RECT 102.235 177.980 104.810 178.235 ;
        RECT 105.515 178.190 105.805 178.930 ;
        RECT 105.975 178.375 106.230 179.100 ;
        RECT 106.415 178.205 106.675 178.930 ;
        RECT 106.845 178.375 107.090 179.100 ;
        RECT 107.275 178.205 107.535 178.930 ;
        RECT 107.705 178.375 107.950 179.100 ;
        RECT 108.135 178.205 108.395 178.930 ;
        RECT 108.565 178.375 108.810 179.100 ;
        RECT 108.980 178.205 109.240 178.930 ;
        RECT 109.410 178.375 109.670 179.100 ;
        RECT 109.840 178.205 110.100 178.930 ;
        RECT 110.270 178.375 110.530 179.100 ;
        RECT 110.700 178.205 110.960 178.930 ;
        RECT 111.130 178.375 111.390 179.100 ;
        RECT 111.560 178.205 111.820 178.930 ;
        RECT 111.990 178.305 112.250 179.100 ;
        RECT 106.415 178.190 111.820 178.205 ;
        RECT 102.235 177.795 102.405 177.980 ;
        RECT 101.725 177.465 102.405 177.795 ;
        RECT 102.575 177.465 102.910 177.795 ;
        RECT 103.080 177.745 103.370 177.795 ;
        RECT 103.080 177.575 103.375 177.745 ;
        RECT 103.080 177.465 103.370 177.575 ;
        RECT 103.660 177.465 104.020 177.795 ;
        RECT 104.190 177.295 104.370 177.980 ;
        RECT 105.075 177.965 111.820 178.190 ;
        RECT 104.540 177.465 104.815 177.795 ;
        RECT 105.075 177.375 106.240 177.965 ;
        RECT 112.420 177.795 112.670 178.930 ;
        RECT 112.850 178.295 113.110 179.105 ;
        RECT 113.285 177.795 113.530 178.935 ;
        RECT 113.710 178.295 114.005 179.105 ;
        RECT 114.200 178.120 114.525 179.105 ;
        RECT 115.095 178.475 115.355 178.935 ;
        RECT 115.525 178.655 116.375 179.105 ;
        RECT 114.710 178.085 114.915 178.455 ;
        RECT 115.095 178.255 116.215 178.475 ;
        RECT 106.410 177.545 113.530 177.795 ;
        RECT 101.360 177.085 102.180 177.255 ;
        RECT 102.750 177.105 104.020 177.295 ;
        RECT 101.350 176.555 101.680 176.915 ;
        RECT 101.850 176.725 102.180 177.085 ;
        RECT 102.350 176.555 102.585 176.995 ;
        RECT 103.175 176.555 103.510 176.935 ;
        RECT 104.190 176.895 104.805 177.295 ;
        RECT 105.075 177.205 111.820 177.375 ;
        RECT 104.470 176.725 104.805 176.895 ;
        RECT 105.075 176.555 105.375 177.035 ;
        RECT 105.545 176.750 105.805 177.205 ;
        RECT 105.975 176.555 106.235 177.035 ;
        RECT 106.415 176.750 106.675 177.205 ;
        RECT 106.845 176.555 107.095 177.035 ;
        RECT 107.275 176.750 107.535 177.205 ;
        RECT 107.705 176.555 107.955 177.035 ;
        RECT 108.135 176.750 108.395 177.205 ;
        RECT 108.565 176.555 108.810 177.035 ;
        RECT 108.980 176.750 109.255 177.205 ;
        RECT 109.425 176.555 109.670 177.035 ;
        RECT 109.840 176.750 110.100 177.205 ;
        RECT 110.270 176.555 110.530 177.035 ;
        RECT 110.700 176.750 110.960 177.205 ;
        RECT 111.130 176.555 111.390 177.035 ;
        RECT 111.560 176.750 111.820 177.205 ;
        RECT 111.990 176.555 112.250 177.115 ;
        RECT 112.420 176.735 112.670 177.545 ;
        RECT 112.850 176.555 113.110 177.080 ;
        RECT 113.280 176.735 113.530 177.545 ;
        RECT 113.700 177.235 114.015 177.795 ;
        RECT 114.195 177.465 114.455 177.920 ;
        RECT 114.705 177.915 114.915 178.085 ;
        RECT 114.710 177.870 114.915 177.915 ;
        RECT 114.710 177.495 115.295 177.870 ;
        RECT 115.465 177.480 115.875 178.085 ;
        RECT 116.045 177.800 116.215 178.255 ;
        RECT 116.045 177.310 116.375 177.800 ;
        RECT 114.200 177.105 115.355 177.295 ;
        RECT 113.710 176.555 114.015 177.065 ;
        RECT 114.200 176.965 114.475 177.105 ;
        RECT 115.145 176.935 115.355 177.105 ;
        RECT 115.525 177.105 116.375 177.310 ;
        RECT 114.645 176.555 114.975 176.935 ;
        RECT 115.525 176.725 115.855 177.105 ;
        RECT 116.045 176.555 116.375 176.935 ;
        RECT 116.545 176.725 116.790 178.935 ;
        RECT 116.975 178.105 117.230 179.105 ;
        RECT 117.405 177.940 117.695 179.105 ;
        RECT 118.030 178.140 118.360 178.935 ;
        RECT 118.530 178.320 118.770 179.105 ;
        RECT 119.330 178.515 120.085 178.935 ;
        RECT 118.940 178.345 120.405 178.515 ;
        RECT 118.940 178.140 119.110 178.345 ;
        RECT 118.030 177.965 119.110 178.140 ;
        RECT 118.325 177.915 119.110 177.965 ;
        RECT 117.865 177.445 118.125 177.795 ;
        RECT 116.975 176.555 117.215 177.355 ;
        RECT 117.405 176.555 117.695 177.280 ;
        RECT 118.325 177.275 118.495 177.915 ;
        RECT 119.280 177.745 119.570 178.175 ;
        RECT 118.665 177.545 119.010 177.745 ;
        RECT 119.180 177.545 119.570 177.745 ;
        RECT 119.760 177.755 120.065 178.175 ;
        RECT 120.235 178.095 120.405 178.345 ;
        RECT 120.575 178.265 120.905 179.105 ;
        RECT 121.075 178.515 121.325 178.935 ;
        RECT 121.495 178.685 121.835 179.105 ;
        RECT 121.075 178.345 121.835 178.515 ;
        RECT 120.235 177.925 121.195 178.095 ;
        RECT 121.025 177.755 121.195 177.925 ;
        RECT 119.760 177.545 120.245 177.755 ;
        RECT 120.415 177.545 120.855 177.755 ;
        RECT 121.025 177.545 121.355 177.755 ;
        RECT 121.525 177.375 121.835 178.345 ;
        RECT 122.475 178.295 122.770 179.105 ;
        RECT 122.950 177.795 123.195 178.935 ;
        RECT 123.370 178.295 123.630 179.105 ;
        RECT 124.230 179.100 130.505 179.105 ;
        RECT 123.810 177.795 124.060 178.930 ;
        RECT 124.230 178.305 124.490 179.100 ;
        RECT 124.660 178.205 124.920 178.930 ;
        RECT 125.090 178.375 125.350 179.100 ;
        RECT 125.520 178.205 125.780 178.930 ;
        RECT 125.950 178.375 126.210 179.100 ;
        RECT 126.380 178.205 126.640 178.930 ;
        RECT 126.810 178.375 127.070 179.100 ;
        RECT 127.240 178.205 127.500 178.930 ;
        RECT 127.670 178.375 127.915 179.100 ;
        RECT 128.085 178.205 128.345 178.930 ;
        RECT 128.530 178.375 128.775 179.100 ;
        RECT 128.945 178.205 129.205 178.930 ;
        RECT 129.390 178.375 129.635 179.100 ;
        RECT 129.805 178.205 130.065 178.930 ;
        RECT 130.250 178.375 130.505 179.100 ;
        RECT 124.660 178.190 130.065 178.205 ;
        RECT 130.675 178.190 130.965 178.930 ;
        RECT 131.135 178.360 131.405 179.105 ;
        RECT 124.660 177.965 131.405 178.190 ;
        RECT 131.665 177.965 131.995 179.105 ;
        RECT 132.165 178.475 132.520 178.935 ;
        RECT 132.690 178.645 133.265 179.105 ;
        RECT 133.435 178.475 133.765 178.935 ;
        RECT 132.165 178.305 133.765 178.475 ;
        RECT 133.965 178.305 134.220 179.105 ;
        RECT 134.905 178.515 135.145 178.905 ;
        RECT 135.315 178.695 135.665 179.105 ;
        RECT 132.165 177.965 132.440 178.305 ;
        RECT 117.950 177.105 118.495 177.275 ;
        RECT 118.865 177.205 120.565 177.375 ;
        RECT 118.865 177.115 119.250 177.205 ;
        RECT 117.950 176.725 118.280 177.105 ;
        RECT 118.450 176.765 119.635 176.935 ;
        RECT 119.895 176.555 120.065 177.025 ;
        RECT 120.235 176.740 120.565 177.205 ;
        RECT 120.735 176.555 120.905 177.375 ;
        RECT 121.075 177.205 121.835 177.375 ;
        RECT 122.465 177.235 122.780 177.795 ;
        RECT 122.950 177.545 130.070 177.795 ;
        RECT 121.075 176.735 121.405 177.205 ;
        RECT 121.575 176.555 121.745 177.035 ;
        RECT 122.465 176.555 122.770 177.065 ;
        RECT 122.950 176.735 123.200 177.545 ;
        RECT 123.370 176.555 123.630 177.080 ;
        RECT 123.810 176.735 124.060 177.545 ;
        RECT 130.240 177.375 131.405 177.965 ;
        RECT 132.620 177.745 132.810 178.125 ;
        RECT 131.665 177.545 132.810 177.745 ;
        RECT 132.990 177.375 133.270 178.305 ;
        RECT 134.390 178.135 134.690 178.330 ;
        RECT 134.905 178.315 135.655 178.515 ;
        RECT 133.440 177.965 134.690 178.135 ;
        RECT 133.440 177.545 133.770 177.965 ;
        RECT 134.000 177.465 134.345 177.795 ;
        RECT 124.660 177.205 131.405 177.375 ;
        RECT 124.230 176.555 124.490 177.115 ;
        RECT 124.660 176.750 124.920 177.205 ;
        RECT 125.090 176.555 125.350 177.035 ;
        RECT 125.520 176.750 125.780 177.205 ;
        RECT 125.950 176.555 126.210 177.035 ;
        RECT 126.380 176.750 126.640 177.205 ;
        RECT 126.810 176.555 127.055 177.035 ;
        RECT 127.225 176.750 127.500 177.205 ;
        RECT 127.670 176.555 127.915 177.035 ;
        RECT 128.085 176.750 128.345 177.205 ;
        RECT 128.525 176.555 128.775 177.035 ;
        RECT 128.945 176.750 129.205 177.205 ;
        RECT 129.385 176.555 129.635 177.035 ;
        RECT 129.805 176.750 130.065 177.205 ;
        RECT 130.245 176.555 130.505 177.035 ;
        RECT 130.675 176.750 130.935 177.205 ;
        RECT 131.665 177.165 132.775 177.375 ;
        RECT 131.105 176.555 131.405 177.035 ;
        RECT 131.665 176.725 132.015 177.165 ;
        RECT 132.185 176.555 132.355 176.995 ;
        RECT 132.525 176.935 132.775 177.165 ;
        RECT 132.945 177.275 133.270 177.375 ;
        RECT 132.945 177.105 133.275 177.275 ;
        RECT 133.445 176.935 133.720 177.375 ;
        RECT 134.520 177.310 134.690 177.965 ;
        RECT 132.525 176.725 133.720 176.935 ;
        RECT 133.955 176.555 134.285 177.295 ;
        RECT 134.455 176.980 134.690 177.310 ;
        RECT 134.905 176.795 135.135 178.135 ;
        RECT 135.315 177.635 135.655 178.315 ;
        RECT 135.835 177.815 136.165 178.925 ;
        RECT 136.335 178.455 136.515 178.925 ;
        RECT 136.685 178.625 137.015 179.105 ;
        RECT 137.190 178.455 137.360 178.925 ;
        RECT 136.335 178.255 137.360 178.455 ;
        RECT 135.315 176.735 135.545 177.635 ;
        RECT 135.835 177.515 136.380 177.815 ;
        RECT 135.745 176.555 135.990 177.335 ;
        RECT 136.160 177.285 136.380 177.515 ;
        RECT 136.550 177.465 136.975 178.085 ;
        RECT 137.170 177.465 137.430 178.085 ;
        RECT 137.625 177.965 137.910 179.105 ;
        RECT 137.640 177.285 137.900 177.795 ;
        RECT 136.160 177.095 137.900 177.285 ;
        RECT 136.160 176.735 136.590 177.095 ;
        RECT 137.170 176.555 137.900 176.925 ;
        RECT 138.100 176.735 138.380 178.925 ;
        RECT 138.565 178.015 139.775 179.105 ;
        RECT 138.565 177.475 139.085 178.015 ;
        RECT 139.255 177.305 139.775 177.845 ;
        RECT 138.565 176.555 139.775 177.305 ;
        RECT 27.160 176.385 139.860 176.555 ;
        RECT 27.245 175.635 28.455 176.385 ;
        RECT 28.625 175.840 33.970 176.385 ;
        RECT 34.145 175.840 39.490 176.385 ;
        RECT 27.245 175.095 27.765 175.635 ;
        RECT 27.935 174.925 28.455 175.465 ;
        RECT 30.210 175.010 30.550 175.840 ;
        RECT 27.245 173.835 28.455 174.925 ;
        RECT 32.030 174.270 32.380 175.520 ;
        RECT 35.730 175.010 36.070 175.840 ;
        RECT 39.665 175.615 41.335 176.385 ;
        RECT 41.510 175.880 41.845 176.385 ;
        RECT 42.015 175.815 42.255 176.190 ;
        RECT 42.535 176.055 42.705 176.200 ;
        RECT 42.535 175.860 42.910 176.055 ;
        RECT 43.270 175.890 43.665 176.385 ;
        RECT 37.550 174.270 37.900 175.520 ;
        RECT 39.665 175.095 40.415 175.615 ;
        RECT 40.585 174.925 41.335 175.445 ;
        RECT 28.625 173.835 33.970 174.270 ;
        RECT 34.145 173.835 39.490 174.270 ;
        RECT 39.665 173.835 41.335 174.925 ;
        RECT 41.565 174.855 41.865 175.705 ;
        RECT 42.035 175.665 42.255 175.815 ;
        RECT 42.035 175.335 42.570 175.665 ;
        RECT 42.740 175.525 42.910 175.860 ;
        RECT 43.835 175.695 44.075 176.215 ;
        RECT 44.270 175.985 44.605 176.385 ;
        RECT 44.775 175.815 44.980 176.215 ;
        RECT 45.190 175.905 45.465 176.385 ;
        RECT 45.675 175.885 45.935 176.215 ;
        RECT 42.035 174.685 42.270 175.335 ;
        RECT 42.740 175.165 43.725 175.525 ;
        RECT 41.595 174.455 42.270 174.685 ;
        RECT 42.440 175.145 43.725 175.165 ;
        RECT 42.440 174.995 43.300 175.145 ;
        RECT 43.900 175.025 44.075 175.695 ;
        RECT 41.595 174.025 41.765 174.455 ;
        RECT 41.935 173.835 42.265 174.285 ;
        RECT 42.440 174.050 42.725 174.995 ;
        RECT 43.865 174.890 44.075 175.025 ;
        RECT 42.900 174.515 43.595 174.825 ;
        RECT 42.905 173.835 43.590 174.305 ;
        RECT 43.770 174.105 44.075 174.890 ;
        RECT 44.295 175.645 44.980 175.815 ;
        RECT 44.295 174.615 44.635 175.645 ;
        RECT 44.805 174.975 45.055 175.475 ;
        RECT 45.235 175.145 45.595 175.725 ;
        RECT 45.765 174.975 45.935 175.885 ;
        RECT 46.105 175.635 47.315 176.385 ;
        RECT 47.485 175.925 48.045 176.215 ;
        RECT 48.215 175.925 48.465 176.385 ;
        RECT 46.105 175.095 46.625 175.635 ;
        RECT 44.805 174.805 45.935 174.975 ;
        RECT 46.795 174.925 47.315 175.465 ;
        RECT 44.295 174.440 44.960 174.615 ;
        RECT 44.270 173.835 44.605 174.260 ;
        RECT 44.775 174.035 44.960 174.440 ;
        RECT 45.165 173.835 45.495 174.615 ;
        RECT 45.665 174.035 45.935 174.805 ;
        RECT 46.105 173.835 47.315 174.925 ;
        RECT 47.485 174.555 47.735 175.925 ;
        RECT 49.085 175.755 49.415 176.115 ;
        RECT 49.790 175.985 50.125 176.385 ;
        RECT 50.295 175.815 50.500 176.215 ;
        RECT 50.710 175.905 50.985 176.385 ;
        RECT 51.195 175.885 51.455 176.215 ;
        RECT 48.025 175.565 49.415 175.755 ;
        RECT 49.815 175.645 50.500 175.815 ;
        RECT 48.025 175.475 48.195 175.565 ;
        RECT 47.905 175.145 48.195 175.475 ;
        RECT 48.365 175.145 48.705 175.395 ;
        RECT 48.925 175.145 49.600 175.395 ;
        RECT 48.025 174.895 48.195 175.145 ;
        RECT 48.025 174.725 48.965 174.895 ;
        RECT 49.335 174.785 49.600 175.145 ;
        RECT 47.485 174.005 47.945 174.555 ;
        RECT 48.135 173.835 48.465 174.555 ;
        RECT 48.665 174.175 48.965 174.725 ;
        RECT 49.815 174.615 50.155 175.645 ;
        RECT 50.325 174.975 50.575 175.475 ;
        RECT 50.755 175.145 51.115 175.725 ;
        RECT 51.285 174.975 51.455 175.885 ;
        RECT 51.625 175.635 52.835 176.385 ;
        RECT 53.005 175.660 53.295 176.385 ;
        RECT 53.465 175.840 58.810 176.385 ;
        RECT 51.625 175.095 52.145 175.635 ;
        RECT 50.325 174.805 51.455 174.975 ;
        RECT 52.315 174.925 52.835 175.465 ;
        RECT 55.050 175.010 55.390 175.840 ;
        RECT 58.985 175.585 59.295 176.385 ;
        RECT 59.500 175.585 60.195 176.215 ;
        RECT 60.365 175.585 60.675 176.385 ;
        RECT 60.880 175.585 61.575 176.215 ;
        RECT 49.135 173.835 49.415 174.505 ;
        RECT 49.815 174.440 50.480 174.615 ;
        RECT 49.790 173.835 50.125 174.260 ;
        RECT 50.295 174.035 50.480 174.440 ;
        RECT 50.685 173.835 51.015 174.615 ;
        RECT 51.185 174.035 51.455 174.805 ;
        RECT 51.625 173.835 52.835 174.925 ;
        RECT 53.005 173.835 53.295 175.000 ;
        RECT 56.870 174.270 57.220 175.520 ;
        RECT 58.995 175.145 59.330 175.415 ;
        RECT 59.500 174.985 59.670 175.585 ;
        RECT 59.840 175.145 60.175 175.395 ;
        RECT 60.375 175.145 60.710 175.415 ;
        RECT 60.880 174.985 61.050 175.585 ;
        RECT 61.755 175.575 62.025 176.385 ;
        RECT 62.195 175.575 62.525 176.215 ;
        RECT 62.695 175.575 62.935 176.385 ;
        RECT 63.160 175.645 63.775 176.215 ;
        RECT 63.945 175.875 64.160 176.385 ;
        RECT 64.390 175.875 64.670 176.205 ;
        RECT 64.850 175.875 65.090 176.385 ;
        RECT 61.220 175.145 61.555 175.395 ;
        RECT 61.745 175.145 62.095 175.395 ;
        RECT 53.465 173.835 58.810 174.270 ;
        RECT 58.985 173.835 59.265 174.975 ;
        RECT 59.435 174.005 59.765 174.985 ;
        RECT 59.935 173.835 60.195 174.975 ;
        RECT 60.365 173.835 60.645 174.975 ;
        RECT 60.815 174.005 61.145 174.985 ;
        RECT 62.265 174.975 62.435 175.575 ;
        RECT 62.605 175.145 62.955 175.395 ;
        RECT 61.315 173.835 61.575 174.975 ;
        RECT 61.755 173.835 62.085 174.975 ;
        RECT 62.265 174.805 62.945 174.975 ;
        RECT 62.615 174.020 62.945 174.805 ;
        RECT 63.160 174.625 63.475 175.645 ;
        RECT 63.645 174.975 63.815 175.475 ;
        RECT 64.065 175.145 64.330 175.705 ;
        RECT 64.500 174.975 64.670 175.875 ;
        RECT 65.975 175.835 66.145 176.215 ;
        RECT 66.325 176.005 66.655 176.385 ;
        RECT 64.840 175.145 65.195 175.705 ;
        RECT 65.975 175.665 66.640 175.835 ;
        RECT 66.835 175.710 67.095 176.215 ;
        RECT 65.905 175.115 66.245 175.485 ;
        RECT 66.470 175.410 66.640 175.665 ;
        RECT 66.470 175.080 66.745 175.410 ;
        RECT 63.645 174.805 65.070 174.975 ;
        RECT 66.470 174.935 66.640 175.080 ;
        RECT 63.160 174.005 63.695 174.625 ;
        RECT 63.865 173.835 64.195 174.635 ;
        RECT 64.680 174.630 65.070 174.805 ;
        RECT 65.965 174.765 66.640 174.935 ;
        RECT 66.915 174.910 67.095 175.710 ;
        RECT 67.285 175.655 67.575 176.385 ;
        RECT 67.275 175.145 67.575 175.475 ;
        RECT 67.755 175.455 67.985 176.095 ;
        RECT 68.165 175.835 68.475 176.205 ;
        RECT 68.655 176.015 69.325 176.385 ;
        RECT 68.165 175.635 69.395 175.835 ;
        RECT 67.755 175.145 68.280 175.455 ;
        RECT 68.460 175.145 68.925 175.455 ;
        RECT 69.105 174.965 69.395 175.635 ;
        RECT 65.965 174.005 66.145 174.765 ;
        RECT 66.325 173.835 66.655 174.595 ;
        RECT 66.825 174.005 67.095 174.910 ;
        RECT 67.285 174.725 68.445 174.965 ;
        RECT 67.285 174.015 67.545 174.725 ;
        RECT 67.715 173.835 68.045 174.545 ;
        RECT 68.215 174.015 68.445 174.725 ;
        RECT 68.625 174.745 69.395 174.965 ;
        RECT 68.625 174.015 68.895 174.745 ;
        RECT 69.075 173.835 69.415 174.565 ;
        RECT 69.585 174.015 69.845 176.205 ;
        RECT 70.485 174.005 71.235 176.215 ;
        RECT 71.495 175.835 71.665 176.215 ;
        RECT 71.845 176.005 72.175 176.385 ;
        RECT 71.495 175.665 72.160 175.835 ;
        RECT 72.355 175.710 72.615 176.215 ;
        RECT 71.425 175.115 71.765 175.485 ;
        RECT 71.990 175.410 72.160 175.665 ;
        RECT 71.990 175.080 72.265 175.410 ;
        RECT 71.990 174.935 72.160 175.080 ;
        RECT 71.485 174.765 72.160 174.935 ;
        RECT 72.435 174.910 72.615 175.710 ;
        RECT 72.875 175.835 73.045 176.215 ;
        RECT 73.225 176.005 73.555 176.385 ;
        RECT 72.875 175.665 73.540 175.835 ;
        RECT 73.735 175.710 73.995 176.215 ;
        RECT 72.805 175.115 73.135 175.485 ;
        RECT 73.370 175.410 73.540 175.665 ;
        RECT 73.370 175.080 73.655 175.410 ;
        RECT 73.370 174.935 73.540 175.080 ;
        RECT 71.485 174.005 71.665 174.765 ;
        RECT 71.845 173.835 72.175 174.595 ;
        RECT 72.345 174.005 72.615 174.910 ;
        RECT 72.875 174.765 73.540 174.935 ;
        RECT 73.825 174.910 73.995 175.710 ;
        RECT 72.875 174.005 73.045 174.765 ;
        RECT 73.225 173.835 73.555 174.595 ;
        RECT 73.725 174.005 73.995 174.910 ;
        RECT 74.165 174.005 74.915 176.215 ;
        RECT 75.555 175.885 75.885 176.385 ;
        RECT 76.085 175.815 76.255 176.165 ;
        RECT 76.455 175.985 76.785 176.385 ;
        RECT 76.955 175.815 77.125 176.165 ;
        RECT 77.295 175.985 77.675 176.385 ;
        RECT 75.550 175.145 75.900 175.715 ;
        RECT 76.085 175.645 77.695 175.815 ;
        RECT 77.865 175.710 78.135 176.055 ;
        RECT 77.525 175.475 77.695 175.645 ;
        RECT 76.070 175.025 76.780 175.475 ;
        RECT 76.950 175.145 77.355 175.475 ;
        RECT 77.525 175.145 77.795 175.475 ;
        RECT 75.550 174.685 75.870 174.975 ;
        RECT 76.065 174.855 76.780 175.025 ;
        RECT 77.525 174.975 77.695 175.145 ;
        RECT 77.965 174.975 78.135 175.710 ;
        RECT 78.765 175.660 79.055 176.385 ;
        RECT 79.225 176.005 80.115 176.175 ;
        RECT 79.225 175.450 79.775 175.835 ;
        RECT 79.945 175.280 80.115 176.005 ;
        RECT 79.225 175.210 80.115 175.280 ;
        RECT 80.285 175.680 80.505 176.165 ;
        RECT 80.675 175.845 80.925 176.385 ;
        RECT 81.095 175.735 81.355 176.215 ;
        RECT 80.285 175.255 80.615 175.680 ;
        RECT 79.225 175.185 80.120 175.210 ;
        RECT 79.225 175.170 80.130 175.185 ;
        RECT 79.225 175.155 80.135 175.170 ;
        RECT 79.225 175.150 80.145 175.155 ;
        RECT 79.225 175.140 80.150 175.150 ;
        RECT 79.225 175.130 80.155 175.140 ;
        RECT 79.225 175.125 80.165 175.130 ;
        RECT 79.225 175.115 80.175 175.125 ;
        RECT 79.225 175.110 80.185 175.115 ;
        RECT 76.970 174.805 77.695 174.975 ;
        RECT 76.970 174.685 77.140 174.805 ;
        RECT 75.550 174.515 77.140 174.685 ;
        RECT 75.550 174.055 77.205 174.345 ;
        RECT 77.375 173.835 77.655 174.635 ;
        RECT 77.865 174.005 78.135 174.975 ;
        RECT 78.765 173.835 79.055 175.000 ;
        RECT 79.225 174.660 79.485 175.110 ;
        RECT 79.850 175.105 80.185 175.110 ;
        RECT 79.850 175.100 80.200 175.105 ;
        RECT 79.850 175.090 80.215 175.100 ;
        RECT 79.850 175.085 80.240 175.090 ;
        RECT 80.785 175.085 81.015 175.480 ;
        RECT 79.850 175.080 81.015 175.085 ;
        RECT 79.880 175.045 81.015 175.080 ;
        RECT 79.915 175.020 81.015 175.045 ;
        RECT 79.945 174.990 81.015 175.020 ;
        RECT 79.965 174.960 81.015 174.990 ;
        RECT 79.985 174.930 81.015 174.960 ;
        RECT 80.055 174.920 81.015 174.930 ;
        RECT 80.080 174.910 81.015 174.920 ;
        RECT 80.100 174.895 81.015 174.910 ;
        RECT 80.120 174.880 81.015 174.895 ;
        RECT 80.125 174.870 80.910 174.880 ;
        RECT 80.140 174.835 80.910 174.870 ;
        RECT 79.655 174.515 79.985 174.760 ;
        RECT 80.155 174.585 80.910 174.835 ;
        RECT 81.185 174.705 81.355 175.735 ;
        RECT 81.615 175.835 81.785 176.215 ;
        RECT 81.965 176.005 82.295 176.385 ;
        RECT 81.615 175.665 82.280 175.835 ;
        RECT 82.475 175.710 82.735 176.215 ;
        RECT 81.545 175.115 81.885 175.485 ;
        RECT 82.110 175.410 82.280 175.665 ;
        RECT 82.110 175.080 82.385 175.410 ;
        RECT 82.110 174.935 82.280 175.080 ;
        RECT 79.655 174.490 79.840 174.515 ;
        RECT 79.225 174.390 79.840 174.490 ;
        RECT 79.225 173.835 79.830 174.390 ;
        RECT 80.005 174.005 80.485 174.345 ;
        RECT 80.655 173.835 80.910 174.380 ;
        RECT 81.080 174.005 81.355 174.705 ;
        RECT 81.605 174.765 82.280 174.935 ;
        RECT 82.555 174.910 82.735 175.710 ;
        RECT 83.455 175.835 83.625 176.215 ;
        RECT 83.805 176.005 84.135 176.385 ;
        RECT 83.455 175.665 84.120 175.835 ;
        RECT 84.315 175.710 84.575 176.215 ;
        RECT 83.385 175.115 83.725 175.485 ;
        RECT 83.950 175.410 84.120 175.665 ;
        RECT 83.950 175.080 84.225 175.410 ;
        RECT 83.950 174.935 84.120 175.080 ;
        RECT 81.605 174.005 81.785 174.765 ;
        RECT 81.965 173.835 82.295 174.595 ;
        RECT 82.465 174.005 82.735 174.910 ;
        RECT 83.445 174.765 84.120 174.935 ;
        RECT 84.395 174.910 84.575 175.710 ;
        RECT 84.835 175.735 85.005 176.215 ;
        RECT 85.175 175.905 85.505 176.385 ;
        RECT 85.730 175.965 87.265 176.215 ;
        RECT 85.730 175.735 85.900 175.965 ;
        RECT 84.835 175.565 85.900 175.735 ;
        RECT 86.080 175.395 86.360 175.795 ;
        RECT 84.750 175.185 85.100 175.395 ;
        RECT 85.270 175.195 85.715 175.395 ;
        RECT 85.885 175.195 86.360 175.395 ;
        RECT 86.630 175.395 86.915 175.795 ;
        RECT 87.095 175.735 87.265 175.965 ;
        RECT 87.435 175.905 87.765 176.385 ;
        RECT 87.980 175.885 88.235 176.215 ;
        RECT 88.050 175.805 88.235 175.885 ;
        RECT 87.095 175.565 87.895 175.735 ;
        RECT 86.630 175.195 86.960 175.395 ;
        RECT 87.130 175.365 87.495 175.395 ;
        RECT 87.130 175.195 87.505 175.365 ;
        RECT 87.725 175.015 87.895 175.565 ;
        RECT 83.445 174.005 83.625 174.765 ;
        RECT 83.805 173.835 84.135 174.595 ;
        RECT 84.305 174.005 84.575 174.910 ;
        RECT 84.835 174.845 87.895 175.015 ;
        RECT 84.835 174.005 85.005 174.845 ;
        RECT 88.065 174.685 88.235 175.805 ;
        RECT 88.435 175.655 88.735 176.385 ;
        RECT 88.915 175.475 89.145 176.095 ;
        RECT 89.345 175.825 89.570 176.205 ;
        RECT 89.740 175.995 90.070 176.385 ;
        RECT 90.290 175.985 90.620 176.385 ;
        RECT 89.345 175.645 89.675 175.825 ;
        RECT 90.790 175.815 90.960 176.085 ;
        RECT 91.130 175.875 91.445 176.385 ;
        RECT 91.675 175.875 91.965 176.215 ;
        RECT 92.135 175.875 92.375 176.385 ;
        RECT 92.615 175.915 92.905 176.385 ;
        RECT 88.440 175.145 88.735 175.475 ;
        RECT 88.915 175.145 89.330 175.475 ;
        RECT 89.500 174.975 89.675 175.645 ;
        RECT 89.845 175.145 90.085 175.795 ;
        RECT 90.265 175.645 90.960 175.815 ;
        RECT 88.025 174.675 88.235 174.685 ;
        RECT 85.175 174.175 85.505 174.675 ;
        RECT 85.675 174.435 87.310 174.675 ;
        RECT 85.675 174.345 85.905 174.435 ;
        RECT 86.015 174.175 86.345 174.215 ;
        RECT 85.175 174.005 86.345 174.175 ;
        RECT 86.535 173.835 86.890 174.255 ;
        RECT 87.060 174.005 87.310 174.435 ;
        RECT 87.480 173.835 87.810 174.595 ;
        RECT 87.980 174.005 88.235 174.675 ;
        RECT 88.435 174.615 89.330 174.945 ;
        RECT 89.500 174.785 90.085 174.975 ;
        RECT 88.435 174.445 89.640 174.615 ;
        RECT 88.435 174.015 88.765 174.445 ;
        RECT 88.945 173.835 89.140 174.275 ;
        RECT 89.310 174.015 89.640 174.445 ;
        RECT 89.810 174.015 90.085 174.785 ;
        RECT 90.265 174.635 90.695 175.645 ;
        RECT 90.865 174.975 91.035 175.475 ;
        RECT 91.205 175.145 91.615 175.705 ;
        RECT 91.785 174.975 91.965 175.875 ;
        RECT 93.075 175.745 93.405 176.215 ;
        RECT 93.575 175.915 93.745 176.385 ;
        RECT 93.915 175.745 94.245 176.215 ;
        RECT 93.075 175.735 94.245 175.745 ;
        RECT 92.135 175.365 92.330 175.705 ;
        RECT 92.645 175.565 94.245 175.735 ;
        RECT 94.415 175.565 94.690 176.385 ;
        RECT 94.915 175.915 95.205 176.385 ;
        RECT 95.375 175.745 95.705 176.215 ;
        RECT 95.875 175.915 96.045 176.385 ;
        RECT 96.215 175.745 96.545 176.215 ;
        RECT 95.375 175.735 96.545 175.745 ;
        RECT 94.945 175.565 96.545 175.735 ;
        RECT 96.715 175.565 96.990 176.385 ;
        RECT 97.190 175.630 97.425 175.960 ;
        RECT 97.595 175.645 97.925 176.385 ;
        RECT 98.160 176.005 99.355 176.215 ;
        RECT 92.645 175.365 92.860 175.565 ;
        RECT 92.135 175.195 92.335 175.365 ;
        RECT 92.625 175.195 92.860 175.365 ;
        RECT 93.030 175.195 93.800 175.395 ;
        RECT 93.970 175.195 94.690 175.395 ;
        RECT 92.135 175.145 92.330 175.195 ;
        RECT 92.645 175.025 92.860 175.195 ;
        RECT 94.945 175.025 95.160 175.565 ;
        RECT 95.330 175.195 96.100 175.395 ;
        RECT 96.270 175.195 96.990 175.395 ;
        RECT 90.865 174.805 92.325 174.975 ;
        RECT 92.645 174.805 93.405 175.025 ;
        RECT 90.265 174.465 91.040 174.635 ;
        RECT 90.370 173.835 90.540 174.295 ;
        RECT 90.710 174.005 91.040 174.465 ;
        RECT 91.210 173.835 91.380 174.635 ;
        RECT 91.965 174.630 92.325 174.805 ;
        RECT 92.605 174.175 92.905 174.635 ;
        RECT 93.075 174.345 93.405 174.805 ;
        RECT 93.575 174.805 94.690 175.015 ;
        RECT 94.945 174.805 95.705 175.025 ;
        RECT 93.575 174.175 93.745 174.805 ;
        RECT 92.605 174.005 93.745 174.175 ;
        RECT 93.915 173.835 94.245 174.635 ;
        RECT 94.415 174.005 94.690 174.805 ;
        RECT 94.905 174.175 95.205 174.635 ;
        RECT 95.375 174.345 95.705 174.805 ;
        RECT 95.875 174.805 96.990 175.015 ;
        RECT 95.875 174.175 96.045 174.805 ;
        RECT 94.905 174.005 96.045 174.175 ;
        RECT 96.215 173.835 96.545 174.635 ;
        RECT 96.715 174.005 96.990 174.805 ;
        RECT 97.190 174.975 97.360 175.630 ;
        RECT 98.160 175.565 98.435 176.005 ;
        RECT 98.605 175.665 98.935 175.835 ;
        RECT 98.610 175.565 98.935 175.665 ;
        RECT 99.105 175.775 99.355 176.005 ;
        RECT 99.525 175.945 99.695 176.385 ;
        RECT 99.865 175.775 100.215 176.215 ;
        RECT 99.105 175.565 100.215 175.775 ;
        RECT 101.315 175.660 101.645 176.170 ;
        RECT 101.815 175.985 102.145 176.385 ;
        RECT 103.195 175.815 103.525 176.155 ;
        RECT 103.695 175.985 104.025 176.385 ;
        RECT 97.535 175.145 97.880 175.475 ;
        RECT 98.110 174.975 98.440 175.395 ;
        RECT 97.190 174.805 98.440 174.975 ;
        RECT 97.190 174.610 97.490 174.805 ;
        RECT 98.610 174.635 98.890 175.565 ;
        RECT 99.070 175.195 100.215 175.395 ;
        RECT 99.070 174.815 99.260 175.195 ;
        RECT 99.440 174.635 99.715 174.975 ;
        RECT 97.660 173.835 97.915 174.635 ;
        RECT 98.115 174.465 99.715 174.635 ;
        RECT 98.115 174.005 98.445 174.465 ;
        RECT 98.615 173.835 99.190 174.295 ;
        RECT 99.360 174.005 99.715 174.465 ;
        RECT 99.885 173.835 100.215 174.975 ;
        RECT 101.315 174.895 101.505 175.660 ;
        RECT 101.815 175.645 104.180 175.815 ;
        RECT 104.525 175.660 104.815 176.385 ;
        RECT 104.985 175.885 105.285 176.215 ;
        RECT 105.455 175.905 105.730 176.385 ;
        RECT 101.815 175.475 101.985 175.645 ;
        RECT 101.675 175.145 101.985 175.475 ;
        RECT 102.155 175.145 102.460 175.475 ;
        RECT 101.315 174.045 101.645 174.895 ;
        RECT 101.815 173.835 102.065 174.975 ;
        RECT 102.245 174.815 102.460 175.145 ;
        RECT 102.635 174.815 102.920 175.475 ;
        RECT 103.115 174.815 103.380 175.475 ;
        RECT 103.595 174.815 103.840 175.475 ;
        RECT 104.010 174.645 104.180 175.645 ;
        RECT 102.255 174.475 103.545 174.645 ;
        RECT 102.255 174.055 102.505 174.475 ;
        RECT 102.735 173.835 103.065 174.305 ;
        RECT 103.295 174.055 103.545 174.475 ;
        RECT 103.725 174.475 104.180 174.645 ;
        RECT 103.725 174.045 104.055 174.475 ;
        RECT 104.525 173.835 104.815 175.000 ;
        RECT 104.985 174.975 105.155 175.885 ;
        RECT 105.910 175.735 106.205 176.125 ;
        RECT 106.375 175.905 106.630 176.385 ;
        RECT 106.805 175.735 107.065 176.125 ;
        RECT 107.235 175.905 107.515 176.385 ;
        RECT 105.325 175.145 105.675 175.715 ;
        RECT 105.910 175.565 107.560 175.735 ;
        RECT 107.750 175.565 108.045 176.385 ;
        RECT 108.215 175.835 108.435 176.215 ;
        RECT 108.605 176.025 109.455 176.385 ;
        RECT 105.845 175.225 106.985 175.395 ;
        RECT 105.845 174.975 106.015 175.225 ;
        RECT 107.155 175.055 107.560 175.565 ;
        RECT 104.985 174.805 106.015 174.975 ;
        RECT 106.805 174.885 107.560 175.055 ;
        RECT 104.985 174.005 105.295 174.805 ;
        RECT 106.805 174.635 107.065 174.885 ;
        RECT 105.465 173.835 105.775 174.635 ;
        RECT 105.945 174.465 107.065 174.635 ;
        RECT 105.945 174.005 106.205 174.465 ;
        RECT 106.375 173.835 106.630 174.295 ;
        RECT 106.805 174.005 107.065 174.465 ;
        RECT 107.235 173.835 107.520 174.705 ;
        RECT 107.750 173.835 108.045 174.980 ;
        RECT 108.215 174.135 108.445 175.835 ;
        RECT 109.935 175.775 110.265 176.195 ;
        RECT 110.470 175.945 110.745 176.385 ;
        RECT 110.915 175.775 111.245 176.195 ;
        RECT 111.425 175.875 111.730 176.385 ;
        RECT 108.660 175.595 111.245 175.775 ;
        RECT 108.660 174.980 108.970 175.595 ;
        RECT 109.140 175.195 109.470 175.425 ;
        RECT 109.640 175.195 110.110 175.425 ;
        RECT 110.280 175.365 110.730 175.425 ;
        RECT 110.280 175.195 110.735 175.365 ;
        RECT 110.920 175.195 111.255 175.425 ;
        RECT 111.425 175.145 111.740 175.705 ;
        RECT 111.910 175.395 112.160 176.205 ;
        RECT 112.330 175.860 112.590 176.385 ;
        RECT 112.770 175.395 113.020 176.205 ;
        RECT 113.190 175.825 113.450 176.385 ;
        RECT 113.620 175.735 113.880 176.190 ;
        RECT 114.050 175.905 114.310 176.385 ;
        RECT 114.480 175.735 114.740 176.190 ;
        RECT 114.910 175.905 115.170 176.385 ;
        RECT 115.340 175.735 115.600 176.190 ;
        RECT 115.770 175.905 116.015 176.385 ;
        RECT 116.185 175.735 116.460 176.190 ;
        RECT 116.630 175.905 116.875 176.385 ;
        RECT 117.045 175.735 117.305 176.190 ;
        RECT 117.485 175.905 117.735 176.385 ;
        RECT 117.905 175.735 118.165 176.190 ;
        RECT 118.345 175.905 118.595 176.385 ;
        RECT 118.765 175.735 119.025 176.190 ;
        RECT 119.205 175.905 119.465 176.385 ;
        RECT 119.635 175.735 119.895 176.190 ;
        RECT 120.065 175.905 120.365 176.385 ;
        RECT 120.715 175.905 121.015 176.385 ;
        RECT 121.185 175.735 121.445 176.190 ;
        RECT 121.615 175.905 121.875 176.385 ;
        RECT 122.055 175.735 122.315 176.190 ;
        RECT 122.485 175.905 122.735 176.385 ;
        RECT 122.915 175.735 123.175 176.190 ;
        RECT 123.345 175.905 123.595 176.385 ;
        RECT 123.775 175.735 124.035 176.190 ;
        RECT 124.205 175.905 124.450 176.385 ;
        RECT 124.620 175.735 124.895 176.190 ;
        RECT 125.065 175.905 125.310 176.385 ;
        RECT 125.480 175.735 125.740 176.190 ;
        RECT 125.910 175.905 126.170 176.385 ;
        RECT 126.340 175.735 126.600 176.190 ;
        RECT 126.770 175.905 127.030 176.385 ;
        RECT 127.200 175.735 127.460 176.190 ;
        RECT 127.630 175.825 127.890 176.385 ;
        RECT 113.620 175.565 120.365 175.735 ;
        RECT 111.910 175.145 119.030 175.395 ;
        RECT 119.200 175.365 120.365 175.565 ;
        RECT 120.715 175.565 127.460 175.735 ;
        RECT 119.200 175.195 120.395 175.365 ;
        RECT 108.660 174.810 111.245 174.980 ;
        RECT 108.660 173.835 108.915 174.640 ;
        RECT 109.115 174.450 110.455 174.630 ;
        RECT 109.115 174.005 109.445 174.450 ;
        RECT 109.615 173.835 109.890 174.280 ;
        RECT 110.125 174.005 110.455 174.450 ;
        RECT 110.915 174.145 111.245 174.810 ;
        RECT 111.435 173.835 111.730 174.645 ;
        RECT 111.910 174.005 112.155 175.145 ;
        RECT 112.330 173.835 112.590 174.645 ;
        RECT 112.770 174.010 113.020 175.145 ;
        RECT 119.200 174.975 120.365 175.195 ;
        RECT 113.620 174.750 120.365 174.975 ;
        RECT 120.715 174.975 121.880 175.565 ;
        RECT 128.060 175.395 128.310 176.205 ;
        RECT 128.490 175.860 128.750 176.385 ;
        RECT 128.920 175.395 129.170 176.205 ;
        RECT 129.350 175.875 129.655 176.385 ;
        RECT 122.050 175.145 129.170 175.395 ;
        RECT 129.340 175.145 129.655 175.705 ;
        RECT 130.285 175.660 130.575 176.385 ;
        RECT 130.750 175.755 131.085 176.215 ;
        RECT 131.255 175.925 131.450 176.385 ;
        RECT 131.695 176.005 133.720 176.215 ;
        RECT 130.750 175.565 131.440 175.755 ;
        RECT 131.695 175.565 131.945 176.005 ;
        RECT 132.115 175.565 133.300 175.835 ;
        RECT 133.470 175.755 133.720 176.005 ;
        RECT 133.890 175.925 134.060 176.385 ;
        RECT 134.230 175.755 134.560 176.215 ;
        RECT 134.730 175.925 134.970 176.385 ;
        RECT 135.180 175.755 135.510 176.215 ;
        RECT 133.470 175.565 135.510 175.755 ;
        RECT 136.270 175.645 136.605 176.385 ;
        RECT 131.270 175.395 131.440 175.565 ;
        RECT 130.770 175.195 131.100 175.395 ;
        RECT 131.270 175.195 132.865 175.395 ;
        RECT 120.715 174.750 127.460 174.975 ;
        RECT 113.620 174.735 119.025 174.750 ;
        RECT 113.190 173.840 113.450 174.635 ;
        RECT 113.620 174.010 113.880 174.735 ;
        RECT 114.050 173.840 114.310 174.565 ;
        RECT 114.480 174.010 114.740 174.735 ;
        RECT 114.910 173.840 115.170 174.565 ;
        RECT 115.340 174.010 115.600 174.735 ;
        RECT 115.770 173.840 116.030 174.565 ;
        RECT 116.200 174.010 116.460 174.735 ;
        RECT 116.630 173.840 116.875 174.565 ;
        RECT 117.045 174.010 117.305 174.735 ;
        RECT 117.490 173.840 117.735 174.565 ;
        RECT 117.905 174.010 118.165 174.735 ;
        RECT 118.350 173.840 118.595 174.565 ;
        RECT 118.765 174.010 119.025 174.735 ;
        RECT 119.210 173.840 119.465 174.565 ;
        RECT 119.635 174.010 119.925 174.750 ;
        RECT 113.190 173.835 119.465 173.840 ;
        RECT 120.095 173.835 120.365 174.580 ;
        RECT 120.715 173.835 120.985 174.580 ;
        RECT 121.155 174.010 121.445 174.750 ;
        RECT 122.055 174.735 127.460 174.750 ;
        RECT 121.615 173.840 121.870 174.565 ;
        RECT 122.055 174.010 122.315 174.735 ;
        RECT 122.485 173.840 122.730 174.565 ;
        RECT 122.915 174.010 123.175 174.735 ;
        RECT 123.345 173.840 123.590 174.565 ;
        RECT 123.775 174.010 124.035 174.735 ;
        RECT 124.205 173.840 124.450 174.565 ;
        RECT 124.620 174.010 124.880 174.735 ;
        RECT 125.050 173.840 125.310 174.565 ;
        RECT 125.480 174.010 125.740 174.735 ;
        RECT 125.910 173.840 126.170 174.565 ;
        RECT 126.340 174.010 126.600 174.735 ;
        RECT 126.770 173.840 127.030 174.565 ;
        RECT 127.200 174.010 127.460 174.735 ;
        RECT 127.630 173.840 127.890 174.635 ;
        RECT 128.060 174.010 128.310 175.145 ;
        RECT 121.615 173.835 127.890 173.840 ;
        RECT 128.490 173.835 128.750 174.645 ;
        RECT 128.925 174.005 129.170 175.145 ;
        RECT 131.270 175.025 131.440 175.195 ;
        RECT 133.035 175.025 133.300 175.565 ;
        RECT 136.775 175.475 136.990 176.170 ;
        RECT 137.180 175.645 137.530 176.170 ;
        RECT 137.700 175.645 138.395 176.215 ;
        RECT 137.325 175.475 137.530 175.645 ;
        RECT 133.815 175.195 135.600 175.395 ;
        RECT 136.290 175.145 136.575 175.475 ;
        RECT 136.775 175.145 137.155 175.475 ;
        RECT 137.325 175.145 137.635 175.475 ;
        RECT 129.350 173.835 129.645 174.645 ;
        RECT 130.285 173.835 130.575 175.000 ;
        RECT 130.750 174.805 131.440 175.025 ;
        RECT 130.750 174.005 131.085 174.805 ;
        RECT 131.630 174.635 131.945 175.025 ;
        RECT 131.255 173.835 131.945 174.635 ;
        RECT 132.115 174.805 134.980 175.025 ;
        RECT 137.805 174.975 137.975 175.645 ;
        RECT 138.565 175.635 139.775 176.385 ;
        RECT 132.115 174.005 132.445 174.805 ;
        RECT 132.615 173.835 132.785 174.635 ;
        RECT 132.955 174.005 133.300 174.805 ;
        RECT 133.470 173.835 133.640 174.635 ;
        RECT 133.810 174.005 134.140 174.805 ;
        RECT 134.310 173.835 134.480 174.635 ;
        RECT 134.650 174.005 134.980 174.805 ;
        RECT 135.180 173.835 135.510 174.975 ;
        RECT 136.265 173.835 136.525 174.975 ;
        RECT 136.695 174.805 137.975 174.975 ;
        RECT 138.155 174.805 138.395 175.475 ;
        RECT 138.565 174.925 139.085 175.465 ;
        RECT 139.255 175.095 139.775 175.635 ;
        RECT 136.695 174.005 137.025 174.805 ;
        RECT 137.195 173.835 137.365 174.635 ;
        RECT 137.565 174.005 137.895 174.805 ;
        RECT 138.095 173.835 138.375 174.635 ;
        RECT 138.565 173.835 139.775 174.925 ;
        RECT 27.160 173.665 139.860 173.835 ;
        RECT 27.245 172.575 28.455 173.665 ;
        RECT 28.625 173.230 33.970 173.665 ;
        RECT 34.145 173.230 39.490 173.665 ;
        RECT 27.245 171.865 27.765 172.405 ;
        RECT 27.935 172.035 28.455 172.575 ;
        RECT 27.245 171.115 28.455 171.865 ;
        RECT 30.210 171.660 30.550 172.490 ;
        RECT 32.030 171.980 32.380 173.230 ;
        RECT 35.730 171.660 36.070 172.490 ;
        RECT 37.550 171.980 37.900 173.230 ;
        RECT 40.125 172.500 40.415 173.665 ;
        RECT 40.585 173.230 45.930 173.665 ;
        RECT 46.105 173.230 51.450 173.665 ;
        RECT 51.625 173.230 56.970 173.665 ;
        RECT 28.625 171.115 33.970 171.660 ;
        RECT 34.145 171.115 39.490 171.660 ;
        RECT 40.125 171.115 40.415 171.840 ;
        RECT 42.170 171.660 42.510 172.490 ;
        RECT 43.990 171.980 44.340 173.230 ;
        RECT 47.690 171.660 48.030 172.490 ;
        RECT 49.510 171.980 49.860 173.230 ;
        RECT 53.210 171.660 53.550 172.490 ;
        RECT 55.030 171.980 55.380 173.230 ;
        RECT 57.145 172.575 58.355 173.665 ;
        RECT 57.145 171.865 57.665 172.405 ;
        RECT 57.835 172.035 58.355 172.575 ;
        RECT 58.545 172.775 58.805 173.485 ;
        RECT 58.975 172.955 59.305 173.665 ;
        RECT 59.475 172.775 59.705 173.485 ;
        RECT 58.545 172.535 59.705 172.775 ;
        RECT 59.885 172.755 60.155 173.485 ;
        RECT 60.335 172.935 60.675 173.665 ;
        RECT 59.885 172.535 60.655 172.755 ;
        RECT 58.535 172.025 58.835 172.355 ;
        RECT 59.015 172.045 59.540 172.355 ;
        RECT 59.720 172.045 60.185 172.355 ;
        RECT 40.585 171.115 45.930 171.660 ;
        RECT 46.105 171.115 51.450 171.660 ;
        RECT 51.625 171.115 56.970 171.660 ;
        RECT 57.145 171.115 58.355 171.865 ;
        RECT 58.545 171.115 58.835 171.845 ;
        RECT 59.015 171.405 59.245 172.045 ;
        RECT 60.365 171.865 60.655 172.535 ;
        RECT 59.425 171.665 60.655 171.865 ;
        RECT 59.425 171.295 59.735 171.665 ;
        RECT 59.915 171.115 60.585 171.485 ;
        RECT 60.845 171.295 61.105 173.485 ;
        RECT 61.295 173.055 61.625 173.485 ;
        RECT 61.805 173.225 62.000 173.665 ;
        RECT 62.170 173.055 62.500 173.485 ;
        RECT 61.295 172.885 62.500 173.055 ;
        RECT 61.295 172.555 62.190 172.885 ;
        RECT 62.670 172.715 62.945 173.485 ;
        RECT 62.360 172.525 62.945 172.715 ;
        RECT 64.055 173.055 64.385 173.485 ;
        RECT 64.565 173.225 64.760 173.665 ;
        RECT 64.930 173.055 65.260 173.485 ;
        RECT 64.055 172.885 65.260 173.055 ;
        RECT 64.055 172.555 64.950 172.885 ;
        RECT 65.430 172.715 65.705 173.485 ;
        RECT 65.120 172.525 65.705 172.715 ;
        RECT 61.300 172.025 61.595 172.355 ;
        RECT 61.775 172.025 62.190 172.355 ;
        RECT 61.295 171.115 61.595 171.845 ;
        RECT 61.775 171.405 62.005 172.025 ;
        RECT 62.360 171.855 62.535 172.525 ;
        RECT 62.205 171.675 62.535 171.855 ;
        RECT 62.705 171.705 62.945 172.355 ;
        RECT 64.060 172.025 64.355 172.355 ;
        RECT 64.535 172.025 64.950 172.355 ;
        RECT 62.205 171.295 62.430 171.675 ;
        RECT 62.600 171.115 62.930 171.505 ;
        RECT 64.055 171.115 64.355 171.845 ;
        RECT 64.535 171.405 64.765 172.025 ;
        RECT 65.120 171.855 65.295 172.525 ;
        RECT 65.885 172.500 66.175 173.665 ;
        RECT 66.345 172.485 66.665 173.665 ;
        RECT 66.835 172.645 67.035 173.435 ;
        RECT 67.360 172.835 67.745 173.495 ;
        RECT 68.140 172.905 68.925 173.665 ;
        RECT 67.335 172.735 67.745 172.835 ;
        RECT 66.835 172.475 67.165 172.645 ;
        RECT 67.335 172.525 68.945 172.735 ;
        RECT 66.985 172.355 67.165 172.475 ;
        RECT 64.965 171.675 65.295 171.855 ;
        RECT 65.465 171.705 65.705 172.355 ;
        RECT 66.345 172.105 66.810 172.305 ;
        RECT 66.985 172.105 67.315 172.355 ;
        RECT 67.485 172.305 67.950 172.355 ;
        RECT 67.485 172.135 67.955 172.305 ;
        RECT 67.485 172.105 67.950 172.135 ;
        RECT 68.145 172.105 68.500 172.355 ;
        RECT 68.670 171.925 68.945 172.525 ;
        RECT 64.965 171.295 65.190 171.675 ;
        RECT 65.360 171.115 65.690 171.505 ;
        RECT 65.885 171.115 66.175 171.840 ;
        RECT 66.345 171.725 67.525 171.895 ;
        RECT 66.345 171.310 66.685 171.725 ;
        RECT 66.855 171.115 67.025 171.555 ;
        RECT 67.195 171.505 67.525 171.725 ;
        RECT 67.695 171.745 68.945 171.925 ;
        RECT 67.695 171.675 68.060 171.745 ;
        RECT 67.195 171.325 68.445 171.505 ;
        RECT 68.715 171.115 68.885 171.575 ;
        RECT 69.115 171.395 69.395 173.495 ;
        RECT 69.565 172.485 69.885 173.665 ;
        RECT 70.055 172.645 70.255 173.435 ;
        RECT 70.580 172.835 70.965 173.495 ;
        RECT 71.360 172.905 72.145 173.665 ;
        RECT 70.555 172.735 70.965 172.835 ;
        RECT 70.055 172.475 70.385 172.645 ;
        RECT 70.555 172.525 72.165 172.735 ;
        RECT 70.205 172.355 70.385 172.475 ;
        RECT 69.565 172.105 70.030 172.305 ;
        RECT 70.205 172.105 70.535 172.355 ;
        RECT 70.705 172.305 71.170 172.355 ;
        RECT 70.705 172.135 71.175 172.305 ;
        RECT 70.705 172.105 71.170 172.135 ;
        RECT 71.365 172.105 71.720 172.355 ;
        RECT 71.890 171.925 72.165 172.525 ;
        RECT 69.565 171.725 70.745 171.895 ;
        RECT 69.565 171.310 69.905 171.725 ;
        RECT 70.075 171.115 70.245 171.555 ;
        RECT 70.415 171.505 70.745 171.725 ;
        RECT 70.915 171.745 72.165 171.925 ;
        RECT 70.915 171.675 71.280 171.745 ;
        RECT 70.415 171.325 71.665 171.505 ;
        RECT 71.935 171.115 72.105 171.575 ;
        RECT 72.335 171.395 72.615 173.495 ;
        RECT 73.245 173.110 73.850 173.665 ;
        RECT 74.025 173.155 74.505 173.495 ;
        RECT 74.675 173.120 74.930 173.665 ;
        RECT 73.245 173.010 73.860 173.110 ;
        RECT 73.675 172.985 73.860 173.010 ;
        RECT 73.245 172.390 73.505 172.840 ;
        RECT 73.675 172.740 74.005 172.985 ;
        RECT 74.175 172.665 74.930 172.915 ;
        RECT 75.100 172.795 75.375 173.495 ;
        RECT 74.160 172.630 74.930 172.665 ;
        RECT 74.145 172.620 74.930 172.630 ;
        RECT 74.140 172.605 75.035 172.620 ;
        RECT 74.120 172.590 75.035 172.605 ;
        RECT 74.100 172.580 75.035 172.590 ;
        RECT 74.075 172.570 75.035 172.580 ;
        RECT 74.005 172.540 75.035 172.570 ;
        RECT 73.985 172.510 75.035 172.540 ;
        RECT 73.965 172.480 75.035 172.510 ;
        RECT 73.935 172.455 75.035 172.480 ;
        RECT 73.900 172.420 75.035 172.455 ;
        RECT 73.870 172.415 75.035 172.420 ;
        RECT 73.870 172.410 74.260 172.415 ;
        RECT 73.870 172.400 74.235 172.410 ;
        RECT 73.870 172.395 74.220 172.400 ;
        RECT 73.870 172.390 74.205 172.395 ;
        RECT 73.245 172.385 74.205 172.390 ;
        RECT 73.245 172.375 74.195 172.385 ;
        RECT 73.245 172.370 74.185 172.375 ;
        RECT 73.245 172.360 74.175 172.370 ;
        RECT 73.245 172.350 74.170 172.360 ;
        RECT 73.245 172.345 74.165 172.350 ;
        RECT 73.245 172.330 74.155 172.345 ;
        RECT 73.245 172.315 74.150 172.330 ;
        RECT 73.245 172.290 74.140 172.315 ;
        RECT 73.245 172.220 74.135 172.290 ;
        RECT 73.245 171.665 73.795 172.050 ;
        RECT 73.965 171.495 74.135 172.220 ;
        RECT 73.245 171.325 74.135 171.495 ;
        RECT 74.305 171.820 74.635 172.245 ;
        RECT 74.805 172.020 75.035 172.415 ;
        RECT 74.305 171.795 74.555 171.820 ;
        RECT 74.305 171.335 74.525 171.795 ;
        RECT 75.205 171.765 75.375 172.795 ;
        RECT 75.545 172.485 75.865 173.665 ;
        RECT 76.035 172.645 76.235 173.435 ;
        RECT 76.560 172.835 76.945 173.495 ;
        RECT 77.340 172.905 78.125 173.665 ;
        RECT 76.535 172.735 76.945 172.835 ;
        RECT 76.035 172.475 76.365 172.645 ;
        RECT 76.535 172.525 78.145 172.735 ;
        RECT 76.185 172.355 76.365 172.475 ;
        RECT 75.545 172.105 76.010 172.305 ;
        RECT 76.185 172.105 76.515 172.355 ;
        RECT 76.685 172.305 77.150 172.355 ;
        RECT 76.685 172.135 77.155 172.305 ;
        RECT 76.685 172.105 77.150 172.135 ;
        RECT 77.345 172.105 77.700 172.355 ;
        RECT 77.870 171.925 78.145 172.525 ;
        RECT 74.695 171.115 74.945 171.655 ;
        RECT 75.115 171.285 75.375 171.765 ;
        RECT 75.545 171.725 76.725 171.895 ;
        RECT 75.545 171.310 75.885 171.725 ;
        RECT 76.055 171.115 76.225 171.555 ;
        RECT 76.395 171.505 76.725 171.725 ;
        RECT 76.895 171.745 78.145 171.925 ;
        RECT 76.895 171.675 77.260 171.745 ;
        RECT 76.395 171.325 77.645 171.505 ;
        RECT 77.915 171.115 78.085 171.575 ;
        RECT 78.315 171.395 78.595 173.495 ;
        RECT 78.765 173.155 79.955 173.445 ;
        RECT 78.785 172.815 79.955 172.985 ;
        RECT 80.125 172.865 80.405 173.665 ;
        RECT 78.785 172.525 79.110 172.815 ;
        RECT 79.785 172.695 79.955 172.815 ;
        RECT 79.280 172.355 79.475 172.645 ;
        RECT 79.785 172.525 80.445 172.695 ;
        RECT 80.615 172.525 80.890 173.495 ;
        RECT 81.075 172.865 81.405 173.665 ;
        RECT 81.585 173.325 83.015 173.495 ;
        RECT 81.585 172.695 81.835 173.325 ;
        RECT 80.275 172.355 80.445 172.525 ;
        RECT 78.765 172.025 79.110 172.355 ;
        RECT 79.280 172.025 80.105 172.355 ;
        RECT 80.275 172.025 80.550 172.355 ;
        RECT 80.275 171.855 80.445 172.025 ;
        RECT 78.780 171.685 80.445 171.855 ;
        RECT 80.720 171.790 80.890 172.525 ;
        RECT 78.780 171.335 79.035 171.685 ;
        RECT 79.205 171.115 79.535 171.515 ;
        RECT 79.705 171.335 79.875 171.685 ;
        RECT 80.045 171.115 80.425 171.515 ;
        RECT 80.615 171.445 80.890 171.790 ;
        RECT 81.065 172.525 81.835 172.695 ;
        RECT 81.065 171.855 81.235 172.525 ;
        RECT 81.405 172.025 81.810 172.355 ;
        RECT 82.025 172.025 82.275 173.155 ;
        RECT 82.475 172.355 82.675 173.155 ;
        RECT 82.845 172.645 83.015 173.325 ;
        RECT 83.185 172.815 83.500 173.665 ;
        RECT 83.675 172.865 84.115 173.495 ;
        RECT 82.845 172.475 83.635 172.645 ;
        RECT 82.475 172.025 82.720 172.355 ;
        RECT 82.905 172.025 83.295 172.305 ;
        RECT 83.465 172.025 83.635 172.475 ;
        RECT 83.805 171.855 84.115 172.865 ;
        RECT 84.500 172.565 84.830 173.665 ;
        RECT 85.305 173.065 85.630 173.495 ;
        RECT 85.800 173.245 86.130 173.665 ;
        RECT 86.875 173.235 87.285 173.665 ;
        RECT 85.305 172.895 87.285 173.065 ;
        RECT 85.305 172.485 86.010 172.895 ;
        RECT 84.285 172.105 84.930 172.315 ;
        RECT 85.100 172.105 85.670 172.315 ;
        RECT 81.065 171.285 81.555 171.855 ;
        RECT 81.725 171.685 82.885 171.855 ;
        RECT 81.725 171.285 81.955 171.685 ;
        RECT 82.125 171.115 82.545 171.515 ;
        RECT 82.715 171.285 82.885 171.685 ;
        RECT 83.055 171.115 83.505 171.855 ;
        RECT 83.675 171.295 84.115 171.855 ;
        RECT 84.440 171.765 85.610 171.935 ;
        RECT 84.440 171.300 84.770 171.765 ;
        RECT 84.940 171.115 85.110 171.585 ;
        RECT 85.280 171.285 85.610 171.765 ;
        RECT 85.840 171.285 86.010 172.485 ;
        RECT 86.180 172.555 86.805 172.725 ;
        RECT 86.180 171.855 86.350 172.555 ;
        RECT 87.020 172.355 87.285 172.895 ;
        RECT 87.455 172.510 87.795 173.495 ;
        RECT 87.965 173.155 89.155 173.445 ;
        RECT 87.985 172.815 89.155 172.985 ;
        RECT 89.325 172.865 89.605 173.665 ;
        RECT 87.985 172.525 88.310 172.815 ;
        RECT 88.985 172.695 89.155 172.815 ;
        RECT 86.520 172.025 86.850 172.355 ;
        RECT 87.020 172.025 87.370 172.355 ;
        RECT 87.540 171.855 87.795 172.510 ;
        RECT 88.480 172.355 88.675 172.645 ;
        RECT 88.985 172.525 89.645 172.695 ;
        RECT 89.815 172.525 90.090 173.495 ;
        RECT 90.325 172.525 90.535 173.665 ;
        RECT 89.475 172.355 89.645 172.525 ;
        RECT 87.965 172.025 88.310 172.355 ;
        RECT 88.480 172.025 89.305 172.355 ;
        RECT 89.475 172.025 89.750 172.355 ;
        RECT 89.475 171.855 89.645 172.025 ;
        RECT 86.180 171.685 86.720 171.855 ;
        RECT 86.550 171.480 86.720 171.685 ;
        RECT 87.000 171.115 87.170 171.855 ;
        RECT 87.435 171.480 87.795 171.855 ;
        RECT 87.980 171.685 89.645 171.855 ;
        RECT 89.920 171.790 90.090 172.525 ;
        RECT 90.705 172.515 91.035 173.495 ;
        RECT 91.205 172.525 91.435 173.665 ;
        RECT 87.565 171.455 87.735 171.480 ;
        RECT 87.980 171.335 88.235 171.685 ;
        RECT 88.405 171.115 88.735 171.515 ;
        RECT 88.905 171.335 89.075 171.685 ;
        RECT 89.245 171.115 89.625 171.515 ;
        RECT 89.815 171.445 90.090 171.790 ;
        RECT 90.325 171.115 90.535 171.935 ;
        RECT 90.705 171.915 90.955 172.515 ;
        RECT 91.645 172.500 91.935 173.665 ;
        RECT 92.125 172.825 92.455 173.665 ;
        RECT 92.625 172.645 92.970 173.400 ;
        RECT 93.145 173.055 93.490 173.495 ;
        RECT 93.700 173.285 94.030 173.665 ;
        RECT 94.215 173.055 94.450 173.495 ;
        RECT 94.620 173.225 94.950 173.665 ;
        RECT 93.145 172.815 95.155 173.055 ;
        RECT 91.125 172.105 91.455 172.355 ;
        RECT 92.125 172.035 92.455 172.645 ;
        RECT 92.625 172.025 93.255 172.645 ;
        RECT 93.425 172.025 93.715 172.645 ;
        RECT 90.705 171.285 91.035 171.915 ;
        RECT 91.205 171.115 91.435 171.935 ;
        RECT 91.645 171.115 91.935 171.840 ;
        RECT 92.125 171.655 93.490 171.855 ;
        RECT 92.125 171.285 92.455 171.655 ;
        RECT 92.625 171.115 92.955 171.485 ;
        RECT 93.145 171.285 93.490 171.655 ;
        RECT 93.885 171.285 94.215 172.645 ;
        RECT 94.425 172.105 94.755 172.645 ;
        RECT 94.925 171.915 95.155 172.815 ;
        RECT 94.550 171.285 95.155 171.915 ;
        RECT 95.805 172.610 96.110 173.395 ;
        RECT 96.290 173.195 96.975 173.665 ;
        RECT 96.285 172.675 96.980 172.985 ;
        RECT 95.805 171.805 95.980 172.610 ;
        RECT 97.155 172.505 97.440 173.450 ;
        RECT 97.615 173.215 97.945 173.665 ;
        RECT 98.115 173.045 98.285 173.475 ;
        RECT 96.580 172.355 97.440 172.505 ;
        RECT 96.155 172.335 97.440 172.355 ;
        RECT 97.610 172.815 98.285 173.045 ;
        RECT 98.545 173.235 98.885 173.495 ;
        RECT 96.155 171.975 97.140 172.335 ;
        RECT 97.610 172.165 97.845 172.815 ;
        RECT 95.805 171.285 96.045 171.805 ;
        RECT 96.970 171.640 97.140 171.975 ;
        RECT 97.310 171.835 97.845 172.165 ;
        RECT 97.625 171.685 97.845 171.835 ;
        RECT 98.015 171.795 98.315 172.645 ;
        RECT 98.545 171.835 98.805 173.235 ;
        RECT 99.055 172.865 99.385 173.665 ;
        RECT 99.850 172.695 100.100 173.495 ;
        RECT 100.285 172.945 100.615 173.665 ;
        RECT 100.835 172.695 101.085 173.495 ;
        RECT 101.255 173.285 101.590 173.665 ;
        RECT 98.995 172.525 101.185 172.695 ;
        RECT 98.995 172.355 99.310 172.525 ;
        RECT 98.980 172.105 99.310 172.355 ;
        RECT 96.215 171.115 96.610 171.610 ;
        RECT 96.970 171.445 97.345 171.640 ;
        RECT 97.175 171.300 97.345 171.445 ;
        RECT 97.625 171.310 97.865 171.685 ;
        RECT 98.035 171.115 98.370 171.620 ;
        RECT 98.545 171.325 98.885 171.835 ;
        RECT 99.055 171.115 99.325 171.915 ;
        RECT 99.505 171.385 99.785 172.355 ;
        RECT 99.965 171.385 100.265 172.355 ;
        RECT 100.445 171.390 100.795 172.355 ;
        RECT 101.015 171.615 101.185 172.525 ;
        RECT 101.355 171.795 101.595 173.105 ;
        RECT 101.775 172.855 102.070 173.665 ;
        RECT 102.250 172.355 102.495 173.495 ;
        RECT 102.670 172.855 102.930 173.665 ;
        RECT 103.530 173.660 109.805 173.665 ;
        RECT 103.110 172.355 103.360 173.490 ;
        RECT 103.530 172.865 103.790 173.660 ;
        RECT 103.960 172.765 104.220 173.490 ;
        RECT 104.390 172.935 104.650 173.660 ;
        RECT 104.820 172.765 105.080 173.490 ;
        RECT 105.250 172.935 105.510 173.660 ;
        RECT 105.680 172.765 105.940 173.490 ;
        RECT 106.110 172.935 106.370 173.660 ;
        RECT 106.540 172.765 106.800 173.490 ;
        RECT 106.970 172.935 107.215 173.660 ;
        RECT 107.385 172.765 107.645 173.490 ;
        RECT 107.830 172.935 108.075 173.660 ;
        RECT 108.245 172.765 108.505 173.490 ;
        RECT 108.690 172.935 108.935 173.660 ;
        RECT 109.105 172.765 109.365 173.490 ;
        RECT 109.550 172.935 109.805 173.660 ;
        RECT 103.960 172.750 109.365 172.765 ;
        RECT 109.975 172.750 110.265 173.490 ;
        RECT 110.435 172.920 110.705 173.665 ;
        RECT 103.960 172.525 110.705 172.750 ;
        RECT 101.765 171.795 102.080 172.355 ;
        RECT 102.250 172.105 109.370 172.355 ;
        RECT 101.015 171.285 101.510 171.615 ;
        RECT 101.765 171.115 102.070 171.625 ;
        RECT 102.250 171.295 102.500 172.105 ;
        RECT 102.670 171.115 102.930 171.640 ;
        RECT 103.110 171.295 103.360 172.105 ;
        RECT 109.540 171.935 110.705 172.525 ;
        RECT 111.055 172.475 111.225 173.665 ;
        RECT 111.395 172.575 111.725 173.495 ;
        RECT 111.555 172.305 111.725 172.575 ;
        RECT 111.915 172.645 112.245 173.495 ;
        RECT 112.415 172.815 112.585 173.665 ;
        RECT 112.755 172.645 113.085 173.495 ;
        RECT 113.255 172.815 113.425 173.665 ;
        RECT 113.595 172.645 113.925 173.495 ;
        RECT 114.095 172.865 114.265 173.665 ;
        RECT 114.435 172.645 114.765 173.495 ;
        RECT 114.935 172.865 115.105 173.665 ;
        RECT 115.275 172.645 115.605 173.495 ;
        RECT 115.775 172.865 115.945 173.665 ;
        RECT 116.115 172.645 116.445 173.495 ;
        RECT 116.615 172.865 116.785 173.665 ;
        RECT 111.915 172.475 113.425 172.645 ;
        RECT 113.595 172.475 117.235 172.645 ;
        RECT 117.405 172.500 117.695 173.665 ;
        RECT 117.875 172.855 118.170 173.665 ;
        RECT 113.255 172.305 113.425 172.475 ;
        RECT 110.965 172.105 111.385 172.305 ;
        RECT 111.555 172.105 113.085 172.305 ;
        RECT 113.255 172.105 116.640 172.305 ;
        RECT 111.555 171.935 111.725 172.105 ;
        RECT 113.255 171.935 113.425 172.105 ;
        RECT 116.850 171.935 117.235 172.475 ;
        RECT 118.350 172.355 118.595 173.495 ;
        RECT 118.770 172.855 119.030 173.665 ;
        RECT 119.630 173.660 125.905 173.665 ;
        RECT 119.210 172.355 119.460 173.490 ;
        RECT 119.630 172.865 119.890 173.660 ;
        RECT 120.060 172.765 120.320 173.490 ;
        RECT 120.490 172.935 120.750 173.660 ;
        RECT 120.920 172.765 121.180 173.490 ;
        RECT 121.350 172.935 121.610 173.660 ;
        RECT 121.780 172.765 122.040 173.490 ;
        RECT 122.210 172.935 122.470 173.660 ;
        RECT 122.640 172.765 122.900 173.490 ;
        RECT 123.070 172.935 123.315 173.660 ;
        RECT 123.485 172.765 123.745 173.490 ;
        RECT 123.930 172.935 124.175 173.660 ;
        RECT 124.345 172.765 124.605 173.490 ;
        RECT 124.790 172.935 125.035 173.660 ;
        RECT 125.205 172.765 125.465 173.490 ;
        RECT 125.650 172.935 125.905 173.660 ;
        RECT 120.060 172.750 125.465 172.765 ;
        RECT 126.075 172.750 126.365 173.490 ;
        RECT 126.535 172.920 126.805 173.665 ;
        RECT 127.075 172.855 127.370 173.665 ;
        RECT 120.060 172.525 126.805 172.750 ;
        RECT 103.960 171.765 110.705 171.935 ;
        RECT 103.530 171.115 103.790 171.675 ;
        RECT 103.960 171.310 104.220 171.765 ;
        RECT 104.390 171.115 104.650 171.595 ;
        RECT 104.820 171.310 105.080 171.765 ;
        RECT 105.250 171.115 105.510 171.595 ;
        RECT 105.680 171.310 105.940 171.765 ;
        RECT 106.110 171.115 106.355 171.595 ;
        RECT 106.525 171.310 106.800 171.765 ;
        RECT 106.970 171.115 107.215 171.595 ;
        RECT 107.385 171.310 107.645 171.765 ;
        RECT 107.825 171.115 108.075 171.595 ;
        RECT 108.245 171.310 108.505 171.765 ;
        RECT 108.685 171.115 108.935 171.595 ;
        RECT 109.105 171.310 109.365 171.765 ;
        RECT 109.545 171.115 109.805 171.595 ;
        RECT 109.975 171.310 110.235 171.765 ;
        RECT 110.405 171.115 110.705 171.595 ;
        RECT 111.055 171.115 111.225 171.935 ;
        RECT 111.395 171.290 111.725 171.935 ;
        RECT 111.915 171.765 113.425 171.935 ;
        RECT 113.595 171.765 117.235 171.935 ;
        RECT 111.915 171.290 112.245 171.765 ;
        RECT 112.415 171.115 112.585 171.595 ;
        RECT 112.755 171.290 113.085 171.765 ;
        RECT 113.255 171.115 113.425 171.595 ;
        RECT 113.595 171.290 113.925 171.765 ;
        RECT 114.095 171.115 114.265 171.595 ;
        RECT 114.435 171.290 114.765 171.765 ;
        RECT 114.935 171.115 115.105 171.595 ;
        RECT 115.275 171.290 115.605 171.765 ;
        RECT 115.775 171.115 115.945 171.595 ;
        RECT 116.115 171.290 116.445 171.765 ;
        RECT 116.615 171.115 116.785 171.595 ;
        RECT 117.405 171.115 117.695 171.840 ;
        RECT 117.865 171.795 118.180 172.355 ;
        RECT 118.350 172.105 125.470 172.355 ;
        RECT 117.865 171.115 118.170 171.625 ;
        RECT 118.350 171.295 118.600 172.105 ;
        RECT 118.770 171.115 119.030 171.640 ;
        RECT 119.210 171.295 119.460 172.105 ;
        RECT 125.640 171.935 126.805 172.525 ;
        RECT 127.550 172.355 127.795 173.495 ;
        RECT 127.970 172.855 128.230 173.665 ;
        RECT 128.830 173.660 135.105 173.665 ;
        RECT 128.410 172.355 128.660 173.490 ;
        RECT 128.830 172.865 129.090 173.660 ;
        RECT 129.260 172.765 129.520 173.490 ;
        RECT 129.690 172.935 129.950 173.660 ;
        RECT 130.120 172.765 130.380 173.490 ;
        RECT 130.550 172.935 130.810 173.660 ;
        RECT 130.980 172.765 131.240 173.490 ;
        RECT 131.410 172.935 131.670 173.660 ;
        RECT 131.840 172.765 132.100 173.490 ;
        RECT 132.270 172.935 132.515 173.660 ;
        RECT 132.685 172.765 132.945 173.490 ;
        RECT 133.130 172.935 133.375 173.660 ;
        RECT 133.545 172.765 133.805 173.490 ;
        RECT 133.990 172.935 134.235 173.660 ;
        RECT 134.405 172.765 134.665 173.490 ;
        RECT 134.850 172.935 135.105 173.660 ;
        RECT 129.260 172.750 134.665 172.765 ;
        RECT 135.275 172.750 135.565 173.490 ;
        RECT 135.735 172.920 136.005 173.665 ;
        RECT 129.260 172.525 136.005 172.750 ;
        RECT 136.450 172.695 136.840 172.870 ;
        RECT 137.325 172.865 137.655 173.665 ;
        RECT 137.825 172.875 138.360 173.495 ;
        RECT 136.450 172.525 137.875 172.695 ;
        RECT 120.060 171.765 126.805 171.935 ;
        RECT 127.065 171.795 127.380 172.355 ;
        RECT 127.550 172.105 134.670 172.355 ;
        RECT 119.630 171.115 119.890 171.675 ;
        RECT 120.060 171.310 120.320 171.765 ;
        RECT 120.490 171.115 120.750 171.595 ;
        RECT 120.920 171.310 121.180 171.765 ;
        RECT 121.350 171.115 121.610 171.595 ;
        RECT 121.780 171.310 122.040 171.765 ;
        RECT 122.210 171.115 122.455 171.595 ;
        RECT 122.625 171.310 122.900 171.765 ;
        RECT 123.070 171.115 123.315 171.595 ;
        RECT 123.485 171.310 123.745 171.765 ;
        RECT 123.925 171.115 124.175 171.595 ;
        RECT 124.345 171.310 124.605 171.765 ;
        RECT 124.785 171.115 125.035 171.595 ;
        RECT 125.205 171.310 125.465 171.765 ;
        RECT 125.645 171.115 125.905 171.595 ;
        RECT 126.075 171.310 126.335 171.765 ;
        RECT 126.505 171.115 126.805 171.595 ;
        RECT 127.065 171.115 127.370 171.625 ;
        RECT 127.550 171.295 127.800 172.105 ;
        RECT 127.970 171.115 128.230 171.640 ;
        RECT 128.410 171.295 128.660 172.105 ;
        RECT 134.840 171.935 136.005 172.525 ;
        RECT 129.260 171.765 136.005 171.935 ;
        RECT 136.325 171.795 136.680 172.355 ;
        RECT 128.830 171.115 129.090 171.675 ;
        RECT 129.260 171.310 129.520 171.765 ;
        RECT 129.690 171.115 129.950 171.595 ;
        RECT 130.120 171.310 130.380 171.765 ;
        RECT 130.550 171.115 130.810 171.595 ;
        RECT 130.980 171.310 131.240 171.765 ;
        RECT 131.410 171.115 131.655 171.595 ;
        RECT 131.825 171.310 132.100 171.765 ;
        RECT 132.270 171.115 132.515 171.595 ;
        RECT 132.685 171.310 132.945 171.765 ;
        RECT 133.125 171.115 133.375 171.595 ;
        RECT 133.545 171.310 133.805 171.765 ;
        RECT 133.985 171.115 134.235 171.595 ;
        RECT 134.405 171.310 134.665 171.765 ;
        RECT 134.845 171.115 135.105 171.595 ;
        RECT 135.275 171.310 135.535 171.765 ;
        RECT 136.850 171.625 137.020 172.525 ;
        RECT 137.190 171.795 137.455 172.355 ;
        RECT 137.705 172.025 137.875 172.525 ;
        RECT 138.045 171.855 138.360 172.875 ;
        RECT 138.565 172.575 139.775 173.665 ;
        RECT 138.565 172.035 139.085 172.575 ;
        RECT 139.255 171.865 139.775 172.405 ;
        RECT 135.705 171.115 136.005 171.595 ;
        RECT 136.430 171.115 136.670 171.625 ;
        RECT 136.850 171.295 137.130 171.625 ;
        RECT 137.360 171.115 137.575 171.625 ;
        RECT 137.745 171.285 138.360 171.855 ;
        RECT 138.565 171.115 139.775 171.865 ;
        RECT 27.160 170.945 139.860 171.115 ;
        RECT 27.245 170.195 28.455 170.945 ;
        RECT 28.805 170.285 29.145 170.945 ;
        RECT 27.245 169.655 27.765 170.195 ;
        RECT 27.935 169.485 28.455 170.025 ;
        RECT 27.245 168.395 28.455 169.485 ;
        RECT 28.625 168.565 29.145 170.115 ;
        RECT 29.315 169.290 29.835 170.775 ;
        RECT 30.005 170.400 35.350 170.945 ;
        RECT 35.525 170.400 40.870 170.945 ;
        RECT 41.045 170.400 46.390 170.945 ;
        RECT 46.565 170.400 51.910 170.945 ;
        RECT 31.590 169.570 31.930 170.400 ;
        RECT 29.315 168.395 29.645 169.120 ;
        RECT 33.410 168.830 33.760 170.080 ;
        RECT 37.110 169.570 37.450 170.400 ;
        RECT 38.930 168.830 39.280 170.080 ;
        RECT 42.630 169.570 42.970 170.400 ;
        RECT 44.450 168.830 44.800 170.080 ;
        RECT 48.150 169.570 48.490 170.400 ;
        RECT 53.005 170.220 53.295 170.945 ;
        RECT 53.465 170.195 54.675 170.945 ;
        RECT 49.970 168.830 50.320 170.080 ;
        RECT 53.465 169.655 53.985 170.195 ;
        RECT 54.850 170.105 55.110 170.945 ;
        RECT 55.285 170.200 55.540 170.775 ;
        RECT 55.710 170.565 56.040 170.945 ;
        RECT 56.255 170.395 56.425 170.775 ;
        RECT 55.710 170.225 56.425 170.395 ;
        RECT 56.690 170.375 57.010 170.775 ;
        RECT 30.005 168.395 35.350 168.830 ;
        RECT 35.525 168.395 40.870 168.830 ;
        RECT 41.045 168.395 46.390 168.830 ;
        RECT 46.565 168.395 51.910 168.830 ;
        RECT 53.005 168.395 53.295 169.560 ;
        RECT 54.155 169.485 54.675 170.025 ;
        RECT 53.465 168.395 54.675 169.485 ;
        RECT 54.850 168.395 55.110 169.545 ;
        RECT 55.285 169.470 55.455 170.200 ;
        RECT 55.710 170.035 55.880 170.225 ;
        RECT 55.625 169.705 55.880 170.035 ;
        RECT 55.710 169.495 55.880 169.705 ;
        RECT 56.160 169.675 56.515 170.045 ;
        RECT 56.690 169.585 56.860 170.375 ;
        RECT 57.180 170.125 57.490 170.945 ;
        RECT 57.660 170.315 57.990 170.775 ;
        RECT 58.160 170.485 58.410 170.945 ;
        RECT 58.600 170.565 60.650 170.775 ;
        RECT 58.600 170.315 59.350 170.395 ;
        RECT 57.660 170.125 59.350 170.315 ;
        RECT 59.520 170.125 59.690 170.565 ;
        RECT 61.375 170.395 61.545 170.775 ;
        RECT 61.760 170.565 62.090 170.945 ;
        RECT 59.860 170.125 60.650 170.395 ;
        RECT 61.375 170.225 62.090 170.395 ;
        RECT 57.030 169.755 57.380 169.955 ;
        RECT 57.660 169.755 58.340 169.955 ;
        RECT 58.550 169.755 59.740 169.955 ;
        RECT 59.920 169.585 60.250 169.955 ;
        RECT 55.285 168.565 55.540 169.470 ;
        RECT 55.710 169.325 56.425 169.495 ;
        RECT 55.710 168.395 56.040 169.155 ;
        RECT 56.255 168.565 56.425 169.325 ;
        RECT 56.690 169.415 60.250 169.585 ;
        RECT 56.690 168.965 56.860 169.415 ;
        RECT 60.450 169.245 60.650 170.125 ;
        RECT 61.285 169.675 61.640 170.045 ;
        RECT 61.920 170.035 62.090 170.225 ;
        RECT 62.260 170.200 62.515 170.775 ;
        RECT 61.920 169.705 62.175 170.035 ;
        RECT 61.920 169.495 62.090 169.705 ;
        RECT 56.690 168.565 57.010 168.965 ;
        RECT 57.180 168.395 57.490 169.195 ;
        RECT 57.660 169.075 60.650 169.245 ;
        RECT 57.660 169.025 58.830 169.075 ;
        RECT 57.660 168.565 57.990 169.025 ;
        RECT 58.160 168.395 58.330 168.855 ;
        RECT 58.500 168.565 58.830 169.025 ;
        RECT 59.860 169.025 60.650 169.075 ;
        RECT 61.375 169.325 62.090 169.495 ;
        RECT 62.345 169.470 62.515 170.200 ;
        RECT 62.690 170.105 62.950 170.945 ;
        RECT 63.220 170.005 63.390 170.945 ;
        RECT 63.560 170.270 63.835 170.615 ;
        RECT 64.025 170.545 64.405 170.945 ;
        RECT 64.575 170.375 64.745 170.725 ;
        RECT 64.915 170.545 65.245 170.945 ;
        RECT 65.445 170.375 65.615 170.725 ;
        RECT 65.790 170.545 66.145 170.945 ;
        RECT 66.390 170.375 66.560 170.580 ;
        RECT 59.000 168.395 59.250 168.855 ;
        RECT 59.440 168.395 59.690 168.855 ;
        RECT 59.860 168.565 60.110 169.025 ;
        RECT 60.360 168.395 60.650 168.855 ;
        RECT 61.375 168.565 61.545 169.325 ;
        RECT 61.760 168.395 62.090 169.155 ;
        RECT 62.260 168.565 62.515 169.470 ;
        RECT 62.690 168.395 62.950 169.545 ;
        RECT 63.220 168.395 63.390 169.590 ;
        RECT 63.560 169.535 63.730 170.270 ;
        RECT 64.005 170.205 65.615 170.375 ;
        RECT 66.040 170.205 66.560 170.375 ;
        RECT 66.810 170.205 66.980 170.945 ;
        RECT 67.235 170.205 67.555 170.580 ;
        RECT 67.730 170.565 69.780 170.775 ;
        RECT 64.005 170.035 64.175 170.205 ;
        RECT 63.900 169.705 64.175 170.035 ;
        RECT 64.345 169.705 65.000 170.035 ;
        RECT 64.005 169.535 64.175 169.705 ;
        RECT 65.220 169.615 65.390 170.035 ;
        RECT 66.040 169.955 66.230 170.205 ;
        RECT 65.785 169.785 66.230 169.955 ;
        RECT 63.560 168.565 63.835 169.535 ;
        RECT 64.005 169.365 64.665 169.535 ;
        RECT 65.220 169.445 65.870 169.615 ;
        RECT 64.495 169.245 64.665 169.365 ;
        RECT 64.045 168.395 64.325 169.195 ;
        RECT 64.495 169.075 65.530 169.245 ;
        RECT 64.495 168.575 65.135 168.905 ;
        RECT 65.360 168.825 65.530 169.075 ;
        RECT 65.700 169.165 65.870 169.445 ;
        RECT 66.040 169.505 66.230 169.785 ;
        RECT 66.400 169.705 66.690 170.035 ;
        RECT 66.040 169.335 66.645 169.505 ;
        RECT 66.860 169.335 67.210 170.035 ;
        RECT 67.380 169.165 67.555 170.205 ;
        RECT 65.700 168.995 67.555 169.165 ;
        RECT 67.730 170.125 68.520 170.395 ;
        RECT 68.690 170.125 68.860 170.565 ;
        RECT 69.970 170.485 70.220 170.945 ;
        RECT 69.030 170.315 69.780 170.395 ;
        RECT 70.390 170.315 70.720 170.775 ;
        RECT 69.030 170.125 70.720 170.315 ;
        RECT 70.890 170.125 71.200 170.945 ;
        RECT 71.370 170.375 71.690 170.775 ;
        RECT 67.730 169.245 67.930 170.125 ;
        RECT 68.130 169.585 68.460 169.955 ;
        RECT 68.640 169.755 69.830 169.955 ;
        RECT 70.040 169.755 70.720 169.955 ;
        RECT 71.000 169.755 71.350 169.955 ;
        RECT 71.520 169.585 71.690 170.375 ;
        RECT 72.875 170.395 73.045 170.775 ;
        RECT 73.225 170.565 73.555 170.945 ;
        RECT 72.875 170.225 73.540 170.395 ;
        RECT 73.735 170.270 73.995 170.775 ;
        RECT 74.165 170.565 75.055 170.735 ;
        RECT 72.805 169.675 73.135 170.045 ;
        RECT 73.370 169.970 73.540 170.225 ;
        RECT 68.130 169.415 71.690 169.585 ;
        RECT 73.370 169.640 73.655 169.970 ;
        RECT 73.370 169.495 73.540 169.640 ;
        RECT 67.730 169.075 70.720 169.245 ;
        RECT 67.730 169.025 68.520 169.075 ;
        RECT 65.360 168.655 66.105 168.825 ;
        RECT 66.795 168.395 67.125 168.825 ;
        RECT 67.295 168.575 67.555 168.995 ;
        RECT 67.730 168.395 68.020 168.855 ;
        RECT 68.270 168.565 68.520 169.025 ;
        RECT 69.550 169.025 70.720 169.075 ;
        RECT 68.690 168.395 68.940 168.855 ;
        RECT 69.130 168.395 69.380 168.855 ;
        RECT 69.550 168.565 69.880 169.025 ;
        RECT 70.050 168.395 70.220 168.855 ;
        RECT 70.390 168.565 70.720 169.025 ;
        RECT 70.890 168.395 71.200 169.195 ;
        RECT 71.520 168.965 71.690 169.415 ;
        RECT 71.370 168.565 71.690 168.965 ;
        RECT 72.875 169.325 73.540 169.495 ;
        RECT 73.825 169.470 73.995 170.270 ;
        RECT 74.165 170.010 74.715 170.395 ;
        RECT 74.885 169.840 75.055 170.565 ;
        RECT 72.875 168.565 73.045 169.325 ;
        RECT 73.225 168.395 73.555 169.155 ;
        RECT 73.725 168.565 73.995 169.470 ;
        RECT 74.165 169.770 75.055 169.840 ;
        RECT 75.225 170.240 75.445 170.725 ;
        RECT 75.615 170.405 75.865 170.945 ;
        RECT 76.035 170.295 76.295 170.775 ;
        RECT 76.465 170.565 77.355 170.735 ;
        RECT 75.225 169.815 75.555 170.240 ;
        RECT 74.165 169.745 75.060 169.770 ;
        RECT 74.165 169.730 75.070 169.745 ;
        RECT 74.165 169.715 75.075 169.730 ;
        RECT 74.165 169.710 75.085 169.715 ;
        RECT 74.165 169.700 75.090 169.710 ;
        RECT 74.165 169.690 75.095 169.700 ;
        RECT 74.165 169.685 75.105 169.690 ;
        RECT 74.165 169.675 75.115 169.685 ;
        RECT 74.165 169.670 75.125 169.675 ;
        RECT 74.165 169.220 74.425 169.670 ;
        RECT 74.790 169.665 75.125 169.670 ;
        RECT 74.790 169.660 75.140 169.665 ;
        RECT 74.790 169.650 75.155 169.660 ;
        RECT 74.790 169.645 75.180 169.650 ;
        RECT 75.725 169.645 75.955 170.040 ;
        RECT 74.790 169.640 75.955 169.645 ;
        RECT 74.820 169.605 75.955 169.640 ;
        RECT 74.855 169.580 75.955 169.605 ;
        RECT 74.885 169.550 75.955 169.580 ;
        RECT 74.905 169.520 75.955 169.550 ;
        RECT 74.925 169.490 75.955 169.520 ;
        RECT 74.995 169.480 75.955 169.490 ;
        RECT 75.020 169.470 75.955 169.480 ;
        RECT 75.040 169.455 75.955 169.470 ;
        RECT 75.060 169.440 75.955 169.455 ;
        RECT 75.065 169.430 75.850 169.440 ;
        RECT 75.080 169.395 75.850 169.430 ;
        RECT 74.595 169.075 74.925 169.320 ;
        RECT 75.095 169.145 75.850 169.395 ;
        RECT 76.125 169.265 76.295 170.295 ;
        RECT 76.465 170.010 77.015 170.395 ;
        RECT 77.185 169.840 77.355 170.565 ;
        RECT 74.595 169.050 74.780 169.075 ;
        RECT 74.165 168.950 74.780 169.050 ;
        RECT 74.165 168.395 74.770 168.950 ;
        RECT 74.945 168.565 75.425 168.905 ;
        RECT 75.595 168.395 75.850 168.940 ;
        RECT 76.020 168.565 76.295 169.265 ;
        RECT 76.465 169.770 77.355 169.840 ;
        RECT 77.525 170.240 77.745 170.725 ;
        RECT 77.915 170.405 78.165 170.945 ;
        RECT 78.335 170.295 78.595 170.775 ;
        RECT 77.525 169.815 77.855 170.240 ;
        RECT 76.465 169.745 77.360 169.770 ;
        RECT 76.465 169.730 77.370 169.745 ;
        RECT 76.465 169.715 77.375 169.730 ;
        RECT 76.465 169.710 77.385 169.715 ;
        RECT 76.465 169.700 77.390 169.710 ;
        RECT 76.465 169.690 77.395 169.700 ;
        RECT 76.465 169.685 77.405 169.690 ;
        RECT 76.465 169.675 77.415 169.685 ;
        RECT 76.465 169.670 77.425 169.675 ;
        RECT 76.465 169.220 76.725 169.670 ;
        RECT 77.090 169.665 77.425 169.670 ;
        RECT 77.090 169.660 77.440 169.665 ;
        RECT 77.090 169.650 77.455 169.660 ;
        RECT 77.090 169.645 77.480 169.650 ;
        RECT 78.025 169.645 78.255 170.040 ;
        RECT 77.090 169.640 78.255 169.645 ;
        RECT 77.120 169.605 78.255 169.640 ;
        RECT 77.155 169.580 78.255 169.605 ;
        RECT 77.185 169.550 78.255 169.580 ;
        RECT 77.205 169.520 78.255 169.550 ;
        RECT 77.225 169.490 78.255 169.520 ;
        RECT 77.295 169.480 78.255 169.490 ;
        RECT 77.320 169.470 78.255 169.480 ;
        RECT 77.340 169.455 78.255 169.470 ;
        RECT 77.360 169.440 78.255 169.455 ;
        RECT 77.365 169.430 78.150 169.440 ;
        RECT 77.380 169.395 78.150 169.430 ;
        RECT 76.895 169.075 77.225 169.320 ;
        RECT 77.395 169.145 78.150 169.395 ;
        RECT 78.425 169.265 78.595 170.295 ;
        RECT 78.765 170.220 79.055 170.945 ;
        RECT 79.380 170.295 79.710 170.760 ;
        RECT 79.880 170.475 80.050 170.945 ;
        RECT 80.220 170.295 80.550 170.775 ;
        RECT 79.380 170.125 80.550 170.295 ;
        RECT 79.225 169.745 79.870 169.955 ;
        RECT 80.040 169.745 80.610 169.955 ;
        RECT 80.780 169.575 80.950 170.775 ;
        RECT 81.490 170.375 81.660 170.580 ;
        RECT 76.895 169.050 77.080 169.075 ;
        RECT 76.465 168.950 77.080 169.050 ;
        RECT 76.465 168.395 77.070 168.950 ;
        RECT 77.245 168.565 77.725 168.905 ;
        RECT 77.895 168.395 78.150 168.940 ;
        RECT 78.320 168.565 78.595 169.265 ;
        RECT 78.765 168.395 79.055 169.560 ;
        RECT 79.440 168.395 79.770 169.495 ;
        RECT 80.245 169.165 80.950 169.575 ;
        RECT 81.120 170.205 81.660 170.375 ;
        RECT 81.940 170.205 82.110 170.945 ;
        RECT 82.505 170.580 82.675 170.605 ;
        RECT 82.375 170.205 82.735 170.580 ;
        RECT 81.120 169.505 81.290 170.205 ;
        RECT 81.460 169.705 81.790 170.035 ;
        RECT 81.960 169.705 82.310 170.035 ;
        RECT 81.120 169.335 81.745 169.505 ;
        RECT 81.960 169.165 82.225 169.705 ;
        RECT 82.480 169.550 82.735 170.205 ;
        RECT 80.245 168.995 82.225 169.165 ;
        RECT 80.245 168.565 80.570 168.995 ;
        RECT 80.740 168.395 81.070 168.815 ;
        RECT 81.815 168.395 82.225 168.825 ;
        RECT 82.395 168.565 82.735 169.550 ;
        RECT 82.905 170.445 83.165 170.775 ;
        RECT 83.375 170.465 83.650 170.945 ;
        RECT 82.905 169.535 83.075 170.445 ;
        RECT 83.860 170.375 84.065 170.775 ;
        RECT 84.235 170.545 84.570 170.945 ;
        RECT 84.745 170.445 85.005 170.775 ;
        RECT 85.215 170.465 85.490 170.945 ;
        RECT 83.245 169.705 83.605 170.285 ;
        RECT 83.860 170.205 84.545 170.375 ;
        RECT 83.785 169.535 84.035 170.035 ;
        RECT 82.905 169.365 84.035 169.535 ;
        RECT 82.905 168.595 83.175 169.365 ;
        RECT 84.205 169.175 84.545 170.205 ;
        RECT 83.345 168.395 83.675 169.175 ;
        RECT 83.880 169.000 84.545 169.175 ;
        RECT 84.745 169.535 84.915 170.445 ;
        RECT 85.700 170.375 85.905 170.775 ;
        RECT 86.075 170.545 86.410 170.945 ;
        RECT 86.585 170.485 87.145 170.775 ;
        RECT 87.315 170.485 87.565 170.945 ;
        RECT 85.085 169.705 85.445 170.285 ;
        RECT 85.700 170.205 86.385 170.375 ;
        RECT 85.625 169.535 85.875 170.035 ;
        RECT 84.745 169.365 85.875 169.535 ;
        RECT 83.880 168.595 84.065 169.000 ;
        RECT 84.235 168.395 84.570 168.820 ;
        RECT 84.745 168.595 85.015 169.365 ;
        RECT 86.045 169.175 86.385 170.205 ;
        RECT 85.185 168.395 85.515 169.175 ;
        RECT 85.720 169.000 86.385 169.175 ;
        RECT 86.585 169.115 86.835 170.485 ;
        RECT 88.185 170.315 88.515 170.675 ;
        RECT 87.125 170.125 88.515 170.315 ;
        RECT 88.975 170.395 89.145 170.775 ;
        RECT 89.315 170.565 89.645 170.945 ;
        RECT 88.975 170.225 89.470 170.395 ;
        RECT 87.125 170.035 87.295 170.125 ;
        RECT 87.005 169.705 87.295 170.035 ;
        RECT 87.465 169.705 87.805 169.955 ;
        RECT 88.025 169.705 88.700 169.955 ;
        RECT 87.125 169.455 87.295 169.705 ;
        RECT 87.125 169.285 88.065 169.455 ;
        RECT 88.435 169.345 88.700 169.705 ;
        RECT 88.950 169.585 89.130 170.035 ;
        RECT 88.945 169.415 89.130 169.585 ;
        RECT 88.950 169.395 89.130 169.415 ;
        RECT 85.720 168.595 85.905 169.000 ;
        RECT 86.075 168.395 86.410 168.820 ;
        RECT 86.585 168.565 87.045 169.115 ;
        RECT 87.235 168.395 87.565 169.115 ;
        RECT 87.765 168.735 88.065 169.285 ;
        RECT 89.300 169.145 89.470 170.225 ;
        RECT 89.815 169.485 90.040 170.775 ;
        RECT 90.210 170.565 90.540 170.945 ;
        RECT 90.810 170.395 90.980 170.775 ;
        RECT 91.710 170.605 91.975 170.610 ;
        RECT 91.705 170.435 91.975 170.605 ;
        RECT 90.215 170.225 91.205 170.395 ;
        RECT 90.215 169.705 90.385 170.225 ;
        RECT 90.555 169.705 90.865 170.035 ;
        RECT 89.790 169.315 90.120 169.485 ;
        RECT 90.555 169.145 90.725 169.705 ;
        RECT 88.235 168.395 88.515 169.065 ;
        RECT 88.975 168.975 90.725 169.145 ;
        RECT 91.035 169.115 91.205 170.225 ;
        RECT 91.710 169.755 91.975 170.435 ;
        RECT 91.375 169.455 91.545 169.630 ;
        RECT 92.150 169.625 92.455 170.605 ;
        RECT 92.635 170.445 92.885 170.945 ;
        RECT 93.055 170.445 93.315 170.775 ;
        RECT 92.625 169.725 92.975 170.265 ;
        RECT 91.375 169.285 92.555 169.455 ;
        RECT 92.385 169.115 92.555 169.285 ;
        RECT 93.145 169.115 93.315 170.445 ;
        RECT 93.505 170.405 93.835 170.775 ;
        RECT 94.005 170.575 94.335 170.945 ;
        RECT 94.525 170.405 94.870 170.775 ;
        RECT 93.505 170.205 94.870 170.405 ;
        RECT 93.505 169.415 93.835 170.025 ;
        RECT 94.005 169.415 94.635 170.035 ;
        RECT 94.805 169.415 95.095 170.035 ;
        RECT 95.265 169.415 95.595 170.775 ;
        RECT 95.930 170.145 96.535 170.775 ;
        RECT 95.805 169.415 96.135 169.955 ;
        RECT 88.975 168.565 89.145 168.975 ;
        RECT 91.035 168.945 92.215 169.115 ;
        RECT 92.385 168.945 93.315 169.115 ;
        RECT 89.315 168.395 89.645 168.775 ;
        RECT 90.290 168.395 90.960 168.775 ;
        RECT 91.195 168.565 91.365 168.945 ;
        RECT 91.535 168.395 91.875 168.775 ;
        RECT 92.045 168.565 92.215 168.945 ;
        RECT 92.555 168.395 92.885 168.775 ;
        RECT 93.055 168.565 93.315 168.945 ;
        RECT 93.505 168.395 93.835 169.235 ;
        RECT 94.005 168.660 94.350 169.415 ;
        RECT 96.305 169.245 96.535 170.145 ;
        RECT 96.905 170.315 97.235 170.675 ;
        RECT 97.865 170.485 98.115 170.945 ;
        RECT 98.285 170.485 98.835 170.775 ;
        RECT 96.905 170.125 98.295 170.315 ;
        RECT 98.125 170.035 98.295 170.125 ;
        RECT 96.705 169.705 97.395 169.955 ;
        RECT 97.625 169.705 97.955 169.955 ;
        RECT 98.125 169.705 98.415 170.035 ;
        RECT 96.705 169.265 97.020 169.705 ;
        RECT 98.125 169.455 98.295 169.705 ;
        RECT 97.355 169.285 98.295 169.455 ;
        RECT 94.525 169.005 96.535 169.245 ;
        RECT 94.525 168.565 94.870 169.005 ;
        RECT 95.080 168.395 95.410 168.775 ;
        RECT 95.595 168.565 95.830 169.005 ;
        RECT 96.000 168.395 96.330 168.835 ;
        RECT 96.905 168.395 97.185 169.065 ;
        RECT 97.355 168.735 97.655 169.285 ;
        RECT 98.585 169.115 98.835 170.485 ;
        RECT 99.005 170.145 99.295 170.945 ;
        RECT 99.515 170.475 99.805 170.945 ;
        RECT 99.975 170.305 100.305 170.775 ;
        RECT 100.475 170.475 101.185 170.945 ;
        RECT 101.355 170.305 101.685 170.775 ;
        RECT 101.855 170.475 102.025 170.945 ;
        RECT 102.195 170.305 102.525 170.775 ;
        RECT 99.465 170.125 102.525 170.305 ;
        RECT 102.695 170.125 102.970 170.945 ;
        RECT 103.235 170.395 103.405 170.775 ;
        RECT 103.585 170.565 103.915 170.945 ;
        RECT 103.235 170.225 103.900 170.395 ;
        RECT 104.095 170.270 104.355 170.775 ;
        RECT 99.465 169.575 99.925 170.125 ;
        RECT 100.095 169.745 100.685 169.955 ;
        RECT 100.875 169.745 101.925 169.955 ;
        RECT 102.095 169.745 102.925 169.955 ;
        RECT 97.865 168.395 98.195 169.115 ;
        RECT 98.385 168.565 98.835 169.115 ;
        RECT 99.005 168.395 99.295 169.535 ;
        RECT 99.465 169.405 100.225 169.575 ;
        RECT 100.420 169.405 100.685 169.745 ;
        RECT 103.165 169.675 103.495 170.045 ;
        RECT 103.730 169.970 103.900 170.225 ;
        RECT 103.730 169.640 104.015 169.970 ;
        RECT 100.975 169.405 102.910 169.575 ;
        RECT 103.730 169.495 103.900 169.640 ;
        RECT 99.595 168.735 99.845 169.235 ;
        RECT 100.015 168.905 100.225 169.405 ;
        RECT 100.435 168.735 100.645 169.235 ;
        RECT 100.975 168.905 101.225 169.405 ;
        RECT 101.395 168.735 101.645 169.235 ;
        RECT 99.595 168.565 101.645 168.735 ;
        RECT 101.815 168.565 102.065 169.405 ;
        RECT 102.235 168.395 102.485 169.235 ;
        RECT 102.655 168.565 102.910 169.405 ;
        RECT 103.235 169.325 103.900 169.495 ;
        RECT 104.185 169.470 104.355 170.270 ;
        RECT 104.525 170.220 104.815 170.945 ;
        RECT 104.985 170.335 105.335 170.775 ;
        RECT 105.505 170.505 105.675 170.945 ;
        RECT 105.845 170.565 107.040 170.775 ;
        RECT 105.845 170.335 106.095 170.565 ;
        RECT 104.985 170.125 106.095 170.335 ;
        RECT 106.265 170.125 106.595 170.395 ;
        RECT 106.765 170.125 107.040 170.565 ;
        RECT 107.275 170.205 107.605 170.945 ;
        RECT 107.775 170.190 108.010 170.520 ;
        RECT 106.310 170.095 106.595 170.125 ;
        RECT 104.985 169.755 106.130 169.955 ;
        RECT 105.940 169.585 106.130 169.755 ;
        RECT 103.235 168.565 103.405 169.325 ;
        RECT 103.585 168.395 103.915 169.155 ;
        RECT 104.085 168.565 104.355 169.470 ;
        RECT 104.525 168.395 104.815 169.560 ;
        RECT 104.985 168.395 105.315 169.535 ;
        RECT 105.485 169.195 105.760 169.535 ;
        RECT 105.940 169.415 106.135 169.585 ;
        RECT 105.940 169.375 106.130 169.415 ;
        RECT 106.310 169.195 106.590 170.095 ;
        RECT 106.760 169.535 107.090 169.955 ;
        RECT 107.320 169.705 107.665 170.035 ;
        RECT 107.840 169.535 108.010 170.190 ;
        RECT 106.760 169.365 108.010 169.535 ;
        RECT 105.485 169.025 107.085 169.195 ;
        RECT 105.485 168.565 105.840 169.025 ;
        RECT 106.010 168.395 106.585 168.855 ;
        RECT 106.755 168.565 107.085 169.025 ;
        RECT 107.285 168.395 107.540 169.195 ;
        RECT 107.710 169.170 108.010 169.365 ;
        RECT 108.205 170.445 108.505 170.775 ;
        RECT 108.675 170.465 108.950 170.945 ;
        RECT 108.205 169.535 108.375 170.445 ;
        RECT 109.130 170.295 109.425 170.685 ;
        RECT 109.595 170.465 109.850 170.945 ;
        RECT 110.025 170.295 110.285 170.685 ;
        RECT 110.455 170.465 110.735 170.945 ;
        RECT 110.965 170.435 111.270 170.945 ;
        RECT 108.545 169.705 108.895 170.275 ;
        RECT 109.130 170.125 110.780 170.295 ;
        RECT 109.065 169.785 110.205 169.955 ;
        RECT 109.065 169.535 109.235 169.785 ;
        RECT 110.375 169.615 110.780 170.125 ;
        RECT 110.965 169.705 111.280 170.265 ;
        RECT 111.450 169.955 111.700 170.765 ;
        RECT 111.870 170.420 112.130 170.945 ;
        RECT 112.310 169.955 112.560 170.765 ;
        RECT 112.730 170.385 112.990 170.945 ;
        RECT 113.160 170.295 113.420 170.750 ;
        RECT 113.590 170.465 113.850 170.945 ;
        RECT 114.020 170.295 114.280 170.750 ;
        RECT 114.450 170.465 114.710 170.945 ;
        RECT 114.880 170.295 115.140 170.750 ;
        RECT 115.310 170.465 115.555 170.945 ;
        RECT 115.725 170.295 116.000 170.750 ;
        RECT 116.170 170.465 116.415 170.945 ;
        RECT 116.585 170.295 116.845 170.750 ;
        RECT 117.025 170.465 117.275 170.945 ;
        RECT 117.445 170.295 117.705 170.750 ;
        RECT 117.885 170.465 118.135 170.945 ;
        RECT 118.305 170.295 118.565 170.750 ;
        RECT 118.745 170.465 119.005 170.945 ;
        RECT 119.175 170.295 119.435 170.750 ;
        RECT 119.605 170.465 119.905 170.945 ;
        RECT 120.255 170.465 120.555 170.945 ;
        RECT 120.725 170.295 120.985 170.750 ;
        RECT 121.155 170.465 121.415 170.945 ;
        RECT 121.595 170.295 121.855 170.750 ;
        RECT 122.025 170.465 122.275 170.945 ;
        RECT 122.455 170.295 122.715 170.750 ;
        RECT 122.885 170.465 123.135 170.945 ;
        RECT 123.315 170.295 123.575 170.750 ;
        RECT 123.745 170.465 123.990 170.945 ;
        RECT 124.160 170.295 124.435 170.750 ;
        RECT 124.605 170.465 124.850 170.945 ;
        RECT 125.020 170.295 125.280 170.750 ;
        RECT 125.450 170.465 125.710 170.945 ;
        RECT 125.880 170.295 126.140 170.750 ;
        RECT 126.310 170.465 126.570 170.945 ;
        RECT 126.740 170.295 127.000 170.750 ;
        RECT 127.170 170.385 127.430 170.945 ;
        RECT 113.160 170.125 119.905 170.295 ;
        RECT 111.450 169.705 118.570 169.955 ;
        RECT 108.205 169.365 109.235 169.535 ;
        RECT 110.025 169.445 110.780 169.615 ;
        RECT 108.205 168.565 108.515 169.365 ;
        RECT 110.025 169.195 110.285 169.445 ;
        RECT 108.685 168.395 108.995 169.195 ;
        RECT 109.165 169.025 110.285 169.195 ;
        RECT 109.165 168.565 109.425 169.025 ;
        RECT 109.595 168.395 109.850 168.855 ;
        RECT 110.025 168.565 110.285 169.025 ;
        RECT 110.455 168.395 110.740 169.265 ;
        RECT 110.975 168.395 111.270 169.205 ;
        RECT 111.450 168.565 111.695 169.705 ;
        RECT 111.870 168.395 112.130 169.205 ;
        RECT 112.310 168.570 112.560 169.705 ;
        RECT 118.740 169.535 119.905 170.125 ;
        RECT 120.255 170.125 127.000 170.295 ;
        RECT 120.255 169.925 121.420 170.125 ;
        RECT 127.600 169.955 127.850 170.765 ;
        RECT 128.030 170.420 128.290 170.945 ;
        RECT 128.460 169.955 128.710 170.765 ;
        RECT 128.890 170.435 129.195 170.945 ;
        RECT 120.225 169.755 121.420 169.925 ;
        RECT 113.160 169.310 119.905 169.535 ;
        RECT 120.255 169.535 121.420 169.755 ;
        RECT 121.590 169.705 128.710 169.955 ;
        RECT 128.880 169.705 129.195 170.265 ;
        RECT 130.285 170.220 130.575 170.945 ;
        RECT 120.255 169.310 127.000 169.535 ;
        RECT 113.160 169.295 118.565 169.310 ;
        RECT 112.730 168.400 112.990 169.195 ;
        RECT 113.160 168.570 113.420 169.295 ;
        RECT 113.590 168.400 113.850 169.125 ;
        RECT 114.020 168.570 114.280 169.295 ;
        RECT 114.450 168.400 114.710 169.125 ;
        RECT 114.880 168.570 115.140 169.295 ;
        RECT 115.310 168.400 115.570 169.125 ;
        RECT 115.740 168.570 116.000 169.295 ;
        RECT 116.170 168.400 116.415 169.125 ;
        RECT 116.585 168.570 116.845 169.295 ;
        RECT 117.030 168.400 117.275 169.125 ;
        RECT 117.445 168.570 117.705 169.295 ;
        RECT 117.890 168.400 118.135 169.125 ;
        RECT 118.305 168.570 118.565 169.295 ;
        RECT 118.750 168.400 119.005 169.125 ;
        RECT 119.175 168.570 119.465 169.310 ;
        RECT 112.730 168.395 119.005 168.400 ;
        RECT 119.635 168.395 119.905 169.140 ;
        RECT 120.255 168.395 120.525 169.140 ;
        RECT 120.695 168.570 120.985 169.310 ;
        RECT 121.595 169.295 127.000 169.310 ;
        RECT 121.155 168.400 121.410 169.125 ;
        RECT 121.595 168.570 121.855 169.295 ;
        RECT 122.025 168.400 122.270 169.125 ;
        RECT 122.455 168.570 122.715 169.295 ;
        RECT 122.885 168.400 123.130 169.125 ;
        RECT 123.315 168.570 123.575 169.295 ;
        RECT 123.745 168.400 123.990 169.125 ;
        RECT 124.160 168.570 124.420 169.295 ;
        RECT 124.590 168.400 124.850 169.125 ;
        RECT 125.020 168.570 125.280 169.295 ;
        RECT 125.450 168.400 125.710 169.125 ;
        RECT 125.880 168.570 126.140 169.295 ;
        RECT 126.310 168.400 126.570 169.125 ;
        RECT 126.740 168.570 127.000 169.295 ;
        RECT 127.170 168.400 127.430 169.195 ;
        RECT 127.600 168.570 127.850 169.705 ;
        RECT 121.155 168.395 127.430 168.400 ;
        RECT 128.030 168.395 128.290 169.205 ;
        RECT 128.465 168.565 128.710 169.705 ;
        RECT 128.890 168.395 129.185 169.205 ;
        RECT 130.285 168.395 130.575 169.560 ;
        RECT 130.765 169.365 130.995 170.705 ;
        RECT 131.175 169.865 131.405 170.765 ;
        RECT 131.605 170.165 131.850 170.945 ;
        RECT 132.020 170.405 132.450 170.765 ;
        RECT 133.030 170.575 133.760 170.945 ;
        RECT 132.020 170.215 133.760 170.405 ;
        RECT 132.020 169.985 132.240 170.215 ;
        RECT 131.175 169.185 131.515 169.865 ;
        RECT 130.765 168.985 131.515 169.185 ;
        RECT 131.695 169.685 132.240 169.985 ;
        RECT 130.765 168.595 131.005 168.985 ;
        RECT 131.175 168.395 131.525 168.805 ;
        RECT 131.695 168.575 132.025 169.685 ;
        RECT 132.410 169.415 132.835 170.035 ;
        RECT 133.030 169.415 133.290 170.035 ;
        RECT 133.500 169.705 133.760 170.215 ;
        RECT 132.195 169.045 133.220 169.245 ;
        RECT 132.195 168.575 132.375 169.045 ;
        RECT 132.545 168.395 132.875 168.875 ;
        RECT 133.050 168.575 133.220 169.045 ;
        RECT 133.485 168.395 133.770 169.535 ;
        RECT 133.960 168.575 134.240 170.765 ;
        RECT 134.445 169.365 134.675 170.705 ;
        RECT 134.855 169.865 135.085 170.765 ;
        RECT 135.285 170.165 135.530 170.945 ;
        RECT 135.700 170.405 136.130 170.765 ;
        RECT 136.710 170.575 137.440 170.945 ;
        RECT 135.700 170.215 137.440 170.405 ;
        RECT 135.700 169.985 135.920 170.215 ;
        RECT 134.855 169.185 135.195 169.865 ;
        RECT 134.445 168.985 135.195 169.185 ;
        RECT 135.375 169.685 135.920 169.985 ;
        RECT 134.445 168.595 134.685 168.985 ;
        RECT 134.855 168.395 135.205 168.805 ;
        RECT 135.375 168.575 135.705 169.685 ;
        RECT 136.090 169.415 136.515 170.035 ;
        RECT 136.710 169.415 136.970 170.035 ;
        RECT 137.180 169.705 137.440 170.215 ;
        RECT 135.875 169.045 136.900 169.245 ;
        RECT 135.875 168.575 136.055 169.045 ;
        RECT 136.225 168.395 136.555 168.875 ;
        RECT 136.730 168.575 136.900 169.045 ;
        RECT 137.165 168.395 137.450 169.535 ;
        RECT 137.640 168.575 137.920 170.765 ;
        RECT 138.565 170.195 139.775 170.945 ;
        RECT 138.565 169.485 139.085 170.025 ;
        RECT 139.255 169.655 139.775 170.195 ;
        RECT 138.565 168.395 139.775 169.485 ;
        RECT 27.160 168.225 139.860 168.395 ;
        RECT 27.245 167.135 28.455 168.225 ;
        RECT 28.625 167.790 33.970 168.225 ;
        RECT 34.145 167.790 39.490 168.225 ;
        RECT 27.245 166.425 27.765 166.965 ;
        RECT 27.935 166.595 28.455 167.135 ;
        RECT 27.245 165.675 28.455 166.425 ;
        RECT 30.210 166.220 30.550 167.050 ;
        RECT 32.030 166.540 32.380 167.790 ;
        RECT 35.730 166.220 36.070 167.050 ;
        RECT 37.550 166.540 37.900 167.790 ;
        RECT 40.125 167.060 40.415 168.225 ;
        RECT 41.585 167.295 41.765 168.055 ;
        RECT 41.945 167.465 42.275 168.225 ;
        RECT 41.585 167.125 42.260 167.295 ;
        RECT 42.445 167.150 42.715 168.055 ;
        RECT 42.090 166.980 42.260 167.125 ;
        RECT 41.525 166.575 41.865 166.945 ;
        RECT 42.090 166.650 42.365 166.980 ;
        RECT 28.625 165.675 33.970 166.220 ;
        RECT 34.145 165.675 39.490 166.220 ;
        RECT 40.125 165.675 40.415 166.400 ;
        RECT 42.090 166.395 42.260 166.650 ;
        RECT 41.595 166.225 42.260 166.395 ;
        RECT 42.535 166.350 42.715 167.150 ;
        RECT 42.885 167.135 44.555 168.225 ;
        RECT 41.595 165.845 41.765 166.225 ;
        RECT 41.945 165.675 42.275 166.055 ;
        RECT 42.455 165.845 42.715 166.350 ;
        RECT 42.885 166.445 43.635 166.965 ;
        RECT 43.805 166.615 44.555 167.135 ;
        RECT 44.815 167.295 44.985 168.055 ;
        RECT 45.165 167.465 45.495 168.225 ;
        RECT 44.815 167.125 45.480 167.295 ;
        RECT 45.665 167.150 45.935 168.055 ;
        RECT 45.310 166.980 45.480 167.125 ;
        RECT 44.745 166.575 45.075 166.945 ;
        RECT 45.310 166.650 45.595 166.980 ;
        RECT 42.885 165.675 44.555 166.445 ;
        RECT 45.310 166.395 45.480 166.650 ;
        RECT 44.815 166.225 45.480 166.395 ;
        RECT 45.765 166.350 45.935 167.150 ;
        RECT 46.105 167.135 47.775 168.225 ;
        RECT 44.815 165.845 44.985 166.225 ;
        RECT 45.165 165.675 45.495 166.055 ;
        RECT 45.675 165.845 45.935 166.350 ;
        RECT 46.105 166.445 46.855 166.965 ;
        RECT 47.025 166.615 47.775 167.135 ;
        RECT 48.035 167.295 48.205 168.055 ;
        RECT 48.420 167.465 48.750 168.225 ;
        RECT 48.035 167.125 48.750 167.295 ;
        RECT 48.920 167.150 49.175 168.055 ;
        RECT 47.945 166.575 48.300 166.945 ;
        RECT 48.580 166.915 48.750 167.125 ;
        RECT 48.580 166.585 48.835 166.915 ;
        RECT 46.105 165.675 47.775 166.445 ;
        RECT 48.580 166.395 48.750 166.585 ;
        RECT 49.005 166.420 49.175 167.150 ;
        RECT 49.350 167.075 49.610 168.225 ;
        RECT 50.325 167.295 50.505 168.055 ;
        RECT 50.685 167.465 51.015 168.225 ;
        RECT 50.325 167.125 51.000 167.295 ;
        RECT 51.185 167.150 51.455 168.055 ;
        RECT 50.830 166.980 51.000 167.125 ;
        RECT 50.265 166.575 50.605 166.945 ;
        RECT 50.830 166.650 51.105 166.980 ;
        RECT 48.035 166.225 48.750 166.395 ;
        RECT 48.035 165.845 48.205 166.225 ;
        RECT 48.420 165.675 48.750 166.055 ;
        RECT 48.920 165.845 49.175 166.420 ;
        RECT 49.350 165.675 49.610 166.515 ;
        RECT 50.830 166.395 51.000 166.650 ;
        RECT 50.335 166.225 51.000 166.395 ;
        RECT 51.275 166.350 51.455 167.150 ;
        RECT 51.705 167.295 51.885 168.055 ;
        RECT 52.065 167.465 52.395 168.225 ;
        RECT 51.705 167.125 52.380 167.295 ;
        RECT 52.565 167.150 52.835 168.055 ;
        RECT 52.210 166.980 52.380 167.125 ;
        RECT 51.645 166.575 51.985 166.945 ;
        RECT 52.210 166.650 52.485 166.980 ;
        RECT 52.210 166.395 52.380 166.650 ;
        RECT 50.335 165.845 50.505 166.225 ;
        RECT 50.685 165.675 51.015 166.055 ;
        RECT 51.195 165.845 51.455 166.350 ;
        RECT 51.715 166.225 52.380 166.395 ;
        RECT 52.655 166.350 52.835 167.150 ;
        RECT 53.005 167.060 53.295 168.225 ;
        RECT 54.465 167.295 54.645 168.055 ;
        RECT 54.825 167.465 55.155 168.225 ;
        RECT 54.465 167.125 55.140 167.295 ;
        RECT 55.325 167.150 55.595 168.055 ;
        RECT 54.970 166.980 55.140 167.125 ;
        RECT 54.405 166.575 54.745 166.945 ;
        RECT 54.970 166.650 55.245 166.980 ;
        RECT 51.715 165.845 51.885 166.225 ;
        RECT 52.065 165.675 52.395 166.055 ;
        RECT 52.575 165.845 52.835 166.350 ;
        RECT 53.005 165.675 53.295 166.400 ;
        RECT 54.970 166.395 55.140 166.650 ;
        RECT 54.475 166.225 55.140 166.395 ;
        RECT 55.415 166.350 55.595 167.150 ;
        RECT 54.475 165.845 54.645 166.225 ;
        RECT 54.825 165.675 55.155 166.055 ;
        RECT 55.335 165.845 55.595 166.350 ;
        RECT 55.765 167.625 56.025 168.045 ;
        RECT 56.195 167.795 56.525 168.225 ;
        RECT 57.190 167.795 57.935 167.965 ;
        RECT 55.765 167.455 57.595 167.625 ;
        RECT 55.765 166.415 55.935 167.455 ;
        RECT 56.105 166.585 56.455 167.285 ;
        RECT 56.670 167.115 57.255 167.285 ;
        RECT 56.625 166.585 56.915 166.915 ;
        RECT 57.085 166.835 57.255 167.115 ;
        RECT 57.425 167.175 57.595 167.455 ;
        RECT 57.765 167.545 57.935 167.795 ;
        RECT 58.160 167.715 58.800 168.045 ;
        RECT 57.765 167.375 58.800 167.545 ;
        RECT 58.970 167.425 59.250 168.225 ;
        RECT 58.630 167.255 58.800 167.375 ;
        RECT 57.425 167.005 58.075 167.175 ;
        RECT 58.630 167.085 59.290 167.255 ;
        RECT 59.460 167.085 59.735 168.055 ;
        RECT 57.085 166.665 57.510 166.835 ;
        RECT 57.085 166.415 57.255 166.665 ;
        RECT 57.905 166.585 58.075 167.005 ;
        RECT 59.120 166.915 59.290 167.085 ;
        RECT 58.295 166.585 58.950 166.915 ;
        RECT 59.120 166.585 59.395 166.915 ;
        RECT 59.120 166.415 59.290 166.585 ;
        RECT 55.765 166.040 56.080 166.415 ;
        RECT 56.335 165.675 56.505 166.415 ;
        RECT 56.755 166.245 57.255 166.415 ;
        RECT 57.695 166.245 59.290 166.415 ;
        RECT 59.565 166.350 59.735 167.085 ;
        RECT 59.910 167.075 60.170 168.225 ;
        RECT 60.345 167.150 60.600 168.055 ;
        RECT 60.770 167.465 61.100 168.225 ;
        RECT 61.315 167.295 61.485 168.055 ;
        RECT 56.755 166.040 56.925 166.245 ;
        RECT 57.150 165.675 57.525 166.075 ;
        RECT 57.695 165.895 57.865 166.245 ;
        RECT 58.050 165.675 58.380 166.075 ;
        RECT 58.550 165.895 58.720 166.245 ;
        RECT 58.890 165.675 59.270 166.075 ;
        RECT 59.460 166.005 59.735 166.350 ;
        RECT 59.910 165.675 60.170 166.515 ;
        RECT 60.345 166.420 60.515 167.150 ;
        RECT 60.770 167.125 61.485 167.295 ;
        RECT 61.745 167.255 62.015 168.025 ;
        RECT 62.185 167.445 62.515 168.225 ;
        RECT 62.720 167.620 62.905 168.025 ;
        RECT 63.075 167.800 63.410 168.225 ;
        RECT 62.720 167.445 63.385 167.620 ;
        RECT 60.770 166.915 60.940 167.125 ;
        RECT 61.745 167.085 62.875 167.255 ;
        RECT 60.685 166.585 60.940 166.915 ;
        RECT 60.345 165.845 60.600 166.420 ;
        RECT 60.770 166.395 60.940 166.585 ;
        RECT 61.220 166.575 61.575 166.945 ;
        RECT 60.770 166.225 61.485 166.395 ;
        RECT 60.770 165.675 61.100 166.055 ;
        RECT 61.315 165.845 61.485 166.225 ;
        RECT 61.745 166.175 61.915 167.085 ;
        RECT 62.085 166.335 62.445 166.915 ;
        RECT 62.625 166.585 62.875 167.085 ;
        RECT 63.045 166.415 63.385 167.445 ;
        RECT 64.585 167.295 64.765 168.055 ;
        RECT 64.945 167.465 65.275 168.225 ;
        RECT 64.585 167.125 65.260 167.295 ;
        RECT 65.445 167.150 65.715 168.055 ;
        RECT 65.090 166.980 65.260 167.125 ;
        RECT 64.525 166.575 64.865 166.945 ;
        RECT 65.090 166.650 65.365 166.980 ;
        RECT 62.700 166.245 63.385 166.415 ;
        RECT 65.090 166.395 65.260 166.650 ;
        RECT 61.745 165.845 62.005 166.175 ;
        RECT 62.215 165.675 62.490 166.155 ;
        RECT 62.700 165.845 62.905 166.245 ;
        RECT 64.595 166.225 65.260 166.395 ;
        RECT 65.535 166.350 65.715 167.150 ;
        RECT 65.885 167.060 66.175 168.225 ;
        RECT 66.350 167.075 66.610 168.225 ;
        RECT 66.785 167.150 67.040 168.055 ;
        RECT 67.210 167.465 67.540 168.225 ;
        RECT 67.755 167.295 67.925 168.055 ;
        RECT 63.075 165.675 63.410 166.075 ;
        RECT 64.595 165.845 64.765 166.225 ;
        RECT 64.945 165.675 65.275 166.055 ;
        RECT 65.455 165.845 65.715 166.350 ;
        RECT 65.885 165.675 66.175 166.400 ;
        RECT 66.350 165.675 66.610 166.515 ;
        RECT 66.785 166.420 66.955 167.150 ;
        RECT 67.210 167.125 67.925 167.295 ;
        RECT 69.195 167.295 69.365 168.055 ;
        RECT 69.545 167.465 69.875 168.225 ;
        RECT 69.195 167.125 69.860 167.295 ;
        RECT 70.045 167.150 70.315 168.055 ;
        RECT 67.210 166.915 67.380 167.125 ;
        RECT 69.690 166.980 69.860 167.125 ;
        RECT 67.125 166.585 67.380 166.915 ;
        RECT 66.785 165.845 67.040 166.420 ;
        RECT 67.210 166.395 67.380 166.585 ;
        RECT 67.660 166.575 68.015 166.945 ;
        RECT 69.125 166.575 69.455 166.945 ;
        RECT 69.690 166.650 69.975 166.980 ;
        RECT 69.690 166.395 69.860 166.650 ;
        RECT 67.210 166.225 67.925 166.395 ;
        RECT 67.210 165.675 67.540 166.055 ;
        RECT 67.755 165.845 67.925 166.225 ;
        RECT 69.195 166.225 69.860 166.395 ;
        RECT 70.145 166.350 70.315 167.150 ;
        RECT 70.565 167.295 70.745 168.055 ;
        RECT 70.925 167.465 71.255 168.225 ;
        RECT 70.565 167.125 71.240 167.295 ;
        RECT 71.425 167.150 71.695 168.055 ;
        RECT 71.070 166.980 71.240 167.125 ;
        RECT 70.505 166.575 70.845 166.945 ;
        RECT 71.070 166.650 71.345 166.980 ;
        RECT 71.070 166.395 71.240 166.650 ;
        RECT 69.195 165.845 69.365 166.225 ;
        RECT 69.545 165.675 69.875 166.055 ;
        RECT 70.055 165.845 70.315 166.350 ;
        RECT 70.575 166.225 71.240 166.395 ;
        RECT 71.515 166.350 71.695 167.150 ;
        RECT 71.875 167.085 72.205 168.225 ;
        RECT 72.735 167.255 73.065 168.040 ;
        RECT 72.385 167.085 73.065 167.255 ;
        RECT 73.325 167.295 73.505 168.055 ;
        RECT 73.685 167.465 74.015 168.225 ;
        RECT 73.325 167.125 74.000 167.295 ;
        RECT 74.185 167.150 74.455 168.055 ;
        RECT 71.865 166.665 72.215 166.915 ;
        RECT 72.385 166.485 72.555 167.085 ;
        RECT 73.830 166.980 74.000 167.125 ;
        RECT 72.725 166.665 73.075 166.915 ;
        RECT 73.265 166.575 73.605 166.945 ;
        RECT 73.830 166.650 74.105 166.980 ;
        RECT 70.575 165.845 70.745 166.225 ;
        RECT 70.925 165.675 71.255 166.055 ;
        RECT 71.435 165.845 71.695 166.350 ;
        RECT 71.875 165.675 72.145 166.485 ;
        RECT 72.315 165.845 72.645 166.485 ;
        RECT 72.815 165.675 73.055 166.485 ;
        RECT 73.830 166.395 74.000 166.650 ;
        RECT 73.335 166.225 74.000 166.395 ;
        RECT 74.275 166.350 74.455 167.150 ;
        RECT 74.705 167.295 74.885 168.055 ;
        RECT 75.065 167.465 75.395 168.225 ;
        RECT 74.705 167.125 75.380 167.295 ;
        RECT 75.565 167.150 75.835 168.055 ;
        RECT 75.210 166.980 75.380 167.125 ;
        RECT 74.645 166.575 74.985 166.945 ;
        RECT 75.210 166.650 75.485 166.980 ;
        RECT 75.210 166.395 75.380 166.650 ;
        RECT 73.335 165.845 73.505 166.225 ;
        RECT 73.685 165.675 74.015 166.055 ;
        RECT 74.195 165.845 74.455 166.350 ;
        RECT 74.715 166.225 75.380 166.395 ;
        RECT 75.655 166.350 75.835 167.150 ;
        RECT 76.085 167.295 76.265 168.055 ;
        RECT 76.445 167.465 76.775 168.225 ;
        RECT 76.085 167.125 76.760 167.295 ;
        RECT 76.945 167.150 77.215 168.055 ;
        RECT 76.590 166.980 76.760 167.125 ;
        RECT 76.025 166.575 76.365 166.945 ;
        RECT 76.590 166.650 76.865 166.980 ;
        RECT 76.590 166.395 76.760 166.650 ;
        RECT 74.715 165.845 74.885 166.225 ;
        RECT 75.065 165.675 75.395 166.055 ;
        RECT 75.575 165.845 75.835 166.350 ;
        RECT 76.095 166.225 76.760 166.395 ;
        RECT 77.035 166.350 77.215 167.150 ;
        RECT 77.465 167.295 77.645 168.055 ;
        RECT 77.825 167.465 78.155 168.225 ;
        RECT 77.465 167.125 78.140 167.295 ;
        RECT 78.325 167.150 78.595 168.055 ;
        RECT 77.970 166.980 78.140 167.125 ;
        RECT 77.405 166.575 77.745 166.945 ;
        RECT 77.970 166.650 78.245 166.980 ;
        RECT 77.970 166.395 78.140 166.650 ;
        RECT 76.095 165.845 76.265 166.225 ;
        RECT 76.445 165.675 76.775 166.055 ;
        RECT 76.955 165.845 77.215 166.350 ;
        RECT 77.475 166.225 78.140 166.395 ;
        RECT 78.415 166.350 78.595 167.150 ;
        RECT 78.765 167.060 79.055 168.225 ;
        RECT 80.235 167.295 80.405 168.055 ;
        RECT 80.620 167.465 80.950 168.225 ;
        RECT 80.235 167.125 80.950 167.295 ;
        RECT 81.120 167.150 81.375 168.055 ;
        RECT 80.145 166.575 80.500 166.945 ;
        RECT 80.780 166.915 80.950 167.125 ;
        RECT 80.780 166.585 81.035 166.915 ;
        RECT 77.475 165.845 77.645 166.225 ;
        RECT 77.825 165.675 78.155 166.055 ;
        RECT 78.335 165.845 78.595 166.350 ;
        RECT 78.765 165.675 79.055 166.400 ;
        RECT 80.780 166.395 80.950 166.585 ;
        RECT 81.205 166.420 81.375 167.150 ;
        RECT 81.550 167.075 81.810 168.225 ;
        RECT 81.990 167.075 82.250 168.225 ;
        RECT 82.425 167.150 82.680 168.055 ;
        RECT 82.850 167.465 83.180 168.225 ;
        RECT 83.395 167.295 83.565 168.055 ;
        RECT 84.320 167.425 84.570 168.225 ;
        RECT 84.740 167.595 85.070 168.055 ;
        RECT 85.240 167.765 85.455 168.225 ;
        RECT 84.740 167.425 85.910 167.595 ;
        RECT 80.235 166.225 80.950 166.395 ;
        RECT 80.235 165.845 80.405 166.225 ;
        RECT 80.620 165.675 80.950 166.055 ;
        RECT 81.120 165.845 81.375 166.420 ;
        RECT 81.550 165.675 81.810 166.515 ;
        RECT 81.990 165.675 82.250 166.515 ;
        RECT 82.425 166.420 82.595 167.150 ;
        RECT 82.850 167.125 83.565 167.295 ;
        RECT 83.830 167.255 84.110 167.415 ;
        RECT 82.850 166.915 83.020 167.125 ;
        RECT 83.830 167.085 85.165 167.255 ;
        RECT 82.765 166.585 83.020 166.915 ;
        RECT 82.425 165.845 82.680 166.420 ;
        RECT 82.850 166.395 83.020 166.585 ;
        RECT 83.300 166.575 83.655 166.945 ;
        RECT 84.995 166.915 85.165 167.085 ;
        RECT 83.830 166.665 84.180 166.905 ;
        RECT 84.350 166.665 84.825 166.905 ;
        RECT 84.995 166.665 85.370 166.915 ;
        RECT 84.995 166.495 85.165 166.665 ;
        RECT 82.850 166.225 83.565 166.395 ;
        RECT 82.850 165.675 83.180 166.055 ;
        RECT 83.395 165.845 83.565 166.225 ;
        RECT 83.830 166.325 85.165 166.495 ;
        RECT 83.830 166.115 84.100 166.325 ;
        RECT 85.540 166.135 85.910 167.425 ;
        RECT 86.145 167.335 86.405 168.045 ;
        RECT 86.575 167.515 86.905 168.225 ;
        RECT 87.075 167.335 87.305 168.045 ;
        RECT 86.145 167.095 87.305 167.335 ;
        RECT 87.485 167.315 87.755 168.045 ;
        RECT 87.935 167.495 88.275 168.225 ;
        RECT 87.485 167.095 88.255 167.315 ;
        RECT 86.135 166.585 86.435 166.915 ;
        RECT 86.615 166.605 87.140 166.915 ;
        RECT 87.320 166.605 87.785 166.915 ;
        RECT 84.320 165.675 84.650 166.135 ;
        RECT 85.160 165.845 85.910 166.135 ;
        RECT 86.145 165.675 86.435 166.405 ;
        RECT 86.615 165.965 86.845 166.605 ;
        RECT 87.965 166.425 88.255 167.095 ;
        RECT 87.025 166.225 88.255 166.425 ;
        RECT 87.025 165.855 87.335 166.225 ;
        RECT 87.515 165.675 88.185 166.045 ;
        RECT 88.445 165.855 88.705 168.045 ;
        RECT 88.885 167.215 89.145 168.225 ;
        RECT 89.315 167.385 89.590 168.055 ;
        RECT 89.315 167.035 89.485 167.385 ;
        RECT 89.790 167.380 90.005 168.225 ;
        RECT 90.190 167.715 90.665 168.055 ;
        RECT 90.845 167.720 91.475 168.225 ;
        RECT 90.845 167.545 91.035 167.720 ;
        RECT 90.230 167.185 90.480 167.480 ;
        RECT 90.705 167.355 91.035 167.545 ;
        RECT 91.205 167.185 91.460 167.550 ;
        RECT 88.885 166.515 89.500 167.035 ;
        RECT 89.670 167.015 91.460 167.185 ;
        RECT 91.645 167.060 91.935 168.225 ;
        RECT 92.655 167.480 92.925 168.225 ;
        RECT 93.555 168.220 99.830 168.225 ;
        RECT 93.095 167.310 93.385 168.050 ;
        RECT 93.555 167.495 93.810 168.220 ;
        RECT 93.995 167.325 94.255 168.050 ;
        RECT 94.425 167.495 94.670 168.220 ;
        RECT 94.855 167.325 95.115 168.050 ;
        RECT 95.285 167.495 95.530 168.220 ;
        RECT 95.715 167.325 95.975 168.050 ;
        RECT 96.145 167.495 96.390 168.220 ;
        RECT 96.560 167.325 96.820 168.050 ;
        RECT 96.990 167.495 97.250 168.220 ;
        RECT 97.420 167.325 97.680 168.050 ;
        RECT 97.850 167.495 98.110 168.220 ;
        RECT 98.280 167.325 98.540 168.050 ;
        RECT 98.710 167.495 98.970 168.220 ;
        RECT 99.140 167.325 99.400 168.050 ;
        RECT 99.570 167.425 99.830 168.220 ;
        RECT 93.995 167.310 99.400 167.325 ;
        RECT 92.655 167.085 99.400 167.310 ;
        RECT 89.670 166.585 89.900 167.015 ;
        RECT 88.885 165.675 89.160 166.335 ;
        RECT 89.330 166.305 89.500 166.515 ;
        RECT 90.085 166.340 90.495 166.835 ;
        RECT 89.330 165.845 89.580 166.305 ;
        RECT 89.755 165.675 90.085 166.170 ;
        RECT 90.265 165.895 90.495 166.340 ;
        RECT 90.665 166.160 90.920 167.015 ;
        RECT 91.090 166.355 91.475 166.835 ;
        RECT 92.655 166.495 93.820 167.085 ;
        RECT 100.000 166.915 100.250 168.050 ;
        RECT 100.430 167.415 100.690 168.225 ;
        RECT 100.865 166.915 101.110 168.055 ;
        RECT 101.290 167.415 101.585 168.225 ;
        RECT 101.765 167.085 102.055 168.225 ;
        RECT 102.225 167.505 102.675 168.055 ;
        RECT 102.865 167.505 103.195 168.225 ;
        RECT 93.990 166.665 101.110 166.915 ;
        RECT 90.665 165.895 91.455 166.160 ;
        RECT 91.645 165.675 91.935 166.400 ;
        RECT 92.655 166.325 99.400 166.495 ;
        RECT 92.655 165.675 92.955 166.155 ;
        RECT 93.125 165.870 93.385 166.325 ;
        RECT 93.555 165.675 93.815 166.155 ;
        RECT 93.995 165.870 94.255 166.325 ;
        RECT 94.425 165.675 94.675 166.155 ;
        RECT 94.855 165.870 95.115 166.325 ;
        RECT 95.285 165.675 95.535 166.155 ;
        RECT 95.715 165.870 95.975 166.325 ;
        RECT 96.145 165.675 96.390 166.155 ;
        RECT 96.560 165.870 96.835 166.325 ;
        RECT 97.005 165.675 97.250 166.155 ;
        RECT 97.420 165.870 97.680 166.325 ;
        RECT 97.850 165.675 98.110 166.155 ;
        RECT 98.280 165.870 98.540 166.325 ;
        RECT 98.710 165.675 98.970 166.155 ;
        RECT 99.140 165.870 99.400 166.325 ;
        RECT 99.570 165.675 99.830 166.235 ;
        RECT 100.000 165.855 100.250 166.665 ;
        RECT 100.430 165.675 100.690 166.200 ;
        RECT 100.860 165.855 101.110 166.665 ;
        RECT 101.280 166.355 101.595 166.915 ;
        RECT 101.290 165.675 101.595 166.185 ;
        RECT 101.765 165.675 102.055 166.475 ;
        RECT 102.225 166.135 102.475 167.505 ;
        RECT 103.405 167.335 103.705 167.885 ;
        RECT 103.875 167.555 104.155 168.225 ;
        RECT 102.765 167.165 103.705 167.335 ;
        RECT 102.765 166.915 102.935 167.165 ;
        RECT 104.040 166.915 104.355 167.355 ;
        RECT 104.525 167.060 104.815 168.225 ;
        RECT 105.045 167.525 105.265 168.055 ;
        RECT 105.435 167.715 105.765 168.225 ;
        RECT 105.935 167.525 106.160 168.055 ;
        RECT 105.045 167.260 106.160 167.525 ;
        RECT 106.330 167.510 106.645 168.055 ;
        RECT 106.835 167.810 107.165 168.225 ;
        RECT 106.330 167.280 107.165 167.510 ;
        RECT 102.645 166.585 102.935 166.915 ;
        RECT 103.105 166.665 103.435 166.915 ;
        RECT 103.665 166.665 104.355 166.915 ;
        RECT 102.765 166.495 102.935 166.585 ;
        RECT 102.765 166.305 104.155 166.495 ;
        RECT 102.225 165.845 102.775 166.135 ;
        RECT 102.945 165.675 103.195 166.135 ;
        RECT 103.825 165.945 104.155 166.305 ;
        RECT 104.525 165.675 104.815 166.400 ;
        RECT 104.995 166.340 105.310 166.915 ;
        RECT 104.985 165.675 105.315 166.155 ;
        RECT 105.500 165.955 105.880 166.915 ;
        RECT 106.330 166.585 106.655 167.000 ;
        RECT 106.825 166.585 107.165 167.280 ;
        RECT 106.825 166.415 106.995 166.585 ;
        RECT 107.335 166.415 107.565 168.055 ;
        RECT 107.735 167.255 108.025 168.225 ;
        RECT 108.210 167.835 108.545 168.055 ;
        RECT 109.550 167.845 109.905 168.225 ;
        RECT 108.210 167.215 108.465 167.835 ;
        RECT 108.715 167.675 108.945 167.715 ;
        RECT 110.075 167.675 110.325 168.055 ;
        RECT 108.715 167.475 110.325 167.675 ;
        RECT 108.715 167.385 108.900 167.475 ;
        RECT 109.490 167.465 110.325 167.475 ;
        RECT 110.575 167.445 110.825 168.225 ;
        RECT 110.995 167.375 111.255 168.055 ;
        RECT 109.055 167.275 109.385 167.305 ;
        RECT 109.055 167.215 110.855 167.275 ;
        RECT 108.210 167.105 110.915 167.215 ;
        RECT 108.210 167.045 109.385 167.105 ;
        RECT 110.715 167.070 110.915 167.105 ;
        RECT 108.205 166.665 108.695 166.865 ;
        RECT 108.885 166.665 109.360 166.875 ;
        RECT 106.255 166.245 106.995 166.415 ;
        RECT 106.255 165.845 106.445 166.245 ;
        RECT 107.165 166.225 107.565 166.415 ;
        RECT 106.665 165.675 106.995 166.035 ;
        RECT 107.165 165.845 107.355 166.225 ;
        RECT 107.525 165.675 107.855 166.055 ;
        RECT 108.210 165.675 108.665 166.440 ;
        RECT 109.140 166.265 109.360 166.665 ;
        RECT 109.605 166.665 109.935 166.875 ;
        RECT 109.605 166.265 109.815 166.665 ;
        RECT 110.105 166.630 110.515 166.935 ;
        RECT 110.745 166.495 110.915 167.070 ;
        RECT 110.645 166.375 110.915 166.495 ;
        RECT 110.070 166.330 110.915 166.375 ;
        RECT 110.070 166.205 110.825 166.330 ;
        RECT 110.070 166.055 110.240 166.205 ;
        RECT 111.085 166.175 111.255 167.375 ;
        RECT 108.940 165.845 110.240 166.055 ;
        RECT 110.495 165.675 110.825 166.035 ;
        RECT 110.995 165.845 111.255 166.175 ;
        RECT 111.425 165.955 111.705 168.055 ;
        RECT 111.895 167.465 112.680 168.225 ;
        RECT 113.075 167.395 113.460 168.055 ;
        RECT 113.075 167.295 113.485 167.395 ;
        RECT 111.875 167.085 113.485 167.295 ;
        RECT 113.785 167.205 113.985 167.995 ;
        RECT 111.875 166.485 112.150 167.085 ;
        RECT 113.655 167.035 113.985 167.205 ;
        RECT 114.155 167.045 114.475 168.225 ;
        RECT 114.700 167.355 114.985 168.225 ;
        RECT 115.155 167.595 115.415 168.055 ;
        RECT 115.590 167.765 115.845 168.225 ;
        RECT 116.015 167.595 116.275 168.055 ;
        RECT 115.155 167.425 116.275 167.595 ;
        RECT 116.445 167.425 116.755 168.225 ;
        RECT 115.155 167.175 115.415 167.425 ;
        RECT 116.925 167.255 117.235 168.055 ;
        RECT 113.655 166.915 113.835 167.035 ;
        RECT 112.320 166.665 112.675 166.915 ;
        RECT 112.870 166.865 113.335 166.915 ;
        RECT 112.865 166.695 113.335 166.865 ;
        RECT 112.870 166.665 113.335 166.695 ;
        RECT 113.505 166.665 113.835 166.915 ;
        RECT 114.660 167.005 115.415 167.175 ;
        RECT 116.205 167.085 117.235 167.255 ;
        RECT 114.010 166.665 114.475 166.865 ;
        RECT 114.660 166.495 115.065 167.005 ;
        RECT 116.205 166.835 116.375 167.085 ;
        RECT 115.235 166.665 116.375 166.835 ;
        RECT 111.875 166.305 113.125 166.485 ;
        RECT 112.760 166.235 113.125 166.305 ;
        RECT 113.295 166.285 114.475 166.455 ;
        RECT 114.660 166.325 116.310 166.495 ;
        RECT 116.545 166.345 116.895 166.915 ;
        RECT 111.935 165.675 112.105 166.135 ;
        RECT 113.295 166.065 113.625 166.285 ;
        RECT 112.375 165.885 113.625 166.065 ;
        RECT 113.795 165.675 113.965 166.115 ;
        RECT 114.135 165.870 114.475 166.285 ;
        RECT 114.705 165.675 114.985 166.155 ;
        RECT 115.155 165.935 115.415 166.325 ;
        RECT 115.590 165.675 115.845 166.155 ;
        RECT 116.015 165.935 116.310 166.325 ;
        RECT 117.065 166.175 117.235 167.085 ;
        RECT 117.405 167.060 117.695 168.225 ;
        RECT 117.955 167.295 118.125 168.055 ;
        RECT 118.340 167.465 118.670 168.225 ;
        RECT 117.955 167.125 118.670 167.295 ;
        RECT 118.840 167.150 119.095 168.055 ;
        RECT 117.865 166.575 118.220 166.945 ;
        RECT 118.500 166.915 118.670 167.125 ;
        RECT 118.500 166.585 118.755 166.915 ;
        RECT 116.490 165.675 116.765 166.155 ;
        RECT 116.935 165.845 117.235 166.175 ;
        RECT 117.405 165.675 117.695 166.400 ;
        RECT 118.500 166.395 118.670 166.585 ;
        RECT 118.925 166.420 119.095 167.150 ;
        RECT 119.270 167.075 119.530 168.225 ;
        RECT 119.715 167.415 120.010 168.225 ;
        RECT 120.190 166.915 120.435 168.055 ;
        RECT 120.610 167.415 120.870 168.225 ;
        RECT 121.470 168.220 127.745 168.225 ;
        RECT 121.050 166.915 121.300 168.050 ;
        RECT 121.470 167.425 121.730 168.220 ;
        RECT 121.900 167.325 122.160 168.050 ;
        RECT 122.330 167.495 122.590 168.220 ;
        RECT 122.760 167.325 123.020 168.050 ;
        RECT 123.190 167.495 123.450 168.220 ;
        RECT 123.620 167.325 123.880 168.050 ;
        RECT 124.050 167.495 124.310 168.220 ;
        RECT 124.480 167.325 124.740 168.050 ;
        RECT 124.910 167.495 125.155 168.220 ;
        RECT 125.325 167.325 125.585 168.050 ;
        RECT 125.770 167.495 126.015 168.220 ;
        RECT 126.185 167.325 126.445 168.050 ;
        RECT 126.630 167.495 126.875 168.220 ;
        RECT 127.045 167.325 127.305 168.050 ;
        RECT 127.490 167.495 127.745 168.220 ;
        RECT 121.900 167.310 127.305 167.325 ;
        RECT 127.915 167.310 128.205 168.050 ;
        RECT 128.375 167.480 128.645 168.225 ;
        RECT 121.900 167.205 128.645 167.310 ;
        RECT 121.900 167.085 128.675 167.205 ;
        RECT 127.480 167.035 128.675 167.085 ;
        RECT 128.905 167.150 129.175 168.055 ;
        RECT 129.345 167.465 129.675 168.225 ;
        RECT 129.855 167.295 130.035 168.055 ;
        RECT 117.955 166.225 118.670 166.395 ;
        RECT 117.955 165.845 118.125 166.225 ;
        RECT 118.340 165.675 118.670 166.055 ;
        RECT 118.840 165.845 119.095 166.420 ;
        RECT 119.270 165.675 119.530 166.515 ;
        RECT 119.705 166.355 120.020 166.915 ;
        RECT 120.190 166.665 127.310 166.915 ;
        RECT 119.705 165.675 120.010 166.185 ;
        RECT 120.190 165.855 120.440 166.665 ;
        RECT 120.610 165.675 120.870 166.200 ;
        RECT 121.050 165.855 121.300 166.665 ;
        RECT 127.480 166.495 128.645 167.035 ;
        RECT 121.900 166.325 128.645 166.495 ;
        RECT 128.905 166.350 129.085 167.150 ;
        RECT 129.360 167.125 130.035 167.295 ;
        RECT 129.360 166.980 129.530 167.125 ;
        RECT 130.285 167.060 130.575 168.225 ;
        RECT 130.745 167.505 131.205 168.055 ;
        RECT 131.395 167.505 131.725 168.225 ;
        RECT 129.255 166.650 129.530 166.980 ;
        RECT 129.360 166.395 129.530 166.650 ;
        RECT 129.755 166.575 130.095 166.945 ;
        RECT 121.470 165.675 121.730 166.235 ;
        RECT 121.900 165.870 122.160 166.325 ;
        RECT 122.330 165.675 122.590 166.155 ;
        RECT 122.760 165.870 123.020 166.325 ;
        RECT 123.190 165.675 123.450 166.155 ;
        RECT 123.620 165.870 123.880 166.325 ;
        RECT 124.050 165.675 124.295 166.155 ;
        RECT 124.465 165.870 124.740 166.325 ;
        RECT 124.910 165.675 125.155 166.155 ;
        RECT 125.325 165.870 125.585 166.325 ;
        RECT 125.765 165.675 126.015 166.155 ;
        RECT 126.185 165.870 126.445 166.325 ;
        RECT 126.625 165.675 126.875 166.155 ;
        RECT 127.045 165.870 127.305 166.325 ;
        RECT 127.485 165.675 127.745 166.155 ;
        RECT 127.915 165.870 128.175 166.325 ;
        RECT 128.345 165.675 128.645 166.155 ;
        RECT 128.905 165.845 129.165 166.350 ;
        RECT 129.360 166.225 130.025 166.395 ;
        RECT 129.345 165.675 129.675 166.055 ;
        RECT 129.855 165.845 130.025 166.225 ;
        RECT 130.285 165.675 130.575 166.400 ;
        RECT 130.745 166.135 130.995 167.505 ;
        RECT 131.925 167.335 132.225 167.885 ;
        RECT 132.395 167.555 132.675 168.225 ;
        RECT 133.065 167.635 133.305 168.025 ;
        RECT 133.475 167.815 133.825 168.225 ;
        RECT 133.065 167.435 133.815 167.635 ;
        RECT 131.285 167.165 132.225 167.335 ;
        RECT 131.285 166.915 131.455 167.165 ;
        RECT 132.595 166.915 132.860 167.275 ;
        RECT 131.165 166.585 131.455 166.915 ;
        RECT 131.625 166.665 131.965 166.915 ;
        RECT 132.185 166.665 132.860 166.915 ;
        RECT 131.285 166.495 131.455 166.585 ;
        RECT 131.285 166.305 132.675 166.495 ;
        RECT 130.745 165.845 131.305 166.135 ;
        RECT 131.475 165.675 131.725 166.135 ;
        RECT 132.345 165.945 132.675 166.305 ;
        RECT 133.065 165.915 133.295 167.255 ;
        RECT 133.475 166.755 133.815 167.435 ;
        RECT 133.995 166.935 134.325 168.045 ;
        RECT 134.495 167.575 134.675 168.045 ;
        RECT 134.845 167.745 135.175 168.225 ;
        RECT 135.350 167.575 135.520 168.045 ;
        RECT 134.495 167.375 135.520 167.575 ;
        RECT 133.475 165.855 133.705 166.755 ;
        RECT 133.995 166.635 134.540 166.935 ;
        RECT 133.905 165.675 134.150 166.455 ;
        RECT 134.320 166.405 134.540 166.635 ;
        RECT 134.710 166.585 135.135 167.205 ;
        RECT 135.330 166.585 135.590 167.205 ;
        RECT 135.785 167.085 136.070 168.225 ;
        RECT 135.800 166.405 136.060 166.915 ;
        RECT 134.320 166.215 136.060 166.405 ;
        RECT 134.320 165.855 134.750 166.215 ;
        RECT 135.330 165.675 136.060 166.045 ;
        RECT 136.260 165.855 136.540 168.045 ;
        RECT 136.815 167.295 136.985 168.055 ;
        RECT 137.200 167.465 137.530 168.225 ;
        RECT 136.815 167.125 137.530 167.295 ;
        RECT 137.700 167.150 137.955 168.055 ;
        RECT 136.725 166.575 137.080 166.945 ;
        RECT 137.360 166.915 137.530 167.125 ;
        RECT 137.360 166.585 137.615 166.915 ;
        RECT 137.360 166.395 137.530 166.585 ;
        RECT 137.785 166.420 137.955 167.150 ;
        RECT 138.130 167.075 138.390 168.225 ;
        RECT 138.565 167.135 139.775 168.225 ;
        RECT 138.565 166.595 139.085 167.135 ;
        RECT 136.815 166.225 137.530 166.395 ;
        RECT 136.815 165.845 136.985 166.225 ;
        RECT 137.200 165.675 137.530 166.055 ;
        RECT 137.700 165.845 137.955 166.420 ;
        RECT 138.130 165.675 138.390 166.515 ;
        RECT 139.255 166.425 139.775 166.965 ;
        RECT 138.565 165.675 139.775 166.425 ;
        RECT 27.160 165.505 139.860 165.675 ;
      LAYER met1 ;
        RECT 82.890 210.370 83.210 210.430 ;
        RECT 118.310 210.370 118.630 210.430 ;
        RECT 82.890 210.230 118.630 210.370 ;
        RECT 82.890 210.170 83.210 210.230 ;
        RECT 118.310 210.170 118.630 210.230 ;
        RECT 89.790 210.030 90.110 210.090 ;
        RECT 129.350 210.030 129.670 210.090 ;
        RECT 89.790 209.890 129.670 210.030 ;
        RECT 89.790 209.830 90.110 209.890 ;
        RECT 129.350 209.830 129.670 209.890 ;
        RECT 64.950 209.690 65.270 209.750 ;
        RECT 95.770 209.690 96.090 209.750 ;
        RECT 64.950 209.550 96.090 209.690 ;
        RECT 64.950 209.490 65.270 209.550 ;
        RECT 95.770 209.490 96.090 209.550 ;
        RECT 125.670 209.690 125.990 209.750 ;
        RECT 129.810 209.690 130.130 209.750 ;
        RECT 125.670 209.550 130.130 209.690 ;
        RECT 125.670 209.490 125.990 209.550 ;
        RECT 129.810 209.490 130.130 209.550 ;
        RECT 27.160 208.870 139.860 209.350 ;
        RECT 75.070 208.670 75.390 208.730 ;
        RECT 75.545 208.670 75.835 208.715 ;
        RECT 75.070 208.530 75.835 208.670 ;
        RECT 75.070 208.470 75.390 208.530 ;
        RECT 75.545 208.485 75.835 208.530 ;
        RECT 87.030 208.470 87.350 208.730 ;
        RECT 89.330 208.470 89.650 208.730 ;
        RECT 90.250 208.470 90.570 208.730 ;
        RECT 93.485 208.670 93.775 208.715 ;
        RECT 100.830 208.670 101.150 208.730 ;
        RECT 93.485 208.530 101.150 208.670 ;
        RECT 93.485 208.485 93.775 208.530 ;
        RECT 100.830 208.470 101.150 208.530 ;
        RECT 104.510 208.670 104.830 208.730 ;
        RECT 109.125 208.670 109.415 208.715 ;
        RECT 104.510 208.530 109.415 208.670 ;
        RECT 104.510 208.470 104.830 208.530 ;
        RECT 109.125 208.485 109.415 208.530 ;
        RECT 111.870 208.670 112.190 208.730 ;
        RECT 112.805 208.670 113.095 208.715 ;
        RECT 111.870 208.530 113.095 208.670 ;
        RECT 111.870 208.470 112.190 208.530 ;
        RECT 112.805 208.485 113.095 208.530 ;
        RECT 115.090 208.670 115.410 208.730 ;
        RECT 116.025 208.670 116.315 208.715 ;
        RECT 115.090 208.530 116.315 208.670 ;
        RECT 115.090 208.470 115.410 208.530 ;
        RECT 116.025 208.485 116.315 208.530 ;
        RECT 118.770 208.670 119.090 208.730 ;
        RECT 119.245 208.670 119.535 208.715 ;
        RECT 118.770 208.530 119.535 208.670 ;
        RECT 118.770 208.470 119.090 208.530 ;
        RECT 119.245 208.485 119.535 208.530 ;
        RECT 126.605 208.670 126.895 208.715 ;
        RECT 127.510 208.670 127.830 208.730 ;
        RECT 126.605 208.530 127.830 208.670 ;
        RECT 126.605 208.485 126.895 208.530 ;
        RECT 127.510 208.470 127.830 208.530 ;
        RECT 127.970 208.470 128.290 208.730 ;
        RECT 128.430 208.670 128.750 208.730 ;
        RECT 136.725 208.670 137.015 208.715 ;
        RECT 128.430 208.530 137.015 208.670 ;
        RECT 128.430 208.470 128.750 208.530 ;
        RECT 136.725 208.485 137.015 208.530 ;
        RECT 86.110 208.330 86.430 208.390 ;
        RECT 83.670 208.190 86.430 208.330 ;
        RECT 30.005 207.990 30.295 208.035 ;
        RECT 35.510 207.990 35.830 208.050 ;
        RECT 30.005 207.850 35.830 207.990 ;
        RECT 30.005 207.805 30.295 207.850 ;
        RECT 35.510 207.790 35.830 207.850 ;
        RECT 56.670 207.790 56.990 208.050 ;
        RECT 66.790 207.990 67.110 208.050 ;
        RECT 67.265 207.990 67.555 208.035 ;
        RECT 66.790 207.850 67.555 207.990 ;
        RECT 66.790 207.790 67.110 207.850 ;
        RECT 67.265 207.805 67.555 207.850 ;
        RECT 75.530 207.790 75.850 208.050 ;
        RECT 81.525 207.990 81.815 208.035 ;
        RECT 83.670 207.990 83.810 208.190 ;
        RECT 86.110 208.130 86.430 208.190 ;
        RECT 81.525 207.850 83.810 207.990 ;
        RECT 81.525 207.805 81.815 207.850 ;
        RECT 84.745 207.805 85.035 208.035 ;
        RECT 85.205 207.990 85.495 208.035 ;
        RECT 87.120 207.990 87.260 208.470 ;
        RECT 95.770 208.130 96.090 208.390 ;
        RECT 96.705 208.330 96.995 208.375 ;
        RECT 97.610 208.330 97.930 208.390 ;
        RECT 96.705 208.190 97.930 208.330 ;
        RECT 100.920 208.330 101.060 208.470 ;
        RECT 108.205 208.330 108.495 208.375 ;
        RECT 108.650 208.330 108.970 208.390 ;
        RECT 134.410 208.330 134.730 208.390 ;
        RECT 100.920 208.190 107.960 208.330 ;
        RECT 96.705 208.145 96.995 208.190 ;
        RECT 97.610 208.130 97.930 208.190 ;
        RECT 85.205 207.850 87.260 207.990 ;
        RECT 85.205 207.805 85.495 207.850 ;
        RECT 27.230 207.650 27.550 207.710 ;
        RECT 30.465 207.650 30.755 207.695 ;
        RECT 27.230 207.510 30.755 207.650 ;
        RECT 27.230 207.450 27.550 207.510 ;
        RECT 30.465 207.465 30.755 207.510 ;
        RECT 57.130 207.450 57.450 207.710 ;
        RECT 57.590 207.450 57.910 207.710 ;
        RECT 77.370 207.650 77.690 207.710 ;
        RECT 77.845 207.650 78.135 207.695 ;
        RECT 77.370 207.510 78.135 207.650 ;
        RECT 77.370 207.450 77.690 207.510 ;
        RECT 77.845 207.465 78.135 207.510 ;
        RECT 83.365 207.650 83.655 207.695 ;
        RECT 84.820 207.650 84.960 207.805 ;
        RECT 88.410 207.790 88.730 208.050 ;
        RECT 91.185 207.990 91.475 208.035 ;
        RECT 92.090 207.990 92.410 208.050 ;
        RECT 91.185 207.850 92.410 207.990 ;
        RECT 91.185 207.805 91.475 207.850 ;
        RECT 92.090 207.790 92.410 207.850 ;
        RECT 92.565 207.990 92.855 208.035 ;
        RECT 95.310 207.990 95.630 208.050 ;
        RECT 97.165 207.990 97.455 208.035 ;
        RECT 92.565 207.850 95.630 207.990 ;
        RECT 92.565 207.805 92.855 207.850 ;
        RECT 95.310 207.790 95.630 207.850 ;
        RECT 95.860 207.850 97.455 207.990 ;
        RECT 94.850 207.650 95.170 207.710 ;
        RECT 83.365 207.510 95.170 207.650 ;
        RECT 83.365 207.465 83.655 207.510 ;
        RECT 94.850 207.450 95.170 207.510 ;
        RECT 79.670 207.310 79.990 207.370 ;
        RECT 82.445 207.310 82.735 207.355 ;
        RECT 95.860 207.310 96.000 207.850 ;
        RECT 97.165 207.805 97.455 207.850 ;
        RECT 98.990 207.990 99.310 208.050 ;
        RECT 99.465 207.990 99.755 208.035 ;
        RECT 98.990 207.850 99.755 207.990 ;
        RECT 98.990 207.790 99.310 207.850 ;
        RECT 99.465 207.805 99.755 207.850 ;
        RECT 100.370 207.990 100.690 208.050 ;
        RECT 106.350 207.990 106.670 208.050 ;
        RECT 107.820 208.035 107.960 208.190 ;
        RECT 108.205 208.190 115.320 208.330 ;
        RECT 108.205 208.145 108.495 208.190 ;
        RECT 108.650 208.130 108.970 208.190 ;
        RECT 100.370 207.850 106.670 207.990 ;
        RECT 100.370 207.790 100.690 207.850 ;
        RECT 106.350 207.790 106.670 207.850 ;
        RECT 107.285 207.805 107.575 208.035 ;
        RECT 107.745 207.805 108.035 208.035 ;
        RECT 100.845 207.650 101.135 207.695 ;
        RECT 104.510 207.650 104.830 207.710 ;
        RECT 107.360 207.650 107.500 207.805 ;
        RECT 110.030 207.790 110.350 208.050 ;
        RECT 111.500 208.035 111.640 208.190 ;
        RECT 111.425 207.805 111.715 208.035 ;
        RECT 113.725 207.805 114.015 208.035 ;
        RECT 113.800 207.650 113.940 207.805 ;
        RECT 114.170 207.790 114.490 208.050 ;
        RECT 115.180 208.035 115.320 208.190 ;
        RECT 117.020 208.190 134.730 208.330 ;
        RECT 117.020 208.035 117.160 208.190 ;
        RECT 134.410 208.130 134.730 208.190 ;
        RECT 115.105 207.805 115.395 208.035 ;
        RECT 116.945 207.805 117.235 208.035 ;
        RECT 120.165 207.990 120.455 208.035 ;
        RECT 120.165 207.850 121.300 207.990 ;
        RECT 120.165 207.805 120.455 207.850 ;
        RECT 121.160 207.650 121.300 207.850 ;
        RECT 121.530 207.790 121.850 208.050 ;
        RECT 125.670 207.790 125.990 208.050 ;
        RECT 127.050 207.790 127.370 208.050 ;
        RECT 127.970 207.990 128.290 208.050 ;
        RECT 128.445 207.990 128.735 208.035 ;
        RECT 127.970 207.850 128.735 207.990 ;
        RECT 127.970 207.790 128.290 207.850 ;
        RECT 128.445 207.805 128.735 207.850 ;
        RECT 131.190 207.790 131.510 208.050 ;
        RECT 137.630 207.790 137.950 208.050 ;
        RECT 124.750 207.650 125.070 207.710 ;
        RECT 133.045 207.650 133.335 207.695 ;
        RECT 100.845 207.510 107.040 207.650 ;
        RECT 107.360 207.510 110.720 207.650 ;
        RECT 113.800 207.510 120.840 207.650 ;
        RECT 121.160 207.510 124.520 207.650 ;
        RECT 100.845 207.465 101.135 207.510 ;
        RECT 104.510 207.450 104.830 207.510 ;
        RECT 79.670 207.170 96.000 207.310 ;
        RECT 96.230 207.310 96.550 207.370 ;
        RECT 98.070 207.310 98.390 207.370 ;
        RECT 104.050 207.310 104.370 207.370 ;
        RECT 96.230 207.170 104.370 207.310 ;
        RECT 79.670 207.110 79.990 207.170 ;
        RECT 82.445 207.125 82.735 207.170 ;
        RECT 96.230 207.110 96.550 207.170 ;
        RECT 98.070 207.110 98.390 207.170 ;
        RECT 104.050 207.110 104.370 207.170 ;
        RECT 105.430 207.310 105.750 207.370 ;
        RECT 106.365 207.310 106.655 207.355 ;
        RECT 105.430 207.170 106.655 207.310 ;
        RECT 106.900 207.310 107.040 207.510 ;
        RECT 108.190 207.310 108.510 207.370 ;
        RECT 110.580 207.355 110.720 207.510 ;
        RECT 120.700 207.355 120.840 207.510 ;
        RECT 106.900 207.170 108.510 207.310 ;
        RECT 105.430 207.110 105.750 207.170 ;
        RECT 106.365 207.125 106.655 207.170 ;
        RECT 108.190 207.110 108.510 207.170 ;
        RECT 110.505 207.125 110.795 207.355 ;
        RECT 111.040 207.170 118.310 207.310 ;
        RECT 25.390 206.970 25.710 207.030 ;
        RECT 29.085 206.970 29.375 207.015 ;
        RECT 25.390 206.830 29.375 206.970 ;
        RECT 25.390 206.770 25.710 206.830 ;
        RECT 29.085 206.785 29.375 206.830 ;
        RECT 52.990 206.970 53.310 207.030 ;
        RECT 54.845 206.970 55.135 207.015 ;
        RECT 52.990 206.830 55.135 206.970 ;
        RECT 52.990 206.770 53.310 206.830 ;
        RECT 54.845 206.785 55.135 206.830 ;
        RECT 68.170 206.770 68.490 207.030 ;
        RECT 72.310 206.970 72.630 207.030 ;
        RECT 74.625 206.970 74.915 207.015 ;
        RECT 72.310 206.830 74.915 206.970 ;
        RECT 72.310 206.770 72.630 206.830 ;
        RECT 74.625 206.785 74.915 206.830 ;
        RECT 77.385 206.970 77.675 207.015 ;
        RECT 80.130 206.970 80.450 207.030 ;
        RECT 77.385 206.830 80.450 206.970 ;
        RECT 77.385 206.785 77.675 206.830 ;
        RECT 80.130 206.770 80.450 206.830 ;
        RECT 83.825 206.970 84.115 207.015 ;
        RECT 84.270 206.970 84.590 207.030 ;
        RECT 83.825 206.830 84.590 206.970 ;
        RECT 83.825 206.785 84.115 206.830 ;
        RECT 84.270 206.770 84.590 206.830 ;
        RECT 86.125 206.970 86.415 207.015 ;
        RECT 90.250 206.970 90.570 207.030 ;
        RECT 86.125 206.830 90.570 206.970 ;
        RECT 86.125 206.785 86.415 206.830 ;
        RECT 90.250 206.770 90.570 206.830 ;
        RECT 94.865 206.970 95.155 207.015 ;
        RECT 95.310 206.970 95.630 207.030 ;
        RECT 94.865 206.830 95.630 206.970 ;
        RECT 94.865 206.785 95.155 206.830 ;
        RECT 95.310 206.770 95.630 206.830 ;
        RECT 103.130 206.970 103.450 207.030 ;
        RECT 105.890 206.970 106.210 207.030 ;
        RECT 111.040 206.970 111.180 207.170 ;
        RECT 103.130 206.830 111.180 206.970 ;
        RECT 112.330 206.970 112.650 207.030 ;
        RECT 115.105 206.970 115.395 207.015 ;
        RECT 112.330 206.830 115.395 206.970 ;
        RECT 118.170 206.970 118.310 207.170 ;
        RECT 120.625 207.125 120.915 207.355 ;
        RECT 124.380 207.310 124.520 207.510 ;
        RECT 124.750 207.510 133.335 207.650 ;
        RECT 124.750 207.450 125.070 207.510 ;
        RECT 133.045 207.465 133.335 207.510 ;
        RECT 135.790 207.310 136.110 207.370 ;
        RECT 124.380 207.170 136.110 207.310 ;
        RECT 135.790 207.110 136.110 207.170 ;
        RECT 121.530 206.970 121.850 207.030 ;
        RECT 118.170 206.830 121.850 206.970 ;
        RECT 103.130 206.770 103.450 206.830 ;
        RECT 105.890 206.770 106.210 206.830 ;
        RECT 112.330 206.770 112.650 206.830 ;
        RECT 115.105 206.785 115.395 206.830 ;
        RECT 121.530 206.770 121.850 206.830 ;
        RECT 122.910 206.970 123.230 207.030 ;
        RECT 129.365 206.970 129.655 207.015 ;
        RECT 122.910 206.830 129.655 206.970 ;
        RECT 122.910 206.770 123.230 206.830 ;
        RECT 129.365 206.785 129.655 206.830 ;
        RECT 27.160 206.150 139.860 206.630 ;
        RECT 35.510 205.750 35.830 206.010 ;
        RECT 52.070 205.950 52.390 206.010 ;
        RECT 43.420 205.810 52.390 205.950 ;
        RECT 39.205 205.610 39.495 205.655 ;
        RECT 40.585 205.610 40.875 205.655 ;
        RECT 39.205 205.470 40.875 205.610 ;
        RECT 39.205 205.425 39.495 205.470 ;
        RECT 40.585 205.425 40.875 205.470 ;
        RECT 29.990 204.730 30.310 204.990 ;
        RECT 36.430 204.730 36.750 204.990 ;
        RECT 37.810 204.730 38.130 204.990 ;
        RECT 38.270 204.730 38.590 204.990 ;
        RECT 39.650 204.930 39.970 204.990 ;
        RECT 43.420 204.930 43.560 205.810 ;
        RECT 52.070 205.750 52.390 205.810 ;
        RECT 53.910 205.950 54.230 206.010 ;
        RECT 57.590 205.950 57.910 206.010 ;
        RECT 53.910 205.810 57.910 205.950 ;
        RECT 53.910 205.750 54.230 205.810 ;
        RECT 57.590 205.750 57.910 205.810 ;
        RECT 74.165 205.950 74.455 205.995 ;
        RECT 77.370 205.950 77.690 206.010 ;
        RECT 74.165 205.810 77.690 205.950 ;
        RECT 74.165 205.765 74.455 205.810 ;
        RECT 77.370 205.750 77.690 205.810 ;
        RECT 80.130 205.750 80.450 206.010 ;
        RECT 88.870 205.950 89.190 206.010 ;
        RECT 89.345 205.950 89.635 205.995 ;
        RECT 88.870 205.810 89.635 205.950 ;
        RECT 88.870 205.750 89.190 205.810 ;
        RECT 89.345 205.765 89.635 205.810 ;
        RECT 92.090 205.750 92.410 206.010 ;
        RECT 93.930 205.950 94.250 206.010 ;
        RECT 98.530 205.950 98.850 206.010 ;
        RECT 93.930 205.810 98.850 205.950 ;
        RECT 93.930 205.750 94.250 205.810 ;
        RECT 98.530 205.750 98.850 205.810 ;
        RECT 99.910 205.950 100.230 206.010 ;
        RECT 100.845 205.950 101.135 205.995 ;
        RECT 99.910 205.810 101.135 205.950 ;
        RECT 99.910 205.750 100.230 205.810 ;
        RECT 100.845 205.765 101.135 205.810 ;
        RECT 101.765 205.950 102.055 205.995 ;
        RECT 110.030 205.950 110.350 206.010 ;
        RECT 101.765 205.810 110.350 205.950 ;
        RECT 101.765 205.765 102.055 205.810 ;
        RECT 110.030 205.750 110.350 205.810 ;
        RECT 110.490 205.750 110.810 206.010 ;
        RECT 113.250 205.950 113.570 206.010 ;
        RECT 116.485 205.950 116.775 205.995 ;
        RECT 113.250 205.810 116.775 205.950 ;
        RECT 113.250 205.750 113.570 205.810 ;
        RECT 116.485 205.765 116.775 205.810 ;
        RECT 123.845 205.950 124.135 205.995 ;
        RECT 131.190 205.950 131.510 206.010 ;
        RECT 123.845 205.810 131.510 205.950 ;
        RECT 123.845 205.765 124.135 205.810 ;
        RECT 131.190 205.750 131.510 205.810 ;
        RECT 134.410 205.750 134.730 206.010 ;
        RECT 135.790 205.750 136.110 206.010 ;
        RECT 50.245 205.610 50.535 205.655 ;
        RECT 50.245 205.470 57.360 205.610 ;
        RECT 50.245 205.425 50.535 205.470 ;
        RECT 43.805 205.270 44.095 205.315 ;
        RECT 51.150 205.270 51.470 205.330 ;
        RECT 43.805 205.130 51.470 205.270 ;
        RECT 43.805 205.085 44.095 205.130 ;
        RECT 51.150 205.070 51.470 205.130 ;
        RECT 52.530 205.270 52.850 205.330 ;
        RECT 52.530 205.130 53.680 205.270 ;
        RECT 52.530 205.070 52.850 205.130 ;
        RECT 39.650 204.790 43.560 204.930 ;
        RECT 51.625 204.930 51.915 204.975 ;
        RECT 52.085 204.930 52.375 204.975 ;
        RECT 51.625 204.790 52.375 204.930 ;
        RECT 39.650 204.730 39.970 204.790 ;
        RECT 51.625 204.745 51.915 204.790 ;
        RECT 52.085 204.745 52.375 204.790 ;
        RECT 52.990 204.730 53.310 204.990 ;
        RECT 53.540 204.975 53.680 205.130 ;
        RECT 54.370 205.070 54.690 205.330 ;
        RECT 53.465 204.745 53.755 204.975 ;
        RECT 54.845 204.745 55.135 204.975 ;
        RECT 57.220 204.930 57.360 205.470 ;
        RECT 57.680 205.270 57.820 205.750 ;
        RECT 64.030 205.410 64.350 205.670 ;
        RECT 87.490 205.610 87.810 205.670 ;
        RECT 77.460 205.470 87.810 205.610 ;
        RECT 58.065 205.270 58.355 205.315 ;
        RECT 57.680 205.130 58.355 205.270 ;
        RECT 58.065 205.085 58.355 205.130 ;
        RECT 64.045 204.930 64.335 204.975 ;
        RECT 57.220 204.790 64.335 204.930 ;
        RECT 64.045 204.745 64.335 204.790 ;
        RECT 36.905 204.590 37.195 204.635 ;
        RECT 47.930 204.590 48.250 204.650 ;
        RECT 36.905 204.450 48.250 204.590 ;
        RECT 36.905 204.405 37.195 204.450 ;
        RECT 47.930 204.390 48.250 204.450 ;
        RECT 50.230 204.390 50.550 204.650 ;
        RECT 50.690 204.590 51.010 204.650 ;
        RECT 54.920 204.590 55.060 204.745 ;
        RECT 64.950 204.730 65.270 204.990 ;
        RECT 65.410 204.730 65.730 204.990 ;
        RECT 66.790 204.730 67.110 204.990 ;
        RECT 68.185 204.745 68.475 204.975 ;
        RECT 75.530 204.930 75.820 204.975 ;
        RECT 77.460 204.930 77.600 205.470 ;
        RECT 87.490 205.410 87.810 205.470 ;
        RECT 88.410 205.610 88.730 205.670 ;
        RECT 111.425 205.610 111.715 205.655 ;
        RECT 88.410 205.470 111.715 205.610 ;
        RECT 88.410 205.410 88.730 205.470 ;
        RECT 111.425 205.425 111.715 205.470 ;
        RECT 115.105 205.610 115.395 205.655 ;
        RECT 137.630 205.610 137.950 205.670 ;
        RECT 115.105 205.470 137.950 205.610 ;
        RECT 115.105 205.425 115.395 205.470 ;
        RECT 137.630 205.410 137.950 205.470 ;
        RECT 81.510 205.270 81.830 205.330 ;
        RECT 82.905 205.270 83.195 205.315 ;
        RECT 81.510 205.130 83.195 205.270 ;
        RECT 81.510 205.070 81.830 205.130 ;
        RECT 82.905 205.085 83.195 205.130 ;
        RECT 83.810 205.270 84.130 205.330 ;
        RECT 92.550 205.270 92.870 205.330 ;
        RECT 103.130 205.270 103.450 205.330 ;
        RECT 83.810 205.130 90.940 205.270 ;
        RECT 83.810 205.070 84.130 205.130 ;
        RECT 75.530 204.790 77.600 204.930 ;
        RECT 75.530 204.745 75.820 204.790 ;
        RECT 50.690 204.450 55.060 204.590 ;
        RECT 57.145 204.590 57.435 204.635 ;
        RECT 63.570 204.590 63.890 204.650 ;
        RECT 57.145 204.450 63.890 204.590 ;
        RECT 50.690 204.390 51.010 204.450 ;
        RECT 57.145 204.405 57.435 204.450 ;
        RECT 63.570 204.390 63.890 204.450 ;
        RECT 65.870 204.590 66.190 204.650 ;
        RECT 68.260 204.590 68.400 204.745 ;
        RECT 77.830 204.730 78.150 204.990 ;
        RECT 84.745 204.930 85.035 204.975 ;
        RECT 85.190 204.930 85.510 204.990 ;
        RECT 78.380 204.790 83.810 204.930 ;
        RECT 65.870 204.450 68.400 204.590 ;
        RECT 71.390 204.590 71.710 204.650 ;
        RECT 72.325 204.590 72.615 204.635 ;
        RECT 71.390 204.450 72.615 204.590 ;
        RECT 65.870 204.390 66.190 204.450 ;
        RECT 71.390 204.390 71.710 204.450 ;
        RECT 72.325 204.405 72.615 204.450 ;
        RECT 73.245 204.590 73.535 204.635 ;
        RECT 75.070 204.590 75.390 204.650 ;
        RECT 73.245 204.450 75.760 204.590 ;
        RECT 73.245 204.405 73.535 204.450 ;
        RECT 75.070 204.390 75.390 204.450 ;
        RECT 25.390 204.250 25.710 204.310 ;
        RECT 29.085 204.250 29.375 204.295 ;
        RECT 25.390 204.110 29.375 204.250 ;
        RECT 25.390 204.050 25.710 204.110 ;
        RECT 29.085 204.065 29.375 204.110 ;
        RECT 41.490 204.250 41.810 204.310 ;
        RECT 42.425 204.250 42.715 204.295 ;
        RECT 41.490 204.110 42.715 204.250 ;
        RECT 41.490 204.050 41.810 204.110 ;
        RECT 42.425 204.065 42.715 204.110 ;
        RECT 42.870 204.050 43.190 204.310 ;
        RECT 49.310 204.250 49.630 204.310 ;
        RECT 51.165 204.250 51.455 204.295 ;
        RECT 49.310 204.110 51.455 204.250 ;
        RECT 49.310 204.050 49.630 204.110 ;
        RECT 51.165 204.065 51.455 204.110 ;
        RECT 51.610 204.250 51.930 204.310 ;
        RECT 55.305 204.250 55.595 204.295 ;
        RECT 51.610 204.110 55.595 204.250 ;
        RECT 51.610 204.050 51.930 204.110 ;
        RECT 55.305 204.065 55.595 204.110 ;
        RECT 57.605 204.250 57.895 204.295 ;
        RECT 58.050 204.250 58.370 204.310 ;
        RECT 57.605 204.110 58.370 204.250 ;
        RECT 57.605 204.065 57.895 204.110 ;
        RECT 58.050 204.050 58.370 204.110 ;
        RECT 67.250 204.050 67.570 204.310 ;
        RECT 69.105 204.250 69.395 204.295 ;
        RECT 69.550 204.250 69.870 204.310 ;
        RECT 69.105 204.110 69.870 204.250 ;
        RECT 69.105 204.065 69.395 204.110 ;
        RECT 69.550 204.050 69.870 204.110 ;
        RECT 74.610 204.050 74.930 204.310 ;
        RECT 75.620 204.295 75.760 204.450 ;
        RECT 75.545 204.250 75.835 204.295 ;
        RECT 78.380 204.250 78.520 204.790 ;
        RECT 80.590 204.590 80.910 204.650 ;
        RECT 82.445 204.590 82.735 204.635 ;
        RECT 80.590 204.450 82.735 204.590 ;
        RECT 83.670 204.590 83.810 204.790 ;
        RECT 84.745 204.790 85.510 204.930 ;
        RECT 84.745 204.745 85.035 204.790 ;
        RECT 85.190 204.730 85.510 204.790 ;
        RECT 85.650 204.730 85.970 204.990 ;
        RECT 86.585 204.930 86.875 204.975 ;
        RECT 87.950 204.930 88.270 204.990 ;
        RECT 86.585 204.790 88.270 204.930 ;
        RECT 86.585 204.745 86.875 204.790 ;
        RECT 87.950 204.730 88.270 204.790 ;
        RECT 88.870 204.930 89.190 204.990 ;
        RECT 90.265 204.930 90.555 204.975 ;
        RECT 88.870 204.790 90.555 204.930 ;
        RECT 90.800 204.930 90.940 205.130 ;
        RECT 92.550 205.130 99.220 205.270 ;
        RECT 92.550 205.070 92.870 205.130 ;
        RECT 93.025 204.930 93.315 204.975 ;
        RECT 90.800 204.790 93.315 204.930 ;
        RECT 88.870 204.730 89.190 204.790 ;
        RECT 90.265 204.745 90.555 204.790 ;
        RECT 93.025 204.745 93.315 204.790 ;
        RECT 93.930 204.730 94.250 204.990 ;
        RECT 94.405 204.930 94.695 204.975 ;
        RECT 94.850 204.930 95.170 204.990 ;
        RECT 94.405 204.790 95.170 204.930 ;
        RECT 94.405 204.745 94.695 204.790 ;
        RECT 94.850 204.730 95.170 204.790 ;
        RECT 95.325 204.930 95.615 204.975 ;
        RECT 95.325 204.790 96.920 204.930 ;
        RECT 95.325 204.745 95.615 204.790 ;
        RECT 88.410 204.590 88.730 204.650 ;
        RECT 83.670 204.450 88.730 204.590 ;
        RECT 80.590 204.390 80.910 204.450 ;
        RECT 82.445 204.405 82.735 204.450 ;
        RECT 88.410 204.390 88.730 204.450 ;
        RECT 75.545 204.110 78.520 204.250 ;
        RECT 81.985 204.250 82.275 204.295 ;
        RECT 83.350 204.250 83.670 204.310 ;
        RECT 81.985 204.110 83.670 204.250 ;
        RECT 75.545 204.065 75.835 204.110 ;
        RECT 81.985 204.065 82.275 204.110 ;
        RECT 83.350 204.050 83.670 204.110 ;
        RECT 84.730 204.050 85.050 204.310 ;
        RECT 86.570 204.250 86.890 204.310 ;
        RECT 87.045 204.250 87.335 204.295 ;
        RECT 86.570 204.110 87.335 204.250 ;
        RECT 86.570 204.050 86.890 204.110 ;
        RECT 87.045 204.065 87.335 204.110 ;
        RECT 91.185 204.250 91.475 204.295 ;
        RECT 92.550 204.250 92.870 204.310 ;
        RECT 91.185 204.110 92.870 204.250 ;
        RECT 91.185 204.065 91.475 204.110 ;
        RECT 92.550 204.050 92.870 204.110 ;
        RECT 93.930 204.250 94.250 204.310 ;
        RECT 95.400 204.250 95.540 204.745 ;
        RECT 96.230 204.390 96.550 204.650 ;
        RECT 96.780 204.310 96.920 204.790 ;
        RECT 97.610 204.730 97.930 204.990 ;
        RECT 98.070 204.730 98.390 204.990 ;
        RECT 99.080 204.930 99.220 205.130 ;
        RECT 103.130 205.130 105.200 205.270 ;
        RECT 103.130 205.070 103.450 205.130 ;
        RECT 102.685 204.930 102.975 204.975 ;
        RECT 99.080 204.790 102.975 204.930 ;
        RECT 102.685 204.745 102.975 204.790 ;
        RECT 104.050 204.730 104.370 204.990 ;
        RECT 105.060 204.975 105.200 205.130 ;
        RECT 105.890 205.070 106.210 205.330 ;
        RECT 107.285 205.270 107.575 205.315 ;
        RECT 107.730 205.270 108.050 205.330 ;
        RECT 111.870 205.270 112.190 205.330 ;
        RECT 107.285 205.130 108.050 205.270 ;
        RECT 107.285 205.085 107.575 205.130 ;
        RECT 107.730 205.070 108.050 205.130 ;
        RECT 108.280 205.130 112.190 205.270 ;
        RECT 108.280 204.990 108.420 205.130 ;
        RECT 111.870 205.070 112.190 205.130 ;
        RECT 114.630 205.270 114.950 205.330 ;
        RECT 126.590 205.270 126.910 205.330 ;
        RECT 114.630 205.130 118.540 205.270 ;
        RECT 114.630 205.070 114.950 205.130 ;
        RECT 104.955 204.745 105.245 204.975 ;
        RECT 105.430 204.730 105.750 204.990 ;
        RECT 106.350 204.930 106.670 204.990 ;
        RECT 106.350 204.790 107.960 204.930 ;
        RECT 106.350 204.730 106.670 204.790 ;
        RECT 93.930 204.110 95.540 204.250 ;
        RECT 93.930 204.050 94.250 204.110 ;
        RECT 96.690 204.050 97.010 204.310 ;
        RECT 97.700 204.250 97.840 204.730 ;
        RECT 99.005 204.590 99.295 204.635 ;
        RECT 100.370 204.590 100.690 204.650 ;
        RECT 99.005 204.450 100.690 204.590 ;
        RECT 99.005 204.405 99.295 204.450 ;
        RECT 100.370 204.390 100.690 204.450 ;
        RECT 101.075 204.590 101.365 204.635 ;
        RECT 102.210 204.590 102.530 204.650 ;
        RECT 101.075 204.450 102.530 204.590 ;
        RECT 101.075 204.405 101.365 204.450 ;
        RECT 102.210 204.390 102.530 204.450 ;
        RECT 104.525 204.590 104.815 204.635 ;
        RECT 104.525 204.450 105.200 204.590 ;
        RECT 104.525 204.405 104.815 204.450 ;
        RECT 105.060 204.420 105.200 204.450 ;
        RECT 105.890 204.420 106.210 204.650 ;
        RECT 107.820 204.590 107.960 204.790 ;
        RECT 108.190 204.730 108.510 204.990 ;
        RECT 108.650 204.730 108.970 204.990 ;
        RECT 110.030 204.930 110.350 204.990 ;
        RECT 112.345 204.930 112.635 204.975 ;
        RECT 110.030 204.790 112.635 204.930 ;
        RECT 110.030 204.730 110.350 204.790 ;
        RECT 112.345 204.745 112.635 204.790 ;
        RECT 112.790 204.730 113.110 204.990 ;
        RECT 113.725 204.930 114.015 204.975 ;
        RECT 113.340 204.790 114.015 204.930 ;
        RECT 109.585 204.590 109.875 204.635 ;
        RECT 107.820 204.450 109.875 204.590 ;
        RECT 105.060 204.390 106.210 204.420 ;
        RECT 109.585 204.405 109.875 204.450 ;
        RECT 110.950 204.590 111.270 204.650 ;
        RECT 113.340 204.590 113.480 204.790 ;
        RECT 113.725 204.745 114.015 204.790 ;
        RECT 114.170 204.730 114.490 204.990 ;
        RECT 116.010 204.730 116.330 204.990 ;
        RECT 116.945 204.930 117.235 204.975 ;
        RECT 117.390 204.930 117.710 204.990 ;
        RECT 116.945 204.790 117.710 204.930 ;
        RECT 116.945 204.745 117.235 204.790 ;
        RECT 117.390 204.730 117.710 204.790 ;
        RECT 117.850 204.730 118.170 204.990 ;
        RECT 118.400 204.975 118.540 205.130 ;
        RECT 122.080 205.130 126.910 205.270 ;
        RECT 118.330 204.745 118.620 204.975 ;
        RECT 120.610 204.730 120.930 204.990 ;
        RECT 121.530 204.975 121.850 204.990 ;
        RECT 122.080 204.975 122.220 205.130 ;
        RECT 126.590 205.070 126.910 205.130 ;
        RECT 133.030 205.270 133.350 205.330 ;
        RECT 133.030 205.130 136.940 205.270 ;
        RECT 133.030 205.070 133.350 205.130 ;
        RECT 122.910 204.975 123.230 204.990 ;
        RECT 121.365 204.745 121.850 204.975 ;
        RECT 122.005 204.745 122.295 204.975 ;
        RECT 122.910 204.745 123.240 204.975 ;
        RECT 131.190 204.930 131.510 204.990 ;
        RECT 124.840 204.790 131.510 204.930 ;
        RECT 121.530 204.730 121.850 204.745 ;
        RECT 122.910 204.730 123.230 204.745 ;
        RECT 110.950 204.450 113.480 204.590 ;
        RECT 116.470 204.590 116.790 204.650 ;
        RECT 122.465 204.590 122.755 204.635 ;
        RECT 124.840 204.590 124.980 204.790 ;
        RECT 131.190 204.730 131.510 204.790 ;
        RECT 135.330 204.730 135.650 204.990 ;
        RECT 136.800 204.975 136.940 205.130 ;
        RECT 136.725 204.745 137.015 204.975 ;
        RECT 116.470 204.450 121.580 204.590 ;
        RECT 110.950 204.390 111.270 204.450 ;
        RECT 116.470 204.390 116.790 204.450 ;
        RECT 103.590 204.250 103.910 204.310 ;
        RECT 105.060 204.280 106.120 204.390 ;
        RECT 97.700 204.110 103.910 204.250 ;
        RECT 103.590 204.050 103.910 204.110 ;
        RECT 109.110 204.250 109.430 204.310 ;
        RECT 110.505 204.250 110.795 204.295 ;
        RECT 109.110 204.110 110.795 204.250 ;
        RECT 109.110 204.050 109.430 204.110 ;
        RECT 110.505 204.065 110.795 204.110 ;
        RECT 113.710 204.250 114.030 204.310 ;
        RECT 116.010 204.250 116.330 204.310 ;
        RECT 118.770 204.250 119.090 204.310 ;
        RECT 113.710 204.110 119.090 204.250 ;
        RECT 113.710 204.050 114.030 204.110 ;
        RECT 116.010 204.050 116.330 204.110 ;
        RECT 118.770 204.050 119.090 204.110 ;
        RECT 119.230 204.250 119.550 204.310 ;
        RECT 119.705 204.250 119.995 204.295 ;
        RECT 119.230 204.110 119.995 204.250 ;
        RECT 121.440 204.250 121.580 204.450 ;
        RECT 122.465 204.450 124.980 204.590 ;
        RECT 122.465 204.405 122.755 204.450 ;
        RECT 125.210 204.390 125.530 204.650 ;
        RECT 137.185 204.590 137.475 204.635 ;
        RECT 125.760 204.450 137.475 204.590 ;
        RECT 122.910 204.250 123.230 204.310 ;
        RECT 121.440 204.110 123.230 204.250 ;
        RECT 119.230 204.050 119.550 204.110 ;
        RECT 119.705 204.065 119.995 204.110 ;
        RECT 122.910 204.050 123.230 204.110 ;
        RECT 124.750 204.250 125.070 204.310 ;
        RECT 125.760 204.250 125.900 204.450 ;
        RECT 137.185 204.405 137.475 204.450 ;
        RECT 124.750 204.110 125.900 204.250 ;
        RECT 124.750 204.050 125.070 204.110 ;
        RECT 131.650 204.050 131.970 204.310 ;
        RECT 27.160 203.430 139.860 203.910 ;
        RECT 29.990 203.230 30.310 203.290 ;
        RECT 31.385 203.230 31.675 203.275 ;
        RECT 29.990 203.090 31.675 203.230 ;
        RECT 29.990 203.030 30.310 203.090 ;
        RECT 31.385 203.045 31.675 203.090 ;
        RECT 37.810 203.230 38.130 203.290 ;
        RECT 40.125 203.230 40.415 203.275 ;
        RECT 37.810 203.090 40.415 203.230 ;
        RECT 37.810 203.030 38.130 203.090 ;
        RECT 40.125 203.045 40.415 203.090 ;
        RECT 41.490 203.230 41.810 203.290 ;
        RECT 42.425 203.230 42.715 203.275 ;
        RECT 41.490 203.090 42.715 203.230 ;
        RECT 41.490 203.030 41.810 203.090 ;
        RECT 42.425 203.045 42.715 203.090 ;
        RECT 49.310 203.030 49.630 203.290 ;
        RECT 51.150 203.230 51.470 203.290 ;
        RECT 53.910 203.230 54.230 203.290 ;
        RECT 49.860 203.090 54.230 203.230 ;
        RECT 41.965 202.890 42.255 202.935 ;
        RECT 42.870 202.890 43.190 202.950 ;
        RECT 44.265 202.890 44.555 202.935 ;
        RECT 41.965 202.750 44.555 202.890 ;
        RECT 41.965 202.705 42.255 202.750 ;
        RECT 42.870 202.690 43.190 202.750 ;
        RECT 44.265 202.705 44.555 202.750 ;
        RECT 44.710 202.890 45.030 202.950 ;
        RECT 46.105 202.890 46.395 202.935 ;
        RECT 44.710 202.750 46.395 202.890 ;
        RECT 44.710 202.690 45.030 202.750 ;
        RECT 46.105 202.705 46.395 202.750 ;
        RECT 47.470 202.890 47.790 202.950 ;
        RECT 49.860 202.890 50.000 203.090 ;
        RECT 51.150 203.030 51.470 203.090 ;
        RECT 53.910 203.030 54.230 203.090 ;
        RECT 57.605 203.230 57.895 203.275 ;
        RECT 59.430 203.230 59.750 203.290 ;
        RECT 57.605 203.090 59.750 203.230 ;
        RECT 57.605 203.045 57.895 203.090 ;
        RECT 59.430 203.030 59.750 203.090 ;
        RECT 65.410 203.030 65.730 203.290 ;
        RECT 82.430 203.230 82.750 203.290 ;
        RECT 83.810 203.230 84.130 203.290 ;
        RECT 82.430 203.090 84.130 203.230 ;
        RECT 82.430 203.030 82.750 203.090 ;
        RECT 83.810 203.030 84.130 203.090 ;
        RECT 84.270 203.230 84.590 203.290 ;
        RECT 89.330 203.230 89.650 203.290 ;
        RECT 84.270 203.090 89.650 203.230 ;
        RECT 84.270 203.030 84.590 203.090 ;
        RECT 89.330 203.030 89.650 203.090 ;
        RECT 91.645 203.230 91.935 203.275 ;
        RECT 110.950 203.230 111.270 203.290 ;
        RECT 91.645 203.090 111.270 203.230 ;
        RECT 91.645 203.045 91.935 203.090 ;
        RECT 110.950 203.030 111.270 203.090 ;
        RECT 112.345 203.230 112.635 203.275 ;
        RECT 117.850 203.230 118.170 203.290 ;
        RECT 112.345 203.090 118.170 203.230 ;
        RECT 112.345 203.045 112.635 203.090 ;
        RECT 117.850 203.030 118.170 203.090 ;
        RECT 126.590 203.030 126.910 203.290 ;
        RECT 127.050 203.230 127.370 203.290 ;
        RECT 130.730 203.230 131.050 203.290 ;
        RECT 127.050 203.090 131.050 203.230 ;
        RECT 127.050 203.030 127.370 203.090 ;
        RECT 130.730 203.030 131.050 203.090 ;
        RECT 47.470 202.750 50.000 202.890 ;
        RECT 50.230 202.890 50.550 202.950 ;
        RECT 52.545 202.890 52.835 202.935 ;
        RECT 62.205 202.890 62.495 202.935 ;
        RECT 67.250 202.890 67.570 202.950 ;
        RECT 50.230 202.750 52.300 202.890 ;
        RECT 47.470 202.690 47.790 202.750 ;
        RECT 50.230 202.690 50.550 202.750 ;
        RECT 32.305 202.550 32.595 202.595 ;
        RECT 32.750 202.550 33.070 202.610 ;
        RECT 32.305 202.410 33.070 202.550 ;
        RECT 32.305 202.365 32.595 202.410 ;
        RECT 32.750 202.350 33.070 202.410 ;
        RECT 38.270 202.550 38.590 202.610 ;
        RECT 45.185 202.550 45.475 202.595 ;
        RECT 45.630 202.550 45.950 202.610 ;
        RECT 38.270 202.410 44.020 202.550 ;
        RECT 38.270 202.350 38.590 202.410 ;
        RECT 41.030 202.210 41.350 202.270 ;
        RECT 42.885 202.210 43.175 202.255 ;
        RECT 41.030 202.070 43.175 202.210 ;
        RECT 43.880 202.210 44.020 202.410 ;
        RECT 45.185 202.410 45.950 202.550 ;
        RECT 45.185 202.365 45.475 202.410 ;
        RECT 45.630 202.350 45.950 202.410 ;
        RECT 48.390 202.350 48.710 202.610 ;
        RECT 49.785 202.550 50.075 202.595 ;
        RECT 50.690 202.550 51.010 202.610 ;
        RECT 49.785 202.410 51.010 202.550 ;
        RECT 49.785 202.365 50.075 202.410 ;
        RECT 49.860 202.210 50.000 202.365 ;
        RECT 50.690 202.350 51.010 202.410 ;
        RECT 51.165 202.365 51.455 202.595 ;
        RECT 43.880 202.070 50.000 202.210 ;
        RECT 51.240 202.210 51.380 202.365 ;
        RECT 51.610 202.350 51.930 202.610 ;
        RECT 52.160 202.550 52.300 202.750 ;
        RECT 52.545 202.750 60.120 202.890 ;
        RECT 52.545 202.705 52.835 202.750 ;
        RECT 59.980 202.595 60.120 202.750 ;
        RECT 62.205 202.750 67.570 202.890 ;
        RECT 62.205 202.705 62.495 202.750 ;
        RECT 67.250 202.690 67.570 202.750 ;
        RECT 69.090 202.690 69.410 202.950 ;
        RECT 70.485 202.890 70.775 202.935 ;
        RECT 70.485 202.750 77.140 202.890 ;
        RECT 70.485 202.705 70.775 202.750 ;
        RECT 77.000 202.610 77.140 202.750 ;
        RECT 87.120 202.750 89.100 202.890 ;
        RECT 52.160 202.410 59.660 202.550 ;
        RECT 52.070 202.210 52.390 202.270 ;
        RECT 55.290 202.210 55.610 202.270 ;
        RECT 51.240 202.070 55.610 202.210 ;
        RECT 41.030 202.010 41.350 202.070 ;
        RECT 42.885 202.025 43.175 202.070 ;
        RECT 42.960 201.870 43.100 202.025 ;
        RECT 52.070 202.010 52.390 202.070 ;
        RECT 55.290 202.010 55.610 202.070 ;
        RECT 58.050 202.010 58.370 202.270 ;
        RECT 58.510 202.010 58.830 202.270 ;
        RECT 59.520 202.210 59.660 202.410 ;
        RECT 59.905 202.365 60.195 202.595 ;
        RECT 60.350 202.350 60.670 202.610 ;
        RECT 61.285 202.365 61.575 202.595 ;
        RECT 63.585 202.365 63.875 202.595 ;
        RECT 64.505 202.550 64.795 202.595 ;
        RECT 65.410 202.550 65.730 202.610 ;
        RECT 64.505 202.410 65.730 202.550 ;
        RECT 64.505 202.365 64.795 202.410 ;
        RECT 61.360 202.210 61.500 202.365 ;
        RECT 61.730 202.210 62.050 202.270 ;
        RECT 59.520 202.070 62.050 202.210 ;
        RECT 61.730 202.010 62.050 202.070 ;
        RECT 62.650 202.210 62.970 202.270 ;
        RECT 63.660 202.210 63.800 202.365 ;
        RECT 65.410 202.350 65.730 202.410 ;
        RECT 69.550 202.550 69.870 202.610 ;
        RECT 70.025 202.550 70.315 202.595 ;
        RECT 69.550 202.410 70.315 202.550 ;
        RECT 69.550 202.350 69.870 202.410 ;
        RECT 70.025 202.365 70.315 202.410 ;
        RECT 72.785 202.550 73.075 202.595 ;
        RECT 74.165 202.550 74.455 202.595 ;
        RECT 72.785 202.410 74.455 202.550 ;
        RECT 72.785 202.365 73.075 202.410 ;
        RECT 74.165 202.365 74.455 202.410 ;
        RECT 74.610 202.550 74.930 202.610 ;
        RECT 75.085 202.550 75.375 202.595 ;
        RECT 74.610 202.410 75.375 202.550 ;
        RECT 62.650 202.070 64.720 202.210 ;
        RECT 62.650 202.010 62.970 202.070 ;
        RECT 47.470 201.870 47.790 201.930 ;
        RECT 42.960 201.730 47.790 201.870 ;
        RECT 47.470 201.670 47.790 201.730 ;
        RECT 50.245 201.870 50.535 201.915 ;
        RECT 55.765 201.870 56.055 201.915 ;
        RECT 50.245 201.730 56.055 201.870 ;
        RECT 58.140 201.870 58.280 202.010 ;
        RECT 64.045 201.870 64.335 201.915 ;
        RECT 58.140 201.730 64.335 201.870 ;
        RECT 64.580 201.870 64.720 202.070 ;
        RECT 66.330 202.010 66.650 202.270 ;
        RECT 66.805 202.025 67.095 202.255 ;
        RECT 66.880 201.870 67.020 202.025 ;
        RECT 67.250 202.010 67.570 202.270 ;
        RECT 67.710 202.010 68.030 202.270 ;
        RECT 71.405 202.210 71.695 202.255 ;
        RECT 71.850 202.210 72.170 202.270 ;
        RECT 71.405 202.070 72.170 202.210 ;
        RECT 74.240 202.210 74.380 202.365 ;
        RECT 74.610 202.350 74.930 202.410 ;
        RECT 75.085 202.365 75.375 202.410 ;
        RECT 75.990 202.350 76.310 202.610 ;
        RECT 76.910 202.350 77.230 202.610 ;
        RECT 77.370 202.350 77.690 202.610 ;
        RECT 78.290 202.350 78.610 202.610 ;
        RECT 80.590 202.550 80.910 202.610 ;
        RECT 82.905 202.550 83.195 202.595 ;
        RECT 80.590 202.410 83.195 202.550 ;
        RECT 80.590 202.350 80.910 202.410 ;
        RECT 82.905 202.365 83.195 202.410 ;
        RECT 83.350 202.350 83.670 202.610 ;
        RECT 74.240 202.070 74.840 202.210 ;
        RECT 71.405 202.025 71.695 202.070 ;
        RECT 71.850 202.010 72.170 202.070 ;
        RECT 74.700 201.870 74.840 202.070 ;
        RECT 75.530 202.010 75.850 202.270 ;
        RECT 81.985 202.210 82.275 202.255 ;
        RECT 87.120 202.210 87.260 202.750 ;
        RECT 87.505 202.365 87.795 202.595 ;
        RECT 81.985 202.070 87.260 202.210 ;
        RECT 81.985 202.025 82.275 202.070 ;
        RECT 82.430 201.870 82.750 201.930 ;
        RECT 87.580 201.870 87.720 202.365 ;
        RECT 88.960 202.270 89.100 202.750 ;
        RECT 93.930 202.690 94.250 202.950 ;
        RECT 94.850 202.935 95.170 202.950 ;
        RECT 94.635 202.705 95.170 202.935 ;
        RECT 94.850 202.690 95.170 202.705 ;
        RECT 97.610 202.690 97.930 202.950 ;
        RECT 98.070 202.935 98.390 202.950 ;
        RECT 98.070 202.705 98.505 202.935 ;
        RECT 98.990 202.890 99.310 202.950 ;
        RECT 99.465 202.890 99.755 202.935 ;
        RECT 104.510 202.890 104.830 202.950 ;
        RECT 98.990 202.750 99.755 202.890 ;
        RECT 98.070 202.690 98.390 202.705 ;
        RECT 98.990 202.690 99.310 202.750 ;
        RECT 99.465 202.705 99.755 202.750 ;
        RECT 100.460 202.750 104.830 202.890 ;
        RECT 90.265 202.550 90.555 202.595 ;
        RECT 90.710 202.550 91.030 202.610 ;
        RECT 90.265 202.410 91.030 202.550 ;
        RECT 90.265 202.365 90.555 202.410 ;
        RECT 90.710 202.350 91.030 202.410 ;
        RECT 93.025 202.365 93.315 202.595 ;
        RECT 87.950 202.010 88.270 202.270 ;
        RECT 88.870 202.010 89.190 202.270 ;
        RECT 64.580 201.730 74.380 201.870 ;
        RECT 74.700 201.730 82.750 201.870 ;
        RECT 50.245 201.685 50.535 201.730 ;
        RECT 55.765 201.685 56.055 201.730 ;
        RECT 64.045 201.685 64.335 201.730 ;
        RECT 44.710 201.530 45.030 201.590 ;
        RECT 71.390 201.530 71.710 201.590 ;
        RECT 44.710 201.390 71.710 201.530 ;
        RECT 44.710 201.330 45.030 201.390 ;
        RECT 71.390 201.330 71.710 201.390 ;
        RECT 71.865 201.530 72.155 201.575 ;
        RECT 72.310 201.530 72.630 201.590 ;
        RECT 71.865 201.390 72.630 201.530 ;
        RECT 71.865 201.345 72.155 201.390 ;
        RECT 72.310 201.330 72.630 201.390 ;
        RECT 73.690 201.330 74.010 201.590 ;
        RECT 74.240 201.530 74.380 201.730 ;
        RECT 82.430 201.670 82.750 201.730 ;
        RECT 83.670 201.730 87.720 201.870 ;
        RECT 93.100 201.870 93.240 202.365 ;
        RECT 93.470 202.350 93.790 202.610 ;
        RECT 95.770 202.550 96.090 202.610 ;
        RECT 100.460 202.595 100.600 202.750 ;
        RECT 104.510 202.690 104.830 202.750 ;
        RECT 106.350 202.890 106.670 202.950 ;
        RECT 107.515 202.890 107.805 202.935 ;
        RECT 106.350 202.750 107.805 202.890 ;
        RECT 106.350 202.690 106.670 202.750 ;
        RECT 107.515 202.705 107.805 202.750 ;
        RECT 108.190 202.690 108.510 202.950 ;
        RECT 108.650 202.690 108.970 202.950 ;
        RECT 110.045 202.890 110.335 202.935 ;
        RECT 112.790 202.890 113.110 202.950 ;
        RECT 116.010 202.890 116.330 202.950 ;
        RECT 110.045 202.750 116.330 202.890 ;
        RECT 110.045 202.705 110.335 202.750 ;
        RECT 112.790 202.690 113.110 202.750 ;
        RECT 116.010 202.690 116.330 202.750 ;
        RECT 96.705 202.550 96.995 202.595 ;
        RECT 95.770 202.410 96.995 202.550 ;
        RECT 95.770 202.350 96.090 202.410 ;
        RECT 96.705 202.365 96.995 202.410 ;
        RECT 97.165 202.365 97.455 202.595 ;
        RECT 100.385 202.365 100.675 202.595 ;
        RECT 93.930 202.210 94.250 202.270 ;
        RECT 95.325 202.210 95.615 202.255 ;
        RECT 93.930 202.070 95.615 202.210 ;
        RECT 97.240 202.210 97.380 202.365 ;
        RECT 100.830 202.350 101.150 202.610 ;
        RECT 103.130 202.350 103.450 202.610 ;
        RECT 103.590 202.550 103.910 202.610 ;
        RECT 103.590 202.410 104.710 202.550 ;
        RECT 103.590 202.350 103.910 202.410 ;
        RECT 99.005 202.210 99.295 202.255 ;
        RECT 101.750 202.210 102.070 202.270 ;
        RECT 97.240 202.070 98.530 202.210 ;
        RECT 93.930 202.010 94.250 202.070 ;
        RECT 95.325 202.025 95.615 202.070 ;
        RECT 94.850 201.870 95.170 201.930 ;
        RECT 93.100 201.730 95.170 201.870 ;
        RECT 95.400 201.870 95.540 202.025 ;
        RECT 97.150 201.870 97.470 201.930 ;
        RECT 95.400 201.730 97.470 201.870 ;
        RECT 98.390 201.870 98.530 202.070 ;
        RECT 99.005 202.070 102.070 202.210 ;
        RECT 99.005 202.025 99.295 202.070 ;
        RECT 101.750 202.010 102.070 202.070 ;
        RECT 102.225 202.210 102.515 202.255 ;
        RECT 104.050 202.210 104.370 202.270 ;
        RECT 102.225 202.070 104.370 202.210 ;
        RECT 104.570 202.210 104.710 202.410 ;
        RECT 104.970 202.350 105.290 202.610 ;
        RECT 106.810 202.350 107.130 202.610 ;
        RECT 109.125 202.365 109.415 202.595 ;
        RECT 109.570 202.550 109.890 202.610 ;
        RECT 110.505 202.550 110.795 202.595 ;
        RECT 109.570 202.410 110.795 202.550 ;
        RECT 109.200 202.210 109.340 202.365 ;
        RECT 109.570 202.350 109.890 202.410 ;
        RECT 110.505 202.365 110.795 202.410 ;
        RECT 111.425 202.365 111.715 202.595 ;
        RECT 112.330 202.550 112.650 202.610 ;
        RECT 117.940 202.550 118.080 203.030 ;
        RECT 121.545 202.890 121.835 202.935 ;
        RECT 126.130 202.890 126.450 202.950 ;
        RECT 121.545 202.750 126.450 202.890 ;
        RECT 121.545 202.705 121.835 202.750 ;
        RECT 126.130 202.690 126.450 202.750 ;
        RECT 122.925 202.550 123.215 202.595 ;
        RECT 127.140 202.550 127.280 203.030 ;
        RECT 128.890 202.890 129.210 202.950 ;
        RECT 131.205 202.890 131.495 202.935 ;
        RECT 128.890 202.750 131.495 202.890 ;
        RECT 128.890 202.690 129.210 202.750 ;
        RECT 131.205 202.705 131.495 202.750 ;
        RECT 112.330 202.410 114.400 202.550 ;
        RECT 117.940 202.410 123.215 202.550 ;
        RECT 104.570 202.070 109.340 202.210 ;
        RECT 102.225 202.025 102.515 202.070 ;
        RECT 104.050 202.010 104.370 202.070 ;
        RECT 99.450 201.870 99.770 201.930 ;
        RECT 101.290 201.870 101.610 201.930 ;
        RECT 105.430 201.870 105.750 201.930 ;
        RECT 105.905 201.870 106.195 201.915 ;
        RECT 111.500 201.870 111.640 202.365 ;
        RECT 112.330 202.350 112.650 202.410 ;
        RECT 112.805 202.210 113.095 202.255 ;
        RECT 98.390 201.730 98.760 201.870 ;
        RECT 77.370 201.530 77.690 201.590 ;
        RECT 74.240 201.390 77.690 201.530 ;
        RECT 77.370 201.330 77.690 201.390 ;
        RECT 77.845 201.530 78.135 201.575 ;
        RECT 81.050 201.530 81.370 201.590 ;
        RECT 83.670 201.530 83.810 201.730 ;
        RECT 94.850 201.670 95.170 201.730 ;
        RECT 97.150 201.670 97.470 201.730 ;
        RECT 77.845 201.390 83.810 201.530 ;
        RECT 84.270 201.530 84.590 201.590 ;
        RECT 85.205 201.530 85.495 201.575 ;
        RECT 84.270 201.390 85.495 201.530 ;
        RECT 77.845 201.345 78.135 201.390 ;
        RECT 81.050 201.330 81.370 201.390 ;
        RECT 84.270 201.330 84.590 201.390 ;
        RECT 85.205 201.345 85.495 201.390 ;
        RECT 85.665 201.530 85.955 201.575 ;
        RECT 86.110 201.530 86.430 201.590 ;
        RECT 85.665 201.390 86.430 201.530 ;
        RECT 85.665 201.345 85.955 201.390 ;
        RECT 86.110 201.330 86.430 201.390 ;
        RECT 92.105 201.530 92.395 201.575 ;
        RECT 93.010 201.530 93.330 201.590 ;
        RECT 92.105 201.390 93.330 201.530 ;
        RECT 92.105 201.345 92.395 201.390 ;
        RECT 93.010 201.330 93.330 201.390 ;
        RECT 95.770 201.330 96.090 201.590 ;
        RECT 98.620 201.530 98.760 201.730 ;
        RECT 99.450 201.730 106.195 201.870 ;
        RECT 99.450 201.670 99.770 201.730 ;
        RECT 101.290 201.670 101.610 201.730 ;
        RECT 105.430 201.670 105.750 201.730 ;
        RECT 105.905 201.685 106.195 201.730 ;
        RECT 108.740 201.730 111.640 201.870 ;
        RECT 112.420 202.070 113.095 202.210 ;
        RECT 114.260 202.210 114.400 202.410 ;
        RECT 122.925 202.365 123.215 202.410 ;
        RECT 125.300 202.410 127.280 202.550 ;
        RECT 127.510 202.550 127.830 202.610 ;
        RECT 129.365 202.550 129.655 202.595 ;
        RECT 127.510 202.410 129.655 202.550 ;
        RECT 125.300 202.255 125.440 202.410 ;
        RECT 127.510 202.350 127.830 202.410 ;
        RECT 129.365 202.365 129.655 202.410 ;
        RECT 134.425 202.550 134.715 202.595 ;
        RECT 134.870 202.550 135.190 202.610 ;
        RECT 134.425 202.410 135.190 202.550 ;
        RECT 134.425 202.365 134.715 202.410 ;
        RECT 134.870 202.350 135.190 202.410 ;
        RECT 136.250 202.350 136.570 202.610 ;
        RECT 136.710 202.350 137.030 202.610 ;
        RECT 122.465 202.210 122.755 202.255 ;
        RECT 114.260 202.070 122.755 202.210 ;
        RECT 108.740 201.590 108.880 201.730 ;
        RECT 112.420 201.590 112.560 202.070 ;
        RECT 112.805 202.025 113.095 202.070 ;
        RECT 122.465 202.025 122.755 202.070 ;
        RECT 125.225 202.025 125.515 202.255 ;
        RECT 131.190 202.210 131.510 202.270 ;
        RECT 131.190 202.070 132.110 202.210 ;
        RECT 131.190 202.010 131.510 202.070 ;
        RECT 114.170 201.870 114.490 201.930 ;
        RECT 131.970 201.870 132.110 202.070 ;
        RECT 135.345 201.870 135.635 201.915 ;
        RECT 114.170 201.730 131.420 201.870 ;
        RECT 131.970 201.730 135.635 201.870 ;
        RECT 114.170 201.670 114.490 201.730 ;
        RECT 131.280 201.590 131.420 201.730 ;
        RECT 135.345 201.685 135.635 201.730 ;
        RECT 99.910 201.530 100.230 201.590 ;
        RECT 100.830 201.530 101.150 201.590 ;
        RECT 98.620 201.390 101.150 201.530 ;
        RECT 99.910 201.330 100.230 201.390 ;
        RECT 100.830 201.330 101.150 201.390 ;
        RECT 102.670 201.530 102.990 201.590 ;
        RECT 104.065 201.530 104.355 201.575 ;
        RECT 108.650 201.530 108.970 201.590 ;
        RECT 102.670 201.390 108.970 201.530 ;
        RECT 102.670 201.330 102.990 201.390 ;
        RECT 104.065 201.345 104.355 201.390 ;
        RECT 108.650 201.330 108.970 201.390 ;
        RECT 112.330 201.330 112.650 201.590 ;
        RECT 114.630 201.530 114.950 201.590 ;
        RECT 123.370 201.530 123.690 201.590 ;
        RECT 114.630 201.390 123.690 201.530 ;
        RECT 114.630 201.330 114.950 201.390 ;
        RECT 123.370 201.330 123.690 201.390 ;
        RECT 123.830 201.530 124.150 201.590 ;
        RECT 124.750 201.530 125.070 201.590 ;
        RECT 123.830 201.390 125.070 201.530 ;
        RECT 123.830 201.330 124.150 201.390 ;
        RECT 124.750 201.330 125.070 201.390 ;
        RECT 131.190 201.530 131.510 201.590 ;
        RECT 133.965 201.530 134.255 201.575 ;
        RECT 131.190 201.390 134.255 201.530 ;
        RECT 131.190 201.330 131.510 201.390 ;
        RECT 133.965 201.345 134.255 201.390 ;
        RECT 137.645 201.530 137.935 201.575 ;
        RECT 138.090 201.530 138.410 201.590 ;
        RECT 137.645 201.390 138.410 201.530 ;
        RECT 137.645 201.345 137.935 201.390 ;
        RECT 138.090 201.330 138.410 201.390 ;
        RECT 27.160 200.710 139.860 201.190 ;
        RECT 38.270 200.510 38.590 200.570 ;
        RECT 39.205 200.510 39.495 200.555 ;
        RECT 38.270 200.370 39.495 200.510 ;
        RECT 38.270 200.310 38.590 200.370 ;
        RECT 39.205 200.325 39.495 200.370 ;
        RECT 47.025 200.510 47.315 200.555 ;
        RECT 48.390 200.510 48.710 200.570 ;
        RECT 47.025 200.370 48.710 200.510 ;
        RECT 47.025 200.325 47.315 200.370 ;
        RECT 48.390 200.310 48.710 200.370 ;
        RECT 54.370 200.510 54.690 200.570 ;
        RECT 54.845 200.510 55.135 200.555 ;
        RECT 60.350 200.510 60.670 200.570 ;
        RECT 54.370 200.370 55.135 200.510 ;
        RECT 54.370 200.310 54.690 200.370 ;
        RECT 54.845 200.325 55.135 200.370 ;
        RECT 55.380 200.370 60.670 200.510 ;
        RECT 48.850 200.170 49.170 200.230 ;
        RECT 49.325 200.170 49.615 200.215 ;
        RECT 48.850 200.030 49.615 200.170 ;
        RECT 48.850 199.970 49.170 200.030 ;
        RECT 49.325 199.985 49.615 200.030 ;
        RECT 52.545 200.170 52.835 200.215 ;
        RECT 52.990 200.170 53.310 200.230 ;
        RECT 55.380 200.170 55.520 200.370 ;
        RECT 60.350 200.310 60.670 200.370 ;
        RECT 67.250 200.510 67.570 200.570 ;
        RECT 67.250 200.370 70.010 200.510 ;
        RECT 67.250 200.310 67.570 200.370 ;
        RECT 63.125 200.170 63.415 200.215 ;
        RECT 52.545 200.030 55.520 200.170 ;
        RECT 57.220 200.030 63.415 200.170 ;
        RECT 52.545 199.985 52.835 200.030 ;
        RECT 52.990 199.970 53.310 200.030 ;
        RECT 57.220 199.890 57.360 200.030 ;
        RECT 63.125 199.985 63.415 200.030 ;
        RECT 64.030 200.170 64.350 200.230 ;
        RECT 69.105 200.170 69.395 200.215 ;
        RECT 64.030 200.030 69.395 200.170 ;
        RECT 69.870 200.170 70.010 200.370 ;
        RECT 70.930 200.310 71.250 200.570 ;
        RECT 77.830 200.510 78.150 200.570 ;
        RECT 80.145 200.510 80.435 200.555 ;
        RECT 77.830 200.370 80.435 200.510 ;
        RECT 77.830 200.310 78.150 200.370 ;
        RECT 80.145 200.325 80.435 200.370 ;
        RECT 88.870 200.510 89.190 200.570 ;
        RECT 95.325 200.510 95.615 200.555 ;
        RECT 108.205 200.510 108.495 200.555 ;
        RECT 113.250 200.510 113.570 200.570 ;
        RECT 88.870 200.370 95.615 200.510 ;
        RECT 88.870 200.310 89.190 200.370 ;
        RECT 95.325 200.325 95.615 200.370 ;
        RECT 95.860 200.370 113.570 200.510 ;
        RECT 78.290 200.170 78.610 200.230 ;
        RECT 69.870 200.030 78.610 200.170 ;
        RECT 64.030 199.970 64.350 200.030 ;
        RECT 69.105 199.985 69.395 200.030 ;
        RECT 78.290 199.970 78.610 200.030 ;
        RECT 79.225 200.170 79.515 200.215 ;
        RECT 83.350 200.170 83.670 200.230 ;
        RECT 79.225 200.030 83.670 200.170 ;
        RECT 79.225 199.985 79.515 200.030 ;
        RECT 83.350 199.970 83.670 200.030 ;
        RECT 86.110 199.970 86.430 200.230 ;
        RECT 90.710 200.170 91.030 200.230 ;
        RECT 95.860 200.170 96.000 200.370 ;
        RECT 108.205 200.325 108.495 200.370 ;
        RECT 113.250 200.310 113.570 200.370 ;
        RECT 116.930 200.510 117.250 200.570 ;
        RECT 126.590 200.510 126.910 200.570 ;
        RECT 116.930 200.370 126.910 200.510 ;
        RECT 116.930 200.310 117.250 200.370 ;
        RECT 126.590 200.310 126.910 200.370 ;
        RECT 127.970 200.510 128.290 200.570 ;
        RECT 127.970 200.370 138.320 200.510 ;
        RECT 127.970 200.310 128.290 200.370 ;
        RECT 90.710 200.030 96.000 200.170 ;
        RECT 100.845 200.170 101.135 200.215 ;
        RECT 111.870 200.170 112.190 200.230 ;
        RECT 100.845 200.030 112.190 200.170 ;
        RECT 90.710 199.970 91.030 200.030 ;
        RECT 100.845 199.985 101.135 200.030 ;
        RECT 111.870 199.970 112.190 200.030 ;
        RECT 120.150 200.170 120.470 200.230 ;
        RECT 123.370 200.170 123.690 200.230 ;
        RECT 120.150 200.030 123.690 200.170 ;
        RECT 120.150 199.970 120.470 200.030 ;
        RECT 123.370 199.970 123.690 200.030 ;
        RECT 125.670 199.970 125.990 200.230 ;
        RECT 133.045 200.170 133.335 200.215 ;
        RECT 131.970 200.030 133.335 200.170 ;
        RECT 44.725 199.830 45.015 199.875 ;
        RECT 54.830 199.830 55.150 199.890 ;
        RECT 38.820 199.690 45.015 199.830 ;
        RECT 36.430 199.490 36.750 199.550 ;
        RECT 38.820 199.535 38.960 199.690 ;
        RECT 38.745 199.490 39.035 199.535 ;
        RECT 36.430 199.350 39.035 199.490 ;
        RECT 36.430 199.290 36.750 199.350 ;
        RECT 38.745 199.305 39.035 199.350 ;
        RECT 39.190 199.490 39.510 199.550 ;
        RECT 42.500 199.535 42.640 199.690 ;
        RECT 44.725 199.645 45.015 199.690 ;
        RECT 46.640 199.690 55.150 199.830 ;
        RECT 46.640 199.535 46.780 199.690 ;
        RECT 54.830 199.630 55.150 199.690 ;
        RECT 57.130 199.630 57.450 199.890 ;
        RECT 57.605 199.830 57.895 199.875 ;
        RECT 58.510 199.830 58.830 199.890 ;
        RECT 57.605 199.690 58.830 199.830 ;
        RECT 57.605 199.645 57.895 199.690 ;
        RECT 39.665 199.490 39.955 199.535 ;
        RECT 41.965 199.490 42.255 199.535 ;
        RECT 39.190 199.350 42.255 199.490 ;
        RECT 39.190 199.290 39.510 199.350 ;
        RECT 39.665 199.305 39.955 199.350 ;
        RECT 41.965 199.305 42.255 199.350 ;
        RECT 42.425 199.305 42.715 199.535 ;
        RECT 45.185 199.490 45.475 199.535 ;
        RECT 46.565 199.490 46.855 199.535 ;
        RECT 45.185 199.350 46.855 199.490 ;
        RECT 45.185 199.305 45.475 199.350 ;
        RECT 46.565 199.305 46.855 199.350 ;
        RECT 42.040 198.810 42.180 199.305 ;
        RECT 47.470 199.290 47.790 199.550 ;
        RECT 47.930 199.290 48.250 199.550 ;
        RECT 48.405 199.490 48.695 199.535 ;
        RECT 49.770 199.490 50.090 199.550 ;
        RECT 48.405 199.350 50.090 199.490 ;
        RECT 48.405 199.305 48.695 199.350 ;
        RECT 49.770 199.290 50.090 199.350 ;
        RECT 56.670 199.290 56.990 199.550 ;
        RECT 43.330 198.950 43.650 199.210 ;
        RECT 49.325 199.150 49.615 199.195 ;
        RECT 50.230 199.150 50.550 199.210 ;
        RECT 49.325 199.010 50.550 199.150 ;
        RECT 49.325 198.965 49.615 199.010 ;
        RECT 50.230 198.950 50.550 199.010 ;
        RECT 53.465 198.965 53.755 199.195 ;
        RECT 54.370 199.150 54.690 199.210 ;
        RECT 57.680 199.150 57.820 199.645 ;
        RECT 58.510 199.630 58.830 199.690 ;
        RECT 65.870 199.830 66.190 199.890 ;
        RECT 70.025 199.830 70.315 199.875 ;
        RECT 73.690 199.830 74.010 199.890 ;
        RECT 65.870 199.690 68.860 199.830 ;
        RECT 65.870 199.630 66.190 199.690 ;
        RECT 68.720 199.550 68.860 199.690 ;
        RECT 70.025 199.690 74.010 199.830 ;
        RECT 70.025 199.645 70.315 199.690 ;
        RECT 73.690 199.630 74.010 199.690 ;
        RECT 74.150 199.830 74.470 199.890 ;
        RECT 74.150 199.690 79.900 199.830 ;
        RECT 74.150 199.630 74.470 199.690 ;
        RECT 62.650 199.290 62.970 199.550 ;
        RECT 63.585 199.490 63.875 199.535 ;
        RECT 66.330 199.490 66.650 199.550 ;
        RECT 67.250 199.490 67.570 199.550 ;
        RECT 63.585 199.350 67.570 199.490 ;
        RECT 63.585 199.305 63.875 199.350 ;
        RECT 66.330 199.290 66.650 199.350 ;
        RECT 67.250 199.290 67.570 199.350 ;
        RECT 68.630 199.290 68.950 199.550 ;
        RECT 77.370 199.490 77.690 199.550 ;
        RECT 79.760 199.535 79.900 199.690 ;
        RECT 81.050 199.630 81.370 199.890 ;
        RECT 81.510 199.830 81.830 199.890 ;
        RECT 82.905 199.830 83.195 199.875 ;
        RECT 87.950 199.830 88.270 199.890 ;
        RECT 98.530 199.830 98.850 199.890 ;
        RECT 101.290 199.830 101.610 199.890 ;
        RECT 112.330 199.830 112.650 199.890 ;
        RECT 81.510 199.690 83.195 199.830 ;
        RECT 81.510 199.630 81.830 199.690 ;
        RECT 82.905 199.645 83.195 199.690 ;
        RECT 86.200 199.690 88.270 199.830 ;
        RECT 78.765 199.490 79.055 199.535 ;
        RECT 77.370 199.350 79.055 199.490 ;
        RECT 77.370 199.290 77.690 199.350 ;
        RECT 78.765 199.305 79.055 199.350 ;
        RECT 79.685 199.490 79.975 199.535 ;
        RECT 80.130 199.490 80.450 199.550 ;
        RECT 79.685 199.350 80.450 199.490 ;
        RECT 81.140 199.490 81.280 199.630 ;
        RECT 81.985 199.490 82.275 199.535 ;
        RECT 81.140 199.350 82.275 199.490 ;
        RECT 79.685 199.305 79.975 199.350 ;
        RECT 80.130 199.290 80.450 199.350 ;
        RECT 81.985 199.305 82.275 199.350 ;
        RECT 83.350 199.490 83.670 199.550 ;
        RECT 85.205 199.490 85.495 199.535 ;
        RECT 83.350 199.350 85.495 199.490 ;
        RECT 83.350 199.290 83.670 199.350 ;
        RECT 85.205 199.305 85.495 199.350 ;
        RECT 85.650 199.290 85.970 199.550 ;
        RECT 79.210 199.150 79.530 199.210 ;
        RECT 54.370 199.010 57.820 199.150 ;
        RECT 58.140 199.010 79.530 199.150 ;
        RECT 47.470 198.810 47.790 198.870 ;
        RECT 42.040 198.670 47.790 198.810 ;
        RECT 47.470 198.610 47.790 198.670 ;
        RECT 48.390 198.810 48.710 198.870 ;
        RECT 53.540 198.810 53.680 198.965 ;
        RECT 54.370 198.950 54.690 199.010 ;
        RECT 48.390 198.670 53.680 198.810 ;
        RECT 57.130 198.810 57.450 198.870 ;
        RECT 58.140 198.810 58.280 199.010 ;
        RECT 79.210 198.950 79.530 199.010 ;
        RECT 81.050 199.150 81.370 199.210 ;
        RECT 82.445 199.150 82.735 199.195 ;
        RECT 86.200 199.150 86.340 199.690 ;
        RECT 87.950 199.630 88.270 199.690 ;
        RECT 95.860 199.690 96.920 199.830 ;
        RECT 86.585 199.305 86.875 199.535 ;
        RECT 81.050 199.010 86.340 199.150 ;
        RECT 86.660 199.150 86.800 199.305 ;
        RECT 87.490 199.290 87.810 199.550 ;
        RECT 88.425 199.490 88.715 199.535 ;
        RECT 88.870 199.490 89.190 199.550 ;
        RECT 88.425 199.350 89.190 199.490 ;
        RECT 88.425 199.305 88.715 199.350 ;
        RECT 88.870 199.290 89.190 199.350 ;
        RECT 93.010 199.290 93.330 199.550 ;
        RECT 94.405 199.490 94.695 199.535 ;
        RECT 95.860 199.490 96.000 199.690 ;
        RECT 96.780 199.535 96.920 199.690 ;
        RECT 98.530 199.690 101.610 199.830 ;
        RECT 98.530 199.630 98.850 199.690 ;
        RECT 94.405 199.350 96.000 199.490 ;
        RECT 96.705 199.490 96.995 199.535 ;
        RECT 98.085 199.490 98.375 199.535 ;
        RECT 99.450 199.490 99.770 199.550 ;
        RECT 100.000 199.535 100.140 199.690 ;
        RECT 101.290 199.630 101.610 199.690 ;
        RECT 101.840 199.690 112.650 199.830 ;
        RECT 101.840 199.535 101.980 199.690 ;
        RECT 96.705 199.350 97.840 199.490 ;
        RECT 94.405 199.305 94.695 199.350 ;
        RECT 96.705 199.305 96.995 199.350 ;
        RECT 87.965 199.150 88.255 199.195 ;
        RECT 86.660 199.010 88.255 199.150 ;
        RECT 81.050 198.950 81.370 199.010 ;
        RECT 82.445 198.965 82.735 199.010 ;
        RECT 87.965 198.965 88.255 199.010 ;
        RECT 95.310 198.950 95.630 199.210 ;
        RECT 57.130 198.670 58.280 198.810 ;
        RECT 63.110 198.810 63.430 198.870 ;
        RECT 65.410 198.810 65.730 198.870 ;
        RECT 63.110 198.670 65.730 198.810 ;
        RECT 48.390 198.610 48.710 198.670 ;
        RECT 57.130 198.610 57.450 198.670 ;
        RECT 63.110 198.610 63.430 198.670 ;
        RECT 65.410 198.610 65.730 198.670 ;
        RECT 71.390 198.810 71.710 198.870 ;
        RECT 83.350 198.810 83.670 198.870 ;
        RECT 71.390 198.670 83.670 198.810 ;
        RECT 71.390 198.610 71.710 198.670 ;
        RECT 83.350 198.610 83.670 198.670 ;
        RECT 84.285 198.810 84.575 198.855 ;
        RECT 87.030 198.810 87.350 198.870 ;
        RECT 84.285 198.670 87.350 198.810 ;
        RECT 84.285 198.625 84.575 198.670 ;
        RECT 87.030 198.610 87.350 198.670 ;
        RECT 88.410 198.810 88.730 198.870 ;
        RECT 92.105 198.810 92.395 198.855 ;
        RECT 88.410 198.670 92.395 198.810 ;
        RECT 88.410 198.610 88.730 198.670 ;
        RECT 92.105 198.625 92.395 198.670 ;
        RECT 93.930 198.810 94.250 198.870 ;
        RECT 96.245 198.810 96.535 198.855 ;
        RECT 93.930 198.670 96.535 198.810 ;
        RECT 93.930 198.610 94.250 198.670 ;
        RECT 96.245 198.625 96.535 198.670 ;
        RECT 97.150 198.610 97.470 198.870 ;
        RECT 97.700 198.810 97.840 199.350 ;
        RECT 98.085 199.350 99.770 199.490 ;
        RECT 98.085 199.305 98.375 199.350 ;
        RECT 99.450 199.290 99.770 199.350 ;
        RECT 99.925 199.305 100.215 199.535 ;
        RECT 101.765 199.305 102.055 199.535 ;
        RECT 103.605 199.305 103.895 199.535 ;
        RECT 98.530 198.950 98.850 199.210 ;
        RECT 99.005 199.150 99.295 199.195 ;
        RECT 102.670 199.150 102.990 199.210 ;
        RECT 99.005 199.010 102.990 199.150 ;
        RECT 103.680 199.150 103.820 199.305 ;
        RECT 105.430 199.290 105.750 199.550 ;
        RECT 105.890 199.290 106.210 199.550 ;
        RECT 107.285 199.490 107.575 199.535 ;
        RECT 108.650 199.490 108.970 199.550 ;
        RECT 107.285 199.350 108.970 199.490 ;
        RECT 107.285 199.305 107.575 199.350 ;
        RECT 108.650 199.290 108.970 199.350 ;
        RECT 109.110 199.290 109.430 199.550 ;
        RECT 110.030 199.290 110.350 199.550 ;
        RECT 110.965 199.490 111.255 199.535 ;
        RECT 111.410 199.490 111.730 199.550 ;
        RECT 111.960 199.535 112.100 199.690 ;
        RECT 112.330 199.630 112.650 199.690 ;
        RECT 112.805 199.830 113.095 199.875 ;
        RECT 114.170 199.830 114.490 199.890 ;
        RECT 112.805 199.690 114.490 199.830 ;
        RECT 112.805 199.645 113.095 199.690 ;
        RECT 114.170 199.630 114.490 199.690 ;
        RECT 114.630 199.630 114.950 199.890 ;
        RECT 115.105 199.830 115.395 199.875 ;
        RECT 125.760 199.830 125.900 199.970 ;
        RECT 115.105 199.690 125.900 199.830 ;
        RECT 127.510 199.830 127.830 199.890 ;
        RECT 131.970 199.830 132.110 200.030 ;
        RECT 133.045 199.985 133.335 200.030 ;
        RECT 127.510 199.690 132.110 199.830 ;
        RECT 135.790 199.830 136.110 199.890 ;
        RECT 136.725 199.830 137.015 199.875 ;
        RECT 135.790 199.690 137.015 199.830 ;
        RECT 115.105 199.645 115.395 199.690 ;
        RECT 127.510 199.630 127.830 199.690 ;
        RECT 135.790 199.630 136.110 199.690 ;
        RECT 136.725 199.645 137.015 199.690 ;
        RECT 110.965 199.350 111.730 199.490 ;
        RECT 110.965 199.305 111.255 199.350 ;
        RECT 111.410 199.290 111.730 199.350 ;
        RECT 111.885 199.305 112.175 199.535 ;
        RECT 113.710 199.490 114.030 199.550 ;
        RECT 112.880 199.350 114.030 199.490 ;
        RECT 103.680 199.010 105.200 199.150 ;
        RECT 99.005 198.965 99.295 199.010 ;
        RECT 102.670 198.950 102.990 199.010 ;
        RECT 104.525 198.810 104.815 198.855 ;
        RECT 97.700 198.670 104.815 198.810 ;
        RECT 105.060 198.810 105.200 199.010 ;
        RECT 106.350 198.950 106.670 199.210 ;
        RECT 112.330 199.150 112.650 199.210 ;
        RECT 106.900 199.010 112.650 199.150 ;
        RECT 106.900 198.810 107.040 199.010 ;
        RECT 112.330 198.950 112.650 199.010 ;
        RECT 105.060 198.670 107.040 198.810 ;
        RECT 111.425 198.810 111.715 198.855 ;
        RECT 112.880 198.810 113.020 199.350 ;
        RECT 113.710 199.290 114.030 199.350 ;
        RECT 115.550 199.290 115.870 199.550 ;
        RECT 116.025 199.490 116.315 199.535 ;
        RECT 116.470 199.490 116.790 199.550 ;
        RECT 116.025 199.350 116.790 199.490 ;
        RECT 116.025 199.305 116.315 199.350 ;
        RECT 116.470 199.290 116.790 199.350 ;
        RECT 116.930 199.290 117.250 199.550 ;
        RECT 122.465 199.490 122.755 199.535 ;
        RECT 117.480 199.350 122.755 199.490 ;
        RECT 113.250 199.150 113.570 199.210 ;
        RECT 117.480 199.150 117.620 199.350 ;
        RECT 122.465 199.305 122.755 199.350 ;
        RECT 122.925 199.305 123.215 199.535 ;
        RECT 113.250 199.010 117.620 199.150 ;
        RECT 123.000 199.150 123.140 199.305 ;
        RECT 123.370 199.290 123.690 199.550 ;
        RECT 125.685 199.490 125.975 199.535 ;
        RECT 127.970 199.490 128.290 199.550 ;
        RECT 125.685 199.350 128.290 199.490 ;
        RECT 125.685 199.305 125.975 199.350 ;
        RECT 127.970 199.290 128.290 199.350 ;
        RECT 137.630 199.290 137.950 199.550 ;
        RECT 138.180 199.535 138.320 200.370 ;
        RECT 138.105 199.305 138.395 199.535 ;
        RECT 124.290 199.150 124.610 199.210 ;
        RECT 126.605 199.150 126.895 199.195 ;
        RECT 123.000 199.010 123.600 199.150 ;
        RECT 113.250 198.950 113.570 199.010 ;
        RECT 123.460 198.870 123.600 199.010 ;
        RECT 124.290 199.010 126.895 199.150 ;
        RECT 124.290 198.950 124.610 199.010 ;
        RECT 126.605 198.965 126.895 199.010 ;
        RECT 135.330 199.150 135.650 199.210 ;
        RECT 136.725 199.150 137.015 199.195 ;
        RECT 135.330 199.010 137.015 199.150 ;
        RECT 135.330 198.950 135.650 199.010 ;
        RECT 136.725 198.965 137.015 199.010 ;
        RECT 111.425 198.670 113.020 198.810 ;
        RECT 113.725 198.810 114.015 198.855 ;
        RECT 121.070 198.810 121.390 198.870 ;
        RECT 113.725 198.670 121.390 198.810 ;
        RECT 104.525 198.625 104.815 198.670 ;
        RECT 111.425 198.625 111.715 198.670 ;
        RECT 113.725 198.625 114.015 198.670 ;
        RECT 121.070 198.610 121.390 198.670 ;
        RECT 123.370 198.610 123.690 198.870 ;
        RECT 124.750 198.610 125.070 198.870 ;
        RECT 125.670 198.810 125.990 198.870 ;
        RECT 131.650 198.810 131.970 198.870 ;
        RECT 125.670 198.670 131.970 198.810 ;
        RECT 125.670 198.610 125.990 198.670 ;
        RECT 131.650 198.610 131.970 198.670 ;
        RECT 135.790 198.610 136.110 198.870 ;
        RECT 27.160 197.990 139.860 198.470 ;
        RECT 44.710 197.790 45.030 197.850 ;
        RECT 46.090 197.790 46.410 197.850 ;
        RECT 44.710 197.650 46.410 197.790 ;
        RECT 44.710 197.590 45.030 197.650 ;
        RECT 46.090 197.590 46.410 197.650 ;
        RECT 66.790 197.590 67.110 197.850 ;
        RECT 67.710 197.590 68.030 197.850 ;
        RECT 68.170 197.790 68.490 197.850 ;
        RECT 69.550 197.790 69.870 197.850 ;
        RECT 71.865 197.790 72.155 197.835 ;
        RECT 68.170 197.650 69.320 197.790 ;
        RECT 68.170 197.590 68.490 197.650 ;
        RECT 36.445 197.450 36.735 197.495 ;
        RECT 41.045 197.450 41.335 197.495 ;
        RECT 45.170 197.450 45.490 197.510 ;
        RECT 36.445 197.310 45.490 197.450 ;
        RECT 36.445 197.265 36.735 197.310 ;
        RECT 41.045 197.265 41.335 197.310 ;
        RECT 45.170 197.250 45.490 197.310 ;
        RECT 50.230 197.450 50.550 197.510 ;
        RECT 52.525 197.450 52.815 197.495 ;
        RECT 50.230 197.310 52.815 197.450 ;
        RECT 50.230 197.250 50.550 197.310 ;
        RECT 52.525 197.265 52.815 197.310 ;
        RECT 56.670 197.450 56.990 197.510 ;
        RECT 60.810 197.450 61.130 197.510 ;
        RECT 56.670 197.310 61.130 197.450 ;
        RECT 56.670 197.250 56.990 197.310 ;
        RECT 60.810 197.250 61.130 197.310 ;
        RECT 62.650 197.450 62.970 197.510 ;
        RECT 69.180 197.450 69.320 197.650 ;
        RECT 69.550 197.650 72.155 197.790 ;
        RECT 69.550 197.590 69.870 197.650 ;
        RECT 71.865 197.605 72.155 197.650 ;
        RECT 81.050 197.590 81.370 197.850 ;
        RECT 81.510 197.790 81.830 197.850 ;
        RECT 93.515 197.790 93.805 197.835 ;
        RECT 95.310 197.790 95.630 197.850 ;
        RECT 98.085 197.790 98.375 197.835 ;
        RECT 81.510 197.650 93.805 197.790 ;
        RECT 81.510 197.590 81.830 197.650 ;
        RECT 93.515 197.605 93.805 197.650 ;
        RECT 94.020 197.650 98.375 197.790 ;
        RECT 72.325 197.450 72.615 197.495 ;
        RECT 62.650 197.310 67.020 197.450 ;
        RECT 69.180 197.310 72.615 197.450 ;
        RECT 62.650 197.250 62.970 197.310 ;
        RECT 36.905 197.110 37.195 197.155 ;
        RECT 37.350 197.110 37.670 197.170 ;
        RECT 40.585 197.110 40.875 197.155 ;
        RECT 36.905 196.970 40.875 197.110 ;
        RECT 36.905 196.925 37.195 196.970 ;
        RECT 37.350 196.910 37.670 196.970 ;
        RECT 40.585 196.925 40.875 196.970 ;
        RECT 48.390 197.110 48.710 197.170 ;
        RECT 49.785 197.110 50.075 197.155 ;
        RECT 48.390 196.970 50.075 197.110 ;
        RECT 48.390 196.910 48.710 196.970 ;
        RECT 49.785 196.925 50.075 196.970 ;
        RECT 51.165 196.925 51.455 197.155 ;
        RECT 51.625 197.110 51.915 197.155 ;
        RECT 52.990 197.110 53.310 197.170 ;
        RECT 51.625 196.970 53.310 197.110 ;
        RECT 51.625 196.925 51.915 196.970 ;
        RECT 35.985 196.770 36.275 196.815 ;
        RECT 39.665 196.770 39.955 196.815 ;
        RECT 41.030 196.770 41.350 196.830 ;
        RECT 35.985 196.630 41.350 196.770 ;
        RECT 35.985 196.585 36.275 196.630 ;
        RECT 39.665 196.585 39.955 196.630 ;
        RECT 41.030 196.570 41.350 196.630 ;
        RECT 44.710 196.770 45.030 196.830 ;
        RECT 51.240 196.770 51.380 196.925 ;
        RECT 52.990 196.910 53.310 196.970 ;
        RECT 64.950 196.910 65.270 197.170 ;
        RECT 65.410 197.110 65.730 197.170 ;
        RECT 66.880 197.155 67.020 197.310 ;
        RECT 68.260 197.265 68.860 197.280 ;
        RECT 72.325 197.265 72.615 197.310 ;
        RECT 79.210 197.450 79.530 197.510 ;
        RECT 93.025 197.450 93.315 197.495 ;
        RECT 94.020 197.450 94.160 197.650 ;
        RECT 95.310 197.590 95.630 197.650 ;
        RECT 98.085 197.605 98.375 197.650 ;
        RECT 103.590 197.790 103.910 197.850 ;
        RECT 107.730 197.790 108.050 197.850 ;
        RECT 119.690 197.790 120.010 197.850 ;
        RECT 123.830 197.790 124.150 197.850 ;
        RECT 103.590 197.650 108.050 197.790 ;
        RECT 103.590 197.590 103.910 197.650 ;
        RECT 107.730 197.590 108.050 197.650 ;
        RECT 109.200 197.650 124.150 197.790 ;
        RECT 97.150 197.450 97.470 197.510 ;
        RECT 79.210 197.310 92.780 197.450 ;
        RECT 66.345 197.110 66.635 197.155 ;
        RECT 65.410 196.970 66.635 197.110 ;
        RECT 65.410 196.910 65.730 196.970 ;
        RECT 66.345 196.925 66.635 196.970 ;
        RECT 66.805 196.925 67.095 197.155 ;
        RECT 68.260 197.140 68.940 197.265 ;
        RECT 79.210 197.250 79.530 197.310 ;
        RECT 68.260 197.110 68.400 197.140 ;
        RECT 67.340 196.970 68.400 197.110 ;
        RECT 68.650 197.035 68.940 197.140 ;
        RECT 44.710 196.630 51.380 196.770 ;
        RECT 63.110 196.770 63.430 196.830 ;
        RECT 67.340 196.770 67.480 196.970 ;
        RECT 69.105 196.925 69.395 197.155 ;
        RECT 63.110 196.630 67.480 196.770 ;
        RECT 44.710 196.570 45.030 196.630 ;
        RECT 63.110 196.570 63.430 196.630 ;
        RECT 38.745 196.430 39.035 196.475 ;
        RECT 41.950 196.430 42.270 196.490 ;
        RECT 38.745 196.290 42.270 196.430 ;
        RECT 38.745 196.245 39.035 196.290 ;
        RECT 41.950 196.230 42.270 196.290 ;
        RECT 43.330 196.430 43.650 196.490 ;
        RECT 50.230 196.430 50.550 196.490 ;
        RECT 67.340 196.430 67.480 196.630 ;
        RECT 67.710 196.770 68.030 196.830 ;
        RECT 69.180 196.770 69.320 196.925 ;
        RECT 69.550 196.910 69.870 197.170 ;
        RECT 70.010 197.155 70.330 197.170 ;
        RECT 70.010 196.925 70.445 197.155 ;
        RECT 71.390 197.110 71.710 197.170 ;
        RECT 79.685 197.110 79.975 197.155 ;
        RECT 71.390 196.970 79.975 197.110 ;
        RECT 70.010 196.910 70.330 196.925 ;
        RECT 71.390 196.910 71.710 196.970 ;
        RECT 79.685 196.925 79.975 196.970 ;
        RECT 83.350 196.910 83.670 197.170 ;
        RECT 84.270 196.910 84.590 197.170 ;
        RECT 84.730 196.910 85.050 197.170 ;
        RECT 91.645 197.110 91.935 197.155 ;
        RECT 91.260 196.970 91.935 197.110 ;
        RECT 92.640 197.110 92.780 197.310 ;
        RECT 93.025 197.310 94.160 197.450 ;
        RECT 94.480 197.310 97.470 197.450 ;
        RECT 93.025 197.265 93.315 197.310 ;
        RECT 93.930 197.110 94.250 197.170 ;
        RECT 94.480 197.155 94.620 197.310 ;
        RECT 97.150 197.250 97.470 197.310 ;
        RECT 98.530 197.450 98.850 197.510 ;
        RECT 106.365 197.450 106.655 197.495 ;
        RECT 98.530 197.310 105.200 197.450 ;
        RECT 98.530 197.250 98.850 197.310 ;
        RECT 92.640 196.970 94.250 197.110 ;
        RECT 91.260 196.830 91.400 196.970 ;
        RECT 91.645 196.925 91.935 196.970 ;
        RECT 93.930 196.910 94.250 196.970 ;
        RECT 94.405 196.925 94.695 197.155 ;
        RECT 94.850 196.910 95.170 197.170 ;
        RECT 95.785 196.925 96.075 197.155 ;
        RECT 67.710 196.630 69.320 196.770 ;
        RECT 70.945 196.770 71.235 196.815 ;
        RECT 73.690 196.770 74.010 196.830 ;
        RECT 81.065 196.770 81.355 196.815 ;
        RECT 70.945 196.630 81.355 196.770 ;
        RECT 67.710 196.570 68.030 196.630 ;
        RECT 70.945 196.585 71.235 196.630 ;
        RECT 73.690 196.570 74.010 196.630 ;
        RECT 81.065 196.585 81.355 196.630 ;
        RECT 83.825 196.770 84.115 196.815 ;
        RECT 85.650 196.770 85.970 196.830 ;
        RECT 83.825 196.630 85.970 196.770 ;
        RECT 83.825 196.585 84.115 196.630 ;
        RECT 85.650 196.570 85.970 196.630 ;
        RECT 91.170 196.570 91.490 196.830 ;
        RECT 93.470 196.770 93.790 196.830 ;
        RECT 95.860 196.770 96.000 196.925 ;
        RECT 96.690 196.910 97.010 197.170 ;
        RECT 99.005 197.110 99.295 197.155 ;
        RECT 99.450 197.110 99.770 197.170 ;
        RECT 100.920 197.155 101.060 197.310 ;
        RECT 99.005 196.970 99.770 197.110 ;
        RECT 99.005 196.925 99.295 196.970 ;
        RECT 99.450 196.910 99.770 196.970 ;
        RECT 100.845 196.925 101.135 197.155 ;
        RECT 101.750 196.910 102.070 197.170 ;
        RECT 102.210 197.110 102.530 197.170 ;
        RECT 105.060 197.155 105.200 197.310 ;
        RECT 106.365 197.310 107.960 197.450 ;
        RECT 106.365 197.265 106.655 197.310 ;
        RECT 103.145 197.110 103.435 197.155 ;
        RECT 102.210 196.970 103.435 197.110 ;
        RECT 102.210 196.910 102.530 196.970 ;
        RECT 103.145 196.925 103.435 196.970 ;
        RECT 104.985 197.110 105.275 197.155 ;
        RECT 105.890 197.110 106.210 197.170 ;
        RECT 104.985 196.970 106.210 197.110 ;
        RECT 104.985 196.925 105.275 196.970 ;
        RECT 105.890 196.910 106.210 196.970 ;
        RECT 107.285 196.925 107.575 197.155 ;
        RECT 97.150 196.770 97.470 196.830 ;
        RECT 93.470 196.630 95.540 196.770 ;
        RECT 95.860 196.630 97.470 196.770 ;
        RECT 93.470 196.570 93.790 196.630 ;
        RECT 69.090 196.430 69.410 196.490 ;
        RECT 94.390 196.430 94.710 196.490 ;
        RECT 43.330 196.290 66.100 196.430 ;
        RECT 67.340 196.290 94.710 196.430 ;
        RECT 95.400 196.430 95.540 196.630 ;
        RECT 97.150 196.570 97.470 196.630 ;
        RECT 99.910 196.570 100.230 196.830 ;
        RECT 100.385 196.770 100.675 196.815 ;
        RECT 102.670 196.770 102.990 196.830 ;
        RECT 100.385 196.630 102.990 196.770 ;
        RECT 100.385 196.585 100.675 196.630 ;
        RECT 102.670 196.570 102.990 196.630 ;
        RECT 104.065 196.585 104.355 196.815 ;
        RECT 104.510 196.770 104.830 196.830 ;
        RECT 107.360 196.770 107.500 196.925 ;
        RECT 107.820 196.830 107.960 197.310 ;
        RECT 109.200 197.155 109.340 197.650 ;
        RECT 119.690 197.590 120.010 197.650 ;
        RECT 123.830 197.590 124.150 197.650 ;
        RECT 125.670 197.590 125.990 197.850 ;
        RECT 129.810 197.790 130.130 197.850 ;
        RECT 131.205 197.790 131.495 197.835 ;
        RECT 127.140 197.650 129.080 197.790 ;
        RECT 110.045 197.450 110.335 197.495 ;
        RECT 110.950 197.450 111.270 197.510 ;
        RECT 115.550 197.450 115.870 197.510 ;
        RECT 110.045 197.310 111.270 197.450 ;
        RECT 110.045 197.265 110.335 197.310 ;
        RECT 110.950 197.250 111.270 197.310 ;
        RECT 112.880 197.310 115.870 197.450 ;
        RECT 109.125 196.925 109.415 197.155 ;
        RECT 109.570 197.110 109.890 197.170 ;
        RECT 111.885 197.110 112.175 197.155 ;
        RECT 112.880 197.110 113.020 197.310 ;
        RECT 115.550 197.250 115.870 197.310 ;
        RECT 121.530 197.450 121.850 197.510 ;
        RECT 122.925 197.450 123.215 197.495 ;
        RECT 125.760 197.450 125.900 197.590 ;
        RECT 121.530 197.310 123.215 197.450 ;
        RECT 121.530 197.250 121.850 197.310 ;
        RECT 122.925 197.265 123.215 197.310 ;
        RECT 123.460 197.310 125.900 197.450 ;
        RECT 109.570 196.970 113.020 197.110 ;
        RECT 109.570 196.910 109.890 196.970 ;
        RECT 111.885 196.925 112.175 196.970 ;
        RECT 113.250 196.910 113.570 197.170 ;
        RECT 113.725 197.110 114.015 197.155 ;
        RECT 116.010 197.110 116.330 197.170 ;
        RECT 113.725 196.970 116.330 197.110 ;
        RECT 113.725 196.925 114.015 196.970 ;
        RECT 116.010 196.910 116.330 196.970 ;
        RECT 122.450 196.910 122.770 197.170 ;
        RECT 123.460 197.125 123.600 197.310 ;
        RECT 123.845 197.125 124.135 197.155 ;
        RECT 123.460 196.985 124.135 197.125 ;
        RECT 125.225 197.110 125.515 197.155 ;
        RECT 123.845 196.925 124.135 196.985 ;
        RECT 124.380 196.970 125.515 197.110 ;
        RECT 104.510 196.630 107.500 196.770 ;
        RECT 107.730 196.770 108.050 196.830 ;
        RECT 110.490 196.770 110.810 196.830 ;
        RECT 110.965 196.770 111.255 196.815 ;
        RECT 107.730 196.630 109.800 196.770 ;
        RECT 100.830 196.430 101.150 196.490 ;
        RECT 102.225 196.430 102.515 196.475 ;
        RECT 95.400 196.290 102.515 196.430 ;
        RECT 43.330 196.230 43.650 196.290 ;
        RECT 50.230 196.230 50.550 196.290 ;
        RECT 41.030 196.090 41.350 196.150 ;
        RECT 42.885 196.090 43.175 196.135 ;
        RECT 41.030 195.950 43.175 196.090 ;
        RECT 41.030 195.890 41.350 195.950 ;
        RECT 42.885 195.905 43.175 195.950 ;
        RECT 49.325 196.090 49.615 196.135 ;
        RECT 49.770 196.090 50.090 196.150 ;
        RECT 49.325 195.950 50.090 196.090 ;
        RECT 49.325 195.905 49.615 195.950 ;
        RECT 49.770 195.890 50.090 195.950 ;
        RECT 51.150 196.090 51.470 196.150 ;
        RECT 52.545 196.090 52.835 196.135 ;
        RECT 51.150 195.950 52.835 196.090 ;
        RECT 51.150 195.890 51.470 195.950 ;
        RECT 52.545 195.905 52.835 195.950 ;
        RECT 65.410 195.890 65.730 196.150 ;
        RECT 65.960 196.090 66.100 196.290 ;
        RECT 69.090 196.230 69.410 196.290 ;
        RECT 94.390 196.230 94.710 196.290 ;
        RECT 100.830 196.230 101.150 196.290 ;
        RECT 102.225 196.245 102.515 196.290 ;
        RECT 66.330 196.090 66.650 196.150 ;
        RECT 65.960 195.950 66.650 196.090 ;
        RECT 66.330 195.890 66.650 195.950 ;
        RECT 66.790 196.090 67.110 196.150 ;
        RECT 70.930 196.090 71.250 196.150 ;
        RECT 80.130 196.090 80.450 196.150 ;
        RECT 66.790 195.950 80.450 196.090 ;
        RECT 66.790 195.890 67.110 195.950 ;
        RECT 70.930 195.890 71.250 195.950 ;
        RECT 80.130 195.890 80.450 195.950 ;
        RECT 82.445 196.090 82.735 196.135 ;
        RECT 83.350 196.090 83.670 196.150 ;
        RECT 82.445 195.950 83.670 196.090 ;
        RECT 82.445 195.905 82.735 195.950 ;
        RECT 83.350 195.890 83.670 195.950 ;
        RECT 92.565 196.090 92.855 196.135 ;
        RECT 93.930 196.090 94.250 196.150 ;
        RECT 92.565 195.950 94.250 196.090 ;
        RECT 92.565 195.905 92.855 195.950 ;
        RECT 93.930 195.890 94.250 195.950 ;
        RECT 99.910 196.090 100.230 196.150 ;
        RECT 104.140 196.090 104.280 196.585 ;
        RECT 104.510 196.570 104.830 196.630 ;
        RECT 107.730 196.570 108.050 196.630 ;
        RECT 105.445 196.430 105.735 196.475 ;
        RECT 109.110 196.430 109.430 196.490 ;
        RECT 105.445 196.290 109.430 196.430 ;
        RECT 109.660 196.430 109.800 196.630 ;
        RECT 110.490 196.630 111.255 196.770 ;
        RECT 110.490 196.570 110.810 196.630 ;
        RECT 110.965 196.585 111.255 196.630 ;
        RECT 111.425 196.585 111.715 196.815 ;
        RECT 111.500 196.430 111.640 196.585 ;
        RECT 112.330 196.570 112.650 196.830 ;
        RECT 116.470 196.770 116.790 196.830 ;
        RECT 124.380 196.770 124.520 196.970 ;
        RECT 125.225 196.925 125.515 196.970 ;
        RECT 116.470 196.630 124.520 196.770 ;
        RECT 116.470 196.570 116.790 196.630 ;
        RECT 124.765 196.585 125.055 196.815 ;
        RECT 125.300 196.770 125.440 196.925 ;
        RECT 125.670 196.910 125.990 197.170 ;
        RECT 126.605 197.125 126.895 197.155 ;
        RECT 127.140 197.125 127.280 197.650 ;
        RECT 128.430 197.250 128.750 197.510 ;
        RECT 128.940 197.450 129.080 197.650 ;
        RECT 129.810 197.650 131.495 197.790 ;
        RECT 129.810 197.590 130.130 197.650 ;
        RECT 131.205 197.605 131.495 197.650 ;
        RECT 132.110 197.790 132.430 197.850 ;
        RECT 135.345 197.790 135.635 197.835 ;
        RECT 132.110 197.650 135.635 197.790 ;
        RECT 132.110 197.590 132.430 197.650 ;
        RECT 135.345 197.605 135.635 197.650 ;
        RECT 137.170 197.450 137.490 197.510 ;
        RECT 128.940 197.310 131.420 197.450 ;
        RECT 131.280 197.170 131.420 197.310 ;
        RECT 132.200 197.310 137.490 197.450 ;
        RECT 126.605 196.985 127.280 197.125 ;
        RECT 126.605 196.925 126.895 196.985 ;
        RECT 127.970 196.910 128.290 197.170 ;
        RECT 128.905 196.925 129.195 197.155 ;
        RECT 127.510 196.770 127.830 196.830 ;
        RECT 125.300 196.630 127.830 196.770 ;
        RECT 109.660 196.290 111.640 196.430 ;
        RECT 105.445 196.245 105.735 196.290 ;
        RECT 109.110 196.230 109.430 196.290 ;
        RECT 99.910 195.950 104.280 196.090 ;
        RECT 119.230 196.090 119.550 196.150 ;
        RECT 124.840 196.090 124.980 196.585 ;
        RECT 127.510 196.570 127.830 196.630 ;
        RECT 128.430 196.770 128.750 196.830 ;
        RECT 128.980 196.770 129.120 196.925 ;
        RECT 129.810 196.910 130.130 197.170 ;
        RECT 131.190 196.910 131.510 197.170 ;
        RECT 132.200 197.155 132.340 197.310 ;
        RECT 137.170 197.250 137.490 197.310 ;
        RECT 132.125 196.925 132.415 197.155 ;
        RECT 132.570 196.910 132.890 197.170 ;
        RECT 133.490 196.910 133.810 197.170 ;
        RECT 133.965 196.925 134.255 197.155 ;
        RECT 128.430 196.630 129.120 196.770 ;
        RECT 129.350 196.770 129.670 196.830 ;
        RECT 134.040 196.770 134.180 196.925 ;
        RECT 129.350 196.630 134.180 196.770 ;
        RECT 128.430 196.570 128.750 196.630 ;
        RECT 129.350 196.570 129.670 196.630 ;
        RECT 134.410 196.570 134.730 196.830 ;
        RECT 136.265 196.585 136.555 196.815 ;
        RECT 136.340 196.430 136.480 196.585 ;
        RECT 133.120 196.290 136.480 196.430 ;
        RECT 119.230 195.950 124.980 196.090 ;
        RECT 126.590 196.090 126.910 196.150 ;
        RECT 127.065 196.090 127.355 196.135 ;
        RECT 133.120 196.090 133.260 196.290 ;
        RECT 126.590 195.950 133.260 196.090 ;
        RECT 134.870 196.090 135.190 196.150 ;
        RECT 135.790 196.090 136.110 196.150 ;
        RECT 136.265 196.090 136.555 196.135 ;
        RECT 134.870 195.950 136.555 196.090 ;
        RECT 99.910 195.890 100.230 195.950 ;
        RECT 119.230 195.890 119.550 195.950 ;
        RECT 126.590 195.890 126.910 195.950 ;
        RECT 127.065 195.905 127.355 195.950 ;
        RECT 134.870 195.890 135.190 195.950 ;
        RECT 135.790 195.890 136.110 195.950 ;
        RECT 136.265 195.905 136.555 195.950 ;
        RECT 27.160 195.270 139.860 195.750 ;
        RECT 41.030 194.870 41.350 195.130 ;
        RECT 43.345 195.070 43.635 195.115 ;
        RECT 44.710 195.070 45.030 195.130 ;
        RECT 43.345 194.930 45.030 195.070 ;
        RECT 43.345 194.885 43.635 194.930 ;
        RECT 44.710 194.870 45.030 194.930 ;
        RECT 53.005 195.070 53.295 195.115 ;
        RECT 54.370 195.070 54.690 195.130 ;
        RECT 53.005 194.930 54.690 195.070 ;
        RECT 53.005 194.885 53.295 194.930 ;
        RECT 54.370 194.870 54.690 194.930 ;
        RECT 54.830 195.070 55.150 195.130 ;
        RECT 63.110 195.070 63.430 195.130 ;
        RECT 54.830 194.930 63.430 195.070 ;
        RECT 54.830 194.870 55.150 194.930 ;
        RECT 63.110 194.870 63.430 194.930 ;
        RECT 65.410 195.070 65.730 195.130 ;
        RECT 66.345 195.070 66.635 195.115 ;
        RECT 65.410 194.930 66.635 195.070 ;
        RECT 65.410 194.870 65.730 194.930 ;
        RECT 66.345 194.885 66.635 194.930 ;
        RECT 70.010 194.870 70.330 195.130 ;
        RECT 70.930 195.070 71.250 195.130 ;
        RECT 70.930 194.930 72.080 195.070 ;
        RECT 70.930 194.870 71.250 194.930 ;
        RECT 43.805 194.730 44.095 194.775 ;
        RECT 45.170 194.730 45.490 194.790 ;
        RECT 43.805 194.590 45.490 194.730 ;
        RECT 43.805 194.545 44.095 194.590 ;
        RECT 45.170 194.530 45.490 194.590 ;
        RECT 48.865 194.730 49.155 194.775 ;
        RECT 62.650 194.730 62.970 194.790 ;
        RECT 48.865 194.590 62.970 194.730 ;
        RECT 63.200 194.730 63.340 194.870 ;
        RECT 66.790 194.730 67.110 194.790 ;
        RECT 68.170 194.730 68.490 194.790 ;
        RECT 63.200 194.590 67.110 194.730 ;
        RECT 48.865 194.545 49.155 194.590 ;
        RECT 62.650 194.530 62.970 194.590 ;
        RECT 66.790 194.530 67.110 194.590 ;
        RECT 67.340 194.590 68.490 194.730 ;
        RECT 39.650 194.390 39.970 194.450 ;
        RECT 49.310 194.390 49.630 194.450 ;
        RECT 39.650 194.250 42.180 194.390 ;
        RECT 39.650 194.190 39.970 194.250 ;
        RECT 30.005 194.050 30.295 194.095 ;
        RECT 31.370 194.050 31.690 194.110 ;
        RECT 30.005 193.910 31.690 194.050 ;
        RECT 30.005 193.865 30.295 193.910 ;
        RECT 31.370 193.850 31.690 193.910 ;
        RECT 38.270 194.050 38.590 194.110 ;
        RECT 42.040 194.095 42.180 194.250 ;
        RECT 45.255 194.250 49.630 194.390 ;
        RECT 40.585 194.050 40.875 194.095 ;
        RECT 38.270 193.910 40.875 194.050 ;
        RECT 38.270 193.850 38.590 193.910 ;
        RECT 40.585 193.865 40.875 193.910 ;
        RECT 41.965 193.865 42.255 194.095 ;
        RECT 42.410 193.850 42.730 194.110 ;
        RECT 45.255 194.095 45.395 194.250 ;
        RECT 49.310 194.190 49.630 194.250 ;
        RECT 54.845 194.390 55.135 194.435 ;
        RECT 57.590 194.390 57.910 194.450 ;
        RECT 54.845 194.250 57.910 194.390 ;
        RECT 54.845 194.205 55.135 194.250 ;
        RECT 57.590 194.190 57.910 194.250 ;
        RECT 59.445 194.390 59.735 194.435 ;
        RECT 62.190 194.390 62.510 194.450 ;
        RECT 67.340 194.435 67.480 194.590 ;
        RECT 68.170 194.530 68.490 194.590 ;
        RECT 69.090 194.730 69.410 194.790 ;
        RECT 70.470 194.730 70.790 194.790 ;
        RECT 69.090 194.590 69.780 194.730 ;
        RECT 69.090 194.530 69.410 194.590 ;
        RECT 69.640 194.435 69.780 194.590 ;
        RECT 70.470 194.530 70.930 194.730 ;
        RECT 59.445 194.250 62.510 194.390 ;
        RECT 59.445 194.205 59.735 194.250 ;
        RECT 62.190 194.190 62.510 194.250 ;
        RECT 67.265 194.205 67.555 194.435 ;
        RECT 69.565 194.205 69.855 194.435 ;
        RECT 45.180 193.865 45.470 194.095 ;
        RECT 45.645 194.050 45.935 194.095 ;
        RECT 46.090 194.050 46.410 194.110 ;
        RECT 45.645 193.910 46.410 194.050 ;
        RECT 45.645 193.865 45.935 193.910 ;
        RECT 44.250 193.710 44.570 193.770 ;
        RECT 45.720 193.710 45.860 193.865 ;
        RECT 46.090 193.850 46.410 193.910 ;
        RECT 47.485 194.050 47.775 194.095 ;
        RECT 47.930 194.050 48.250 194.110 ;
        RECT 47.485 193.910 48.250 194.050 ;
        RECT 47.485 193.865 47.775 193.910 ;
        RECT 47.930 193.850 48.250 193.910 ;
        RECT 48.850 193.850 49.170 194.110 ;
        RECT 53.925 193.865 54.215 194.095 ;
        RECT 44.250 193.570 45.860 193.710 ;
        RECT 54.000 193.710 54.140 193.865 ;
        RECT 54.370 193.850 54.690 194.110 ;
        RECT 55.305 193.865 55.595 194.095 ;
        RECT 56.225 194.050 56.515 194.095 ;
        RECT 57.130 194.050 57.450 194.110 ;
        RECT 56.225 193.910 57.450 194.050 ;
        RECT 56.225 193.865 56.515 193.910 ;
        RECT 55.380 193.710 55.520 193.865 ;
        RECT 57.130 193.850 57.450 193.910 ;
        RECT 58.050 193.850 58.370 194.110 ;
        RECT 58.525 194.050 58.815 194.095 ;
        RECT 62.650 194.050 62.970 194.110 ;
        RECT 67.725 194.050 68.015 194.095 ;
        RECT 68.630 194.050 68.950 194.110 ;
        RECT 70.790 194.095 70.930 194.530 ;
        RECT 71.940 194.390 72.080 194.930 ;
        RECT 80.590 194.870 80.910 195.130 ;
        RECT 85.190 195.070 85.510 195.130 ;
        RECT 98.990 195.070 99.310 195.130 ;
        RECT 120.610 195.070 120.930 195.130 ;
        RECT 85.190 194.930 99.310 195.070 ;
        RECT 85.190 194.870 85.510 194.930 ;
        RECT 98.990 194.870 99.310 194.930 ;
        RECT 102.300 194.930 120.930 195.070 ;
        RECT 73.230 194.730 73.550 194.790 ;
        RECT 73.705 194.730 73.995 194.775 ;
        RECT 73.230 194.590 73.995 194.730 ;
        RECT 73.230 194.530 73.550 194.590 ;
        RECT 73.705 194.545 73.995 194.590 ;
        RECT 75.160 194.590 89.560 194.730 ;
        RECT 74.150 194.390 74.470 194.450 ;
        RECT 71.495 194.250 72.080 194.390 ;
        RECT 72.855 194.250 74.470 194.390 ;
        RECT 71.495 194.095 71.635 194.250 ;
        RECT 58.525 193.910 66.100 194.050 ;
        RECT 58.525 193.865 58.815 193.910 ;
        RECT 62.650 193.850 62.970 193.910 ;
        RECT 56.670 193.710 56.990 193.770 ;
        RECT 59.445 193.710 59.735 193.755 ;
        RECT 54.000 193.570 55.060 193.710 ;
        RECT 55.380 193.570 59.735 193.710 ;
        RECT 44.250 193.510 44.570 193.570 ;
        RECT 54.920 193.430 55.060 193.570 ;
        RECT 56.670 193.510 56.990 193.570 ;
        RECT 59.445 193.525 59.735 193.570 ;
        RECT 59.890 193.710 60.210 193.770 ;
        RECT 63.125 193.710 63.415 193.755 ;
        RECT 59.890 193.570 63.415 193.710 ;
        RECT 59.890 193.510 60.210 193.570 ;
        RECT 63.125 193.525 63.415 193.570 ;
        RECT 64.030 193.510 64.350 193.770 ;
        RECT 25.390 193.370 25.710 193.430 ;
        RECT 29.085 193.370 29.375 193.415 ;
        RECT 25.390 193.230 29.375 193.370 ;
        RECT 25.390 193.170 25.710 193.230 ;
        RECT 29.085 193.185 29.375 193.230 ;
        RECT 47.945 193.370 48.235 193.415 ;
        RECT 52.070 193.370 52.390 193.430 ;
        RECT 47.945 193.230 52.390 193.370 ;
        RECT 47.945 193.185 48.235 193.230 ;
        RECT 52.070 193.170 52.390 193.230 ;
        RECT 54.830 193.170 55.150 193.430 ;
        RECT 65.960 193.370 66.100 193.910 ;
        RECT 67.725 193.910 68.950 194.050 ;
        RECT 67.725 193.865 68.015 193.910 ;
        RECT 68.630 193.850 68.950 193.910 ;
        RECT 70.725 193.865 71.015 194.095 ;
        RECT 71.405 193.865 71.695 194.095 ;
        RECT 71.865 194.050 72.155 194.095 ;
        RECT 72.310 194.050 72.630 194.110 ;
        RECT 72.855 194.095 72.995 194.250 ;
        RECT 74.150 194.190 74.470 194.250 ;
        RECT 71.865 193.910 72.630 194.050 ;
        RECT 71.865 193.865 72.155 193.910 ;
        RECT 72.310 193.850 72.630 193.910 ;
        RECT 72.780 193.865 73.070 194.095 ;
        RECT 73.230 194.050 73.550 194.110 ;
        RECT 75.160 194.095 75.300 194.590 ;
        RECT 76.910 194.390 77.230 194.450 ;
        RECT 76.910 194.250 80.820 194.390 ;
        RECT 76.910 194.190 77.230 194.250 ;
        RECT 73.705 194.050 73.995 194.095 ;
        RECT 75.085 194.050 75.375 194.095 ;
        RECT 79.685 194.050 79.975 194.095 ;
        RECT 73.230 193.910 73.995 194.050 ;
        RECT 66.330 193.710 66.650 193.770 ;
        RECT 69.105 193.710 69.395 193.755 ;
        RECT 72.855 193.710 72.995 193.865 ;
        RECT 73.230 193.850 73.550 193.910 ;
        RECT 73.705 193.865 73.995 193.910 ;
        RECT 74.240 193.910 75.375 194.050 ;
        RECT 66.330 193.570 72.995 193.710 ;
        RECT 66.330 193.510 66.650 193.570 ;
        RECT 69.105 193.525 69.395 193.570 ;
        RECT 74.240 193.370 74.380 193.910 ;
        RECT 75.085 193.865 75.375 193.910 ;
        RECT 78.840 193.910 79.975 194.050 ;
        RECT 78.840 193.430 78.980 193.910 ;
        RECT 79.685 193.865 79.975 193.910 ;
        RECT 80.130 193.850 80.450 194.110 ;
        RECT 80.680 194.050 80.820 194.250 ;
        RECT 81.050 194.190 81.370 194.450 ;
        RECT 84.730 194.390 85.050 194.450 ;
        RECT 89.420 194.390 89.560 194.590 ;
        RECT 89.790 194.530 90.110 194.790 ;
        RECT 93.930 194.730 94.250 194.790 ;
        RECT 102.300 194.730 102.440 194.930 ;
        RECT 120.610 194.870 120.930 194.930 ;
        RECT 121.530 195.070 121.850 195.130 ;
        RECT 124.305 195.070 124.595 195.115 ;
        RECT 125.210 195.070 125.530 195.130 ;
        RECT 121.530 194.930 125.530 195.070 ;
        RECT 121.530 194.870 121.850 194.930 ;
        RECT 124.305 194.885 124.595 194.930 ;
        RECT 125.210 194.870 125.530 194.930 ;
        RECT 126.130 195.070 126.450 195.130 ;
        RECT 133.505 195.070 133.795 195.115 ;
        RECT 126.130 194.930 133.795 195.070 ;
        RECT 126.130 194.870 126.450 194.930 ;
        RECT 133.505 194.885 133.795 194.930 ;
        RECT 137.630 194.870 137.950 195.130 ;
        RECT 93.930 194.590 102.440 194.730 ;
        RECT 102.670 194.730 102.990 194.790 ;
        RECT 112.790 194.730 113.110 194.790 ;
        RECT 123.370 194.730 123.690 194.790 ;
        RECT 129.350 194.730 129.670 194.790 ;
        RECT 102.670 194.590 113.110 194.730 ;
        RECT 93.930 194.530 94.250 194.590 ;
        RECT 102.670 194.530 102.990 194.590 ;
        RECT 112.790 194.530 113.110 194.590 ;
        RECT 118.170 194.590 129.670 194.730 ;
        RECT 91.170 194.390 91.490 194.450 ;
        RECT 82.520 194.250 86.800 194.390 ;
        RECT 89.420 194.250 91.490 194.390 ;
        RECT 82.520 194.095 82.660 194.250 ;
        RECT 84.730 194.190 85.050 194.250 ;
        RECT 82.445 194.050 82.735 194.095 ;
        RECT 83.350 194.050 83.670 194.110 ;
        RECT 80.680 193.910 82.735 194.050 ;
        RECT 83.155 193.910 83.670 194.050 ;
        RECT 82.445 193.865 82.735 193.910 ;
        RECT 83.350 193.850 83.670 193.910 ;
        RECT 83.810 193.850 84.130 194.110 ;
        RECT 84.285 193.865 84.575 194.095 ;
        RECT 81.970 193.710 82.290 193.770 ;
        RECT 84.360 193.710 84.500 193.865 ;
        RECT 85.190 193.850 85.510 194.110 ;
        RECT 86.660 194.095 86.800 194.250 ;
        RECT 91.170 194.190 91.490 194.250 ;
        RECT 91.630 194.390 91.950 194.450 ;
        RECT 92.105 194.390 92.395 194.435 ;
        RECT 91.630 194.250 92.395 194.390 ;
        RECT 91.630 194.190 91.950 194.250 ;
        RECT 92.105 194.205 92.395 194.250 ;
        RECT 93.010 194.390 93.330 194.450 ;
        RECT 98.070 194.390 98.390 194.450 ;
        RECT 93.010 194.250 98.390 194.390 ;
        RECT 93.010 194.190 93.330 194.250 ;
        RECT 98.070 194.190 98.390 194.250 ;
        RECT 101.290 194.390 101.610 194.450 ;
        RECT 105.890 194.390 106.210 194.450 ;
        RECT 101.290 194.250 106.210 194.390 ;
        RECT 101.290 194.190 101.610 194.250 ;
        RECT 105.890 194.190 106.210 194.250 ;
        RECT 106.350 194.390 106.670 194.450 ;
        RECT 110.950 194.390 111.270 194.450 ;
        RECT 118.170 194.390 118.310 194.590 ;
        RECT 123.370 194.530 123.690 194.590 ;
        RECT 129.350 194.530 129.670 194.590 ;
        RECT 106.350 194.250 118.310 194.390 ;
        RECT 122.450 194.390 122.770 194.450 ;
        RECT 132.570 194.390 132.890 194.450 ;
        RECT 122.450 194.250 132.890 194.390 ;
        RECT 106.350 194.190 106.670 194.250 ;
        RECT 110.950 194.190 111.270 194.250 ;
        RECT 122.450 194.190 122.770 194.250 ;
        RECT 132.570 194.190 132.890 194.250 ;
        RECT 86.585 193.865 86.875 194.095 ;
        RECT 87.510 193.865 87.800 194.095 ;
        RECT 81.970 193.570 84.500 193.710 ;
        RECT 87.580 193.710 87.720 193.865 ;
        RECT 87.950 193.850 88.270 194.110 ;
        RECT 88.410 194.050 88.730 194.110 ;
        RECT 99.450 194.050 99.770 194.110 ;
        RECT 103.590 194.050 103.910 194.110 ;
        RECT 88.410 193.910 103.910 194.050 ;
        RECT 88.410 193.850 88.730 193.910 ;
        RECT 99.450 193.850 99.770 193.910 ;
        RECT 103.590 193.850 103.910 193.910 ;
        RECT 104.065 194.050 104.355 194.095 ;
        RECT 107.270 194.050 107.590 194.110 ;
        RECT 104.065 193.910 107.590 194.050 ;
        RECT 104.065 193.865 104.355 193.910 ;
        RECT 107.270 193.850 107.590 193.910 ;
        RECT 116.945 194.050 117.235 194.095 ;
        RECT 118.770 194.050 119.090 194.110 ;
        RECT 116.945 193.910 119.090 194.050 ;
        RECT 116.945 193.865 117.235 193.910 ;
        RECT 118.770 193.850 119.090 193.910 ;
        RECT 120.610 194.050 120.930 194.110 ;
        RECT 131.190 194.050 131.510 194.110 ;
        RECT 136.725 194.050 137.015 194.095 ;
        RECT 120.610 193.910 127.735 194.050 ;
        RECT 120.610 193.850 120.930 193.910 ;
        RECT 89.790 193.710 90.110 193.770 ;
        RECT 87.580 193.570 90.110 193.710 ;
        RECT 81.970 193.510 82.290 193.570 ;
        RECT 89.790 193.510 90.110 193.570 ;
        RECT 91.170 193.710 91.490 193.770 ;
        RECT 98.990 193.710 99.310 193.770 ;
        RECT 91.170 193.570 99.310 193.710 ;
        RECT 91.170 193.510 91.490 193.570 ;
        RECT 98.990 193.510 99.310 193.570 ;
        RECT 100.370 193.710 100.690 193.770 ;
        RECT 100.845 193.710 101.135 193.755 ;
        RECT 100.370 193.570 101.135 193.710 ;
        RECT 100.370 193.510 100.690 193.570 ;
        RECT 100.845 193.525 101.135 193.570 ;
        RECT 101.750 193.710 102.070 193.770 ;
        RECT 105.905 193.710 106.195 193.755 ;
        RECT 101.750 193.570 106.195 193.710 ;
        RECT 101.750 193.510 102.070 193.570 ;
        RECT 105.905 193.525 106.195 193.570 ;
        RECT 107.745 193.525 108.035 193.755 ;
        RECT 65.960 193.230 74.380 193.370 ;
        RECT 74.625 193.370 74.915 193.415 ;
        RECT 78.750 193.370 79.070 193.430 ;
        RECT 74.625 193.230 79.070 193.370 ;
        RECT 74.625 193.185 74.915 193.230 ;
        RECT 78.750 193.170 79.070 193.230 ;
        RECT 85.665 193.370 85.955 193.415 ;
        RECT 86.110 193.370 86.430 193.430 ;
        RECT 85.665 193.230 86.430 193.370 ;
        RECT 85.665 193.185 85.955 193.230 ;
        RECT 86.110 193.170 86.430 193.230 ;
        RECT 86.570 193.370 86.890 193.430 ;
        RECT 95.310 193.370 95.630 193.430 ;
        RECT 86.570 193.230 95.630 193.370 ;
        RECT 86.570 193.170 86.890 193.230 ;
        RECT 95.310 193.170 95.630 193.230 ;
        RECT 105.430 193.170 105.750 193.430 ;
        RECT 106.350 193.170 106.670 193.430 ;
        RECT 106.810 193.170 107.130 193.430 ;
        RECT 107.820 193.370 107.960 193.525 ;
        RECT 108.190 193.510 108.510 193.770 ;
        RECT 117.850 193.510 118.170 193.770 ;
        RECT 121.990 193.710 122.310 193.770 ;
        RECT 127.065 193.710 127.355 193.755 ;
        RECT 121.990 193.570 127.355 193.710 ;
        RECT 127.595 193.710 127.735 193.910 ;
        RECT 131.190 193.910 137.015 194.050 ;
        RECT 131.190 193.850 131.510 193.910 ;
        RECT 136.725 193.865 137.015 193.910 ;
        RECT 136.250 193.710 136.570 193.770 ;
        RECT 127.595 193.570 136.570 193.710 ;
        RECT 121.990 193.510 122.310 193.570 ;
        RECT 127.065 193.525 127.355 193.570 ;
        RECT 136.250 193.510 136.570 193.570 ;
        RECT 122.910 193.370 123.230 193.430 ;
        RECT 107.820 193.230 123.230 193.370 ;
        RECT 122.910 193.170 123.230 193.230 ;
        RECT 128.430 193.370 128.750 193.430 ;
        RECT 131.190 193.370 131.510 193.430 ;
        RECT 128.430 193.230 131.510 193.370 ;
        RECT 128.430 193.170 128.750 193.230 ;
        RECT 131.190 193.170 131.510 193.230 ;
        RECT 27.160 192.550 139.860 193.030 ;
        RECT 31.370 192.150 31.690 192.410 ;
        RECT 53.910 192.150 54.230 192.410 ;
        RECT 57.145 192.350 57.435 192.395 ;
        RECT 57.590 192.350 57.910 192.410 ;
        RECT 57.145 192.210 57.910 192.350 ;
        RECT 57.145 192.165 57.435 192.210 ;
        RECT 57.590 192.150 57.910 192.210 ;
        RECT 58.510 192.350 58.830 192.410 ;
        RECT 64.950 192.350 65.270 192.410 ;
        RECT 66.345 192.350 66.635 192.395 ;
        RECT 58.510 192.210 61.960 192.350 ;
        RECT 58.510 192.150 58.830 192.210 ;
        RECT 43.345 192.010 43.635 192.055 ;
        RECT 45.630 192.010 45.950 192.070 ;
        RECT 48.390 192.010 48.710 192.070 ;
        RECT 43.345 191.870 48.710 192.010 ;
        RECT 43.345 191.825 43.635 191.870 ;
        RECT 45.630 191.810 45.950 191.870 ;
        RECT 48.390 191.810 48.710 191.870 ;
        RECT 51.150 191.810 51.470 192.070 ;
        RECT 52.990 192.010 53.310 192.070 ;
        RECT 51.700 191.870 53.310 192.010 ;
        RECT 25.390 191.670 25.710 191.730 ;
        RECT 29.085 191.670 29.375 191.715 ;
        RECT 25.390 191.530 29.375 191.670 ;
        RECT 25.390 191.470 25.710 191.530 ;
        RECT 29.085 191.485 29.375 191.530 ;
        RECT 32.290 191.470 32.610 191.730 ;
        RECT 40.110 191.470 40.430 191.730 ;
        RECT 41.030 191.470 41.350 191.730 ;
        RECT 42.885 191.485 43.175 191.715 ;
        RECT 29.990 191.130 30.310 191.390 ;
        RECT 37.810 191.330 38.130 191.390 ;
        RECT 42.960 191.330 43.100 191.485 ;
        RECT 49.310 191.470 49.630 191.730 ;
        RECT 49.785 191.670 50.075 191.715 ;
        RECT 50.705 191.670 50.995 191.715 ;
        RECT 51.700 191.670 51.840 191.870 ;
        RECT 52.990 191.810 53.310 191.870 ;
        RECT 58.140 191.870 61.500 192.010 ;
        RECT 49.785 191.530 50.460 191.670 ;
        RECT 49.785 191.485 50.075 191.530 ;
        RECT 48.390 191.330 48.710 191.390 ;
        RECT 37.810 191.190 48.710 191.330 ;
        RECT 37.810 191.130 38.130 191.190 ;
        RECT 48.390 191.130 48.710 191.190 ;
        RECT 41.045 190.990 41.335 191.035 ;
        RECT 44.250 190.990 44.570 191.050 ;
        RECT 41.045 190.850 44.570 190.990 ;
        RECT 41.045 190.805 41.335 190.850 ;
        RECT 44.250 190.790 44.570 190.850 ;
        RECT 50.320 190.650 50.460 191.530 ;
        RECT 50.705 191.530 51.840 191.670 ;
        RECT 50.705 191.485 50.995 191.530 ;
        RECT 52.070 191.470 52.390 191.730 ;
        RECT 52.530 191.470 52.850 191.730 ;
        RECT 54.830 191.470 55.150 191.730 ;
        RECT 55.305 191.670 55.595 191.715 ;
        RECT 56.210 191.670 56.530 191.730 ;
        RECT 55.305 191.530 56.530 191.670 ;
        RECT 55.305 191.485 55.595 191.530 ;
        RECT 56.210 191.470 56.530 191.530 ;
        RECT 56.670 191.470 56.990 191.730 ;
        RECT 58.140 191.715 58.280 191.870 ;
        RECT 58.065 191.485 58.355 191.715 ;
        RECT 58.510 191.470 58.830 191.730 ;
        RECT 59.445 191.485 59.735 191.715 ;
        RECT 59.890 191.670 60.210 191.730 ;
        RECT 60.365 191.670 60.655 191.715 ;
        RECT 59.890 191.530 60.655 191.670 ;
        RECT 51.525 191.330 51.815 191.375 ;
        RECT 58.600 191.330 58.740 191.470 ;
        RECT 51.525 191.190 58.740 191.330 ;
        RECT 51.525 191.145 51.815 191.190 ;
        RECT 58.985 191.145 59.275 191.375 ;
        RECT 50.705 190.990 50.995 191.035 ;
        RECT 56.225 190.990 56.515 191.035 ;
        RECT 50.705 190.850 56.515 190.990 ;
        RECT 50.705 190.805 50.995 190.850 ;
        RECT 56.225 190.805 56.515 190.850 ;
        RECT 58.050 190.990 58.370 191.050 ;
        RECT 59.060 190.990 59.200 191.145 ;
        RECT 58.050 190.850 59.200 190.990 ;
        RECT 59.520 190.990 59.660 191.485 ;
        RECT 59.890 191.470 60.210 191.530 ;
        RECT 60.365 191.485 60.655 191.530 ;
        RECT 61.360 191.330 61.500 191.870 ;
        RECT 61.820 191.670 61.960 192.210 ;
        RECT 64.950 192.210 66.635 192.350 ;
        RECT 64.950 192.150 65.270 192.210 ;
        RECT 66.345 192.165 66.635 192.210 ;
        RECT 67.710 192.150 68.030 192.410 ;
        RECT 68.170 192.150 68.490 192.410 ;
        RECT 71.865 192.350 72.155 192.395 ;
        RECT 81.050 192.350 81.370 192.410 ;
        RECT 71.865 192.210 81.370 192.350 ;
        RECT 71.865 192.165 72.155 192.210 ;
        RECT 81.050 192.150 81.370 192.210 ;
        RECT 86.110 192.150 86.430 192.410 ;
        RECT 87.965 192.350 88.255 192.395 ;
        RECT 89.790 192.350 90.110 192.410 ;
        RECT 87.965 192.210 90.110 192.350 ;
        RECT 87.965 192.165 88.255 192.210 ;
        RECT 89.790 192.150 90.110 192.210 ;
        RECT 92.090 192.150 92.410 192.410 ;
        RECT 92.550 192.150 92.870 192.410 ;
        RECT 94.850 192.150 95.170 192.410 ;
        RECT 95.310 192.350 95.630 192.410 ;
        RECT 105.445 192.350 105.735 192.395 ;
        RECT 95.310 192.210 105.735 192.350 ;
        RECT 95.310 192.150 95.630 192.210 ;
        RECT 105.445 192.165 105.735 192.210 ;
        RECT 105.890 192.150 106.210 192.410 ;
        RECT 107.730 192.150 108.050 192.410 ;
        RECT 121.070 192.350 121.390 192.410 ;
        RECT 132.570 192.350 132.890 192.410 ;
        RECT 134.425 192.350 134.715 192.395 ;
        RECT 121.070 192.210 131.880 192.350 ;
        RECT 121.070 192.150 121.390 192.210 ;
        RECT 67.250 191.810 67.570 192.070 ;
        RECT 70.930 192.010 71.250 192.070 ;
        RECT 75.070 192.010 75.390 192.070 ;
        RECT 70.930 191.870 75.390 192.010 ;
        RECT 70.930 191.810 71.250 191.870 ;
        RECT 75.070 191.810 75.390 191.870 ;
        RECT 84.745 192.010 85.035 192.055 ;
        RECT 86.200 192.010 86.340 192.150 ;
        RECT 84.745 191.870 86.340 192.010 ;
        RECT 92.640 192.010 92.780 192.150 ;
        RECT 94.940 192.010 95.080 192.150 ;
        RECT 97.165 192.010 97.455 192.055 ;
        RECT 92.640 191.870 94.750 192.010 ;
        RECT 94.940 191.870 97.455 192.010 ;
        RECT 84.745 191.825 85.035 191.870 ;
        RECT 82.905 191.670 83.195 191.715 ;
        RECT 61.820 191.530 83.195 191.670 ;
        RECT 82.905 191.485 83.195 191.530 ;
        RECT 85.190 191.470 85.510 191.730 ;
        RECT 86.110 191.670 86.430 191.730 ;
        RECT 85.740 191.530 86.430 191.670 ;
        RECT 64.030 191.330 64.350 191.390 ;
        RECT 68.170 191.330 68.490 191.390 ;
        RECT 69.565 191.330 69.855 191.375 ;
        RECT 61.360 191.190 69.855 191.330 ;
        RECT 64.030 191.130 64.350 191.190 ;
        RECT 68.170 191.130 68.490 191.190 ;
        RECT 69.565 191.145 69.855 191.190 ;
        RECT 70.010 191.330 70.330 191.390 ;
        RECT 85.740 191.375 85.880 191.530 ;
        RECT 86.110 191.470 86.430 191.530 ;
        RECT 86.570 191.470 86.890 191.730 ;
        RECT 87.030 191.470 87.350 191.730 ;
        RECT 91.185 191.670 91.475 191.715 ;
        RECT 91.630 191.670 91.950 191.730 ;
        RECT 91.185 191.530 91.950 191.670 ;
        RECT 91.185 191.485 91.475 191.530 ;
        RECT 91.630 191.470 91.950 191.530 ;
        RECT 93.470 191.470 93.790 191.730 ;
        RECT 93.930 191.470 94.250 191.730 ;
        RECT 94.610 191.715 94.750 191.870 ;
        RECT 97.165 191.825 97.455 191.870 ;
        RECT 99.005 192.010 99.295 192.055 ;
        RECT 105.980 192.010 106.120 192.150 ;
        RECT 99.005 191.870 106.120 192.010 ;
        RECT 112.330 192.010 112.650 192.070 ;
        RECT 115.565 192.010 115.855 192.055 ;
        RECT 127.970 192.010 128.290 192.070 ;
        RECT 112.330 191.870 115.855 192.010 ;
        RECT 99.005 191.825 99.295 191.870 ;
        RECT 94.610 191.530 95.030 191.715 ;
        RECT 94.740 191.485 95.030 191.530 ;
        RECT 96.245 191.485 96.535 191.715 ;
        RECT 81.985 191.330 82.275 191.375 ;
        RECT 70.010 191.190 82.275 191.330 ;
        RECT 70.010 191.130 70.330 191.190 ;
        RECT 81.985 191.145 82.275 191.190 ;
        RECT 85.665 191.145 85.955 191.375 ;
        RECT 96.320 191.330 96.460 191.485 ;
        RECT 96.690 191.470 97.010 191.730 ;
        RECT 87.120 191.190 96.460 191.330 ;
        RECT 62.650 190.990 62.970 191.050 ;
        RECT 69.090 190.990 69.410 191.050 ;
        RECT 70.945 190.990 71.235 191.035 ;
        RECT 59.520 190.850 63.110 190.990 ;
        RECT 58.050 190.790 58.370 190.850 ;
        RECT 62.650 190.790 63.110 190.850 ;
        RECT 69.090 190.850 71.235 190.990 ;
        RECT 69.090 190.790 69.410 190.850 ;
        RECT 70.945 190.805 71.235 190.850 ;
        RECT 51.150 190.650 51.470 190.710 ;
        RECT 50.320 190.510 51.470 190.650 ;
        RECT 51.150 190.450 51.470 190.510 ;
        RECT 54.370 190.650 54.690 190.710 ;
        RECT 59.905 190.650 60.195 190.695 ;
        RECT 54.370 190.510 60.195 190.650 ;
        RECT 62.970 190.650 63.110 190.790 ;
        RECT 63.570 190.650 63.890 190.710 ;
        RECT 62.970 190.510 63.890 190.650 ;
        RECT 54.370 190.450 54.690 190.510 ;
        RECT 59.905 190.465 60.195 190.510 ;
        RECT 63.570 190.450 63.890 190.510 ;
        RECT 70.470 190.650 70.790 190.710 ;
        RECT 73.690 190.650 74.010 190.710 ;
        RECT 80.130 190.650 80.450 190.710 ;
        RECT 70.470 190.510 80.450 190.650 ;
        RECT 82.060 190.650 82.200 191.145 ;
        RECT 87.120 191.050 87.260 191.190 ;
        RECT 83.350 190.790 83.670 191.050 ;
        RECT 83.810 190.990 84.130 191.050 ;
        RECT 86.570 190.990 86.890 191.050 ;
        RECT 83.810 190.850 86.890 190.990 ;
        RECT 83.810 190.790 84.130 190.850 ;
        RECT 86.570 190.790 86.890 190.850 ;
        RECT 87.030 190.790 87.350 191.050 ;
        RECT 93.010 190.990 93.330 191.050 ;
        RECT 95.325 190.990 95.615 191.035 ;
        RECT 93.010 190.850 95.615 190.990 ;
        RECT 97.240 190.990 97.380 191.825 ;
        RECT 112.330 191.810 112.650 191.870 ;
        RECT 115.565 191.825 115.855 191.870 ;
        RECT 125.300 191.870 127.740 192.010 ;
        RECT 97.610 191.670 97.930 191.730 ;
        RECT 98.085 191.670 98.375 191.715 ;
        RECT 97.610 191.530 98.375 191.670 ;
        RECT 97.610 191.470 97.930 191.530 ;
        RECT 98.085 191.485 98.375 191.530 ;
        RECT 98.545 191.485 98.835 191.715 ;
        RECT 99.465 191.670 99.755 191.715 ;
        RECT 102.670 191.670 102.990 191.730 ;
        RECT 99.465 191.530 102.990 191.670 ;
        RECT 99.465 191.485 99.755 191.530 ;
        RECT 98.070 190.990 98.390 191.050 ;
        RECT 97.240 190.850 98.390 190.990 ;
        RECT 93.010 190.790 93.330 190.850 ;
        RECT 95.325 190.805 95.615 190.850 ;
        RECT 98.070 190.790 98.390 190.850 ;
        RECT 88.410 190.650 88.730 190.710 ;
        RECT 82.060 190.510 88.730 190.650 ;
        RECT 70.470 190.450 70.790 190.510 ;
        RECT 73.690 190.450 74.010 190.510 ;
        RECT 80.130 190.450 80.450 190.510 ;
        RECT 88.410 190.450 88.730 190.510 ;
        RECT 92.550 190.450 92.870 190.710 ;
        RECT 94.390 190.450 94.710 190.710 ;
        RECT 96.230 190.650 96.550 190.710 ;
        RECT 98.620 190.650 98.760 191.485 ;
        RECT 102.670 191.470 102.990 191.530 ;
        RECT 103.145 191.485 103.435 191.715 ;
        RECT 99.910 191.130 100.230 191.390 ;
        RECT 102.210 191.330 102.530 191.390 ;
        RECT 101.380 191.190 102.530 191.330 ;
        RECT 103.220 191.330 103.360 191.485 ;
        RECT 104.050 191.470 104.370 191.730 ;
        RECT 105.905 191.670 106.195 191.715 ;
        RECT 107.270 191.670 107.590 191.730 ;
        RECT 110.030 191.670 110.350 191.730 ;
        RECT 105.905 191.530 110.350 191.670 ;
        RECT 105.905 191.485 106.195 191.530 ;
        RECT 107.270 191.470 107.590 191.530 ;
        RECT 110.030 191.470 110.350 191.530 ;
        RECT 115.105 191.670 115.395 191.715 ;
        RECT 121.530 191.670 121.850 191.730 ;
        RECT 115.105 191.530 121.850 191.670 ;
        RECT 115.105 191.485 115.395 191.530 ;
        RECT 121.530 191.470 121.850 191.530 ;
        RECT 124.290 191.670 124.610 191.760 ;
        RECT 124.290 191.530 124.775 191.670 ;
        RECT 124.290 191.500 124.610 191.530 ;
        RECT 124.305 191.485 124.595 191.500 ;
        RECT 108.650 191.330 108.970 191.390 ;
        RECT 112.790 191.330 113.110 191.390 ;
        RECT 103.220 191.190 113.110 191.330 ;
        RECT 98.990 190.990 99.310 191.050 ;
        RECT 101.380 191.035 101.520 191.190 ;
        RECT 102.210 191.130 102.530 191.190 ;
        RECT 108.650 191.130 108.970 191.190 ;
        RECT 112.790 191.130 113.110 191.190 ;
        RECT 116.470 191.330 116.790 191.390 ;
        RECT 125.300 191.330 125.440 191.870 ;
        RECT 125.670 191.670 125.990 191.730 ;
        RECT 126.145 191.670 126.435 191.715 ;
        RECT 125.670 191.530 126.435 191.670 ;
        RECT 125.670 191.470 125.990 191.530 ;
        RECT 126.145 191.485 126.435 191.530 ;
        RECT 127.050 191.470 127.370 191.730 ;
        RECT 127.600 191.715 127.740 191.870 ;
        RECT 127.970 191.870 129.120 192.010 ;
        RECT 127.970 191.810 128.290 191.870 ;
        RECT 127.525 191.485 127.815 191.715 ;
        RECT 128.430 191.670 128.750 191.730 ;
        RECT 128.980 191.715 129.120 191.870 ;
        RECT 129.350 191.810 129.670 192.070 ;
        RECT 130.270 191.810 130.590 192.070 ;
        RECT 128.235 191.530 128.750 191.670 ;
        RECT 128.430 191.470 128.750 191.530 ;
        RECT 128.905 191.485 129.195 191.715 ;
        RECT 129.825 191.670 130.115 191.715 ;
        RECT 130.360 191.670 130.500 191.810 ;
        RECT 129.825 191.530 130.500 191.670 ;
        RECT 130.745 191.670 131.035 191.715 ;
        RECT 131.190 191.670 131.510 191.730 ;
        RECT 131.740 191.715 131.880 192.210 ;
        RECT 132.570 192.210 134.715 192.350 ;
        RECT 132.570 192.150 132.890 192.210 ;
        RECT 134.425 192.165 134.715 192.210 ;
        RECT 137.170 192.350 137.490 192.410 ;
        RECT 137.645 192.350 137.935 192.395 ;
        RECT 137.170 192.210 137.935 192.350 ;
        RECT 137.170 192.150 137.490 192.210 ;
        RECT 137.645 192.165 137.935 192.210 ;
        RECT 133.490 192.010 133.810 192.070 ;
        RECT 133.965 192.010 134.255 192.055 ;
        RECT 133.490 191.870 134.255 192.010 ;
        RECT 133.490 191.810 133.810 191.870 ;
        RECT 133.965 191.825 134.255 191.870 ;
        RECT 130.745 191.530 131.510 191.670 ;
        RECT 129.825 191.485 130.115 191.530 ;
        RECT 130.745 191.485 131.035 191.530 ;
        RECT 131.190 191.470 131.510 191.530 ;
        RECT 131.665 191.485 131.955 191.715 ;
        RECT 132.125 191.485 132.415 191.715 ;
        RECT 132.590 191.670 132.880 191.715 ;
        RECT 133.030 191.670 133.350 191.730 ;
        RECT 132.590 191.530 133.350 191.670 ;
        RECT 132.590 191.485 132.880 191.530 ;
        RECT 116.470 191.190 125.440 191.330 ;
        RECT 126.605 191.330 126.895 191.375 ;
        RECT 129.350 191.330 129.670 191.390 ;
        RECT 126.605 191.190 129.670 191.330 ;
        RECT 116.470 191.130 116.790 191.190 ;
        RECT 126.605 191.145 126.895 191.190 ;
        RECT 129.350 191.130 129.670 191.190 ;
        RECT 130.270 191.330 130.590 191.390 ;
        RECT 132.200 191.330 132.340 191.485 ;
        RECT 133.030 191.470 133.350 191.530 ;
        RECT 136.250 191.470 136.570 191.730 ;
        RECT 130.270 191.190 132.340 191.330 ;
        RECT 130.270 191.130 130.590 191.190 ;
        RECT 136.710 191.130 137.030 191.390 ;
        RECT 101.305 190.990 101.595 191.035 ;
        RECT 98.990 190.850 101.595 190.990 ;
        RECT 98.990 190.790 99.310 190.850 ;
        RECT 101.305 190.805 101.595 190.850 ;
        RECT 101.750 190.990 102.070 191.050 ;
        RECT 104.065 190.990 104.355 191.035 ;
        RECT 101.750 190.850 104.355 190.990 ;
        RECT 101.750 190.790 102.070 190.850 ;
        RECT 104.065 190.805 104.355 190.850 ;
        RECT 106.810 190.990 107.130 191.050 ;
        RECT 110.030 190.990 110.350 191.050 ;
        RECT 106.810 190.850 110.350 190.990 ;
        RECT 106.810 190.790 107.130 190.850 ;
        RECT 110.030 190.790 110.350 190.850 ;
        RECT 114.170 190.990 114.490 191.050 ;
        RECT 117.850 190.990 118.170 191.050 ;
        RECT 123.830 190.990 124.150 191.050 ;
        RECT 135.790 190.990 136.110 191.050 ;
        RECT 137.630 190.990 137.950 191.050 ;
        RECT 114.170 190.850 124.150 190.990 ;
        RECT 114.170 190.790 114.490 190.850 ;
        RECT 117.850 190.790 118.170 190.850 ;
        RECT 123.830 190.790 124.150 190.850 ;
        RECT 124.840 190.850 137.950 190.990 ;
        RECT 99.910 190.650 100.230 190.710 ;
        RECT 96.230 190.510 100.230 190.650 ;
        RECT 96.230 190.450 96.550 190.510 ;
        RECT 99.910 190.450 100.230 190.510 ;
        RECT 102.225 190.650 102.515 190.695 ;
        RECT 104.970 190.650 105.290 190.710 ;
        RECT 102.225 190.510 105.290 190.650 ;
        RECT 102.225 190.465 102.515 190.510 ;
        RECT 104.970 190.450 105.290 190.510 ;
        RECT 106.350 190.650 106.670 190.710 ;
        RECT 124.840 190.650 124.980 190.850 ;
        RECT 135.790 190.790 136.110 190.850 ;
        RECT 137.630 190.790 137.950 190.850 ;
        RECT 106.350 190.510 124.980 190.650 ;
        RECT 125.225 190.650 125.515 190.695 ;
        RECT 125.670 190.650 125.990 190.710 ;
        RECT 125.225 190.510 125.990 190.650 ;
        RECT 106.350 190.450 106.670 190.510 ;
        RECT 125.225 190.465 125.515 190.510 ;
        RECT 125.670 190.450 125.990 190.510 ;
        RECT 27.160 189.830 139.860 190.310 ;
        RECT 31.845 189.630 32.135 189.675 ;
        RECT 32.290 189.630 32.610 189.690 ;
        RECT 31.845 189.490 32.610 189.630 ;
        RECT 31.845 189.445 32.135 189.490 ;
        RECT 32.290 189.430 32.610 189.490 ;
        RECT 37.350 189.430 37.670 189.690 ;
        RECT 41.030 189.630 41.350 189.690 ;
        RECT 42.425 189.630 42.715 189.675 ;
        RECT 43.330 189.630 43.650 189.690 ;
        RECT 41.030 189.490 43.650 189.630 ;
        RECT 41.030 189.430 41.350 189.490 ;
        RECT 42.425 189.445 42.715 189.490 ;
        RECT 43.330 189.430 43.650 189.490 ;
        RECT 47.470 189.630 47.790 189.690 ;
        RECT 53.910 189.630 54.230 189.690 ;
        RECT 47.470 189.490 54.230 189.630 ;
        RECT 47.470 189.430 47.790 189.490 ;
        RECT 53.910 189.430 54.230 189.490 ;
        RECT 54.830 189.630 55.150 189.690 ;
        RECT 55.305 189.630 55.595 189.675 ;
        RECT 54.830 189.490 55.595 189.630 ;
        RECT 54.830 189.430 55.150 189.490 ;
        RECT 55.305 189.445 55.595 189.490 ;
        RECT 56.210 189.430 56.530 189.690 ;
        RECT 57.130 189.430 57.450 189.690 ;
        RECT 59.890 189.630 60.210 189.690 ;
        RECT 69.090 189.630 69.410 189.690 ;
        RECT 59.890 189.490 69.410 189.630 ;
        RECT 59.890 189.430 60.210 189.490 ;
        RECT 48.850 189.290 49.170 189.350 ;
        RECT 37.440 189.150 49.170 189.290 ;
        RECT 37.440 188.950 37.580 189.150 ;
        RECT 48.850 189.090 49.170 189.150 ;
        RECT 52.070 189.290 52.390 189.350 ;
        RECT 65.870 189.290 66.190 189.350 ;
        RECT 52.070 189.150 66.190 189.290 ;
        RECT 52.070 189.090 52.390 189.150 ;
        RECT 65.870 189.090 66.190 189.150 ;
        RECT 37.825 188.950 38.115 188.995 ;
        RECT 37.440 188.810 38.115 188.950 ;
        RECT 37.825 188.765 38.115 188.810 ;
        RECT 39.665 188.950 39.955 188.995 ;
        RECT 45.630 188.950 45.950 189.010 ;
        RECT 39.665 188.810 45.950 188.950 ;
        RECT 39.665 188.765 39.955 188.810 ;
        RECT 45.630 188.750 45.950 188.810 ;
        RECT 62.650 188.950 62.970 189.010 ;
        RECT 63.585 188.950 63.875 188.995 ;
        RECT 62.650 188.810 63.875 188.950 ;
        RECT 66.420 188.950 66.560 189.490 ;
        RECT 69.090 189.430 69.410 189.490 ;
        RECT 73.690 189.430 74.010 189.690 ;
        RECT 86.110 189.430 86.430 189.690 ;
        RECT 93.470 189.630 93.790 189.690 ;
        RECT 103.590 189.630 103.910 189.690 ;
        RECT 93.470 189.490 103.910 189.630 ;
        RECT 93.470 189.430 93.790 189.490 ;
        RECT 103.590 189.430 103.910 189.490 ;
        RECT 105.890 189.630 106.210 189.690 ;
        RECT 113.710 189.630 114.030 189.690 ;
        RECT 105.890 189.490 114.030 189.630 ;
        RECT 105.890 189.430 106.210 189.490 ;
        RECT 113.710 189.430 114.030 189.490 ;
        RECT 120.165 189.630 120.455 189.675 ;
        RECT 123.370 189.630 123.690 189.690 ;
        RECT 120.165 189.490 123.690 189.630 ;
        RECT 120.165 189.445 120.455 189.490 ;
        RECT 123.370 189.430 123.690 189.490 ;
        RECT 68.170 189.090 68.490 189.350 ;
        RECT 90.725 189.290 91.015 189.335 ;
        RECT 98.070 189.290 98.390 189.350 ;
        RECT 90.725 189.150 98.390 189.290 ;
        RECT 90.725 189.105 91.015 189.150 ;
        RECT 98.070 189.090 98.390 189.150 ;
        RECT 98.530 189.290 98.850 189.350 ;
        RECT 101.750 189.290 102.070 189.350 ;
        RECT 98.530 189.150 102.070 189.290 ;
        RECT 98.530 189.090 98.850 189.150 ;
        RECT 101.750 189.090 102.070 189.150 ;
        RECT 104.050 189.290 104.370 189.350 ;
        RECT 106.350 189.290 106.670 189.350 ;
        RECT 108.190 189.290 108.510 189.350 ;
        RECT 104.050 189.150 106.670 189.290 ;
        RECT 104.050 189.090 104.370 189.150 ;
        RECT 106.350 189.090 106.670 189.150 ;
        RECT 107.360 189.150 108.510 189.290 ;
        RECT 66.805 188.950 67.095 188.995 ;
        RECT 66.420 188.810 67.095 188.950 ;
        RECT 62.650 188.750 62.970 188.810 ;
        RECT 63.585 188.765 63.875 188.810 ;
        RECT 66.805 188.765 67.095 188.810 ;
        RECT 69.105 188.950 69.395 188.995 ;
        RECT 70.470 188.950 70.790 189.010 ;
        RECT 69.105 188.810 70.790 188.950 ;
        RECT 69.105 188.765 69.395 188.810 ;
        RECT 70.470 188.750 70.790 188.810 ;
        RECT 71.850 188.750 72.170 189.010 ;
        RECT 81.050 188.950 81.370 189.010 ;
        RECT 87.030 188.950 87.350 189.010 ;
        RECT 92.550 188.950 92.870 189.010 ;
        RECT 95.310 188.950 95.630 189.010 ;
        RECT 98.990 188.950 99.310 189.010 ;
        RECT 81.050 188.810 87.350 188.950 ;
        RECT 81.050 188.750 81.370 188.810 ;
        RECT 87.030 188.750 87.350 188.810 ;
        RECT 91.260 188.810 95.630 188.950 ;
        RECT 31.370 188.610 31.690 188.670 ;
        RECT 36.430 188.610 36.750 188.670 ;
        RECT 31.370 188.470 36.750 188.610 ;
        RECT 31.370 188.410 31.690 188.470 ;
        RECT 36.430 188.410 36.750 188.470 ;
        RECT 36.905 188.610 37.195 188.655 ;
        RECT 37.350 188.610 37.670 188.670 ;
        RECT 36.905 188.470 37.670 188.610 ;
        RECT 36.905 188.425 37.195 188.470 ;
        RECT 37.350 188.410 37.670 188.470 ;
        RECT 38.285 188.425 38.575 188.655 ;
        RECT 36.520 188.270 36.660 188.410 ;
        RECT 38.360 188.270 38.500 188.425 ;
        RECT 38.730 188.410 39.050 188.670 ;
        RECT 40.110 188.610 40.430 188.670 ;
        RECT 40.585 188.610 40.875 188.655 ;
        RECT 49.310 188.610 49.630 188.670 ;
        RECT 51.625 188.610 51.915 188.655 ;
        RECT 52.070 188.610 52.390 188.670 ;
        RECT 40.110 188.470 43.100 188.610 ;
        RECT 40.110 188.410 40.430 188.470 ;
        RECT 40.585 188.425 40.875 188.470 ;
        RECT 42.960 188.330 43.100 188.470 ;
        RECT 49.310 188.470 52.390 188.610 ;
        RECT 49.310 188.410 49.630 188.470 ;
        RECT 51.625 188.425 51.915 188.470 ;
        RECT 52.070 188.410 52.390 188.470 ;
        RECT 52.990 188.410 53.310 188.670 ;
        RECT 53.450 188.410 53.770 188.670 ;
        RECT 54.370 188.610 54.690 188.670 ;
        RECT 55.765 188.610 56.055 188.655 ;
        RECT 54.370 188.470 56.055 188.610 ;
        RECT 54.370 188.410 54.690 188.470 ;
        RECT 55.765 188.425 56.055 188.470 ;
        RECT 56.670 188.410 56.990 188.670 ;
        RECT 57.145 188.425 57.435 188.655 ;
        RECT 58.065 188.610 58.355 188.655 ;
        RECT 57.680 188.470 58.355 188.610 ;
        RECT 42.425 188.270 42.715 188.315 ;
        RECT 36.520 188.130 42.715 188.270 ;
        RECT 42.425 188.085 42.715 188.130 ;
        RECT 42.870 188.270 43.190 188.330 ;
        RECT 51.150 188.270 51.470 188.330 ;
        RECT 53.540 188.270 53.680 188.410 ;
        RECT 42.870 188.130 52.300 188.270 ;
        RECT 53.540 188.130 56.440 188.270 ;
        RECT 42.870 188.070 43.190 188.130 ;
        RECT 51.150 188.070 51.470 188.130 ;
        RECT 39.665 187.930 39.955 187.975 ;
        RECT 41.490 187.930 41.810 187.990 ;
        RECT 39.665 187.790 41.810 187.930 ;
        RECT 39.665 187.745 39.955 187.790 ;
        RECT 41.490 187.730 41.810 187.790 ;
        RECT 43.345 187.930 43.635 187.975 ;
        RECT 47.470 187.930 47.790 187.990 ;
        RECT 52.160 187.975 52.300 188.130 ;
        RECT 43.345 187.790 47.790 187.930 ;
        RECT 43.345 187.745 43.635 187.790 ;
        RECT 47.470 187.730 47.790 187.790 ;
        RECT 52.085 187.745 52.375 187.975 ;
        RECT 56.300 187.930 56.440 188.130 ;
        RECT 57.220 187.930 57.360 188.425 ;
        RECT 57.680 188.330 57.820 188.470 ;
        RECT 58.065 188.425 58.355 188.470 ;
        RECT 63.125 188.425 63.415 188.655 ;
        RECT 66.330 188.610 66.650 188.670 ;
        RECT 69.565 188.610 69.855 188.655 ;
        RECT 66.330 188.470 69.855 188.610 ;
        RECT 57.590 188.070 57.910 188.330 ;
        RECT 62.190 188.270 62.510 188.330 ;
        RECT 63.200 188.270 63.340 188.425 ;
        RECT 66.330 188.410 66.650 188.470 ;
        RECT 69.565 188.425 69.855 188.470 ;
        RECT 70.945 188.610 71.235 188.655 ;
        RECT 71.390 188.610 71.710 188.670 ;
        RECT 70.945 188.470 71.710 188.610 ;
        RECT 70.945 188.425 71.235 188.470 ;
        RECT 71.390 188.410 71.710 188.470 ;
        RECT 73.705 188.610 73.995 188.655 ;
        RECT 74.150 188.610 74.470 188.670 ;
        RECT 73.705 188.470 74.470 188.610 ;
        RECT 73.705 188.425 73.995 188.470 ;
        RECT 74.150 188.410 74.470 188.470 ;
        RECT 74.610 188.610 74.930 188.670 ;
        RECT 75.085 188.610 75.375 188.655 ;
        RECT 74.610 188.470 75.375 188.610 ;
        RECT 74.610 188.410 74.930 188.470 ;
        RECT 75.085 188.425 75.375 188.470 ;
        RECT 80.130 188.610 80.450 188.670 ;
        RECT 87.505 188.610 87.795 188.655 ;
        RECT 87.950 188.610 88.270 188.670 ;
        RECT 80.130 188.470 87.260 188.610 ;
        RECT 80.130 188.410 80.450 188.470 ;
        RECT 75.990 188.270 76.310 188.330 ;
        RECT 84.730 188.270 85.050 188.330 ;
        RECT 62.190 188.130 73.000 188.270 ;
        RECT 62.190 188.070 62.510 188.130 ;
        RECT 56.300 187.790 57.360 187.930 ;
        RECT 70.025 187.930 70.315 187.975 ;
        RECT 70.470 187.930 70.790 187.990 ;
        RECT 70.025 187.790 70.790 187.930 ;
        RECT 70.025 187.745 70.315 187.790 ;
        RECT 70.470 187.730 70.790 187.790 ;
        RECT 72.310 187.730 72.630 187.990 ;
        RECT 72.860 187.930 73.000 188.130 ;
        RECT 75.990 188.130 85.050 188.270 ;
        RECT 75.990 188.070 76.310 188.130 ;
        RECT 84.730 188.070 85.050 188.130 ;
        RECT 86.110 188.070 86.430 188.330 ;
        RECT 87.120 188.270 87.260 188.470 ;
        RECT 87.505 188.470 88.270 188.610 ;
        RECT 87.505 188.425 87.795 188.470 ;
        RECT 87.950 188.410 88.270 188.470 ;
        RECT 88.410 188.610 88.730 188.670 ;
        RECT 88.885 188.610 89.175 188.655 ;
        RECT 88.410 188.470 89.175 188.610 ;
        RECT 88.410 188.410 88.730 188.470 ;
        RECT 88.885 188.425 89.175 188.470 ;
        RECT 89.330 188.610 89.650 188.670 ;
        RECT 89.805 188.610 90.095 188.655 ;
        RECT 89.330 188.470 90.095 188.610 ;
        RECT 89.330 188.410 89.650 188.470 ;
        RECT 89.805 188.425 90.095 188.470 ;
        RECT 90.250 188.410 90.570 188.670 ;
        RECT 91.260 188.655 91.400 188.810 ;
        RECT 92.550 188.750 92.870 188.810 ;
        RECT 95.310 188.750 95.630 188.810 ;
        RECT 95.860 188.810 99.310 188.950 ;
        RECT 91.185 188.425 91.475 188.655 ;
        RECT 93.025 188.610 93.315 188.655 ;
        RECT 93.025 188.470 94.620 188.610 ;
        RECT 93.025 188.425 93.315 188.470 ;
        RECT 93.100 188.270 93.240 188.425 ;
        RECT 87.120 188.130 93.240 188.270 ;
        RECT 93.470 188.070 93.790 188.330 ;
        RECT 93.930 188.070 94.250 188.330 ;
        RECT 94.480 188.270 94.620 188.470 ;
        RECT 94.850 188.410 95.170 188.670 ;
        RECT 95.860 188.655 96.000 188.810 ;
        RECT 98.990 188.750 99.310 188.810 ;
        RECT 99.450 188.950 99.770 189.010 ;
        RECT 102.210 188.950 102.530 189.010 ;
        RECT 107.360 188.950 107.500 189.150 ;
        RECT 108.190 189.090 108.510 189.150 ;
        RECT 99.450 188.810 107.500 188.950 ;
        RECT 107.745 188.950 108.035 188.995 ;
        RECT 110.950 188.950 111.270 189.010 ;
        RECT 107.745 188.810 111.270 188.950 ;
        RECT 99.450 188.750 99.770 188.810 ;
        RECT 102.210 188.750 102.530 188.810 ;
        RECT 107.745 188.765 108.035 188.810 ;
        RECT 110.950 188.750 111.270 188.810 ;
        RECT 114.170 188.950 114.490 189.010 ;
        RECT 136.265 188.950 136.555 188.995 ;
        RECT 114.170 188.810 136.555 188.950 ;
        RECT 114.170 188.750 114.490 188.810 ;
        RECT 136.265 188.765 136.555 188.810 ;
        RECT 95.785 188.425 96.075 188.655 ;
        RECT 96.705 188.610 96.995 188.655 ;
        RECT 99.910 188.610 100.230 188.670 ;
        RECT 106.350 188.610 106.670 188.670 ;
        RECT 96.705 188.470 99.680 188.610 ;
        RECT 96.705 188.425 96.995 188.470 ;
        RECT 99.540 188.270 99.680 188.470 ;
        RECT 99.910 188.470 106.670 188.610 ;
        RECT 99.910 188.410 100.230 188.470 ;
        RECT 106.350 188.410 106.670 188.470 ;
        RECT 106.825 188.610 107.115 188.655 ;
        RECT 108.650 188.610 108.970 188.670 ;
        RECT 106.825 188.470 108.970 188.610 ;
        RECT 106.825 188.425 107.115 188.470 ;
        RECT 108.650 188.410 108.970 188.470 ;
        RECT 116.945 188.610 117.235 188.655 ;
        RECT 125.210 188.610 125.530 188.670 ;
        RECT 116.945 188.470 125.530 188.610 ;
        RECT 116.945 188.425 117.235 188.470 ;
        RECT 125.210 188.410 125.530 188.470 ;
        RECT 127.065 188.610 127.355 188.655 ;
        RECT 127.510 188.610 127.830 188.670 ;
        RECT 127.065 188.470 127.830 188.610 ;
        RECT 127.065 188.425 127.355 188.470 ;
        RECT 127.510 188.410 127.830 188.470 ;
        RECT 136.725 188.425 137.015 188.655 ;
        RECT 105.905 188.270 106.195 188.315 ;
        RECT 109.125 188.270 109.415 188.315 ;
        RECT 119.230 188.270 119.550 188.330 ;
        RECT 94.480 188.130 96.920 188.270 ;
        RECT 99.540 188.130 103.360 188.270 ;
        RECT 78.290 187.930 78.610 187.990 ;
        RECT 72.860 187.790 78.610 187.930 ;
        RECT 78.290 187.730 78.610 187.790 ;
        RECT 79.670 187.930 79.990 187.990 ;
        RECT 83.350 187.930 83.670 187.990 ;
        RECT 87.045 187.930 87.335 187.975 ;
        RECT 79.670 187.790 87.335 187.930 ;
        RECT 79.670 187.730 79.990 187.790 ;
        RECT 83.350 187.730 83.670 187.790 ;
        RECT 87.045 187.745 87.335 187.790 ;
        RECT 87.490 187.930 87.810 187.990 ;
        RECT 88.885 187.930 89.175 187.975 ;
        RECT 87.490 187.790 89.175 187.930 ;
        RECT 87.490 187.730 87.810 187.790 ;
        RECT 88.885 187.745 89.175 187.790 ;
        RECT 91.170 187.930 91.490 187.990 ;
        RECT 92.105 187.930 92.395 187.975 ;
        RECT 91.170 187.790 92.395 187.930 ;
        RECT 91.170 187.730 91.490 187.790 ;
        RECT 92.105 187.745 92.395 187.790 ;
        RECT 92.550 187.930 92.870 187.990 ;
        RECT 94.020 187.930 94.160 188.070 ;
        RECT 96.780 187.990 96.920 188.130 ;
        RECT 103.220 187.990 103.360 188.130 ;
        RECT 105.905 188.130 108.420 188.270 ;
        RECT 105.905 188.085 106.195 188.130 ;
        RECT 92.550 187.790 94.160 187.930 ;
        RECT 94.390 187.930 94.710 187.990 ;
        RECT 96.245 187.930 96.535 187.975 ;
        RECT 94.390 187.790 96.535 187.930 ;
        RECT 92.550 187.730 92.870 187.790 ;
        RECT 94.390 187.730 94.710 187.790 ;
        RECT 96.245 187.745 96.535 187.790 ;
        RECT 96.690 187.930 97.010 187.990 ;
        RECT 98.530 187.930 98.850 187.990 ;
        RECT 96.690 187.790 98.850 187.930 ;
        RECT 96.690 187.730 97.010 187.790 ;
        RECT 98.530 187.730 98.850 187.790 ;
        RECT 99.450 187.730 99.770 187.990 ;
        RECT 103.130 187.930 103.450 187.990 ;
        RECT 106.810 187.930 107.130 187.990 ;
        RECT 103.130 187.790 107.130 187.930 ;
        RECT 103.130 187.730 103.450 187.790 ;
        RECT 106.810 187.730 107.130 187.790 ;
        RECT 107.270 187.930 107.590 187.990 ;
        RECT 107.745 187.930 108.035 187.975 ;
        RECT 107.270 187.790 108.035 187.930 ;
        RECT 108.280 187.930 108.420 188.130 ;
        RECT 109.125 188.130 119.550 188.270 ;
        RECT 109.125 188.085 109.415 188.130 ;
        RECT 119.230 188.070 119.550 188.130 ;
        RECT 126.590 188.070 126.910 188.330 ;
        RECT 136.800 188.270 136.940 188.425 ;
        RECT 137.630 188.410 137.950 188.670 ;
        RECT 133.580 188.130 136.940 188.270 ;
        RECT 133.580 187.990 133.720 188.130 ;
        RECT 127.510 187.930 127.830 187.990 ;
        RECT 108.280 187.790 127.830 187.930 ;
        RECT 107.270 187.730 107.590 187.790 ;
        RECT 107.745 187.745 108.035 187.790 ;
        RECT 127.510 187.730 127.830 187.790 ;
        RECT 133.490 187.730 133.810 187.990 ;
        RECT 27.160 187.110 139.860 187.590 ;
        RECT 37.810 186.710 38.130 186.970 ;
        RECT 38.730 186.910 39.050 186.970 ;
        RECT 44.265 186.910 44.555 186.955 ;
        RECT 44.710 186.910 45.030 186.970 ;
        RECT 38.730 186.770 45.030 186.910 ;
        RECT 38.730 186.710 39.050 186.770 ;
        RECT 44.265 186.725 44.555 186.770 ;
        RECT 44.710 186.710 45.030 186.770 ;
        RECT 66.330 186.710 66.650 186.970 ;
        RECT 69.550 186.910 69.870 186.970 ;
        RECT 70.945 186.910 71.235 186.955 ;
        RECT 69.550 186.770 71.235 186.910 ;
        RECT 69.550 186.710 69.870 186.770 ;
        RECT 70.945 186.725 71.235 186.770 ;
        RECT 71.865 186.910 72.155 186.955 ;
        RECT 75.070 186.910 75.390 186.970 ;
        RECT 71.865 186.770 75.390 186.910 ;
        RECT 71.865 186.725 72.155 186.770 ;
        RECT 75.070 186.710 75.390 186.770 ;
        RECT 75.530 186.910 75.850 186.970 ;
        RECT 77.370 186.910 77.690 186.970 ;
        RECT 81.095 186.910 81.385 186.955 ;
        RECT 84.775 186.910 85.065 186.955 ;
        RECT 86.110 186.910 86.430 186.970 ;
        RECT 75.530 186.770 80.440 186.910 ;
        RECT 75.530 186.710 75.850 186.770 ;
        RECT 77.370 186.710 77.690 186.770 ;
        RECT 80.300 186.740 80.440 186.770 ;
        RECT 81.095 186.770 82.660 186.910 ;
        RECT 40.125 186.570 40.415 186.615 ;
        RECT 41.490 186.570 41.810 186.630 ;
        RECT 61.730 186.570 62.050 186.630 ;
        RECT 67.250 186.570 67.570 186.630 ;
        RECT 76.450 186.570 76.770 186.630 ;
        RECT 80.300 186.600 80.820 186.740 ;
        RECT 81.095 186.725 81.385 186.770 ;
        RECT 82.520 186.615 82.660 186.770 ;
        RECT 84.775 186.770 86.430 186.910 ;
        RECT 84.775 186.725 85.065 186.770 ;
        RECT 86.110 186.710 86.430 186.770 ;
        RECT 86.570 186.910 86.890 186.970 ;
        RECT 92.550 186.910 92.870 186.970 ;
        RECT 94.865 186.910 95.155 186.955 ;
        RECT 86.570 186.770 92.870 186.910 ;
        RECT 86.570 186.710 86.890 186.770 ;
        RECT 92.550 186.710 92.870 186.770 ;
        RECT 93.560 186.770 95.155 186.910 ;
        RECT 40.125 186.430 41.810 186.570 ;
        RECT 40.125 186.385 40.415 186.430 ;
        RECT 41.490 186.370 41.810 186.430 ;
        RECT 51.240 186.430 55.980 186.570 ;
        RECT 51.240 186.290 51.380 186.430 ;
        RECT 55.840 186.290 55.980 186.430 ;
        RECT 61.730 186.430 67.020 186.570 ;
        RECT 61.730 186.370 62.050 186.430 ;
        RECT 48.850 186.230 49.170 186.290 ;
        RECT 50.245 186.230 50.535 186.275 ;
        RECT 48.850 186.090 50.535 186.230 ;
        RECT 48.850 186.030 49.170 186.090 ;
        RECT 50.245 186.045 50.535 186.090 ;
        RECT 24.470 185.890 24.790 185.950 ;
        RECT 28.625 185.890 28.915 185.935 ;
        RECT 24.470 185.750 28.915 185.890 ;
        RECT 24.470 185.690 24.790 185.750 ;
        RECT 28.625 185.705 28.915 185.750 ;
        RECT 30.005 185.890 30.295 185.935 ;
        RECT 31.830 185.890 32.150 185.950 ;
        RECT 35.525 185.890 35.815 185.935 ;
        RECT 37.350 185.890 37.670 185.950 ;
        RECT 38.730 185.890 39.050 185.950 ;
        RECT 30.005 185.750 39.050 185.890 ;
        RECT 30.005 185.705 30.295 185.750 ;
        RECT 31.830 185.690 32.150 185.750 ;
        RECT 35.525 185.705 35.815 185.750 ;
        RECT 37.350 185.690 37.670 185.750 ;
        RECT 38.730 185.690 39.050 185.750 ;
        RECT 40.570 185.690 40.890 185.950 ;
        RECT 41.170 185.890 41.460 185.935 ;
        RECT 45.645 185.890 45.935 185.935 ;
        RECT 41.170 185.750 45.935 185.890 ;
        RECT 50.320 185.890 50.460 186.045 ;
        RECT 51.150 186.030 51.470 186.290 ;
        RECT 53.465 186.230 53.755 186.275 ;
        RECT 53.910 186.230 54.230 186.290 ;
        RECT 53.465 186.090 54.230 186.230 ;
        RECT 53.465 186.045 53.755 186.090 ;
        RECT 53.910 186.030 54.230 186.090 ;
        RECT 54.370 186.030 54.690 186.290 ;
        RECT 55.750 186.030 56.070 186.290 ;
        RECT 65.410 186.030 65.730 186.290 ;
        RECT 65.870 186.230 66.190 186.290 ;
        RECT 66.345 186.230 66.635 186.275 ;
        RECT 65.870 186.090 66.635 186.230 ;
        RECT 66.880 186.230 67.020 186.430 ;
        RECT 67.250 186.430 69.320 186.570 ;
        RECT 67.250 186.370 67.570 186.430 ;
        RECT 68.645 186.230 68.935 186.275 ;
        RECT 66.880 186.090 68.935 186.230 ;
        RECT 69.180 186.230 69.320 186.430 ;
        RECT 74.240 186.430 76.770 186.570 ;
        RECT 80.680 186.570 80.820 186.600 ;
        RECT 81.525 186.570 81.815 186.615 ;
        RECT 80.680 186.430 81.815 186.570 ;
        RECT 70.960 186.230 71.250 186.275 ;
        RECT 69.180 186.090 71.250 186.230 ;
        RECT 65.870 186.030 66.190 186.090 ;
        RECT 66.345 186.045 66.635 186.090 ;
        RECT 68.645 186.045 68.935 186.090 ;
        RECT 70.960 186.045 71.250 186.090 ;
        RECT 55.290 185.890 55.610 185.950 ;
        RECT 50.320 185.750 55.610 185.890 ;
        RECT 68.720 185.890 68.860 186.045 ;
        RECT 73.690 186.030 74.010 186.290 ;
        RECT 74.240 186.275 74.380 186.430 ;
        RECT 76.450 186.370 76.770 186.430 ;
        RECT 81.525 186.385 81.815 186.430 ;
        RECT 82.445 186.385 82.735 186.615 ;
        RECT 84.270 186.570 84.590 186.630 ;
        RECT 90.250 186.570 90.570 186.630 ;
        RECT 93.560 186.615 93.700 186.770 ;
        RECT 94.865 186.725 95.155 186.770 ;
        RECT 97.150 186.910 97.470 186.970 ;
        RECT 133.950 186.910 134.270 186.970 ;
        RECT 134.425 186.910 134.715 186.955 ;
        RECT 97.150 186.770 132.110 186.910 ;
        RECT 97.150 186.710 97.470 186.770 ;
        RECT 93.485 186.570 93.775 186.615 ;
        RECT 84.270 186.430 90.570 186.570 ;
        RECT 84.270 186.370 84.590 186.430 ;
        RECT 90.250 186.370 90.570 186.430 ;
        RECT 91.720 186.430 93.775 186.570 ;
        RECT 74.165 186.045 74.455 186.275 ;
        RECT 74.625 186.230 74.915 186.275 ;
        RECT 75.070 186.230 75.390 186.290 ;
        RECT 74.625 186.090 75.390 186.230 ;
        RECT 74.625 186.045 74.915 186.090 ;
        RECT 75.070 186.030 75.390 186.090 ;
        RECT 75.530 186.030 75.850 186.290 ;
        RECT 75.990 186.030 76.310 186.290 ;
        RECT 76.910 186.030 77.230 186.290 ;
        RECT 77.830 186.030 78.150 186.290 ;
        RECT 79.210 186.030 79.530 186.290 ;
        RECT 79.670 186.260 79.990 186.290 ;
        RECT 80.145 186.260 80.435 186.325 ;
        RECT 79.670 186.120 80.435 186.260 ;
        RECT 79.670 186.030 79.990 186.120 ;
        RECT 80.145 186.095 80.435 186.120 ;
        RECT 80.605 186.240 80.895 186.275 ;
        RECT 80.605 186.100 81.280 186.240 ;
        RECT 80.605 186.045 80.895 186.100 ;
        RECT 73.780 185.890 73.920 186.030 ;
        RECT 76.450 185.890 76.770 185.950 ;
        RECT 68.720 185.750 73.460 185.890 ;
        RECT 73.780 185.750 76.770 185.890 ;
        RECT 41.170 185.705 41.460 185.750 ;
        RECT 45.645 185.705 45.935 185.750 ;
        RECT 36.430 185.550 36.750 185.610 ;
        RECT 36.905 185.550 37.195 185.595 ;
        RECT 40.110 185.550 40.430 185.610 ;
        RECT 41.245 185.550 41.385 185.705 ;
        RECT 55.290 185.690 55.610 185.750 ;
        RECT 42.425 185.550 42.715 185.595 ;
        RECT 43.330 185.550 43.650 185.610 ;
        RECT 36.430 185.410 41.385 185.550 ;
        RECT 41.580 185.410 43.650 185.550 ;
        RECT 36.430 185.350 36.750 185.410 ;
        RECT 36.905 185.365 37.195 185.410 ;
        RECT 40.110 185.350 40.430 185.410 ;
        RECT 41.030 185.210 41.350 185.270 ;
        RECT 41.580 185.210 41.720 185.410 ;
        RECT 42.425 185.365 42.715 185.410 ;
        RECT 43.330 185.350 43.650 185.410 ;
        RECT 44.710 185.550 45.030 185.610 ;
        RECT 47.025 185.550 47.315 185.595 ;
        RECT 52.990 185.550 53.310 185.610 ;
        RECT 54.370 185.550 54.690 185.610 ;
        RECT 68.170 185.550 68.490 185.610 ;
        RECT 44.710 185.410 47.315 185.550 ;
        RECT 44.710 185.350 45.030 185.410 ;
        RECT 47.025 185.365 47.315 185.410 ;
        RECT 47.560 185.410 54.690 185.550 ;
        RECT 41.030 185.070 41.720 185.210 ;
        RECT 41.030 185.010 41.350 185.070 ;
        RECT 41.950 185.010 42.270 185.270 ;
        RECT 42.870 185.210 43.190 185.270 ;
        RECT 44.265 185.210 44.555 185.255 ;
        RECT 42.870 185.070 44.555 185.210 ;
        RECT 42.870 185.010 43.190 185.070 ;
        RECT 44.265 185.025 44.555 185.070 ;
        RECT 45.170 185.210 45.490 185.270 ;
        RECT 47.560 185.210 47.700 185.410 ;
        RECT 52.990 185.350 53.310 185.410 ;
        RECT 54.370 185.350 54.690 185.410 ;
        RECT 54.920 185.410 68.490 185.550 ;
        RECT 45.170 185.070 47.700 185.210 ;
        RECT 47.945 185.210 48.235 185.255 ;
        RECT 48.850 185.210 49.170 185.270 ;
        RECT 47.945 185.070 49.170 185.210 ;
        RECT 45.170 185.010 45.490 185.070 ;
        RECT 47.945 185.025 48.235 185.070 ;
        RECT 48.850 185.010 49.170 185.070 ;
        RECT 49.310 185.010 49.630 185.270 ;
        RECT 51.610 185.210 51.930 185.270 ;
        RECT 54.920 185.210 55.060 185.410 ;
        RECT 68.170 185.350 68.490 185.410 ;
        RECT 69.105 185.550 69.395 185.595 ;
        RECT 72.325 185.550 72.615 185.595 ;
        RECT 69.105 185.410 72.615 185.550 ;
        RECT 73.320 185.550 73.460 185.750 ;
        RECT 76.450 185.690 76.770 185.750 ;
        RECT 80.130 185.890 80.450 185.950 ;
        RECT 81.140 185.890 81.280 186.100 ;
        RECT 81.985 186.045 82.275 186.275 ;
        RECT 80.130 185.750 81.280 185.890 ;
        RECT 82.060 185.890 82.200 186.045 ;
        RECT 83.350 186.030 83.670 186.290 ;
        RECT 83.810 186.030 84.130 186.290 ;
        RECT 84.730 186.230 85.050 186.290 ;
        RECT 91.720 186.275 91.860 186.430 ;
        RECT 93.485 186.385 93.775 186.430 ;
        RECT 95.310 186.570 95.630 186.630 ;
        RECT 96.245 186.570 96.535 186.615 ;
        RECT 95.310 186.430 96.535 186.570 ;
        RECT 95.310 186.370 95.630 186.430 ;
        RECT 96.245 186.385 96.535 186.430 ;
        RECT 96.705 186.570 96.995 186.615 ;
        RECT 99.450 186.570 99.770 186.630 ;
        RECT 96.705 186.430 99.770 186.570 ;
        RECT 96.705 186.385 96.995 186.430 ;
        RECT 99.450 186.370 99.770 186.430 ;
        RECT 99.910 186.570 100.230 186.630 ;
        RECT 110.505 186.570 110.795 186.615 ;
        RECT 99.910 186.430 110.795 186.570 ;
        RECT 99.910 186.370 100.230 186.430 ;
        RECT 110.505 186.385 110.795 186.430 ;
        RECT 111.410 186.370 111.730 186.630 ;
        RECT 119.690 186.370 120.010 186.630 ;
        RECT 128.445 186.570 128.735 186.615 ;
        RECT 129.350 186.570 129.670 186.630 ;
        RECT 128.445 186.430 129.670 186.570 ;
        RECT 131.970 186.570 132.110 186.770 ;
        RECT 133.950 186.770 134.715 186.910 ;
        RECT 133.950 186.710 134.270 186.770 ;
        RECT 134.425 186.725 134.715 186.770 ;
        RECT 136.710 186.910 137.030 186.970 ;
        RECT 137.645 186.910 137.935 186.955 ;
        RECT 136.710 186.770 137.935 186.910 ;
        RECT 136.710 186.710 137.030 186.770 ;
        RECT 137.645 186.725 137.935 186.770 ;
        RECT 131.970 186.430 136.480 186.570 ;
        RECT 128.445 186.385 128.735 186.430 ;
        RECT 129.350 186.370 129.670 186.430 ;
        RECT 85.205 186.230 85.495 186.275 ;
        RECT 84.730 186.090 85.495 186.230 ;
        RECT 84.730 186.030 85.050 186.090 ;
        RECT 85.205 186.045 85.495 186.090 ;
        RECT 85.665 186.230 85.955 186.275 ;
        RECT 89.345 186.230 89.635 186.275 ;
        RECT 85.665 186.090 89.635 186.230 ;
        RECT 85.665 186.045 85.955 186.090 ;
        RECT 89.345 186.045 89.635 186.090 ;
        RECT 90.725 186.045 91.015 186.275 ;
        RECT 91.645 186.045 91.935 186.275 ;
        RECT 92.105 186.230 92.395 186.275 ;
        RECT 92.550 186.230 92.870 186.290 ;
        RECT 92.105 186.090 92.870 186.230 ;
        RECT 92.105 186.045 92.395 186.090 ;
        RECT 84.270 185.890 84.590 185.950 ;
        RECT 82.060 185.750 84.590 185.890 ;
        RECT 80.130 185.690 80.450 185.750 ;
        RECT 84.270 185.690 84.590 185.750 ;
        RECT 86.125 185.705 86.415 185.935 ;
        RECT 87.965 185.705 88.255 185.935 ;
        RECT 88.425 185.890 88.715 185.935 ;
        RECT 90.250 185.890 90.570 185.950 ;
        RECT 88.425 185.750 90.570 185.890 ;
        RECT 90.800 185.890 90.940 186.045 ;
        RECT 92.180 185.890 92.320 186.045 ;
        RECT 92.550 186.030 92.870 186.090 ;
        RECT 93.025 186.045 93.315 186.275 ;
        RECT 94.125 186.230 94.415 186.275 ;
        RECT 94.125 186.090 95.540 186.230 ;
        RECT 94.125 186.045 94.415 186.090 ;
        RECT 90.800 185.750 92.320 185.890 ;
        RECT 88.425 185.705 88.715 185.750 ;
        RECT 73.690 185.550 74.010 185.610 ;
        RECT 80.220 185.550 80.360 185.690 ;
        RECT 73.320 185.410 80.360 185.550 ;
        RECT 85.650 185.550 85.970 185.610 ;
        RECT 86.200 185.550 86.340 185.705 ;
        RECT 85.650 185.410 86.340 185.550 ;
        RECT 88.040 185.550 88.180 185.705 ;
        RECT 90.250 185.690 90.570 185.750 ;
        RECT 93.100 185.610 93.240 186.045 ;
        RECT 95.400 185.890 95.540 186.090 ;
        RECT 95.770 186.030 96.090 186.290 ;
        RECT 97.150 186.230 97.470 186.290 ;
        RECT 97.625 186.230 97.915 186.275 ;
        RECT 98.085 186.230 98.375 186.275 ;
        RECT 97.150 186.090 98.375 186.230 ;
        RECT 97.150 186.030 97.470 186.090 ;
        RECT 97.625 186.045 97.915 186.090 ;
        RECT 98.085 186.045 98.375 186.090 ;
        RECT 98.990 186.030 99.310 186.290 ;
        RECT 100.845 186.045 101.135 186.275 ;
        RECT 101.765 186.230 102.055 186.275 ;
        RECT 102.685 186.230 102.975 186.275 ;
        RECT 101.765 186.090 102.975 186.230 ;
        RECT 101.765 186.045 102.055 186.090 ;
        RECT 102.685 186.045 102.975 186.090 ;
        RECT 96.690 185.890 97.010 185.950 ;
        RECT 95.400 185.750 97.010 185.890 ;
        RECT 96.690 185.690 97.010 185.750 ;
        RECT 98.530 185.890 98.850 185.950 ;
        RECT 99.465 185.890 99.755 185.935 ;
        RECT 98.530 185.750 99.755 185.890 ;
        RECT 98.530 185.690 98.850 185.750 ;
        RECT 99.465 185.705 99.755 185.750 ;
        RECT 99.925 185.705 100.215 185.935 ;
        RECT 100.920 185.890 101.060 186.045 ;
        RECT 103.130 186.030 103.450 186.290 ;
        RECT 104.065 186.045 104.355 186.275 ;
        RECT 104.985 186.045 105.275 186.275 ;
        RECT 105.905 186.230 106.195 186.275 ;
        RECT 111.500 186.230 111.640 186.370 ;
        RECT 105.905 186.090 111.640 186.230 ;
        RECT 112.330 186.230 112.650 186.290 ;
        RECT 128.905 186.230 129.195 186.275 ;
        RECT 112.330 186.090 129.195 186.230 ;
        RECT 105.905 186.045 106.195 186.090 ;
        RECT 104.140 185.890 104.280 186.045 ;
        RECT 100.920 185.750 101.980 185.890 ;
        RECT 91.185 185.550 91.475 185.595 ;
        RECT 88.040 185.410 91.475 185.550 ;
        RECT 69.105 185.365 69.395 185.410 ;
        RECT 72.325 185.365 72.615 185.410 ;
        RECT 73.690 185.350 74.010 185.410 ;
        RECT 85.650 185.350 85.970 185.410 ;
        RECT 51.610 185.070 55.060 185.210 ;
        RECT 56.685 185.210 56.975 185.255 ;
        RECT 74.610 185.210 74.930 185.270 ;
        RECT 56.685 185.070 74.930 185.210 ;
        RECT 51.610 185.010 51.930 185.070 ;
        RECT 56.685 185.025 56.975 185.070 ;
        RECT 74.610 185.010 74.930 185.070 ;
        RECT 76.450 185.210 76.770 185.270 ;
        RECT 79.685 185.210 79.975 185.255 ;
        RECT 76.450 185.070 79.975 185.210 ;
        RECT 76.450 185.010 76.770 185.070 ;
        RECT 79.685 185.025 79.975 185.070 ;
        RECT 82.430 185.010 82.750 185.270 ;
        RECT 83.350 185.210 83.670 185.270 ;
        RECT 88.040 185.210 88.180 185.410 ;
        RECT 91.185 185.365 91.475 185.410 ;
        RECT 93.010 185.350 93.330 185.610 ;
        RECT 94.390 185.550 94.710 185.610 ;
        RECT 96.230 185.550 96.550 185.610 ;
        RECT 94.390 185.410 96.550 185.550 ;
        RECT 94.390 185.350 94.710 185.410 ;
        RECT 96.230 185.350 96.550 185.410 ;
        RECT 97.150 185.550 97.470 185.610 ;
        RECT 100.000 185.550 100.140 185.705 ;
        RECT 101.840 185.610 101.980 185.750 ;
        RECT 103.220 185.750 104.280 185.890 ;
        RECT 105.060 185.890 105.200 186.045 ;
        RECT 112.330 186.030 112.650 186.090 ;
        RECT 128.905 186.045 129.195 186.090 ;
        RECT 129.825 186.045 130.115 186.275 ;
        RECT 105.060 185.750 106.120 185.890 ;
        RECT 103.220 185.610 103.360 185.750 ;
        RECT 105.980 185.610 106.120 185.750 ;
        RECT 107.270 185.690 107.590 185.950 ;
        RECT 107.745 185.890 108.035 185.935 ;
        RECT 108.190 185.890 108.510 185.950 ;
        RECT 107.745 185.750 108.510 185.890 ;
        RECT 107.745 185.705 108.035 185.750 ;
        RECT 108.190 185.690 108.510 185.750 ;
        RECT 109.585 185.890 109.875 185.935 ;
        RECT 111.410 185.890 111.730 185.950 ;
        RECT 109.585 185.750 111.730 185.890 ;
        RECT 109.585 185.705 109.875 185.750 ;
        RECT 111.410 185.690 111.730 185.750 ;
        RECT 113.710 185.890 114.030 185.950 ;
        RECT 129.900 185.890 130.040 186.045 ;
        RECT 130.730 186.030 131.050 186.290 ;
        RECT 132.110 186.030 132.430 186.290 ;
        RECT 136.340 186.275 136.480 186.430 ;
        RECT 133.045 186.045 133.335 186.275 ;
        RECT 136.265 186.045 136.555 186.275 ;
        RECT 113.710 185.750 130.040 185.890 ;
        RECT 113.710 185.690 114.030 185.750 ;
        RECT 132.570 185.690 132.890 185.950 ;
        RECT 97.150 185.410 100.140 185.550 ;
        RECT 97.150 185.350 97.470 185.410 ;
        RECT 101.750 185.350 102.070 185.610 ;
        RECT 103.130 185.350 103.450 185.610 ;
        RECT 104.065 185.550 104.355 185.595 ;
        RECT 104.510 185.550 104.830 185.610 ;
        RECT 104.065 185.410 104.830 185.550 ;
        RECT 104.065 185.365 104.355 185.410 ;
        RECT 104.510 185.350 104.830 185.410 ;
        RECT 105.890 185.350 106.210 185.610 ;
        RECT 106.365 185.550 106.655 185.595 ;
        RECT 117.850 185.550 118.170 185.610 ;
        RECT 106.365 185.410 118.170 185.550 ;
        RECT 106.365 185.365 106.655 185.410 ;
        RECT 117.850 185.350 118.170 185.410 ;
        RECT 121.530 185.550 121.850 185.610 ;
        RECT 133.120 185.550 133.260 186.045 ;
        RECT 136.710 185.690 137.030 185.950 ;
        RECT 121.530 185.410 133.260 185.550 ;
        RECT 121.530 185.350 121.850 185.410 ;
        RECT 83.350 185.070 88.180 185.210 ;
        RECT 83.350 185.010 83.670 185.070 ;
        RECT 92.090 185.010 92.410 185.270 ;
        RECT 92.550 185.210 92.870 185.270 ;
        RECT 95.770 185.210 96.090 185.270 ;
        RECT 104.970 185.210 105.290 185.270 ;
        RECT 92.550 185.070 105.290 185.210 ;
        RECT 92.550 185.010 92.870 185.070 ;
        RECT 95.770 185.010 96.090 185.070 ;
        RECT 104.970 185.010 105.290 185.070 ;
        RECT 105.445 185.210 105.735 185.255 ;
        RECT 111.870 185.210 112.190 185.270 ;
        RECT 105.445 185.070 112.190 185.210 ;
        RECT 105.445 185.025 105.735 185.070 ;
        RECT 111.870 185.010 112.190 185.070 ;
        RECT 116.010 185.210 116.330 185.270 ;
        RECT 116.945 185.210 117.235 185.255 ;
        RECT 116.010 185.070 117.235 185.210 ;
        RECT 116.010 185.010 116.330 185.070 ;
        RECT 116.945 185.025 117.235 185.070 ;
        RECT 123.830 185.210 124.150 185.270 ;
        RECT 128.905 185.210 129.195 185.255 ;
        RECT 123.830 185.070 129.195 185.210 ;
        RECT 123.830 185.010 124.150 185.070 ;
        RECT 128.905 185.025 129.195 185.070 ;
        RECT 27.160 184.390 139.860 184.870 ;
        RECT 32.750 184.190 33.070 184.250 ;
        RECT 51.150 184.190 51.470 184.250 ;
        RECT 32.750 184.050 51.470 184.190 ;
        RECT 32.750 183.990 33.070 184.050 ;
        RECT 51.150 183.990 51.470 184.050 ;
        RECT 52.530 184.190 52.850 184.250 ;
        RECT 53.925 184.190 54.215 184.235 ;
        RECT 57.590 184.190 57.910 184.250 ;
        RECT 52.530 184.050 54.215 184.190 ;
        RECT 52.530 183.990 52.850 184.050 ;
        RECT 53.925 184.005 54.215 184.050 ;
        RECT 54.920 184.050 57.910 184.190 ;
        RECT 41.950 183.850 42.270 183.910 ;
        RECT 53.450 183.850 53.770 183.910 ;
        RECT 41.950 183.710 53.770 183.850 ;
        RECT 41.950 183.650 42.270 183.710 ;
        RECT 30.005 183.510 30.295 183.555 ;
        RECT 30.925 183.510 31.215 183.555 ;
        RECT 31.370 183.510 31.690 183.570 ;
        RECT 30.005 183.370 31.690 183.510 ;
        RECT 30.005 183.325 30.295 183.370 ;
        RECT 30.925 183.325 31.215 183.370 ;
        RECT 31.370 183.310 31.690 183.370 ;
        RECT 44.710 183.310 45.030 183.570 ;
        RECT 47.010 183.310 47.330 183.570 ;
        RECT 31.830 182.970 32.150 183.230 ;
        RECT 39.190 183.170 39.510 183.230 ;
        RECT 41.045 183.170 41.335 183.215 ;
        RECT 39.190 183.030 41.335 183.170 ;
        RECT 39.190 182.970 39.510 183.030 ;
        RECT 41.045 182.985 41.335 183.030 ;
        RECT 45.170 183.170 45.490 183.230 ;
        RECT 46.105 183.170 46.395 183.215 ;
        RECT 45.170 183.030 46.395 183.170 ;
        RECT 45.170 182.970 45.490 183.030 ;
        RECT 46.105 182.985 46.395 183.030 ;
        RECT 25.390 182.830 25.710 182.890 ;
        RECT 29.085 182.830 29.375 182.875 ;
        RECT 25.390 182.690 29.375 182.830 ;
        RECT 25.390 182.630 25.710 182.690 ;
        RECT 29.085 182.645 29.375 182.690 ;
        RECT 40.110 182.830 40.430 182.890 ;
        RECT 41.505 182.830 41.795 182.875 ;
        RECT 40.110 182.690 41.795 182.830 ;
        RECT 40.110 182.630 40.430 182.690 ;
        RECT 41.505 182.645 41.795 182.690 ;
        RECT 41.965 182.830 42.255 182.875 ;
        RECT 47.100 182.830 47.240 183.310 ;
        RECT 48.480 183.215 48.620 183.710 ;
        RECT 53.450 183.650 53.770 183.710 ;
        RECT 51.165 183.510 51.455 183.555 ;
        RECT 49.400 183.370 51.455 183.510 ;
        RECT 49.400 183.230 49.540 183.370 ;
        RECT 51.165 183.325 51.455 183.370 ;
        RECT 51.610 183.310 51.930 183.570 ;
        RECT 48.405 182.985 48.695 183.215 ;
        RECT 49.310 182.970 49.630 183.230 ;
        RECT 49.785 183.170 50.075 183.215 ;
        RECT 50.230 183.170 50.550 183.230 ;
        RECT 49.785 183.030 50.550 183.170 ;
        RECT 49.785 182.985 50.075 183.030 ;
        RECT 50.230 182.970 50.550 183.030 ;
        RECT 50.690 182.970 51.010 183.230 ;
        RECT 52.545 183.170 52.835 183.215 ;
        RECT 54.370 183.170 54.690 183.230 ;
        RECT 54.920 183.215 55.060 184.050 ;
        RECT 57.590 183.990 57.910 184.050 ;
        RECT 62.190 183.990 62.510 184.250 ;
        RECT 70.470 183.990 70.790 184.250 ;
        RECT 76.465 184.190 76.755 184.235 ;
        RECT 79.210 184.190 79.530 184.250 ;
        RECT 83.350 184.190 83.670 184.250 ;
        RECT 76.465 184.050 83.670 184.190 ;
        RECT 76.465 184.005 76.755 184.050 ;
        RECT 79.210 183.990 79.530 184.050 ;
        RECT 83.350 183.990 83.670 184.050 ;
        RECT 84.270 183.990 84.590 184.250 ;
        RECT 87.030 184.190 87.350 184.250 ;
        RECT 93.470 184.190 93.790 184.250 ;
        RECT 87.030 184.050 93.790 184.190 ;
        RECT 87.030 183.990 87.350 184.050 ;
        RECT 55.290 183.850 55.610 183.910 ;
        RECT 61.745 183.850 62.035 183.895 ;
        RECT 63.110 183.850 63.430 183.910 ;
        RECT 67.250 183.850 67.570 183.910 ;
        RECT 75.990 183.850 76.310 183.910 ;
        RECT 55.290 183.710 61.040 183.850 ;
        RECT 55.290 183.650 55.610 183.710 ;
        RECT 59.905 183.510 60.195 183.555 ;
        RECT 60.350 183.510 60.670 183.570 ;
        RECT 59.905 183.370 60.670 183.510 ;
        RECT 60.900 183.510 61.040 183.710 ;
        RECT 61.745 183.710 67.570 183.850 ;
        RECT 61.745 183.665 62.035 183.710 ;
        RECT 63.110 183.650 63.430 183.710 ;
        RECT 67.250 183.650 67.570 183.710 ;
        RECT 71.480 183.710 76.310 183.850 ;
        RECT 70.930 183.510 71.250 183.570 ;
        RECT 71.480 183.555 71.620 183.710 ;
        RECT 75.990 183.650 76.310 183.710 ;
        RECT 77.370 183.650 77.690 183.910 ;
        RECT 77.830 183.850 78.150 183.910 ;
        RECT 78.305 183.850 78.595 183.895 ;
        RECT 77.830 183.710 78.595 183.850 ;
        RECT 77.830 183.650 78.150 183.710 ;
        RECT 78.305 183.665 78.595 183.710 ;
        RECT 82.430 183.650 82.750 183.910 ;
        RECT 83.825 183.850 84.115 183.895 ;
        RECT 91.630 183.850 91.950 183.910 ;
        RECT 83.825 183.710 91.950 183.850 ;
        RECT 83.825 183.665 84.115 183.710 ;
        RECT 91.630 183.650 91.950 183.710 ;
        RECT 60.900 183.370 71.250 183.510 ;
        RECT 59.905 183.325 60.195 183.370 ;
        RECT 60.350 183.310 60.670 183.370 ;
        RECT 70.930 183.310 71.250 183.370 ;
        RECT 71.405 183.325 71.695 183.555 ;
        RECT 71.850 183.310 72.170 183.570 ;
        RECT 72.310 183.310 72.630 183.570 ;
        RECT 72.785 183.510 73.075 183.555 ;
        RECT 73.690 183.510 74.010 183.570 ;
        RECT 72.785 183.370 74.010 183.510 ;
        RECT 72.785 183.325 73.075 183.370 ;
        RECT 73.690 183.310 74.010 183.370 ;
        RECT 74.150 183.510 74.470 183.570 ;
        RECT 76.910 183.510 77.230 183.570 ;
        RECT 78.765 183.510 79.055 183.555 ;
        RECT 74.150 183.370 76.220 183.510 ;
        RECT 74.150 183.310 74.470 183.370 ;
        RECT 52.545 183.030 54.690 183.170 ;
        RECT 52.545 182.985 52.835 183.030 ;
        RECT 54.370 182.970 54.690 183.030 ;
        RECT 54.845 182.985 55.135 183.215 ;
        RECT 55.290 182.970 55.610 183.230 ;
        RECT 55.750 183.170 56.070 183.230 ;
        RECT 56.225 183.170 56.515 183.215 ;
        RECT 55.750 183.030 56.515 183.170 ;
        RECT 55.750 182.970 56.070 183.030 ;
        RECT 56.225 182.985 56.515 183.030 ;
        RECT 56.670 182.970 56.990 183.230 ;
        RECT 58.050 183.170 58.370 183.230 ;
        RECT 68.630 183.170 68.950 183.230 ;
        RECT 58.050 183.030 68.950 183.170 ;
        RECT 58.050 182.970 58.370 183.030 ;
        RECT 68.630 182.970 68.950 183.030 ;
        RECT 74.610 182.970 74.930 183.230 ;
        RECT 76.080 183.215 76.220 183.370 ;
        RECT 76.910 183.370 79.055 183.510 ;
        RECT 76.910 183.310 77.230 183.370 ;
        RECT 78.765 183.325 79.055 183.370 ;
        RECT 79.670 183.510 79.990 183.570 ;
        RECT 85.205 183.510 85.495 183.555 ;
        RECT 92.090 183.510 92.410 183.570 ;
        RECT 79.670 183.370 82.200 183.510 ;
        RECT 79.670 183.310 79.990 183.370 ;
        RECT 76.005 182.985 76.295 183.215 ;
        RECT 77.830 182.970 78.150 183.230 ;
        RECT 80.145 183.170 80.435 183.215 ;
        RECT 81.050 183.170 81.370 183.230 ;
        RECT 80.145 183.030 81.370 183.170 ;
        RECT 80.145 182.985 80.435 183.030 ;
        RECT 81.050 182.970 81.370 183.030 ;
        RECT 41.965 182.690 47.240 182.830 ;
        RECT 48.850 182.830 49.170 182.890 ;
        RECT 81.525 182.830 81.815 182.875 ;
        RECT 48.850 182.690 81.815 182.830 ;
        RECT 82.060 182.830 82.200 183.370 ;
        RECT 85.205 183.370 92.410 183.510 ;
        RECT 85.205 183.325 85.495 183.370 ;
        RECT 92.090 183.310 92.410 183.370 ;
        RECT 82.905 183.170 83.195 183.215 ;
        RECT 84.730 183.170 85.050 183.230 ;
        RECT 82.905 183.030 85.050 183.170 ;
        RECT 82.905 182.985 83.195 183.030 ;
        RECT 84.730 182.970 85.050 183.030 ;
        RECT 85.665 182.985 85.955 183.215 ;
        RECT 88.410 183.170 88.730 183.230 ;
        RECT 88.885 183.170 89.175 183.215 ;
        RECT 88.410 183.030 89.175 183.170 ;
        RECT 85.740 182.830 85.880 182.985 ;
        RECT 88.410 182.970 88.730 183.030 ;
        RECT 88.885 182.985 89.175 183.030 ;
        RECT 90.265 183.170 90.555 183.215 ;
        RECT 90.265 183.030 90.940 183.170 ;
        RECT 90.265 182.985 90.555 183.030 ;
        RECT 82.060 182.690 90.480 182.830 ;
        RECT 41.965 182.645 42.255 182.690 ;
        RECT 48.850 182.630 49.170 182.690 ;
        RECT 81.525 182.645 81.815 182.690 ;
        RECT 43.330 182.490 43.650 182.550 ;
        RECT 43.805 182.490 44.095 182.535 ;
        RECT 43.330 182.350 44.095 182.490 ;
        RECT 43.330 182.290 43.650 182.350 ;
        RECT 43.805 182.305 44.095 182.350 ;
        RECT 44.250 182.490 44.570 182.550 ;
        RECT 45.185 182.490 45.475 182.535 ;
        RECT 44.250 182.350 45.475 182.490 ;
        RECT 44.250 182.290 44.570 182.350 ;
        RECT 45.185 182.305 45.475 182.350 ;
        RECT 47.485 182.490 47.775 182.535 ;
        RECT 52.990 182.490 53.310 182.550 ;
        RECT 47.485 182.350 53.310 182.490 ;
        RECT 47.485 182.305 47.775 182.350 ;
        RECT 52.990 182.290 53.310 182.350 ;
        RECT 53.465 182.490 53.755 182.535 ;
        RECT 54.830 182.490 55.150 182.550 ;
        RECT 53.465 182.350 55.150 182.490 ;
        RECT 53.465 182.305 53.755 182.350 ;
        RECT 54.830 182.290 55.150 182.350 ;
        RECT 68.170 182.490 68.490 182.550 ;
        RECT 77.830 182.490 78.150 182.550 ;
        RECT 68.170 182.350 78.150 182.490 ;
        RECT 68.170 182.290 68.490 182.350 ;
        RECT 77.830 182.290 78.150 182.350 ;
        RECT 78.290 182.490 78.610 182.550 ;
        RECT 79.210 182.490 79.530 182.550 ;
        RECT 78.290 182.350 79.530 182.490 ;
        RECT 78.290 182.290 78.610 182.350 ;
        RECT 79.210 182.290 79.530 182.350 ;
        RECT 79.685 182.490 79.975 182.535 ;
        RECT 80.590 182.490 80.910 182.550 ;
        RECT 79.685 182.350 80.910 182.490 ;
        RECT 79.685 182.305 79.975 182.350 ;
        RECT 80.590 182.290 80.910 182.350 ;
        RECT 84.730 182.490 85.050 182.550 ;
        RECT 85.650 182.490 85.970 182.550 ;
        RECT 87.505 182.490 87.795 182.535 ;
        RECT 84.730 182.350 87.795 182.490 ;
        RECT 84.730 182.290 85.050 182.350 ;
        RECT 85.650 182.290 85.970 182.350 ;
        RECT 87.505 182.305 87.795 182.350 ;
        RECT 89.790 182.290 90.110 182.550 ;
        RECT 90.340 182.535 90.480 182.690 ;
        RECT 90.265 182.305 90.555 182.535 ;
        RECT 90.800 182.490 90.940 183.030 ;
        RECT 91.170 182.970 91.490 183.230 ;
        RECT 92.640 182.830 92.780 184.050 ;
        RECT 93.470 183.990 93.790 184.050 ;
        RECT 95.310 184.190 95.630 184.250 ;
        RECT 96.690 184.190 97.010 184.250 ;
        RECT 95.310 184.050 97.010 184.190 ;
        RECT 95.310 183.990 95.630 184.050 ;
        RECT 96.690 183.990 97.010 184.050 ;
        RECT 98.530 184.190 98.850 184.250 ;
        RECT 99.910 184.190 100.230 184.250 ;
        RECT 98.530 184.050 100.230 184.190 ;
        RECT 98.530 183.990 98.850 184.050 ;
        RECT 99.910 183.990 100.230 184.050 ;
        RECT 101.305 184.190 101.595 184.235 ;
        RECT 103.590 184.190 103.910 184.250 ;
        RECT 112.330 184.190 112.650 184.250 ;
        RECT 101.305 184.050 103.910 184.190 ;
        RECT 101.305 184.005 101.595 184.050 ;
        RECT 103.590 183.990 103.910 184.050 ;
        RECT 107.820 184.050 112.650 184.190 ;
        RECT 94.390 183.850 94.710 183.910 ;
        RECT 98.990 183.850 99.310 183.910 ;
        RECT 102.210 183.850 102.530 183.910 ;
        RECT 107.820 183.850 107.960 184.050 ;
        RECT 112.330 183.990 112.650 184.050 ;
        RECT 116.470 183.990 116.790 184.250 ;
        RECT 118.310 184.190 118.630 184.250 ;
        RECT 119.690 184.190 120.010 184.250 ;
        RECT 118.310 184.050 120.010 184.190 ;
        RECT 118.310 183.990 118.630 184.050 ;
        RECT 119.690 183.990 120.010 184.050 ;
        RECT 94.390 183.710 98.300 183.850 ;
        RECT 94.390 183.650 94.710 183.710 ;
        RECT 93.930 183.510 94.250 183.570 ;
        RECT 93.930 183.370 96.000 183.510 ;
        RECT 93.930 183.310 94.250 183.370 ;
        RECT 93.010 183.170 93.330 183.230 ;
        RECT 93.485 183.170 93.775 183.215 ;
        RECT 93.010 183.030 93.775 183.170 ;
        RECT 93.010 182.970 93.330 183.030 ;
        RECT 93.485 182.985 93.775 183.030 ;
        RECT 94.850 183.170 95.170 183.230 ;
        RECT 95.325 183.170 95.615 183.215 ;
        RECT 94.850 183.030 95.615 183.170 ;
        RECT 95.860 183.170 96.000 183.370 ;
        RECT 97.610 183.310 97.930 183.570 ;
        RECT 98.160 183.510 98.300 183.710 ;
        RECT 98.990 183.710 102.530 183.850 ;
        RECT 98.990 183.650 99.310 183.710 ;
        RECT 102.210 183.650 102.530 183.710 ;
        RECT 103.680 183.710 107.960 183.850 ;
        RECT 108.190 183.850 108.510 183.910 ;
        RECT 108.190 183.710 121.300 183.850 ;
        RECT 99.925 183.510 100.215 183.555 ;
        RECT 98.160 183.370 101.520 183.510 ;
        RECT 99.925 183.325 100.215 183.370 ;
        RECT 98.085 183.170 98.375 183.215 ;
        RECT 95.860 183.030 98.375 183.170 ;
        RECT 94.850 182.970 95.170 183.030 ;
        RECT 95.325 182.985 95.615 183.030 ;
        RECT 98.085 182.985 98.375 183.030 ;
        RECT 99.465 183.170 99.755 183.215 ;
        RECT 100.830 183.170 101.150 183.230 ;
        RECT 99.465 183.030 101.150 183.170 ;
        RECT 99.465 182.985 99.755 183.030 ;
        RECT 100.830 182.970 101.150 183.030 ;
        RECT 93.945 182.830 94.235 182.875 ;
        RECT 92.640 182.690 94.235 182.830 ;
        RECT 93.945 182.645 94.235 182.690 ;
        RECT 94.405 182.645 94.695 182.875 ;
        RECT 97.150 182.830 97.470 182.890 ;
        RECT 98.530 182.830 98.850 182.890 ;
        RECT 97.150 182.690 98.850 182.830 ;
        RECT 101.380 182.830 101.520 183.370 ;
        RECT 102.670 182.970 102.990 183.230 ;
        RECT 103.130 182.970 103.450 183.230 ;
        RECT 103.680 183.215 103.820 183.710 ;
        RECT 108.190 183.650 108.510 183.710 ;
        RECT 104.970 183.510 105.290 183.570 ;
        RECT 104.600 183.370 105.290 183.510 ;
        RECT 104.600 183.215 104.740 183.370 ;
        RECT 104.970 183.310 105.290 183.370 ;
        RECT 117.390 183.510 117.710 183.570 ;
        RECT 121.160 183.510 121.300 183.710 ;
        RECT 121.530 183.650 121.850 183.910 ;
        RECT 126.590 183.850 126.910 183.910 ;
        RECT 136.725 183.850 137.015 183.895 ;
        RECT 126.590 183.710 137.015 183.850 ;
        RECT 126.590 183.650 126.910 183.710 ;
        RECT 136.725 183.665 137.015 183.710 ;
        RECT 133.505 183.510 133.795 183.555 ;
        RECT 136.285 183.510 136.575 183.555 ;
        RECT 117.390 183.370 120.840 183.510 ;
        RECT 121.160 183.370 133.260 183.510 ;
        RECT 117.390 183.310 117.710 183.370 ;
        RECT 103.605 182.985 103.895 183.215 ;
        RECT 104.525 182.985 104.815 183.215 ;
        RECT 112.790 183.170 113.110 183.230 ;
        RECT 114.645 183.170 114.935 183.215 ;
        RECT 112.790 183.030 114.935 183.170 ;
        RECT 103.680 182.830 103.820 182.985 ;
        RECT 112.790 182.970 113.110 183.030 ;
        RECT 114.645 182.985 114.935 183.030 ;
        RECT 115.090 183.170 115.410 183.230 ;
        RECT 115.565 183.170 115.855 183.215 ;
        RECT 115.090 183.030 115.855 183.170 ;
        RECT 115.090 182.970 115.410 183.030 ;
        RECT 115.565 182.985 115.855 183.030 ;
        RECT 118.770 182.970 119.090 183.230 ;
        RECT 120.700 183.215 120.840 183.370 ;
        RECT 120.625 182.985 120.915 183.215 ;
        RECT 122.450 182.970 122.770 183.230 ;
        RECT 132.110 182.970 132.430 183.230 ;
        RECT 132.570 182.970 132.890 183.230 ;
        RECT 133.120 183.170 133.260 183.370 ;
        RECT 133.505 183.370 136.575 183.510 ;
        RECT 133.505 183.325 133.795 183.370 ;
        RECT 136.285 183.325 136.575 183.370 ;
        RECT 134.425 183.170 134.715 183.215 ;
        RECT 133.120 183.030 134.715 183.170 ;
        RECT 134.425 182.985 134.715 183.030 ;
        RECT 134.885 182.985 135.175 183.215 ;
        RECT 101.380 182.690 103.820 182.830 ;
        RECT 92.565 182.490 92.855 182.535 ;
        RECT 93.010 182.490 93.330 182.550 ;
        RECT 90.800 182.350 93.330 182.490 ;
        RECT 94.480 182.490 94.620 182.645 ;
        RECT 97.150 182.630 97.470 182.690 ;
        RECT 98.530 182.630 98.850 182.690 ;
        RECT 104.970 182.630 105.290 182.890 ;
        RECT 106.810 182.830 107.130 182.890 ;
        RECT 113.250 182.830 113.570 182.890 ;
        RECT 114.185 182.830 114.475 182.875 ;
        RECT 106.810 182.690 112.095 182.830 ;
        RECT 106.810 182.630 107.130 182.690 ;
        RECT 99.450 182.490 99.770 182.550 ;
        RECT 101.290 182.490 101.610 182.550 ;
        RECT 105.890 182.490 106.210 182.550 ;
        RECT 94.480 182.350 106.210 182.490 ;
        RECT 92.565 182.305 92.855 182.350 ;
        RECT 93.010 182.290 93.330 182.350 ;
        RECT 99.450 182.290 99.770 182.350 ;
        RECT 101.290 182.290 101.610 182.350 ;
        RECT 105.890 182.290 106.210 182.350 ;
        RECT 109.570 182.490 109.890 182.550 ;
        RECT 111.425 182.490 111.715 182.535 ;
        RECT 109.570 182.350 111.715 182.490 ;
        RECT 111.955 182.490 112.095 182.690 ;
        RECT 113.250 182.690 114.475 182.830 ;
        RECT 113.250 182.630 113.570 182.690 ;
        RECT 114.185 182.645 114.475 182.690 ;
        RECT 116.470 182.830 116.790 182.890 ;
        RECT 116.470 182.690 125.900 182.830 ;
        RECT 116.470 182.630 116.790 182.690 ;
        RECT 118.770 182.490 119.090 182.550 ;
        RECT 111.955 182.350 119.090 182.490 ;
        RECT 109.570 182.290 109.890 182.350 ;
        RECT 111.425 182.305 111.715 182.350 ;
        RECT 118.770 182.290 119.090 182.350 ;
        RECT 119.690 182.290 120.010 182.550 ;
        RECT 120.165 182.490 120.455 182.535 ;
        RECT 120.610 182.490 120.930 182.550 ;
        RECT 120.165 182.350 120.930 182.490 ;
        RECT 125.760 182.490 125.900 182.690 ;
        RECT 130.730 182.630 131.050 182.890 ;
        RECT 134.960 182.490 135.100 182.985 ;
        RECT 125.760 182.350 135.100 182.490 ;
        RECT 120.165 182.305 120.455 182.350 ;
        RECT 120.610 182.290 120.930 182.350 ;
        RECT 27.160 181.670 139.860 182.150 ;
        RECT 31.385 181.285 31.675 181.515 ;
        RECT 47.025 181.470 47.315 181.515 ;
        RECT 47.930 181.470 48.250 181.530 ;
        RECT 47.025 181.330 48.250 181.470 ;
        RECT 47.025 181.285 47.315 181.330 ;
        RECT 30.005 180.790 30.295 180.835 ;
        RECT 31.460 180.790 31.600 181.285 ;
        RECT 47.930 181.270 48.250 181.330 ;
        RECT 48.390 181.470 48.710 181.530 ;
        RECT 50.690 181.470 51.010 181.530 ;
        RECT 52.070 181.470 52.390 181.530 ;
        RECT 48.390 181.330 55.980 181.470 ;
        RECT 48.390 181.270 48.710 181.330 ;
        RECT 48.850 181.130 49.170 181.190 ;
        RECT 43.880 180.990 49.170 181.130 ;
        RECT 43.880 180.835 44.020 180.990 ;
        RECT 48.850 180.930 49.170 180.990 ;
        RECT 30.005 180.650 31.600 180.790 ;
        RECT 30.005 180.605 30.295 180.650 ;
        RECT 32.305 180.605 32.595 180.835 ;
        RECT 43.805 180.605 44.095 180.835 ;
        RECT 32.380 180.110 32.520 180.605 ;
        RECT 44.250 180.590 44.570 180.850 ;
        RECT 44.710 180.590 45.030 180.850 ;
        RECT 45.630 180.590 45.950 180.850 ;
        RECT 46.105 180.790 46.395 180.835 ;
        RECT 47.485 180.790 47.775 180.835 ;
        RECT 46.105 180.650 47.775 180.790 ;
        RECT 46.105 180.605 46.395 180.650 ;
        RECT 47.485 180.605 47.775 180.650 ;
        RECT 48.405 180.605 48.695 180.835 ;
        RECT 43.330 180.450 43.650 180.510 ;
        RECT 45.170 180.450 45.490 180.510 ;
        RECT 48.480 180.450 48.620 180.605 ;
        RECT 49.310 180.590 49.630 180.850 ;
        RECT 49.860 180.835 50.000 181.330 ;
        RECT 50.690 181.270 51.010 181.330 ;
        RECT 52.070 181.270 52.390 181.330 ;
        RECT 52.990 181.130 53.310 181.190 ;
        RECT 54.155 181.130 54.445 181.175 ;
        RECT 52.990 180.990 54.445 181.130 ;
        RECT 52.990 180.930 53.310 180.990 ;
        RECT 54.155 180.945 54.445 180.990 ;
        RECT 49.785 180.605 50.075 180.835 ;
        RECT 50.230 180.590 50.550 180.850 ;
        RECT 51.150 180.790 51.470 180.850 ;
        RECT 54.845 180.790 55.135 180.835 ;
        RECT 51.150 180.650 55.135 180.790 ;
        RECT 51.150 180.590 51.470 180.650 ;
        RECT 54.845 180.605 55.135 180.650 ;
        RECT 55.290 180.590 55.610 180.850 ;
        RECT 55.840 180.835 55.980 181.330 ;
        RECT 56.670 181.270 56.990 181.530 ;
        RECT 57.590 181.470 57.910 181.530 ;
        RECT 60.365 181.470 60.655 181.515 ;
        RECT 70.010 181.470 70.330 181.530 ;
        RECT 57.590 181.330 70.330 181.470 ;
        RECT 57.590 181.270 57.910 181.330 ;
        RECT 60.365 181.285 60.655 181.330 ;
        RECT 70.010 181.270 70.330 181.330 ;
        RECT 70.485 181.470 70.775 181.515 ;
        RECT 73.230 181.470 73.550 181.530 ;
        RECT 70.485 181.330 73.550 181.470 ;
        RECT 70.485 181.285 70.775 181.330 ;
        RECT 73.230 181.270 73.550 181.330 ;
        RECT 75.085 181.470 75.375 181.515 ;
        RECT 79.670 181.470 79.990 181.530 ;
        RECT 75.085 181.330 79.990 181.470 ;
        RECT 75.085 181.285 75.375 181.330 ;
        RECT 61.730 181.130 62.050 181.190 ;
        RECT 60.440 180.990 62.050 181.130 ;
        RECT 60.440 180.850 60.580 180.990 ;
        RECT 61.730 180.930 62.050 180.990 ;
        RECT 62.190 180.930 62.510 181.190 ;
        RECT 63.570 181.130 63.890 181.190 ;
        RECT 72.770 181.130 73.090 181.190 ;
        RECT 74.165 181.130 74.455 181.175 ;
        RECT 63.200 180.990 65.640 181.130 ;
        RECT 55.765 180.790 56.055 180.835 ;
        RECT 56.210 180.790 56.530 180.850 ;
        RECT 55.765 180.650 56.530 180.790 ;
        RECT 55.765 180.605 56.055 180.650 ;
        RECT 56.210 180.590 56.530 180.650 ;
        RECT 57.605 180.790 57.895 180.835 ;
        RECT 58.050 180.790 58.370 180.850 ;
        RECT 57.605 180.650 58.370 180.790 ;
        RECT 57.605 180.605 57.895 180.650 ;
        RECT 58.050 180.590 58.370 180.650 ;
        RECT 59.890 180.590 60.210 180.850 ;
        RECT 60.350 180.590 60.670 180.850 ;
        RECT 63.200 180.835 63.340 180.990 ;
        RECT 63.570 180.930 63.890 180.990 ;
        RECT 61.285 180.605 61.575 180.835 ;
        RECT 63.125 180.605 63.415 180.835 ;
        RECT 64.490 180.790 64.810 180.850 ;
        RECT 64.965 180.790 65.255 180.835 ;
        RECT 64.490 180.650 65.255 180.790 ;
        RECT 43.330 180.310 48.620 180.450 ;
        RECT 49.400 180.450 49.540 180.590 ;
        RECT 53.465 180.450 53.755 180.495 ;
        RECT 49.400 180.310 53.755 180.450 ;
        RECT 43.330 180.250 43.650 180.310 ;
        RECT 45.170 180.250 45.490 180.310 ;
        RECT 48.480 180.110 48.620 180.310 ;
        RECT 53.465 180.265 53.755 180.310 ;
        RECT 59.430 180.250 59.750 180.510 ;
        RECT 61.360 180.450 61.500 180.605 ;
        RECT 64.490 180.590 64.810 180.650 ;
        RECT 64.965 180.605 65.255 180.650 ;
        RECT 64.030 180.450 64.350 180.510 ;
        RECT 61.360 180.310 64.350 180.450 ;
        RECT 65.500 180.450 65.640 180.990 ;
        RECT 72.770 180.990 74.455 181.130 ;
        RECT 72.770 180.930 73.090 180.990 ;
        RECT 74.165 180.945 74.455 180.990 ;
        RECT 67.710 180.790 68.030 180.850 ;
        RECT 70.025 180.790 70.315 180.835 ;
        RECT 67.710 180.650 70.315 180.790 ;
        RECT 67.710 180.590 68.030 180.650 ;
        RECT 70.025 180.605 70.315 180.650 ;
        RECT 74.625 180.790 74.915 180.835 ;
        RECT 75.160 180.790 75.300 181.285 ;
        RECT 79.670 181.270 79.990 181.330 ;
        RECT 81.510 181.470 81.830 181.530 ;
        RECT 81.510 181.330 82.660 181.470 ;
        RECT 81.510 181.270 81.830 181.330 ;
        RECT 79.210 181.130 79.530 181.190 ;
        RECT 81.970 181.130 82.290 181.190 ;
        RECT 74.625 180.650 75.300 180.790 ;
        RECT 75.620 180.990 79.530 181.130 ;
        RECT 74.625 180.605 74.915 180.650 ;
        RECT 75.620 180.450 75.760 180.990 ;
        RECT 79.210 180.930 79.530 180.990 ;
        RECT 79.760 180.990 82.290 181.130 ;
        RECT 75.990 180.590 76.310 180.850 ;
        RECT 76.910 180.790 77.230 180.850 ;
        RECT 77.385 180.790 77.675 180.835 ;
        RECT 76.910 180.650 77.675 180.790 ;
        RECT 76.910 180.590 77.230 180.650 ;
        RECT 77.385 180.605 77.675 180.650 ;
        RECT 78.290 180.790 78.610 180.850 ;
        RECT 79.760 180.835 79.900 180.990 ;
        RECT 81.970 180.930 82.290 180.990 ;
        RECT 79.685 180.790 79.975 180.835 ;
        RECT 78.290 180.650 79.975 180.790 ;
        RECT 78.290 180.590 78.610 180.650 ;
        RECT 79.685 180.605 79.975 180.650 ;
        RECT 80.130 180.590 80.450 180.850 ;
        RECT 82.520 180.835 82.660 181.330 ;
        RECT 87.030 181.270 87.350 181.530 ;
        RECT 91.170 181.470 91.490 181.530 ;
        RECT 93.470 181.470 93.790 181.530 ;
        RECT 100.370 181.470 100.690 181.530 ;
        RECT 91.170 181.330 92.780 181.470 ;
        RECT 91.170 181.270 91.490 181.330 ;
        RECT 82.890 181.130 83.210 181.190 ;
        RECT 90.250 181.130 90.570 181.190 ;
        RECT 92.105 181.130 92.395 181.175 ;
        RECT 82.890 180.990 87.720 181.130 ;
        RECT 82.890 180.930 83.210 180.990 ;
        RECT 81.525 180.605 81.815 180.835 ;
        RECT 82.445 180.605 82.735 180.835 ;
        RECT 85.665 180.605 85.955 180.835 ;
        RECT 65.500 180.310 75.760 180.450 ;
        RECT 76.450 180.450 76.770 180.510 ;
        RECT 79.225 180.450 79.515 180.495 ;
        RECT 76.450 180.310 79.515 180.450 ;
        RECT 64.030 180.250 64.350 180.310 ;
        RECT 76.450 180.250 76.770 180.310 ;
        RECT 79.225 180.265 79.515 180.310 ;
        RECT 81.600 180.450 81.740 180.605 ;
        RECT 84.730 180.450 85.050 180.510 ;
        RECT 81.600 180.310 85.050 180.450 ;
        RECT 85.740 180.450 85.880 180.605 ;
        RECT 86.110 180.590 86.430 180.850 ;
        RECT 87.580 180.835 87.720 180.990 ;
        RECT 90.250 180.990 92.395 181.130 ;
        RECT 92.640 181.130 92.780 181.330 ;
        RECT 93.470 181.330 94.620 181.470 ;
        RECT 93.470 181.270 93.790 181.330 ;
        RECT 93.025 181.130 93.315 181.175 ;
        RECT 92.640 180.990 93.315 181.130 ;
        RECT 90.250 180.930 90.570 180.990 ;
        RECT 92.105 180.945 92.395 180.990 ;
        RECT 93.025 180.945 93.315 180.990 ;
        RECT 93.930 180.930 94.250 181.190 ;
        RECT 94.480 181.175 94.620 181.330 ;
        RECT 98.620 181.330 100.690 181.470 ;
        RECT 94.405 180.945 94.695 181.175 ;
        RECT 95.310 181.130 95.630 181.190 ;
        RECT 98.070 181.130 98.390 181.190 ;
        RECT 98.620 181.175 98.760 181.330 ;
        RECT 100.370 181.270 100.690 181.330 ;
        RECT 113.710 181.470 114.030 181.530 ;
        RECT 127.065 181.470 127.355 181.515 ;
        RECT 132.570 181.470 132.890 181.530 ;
        RECT 133.490 181.470 133.810 181.530 ;
        RECT 113.710 181.330 125.900 181.470 ;
        RECT 113.710 181.270 114.030 181.330 ;
        RECT 94.965 180.990 95.630 181.130 ;
        RECT 87.505 180.605 87.795 180.835 ;
        RECT 88.885 180.605 89.175 180.835 ;
        RECT 86.570 180.450 86.890 180.510 ;
        RECT 85.740 180.310 86.890 180.450 ;
        RECT 88.960 180.450 89.100 180.605 ;
        RECT 89.790 180.590 90.110 180.850 ;
        RECT 91.185 180.790 91.475 180.835 ;
        RECT 91.630 180.790 91.950 180.850 ;
        RECT 91.185 180.650 91.950 180.790 ;
        RECT 91.185 180.605 91.475 180.650 ;
        RECT 91.630 180.590 91.950 180.650 ;
        RECT 92.565 180.780 92.855 180.835 ;
        RECT 94.965 180.785 95.105 180.990 ;
        RECT 95.310 180.930 95.630 180.990 ;
        RECT 95.860 180.990 98.390 181.130 ;
        RECT 92.565 180.640 93.240 180.780 ;
        RECT 92.565 180.605 92.855 180.640 ;
        RECT 93.100 180.450 93.240 180.640 ;
        RECT 94.890 180.555 95.180 180.785 ;
        RECT 93.470 180.450 93.790 180.510 ;
        RECT 88.960 180.310 92.320 180.450 ;
        RECT 93.100 180.310 93.790 180.450 ;
        RECT 77.370 180.110 77.690 180.170 ;
        RECT 32.380 179.970 48.160 180.110 ;
        RECT 48.480 179.970 77.690 180.110 ;
        RECT 25.390 179.770 25.710 179.830 ;
        RECT 29.085 179.770 29.375 179.815 ;
        RECT 25.390 179.630 29.375 179.770 ;
        RECT 25.390 179.570 25.710 179.630 ;
        RECT 29.085 179.585 29.375 179.630 ;
        RECT 42.885 179.770 43.175 179.815 ;
        RECT 47.470 179.770 47.790 179.830 ;
        RECT 42.885 179.630 47.790 179.770 ;
        RECT 48.020 179.770 48.160 179.970 ;
        RECT 77.370 179.910 77.690 179.970 ;
        RECT 78.750 180.110 79.070 180.170 ;
        RECT 81.600 180.110 81.740 180.310 ;
        RECT 84.730 180.250 85.050 180.310 ;
        RECT 86.570 180.250 86.890 180.310 ;
        RECT 78.750 179.970 81.740 180.110 ;
        RECT 82.430 180.110 82.750 180.170 ;
        RECT 88.425 180.110 88.715 180.155 ;
        RECT 90.250 180.110 90.570 180.170 ;
        RECT 82.430 179.970 88.715 180.110 ;
        RECT 78.750 179.910 79.070 179.970 ;
        RECT 82.430 179.910 82.750 179.970 ;
        RECT 88.425 179.925 88.715 179.970 ;
        RECT 89.420 179.970 90.570 180.110 ;
        RECT 49.310 179.770 49.630 179.830 ;
        RECT 48.020 179.630 49.630 179.770 ;
        RECT 42.885 179.585 43.175 179.630 ;
        RECT 47.470 179.570 47.790 179.630 ;
        RECT 49.310 179.570 49.630 179.630 ;
        RECT 51.150 179.770 51.470 179.830 ;
        RECT 54.370 179.770 54.690 179.830 ;
        RECT 51.150 179.630 54.690 179.770 ;
        RECT 51.150 179.570 51.470 179.630 ;
        RECT 54.370 179.570 54.690 179.630 ;
        RECT 56.210 179.770 56.530 179.830 ;
        RECT 63.570 179.770 63.890 179.830 ;
        RECT 56.210 179.630 63.890 179.770 ;
        RECT 56.210 179.570 56.530 179.630 ;
        RECT 63.570 179.570 63.890 179.630 ;
        RECT 65.870 179.770 66.190 179.830 ;
        RECT 68.170 179.770 68.490 179.830 ;
        RECT 65.870 179.630 68.490 179.770 ;
        RECT 65.870 179.570 66.190 179.630 ;
        RECT 68.170 179.570 68.490 179.630 ;
        RECT 76.910 179.570 77.230 179.830 ;
        RECT 78.305 179.770 78.595 179.815 ;
        RECT 89.420 179.770 89.560 179.970 ;
        RECT 90.250 179.910 90.570 179.970 ;
        RECT 78.305 179.630 89.560 179.770 ;
        RECT 78.305 179.585 78.595 179.630 ;
        RECT 89.790 179.570 90.110 179.830 ;
        RECT 90.710 179.570 91.030 179.830 ;
        RECT 92.180 179.770 92.320 180.310 ;
        RECT 93.470 180.250 93.790 180.310 ;
        RECT 92.550 180.110 92.870 180.170 ;
        RECT 93.025 180.110 93.315 180.155 ;
        RECT 95.860 180.110 96.000 180.990 ;
        RECT 98.070 180.930 98.390 180.990 ;
        RECT 98.545 180.945 98.835 181.175 ;
        RECT 100.845 181.130 101.135 181.175 ;
        RECT 103.130 181.130 103.450 181.190 ;
        RECT 113.250 181.130 113.570 181.190 ;
        RECT 100.000 180.990 113.570 181.130 ;
        RECT 96.690 180.790 97.010 180.850 ;
        RECT 100.000 180.790 100.140 180.990 ;
        RECT 100.845 180.945 101.135 180.990 ;
        RECT 103.130 180.930 103.450 180.990 ;
        RECT 113.250 180.930 113.570 180.990 ;
        RECT 114.170 180.930 114.490 181.190 ;
        RECT 118.770 181.130 119.090 181.190 ;
        RECT 120.610 181.130 120.930 181.190 ;
        RECT 118.770 180.990 120.930 181.130 ;
        RECT 118.770 180.930 119.090 180.990 ;
        RECT 120.610 180.930 120.930 180.990 ;
        RECT 122.450 181.130 122.770 181.190 ;
        RECT 122.450 180.990 124.520 181.130 ;
        RECT 122.450 180.930 122.770 180.990 ;
        RECT 96.690 180.650 100.140 180.790 ;
        RECT 96.690 180.590 97.010 180.650 ;
        RECT 100.370 180.590 100.690 180.850 ;
        RECT 101.305 180.605 101.595 180.835 ;
        RECT 96.230 180.450 96.550 180.510 ;
        RECT 101.380 180.450 101.520 180.605 ;
        RECT 102.210 180.590 102.530 180.850 ;
        RECT 102.670 180.590 102.990 180.850 ;
        RECT 106.350 180.790 106.670 180.850 ;
        RECT 119.690 180.790 120.010 180.850 ;
        RECT 103.220 180.650 120.010 180.790 ;
        RECT 96.230 180.310 101.520 180.450 ;
        RECT 102.300 180.450 102.440 180.590 ;
        RECT 103.220 180.450 103.360 180.650 ;
        RECT 106.350 180.590 106.670 180.650 ;
        RECT 119.690 180.590 120.010 180.650 ;
        RECT 123.370 180.590 123.690 180.850 ;
        RECT 123.830 180.590 124.150 180.850 ;
        RECT 102.300 180.310 103.360 180.450 ;
        RECT 107.270 180.450 107.590 180.510 ;
        RECT 115.550 180.450 115.870 180.510 ;
        RECT 107.270 180.310 115.870 180.450 ;
        RECT 124.380 180.450 124.520 180.990 ;
        RECT 125.760 180.835 125.900 181.330 ;
        RECT 127.065 181.330 132.890 181.470 ;
        RECT 127.065 181.285 127.355 181.330 ;
        RECT 132.570 181.270 132.890 181.330 ;
        RECT 133.120 181.330 133.810 181.470 ;
        RECT 127.510 181.130 127.830 181.190 ;
        RECT 127.985 181.130 128.275 181.175 ;
        RECT 133.120 181.130 133.260 181.330 ;
        RECT 133.490 181.270 133.810 181.330 ;
        RECT 127.510 180.990 128.275 181.130 ;
        RECT 127.510 180.930 127.830 180.990 ;
        RECT 127.985 180.945 128.275 180.990 ;
        RECT 131.970 180.990 133.260 181.130 ;
        RECT 133.580 180.990 136.480 181.130 ;
        RECT 125.685 180.605 125.975 180.835 ;
        RECT 128.430 180.590 128.750 180.850 ;
        RECT 129.365 180.790 129.655 180.835 ;
        RECT 131.970 180.790 132.110 180.990 ;
        RECT 128.980 180.650 132.110 180.790 ;
        RECT 124.765 180.450 125.055 180.495 ;
        RECT 124.380 180.310 125.055 180.450 ;
        RECT 96.230 180.250 96.550 180.310 ;
        RECT 107.270 180.250 107.590 180.310 ;
        RECT 115.550 180.250 115.870 180.310 ;
        RECT 124.765 180.265 125.055 180.310 ;
        RECT 125.210 180.250 125.530 180.510 ;
        RECT 126.145 180.450 126.435 180.495 ;
        RECT 126.590 180.450 126.910 180.510 ;
        RECT 126.145 180.310 126.910 180.450 ;
        RECT 126.145 180.265 126.435 180.310 ;
        RECT 126.590 180.250 126.910 180.310 ;
        RECT 92.550 179.970 93.315 180.110 ;
        RECT 92.550 179.910 92.870 179.970 ;
        RECT 93.025 179.925 93.315 179.970 ;
        RECT 94.025 179.970 96.000 180.110 ;
        RECT 97.610 180.110 97.930 180.170 ;
        RECT 128.980 180.110 129.120 180.650 ;
        RECT 129.365 180.605 129.655 180.650 ;
        RECT 132.570 180.590 132.890 180.850 ;
        RECT 133.045 180.790 133.335 180.835 ;
        RECT 133.580 180.790 133.720 180.990 ;
        RECT 136.340 180.850 136.480 180.990 ;
        RECT 133.045 180.650 133.720 180.790 ;
        RECT 133.950 180.790 134.270 180.850 ;
        RECT 135.345 180.790 135.635 180.835 ;
        RECT 133.950 180.650 135.635 180.790 ;
        RECT 133.045 180.605 133.335 180.650 ;
        RECT 133.950 180.590 134.270 180.650 ;
        RECT 135.345 180.605 135.635 180.650 ;
        RECT 136.250 180.590 136.570 180.850 ;
        RECT 136.725 180.605 137.015 180.835 ;
        RECT 132.660 180.450 132.800 180.590 ;
        RECT 136.800 180.450 136.940 180.605 ;
        RECT 132.660 180.310 136.940 180.450 ;
        RECT 97.610 179.970 129.120 180.110 ;
        RECT 133.505 180.110 133.795 180.155 ;
        RECT 134.870 180.110 135.190 180.170 ;
        RECT 133.505 179.970 135.190 180.110 ;
        RECT 94.025 179.770 94.165 179.970 ;
        RECT 97.610 179.910 97.930 179.970 ;
        RECT 133.505 179.925 133.795 179.970 ;
        RECT 134.870 179.910 135.190 179.970 ;
        RECT 135.790 179.910 136.110 180.170 ;
        RECT 92.180 179.630 94.165 179.770 ;
        RECT 94.390 179.770 94.710 179.830 ;
        RECT 99.465 179.770 99.755 179.815 ;
        RECT 94.390 179.630 99.755 179.770 ;
        RECT 94.390 179.570 94.710 179.630 ;
        RECT 99.465 179.585 99.755 179.630 ;
        RECT 100.370 179.770 100.690 179.830 ;
        RECT 103.130 179.770 103.450 179.830 ;
        RECT 100.370 179.630 103.450 179.770 ;
        RECT 100.370 179.570 100.690 179.630 ;
        RECT 103.130 179.570 103.450 179.630 ;
        RECT 103.605 179.770 103.895 179.815 ;
        RECT 104.050 179.770 104.370 179.830 ;
        RECT 103.605 179.630 104.370 179.770 ;
        RECT 103.605 179.585 103.895 179.630 ;
        RECT 104.050 179.570 104.370 179.630 ;
        RECT 107.730 179.570 108.050 179.830 ;
        RECT 116.930 179.570 117.250 179.830 ;
        RECT 118.310 179.770 118.630 179.830 ;
        RECT 122.450 179.770 122.770 179.830 ;
        RECT 118.310 179.630 122.770 179.770 ;
        RECT 118.310 179.570 118.630 179.630 ;
        RECT 122.450 179.570 122.770 179.630 ;
        RECT 122.910 179.770 123.230 179.830 ;
        RECT 131.665 179.770 131.955 179.815 ;
        RECT 122.910 179.630 131.955 179.770 ;
        RECT 122.910 179.570 123.230 179.630 ;
        RECT 131.665 179.585 131.955 179.630 ;
        RECT 137.630 179.570 137.950 179.830 ;
        RECT 27.160 178.950 139.860 179.430 ;
        RECT 44.710 178.550 45.030 178.810 ;
        RECT 46.565 178.750 46.855 178.795 ;
        RECT 51.610 178.750 51.930 178.810 ;
        RECT 46.565 178.610 51.930 178.750 ;
        RECT 46.565 178.565 46.855 178.610 ;
        RECT 42.885 178.225 43.175 178.455 ;
        RECT 43.345 178.410 43.635 178.455 ;
        RECT 46.090 178.410 46.410 178.470 ;
        RECT 46.640 178.410 46.780 178.565 ;
        RECT 51.610 178.550 51.930 178.610 ;
        RECT 61.745 178.750 62.035 178.795 ;
        RECT 65.870 178.750 66.190 178.810 ;
        RECT 61.745 178.610 66.190 178.750 ;
        RECT 61.745 178.565 62.035 178.610 ;
        RECT 65.870 178.550 66.190 178.610 ;
        RECT 69.550 178.550 69.870 178.810 ;
        RECT 70.945 178.750 71.235 178.795 ;
        RECT 83.365 178.750 83.655 178.795 ;
        RECT 83.810 178.750 84.130 178.810 ;
        RECT 87.045 178.750 87.335 178.795 ;
        RECT 70.945 178.610 78.980 178.750 ;
        RECT 70.945 178.565 71.235 178.610 ;
        RECT 43.345 178.270 46.780 178.410 ;
        RECT 43.345 178.225 43.635 178.270 ;
        RECT 41.490 178.070 41.810 178.130 ;
        RECT 42.960 178.070 43.100 178.225 ;
        RECT 46.090 178.210 46.410 178.270 ;
        RECT 57.130 178.210 57.450 178.470 ;
        RECT 61.270 178.410 61.590 178.470 ;
        RECT 66.790 178.410 67.110 178.470 ;
        RECT 61.270 178.270 62.880 178.410 ;
        RECT 61.270 178.210 61.590 178.270 ;
        RECT 47.025 178.070 47.315 178.115 ;
        RECT 51.150 178.070 51.470 178.130 ;
        RECT 59.890 178.070 60.210 178.130 ;
        RECT 41.490 177.930 46.320 178.070 ;
        RECT 41.490 177.870 41.810 177.930 ;
        RECT 45.170 177.730 45.490 177.790 ;
        RECT 45.645 177.730 45.935 177.775 ;
        RECT 45.170 177.590 45.935 177.730 ;
        RECT 46.180 177.730 46.320 177.930 ;
        RECT 47.025 177.930 51.470 178.070 ;
        RECT 47.025 177.885 47.315 177.930 ;
        RECT 51.150 177.870 51.470 177.930 ;
        RECT 55.380 177.930 60.210 178.070 ;
        RECT 49.770 177.730 50.090 177.790 ;
        RECT 55.380 177.775 55.520 177.930 ;
        RECT 59.890 177.870 60.210 177.930 ;
        RECT 46.180 177.590 50.090 177.730 ;
        RECT 45.170 177.530 45.490 177.590 ;
        RECT 45.645 177.545 45.935 177.590 ;
        RECT 49.770 177.530 50.090 177.590 ;
        RECT 55.305 177.545 55.595 177.775 ;
        RECT 56.075 177.730 56.365 177.775 ;
        RECT 58.050 177.730 58.370 177.790 ;
        RECT 56.075 177.590 58.370 177.730 ;
        RECT 56.075 177.545 56.365 177.590 ;
        RECT 58.050 177.530 58.370 177.590 ;
        RECT 60.810 177.530 61.130 177.790 ;
        RECT 61.730 177.530 62.050 177.790 ;
        RECT 62.740 177.775 62.880 178.270 ;
        RECT 63.660 178.270 67.940 178.410 ;
        RECT 63.660 177.775 63.800 178.270 ;
        RECT 66.790 178.210 67.110 178.270 ;
        RECT 65.870 178.070 66.190 178.130 ;
        RECT 65.870 177.930 67.020 178.070 ;
        RECT 65.870 177.870 66.190 177.930 ;
        RECT 62.205 177.545 62.495 177.775 ;
        RECT 62.665 177.545 62.955 177.775 ;
        RECT 63.585 177.545 63.875 177.775 ;
        RECT 41.030 177.390 41.350 177.450 ;
        RECT 42.870 177.390 43.190 177.450 ;
        RECT 41.030 177.250 43.190 177.390 ;
        RECT 41.030 177.190 41.350 177.250 ;
        RECT 42.870 177.190 43.190 177.250 ;
        RECT 62.280 177.050 62.420 177.545 ;
        RECT 64.490 177.530 64.810 177.790 ;
        RECT 66.330 177.530 66.650 177.790 ;
        RECT 66.880 177.775 67.020 177.930 ;
        RECT 67.800 177.775 67.940 178.270 ;
        RECT 68.630 178.210 68.950 178.470 ;
        RECT 74.610 178.210 74.930 178.470 ;
        RECT 77.370 178.210 77.690 178.470 ;
        RECT 77.830 178.210 78.150 178.470 ;
        RECT 68.720 178.070 68.860 178.210 ;
        RECT 77.460 178.070 77.600 178.210 ;
        RECT 68.260 177.930 68.860 178.070 ;
        RECT 77.000 177.930 77.600 178.070 ;
        RECT 68.260 177.775 68.400 177.930 ;
        RECT 66.805 177.545 67.095 177.775 ;
        RECT 67.725 177.545 68.015 177.775 ;
        RECT 68.185 177.545 68.475 177.775 ;
        RECT 64.045 177.390 64.335 177.435 ;
        RECT 68.260 177.390 68.400 177.545 ;
        RECT 68.630 177.530 68.950 177.790 ;
        RECT 70.010 177.530 70.330 177.790 ;
        RECT 70.930 177.530 71.250 177.790 ;
        RECT 73.705 177.730 73.995 177.775 ;
        RECT 76.005 177.730 76.295 177.775 ;
        RECT 77.000 177.730 77.140 177.930 ;
        RECT 73.705 177.590 74.105 177.730 ;
        RECT 76.005 177.590 77.140 177.730 ;
        RECT 73.705 177.545 73.995 177.590 ;
        RECT 76.005 177.545 76.295 177.590 ;
        RECT 64.045 177.250 68.400 177.390 ;
        RECT 73.245 177.390 73.535 177.435 ;
        RECT 73.780 177.390 73.920 177.545 ;
        RECT 74.610 177.390 74.930 177.450 ;
        RECT 73.245 177.250 74.930 177.390 ;
        RECT 77.000 177.390 77.140 177.590 ;
        RECT 77.385 177.730 77.675 177.775 ;
        RECT 78.290 177.730 78.610 177.790 ;
        RECT 77.385 177.590 78.610 177.730 ;
        RECT 77.385 177.545 77.675 177.590 ;
        RECT 78.290 177.530 78.610 177.590 ;
        RECT 77.845 177.390 78.135 177.435 ;
        RECT 77.000 177.250 78.135 177.390 ;
        RECT 78.840 177.390 78.980 178.610 ;
        RECT 83.365 178.610 84.130 178.750 ;
        RECT 83.365 178.565 83.655 178.610 ;
        RECT 83.810 178.550 84.130 178.610 ;
        RECT 84.360 178.610 87.335 178.750 ;
        RECT 81.510 178.410 81.830 178.470 ;
        RECT 84.360 178.410 84.500 178.610 ;
        RECT 87.045 178.565 87.335 178.610 ;
        RECT 88.410 178.750 88.730 178.810 ;
        RECT 91.185 178.750 91.475 178.795 ;
        RECT 88.410 178.610 91.475 178.750 ;
        RECT 88.410 178.550 88.730 178.610 ;
        RECT 91.185 178.565 91.475 178.610 ;
        RECT 91.630 178.750 91.950 178.810 ;
        RECT 94.390 178.750 94.710 178.810 ;
        RECT 91.630 178.610 94.710 178.750 ;
        RECT 91.630 178.550 91.950 178.610 ;
        RECT 94.390 178.550 94.710 178.610 ;
        RECT 95.785 178.750 96.075 178.795 ;
        RECT 97.150 178.750 97.470 178.810 ;
        RECT 95.785 178.610 97.470 178.750 ;
        RECT 95.785 178.565 96.075 178.610 ;
        RECT 97.150 178.550 97.470 178.610 ;
        RECT 100.370 178.750 100.690 178.810 ;
        RECT 100.845 178.750 101.135 178.795 ;
        RECT 100.370 178.610 101.135 178.750 ;
        RECT 100.370 178.550 100.690 178.610 ;
        RECT 100.845 178.565 101.135 178.610 ;
        RECT 101.290 178.750 101.610 178.810 ;
        RECT 102.210 178.750 102.530 178.810 ;
        RECT 118.310 178.750 118.630 178.810 ;
        RECT 101.290 178.610 118.630 178.750 ;
        RECT 101.290 178.550 101.610 178.610 ;
        RECT 102.210 178.550 102.530 178.610 ;
        RECT 118.310 178.550 118.630 178.610 ;
        RECT 123.370 178.750 123.690 178.810 ;
        RECT 132.125 178.750 132.415 178.795 ;
        RECT 123.370 178.610 132.415 178.750 ;
        RECT 123.370 178.550 123.690 178.610 ;
        RECT 132.125 178.565 132.415 178.610 ;
        RECT 136.710 178.750 137.030 178.810 ;
        RECT 138.105 178.750 138.395 178.795 ;
        RECT 136.710 178.610 138.395 178.750 ;
        RECT 136.710 178.550 137.030 178.610 ;
        RECT 138.105 178.565 138.395 178.610 ;
        RECT 81.510 178.270 84.500 178.410 ;
        RECT 89.345 178.410 89.635 178.455 ;
        RECT 102.670 178.410 102.990 178.470 ;
        RECT 89.345 178.270 102.990 178.410 ;
        RECT 81.510 178.210 81.830 178.270 ;
        RECT 89.345 178.225 89.635 178.270 ;
        RECT 102.670 178.210 102.990 178.270 ;
        RECT 103.590 178.410 103.910 178.470 ;
        RECT 107.285 178.410 107.575 178.455 ;
        RECT 118.770 178.410 119.090 178.470 ;
        RECT 103.590 178.270 119.090 178.410 ;
        RECT 103.590 178.210 103.910 178.270 ;
        RECT 107.285 178.225 107.575 178.270 ;
        RECT 118.770 178.210 119.090 178.270 ;
        RECT 121.545 178.410 121.835 178.455 ;
        RECT 121.990 178.410 122.310 178.470 ;
        RECT 121.545 178.270 122.310 178.410 ;
        RECT 121.545 178.225 121.835 178.270 ;
        RECT 121.990 178.210 122.310 178.270 ;
        RECT 122.450 178.410 122.770 178.470 ;
        RECT 126.590 178.410 126.910 178.470 ;
        RECT 122.450 178.270 126.910 178.410 ;
        RECT 122.450 178.210 122.770 178.270 ;
        RECT 126.590 178.210 126.910 178.270 ;
        RECT 128.890 178.210 129.210 178.470 ;
        RECT 129.350 178.410 129.670 178.470 ;
        RECT 135.790 178.410 136.110 178.470 ;
        RECT 129.350 178.270 136.110 178.410 ;
        RECT 129.350 178.210 129.670 178.270 ;
        RECT 135.790 178.210 136.110 178.270 ;
        RECT 83.350 178.070 83.670 178.130 ;
        RECT 88.870 178.070 89.190 178.130 ;
        RECT 97.150 178.070 97.470 178.130 ;
        RECT 83.350 177.930 84.960 178.070 ;
        RECT 83.350 177.870 83.670 177.930 ;
        RECT 79.210 177.730 79.530 177.790 ;
        RECT 81.050 177.730 81.370 177.790 ;
        RECT 79.210 177.590 81.370 177.730 ;
        RECT 79.210 177.530 79.530 177.590 ;
        RECT 81.050 177.530 81.370 177.590 ;
        RECT 81.525 177.545 81.815 177.775 ;
        RECT 81.600 177.390 81.740 177.545 ;
        RECT 81.970 177.530 82.290 177.790 ;
        RECT 82.890 177.530 83.210 177.790 ;
        RECT 84.820 177.775 84.960 177.930 ;
        RECT 88.870 177.930 93.240 178.070 ;
        RECT 88.870 177.870 89.190 177.930 ;
        RECT 85.650 177.775 85.970 177.800 ;
        RECT 93.100 177.775 93.240 177.930 ;
        RECT 94.940 177.930 97.470 178.070 ;
        RECT 84.285 177.545 84.575 177.775 ;
        RECT 84.745 177.545 85.035 177.775 ;
        RECT 85.590 177.545 85.970 177.775 ;
        RECT 86.175 177.730 86.465 177.775 ;
        RECT 86.175 177.590 86.800 177.730 ;
        RECT 87.925 177.700 88.215 177.755 ;
        RECT 86.175 177.545 86.465 177.590 ;
        RECT 83.810 177.390 84.130 177.450 ;
        RECT 78.840 177.250 79.440 177.390 ;
        RECT 81.600 177.250 84.130 177.390 ;
        RECT 84.360 177.390 84.500 177.545 ;
        RECT 85.650 177.540 85.970 177.545 ;
        RECT 84.360 177.250 85.420 177.390 ;
        RECT 64.045 177.205 64.335 177.250 ;
        RECT 73.245 177.205 73.535 177.250 ;
        RECT 74.610 177.190 74.930 177.250 ;
        RECT 77.845 177.205 78.135 177.250 ;
        RECT 79.300 177.110 79.440 177.250 ;
        RECT 83.810 177.190 84.130 177.250 ;
        RECT 85.280 177.110 85.420 177.250 ;
        RECT 86.660 177.110 86.800 177.590 ;
        RECT 87.580 177.560 88.215 177.700 ;
        RECT 62.650 177.050 62.970 177.110 ;
        RECT 62.280 176.910 62.970 177.050 ;
        RECT 62.650 176.850 62.970 176.910 ;
        RECT 65.425 177.050 65.715 177.095 ;
        RECT 65.870 177.050 66.190 177.110 ;
        RECT 65.425 176.910 66.190 177.050 ;
        RECT 65.425 176.865 65.715 176.910 ;
        RECT 65.870 176.850 66.190 176.910 ;
        RECT 72.325 177.050 72.615 177.095 ;
        RECT 73.690 177.050 74.010 177.110 ;
        RECT 72.325 176.910 74.010 177.050 ;
        RECT 72.325 176.865 72.615 176.910 ;
        RECT 73.690 176.850 74.010 176.910 ;
        RECT 75.070 176.850 75.390 177.110 ;
        RECT 75.530 177.050 75.850 177.110 ;
        RECT 76.925 177.050 77.215 177.095 ;
        RECT 78.750 177.050 79.070 177.110 ;
        RECT 75.530 176.910 79.070 177.050 ;
        RECT 75.530 176.850 75.850 176.910 ;
        RECT 76.925 176.865 77.215 176.910 ;
        RECT 78.750 176.850 79.070 176.910 ;
        RECT 79.210 176.850 79.530 177.110 ;
        RECT 80.130 177.050 80.450 177.110 ;
        RECT 80.605 177.050 80.895 177.095 ;
        RECT 80.130 176.910 80.895 177.050 ;
        RECT 80.130 176.850 80.450 176.910 ;
        RECT 80.605 176.865 80.895 176.910 ;
        RECT 82.905 177.050 83.195 177.095 ;
        RECT 84.270 177.050 84.590 177.110 ;
        RECT 82.905 176.910 84.590 177.050 ;
        RECT 82.905 176.865 83.195 176.910 ;
        RECT 84.270 176.850 84.590 176.910 ;
        RECT 85.190 176.850 85.510 177.110 ;
        RECT 86.570 176.850 86.890 177.110 ;
        RECT 87.580 177.050 87.720 177.560 ;
        RECT 87.925 177.525 88.215 177.560 ;
        RECT 88.425 177.545 88.715 177.775 ;
        RECT 89.805 177.730 90.095 177.775 ;
        RECT 89.805 177.590 91.860 177.730 ;
        RECT 89.805 177.545 90.095 177.590 ;
        RECT 88.500 177.390 88.640 177.545 ;
        RECT 91.720 177.450 91.860 177.590 ;
        RECT 93.025 177.545 93.315 177.775 ;
        RECT 93.490 177.545 93.780 177.775 ;
        RECT 93.930 177.730 94.250 177.790 ;
        RECT 94.940 177.775 95.080 177.930 ;
        RECT 97.150 177.870 97.470 177.930 ;
        RECT 97.610 177.870 97.930 178.130 ;
        RECT 99.005 178.070 99.295 178.115 ;
        RECT 98.160 177.930 99.295 178.070 ;
        RECT 94.865 177.730 95.155 177.775 ;
        RECT 93.930 177.590 95.155 177.730 ;
        RECT 88.500 177.250 90.020 177.390 ;
        RECT 89.880 177.110 90.020 177.250 ;
        RECT 91.170 177.190 91.490 177.450 ;
        RECT 91.630 177.190 91.950 177.450 ;
        RECT 92.090 177.390 92.410 177.450 ;
        RECT 93.565 177.390 93.705 177.545 ;
        RECT 93.930 177.530 94.250 177.590 ;
        RECT 94.865 177.545 95.155 177.590 ;
        RECT 95.770 177.730 96.090 177.790 ;
        RECT 96.705 177.730 96.995 177.775 ;
        RECT 98.160 177.730 98.300 177.930 ;
        RECT 99.005 177.885 99.295 177.930 ;
        RECT 101.305 178.070 101.595 178.115 ;
        RECT 114.645 178.070 114.935 178.115 ;
        RECT 119.245 178.070 119.535 178.115 ;
        RECT 123.830 178.070 124.150 178.130 ;
        RECT 101.305 177.930 114.935 178.070 ;
        RECT 101.305 177.885 101.595 177.930 ;
        RECT 114.645 177.885 114.935 177.930 ;
        RECT 115.180 177.930 124.150 178.070 ;
        RECT 95.770 177.590 96.995 177.730 ;
        RECT 95.770 177.530 96.090 177.590 ;
        RECT 96.705 177.545 96.995 177.590 ;
        RECT 97.700 177.590 98.300 177.730 ;
        RECT 97.700 177.450 97.840 177.590 ;
        RECT 98.530 177.530 98.850 177.790 ;
        RECT 99.465 177.545 99.755 177.775 ;
        RECT 97.150 177.390 97.470 177.450 ;
        RECT 92.090 177.250 97.470 177.390 ;
        RECT 92.090 177.190 92.410 177.250 ;
        RECT 97.150 177.190 97.470 177.250 ;
        RECT 97.610 177.190 97.930 177.450 ;
        RECT 88.870 177.050 89.190 177.110 ;
        RECT 87.580 176.910 89.190 177.050 ;
        RECT 88.870 176.850 89.190 176.910 ;
        RECT 89.790 176.850 90.110 177.110 ;
        RECT 90.250 176.850 90.570 177.110 ;
        RECT 94.390 177.050 94.710 177.110 ;
        RECT 99.540 177.050 99.680 177.545 ;
        RECT 99.910 177.530 100.230 177.790 ;
        RECT 102.210 177.730 102.530 177.790 ;
        RECT 102.680 177.730 102.970 177.775 ;
        RECT 102.210 177.590 102.970 177.730 ;
        RECT 102.210 177.530 102.530 177.590 ;
        RECT 102.680 177.545 102.970 177.590 ;
        RECT 103.130 177.530 103.450 177.790 ;
        RECT 103.590 177.530 103.910 177.790 ;
        RECT 104.525 177.730 104.815 177.775 ;
        RECT 108.650 177.730 108.970 177.790 ;
        RECT 104.525 177.590 108.970 177.730 ;
        RECT 104.525 177.545 104.815 177.590 ;
        RECT 108.650 177.530 108.970 177.590 ;
        RECT 111.410 177.730 111.730 177.790 ;
        RECT 114.185 177.730 114.475 177.775 ;
        RECT 115.180 177.730 115.320 177.930 ;
        RECT 119.245 177.885 119.535 177.930 ;
        RECT 123.830 177.870 124.150 177.930 ;
        RECT 136.710 177.870 137.030 178.130 ;
        RECT 111.410 177.590 115.320 177.730 ;
        RECT 111.410 177.530 111.730 177.590 ;
        RECT 114.185 177.545 114.475 177.590 ;
        RECT 115.550 177.530 115.870 177.790 ;
        RECT 116.470 177.530 116.790 177.790 ;
        RECT 117.850 177.530 118.170 177.790 ;
        RECT 118.310 177.530 118.630 177.790 ;
        RECT 118.770 177.530 119.090 177.790 ;
        RECT 119.690 177.530 120.010 177.790 ;
        RECT 120.610 177.530 120.930 177.790 ;
        RECT 122.450 177.530 122.770 177.790 ;
        RECT 130.270 177.730 130.590 177.790 ;
        RECT 132.125 177.730 132.415 177.775 ;
        RECT 130.270 177.590 132.415 177.730 ;
        RECT 130.270 177.530 130.590 177.590 ;
        RECT 132.125 177.545 132.415 177.590 ;
        RECT 133.030 177.730 133.350 177.790 ;
        RECT 133.965 177.730 134.255 177.775 ;
        RECT 133.030 177.590 134.255 177.730 ;
        RECT 133.030 177.530 133.350 177.590 ;
        RECT 133.965 177.545 134.255 177.590 ;
        RECT 137.170 177.530 137.490 177.790 ;
        RECT 103.220 177.390 103.360 177.530 ;
        RECT 113.250 177.390 113.570 177.450 ;
        RECT 103.220 177.250 113.570 177.390 ;
        RECT 113.250 177.190 113.570 177.250 ;
        RECT 113.725 177.390 114.015 177.435 ;
        RECT 116.930 177.390 117.250 177.450 ;
        RECT 118.405 177.390 118.545 177.530 ;
        RECT 113.725 177.250 118.545 177.390 ;
        RECT 113.725 177.205 114.015 177.250 ;
        RECT 116.930 177.190 117.250 177.250 ;
        RECT 118.310 177.050 118.630 177.110 ;
        RECT 94.390 176.910 118.630 177.050 ;
        RECT 94.390 176.850 94.710 176.910 ;
        RECT 118.310 176.850 118.630 176.910 ;
        RECT 133.490 177.050 133.810 177.110 ;
        RECT 134.885 177.050 135.175 177.095 ;
        RECT 136.250 177.050 136.570 177.110 ;
        RECT 133.490 176.910 136.570 177.050 ;
        RECT 133.490 176.850 133.810 176.910 ;
        RECT 134.885 176.865 135.175 176.910 ;
        RECT 136.250 176.850 136.570 176.910 ;
        RECT 27.160 176.230 139.860 176.710 ;
        RECT 45.630 176.030 45.950 176.090 ;
        RECT 47.485 176.030 47.775 176.075 ;
        RECT 55.290 176.030 55.610 176.090 ;
        RECT 45.630 175.890 55.610 176.030 ;
        RECT 45.630 175.830 45.950 175.890 ;
        RECT 47.485 175.845 47.775 175.890 ;
        RECT 55.290 175.830 55.610 175.890 ;
        RECT 59.430 175.830 59.750 176.090 ;
        RECT 61.270 176.030 61.590 176.090 ;
        RECT 62.205 176.030 62.495 176.075 ;
        RECT 68.630 176.030 68.950 176.090 ;
        RECT 61.270 175.890 62.495 176.030 ;
        RECT 61.270 175.830 61.590 175.890 ;
        RECT 62.205 175.845 62.495 175.890 ;
        RECT 66.420 175.890 68.950 176.030 ;
        RECT 41.490 175.490 41.810 175.750 ;
        RECT 44.710 175.690 45.030 175.750 ;
        RECT 45.185 175.690 45.475 175.735 ;
        RECT 44.710 175.550 45.475 175.690 ;
        RECT 44.710 175.490 45.030 175.550 ;
        RECT 45.185 175.505 45.475 175.550 ;
        RECT 49.770 175.490 50.090 175.750 ;
        RECT 50.690 175.490 51.010 175.750 ;
        RECT 59.520 175.690 59.660 175.830 ;
        RECT 64.045 175.690 64.335 175.735 ;
        RECT 64.490 175.690 64.810 175.750 ;
        RECT 59.520 175.550 61.960 175.690 ;
        RECT 42.870 175.350 43.190 175.410 ;
        RECT 44.265 175.350 44.555 175.395 ;
        RECT 48.390 175.350 48.710 175.410 ;
        RECT 50.230 175.350 50.550 175.410 ;
        RECT 42.870 175.210 48.710 175.350 ;
        RECT 42.870 175.150 43.190 175.210 ;
        RECT 44.265 175.165 44.555 175.210 ;
        RECT 48.390 175.150 48.710 175.210 ;
        RECT 48.940 175.210 50.550 175.350 ;
        RECT 43.805 175.010 44.095 175.055 ;
        RECT 48.940 175.010 49.080 175.210 ;
        RECT 50.230 175.150 50.550 175.210 ;
        RECT 58.050 175.350 58.370 175.410 ;
        RECT 58.985 175.350 59.275 175.395 ;
        RECT 58.050 175.210 59.275 175.350 ;
        RECT 58.050 175.150 58.370 175.210 ;
        RECT 58.985 175.165 59.275 175.210 ;
        RECT 59.430 175.350 59.750 175.410 ;
        RECT 59.905 175.350 60.195 175.395 ;
        RECT 59.430 175.210 60.195 175.350 ;
        RECT 59.430 175.150 59.750 175.210 ;
        RECT 59.905 175.165 60.195 175.210 ;
        RECT 60.350 175.150 60.670 175.410 ;
        RECT 61.270 175.150 61.590 175.410 ;
        RECT 61.820 175.395 61.960 175.550 ;
        RECT 62.280 175.550 64.810 175.690 ;
        RECT 61.745 175.165 62.035 175.395 ;
        RECT 43.805 174.870 49.080 175.010 ;
        RECT 49.325 175.010 49.615 175.055 ;
        RECT 49.770 175.010 50.090 175.070 ;
        RECT 62.280 175.010 62.420 175.550 ;
        RECT 64.045 175.505 64.335 175.550 ;
        RECT 64.490 175.490 64.810 175.550 ;
        RECT 64.965 175.690 65.255 175.735 ;
        RECT 66.420 175.690 66.560 175.890 ;
        RECT 68.630 175.830 68.950 175.890 ;
        RECT 69.565 176.030 69.855 176.075 ;
        RECT 70.010 176.030 70.330 176.090 ;
        RECT 69.565 175.890 70.330 176.030 ;
        RECT 69.565 175.845 69.855 175.890 ;
        RECT 70.010 175.830 70.330 175.890 ;
        RECT 70.930 176.030 71.250 176.090 ;
        RECT 76.450 176.030 76.770 176.090 ;
        RECT 70.930 175.890 76.770 176.030 ;
        RECT 70.930 175.830 71.250 175.890 ;
        RECT 76.450 175.830 76.770 175.890 ;
        RECT 77.830 176.030 78.150 176.090 ;
        RECT 80.225 176.030 80.515 176.075 ;
        RECT 77.830 175.890 80.515 176.030 ;
        RECT 77.830 175.830 78.150 175.890 ;
        RECT 80.225 175.845 80.515 175.890 ;
        RECT 84.270 176.030 84.590 176.090 ;
        RECT 91.170 176.030 91.490 176.090 ;
        RECT 94.390 176.030 94.710 176.090 ;
        RECT 99.450 176.030 99.770 176.090 ;
        RECT 84.270 175.890 90.940 176.030 ;
        RECT 84.270 175.830 84.590 175.890 ;
        RECT 64.965 175.550 66.560 175.690 ;
        RECT 64.965 175.505 65.255 175.550 ;
        RECT 62.665 175.165 62.955 175.395 ;
        RECT 49.325 174.870 50.090 175.010 ;
        RECT 43.805 174.825 44.095 174.870 ;
        RECT 49.325 174.825 49.615 174.870 ;
        RECT 49.770 174.810 50.090 174.870 ;
        RECT 59.520 174.870 62.420 175.010 ;
        RECT 42.870 174.470 43.190 174.730 ;
        RECT 59.520 174.715 59.660 174.870 ;
        RECT 59.445 174.485 59.735 174.715 ;
        RECT 61.730 174.670 62.050 174.730 ;
        RECT 62.740 174.670 62.880 175.165 ;
        RECT 63.125 174.670 63.415 174.715 ;
        RECT 61.730 174.530 63.415 174.670 ;
        RECT 61.730 174.470 62.050 174.530 ;
        RECT 63.125 174.485 63.415 174.530 ;
        RECT 60.825 174.330 61.115 174.375 ;
        RECT 65.040 174.330 65.180 175.505 ;
        RECT 67.710 175.490 68.030 175.750 ;
        RECT 70.100 175.690 70.240 175.830 ;
        RECT 73.230 175.690 73.550 175.750 ;
        RECT 70.100 175.550 73.550 175.690 ;
        RECT 73.230 175.490 73.550 175.550 ;
        RECT 75.070 175.690 75.390 175.750 ;
        RECT 75.545 175.690 75.835 175.735 ;
        RECT 79.225 175.690 79.515 175.735 ;
        RECT 88.885 175.690 89.175 175.735 ;
        RECT 90.250 175.690 90.570 175.750 ;
        RECT 75.070 175.550 75.835 175.690 ;
        RECT 75.070 175.490 75.390 175.550 ;
        RECT 75.545 175.505 75.835 175.550 ;
        RECT 77.000 175.550 79.515 175.690 ;
        RECT 77.000 175.410 77.140 175.550 ;
        RECT 79.225 175.505 79.515 175.550 ;
        RECT 84.360 175.550 90.570 175.690 ;
        RECT 90.800 175.690 90.940 175.890 ;
        RECT 91.170 175.890 99.770 176.030 ;
        RECT 91.170 175.830 91.490 175.890 ;
        RECT 94.390 175.830 94.710 175.890 ;
        RECT 99.450 175.830 99.770 175.890 ;
        RECT 99.910 176.030 100.230 176.090 ;
        RECT 101.305 176.030 101.595 176.075 ;
        RECT 99.910 175.890 101.595 176.030 ;
        RECT 99.910 175.830 100.230 175.890 ;
        RECT 101.305 175.845 101.595 175.890 ;
        RECT 101.750 176.030 102.070 176.090 ;
        RECT 132.570 176.030 132.890 176.090 ;
        RECT 101.750 175.890 118.310 176.030 ;
        RECT 101.750 175.830 102.070 175.890 ;
        RECT 104.970 175.690 105.290 175.750 ;
        RECT 105.445 175.690 105.735 175.735 ;
        RECT 90.800 175.550 103.820 175.690 ;
        RECT 65.870 175.150 66.190 175.410 ;
        RECT 67.265 175.165 67.555 175.395 ;
        RECT 67.340 175.010 67.480 175.165 ;
        RECT 68.630 175.150 68.950 175.410 ;
        RECT 70.930 175.350 71.250 175.410 ;
        RECT 71.405 175.350 71.695 175.395 ;
        RECT 70.930 175.210 71.695 175.350 ;
        RECT 70.930 175.150 71.250 175.210 ;
        RECT 71.405 175.165 71.695 175.210 ;
        RECT 72.310 175.350 72.630 175.410 ;
        RECT 72.785 175.350 73.075 175.395 ;
        RECT 74.165 175.350 74.455 175.395 ;
        RECT 72.310 175.210 74.455 175.350 ;
        RECT 72.310 175.150 72.630 175.210 ;
        RECT 72.785 175.165 73.075 175.210 ;
        RECT 74.165 175.165 74.455 175.210 ;
        RECT 76.910 175.150 77.230 175.410 ;
        RECT 78.750 175.350 79.070 175.410 ;
        RECT 81.525 175.350 81.815 175.395 ;
        RECT 78.750 175.210 81.815 175.350 ;
        RECT 78.750 175.150 79.070 175.210 ;
        RECT 81.525 175.165 81.815 175.210 ;
        RECT 83.350 175.150 83.670 175.410 ;
        RECT 70.010 175.010 70.330 175.070 ;
        RECT 67.340 174.870 70.330 175.010 ;
        RECT 70.010 174.810 70.330 174.870 ;
        RECT 70.470 175.010 70.790 175.070 ;
        RECT 75.530 175.010 75.850 175.070 ;
        RECT 76.005 175.010 76.295 175.055 ;
        RECT 84.360 175.010 84.500 175.550 ;
        RECT 88.885 175.505 89.175 175.550 ;
        RECT 90.250 175.490 90.570 175.550 ;
        RECT 84.730 175.150 85.050 175.410 ;
        RECT 85.210 175.165 85.500 175.395 ;
        RECT 86.125 175.350 86.415 175.395 ;
        RECT 85.740 175.210 86.415 175.350 ;
        RECT 70.470 174.870 76.295 175.010 ;
        RECT 70.470 174.810 70.790 174.870 ;
        RECT 75.530 174.810 75.850 174.870 ;
        RECT 76.005 174.825 76.295 174.870 ;
        RECT 77.920 174.870 84.500 175.010 ;
        RECT 65.410 174.670 65.730 174.730 ;
        RECT 69.550 174.670 69.870 174.730 ;
        RECT 73.705 174.670 73.995 174.715 ;
        RECT 77.370 174.670 77.690 174.730 ;
        RECT 77.920 174.715 78.060 174.870 ;
        RECT 65.410 174.530 72.995 174.670 ;
        RECT 65.410 174.470 65.730 174.530 ;
        RECT 69.550 174.470 69.870 174.530 ;
        RECT 60.825 174.190 65.180 174.330 ;
        RECT 60.825 174.145 61.115 174.190 ;
        RECT 66.790 174.130 67.110 174.390 ;
        RECT 70.930 174.130 71.250 174.390 ;
        RECT 71.390 174.330 71.710 174.390 ;
        RECT 72.325 174.330 72.615 174.375 ;
        RECT 71.390 174.190 72.615 174.330 ;
        RECT 72.855 174.330 72.995 174.530 ;
        RECT 73.705 174.530 77.690 174.670 ;
        RECT 73.705 174.485 73.995 174.530 ;
        RECT 77.370 174.470 77.690 174.530 ;
        RECT 77.845 174.485 78.135 174.715 ;
        RECT 81.065 174.670 81.355 174.715 ;
        RECT 81.970 174.670 82.290 174.730 ;
        RECT 81.065 174.530 82.290 174.670 ;
        RECT 81.065 174.485 81.355 174.530 ;
        RECT 81.970 174.470 82.290 174.530 ;
        RECT 82.445 174.670 82.735 174.715 ;
        RECT 82.890 174.670 83.210 174.730 ;
        RECT 85.280 174.670 85.420 175.165 ;
        RECT 82.445 174.530 83.210 174.670 ;
        RECT 82.445 174.485 82.735 174.530 ;
        RECT 82.890 174.470 83.210 174.530 ;
        RECT 83.670 174.530 85.420 174.670 ;
        RECT 75.545 174.330 75.835 174.375 ;
        RECT 72.855 174.190 75.835 174.330 ;
        RECT 71.390 174.130 71.710 174.190 ;
        RECT 72.325 174.145 72.615 174.190 ;
        RECT 75.545 174.145 75.835 174.190 ;
        RECT 76.450 174.330 76.770 174.390 ;
        RECT 80.145 174.330 80.435 174.375 ;
        RECT 76.450 174.190 80.435 174.330 ;
        RECT 76.450 174.130 76.770 174.190 ;
        RECT 80.145 174.145 80.435 174.190 ;
        RECT 80.590 174.330 80.910 174.390 ;
        RECT 83.670 174.330 83.810 174.530 ;
        RECT 80.590 174.190 83.810 174.330 ;
        RECT 80.590 174.130 80.910 174.190 ;
        RECT 84.270 174.130 84.590 174.390 ;
        RECT 84.730 174.330 85.050 174.390 ;
        RECT 85.740 174.330 85.880 175.210 ;
        RECT 86.125 175.165 86.415 175.210 ;
        RECT 86.585 175.165 86.875 175.395 ;
        RECT 87.275 175.350 87.565 175.395 ;
        RECT 87.275 175.210 88.180 175.350 ;
        RECT 87.275 175.165 87.565 175.210 ;
        RECT 86.660 175.010 86.800 175.165 ;
        RECT 88.040 175.010 88.180 175.210 ;
        RECT 88.410 175.150 88.730 175.410 ;
        RECT 89.805 175.165 90.095 175.395 ;
        RECT 89.330 175.010 89.650 175.070 ;
        RECT 86.660 174.870 87.260 175.010 ;
        RECT 88.040 174.870 89.650 175.010 ;
        RECT 87.120 174.730 87.260 174.870 ;
        RECT 89.330 174.810 89.650 174.870 ;
        RECT 87.030 174.470 87.350 174.730 ;
        RECT 87.950 174.470 88.270 174.730 ;
        RECT 89.880 174.670 90.020 175.165 ;
        RECT 91.170 175.150 91.490 175.410 ;
        RECT 92.105 175.165 92.395 175.395 ;
        RECT 92.180 175.010 92.320 175.165 ;
        RECT 92.550 175.150 92.870 175.410 ;
        RECT 93.470 175.150 93.790 175.410 ;
        RECT 94.405 175.350 94.695 175.395 ;
        RECT 94.850 175.350 95.170 175.410 ;
        RECT 94.405 175.210 95.170 175.350 ;
        RECT 94.405 175.165 94.695 175.210 ;
        RECT 94.850 175.150 95.170 175.210 ;
        RECT 95.770 175.150 96.090 175.410 ;
        RECT 96.230 175.150 96.550 175.410 ;
        RECT 97.150 175.350 97.470 175.410 ;
        RECT 97.625 175.350 97.915 175.395 ;
        RECT 97.150 175.210 97.915 175.350 ;
        RECT 97.150 175.150 97.470 175.210 ;
        RECT 97.625 175.165 97.915 175.210 ;
        RECT 99.450 175.150 99.770 175.410 ;
        RECT 101.750 175.350 102.070 175.410 ;
        RECT 103.680 175.395 103.820 175.550 ;
        RECT 104.970 175.550 109.800 175.690 ;
        RECT 104.970 175.490 105.290 175.550 ;
        RECT 105.445 175.505 105.735 175.550 ;
        RECT 109.660 175.410 109.800 175.550 ;
        RECT 111.410 175.490 111.730 175.750 ;
        RECT 118.170 175.690 118.310 175.890 ;
        RECT 118.680 175.890 132.890 176.030 ;
        RECT 118.680 175.690 118.820 175.890 ;
        RECT 132.570 175.830 132.890 175.890 ;
        RECT 136.710 175.830 137.030 176.090 ;
        RECT 137.185 175.845 137.475 176.075 ;
        RECT 118.170 175.550 118.820 175.690 ;
        RECT 129.365 175.690 129.655 175.735 ;
        RECT 135.790 175.690 136.110 175.750 ;
        RECT 137.260 175.690 137.400 175.845 ;
        RECT 129.365 175.550 132.110 175.690 ;
        RECT 129.365 175.505 129.655 175.550 ;
        RECT 100.920 175.210 102.070 175.350 ;
        RECT 100.920 175.010 101.060 175.210 ;
        RECT 101.750 175.150 102.070 175.210 ;
        RECT 103.605 175.165 103.895 175.395 ;
        RECT 106.810 175.350 107.130 175.410 ;
        RECT 109.125 175.350 109.415 175.395 ;
        RECT 106.810 175.210 109.415 175.350 ;
        RECT 106.810 175.150 107.130 175.210 ;
        RECT 109.125 175.165 109.415 175.210 ;
        RECT 109.570 175.150 109.890 175.410 ;
        RECT 110.505 175.165 110.795 175.395 ;
        RECT 92.180 174.870 99.220 175.010 ;
        RECT 93.930 174.670 94.250 174.730 ;
        RECT 89.880 174.530 94.250 174.670 ;
        RECT 93.930 174.470 94.250 174.530 ;
        RECT 94.850 174.670 95.170 174.730 ;
        RECT 95.325 174.670 95.615 174.715 ;
        RECT 94.850 174.530 95.615 174.670 ;
        RECT 94.850 174.470 95.170 174.530 ;
        RECT 95.325 174.485 95.615 174.530 ;
        RECT 84.730 174.190 85.880 174.330 ;
        RECT 86.570 174.330 86.890 174.390 ;
        RECT 89.805 174.330 90.095 174.375 ;
        RECT 86.570 174.190 90.095 174.330 ;
        RECT 84.730 174.130 85.050 174.190 ;
        RECT 86.570 174.130 86.890 174.190 ;
        RECT 89.805 174.145 90.095 174.190 ;
        RECT 90.725 174.330 91.015 174.375 ;
        RECT 98.530 174.330 98.850 174.390 ;
        RECT 90.725 174.190 98.850 174.330 ;
        RECT 99.080 174.330 99.220 174.870 ;
        RECT 99.540 174.870 101.060 175.010 ;
        RECT 99.540 174.715 99.680 174.870 ;
        RECT 102.210 174.810 102.530 175.070 ;
        RECT 102.670 174.810 102.990 175.070 ;
        RECT 103.130 174.810 103.450 175.070 ;
        RECT 110.580 175.010 110.720 175.165 ;
        RECT 110.950 175.150 111.270 175.410 ;
        RECT 111.870 175.350 112.190 175.410 ;
        RECT 120.150 175.350 120.470 175.410 ;
        RECT 111.870 175.210 120.470 175.350 ;
        RECT 111.870 175.150 112.190 175.210 ;
        RECT 120.150 175.150 120.470 175.210 ;
        RECT 130.270 175.350 130.590 175.410 ;
        RECT 130.745 175.350 131.035 175.395 ;
        RECT 130.270 175.210 131.035 175.350 ;
        RECT 131.970 175.350 132.110 175.550 ;
        RECT 135.790 175.550 137.400 175.690 ;
        RECT 135.790 175.490 136.110 175.550 ;
        RECT 133.045 175.350 133.335 175.395 ;
        RECT 131.970 175.210 133.335 175.350 ;
        RECT 130.270 175.150 130.590 175.210 ;
        RECT 130.745 175.165 131.035 175.210 ;
        RECT 133.045 175.165 133.335 175.210 ;
        RECT 133.490 175.350 133.810 175.410 ;
        RECT 133.965 175.350 134.255 175.395 ;
        RECT 133.490 175.210 134.255 175.350 ;
        RECT 133.490 175.150 133.810 175.210 ;
        RECT 133.965 175.165 134.255 175.210 ;
        RECT 136.250 175.150 136.570 175.410 ;
        RECT 137.630 175.010 137.950 175.070 ;
        RECT 110.580 174.870 137.950 175.010 ;
        RECT 137.630 174.810 137.950 174.870 ;
        RECT 138.105 174.825 138.395 175.055 ;
        RECT 99.465 174.485 99.755 174.715 ;
        RECT 99.910 174.670 100.230 174.730 ;
        RECT 111.870 174.670 112.190 174.730 ;
        RECT 99.910 174.530 112.190 174.670 ;
        RECT 99.910 174.470 100.230 174.530 ;
        RECT 111.870 174.470 112.190 174.530 ;
        RECT 122.925 174.670 123.215 174.715 ;
        RECT 130.730 174.670 131.050 174.730 ;
        RECT 122.925 174.530 131.050 174.670 ;
        RECT 122.925 174.485 123.215 174.530 ;
        RECT 130.730 174.470 131.050 174.530 ;
        RECT 136.250 174.670 136.570 174.730 ;
        RECT 138.180 174.670 138.320 174.825 ;
        RECT 136.250 174.530 138.320 174.670 ;
        RECT 136.250 174.470 136.570 174.530 ;
        RECT 107.270 174.330 107.590 174.390 ;
        RECT 99.080 174.190 107.590 174.330 ;
        RECT 90.725 174.145 91.015 174.190 ;
        RECT 98.530 174.130 98.850 174.190 ;
        RECT 107.270 174.130 107.590 174.190 ;
        RECT 108.190 174.130 108.510 174.390 ;
        RECT 134.870 174.330 135.190 174.390 ;
        RECT 136.725 174.330 137.015 174.375 ;
        RECT 134.870 174.190 137.015 174.330 ;
        RECT 134.870 174.130 135.190 174.190 ;
        RECT 136.725 174.145 137.015 174.190 ;
        RECT 27.160 173.510 139.860 173.990 ;
        RECT 62.665 173.310 62.955 173.355 ;
        RECT 63.110 173.310 63.430 173.370 ;
        RECT 62.665 173.170 63.430 173.310 ;
        RECT 62.665 173.125 62.955 173.170 ;
        RECT 63.110 173.110 63.430 173.170 ;
        RECT 63.570 173.310 63.890 173.370 ;
        RECT 65.410 173.310 65.730 173.370 ;
        RECT 67.710 173.310 68.030 173.370 ;
        RECT 63.570 173.170 65.730 173.310 ;
        RECT 63.570 173.110 63.890 173.170 ;
        RECT 65.410 173.110 65.730 173.170 ;
        RECT 65.960 173.170 68.030 173.310 ;
        RECT 60.350 172.970 60.670 173.030 ;
        RECT 64.490 172.970 64.810 173.030 ;
        RECT 65.960 172.970 66.100 173.170 ;
        RECT 67.710 173.110 68.030 173.170 ;
        RECT 69.105 173.310 69.395 173.355 ;
        RECT 71.850 173.310 72.170 173.370 ;
        RECT 69.105 173.170 72.170 173.310 ;
        RECT 69.105 173.125 69.395 173.170 ;
        RECT 71.850 173.110 72.170 173.170 ;
        RECT 73.230 173.310 73.550 173.370 ;
        RECT 74.165 173.310 74.455 173.355 ;
        RECT 73.230 173.170 74.455 173.310 ;
        RECT 73.230 173.110 73.550 173.170 ;
        RECT 74.165 173.125 74.455 173.170 ;
        RECT 76.005 173.310 76.295 173.355 ;
        RECT 76.450 173.310 76.770 173.370 ;
        RECT 76.005 173.170 76.770 173.310 ;
        RECT 76.005 173.125 76.295 173.170 ;
        RECT 76.450 173.110 76.770 173.170 ;
        RECT 78.290 173.310 78.610 173.370 ;
        RECT 78.765 173.310 79.055 173.355 ;
        RECT 78.290 173.170 79.055 173.310 ;
        RECT 78.290 173.110 78.610 173.170 ;
        RECT 78.765 173.125 79.055 173.170 ;
        RECT 79.210 173.310 79.530 173.370 ;
        RECT 82.890 173.310 83.210 173.370 ;
        RECT 79.210 173.170 83.210 173.310 ;
        RECT 79.210 173.110 79.530 173.170 ;
        RECT 82.890 173.110 83.210 173.170 ;
        RECT 83.825 173.310 84.115 173.355 ;
        RECT 85.650 173.310 85.970 173.370 ;
        RECT 83.825 173.170 85.970 173.310 ;
        RECT 83.825 173.125 84.115 173.170 ;
        RECT 85.650 173.110 85.970 173.170 ;
        RECT 87.030 173.310 87.350 173.370 ;
        RECT 88.410 173.310 88.730 173.370 ;
        RECT 87.030 173.170 88.730 173.310 ;
        RECT 87.030 173.110 87.350 173.170 ;
        RECT 88.410 173.110 88.730 173.170 ;
        RECT 88.885 173.125 89.175 173.355 ;
        RECT 60.350 172.830 64.260 172.970 ;
        RECT 60.350 172.770 60.670 172.830 ;
        RECT 58.050 172.630 58.370 172.690 ;
        RECT 59.430 172.630 59.750 172.690 ;
        RECT 58.050 172.490 61.500 172.630 ;
        RECT 58.050 172.430 58.370 172.490 ;
        RECT 58.600 172.335 58.740 172.490 ;
        RECT 59.430 172.430 59.750 172.490 ;
        RECT 58.525 172.105 58.815 172.335 ;
        RECT 59.890 172.090 60.210 172.350 ;
        RECT 61.360 172.335 61.500 172.490 ;
        RECT 61.285 172.290 61.575 172.335 ;
        RECT 63.110 172.290 63.430 172.350 ;
        RECT 64.120 172.340 64.260 172.830 ;
        RECT 64.490 172.830 66.100 172.970 ;
        RECT 66.330 172.970 66.650 173.030 ;
        RECT 75.085 172.970 75.375 173.015 ;
        RECT 80.605 172.970 80.895 173.015 ;
        RECT 84.730 172.970 85.050 173.030 ;
        RECT 88.960 172.970 89.100 173.125 ;
        RECT 89.790 173.110 90.110 173.370 ;
        RECT 93.470 173.310 93.790 173.370 ;
        RECT 97.610 173.310 97.930 173.370 ;
        RECT 90.800 173.170 93.240 173.310 ;
        RECT 66.330 172.830 71.160 172.970 ;
        RECT 64.490 172.770 64.810 172.830 ;
        RECT 66.330 172.770 66.650 172.830 ;
        RECT 66.805 172.630 67.095 172.675 ;
        RECT 70.010 172.630 70.330 172.690 ;
        RECT 65.040 172.490 70.330 172.630 ;
        RECT 65.040 172.340 65.180 172.490 ;
        RECT 66.805 172.445 67.095 172.490 ;
        RECT 70.010 172.430 70.330 172.490 ;
        RECT 64.120 172.335 65.180 172.340 ;
        RECT 61.285 172.150 63.430 172.290 ;
        RECT 61.285 172.105 61.575 172.150 ;
        RECT 63.110 172.090 63.430 172.150 ;
        RECT 64.045 172.200 65.180 172.335 ;
        RECT 64.045 172.105 64.335 172.200 ;
        RECT 66.330 172.090 66.650 172.350 ;
        RECT 67.710 172.090 68.030 172.350 ;
        RECT 68.185 172.105 68.475 172.335 ;
        RECT 68.630 172.290 68.950 172.350 ;
        RECT 71.020 172.335 71.160 172.830 ;
        RECT 75.085 172.830 80.440 172.970 ;
        RECT 75.085 172.785 75.375 172.830 ;
        RECT 72.325 172.630 72.615 172.675 ;
        RECT 74.150 172.630 74.470 172.690 ;
        RECT 80.300 172.630 80.440 172.830 ;
        RECT 80.605 172.830 85.050 172.970 ;
        RECT 80.605 172.785 80.895 172.830 ;
        RECT 84.730 172.770 85.050 172.830 ;
        RECT 85.280 172.830 89.100 172.970 ;
        RECT 89.330 172.970 89.650 173.030 ;
        RECT 90.800 173.015 90.940 173.170 ;
        RECT 90.725 172.970 91.015 173.015 ;
        RECT 89.330 172.830 91.015 172.970 ;
        RECT 93.100 172.970 93.240 173.170 ;
        RECT 93.470 173.170 97.930 173.310 ;
        RECT 93.470 173.110 93.790 173.170 ;
        RECT 97.610 173.110 97.930 173.170 ;
        RECT 98.530 173.310 98.850 173.370 ;
        RECT 101.750 173.310 102.070 173.370 ;
        RECT 98.530 173.170 102.070 173.310 ;
        RECT 98.530 173.110 98.850 173.170 ;
        RECT 101.750 173.110 102.070 173.170 ;
        RECT 107.270 173.310 107.590 173.370 ;
        RECT 116.470 173.310 116.790 173.370 ;
        RECT 124.305 173.310 124.595 173.355 ;
        RECT 107.270 173.170 124.595 173.310 ;
        RECT 107.270 173.110 107.590 173.170 ;
        RECT 116.470 173.110 116.790 173.170 ;
        RECT 124.305 173.125 124.595 173.170 ;
        RECT 134.410 173.110 134.730 173.370 ;
        RECT 96.690 172.970 97.010 173.030 ;
        RECT 98.990 172.970 99.310 173.030 ;
        RECT 93.100 172.830 94.620 172.970 ;
        RECT 82.445 172.630 82.735 172.675 ;
        RECT 85.280 172.630 85.420 172.830 ;
        RECT 89.330 172.770 89.650 172.830 ;
        RECT 90.725 172.785 91.015 172.830 ;
        RECT 92.105 172.630 92.395 172.675 ;
        RECT 72.325 172.490 74.470 172.630 ;
        RECT 72.325 172.445 72.615 172.490 ;
        RECT 74.150 172.430 74.470 172.490 ;
        RECT 74.700 172.490 79.900 172.630 ;
        RECT 80.300 172.490 85.420 172.630 ;
        RECT 86.200 172.490 88.180 172.630 ;
        RECT 69.565 172.290 69.855 172.335 ;
        RECT 68.630 172.150 69.855 172.290 ;
        RECT 61.745 171.950 62.035 171.995 ;
        RECT 59.060 171.810 62.035 171.950 ;
        RECT 59.060 171.670 59.200 171.810 ;
        RECT 61.745 171.765 62.035 171.810 ;
        RECT 62.190 171.950 62.510 172.010 ;
        RECT 62.665 171.950 62.955 171.995 ;
        RECT 62.190 171.810 62.955 171.950 ;
        RECT 62.190 171.750 62.510 171.810 ;
        RECT 62.665 171.765 62.955 171.810 ;
        RECT 64.490 171.750 64.810 172.010 ;
        RECT 65.425 171.950 65.715 171.995 ;
        RECT 67.800 171.950 67.940 172.090 ;
        RECT 65.425 171.810 67.940 171.950 ;
        RECT 68.260 171.950 68.400 172.105 ;
        RECT 68.630 172.090 68.950 172.150 ;
        RECT 69.565 172.105 69.855 172.150 ;
        RECT 70.945 172.105 71.235 172.335 ;
        RECT 71.390 172.090 71.710 172.350 ;
        RECT 71.850 172.290 72.170 172.350 ;
        RECT 74.700 172.290 74.840 172.490 ;
        RECT 71.850 172.150 74.840 172.290 ;
        RECT 71.850 172.090 72.170 172.150 ;
        RECT 75.545 172.105 75.835 172.335 ;
        RECT 76.450 172.290 76.770 172.350 ;
        RECT 76.925 172.290 77.215 172.335 ;
        RECT 76.450 172.150 77.215 172.290 ;
        RECT 71.480 171.950 71.620 172.090 ;
        RECT 68.260 171.810 71.620 171.950 ;
        RECT 65.425 171.765 65.715 171.810 ;
        RECT 73.245 171.765 73.535 171.995 ;
        RECT 74.325 171.950 74.615 171.995 ;
        RECT 75.070 171.950 75.390 172.010 ;
        RECT 74.325 171.810 75.390 171.950 ;
        RECT 74.325 171.765 74.615 171.810 ;
        RECT 58.970 171.410 59.290 171.670 ;
        RECT 60.825 171.610 61.115 171.655 ;
        RECT 70.470 171.610 70.790 171.670 ;
        RECT 72.770 171.610 73.090 171.670 ;
        RECT 73.320 171.610 73.460 171.765 ;
        RECT 75.070 171.750 75.390 171.810 ;
        RECT 75.620 171.610 75.760 172.105 ;
        RECT 76.450 172.090 76.770 172.150 ;
        RECT 76.925 172.105 77.215 172.150 ;
        RECT 77.370 172.090 77.690 172.350 ;
        RECT 78.765 172.290 79.055 172.335 ;
        RECT 77.920 172.150 79.055 172.290 ;
        RECT 60.825 171.470 75.760 171.610 ;
        RECT 77.920 171.610 78.060 172.150 ;
        RECT 78.765 172.105 79.055 172.150 ;
        RECT 79.210 172.090 79.530 172.350 ;
        RECT 79.760 172.290 79.900 172.490 ;
        RECT 82.445 172.445 82.735 172.490 ;
        RECT 80.590 172.290 80.910 172.350 ;
        RECT 81.525 172.290 81.815 172.335 ;
        RECT 79.760 172.150 81.815 172.290 ;
        RECT 80.590 172.090 80.910 172.150 ;
        RECT 81.525 172.105 81.815 172.150 ;
        RECT 81.970 172.090 82.290 172.350 ;
        RECT 82.890 172.090 83.210 172.350 ;
        RECT 84.360 172.335 84.500 172.490 ;
        RECT 84.285 172.105 84.575 172.335 ;
        RECT 85.205 172.290 85.495 172.335 ;
        RECT 86.200 172.290 86.340 172.490 ;
        RECT 88.040 172.335 88.180 172.490 ;
        RECT 88.500 172.490 92.395 172.630 ;
        RECT 88.500 172.350 88.640 172.490 ;
        RECT 92.105 172.445 92.395 172.490 ;
        RECT 93.485 172.630 93.775 172.675 ;
        RECT 93.930 172.630 94.250 172.690 ;
        RECT 94.480 172.675 94.620 172.830 ;
        RECT 96.690 172.830 99.310 172.970 ;
        RECT 96.690 172.770 97.010 172.830 ;
        RECT 98.990 172.770 99.310 172.830 ;
        RECT 99.450 172.970 99.770 173.030 ;
        RECT 102.670 172.970 102.990 173.030 ;
        RECT 106.810 172.970 107.130 173.030 ;
        RECT 99.450 172.830 107.130 172.970 ;
        RECT 99.450 172.770 99.770 172.830 ;
        RECT 102.670 172.770 102.990 172.830 ;
        RECT 106.810 172.770 107.130 172.830 ;
        RECT 93.485 172.490 94.250 172.630 ;
        RECT 93.485 172.445 93.775 172.490 ;
        RECT 85.205 172.150 86.340 172.290 ;
        RECT 85.205 172.105 85.495 172.150 ;
        RECT 86.585 172.105 86.875 172.335 ;
        RECT 87.965 172.105 88.255 172.335 ;
        RECT 78.305 171.950 78.595 171.995 ;
        RECT 82.060 171.950 82.200 172.090 ;
        RECT 85.280 171.950 85.420 172.105 ;
        RECT 78.305 171.810 81.740 171.950 ;
        RECT 82.060 171.810 85.420 171.950 ;
        RECT 86.110 171.950 86.430 172.010 ;
        RECT 86.660 171.950 86.800 172.105 ;
        RECT 88.410 172.090 88.730 172.350 ;
        RECT 91.185 172.180 91.475 172.335 ;
        RECT 90.340 172.105 91.475 172.180 ;
        RECT 90.340 172.040 91.400 172.105 ;
        RECT 92.550 172.090 92.870 172.350 ;
        RECT 93.560 172.290 93.700 172.445 ;
        RECT 93.930 172.430 94.250 172.490 ;
        RECT 94.405 172.630 94.695 172.675 ;
        RECT 95.310 172.630 95.630 172.690 ;
        RECT 94.405 172.490 95.630 172.630 ;
        RECT 94.405 172.445 94.695 172.490 ;
        RECT 95.310 172.430 95.630 172.490 ;
        RECT 96.230 172.630 96.550 172.690 ;
        RECT 97.610 172.630 97.930 172.690 ;
        RECT 110.030 172.630 110.350 172.690 ;
        RECT 96.230 172.490 109.800 172.630 ;
        RECT 96.230 172.430 96.550 172.490 ;
        RECT 97.610 172.430 97.930 172.490 ;
        RECT 93.100 172.150 93.700 172.290 ;
        RECT 94.865 172.290 95.155 172.335 ;
        RECT 97.150 172.290 97.470 172.350 ;
        RECT 94.865 172.150 97.470 172.290 ;
        RECT 89.330 171.950 89.650 172.010 ;
        RECT 90.340 171.950 90.480 172.040 ;
        RECT 93.100 171.950 93.240 172.150 ;
        RECT 94.865 172.105 95.155 172.150 ;
        RECT 97.150 172.090 97.470 172.150 ;
        RECT 99.450 172.090 99.770 172.350 ;
        RECT 99.910 172.090 100.230 172.350 ;
        RECT 109.660 172.290 109.800 172.490 ;
        RECT 110.030 172.490 111.180 172.630 ;
        RECT 110.030 172.430 110.350 172.490 ;
        RECT 110.490 172.290 110.810 172.350 ;
        RECT 111.040 172.335 111.180 172.490 ;
        RECT 109.660 172.150 110.810 172.290 ;
        RECT 110.490 172.090 110.810 172.150 ;
        RECT 110.965 172.105 111.255 172.335 ;
        RECT 126.130 172.290 126.450 172.350 ;
        RECT 127.065 172.290 127.355 172.335 ;
        RECT 126.130 172.150 127.355 172.290 ;
        RECT 126.130 172.090 126.450 172.150 ;
        RECT 127.065 172.105 127.355 172.150 ;
        RECT 132.570 172.290 132.890 172.350 ;
        RECT 137.185 172.290 137.475 172.335 ;
        RECT 132.570 172.150 137.475 172.290 ;
        RECT 132.570 172.090 132.890 172.150 ;
        RECT 137.185 172.105 137.475 172.150 ;
        RECT 98.070 171.950 98.390 172.010 ;
        RECT 86.110 171.810 89.100 171.950 ;
        RECT 78.305 171.765 78.595 171.810 ;
        RECT 80.590 171.610 80.910 171.670 ;
        RECT 77.920 171.470 80.910 171.610 ;
        RECT 81.600 171.610 81.740 171.810 ;
        RECT 86.110 171.750 86.430 171.810 ;
        RECT 87.030 171.610 87.350 171.670 ;
        RECT 81.600 171.470 87.350 171.610 ;
        RECT 60.825 171.425 61.115 171.470 ;
        RECT 70.470 171.410 70.790 171.470 ;
        RECT 72.770 171.410 73.090 171.470 ;
        RECT 80.590 171.410 80.910 171.470 ;
        RECT 87.030 171.410 87.350 171.470 ;
        RECT 87.505 171.610 87.795 171.655 ;
        RECT 88.410 171.610 88.730 171.670 ;
        RECT 87.505 171.470 88.730 171.610 ;
        RECT 88.960 171.610 89.100 171.810 ;
        RECT 89.330 171.810 90.480 171.950 ;
        RECT 91.720 171.810 93.240 171.950 ;
        RECT 93.560 171.810 98.390 171.950 ;
        RECT 89.330 171.750 89.650 171.810 ;
        RECT 91.720 171.610 91.860 171.810 ;
        RECT 92.090 171.610 92.410 171.670 ;
        RECT 88.960 171.470 92.410 171.610 ;
        RECT 87.505 171.425 87.795 171.470 ;
        RECT 88.410 171.410 88.730 171.470 ;
        RECT 92.090 171.410 92.410 171.470 ;
        RECT 92.550 171.610 92.870 171.670 ;
        RECT 93.560 171.610 93.700 171.810 ;
        RECT 98.070 171.750 98.390 171.810 ;
        RECT 98.530 171.750 98.850 172.010 ;
        RECT 101.305 171.950 101.595 171.995 ;
        RECT 99.540 171.810 101.595 171.950 ;
        RECT 99.540 171.670 99.680 171.810 ;
        RECT 101.305 171.765 101.595 171.810 ;
        RECT 92.550 171.470 93.700 171.610 ;
        RECT 93.945 171.610 94.235 171.655 ;
        RECT 94.390 171.610 94.710 171.670 ;
        RECT 93.945 171.470 94.710 171.610 ;
        RECT 92.550 171.410 92.870 171.470 ;
        RECT 93.945 171.425 94.235 171.470 ;
        RECT 94.390 171.410 94.710 171.470 ;
        RECT 95.785 171.610 96.075 171.655 ;
        RECT 96.690 171.610 97.010 171.670 ;
        RECT 95.785 171.470 97.010 171.610 ;
        RECT 95.785 171.425 96.075 171.470 ;
        RECT 96.690 171.410 97.010 171.470 ;
        RECT 99.450 171.410 99.770 171.670 ;
        RECT 100.370 171.410 100.690 171.670 ;
        RECT 101.380 171.610 101.520 171.765 ;
        RECT 101.750 171.750 102.070 172.010 ;
        RECT 107.270 171.950 107.590 172.010 ;
        RECT 102.300 171.810 107.590 171.950 ;
        RECT 102.300 171.610 102.440 171.810 ;
        RECT 107.270 171.750 107.590 171.810 ;
        RECT 107.730 171.950 108.050 172.010 ;
        RECT 117.865 171.950 118.155 171.995 ;
        RECT 107.730 171.810 118.155 171.950 ;
        RECT 107.730 171.750 108.050 171.810 ;
        RECT 117.865 171.765 118.155 171.810 ;
        RECT 126.590 171.950 126.910 172.010 ;
        RECT 131.190 171.950 131.510 172.010 ;
        RECT 136.265 171.950 136.555 171.995 ;
        RECT 126.590 171.810 136.555 171.950 ;
        RECT 126.590 171.750 126.910 171.810 ;
        RECT 131.190 171.750 131.510 171.810 ;
        RECT 136.265 171.765 136.555 171.810 ;
        RECT 101.380 171.470 102.440 171.610 ;
        RECT 102.670 171.610 102.990 171.670 ;
        RECT 108.205 171.610 108.495 171.655 ;
        RECT 111.410 171.610 111.730 171.670 ;
        RECT 102.670 171.470 111.730 171.610 ;
        RECT 102.670 171.410 102.990 171.470 ;
        RECT 108.205 171.425 108.495 171.470 ;
        RECT 111.410 171.410 111.730 171.470 ;
        RECT 125.210 171.610 125.530 171.670 ;
        RECT 138.105 171.610 138.395 171.655 ;
        RECT 125.210 171.470 138.395 171.610 ;
        RECT 125.210 171.410 125.530 171.470 ;
        RECT 138.105 171.425 138.395 171.470 ;
        RECT 27.160 170.790 139.860 171.270 ;
        RECT 55.290 170.590 55.610 170.650 ;
        RECT 63.585 170.590 63.875 170.635 ;
        RECT 64.490 170.590 64.810 170.650 ;
        RECT 71.850 170.590 72.170 170.650 ;
        RECT 55.290 170.450 61.960 170.590 ;
        RECT 55.290 170.390 55.610 170.450 ;
        RECT 61.820 170.250 61.960 170.450 ;
        RECT 63.585 170.450 64.810 170.590 ;
        RECT 63.585 170.405 63.875 170.450 ;
        RECT 64.490 170.390 64.810 170.450 ;
        RECT 65.040 170.450 72.170 170.590 ;
        RECT 65.040 170.250 65.180 170.450 ;
        RECT 71.850 170.390 72.170 170.450 ;
        RECT 72.770 170.590 73.090 170.650 ;
        RECT 75.070 170.635 75.390 170.650 ;
        RECT 72.770 170.450 74.380 170.590 ;
        RECT 72.770 170.390 73.090 170.450 ;
        RECT 56.300 170.110 61.500 170.250 ;
        RECT 61.820 170.110 65.180 170.250 ;
        RECT 65.410 170.250 65.730 170.310 ;
        RECT 69.550 170.250 69.870 170.310 ;
        RECT 74.240 170.295 74.380 170.450 ;
        RECT 75.070 170.405 75.455 170.635 ;
        RECT 75.070 170.390 75.390 170.405 ;
        RECT 78.290 170.390 78.610 170.650 ;
        RECT 82.445 170.590 82.735 170.635 ;
        RECT 91.170 170.590 91.490 170.650 ;
        RECT 82.445 170.450 91.490 170.590 ;
        RECT 82.445 170.405 82.735 170.450 ;
        RECT 91.170 170.390 91.490 170.450 ;
        RECT 91.630 170.390 91.950 170.650 ;
        RECT 92.090 170.390 92.410 170.650 ;
        RECT 94.390 170.590 94.710 170.650 ;
        RECT 96.230 170.590 96.550 170.650 ;
        RECT 110.030 170.590 110.350 170.650 ;
        RECT 117.405 170.590 117.695 170.635 ;
        RECT 133.950 170.590 134.270 170.650 ;
        RECT 94.390 170.450 95.080 170.590 ;
        RECT 94.390 170.390 94.710 170.450 ;
        RECT 65.410 170.110 68.860 170.250 ;
        RECT 49.310 169.910 49.630 169.970 ;
        RECT 56.300 169.955 56.440 170.110 ;
        RECT 56.225 169.910 56.515 169.955 ;
        RECT 49.310 169.770 56.515 169.910 ;
        RECT 49.310 169.710 49.630 169.770 ;
        RECT 56.225 169.725 56.515 169.770 ;
        RECT 57.130 169.710 57.450 169.970 ;
        RECT 57.605 169.725 57.895 169.955 ;
        RECT 57.680 169.570 57.820 169.725 ;
        RECT 58.510 169.710 58.830 169.970 ;
        RECT 61.360 169.955 61.500 170.110 ;
        RECT 65.410 170.050 65.730 170.110 ;
        RECT 68.720 169.970 68.860 170.110 ;
        RECT 69.550 170.110 73.920 170.250 ;
        RECT 69.550 170.050 69.870 170.110 ;
        RECT 61.285 169.725 61.575 169.955 ;
        RECT 62.650 169.910 62.970 169.970 ;
        RECT 64.505 169.910 64.795 169.955 ;
        RECT 62.650 169.770 64.795 169.910 ;
        RECT 62.650 169.710 62.970 169.770 ;
        RECT 64.505 169.725 64.795 169.770 ;
        RECT 66.330 169.910 66.650 169.970 ;
        RECT 67.250 169.910 67.570 169.970 ;
        RECT 66.330 169.770 67.570 169.910 ;
        RECT 66.330 169.710 66.650 169.770 ;
        RECT 67.250 169.710 67.570 169.770 ;
        RECT 68.630 169.710 68.950 169.970 ;
        RECT 69.090 169.910 69.410 169.970 ;
        RECT 70.025 169.910 70.315 169.955 ;
        RECT 69.090 169.770 70.315 169.910 ;
        RECT 69.090 169.710 69.410 169.770 ;
        RECT 70.025 169.725 70.315 169.770 ;
        RECT 70.945 169.725 71.235 169.955 ;
        RECT 72.785 169.725 73.075 169.955 ;
        RECT 73.780 169.910 73.920 170.110 ;
        RECT 74.165 170.065 74.455 170.295 ;
        RECT 76.465 170.250 76.755 170.295 ;
        RECT 74.700 170.110 76.755 170.250 ;
        RECT 74.700 169.910 74.840 170.110 ;
        RECT 76.465 170.065 76.755 170.110 ;
        RECT 76.910 170.250 77.230 170.310 ;
        RECT 77.465 170.250 77.755 170.295 ;
        RECT 76.910 170.110 77.755 170.250 ;
        RECT 78.380 170.250 78.520 170.390 ;
        RECT 81.970 170.250 82.290 170.310 ;
        RECT 83.365 170.250 83.655 170.295 ;
        RECT 78.380 170.110 80.360 170.250 ;
        RECT 76.910 170.050 77.230 170.110 ;
        RECT 77.465 170.065 77.755 170.110 ;
        RECT 79.210 169.910 79.530 169.970 ;
        RECT 80.220 169.955 80.360 170.110 ;
        RECT 81.970 170.110 83.655 170.250 ;
        RECT 81.970 170.050 82.290 170.110 ;
        RECT 83.365 170.065 83.655 170.110 ;
        RECT 83.810 170.250 84.130 170.310 ;
        RECT 86.585 170.250 86.875 170.295 ;
        RECT 83.810 170.110 86.875 170.250 ;
        RECT 83.810 170.050 84.130 170.110 ;
        RECT 86.585 170.065 86.875 170.110 ;
        RECT 88.410 170.250 88.730 170.310 ;
        RECT 88.410 170.110 90.940 170.250 ;
        RECT 88.410 170.050 88.730 170.110 ;
        RECT 73.780 169.770 74.840 169.910 ;
        RECT 76.080 169.770 79.530 169.910 ;
        RECT 58.050 169.570 58.370 169.630 ;
        RECT 62.740 169.570 62.880 169.710 ;
        RECT 55.380 169.430 62.880 169.570 ;
        RECT 65.410 169.570 65.730 169.630 ;
        RECT 66.805 169.570 67.095 169.615 ;
        RECT 69.550 169.570 69.870 169.630 ;
        RECT 71.020 169.570 71.160 169.725 ;
        RECT 65.410 169.430 71.160 169.570 ;
        RECT 72.860 169.570 73.000 169.725 ;
        RECT 74.150 169.570 74.470 169.630 ;
        RECT 72.860 169.430 74.470 169.570 ;
        RECT 55.380 169.275 55.520 169.430 ;
        RECT 58.050 169.370 58.370 169.430 ;
        RECT 65.410 169.370 65.730 169.430 ;
        RECT 66.805 169.385 67.095 169.430 ;
        RECT 69.550 169.370 69.870 169.430 ;
        RECT 74.150 169.370 74.470 169.430 ;
        RECT 55.305 169.045 55.595 169.275 ;
        RECT 59.430 169.030 59.750 169.290 ;
        RECT 62.205 169.230 62.495 169.275 ;
        RECT 69.090 169.230 69.410 169.290 ;
        RECT 62.205 169.090 69.410 169.230 ;
        RECT 62.205 169.045 62.495 169.090 ;
        RECT 69.090 169.030 69.410 169.090 ;
        RECT 70.010 169.030 70.330 169.290 ;
        RECT 76.080 169.275 76.220 169.770 ;
        RECT 79.210 169.710 79.530 169.770 ;
        RECT 80.145 169.725 80.435 169.955 ;
        RECT 81.050 169.910 81.370 169.970 ;
        RECT 81.525 169.910 81.815 169.955 ;
        RECT 81.050 169.770 81.815 169.910 ;
        RECT 81.050 169.710 81.370 169.770 ;
        RECT 81.525 169.725 81.815 169.770 ;
        RECT 85.190 169.710 85.510 169.970 ;
        RECT 86.110 169.710 86.430 169.970 ;
        RECT 87.505 169.725 87.795 169.955 ;
        RECT 87.580 169.570 87.720 169.725 ;
        RECT 89.790 169.710 90.110 169.970 ;
        RECT 90.800 169.910 90.940 170.110 ;
        RECT 92.550 170.050 92.870 170.310 ;
        RECT 94.940 169.955 95.080 170.450 ;
        RECT 96.230 170.450 134.270 170.590 ;
        RECT 96.230 170.390 96.550 170.450 ;
        RECT 110.030 170.390 110.350 170.450 ;
        RECT 117.405 170.405 117.695 170.450 ;
        RECT 133.950 170.390 134.270 170.450 ;
        RECT 134.425 170.590 134.715 170.635 ;
        RECT 135.790 170.590 136.110 170.650 ;
        RECT 134.425 170.450 136.110 170.590 ;
        RECT 134.425 170.405 134.715 170.450 ;
        RECT 135.790 170.390 136.110 170.450 ;
        RECT 137.170 170.590 137.490 170.650 ;
        RECT 137.645 170.590 137.935 170.635 ;
        RECT 137.170 170.450 137.935 170.590 ;
        RECT 137.170 170.390 137.490 170.450 ;
        RECT 137.645 170.405 137.935 170.450 ;
        RECT 95.310 170.050 95.630 170.310 ;
        RECT 104.970 170.250 105.290 170.310 ;
        RECT 97.700 170.110 105.290 170.250 ;
        RECT 93.100 169.910 93.730 169.930 ;
        RECT 93.945 169.910 94.235 169.955 ;
        RECT 90.800 169.790 94.235 169.910 ;
        RECT 90.800 169.770 93.240 169.790 ;
        RECT 93.590 169.770 94.235 169.790 ;
        RECT 93.945 169.725 94.235 169.770 ;
        RECT 94.865 169.725 95.155 169.955 ;
        RECT 95.400 169.910 95.540 170.050 ;
        RECT 95.785 169.910 96.075 169.955 ;
        RECT 95.400 169.770 96.075 169.910 ;
        RECT 95.785 169.725 96.075 169.770 ;
        RECT 96.230 169.710 96.550 169.970 ;
        RECT 97.700 169.955 97.840 170.110 ;
        RECT 104.970 170.050 105.290 170.110 ;
        RECT 106.350 170.050 106.670 170.310 ;
        RECT 110.965 170.250 111.255 170.295 ;
        RECT 116.010 170.250 116.330 170.310 ;
        RECT 110.965 170.110 116.330 170.250 ;
        RECT 110.965 170.065 111.255 170.110 ;
        RECT 116.010 170.050 116.330 170.110 ;
        RECT 128.905 170.250 129.195 170.295 ;
        RECT 130.730 170.250 131.050 170.310 ;
        RECT 128.905 170.110 131.050 170.250 ;
        RECT 128.905 170.065 129.195 170.110 ;
        RECT 130.730 170.050 131.050 170.110 ;
        RECT 97.625 169.725 97.915 169.955 ;
        RECT 98.070 169.910 98.390 169.970 ;
        RECT 100.845 169.910 101.135 169.955 ;
        RECT 98.070 169.770 101.135 169.910 ;
        RECT 98.070 169.710 98.390 169.770 ;
        RECT 100.845 169.725 101.135 169.770 ;
        RECT 101.290 169.910 101.610 169.970 ;
        RECT 102.225 169.910 102.515 169.955 ;
        RECT 101.290 169.770 102.515 169.910 ;
        RECT 87.950 169.570 88.270 169.630 ;
        RECT 79.300 169.430 88.270 169.570 ;
        RECT 79.300 169.290 79.440 169.430 ;
        RECT 87.950 169.370 88.270 169.430 ;
        RECT 88.410 169.370 88.730 169.630 ;
        RECT 88.885 169.570 89.175 169.615 ;
        RECT 89.330 169.570 89.650 169.630 ;
        RECT 88.885 169.430 89.650 169.570 ;
        RECT 88.885 169.385 89.175 169.430 ;
        RECT 89.330 169.370 89.650 169.430 ;
        RECT 93.485 169.385 93.775 169.615 ;
        RECT 95.325 169.570 95.615 169.615 ;
        RECT 96.320 169.570 96.460 169.710 ;
        RECT 95.325 169.430 96.460 169.570 ;
        RECT 95.325 169.385 95.615 169.430 ;
        RECT 96.705 169.385 96.995 169.615 ;
        RECT 76.005 169.045 76.295 169.275 ;
        RECT 79.210 169.030 79.530 169.290 ;
        RECT 80.590 169.230 80.910 169.290 ;
        RECT 93.560 169.230 93.700 169.385 ;
        RECT 80.590 169.090 93.700 169.230 ;
        RECT 93.935 169.230 94.255 169.290 ;
        RECT 95.400 169.230 95.540 169.385 ;
        RECT 93.935 169.090 95.540 169.230 ;
        RECT 80.590 169.030 80.910 169.090 ;
        RECT 93.935 169.030 94.255 169.090 ;
        RECT 96.230 169.030 96.550 169.290 ;
        RECT 25.390 168.890 25.710 168.950 ;
        RECT 28.625 168.890 28.915 168.935 ;
        RECT 25.390 168.750 28.915 168.890 ;
        RECT 25.390 168.690 25.710 168.750 ;
        RECT 28.625 168.705 28.915 168.750 ;
        RECT 57.130 168.890 57.450 168.950 ;
        RECT 64.505 168.890 64.795 168.935 ;
        RECT 64.950 168.890 65.270 168.950 ;
        RECT 57.130 168.750 65.270 168.890 ;
        RECT 57.130 168.690 57.450 168.750 ;
        RECT 64.505 168.705 64.795 168.750 ;
        RECT 64.950 168.690 65.270 168.750 ;
        RECT 71.850 168.890 72.170 168.950 ;
        RECT 73.705 168.890 73.995 168.935 ;
        RECT 71.850 168.750 73.995 168.890 ;
        RECT 71.850 168.690 72.170 168.750 ;
        RECT 73.705 168.705 73.995 168.750 ;
        RECT 75.070 168.690 75.390 168.950 ;
        RECT 75.530 168.890 75.850 168.950 ;
        RECT 76.910 168.890 77.230 168.950 ;
        RECT 75.530 168.750 77.230 168.890 ;
        RECT 75.530 168.690 75.850 168.750 ;
        RECT 76.910 168.690 77.230 168.750 ;
        RECT 77.370 168.690 77.690 168.950 ;
        RECT 83.825 168.890 84.115 168.935 ;
        RECT 91.170 168.890 91.490 168.950 ;
        RECT 83.825 168.750 91.490 168.890 ;
        RECT 83.825 168.705 84.115 168.750 ;
        RECT 91.170 168.690 91.490 168.750 ;
        RECT 93.010 168.890 93.330 168.950 ;
        RECT 96.780 168.890 96.920 169.385 ;
        RECT 98.530 169.370 98.850 169.630 ;
        RECT 99.450 169.370 99.770 169.630 ;
        RECT 100.385 169.385 100.675 169.615 ;
        RECT 93.010 168.750 96.920 168.890 ;
        RECT 98.070 168.890 98.390 168.950 ;
        RECT 100.460 168.890 100.600 169.385 ;
        RECT 98.070 168.750 100.600 168.890 ;
        RECT 100.920 168.890 101.060 169.725 ;
        RECT 101.290 169.710 101.610 169.770 ;
        RECT 102.225 169.725 102.515 169.770 ;
        RECT 102.300 169.570 102.440 169.725 ;
        RECT 103.130 169.710 103.450 169.970 ;
        RECT 103.590 169.910 103.910 169.970 ;
        RECT 107.285 169.910 107.575 169.955 ;
        RECT 103.590 169.770 107.575 169.910 ;
        RECT 103.590 169.710 103.910 169.770 ;
        RECT 107.285 169.725 107.575 169.770 ;
        RECT 108.650 169.910 108.970 169.970 ;
        RECT 120.165 169.910 120.455 169.955 ;
        RECT 108.650 169.770 120.455 169.910 ;
        RECT 108.650 169.710 108.970 169.770 ;
        RECT 120.165 169.725 120.455 169.770 ;
        RECT 125.670 169.910 125.990 169.970 ;
        RECT 132.585 169.910 132.875 169.955 ;
        RECT 125.670 169.770 132.875 169.910 ;
        RECT 125.670 169.710 125.990 169.770 ;
        RECT 132.585 169.725 132.875 169.770 ;
        RECT 133.965 169.910 134.255 169.955 ;
        RECT 136.725 169.910 137.015 169.955 ;
        RECT 133.965 169.770 137.015 169.910 ;
        RECT 133.965 169.725 134.255 169.770 ;
        RECT 136.725 169.725 137.015 169.770 ;
        RECT 105.905 169.570 106.195 169.615 ;
        RECT 102.300 169.430 106.195 169.570 ;
        RECT 105.905 169.385 106.195 169.430 ;
        RECT 106.810 169.570 107.130 169.630 ;
        RECT 130.745 169.570 131.035 169.615 ;
        RECT 106.810 169.430 131.035 169.570 ;
        RECT 106.810 169.370 107.130 169.430 ;
        RECT 130.745 169.385 131.035 169.430 ;
        RECT 133.030 169.370 133.350 169.630 ;
        RECT 136.250 169.370 136.570 169.630 ;
        RECT 104.065 169.230 104.355 169.275 ;
        RECT 117.850 169.230 118.170 169.290 ;
        RECT 104.065 169.090 118.170 169.230 ;
        RECT 104.065 169.045 104.355 169.090 ;
        RECT 117.850 169.030 118.170 169.090 ;
        RECT 103.590 168.890 103.910 168.950 ;
        RECT 114.170 168.890 114.490 168.950 ;
        RECT 100.920 168.750 114.490 168.890 ;
        RECT 93.010 168.690 93.330 168.750 ;
        RECT 98.070 168.690 98.390 168.750 ;
        RECT 103.590 168.690 103.910 168.750 ;
        RECT 114.170 168.690 114.490 168.750 ;
        RECT 27.160 168.070 139.860 168.550 ;
        RECT 42.425 167.870 42.715 167.915 ;
        RECT 44.710 167.870 45.030 167.930 ;
        RECT 42.425 167.730 45.030 167.870 ;
        RECT 42.425 167.685 42.715 167.730 ;
        RECT 44.710 167.670 45.030 167.730 ;
        RECT 45.645 167.870 45.935 167.915 ;
        RECT 49.310 167.870 49.630 167.930 ;
        RECT 45.645 167.730 49.630 167.870 ;
        RECT 45.645 167.685 45.935 167.730 ;
        RECT 49.310 167.670 49.630 167.730 ;
        RECT 50.690 167.870 51.010 167.930 ;
        RECT 51.165 167.870 51.455 167.915 ;
        RECT 50.690 167.730 51.455 167.870 ;
        RECT 50.690 167.670 51.010 167.730 ;
        RECT 51.165 167.685 51.455 167.730 ;
        RECT 52.545 167.870 52.835 167.915 ;
        RECT 52.545 167.730 58.280 167.870 ;
        RECT 52.545 167.685 52.835 167.730 ;
        RECT 48.865 167.530 49.155 167.575 ;
        RECT 58.140 167.530 58.280 167.730 ;
        RECT 58.510 167.670 58.830 167.930 ;
        RECT 58.970 167.870 59.290 167.930 ;
        RECT 59.445 167.870 59.735 167.915 ;
        RECT 58.970 167.730 59.735 167.870 ;
        RECT 58.970 167.670 59.290 167.730 ;
        RECT 59.445 167.685 59.735 167.730 ;
        RECT 59.890 167.870 60.210 167.930 ;
        RECT 60.365 167.870 60.655 167.915 ;
        RECT 65.410 167.870 65.730 167.930 ;
        RECT 59.890 167.730 65.730 167.870 ;
        RECT 59.890 167.670 60.210 167.730 ;
        RECT 60.365 167.685 60.655 167.730 ;
        RECT 65.410 167.670 65.730 167.730 ;
        RECT 71.405 167.870 71.695 167.915 ;
        RECT 77.830 167.870 78.150 167.930 ;
        RECT 71.405 167.730 78.150 167.870 ;
        RECT 71.405 167.685 71.695 167.730 ;
        RECT 77.830 167.670 78.150 167.730 ;
        RECT 78.305 167.870 78.595 167.915 ;
        RECT 86.110 167.870 86.430 167.930 ;
        RECT 78.305 167.730 86.430 167.870 ;
        RECT 78.305 167.685 78.595 167.730 ;
        RECT 86.110 167.670 86.430 167.730 ;
        RECT 90.265 167.870 90.555 167.915 ;
        RECT 94.865 167.870 95.155 167.915 ;
        RECT 95.770 167.870 96.090 167.930 ;
        RECT 98.070 167.870 98.390 167.930 ;
        RECT 90.265 167.730 94.620 167.870 ;
        RECT 90.265 167.685 90.555 167.730 ;
        RECT 48.865 167.390 56.900 167.530 ;
        RECT 58.140 167.390 67.940 167.530 ;
        RECT 48.865 167.345 49.155 167.390 ;
        RECT 56.210 166.990 56.530 167.250 ;
        RECT 56.760 167.190 56.900 167.390 ;
        RECT 66.330 167.190 66.650 167.250 ;
        RECT 56.760 167.050 66.650 167.190 ;
        RECT 41.030 166.850 41.350 166.910 ;
        RECT 41.505 166.850 41.795 166.895 ;
        RECT 41.030 166.710 41.795 166.850 ;
        RECT 41.030 166.650 41.350 166.710 ;
        RECT 41.505 166.665 41.795 166.710 ;
        RECT 44.250 166.850 44.570 166.910 ;
        RECT 44.725 166.850 45.015 166.895 ;
        RECT 44.250 166.710 45.015 166.850 ;
        RECT 44.250 166.650 44.570 166.710 ;
        RECT 44.725 166.665 45.015 166.710 ;
        RECT 47.930 166.650 48.250 166.910 ;
        RECT 50.245 166.850 50.535 166.895 ;
        RECT 50.690 166.850 51.010 166.910 ;
        RECT 50.245 166.710 51.010 166.850 ;
        RECT 50.245 166.665 50.535 166.710 ;
        RECT 50.690 166.650 51.010 166.710 ;
        RECT 51.625 166.665 51.915 166.895 ;
        RECT 51.700 166.510 51.840 166.665 ;
        RECT 54.370 166.650 54.690 166.910 ;
        RECT 56.760 166.895 56.900 167.050 ;
        RECT 66.330 166.990 66.650 167.050 ;
        RECT 67.800 166.910 67.940 167.390 ;
        RECT 72.770 167.330 73.090 167.590 ;
        RECT 75.545 167.345 75.835 167.575 ;
        RECT 76.925 167.530 77.215 167.575 ;
        RECT 82.890 167.530 83.210 167.590 ;
        RECT 76.925 167.390 83.210 167.530 ;
        RECT 76.925 167.345 77.215 167.390 ;
        RECT 75.070 167.190 75.390 167.250 ;
        RECT 72.860 167.050 75.390 167.190 ;
        RECT 75.620 167.190 75.760 167.345 ;
        RECT 82.890 167.330 83.210 167.390 ;
        RECT 88.425 167.530 88.715 167.575 ;
        RECT 94.480 167.530 94.620 167.730 ;
        RECT 94.865 167.730 98.390 167.870 ;
        RECT 94.865 167.685 95.155 167.730 ;
        RECT 95.770 167.670 96.090 167.730 ;
        RECT 98.070 167.670 98.390 167.730 ;
        RECT 100.830 167.870 101.150 167.930 ;
        RECT 109.110 167.870 109.430 167.930 ;
        RECT 111.425 167.870 111.715 167.915 ;
        RECT 100.830 167.730 107.960 167.870 ;
        RECT 100.830 167.670 101.150 167.730 ;
        RECT 95.310 167.530 95.630 167.590 ;
        RECT 88.425 167.390 94.340 167.530 ;
        RECT 94.480 167.390 95.630 167.530 ;
        RECT 88.425 167.345 88.715 167.390 ;
        RECT 92.550 167.190 92.870 167.250 ;
        RECT 75.620 167.050 92.870 167.190 ;
        RECT 94.200 167.190 94.340 167.390 ;
        RECT 95.310 167.330 95.630 167.390 ;
        RECT 97.150 167.530 97.470 167.590 ;
        RECT 107.285 167.530 107.575 167.575 ;
        RECT 97.150 167.390 107.575 167.530 ;
        RECT 97.150 167.330 97.470 167.390 ;
        RECT 107.285 167.345 107.575 167.390 ;
        RECT 101.750 167.190 102.070 167.250 ;
        RECT 94.200 167.050 102.070 167.190 ;
        RECT 56.685 166.665 56.975 166.895 ;
        RECT 58.050 166.850 58.370 166.910 ;
        RECT 58.525 166.850 58.815 166.895 ;
        RECT 58.050 166.710 58.815 166.850 ;
        RECT 58.050 166.650 58.370 166.710 ;
        RECT 58.525 166.665 58.815 166.710 ;
        RECT 61.285 166.850 61.575 166.895 ;
        RECT 61.285 166.710 62.880 166.850 ;
        RECT 61.285 166.665 61.575 166.710 ;
        RECT 57.130 166.510 57.450 166.570 ;
        RECT 62.205 166.510 62.495 166.555 ;
        RECT 51.700 166.370 56.900 166.510 ;
        RECT 55.290 165.970 55.610 166.230 ;
        RECT 56.760 166.170 56.900 166.370 ;
        RECT 57.130 166.370 62.495 166.510 ;
        RECT 57.130 166.310 57.450 166.370 ;
        RECT 62.205 166.325 62.495 166.370 ;
        RECT 62.740 166.230 62.880 166.710 ;
        RECT 64.490 166.650 64.810 166.910 ;
        RECT 67.710 166.650 68.030 166.910 ;
        RECT 69.090 166.650 69.410 166.910 ;
        RECT 70.470 166.650 70.790 166.910 ;
        RECT 70.930 166.850 71.250 166.910 ;
        RECT 72.860 166.895 73.000 167.050 ;
        RECT 75.070 166.990 75.390 167.050 ;
        RECT 92.550 166.990 92.870 167.050 ;
        RECT 101.750 166.990 102.070 167.050 ;
        RECT 102.210 166.990 102.530 167.250 ;
        RECT 104.970 167.190 105.290 167.250 ;
        RECT 103.220 167.050 105.290 167.190 ;
        RECT 107.820 167.190 107.960 167.730 ;
        RECT 109.110 167.730 111.715 167.870 ;
        RECT 109.110 167.670 109.430 167.730 ;
        RECT 111.425 167.685 111.715 167.730 ;
        RECT 113.710 167.670 114.030 167.930 ;
        RECT 114.170 167.870 114.490 167.930 ;
        RECT 128.905 167.870 129.195 167.915 ;
        RECT 114.170 167.730 129.195 167.870 ;
        RECT 114.170 167.670 114.490 167.730 ;
        RECT 128.905 167.685 129.195 167.730 ;
        RECT 133.030 167.870 133.350 167.930 ;
        RECT 136.265 167.870 136.555 167.915 ;
        RECT 133.030 167.730 136.555 167.870 ;
        RECT 133.030 167.670 133.350 167.730 ;
        RECT 136.265 167.685 136.555 167.730 ;
        RECT 110.965 167.530 111.255 167.575 ;
        RECT 114.630 167.530 114.950 167.590 ;
        RECT 110.965 167.390 114.950 167.530 ;
        RECT 110.965 167.345 111.255 167.390 ;
        RECT 114.630 167.330 114.950 167.390 ;
        RECT 118.785 167.345 119.075 167.575 ;
        RECT 119.690 167.530 120.010 167.590 ;
        RECT 137.645 167.530 137.935 167.575 ;
        RECT 119.690 167.390 137.935 167.530 ;
        RECT 118.860 167.190 119.000 167.345 ;
        RECT 119.690 167.330 120.010 167.390 ;
        RECT 137.645 167.345 137.935 167.390 ;
        RECT 107.820 167.050 119.000 167.190 ;
        RECT 128.445 167.190 128.735 167.235 ;
        RECT 130.270 167.190 130.590 167.250 ;
        RECT 128.445 167.050 130.590 167.190 ;
        RECT 71.865 166.850 72.155 166.895 ;
        RECT 70.930 166.710 72.155 166.850 ;
        RECT 70.930 166.650 71.250 166.710 ;
        RECT 71.865 166.665 72.155 166.710 ;
        RECT 72.785 166.665 73.075 166.895 ;
        RECT 73.230 166.650 73.550 166.910 ;
        RECT 74.625 166.665 74.915 166.895 ;
        RECT 64.950 166.510 65.270 166.570 ;
        RECT 74.700 166.510 74.840 166.665 ;
        RECT 75.990 166.650 76.310 166.910 ;
        RECT 77.370 166.650 77.690 166.910 ;
        RECT 80.130 166.650 80.450 166.910 ;
        RECT 81.510 166.850 81.830 166.910 ;
        RECT 83.365 166.850 83.655 166.895 ;
        RECT 81.510 166.710 83.655 166.850 ;
        RECT 81.510 166.650 81.830 166.710 ;
        RECT 83.365 166.665 83.655 166.710 ;
        RECT 83.810 166.650 84.130 166.910 ;
        RECT 84.730 166.895 85.050 166.910 ;
        RECT 84.595 166.665 85.050 166.895 ;
        RECT 84.730 166.650 85.050 166.665 ;
        RECT 85.190 166.850 85.510 166.910 ;
        RECT 86.125 166.850 86.415 166.895 ;
        RECT 85.190 166.710 86.415 166.850 ;
        RECT 85.190 166.650 85.510 166.710 ;
        RECT 86.125 166.665 86.415 166.710 ;
        RECT 86.570 166.650 86.890 166.910 ;
        RECT 87.490 166.650 87.810 166.910 ;
        RECT 88.885 166.665 89.175 166.895 ;
        RECT 89.330 166.850 89.650 166.910 ;
        RECT 100.370 166.850 100.690 166.910 ;
        RECT 89.330 166.710 100.690 166.850 ;
        RECT 88.960 166.510 89.100 166.665 ;
        RECT 89.330 166.650 89.650 166.710 ;
        RECT 100.370 166.650 100.690 166.710 ;
        RECT 101.305 166.850 101.595 166.895 ;
        RECT 102.670 166.850 102.990 166.910 ;
        RECT 103.220 166.895 103.360 167.050 ;
        RECT 104.970 166.990 105.290 167.050 ;
        RECT 128.445 167.005 128.735 167.050 ;
        RECT 130.270 166.990 130.590 167.050 ;
        RECT 132.570 166.990 132.890 167.250 ;
        RECT 135.330 166.990 135.650 167.250 ;
        RECT 101.305 166.710 102.990 166.850 ;
        RECT 101.305 166.665 101.595 166.710 ;
        RECT 102.670 166.650 102.990 166.710 ;
        RECT 103.145 166.665 103.435 166.895 ;
        RECT 104.065 166.850 104.355 166.895 ;
        RECT 104.510 166.850 104.830 166.910 ;
        RECT 104.065 166.710 104.830 166.850 ;
        RECT 104.065 166.665 104.355 166.710 ;
        RECT 104.510 166.650 104.830 166.710 ;
        RECT 105.430 166.850 105.750 166.910 ;
        RECT 106.365 166.850 106.655 166.895 ;
        RECT 105.430 166.710 106.655 166.850 ;
        RECT 105.430 166.650 105.750 166.710 ;
        RECT 106.365 166.665 106.655 166.710 ;
        RECT 106.810 166.850 107.130 166.910 ;
        RECT 108.205 166.850 108.495 166.895 ;
        RECT 110.030 166.850 110.350 166.910 ;
        RECT 106.810 166.710 108.495 166.850 ;
        RECT 106.810 166.650 107.130 166.710 ;
        RECT 108.205 166.665 108.495 166.710 ;
        RECT 108.740 166.710 110.350 166.850 ;
        RECT 64.950 166.370 67.020 166.510 ;
        RECT 74.700 166.370 89.100 166.510 ;
        RECT 91.185 166.510 91.475 166.555 ;
        RECT 92.090 166.510 92.410 166.570 ;
        RECT 91.185 166.370 92.410 166.510 ;
        RECT 64.950 166.310 65.270 166.370 ;
        RECT 60.350 166.170 60.670 166.230 ;
        RECT 56.760 166.030 60.670 166.170 ;
        RECT 60.350 165.970 60.670 166.030 ;
        RECT 62.650 165.970 62.970 166.230 ;
        RECT 65.410 165.970 65.730 166.230 ;
        RECT 66.880 166.215 67.020 166.370 ;
        RECT 91.185 166.325 91.475 166.370 ;
        RECT 92.090 166.310 92.410 166.370 ;
        RECT 96.230 166.510 96.550 166.570 ;
        RECT 104.985 166.510 105.275 166.555 ;
        RECT 96.230 166.370 105.275 166.510 ;
        RECT 96.230 166.310 96.550 166.370 ;
        RECT 104.985 166.325 105.275 166.370 ;
        RECT 105.890 166.510 106.210 166.570 ;
        RECT 108.740 166.510 108.880 166.710 ;
        RECT 110.030 166.650 110.350 166.710 ;
        RECT 110.490 166.850 110.810 166.910 ;
        RECT 112.345 166.850 112.635 166.895 ;
        RECT 110.490 166.710 112.635 166.850 ;
        RECT 110.490 166.650 110.810 166.710 ;
        RECT 112.345 166.665 112.635 166.710 ;
        RECT 112.805 166.850 113.095 166.895 ;
        RECT 112.805 166.710 113.940 166.850 ;
        RECT 112.805 166.665 113.095 166.710 ;
        RECT 105.890 166.370 108.880 166.510 ;
        RECT 105.890 166.310 106.210 166.370 ;
        RECT 109.125 166.325 109.415 166.555 ;
        RECT 66.805 165.985 67.095 166.215 ;
        RECT 70.010 165.970 70.330 166.230 ;
        RECT 74.165 166.170 74.455 166.215 ;
        RECT 79.210 166.170 79.530 166.230 ;
        RECT 74.165 166.030 79.530 166.170 ;
        RECT 74.165 165.985 74.455 166.030 ;
        RECT 79.210 165.970 79.530 166.030 ;
        RECT 81.050 165.970 81.370 166.230 ;
        RECT 82.445 166.170 82.735 166.215 ;
        RECT 83.350 166.170 83.670 166.230 ;
        RECT 82.445 166.030 83.670 166.170 ;
        RECT 82.445 165.985 82.735 166.030 ;
        RECT 83.350 165.970 83.670 166.030 ;
        RECT 85.665 166.170 85.955 166.215 ;
        RECT 88.870 166.170 89.190 166.230 ;
        RECT 85.665 166.030 89.190 166.170 ;
        RECT 85.665 165.985 85.955 166.030 ;
        RECT 88.870 165.970 89.190 166.030 ;
        RECT 90.265 166.170 90.555 166.215 ;
        RECT 91.630 166.170 91.950 166.230 ;
        RECT 90.265 166.030 91.950 166.170 ;
        RECT 90.265 165.985 90.555 166.030 ;
        RECT 91.630 165.970 91.950 166.030 ;
        RECT 94.390 166.170 94.710 166.230 ;
        RECT 97.150 166.170 97.470 166.230 ;
        RECT 94.390 166.030 97.470 166.170 ;
        RECT 94.390 165.970 94.710 166.030 ;
        RECT 97.150 165.970 97.470 166.030 ;
        RECT 105.430 165.970 105.750 166.230 ;
        RECT 109.200 166.170 109.340 166.325 ;
        RECT 109.570 166.310 109.890 166.570 ;
        RECT 112.880 166.510 113.020 166.665 ;
        RECT 110.120 166.370 113.020 166.510 ;
        RECT 113.800 166.510 113.940 166.710 ;
        RECT 114.170 166.650 114.490 166.910 ;
        RECT 116.470 166.650 116.790 166.910 ;
        RECT 117.850 166.650 118.170 166.910 ;
        RECT 119.230 166.850 119.550 166.910 ;
        RECT 119.705 166.850 119.995 166.895 ;
        RECT 119.230 166.710 119.995 166.850 ;
        RECT 119.230 166.650 119.550 166.710 ;
        RECT 119.705 166.665 119.995 166.710 ;
        RECT 129.810 166.650 130.130 166.910 ;
        RECT 131.190 166.850 131.510 166.910 ;
        RECT 131.665 166.850 131.955 166.895 ;
        RECT 131.190 166.710 131.955 166.850 ;
        RECT 131.190 166.650 131.510 166.710 ;
        RECT 131.665 166.665 131.955 166.710 ;
        RECT 134.870 166.650 135.190 166.910 ;
        RECT 136.710 166.650 137.030 166.910 ;
        RECT 120.150 166.510 120.470 166.570 ;
        RECT 113.800 166.370 120.470 166.510 ;
        RECT 110.120 166.170 110.260 166.370 ;
        RECT 120.150 166.310 120.470 166.370 ;
        RECT 121.070 166.510 121.390 166.570 ;
        RECT 130.745 166.510 131.035 166.555 ;
        RECT 121.070 166.370 131.035 166.510 ;
        RECT 121.070 166.310 121.390 166.370 ;
        RECT 130.745 166.325 131.035 166.370 ;
        RECT 109.200 166.030 110.260 166.170 ;
        RECT 133.030 165.970 133.350 166.230 ;
        RECT 27.160 165.350 139.860 165.830 ;
        RECT 75.990 165.150 76.310 165.210 ;
        RECT 89.790 165.150 90.110 165.210 ;
        RECT 75.990 165.010 90.110 165.150 ;
        RECT 75.990 164.950 76.310 165.010 ;
        RECT 89.790 164.950 90.110 165.010 ;
        RECT 91.170 165.150 91.490 165.210 ;
        RECT 93.470 165.150 93.790 165.210 ;
        RECT 91.170 165.010 93.790 165.150 ;
        RECT 91.170 164.950 91.490 165.010 ;
        RECT 93.470 164.950 93.790 165.010 ;
        RECT 73.230 164.810 73.550 164.870 ;
        RECT 99.450 164.810 99.770 164.870 ;
        RECT 73.230 164.670 99.770 164.810 ;
        RECT 73.230 164.610 73.550 164.670 ;
        RECT 99.450 164.610 99.770 164.670 ;
        RECT 110.030 164.810 110.350 164.870 ;
        RECT 119.690 164.810 120.010 164.870 ;
        RECT 136.710 164.810 137.030 164.870 ;
        RECT 110.030 164.670 120.010 164.810 ;
        RECT 110.030 164.610 110.350 164.670 ;
        RECT 119.690 164.610 120.010 164.670 ;
        RECT 131.970 164.670 137.030 164.810 ;
        RECT 77.370 164.470 77.690 164.530 ;
        RECT 94.850 164.470 95.170 164.530 ;
        RECT 77.370 164.330 95.170 164.470 ;
        RECT 77.370 164.270 77.690 164.330 ;
        RECT 94.850 164.270 95.170 164.330 ;
        RECT 96.690 164.470 97.010 164.530 ;
        RECT 131.970 164.470 132.110 164.670 ;
        RECT 136.710 164.610 137.030 164.670 ;
        RECT 96.690 164.330 132.110 164.470 ;
        RECT 96.690 164.270 97.010 164.330 ;
        RECT 70.010 164.130 70.330 164.190 ;
        RECT 85.190 164.130 85.510 164.190 ;
        RECT 70.010 163.990 85.510 164.130 ;
        RECT 70.010 163.930 70.330 163.990 ;
        RECT 85.190 163.930 85.510 163.990 ;
        RECT 90.250 164.130 90.570 164.190 ;
        RECT 109.570 164.130 109.890 164.190 ;
        RECT 114.170 164.130 114.490 164.190 ;
        RECT 125.210 164.130 125.530 164.190 ;
        RECT 132.570 164.130 132.890 164.190 ;
        RECT 90.250 163.990 125.530 164.130 ;
        RECT 90.250 163.930 90.570 163.990 ;
        RECT 109.570 163.930 109.890 163.990 ;
        RECT 114.170 163.930 114.490 163.990 ;
        RECT 125.210 163.930 125.530 163.990 ;
        RECT 131.970 163.990 132.890 164.130 ;
        RECT 79.670 163.790 79.990 163.850 ;
        RECT 86.570 163.790 86.890 163.850 ;
        RECT 79.670 163.650 86.890 163.790 ;
        RECT 79.670 163.590 79.990 163.650 ;
        RECT 86.570 163.590 86.890 163.650 ;
        RECT 88.870 163.790 89.190 163.850 ;
        RECT 97.610 163.790 97.930 163.850 ;
        RECT 88.870 163.650 97.930 163.790 ;
        RECT 88.870 163.590 89.190 163.650 ;
        RECT 97.610 163.590 97.930 163.650 ;
        RECT 104.510 163.790 104.830 163.850 ;
        RECT 131.970 163.790 132.110 163.990 ;
        RECT 132.570 163.930 132.890 163.990 ;
        RECT 104.510 163.650 132.110 163.790 ;
        RECT 104.510 163.590 104.830 163.650 ;
        RECT 85.190 163.450 85.510 163.510 ;
        RECT 88.410 163.450 88.730 163.510 ;
        RECT 104.600 163.450 104.740 163.590 ;
        RECT 85.190 163.310 104.740 163.450 ;
        RECT 85.190 163.250 85.510 163.310 ;
        RECT 88.410 163.250 88.730 163.310 ;
        RECT 107.730 163.110 108.050 163.170 ;
        RECT 134.870 163.110 135.190 163.170 ;
        RECT 107.730 162.970 135.190 163.110 ;
        RECT 107.730 162.910 108.050 162.970 ;
        RECT 134.870 162.910 135.190 162.970 ;
        RECT 62.650 162.770 62.970 162.830 ;
        RECT 89.330 162.770 89.650 162.830 ;
        RECT 62.650 162.630 89.650 162.770 ;
        RECT 62.650 162.570 62.970 162.630 ;
        RECT 89.330 162.570 89.650 162.630 ;
        RECT 99.910 162.770 100.230 162.830 ;
        RECT 133.030 162.770 133.350 162.830 ;
        RECT 99.910 162.630 133.350 162.770 ;
        RECT 99.910 162.570 100.230 162.630 ;
        RECT 133.030 162.570 133.350 162.630 ;
        RECT 69.550 162.430 69.870 162.490 ;
        RECT 83.810 162.430 84.130 162.490 ;
        RECT 98.990 162.430 99.310 162.490 ;
        RECT 69.550 162.290 99.310 162.430 ;
        RECT 69.550 162.230 69.870 162.290 ;
        RECT 83.810 162.230 84.130 162.290 ;
        RECT 98.990 162.230 99.310 162.290 ;
        RECT 74.610 161.410 74.930 161.470 ;
        RECT 101.750 161.410 102.070 161.470 ;
        RECT 74.610 161.270 102.070 161.410 ;
        RECT 74.610 161.210 74.930 161.270 ;
        RECT 101.750 161.210 102.070 161.270 ;
        RECT 102.210 161.410 102.530 161.470 ;
        RECT 124.750 161.410 125.070 161.470 ;
        RECT 132.110 161.410 132.430 161.470 ;
        RECT 102.210 161.270 125.070 161.410 ;
        RECT 102.210 161.210 102.530 161.270 ;
        RECT 124.750 161.210 125.070 161.270 ;
        RECT 131.970 161.210 132.430 161.410 ;
        RECT 83.350 161.070 83.670 161.130 ;
        RECT 83.810 161.070 84.130 161.130 ;
        RECT 83.350 160.930 84.130 161.070 ;
        RECT 83.350 160.870 83.670 160.930 ;
        RECT 83.810 160.870 84.130 160.930 ;
        RECT 84.270 161.070 84.590 161.130 ;
        RECT 115.090 161.070 115.410 161.130 ;
        RECT 84.270 160.930 115.410 161.070 ;
        RECT 84.270 160.870 84.590 160.930 ;
        RECT 115.090 160.870 115.410 160.930 ;
        RECT 77.830 160.730 78.150 160.790 ;
        RECT 108.650 160.730 108.970 160.790 ;
        RECT 77.830 160.590 108.970 160.730 ;
        RECT 77.830 160.530 78.150 160.590 ;
        RECT 108.650 160.530 108.970 160.590 ;
        RECT 101.750 160.390 102.070 160.450 ;
        RECT 131.970 160.390 132.110 161.210 ;
        RECT 101.750 160.250 132.110 160.390 ;
        RECT 101.750 160.190 102.070 160.250 ;
        RECT 83.810 159.030 84.130 159.090 ;
        RECT 89.330 159.030 89.650 159.090 ;
        RECT 83.810 158.890 89.650 159.030 ;
        RECT 83.810 158.830 84.130 158.890 ;
        RECT 89.330 158.830 89.650 158.890 ;
        RECT 69.090 158.690 69.410 158.750 ;
        RECT 111.870 158.690 112.190 158.750 ;
        RECT 69.090 158.550 112.190 158.690 ;
        RECT 69.090 158.490 69.410 158.550 ;
        RECT 111.870 158.490 112.190 158.550 ;
        RECT 81.050 158.350 81.370 158.410 ;
        RECT 127.970 158.350 128.290 158.410 ;
        RECT 81.050 158.210 128.290 158.350 ;
        RECT 81.050 158.150 81.370 158.210 ;
        RECT 127.970 158.150 128.290 158.210 ;
        RECT 81.970 158.010 82.290 158.070 ;
        RECT 131.190 158.010 131.510 158.070 ;
        RECT 81.970 157.870 131.510 158.010 ;
        RECT 81.970 157.810 82.290 157.870 ;
        RECT 131.190 157.810 131.510 157.870 ;
        RECT 64.490 157.670 64.810 157.730 ;
        RECT 118.310 157.670 118.630 157.730 ;
        RECT 64.490 157.530 118.630 157.670 ;
        RECT 64.490 157.470 64.810 157.530 ;
        RECT 118.310 157.470 118.630 157.530 ;
        RECT 78.290 157.330 78.610 157.390 ;
        RECT 144.070 157.330 144.390 157.390 ;
        RECT 78.290 157.190 144.390 157.330 ;
        RECT 78.290 157.130 78.610 157.190 ;
        RECT 144.070 157.130 144.390 157.190 ;
        RECT 82.430 155.970 82.750 156.030 ;
        RECT 140.850 155.970 141.170 156.030 ;
        RECT 82.430 155.830 141.170 155.970 ;
        RECT 82.430 155.770 82.750 155.830 ;
        RECT 140.850 155.770 141.170 155.830 ;
        RECT 66.790 155.630 67.110 155.690 ;
        RECT 124.750 155.630 125.070 155.690 ;
        RECT 66.790 155.490 125.070 155.630 ;
        RECT 66.790 155.430 67.110 155.490 ;
        RECT 124.750 155.430 125.070 155.490 ;
        RECT 55.290 155.290 55.610 155.350 ;
        RECT 121.530 155.290 121.850 155.350 ;
        RECT 55.290 155.150 121.850 155.290 ;
        RECT 55.290 155.090 55.610 155.150 ;
        RECT 121.530 155.090 121.850 155.150 ;
      LAYER met2 ;
        RECT 66.810 221.070 67.090 221.570 ;
        RECT 86.130 221.070 86.410 221.570 ;
        RECT 89.350 221.080 89.630 221.570 ;
        RECT 89.880 221.250 90.480 221.390 ;
        RECT 89.880 221.080 90.020 221.250 ;
        RECT 89.350 221.070 90.020 221.080 ;
        RECT 27.250 209.265 27.530 209.635 ;
        RECT 64.980 209.460 65.240 209.780 ;
        RECT 27.320 207.740 27.460 209.265 ;
        RECT 46.010 208.925 47.550 209.295 ;
        RECT 35.540 207.760 35.800 208.080 ;
        RECT 56.700 207.760 56.960 208.080 ;
        RECT 27.260 207.420 27.520 207.740 ;
        RECT 25.420 206.740 25.680 207.060 ;
        RECT 25.480 206.235 25.620 206.740 ;
        RECT 25.410 205.865 25.690 206.235 ;
        RECT 35.600 206.040 35.740 207.760 ;
        RECT 53.020 206.740 53.280 207.060 ;
        RECT 42.710 206.205 44.250 206.575 ;
        RECT 35.540 205.720 35.800 206.040 ;
        RECT 52.100 205.720 52.360 206.040 ;
        RECT 51.180 205.040 51.440 205.360 ;
        RECT 52.160 205.270 52.300 205.720 ;
        RECT 52.560 205.270 52.820 205.360 ;
        RECT 52.160 205.130 52.820 205.270 ;
        RECT 30.020 204.700 30.280 205.020 ;
        RECT 36.460 204.700 36.720 205.020 ;
        RECT 37.840 204.700 38.100 205.020 ;
        RECT 38.300 204.700 38.560 205.020 ;
        RECT 39.680 204.700 39.940 205.020 ;
        RECT 25.420 204.020 25.680 204.340 ;
        RECT 25.480 202.835 25.620 204.020 ;
        RECT 30.080 203.320 30.220 204.700 ;
        RECT 30.020 203.000 30.280 203.320 ;
        RECT 25.410 202.465 25.690 202.835 ;
        RECT 32.780 202.320 33.040 202.640 ;
        RECT 31.400 193.820 31.660 194.140 ;
        RECT 25.420 193.140 25.680 193.460 ;
        RECT 25.480 192.635 25.620 193.140 ;
        RECT 25.410 192.265 25.690 192.635 ;
        RECT 31.460 192.440 31.600 193.820 ;
        RECT 31.400 192.120 31.660 192.440 ;
        RECT 25.420 191.440 25.680 191.760 ;
        RECT 32.320 191.440 32.580 191.760 ;
        RECT 25.480 189.235 25.620 191.440 ;
        RECT 30.020 191.275 30.280 191.420 ;
        RECT 30.010 190.905 30.290 191.275 ;
        RECT 32.380 189.720 32.520 191.440 ;
        RECT 32.320 189.400 32.580 189.720 ;
        RECT 25.410 188.865 25.690 189.235 ;
        RECT 31.400 188.380 31.660 188.700 ;
        RECT 24.500 185.835 24.760 185.980 ;
        RECT 24.490 185.465 24.770 185.835 ;
        RECT 31.460 183.600 31.600 188.380 ;
        RECT 31.860 185.660 32.120 185.980 ;
        RECT 31.400 183.280 31.660 183.600 ;
        RECT 31.920 183.260 32.060 185.660 ;
        RECT 32.840 184.280 32.980 202.320 ;
        RECT 36.520 199.580 36.660 204.700 ;
        RECT 37.900 203.320 38.040 204.700 ;
        RECT 37.840 203.000 38.100 203.320 ;
        RECT 38.360 202.640 38.500 204.700 ;
        RECT 38.300 202.320 38.560 202.640 ;
        RECT 38.360 200.600 38.500 202.320 ;
        RECT 38.300 200.280 38.560 200.600 ;
        RECT 36.460 199.260 36.720 199.580 ;
        RECT 37.380 196.880 37.640 197.200 ;
        RECT 37.440 189.720 37.580 196.880 ;
        RECT 38.360 194.140 38.500 200.280 ;
        RECT 39.220 199.260 39.480 199.580 ;
        RECT 38.300 193.820 38.560 194.140 ;
        RECT 37.840 191.100 38.100 191.420 ;
        RECT 37.380 189.400 37.640 189.720 ;
        RECT 36.460 188.380 36.720 188.700 ;
        RECT 37.380 188.380 37.640 188.700 ;
        RECT 36.520 185.640 36.660 188.380 ;
        RECT 37.440 185.980 37.580 188.380 ;
        RECT 37.900 187.000 38.040 191.100 ;
        RECT 38.760 188.380 39.020 188.700 ;
        RECT 38.820 187.000 38.960 188.380 ;
        RECT 37.840 186.680 38.100 187.000 ;
        RECT 38.760 186.680 39.020 187.000 ;
        RECT 38.820 185.980 38.960 186.680 ;
        RECT 37.380 185.660 37.640 185.980 ;
        RECT 38.760 185.660 39.020 185.980 ;
        RECT 36.460 185.320 36.720 185.640 ;
        RECT 32.780 183.960 33.040 184.280 ;
        RECT 39.280 183.260 39.420 199.260 ;
        RECT 39.740 194.480 39.880 204.700 ;
        RECT 47.960 204.360 48.220 204.680 ;
        RECT 50.260 204.360 50.520 204.680 ;
        RECT 50.720 204.360 50.980 204.680 ;
        RECT 41.520 204.020 41.780 204.340 ;
        RECT 42.900 204.020 43.160 204.340 ;
        RECT 41.580 203.320 41.720 204.020 ;
        RECT 41.520 203.000 41.780 203.320 ;
        RECT 41.060 201.980 41.320 202.300 ;
        RECT 41.120 196.860 41.260 201.980 ;
        RECT 41.060 196.540 41.320 196.860 ;
        RECT 41.060 195.860 41.320 196.180 ;
        RECT 41.120 195.160 41.260 195.860 ;
        RECT 41.060 194.840 41.320 195.160 ;
        RECT 39.680 194.160 39.940 194.480 ;
        RECT 40.140 191.440 40.400 191.760 ;
        RECT 41.060 191.440 41.320 191.760 ;
        RECT 40.200 188.700 40.340 191.440 ;
        RECT 41.120 189.720 41.260 191.440 ;
        RECT 41.060 189.400 41.320 189.720 ;
        RECT 40.140 188.380 40.400 188.700 ;
        RECT 41.580 188.020 41.720 203.000 ;
        RECT 42.960 202.980 43.100 204.020 ;
        RECT 46.010 203.485 47.550 203.855 ;
        RECT 42.900 202.660 43.160 202.980 ;
        RECT 44.740 202.660 45.000 202.980 ;
        RECT 47.500 202.660 47.760 202.980 ;
        RECT 44.800 201.620 44.940 202.660 ;
        RECT 45.660 202.320 45.920 202.640 ;
        RECT 44.740 201.300 45.000 201.620 ;
        RECT 42.710 200.765 44.250 201.135 ;
        RECT 43.360 198.920 43.620 199.240 ;
        RECT 43.420 196.520 43.560 198.920 ;
        RECT 44.800 197.880 44.940 201.300 ;
        RECT 44.740 197.560 45.000 197.880 ;
        RECT 45.200 197.220 45.460 197.540 ;
        RECT 44.740 196.540 45.000 196.860 ;
        RECT 41.980 196.200 42.240 196.520 ;
        RECT 43.360 196.200 43.620 196.520 ;
        RECT 42.040 195.070 42.180 196.200 ;
        RECT 42.710 195.325 44.250 195.695 ;
        RECT 44.800 195.160 44.940 196.540 ;
        RECT 42.040 194.930 42.640 195.070 ;
        RECT 42.500 194.140 42.640 194.930 ;
        RECT 44.740 194.840 45.000 195.160 ;
        RECT 45.260 194.820 45.400 197.220 ;
        RECT 45.200 194.500 45.460 194.820 ;
        RECT 42.440 193.820 42.700 194.140 ;
        RECT 44.280 193.480 44.540 193.800 ;
        RECT 44.340 191.080 44.480 193.480 ;
        RECT 45.720 192.100 45.860 202.320 ;
        RECT 47.560 201.960 47.700 202.660 ;
        RECT 47.500 201.640 47.760 201.960 ;
        RECT 48.020 199.580 48.160 204.360 ;
        RECT 49.340 204.020 49.600 204.340 ;
        RECT 49.400 203.320 49.540 204.020 ;
        RECT 49.340 203.230 49.600 203.320 ;
        RECT 49.340 203.090 50.000 203.230 ;
        RECT 49.340 203.000 49.600 203.090 ;
        RECT 48.420 202.320 48.680 202.640 ;
        RECT 48.480 200.600 48.620 202.320 ;
        RECT 48.420 200.280 48.680 200.600 ;
        RECT 47.500 199.260 47.760 199.580 ;
        RECT 47.960 199.260 48.220 199.580 ;
        RECT 47.560 198.900 47.700 199.260 ;
        RECT 48.480 198.900 48.620 200.280 ;
        RECT 48.880 199.940 49.140 200.260 ;
        RECT 47.500 198.810 47.760 198.900 ;
        RECT 47.500 198.670 48.160 198.810 ;
        RECT 47.500 198.580 47.760 198.670 ;
        RECT 46.010 198.045 47.550 198.415 ;
        RECT 46.120 197.560 46.380 197.880 ;
        RECT 46.180 194.140 46.320 197.560 ;
        RECT 48.020 196.715 48.160 198.670 ;
        RECT 48.420 198.580 48.680 198.900 ;
        RECT 48.480 197.200 48.620 198.580 ;
        RECT 48.420 196.880 48.680 197.200 ;
        RECT 47.950 196.345 48.230 196.715 ;
        RECT 48.940 194.140 49.080 199.940 ;
        RECT 49.860 199.580 50.000 203.090 ;
        RECT 50.320 202.980 50.460 204.360 ;
        RECT 50.260 202.660 50.520 202.980 ;
        RECT 49.800 199.260 50.060 199.580 ;
        RECT 50.320 199.240 50.460 202.660 ;
        RECT 50.780 202.640 50.920 204.360 ;
        RECT 51.240 203.320 51.380 205.040 ;
        RECT 51.640 204.020 51.900 204.340 ;
        RECT 51.180 203.000 51.440 203.320 ;
        RECT 51.700 202.640 51.840 204.020 ;
        RECT 50.720 202.320 50.980 202.640 ;
        RECT 51.640 202.320 51.900 202.640 ;
        RECT 52.160 202.300 52.300 205.130 ;
        RECT 52.560 205.040 52.820 205.130 ;
        RECT 53.080 205.020 53.220 206.740 ;
        RECT 53.940 205.720 54.200 206.040 ;
        RECT 53.020 204.700 53.280 205.020 ;
        RECT 54.000 203.320 54.140 205.720 ;
        RECT 54.400 205.040 54.660 205.360 ;
        RECT 53.940 203.000 54.200 203.320 ;
        RECT 52.100 201.980 52.360 202.300 ;
        RECT 53.020 199.940 53.280 200.260 ;
        RECT 50.260 198.920 50.520 199.240 ;
        RECT 50.320 197.540 50.460 198.920 ;
        RECT 50.260 197.220 50.520 197.540 ;
        RECT 53.080 197.200 53.220 199.940 ;
        RECT 53.020 196.880 53.280 197.200 ;
        RECT 50.260 196.200 50.520 196.520 ;
        RECT 49.800 195.860 50.060 196.180 ;
        RECT 49.340 194.160 49.600 194.480 ;
        RECT 46.120 193.820 46.380 194.140 ;
        RECT 47.960 193.820 48.220 194.140 ;
        RECT 48.880 193.820 49.140 194.140 ;
        RECT 46.010 192.605 47.550 192.975 ;
        RECT 45.660 191.780 45.920 192.100 ;
        RECT 44.280 190.760 44.540 191.080 ;
        RECT 42.710 189.885 44.250 190.255 ;
        RECT 43.360 189.400 43.620 189.720 ;
        RECT 47.500 189.400 47.760 189.720 ;
        RECT 42.900 188.040 43.160 188.360 ;
        RECT 41.520 187.700 41.780 188.020 ;
        RECT 41.520 186.340 41.780 186.660 ;
        RECT 40.600 185.720 40.860 185.980 ;
        RECT 41.580 185.720 41.720 186.340 ;
        RECT 42.960 185.720 43.100 188.040 ;
        RECT 40.600 185.660 41.260 185.720 ;
        RECT 40.140 185.320 40.400 185.640 ;
        RECT 40.660 185.580 41.260 185.660 ;
        RECT 31.860 182.940 32.120 183.260 ;
        RECT 39.220 182.940 39.480 183.260 ;
        RECT 40.200 182.920 40.340 185.320 ;
        RECT 41.120 185.300 41.260 185.580 ;
        RECT 41.580 185.580 43.100 185.720 ;
        RECT 43.420 185.640 43.560 189.400 ;
        RECT 45.660 188.720 45.920 189.040 ;
        RECT 44.740 186.680 45.000 187.000 ;
        RECT 44.800 185.640 44.940 186.680 ;
        RECT 41.060 184.980 41.320 185.300 ;
        RECT 25.420 182.600 25.680 182.920 ;
        RECT 40.140 182.600 40.400 182.920 ;
        RECT 25.480 182.435 25.620 182.600 ;
        RECT 25.410 182.065 25.690 182.435 ;
        RECT 25.420 179.540 25.680 179.860 ;
        RECT 25.480 179.035 25.620 179.540 ;
        RECT 25.410 178.665 25.690 179.035 ;
        RECT 41.120 177.480 41.260 184.980 ;
        RECT 41.580 178.160 41.720 185.580 ;
        RECT 42.960 185.300 43.100 185.580 ;
        RECT 43.360 185.320 43.620 185.640 ;
        RECT 44.740 185.320 45.000 185.640 ;
        RECT 41.980 184.980 42.240 185.300 ;
        RECT 42.900 184.980 43.160 185.300 ;
        RECT 42.040 183.940 42.180 184.980 ;
        RECT 42.710 184.445 44.250 184.815 ;
        RECT 41.980 183.620 42.240 183.940 ;
        RECT 44.800 183.600 44.940 185.320 ;
        RECT 45.200 184.980 45.460 185.300 ;
        RECT 44.740 183.280 45.000 183.600 ;
        RECT 45.260 183.260 45.400 184.980 ;
        RECT 45.200 182.940 45.460 183.260 ;
        RECT 43.360 182.260 43.620 182.580 ;
        RECT 44.280 182.260 44.540 182.580 ;
        RECT 43.420 180.540 43.560 182.260 ;
        RECT 44.340 180.880 44.480 182.260 ;
        RECT 45.720 181.470 45.860 188.720 ;
        RECT 47.560 188.020 47.700 189.400 ;
        RECT 47.500 187.700 47.760 188.020 ;
        RECT 46.010 187.165 47.550 187.535 ;
        RECT 47.030 183.425 47.310 183.795 ;
        RECT 47.040 183.280 47.300 183.425 ;
        RECT 46.010 181.725 47.550 182.095 ;
        RECT 48.020 181.560 48.160 193.820 ;
        RECT 48.410 192.265 48.690 192.635 ;
        RECT 48.480 192.100 48.620 192.265 ;
        RECT 48.420 191.780 48.680 192.100 ;
        RECT 49.400 191.760 49.540 194.160 ;
        RECT 49.860 191.955 50.000 195.860 ;
        RECT 49.340 191.440 49.600 191.760 ;
        RECT 49.790 191.585 50.070 191.955 ;
        RECT 48.420 191.100 48.680 191.420 ;
        RECT 48.480 187.875 48.620 191.100 ;
        RECT 48.880 189.060 49.140 189.380 ;
        RECT 48.410 187.505 48.690 187.875 ;
        RECT 48.940 186.320 49.080 189.060 ;
        RECT 49.400 188.700 49.540 191.440 ;
        RECT 49.340 188.380 49.600 188.700 ;
        RECT 48.880 186.000 49.140 186.320 ;
        RECT 48.880 184.980 49.140 185.300 ;
        RECT 49.340 184.980 49.600 185.300 ;
        RECT 48.940 182.920 49.080 184.980 ;
        RECT 49.400 183.260 49.540 184.980 ;
        RECT 49.340 182.940 49.600 183.260 ;
        RECT 48.880 182.600 49.140 182.920 ;
        RECT 45.720 181.330 46.320 181.470 ;
        RECT 44.280 180.560 44.540 180.880 ;
        RECT 44.740 180.560 45.000 180.880 ;
        RECT 45.660 180.560 45.920 180.880 ;
        RECT 43.360 180.220 43.620 180.540 ;
        RECT 42.710 179.005 44.250 179.375 ;
        RECT 44.800 178.840 44.940 180.560 ;
        RECT 45.200 180.220 45.460 180.540 ;
        RECT 44.740 178.520 45.000 178.840 ;
        RECT 41.520 177.840 41.780 178.160 ;
        RECT 41.060 177.160 41.320 177.480 ;
        RECT 41.580 175.780 41.720 177.840 ;
        RECT 45.260 177.820 45.400 180.220 ;
        RECT 45.200 177.500 45.460 177.820 ;
        RECT 42.900 177.160 43.160 177.480 ;
        RECT 41.520 175.460 41.780 175.780 ;
        RECT 42.960 175.440 43.100 177.160 ;
        RECT 45.720 176.120 45.860 180.560 ;
        RECT 46.180 178.500 46.320 181.330 ;
        RECT 47.960 181.240 48.220 181.560 ;
        RECT 48.420 181.240 48.680 181.560 ;
        RECT 47.500 179.770 47.760 179.860 ;
        RECT 48.480 179.770 48.620 181.240 ;
        RECT 48.940 181.220 49.080 182.600 ;
        RECT 48.880 180.900 49.140 181.220 ;
        RECT 49.340 180.790 49.600 180.880 ;
        RECT 49.860 180.790 50.000 191.585 ;
        RECT 50.320 183.680 50.460 196.200 ;
        RECT 51.180 195.860 51.440 196.180 ;
        RECT 51.240 192.100 51.380 195.860 ;
        RECT 52.100 193.140 52.360 193.460 ;
        RECT 51.180 191.780 51.440 192.100 ;
        RECT 52.160 191.760 52.300 193.140 ;
        RECT 54.000 192.440 54.140 203.000 ;
        RECT 54.460 200.600 54.600 205.040 ;
        RECT 55.320 201.980 55.580 202.300 ;
        RECT 54.400 200.280 54.660 200.600 ;
        RECT 54.860 199.600 55.120 199.920 ;
        RECT 54.400 198.920 54.660 199.240 ;
        RECT 54.460 195.160 54.600 198.920 ;
        RECT 54.920 195.160 55.060 199.600 ;
        RECT 54.400 194.840 54.660 195.160 ;
        RECT 54.860 194.840 55.120 195.160 ;
        RECT 54.400 193.820 54.660 194.140 ;
        RECT 53.940 192.120 54.200 192.440 ;
        RECT 53.020 191.780 53.280 192.100 ;
        RECT 52.100 191.440 52.360 191.760 ;
        RECT 52.560 191.440 52.820 191.760 ;
        RECT 51.180 190.420 51.440 190.740 ;
        RECT 51.240 188.360 51.380 190.420 ;
        RECT 52.160 189.380 52.300 191.440 ;
        RECT 52.100 189.060 52.360 189.380 ;
        RECT 52.100 188.380 52.360 188.700 ;
        RECT 51.180 188.040 51.440 188.360 ;
        RECT 51.180 186.000 51.440 186.320 ;
        RECT 51.240 184.280 51.380 186.000 ;
        RECT 51.640 184.980 51.900 185.300 ;
        RECT 51.180 183.960 51.440 184.280 ;
        RECT 50.320 183.540 51.380 183.680 ;
        RECT 51.700 183.600 51.840 184.980 ;
        RECT 50.320 183.260 50.460 183.540 ;
        RECT 50.260 182.940 50.520 183.260 ;
        RECT 50.720 182.940 50.980 183.260 ;
        RECT 50.780 181.560 50.920 182.940 ;
        RECT 50.720 181.240 50.980 181.560 ;
        RECT 49.340 180.650 50.000 180.790 ;
        RECT 50.250 180.705 50.530 181.075 ;
        RECT 51.240 180.880 51.380 183.540 ;
        RECT 51.640 183.280 51.900 183.600 ;
        RECT 49.340 180.560 49.600 180.650 ;
        RECT 50.260 180.560 50.520 180.705 ;
        RECT 51.180 180.560 51.440 180.880 ;
        RECT 49.400 179.860 49.540 180.560 ;
        RECT 47.500 179.630 48.620 179.770 ;
        RECT 47.500 179.540 47.760 179.630 ;
        RECT 49.340 179.540 49.600 179.860 ;
        RECT 46.120 178.180 46.380 178.500 ;
        RECT 49.800 177.500 50.060 177.820 ;
        RECT 46.010 176.285 47.550 176.655 ;
        RECT 49.860 176.315 50.000 177.500 ;
        RECT 45.660 175.800 45.920 176.120 ;
        RECT 49.790 175.945 50.070 176.315 ;
        RECT 49.860 175.780 50.000 175.945 ;
        RECT 44.740 175.460 45.000 175.780 ;
        RECT 49.800 175.460 50.060 175.780 ;
        RECT 42.900 175.120 43.160 175.440 ;
        RECT 42.960 174.760 43.100 175.120 ;
        RECT 42.900 174.440 43.160 174.760 ;
        RECT 42.710 173.565 44.250 173.935 ;
        RECT 44.800 170.195 44.940 175.460 ;
        RECT 48.420 175.120 48.680 175.440 ;
        RECT 48.480 174.275 48.620 175.120 ;
        RECT 49.860 175.100 50.000 175.460 ;
        RECT 50.320 175.440 50.460 180.560 ;
        RECT 51.180 179.540 51.440 179.860 ;
        RECT 51.240 178.160 51.380 179.540 ;
        RECT 51.700 178.840 51.840 183.280 ;
        RECT 52.160 181.560 52.300 188.380 ;
        RECT 52.620 184.280 52.760 191.440 ;
        RECT 53.080 188.700 53.220 191.780 ;
        RECT 54.460 190.740 54.600 193.820 ;
        RECT 54.860 193.140 55.120 193.460 ;
        RECT 54.920 191.760 55.060 193.140 ;
        RECT 54.860 191.440 55.120 191.760 ;
        RECT 54.400 190.420 54.660 190.740 ;
        RECT 53.940 189.400 54.200 189.720 ;
        RECT 53.020 188.380 53.280 188.700 ;
        RECT 53.480 188.380 53.740 188.700 ;
        RECT 54.000 188.555 54.140 189.400 ;
        RECT 54.460 188.700 54.600 190.420 ;
        RECT 54.920 189.720 55.060 191.440 ;
        RECT 55.380 189.915 55.520 201.980 ;
        RECT 56.760 199.580 56.900 207.760 ;
        RECT 57.160 207.420 57.420 207.740 ;
        RECT 57.620 207.420 57.880 207.740 ;
        RECT 57.220 199.920 57.360 207.420 ;
        RECT 57.680 206.040 57.820 207.420 ;
        RECT 57.620 205.720 57.880 206.040 ;
        RECT 64.060 205.380 64.320 205.700 ;
        RECT 63.600 204.360 63.860 204.680 ;
        RECT 58.080 204.020 58.340 204.340 ;
        RECT 58.140 202.300 58.280 204.020 ;
        RECT 59.460 203.000 59.720 203.320 ;
        RECT 58.080 201.980 58.340 202.300 ;
        RECT 58.540 201.980 58.800 202.300 ;
        RECT 58.600 199.920 58.740 201.980 ;
        RECT 57.160 199.600 57.420 199.920 ;
        RECT 58.540 199.600 58.800 199.920 ;
        RECT 56.700 199.260 56.960 199.580 ;
        RECT 56.760 197.540 56.900 199.260 ;
        RECT 57.160 198.580 57.420 198.900 ;
        RECT 56.700 197.220 56.960 197.540 ;
        RECT 57.220 194.560 57.360 198.580 ;
        RECT 56.300 194.420 57.360 194.560 ;
        RECT 56.300 192.520 56.440 194.420 ;
        RECT 57.620 194.160 57.880 194.480 ;
        RECT 57.160 193.820 57.420 194.140 ;
        RECT 56.700 193.480 56.960 193.800 ;
        RECT 55.840 192.380 56.440 192.520 ;
        RECT 54.860 189.400 55.120 189.720 ;
        RECT 55.310 189.545 55.590 189.915 ;
        RECT 53.080 185.640 53.220 188.380 ;
        RECT 53.020 185.320 53.280 185.640 ;
        RECT 52.560 183.960 52.820 184.280 ;
        RECT 53.540 183.940 53.680 188.380 ;
        RECT 53.930 188.185 54.210 188.555 ;
        RECT 54.400 188.380 54.660 188.700 ;
        RECT 54.000 186.320 54.140 188.185 ;
        RECT 55.840 186.320 55.980 192.380 ;
        RECT 56.760 191.760 56.900 193.480 ;
        RECT 56.240 191.440 56.500 191.760 ;
        RECT 56.700 191.440 56.960 191.760 ;
        RECT 56.300 189.720 56.440 191.440 ;
        RECT 57.220 189.720 57.360 193.820 ;
        RECT 57.680 192.440 57.820 194.160 ;
        RECT 58.080 193.820 58.340 194.140 ;
        RECT 57.620 192.120 57.880 192.440 ;
        RECT 56.240 189.400 56.500 189.720 ;
        RECT 57.160 189.400 57.420 189.720 ;
        RECT 57.680 189.120 57.820 192.120 ;
        RECT 58.140 191.080 58.280 193.820 ;
        RECT 58.540 192.120 58.800 192.440 ;
        RECT 58.600 191.760 58.740 192.120 ;
        RECT 58.540 191.440 58.800 191.760 ;
        RECT 58.080 190.990 58.340 191.080 ;
        RECT 58.080 190.850 58.740 190.990 ;
        RECT 58.080 190.760 58.340 190.850 ;
        RECT 56.760 188.980 57.820 189.120 ;
        RECT 56.760 188.700 56.900 188.980 ;
        RECT 56.700 188.380 56.960 188.700 ;
        RECT 57.610 188.185 57.890 188.555 ;
        RECT 57.620 188.040 57.880 188.185 ;
        RECT 53.940 186.000 54.200 186.320 ;
        RECT 54.400 186.000 54.660 186.320 ;
        RECT 55.780 186.000 56.040 186.320 ;
        RECT 54.460 185.640 54.600 186.000 ;
        RECT 55.320 185.660 55.580 185.980 ;
        RECT 54.400 185.320 54.660 185.640 ;
        RECT 55.380 183.940 55.520 185.660 ;
        RECT 57.620 183.960 57.880 184.280 ;
        RECT 53.480 183.620 53.740 183.940 ;
        RECT 55.320 183.620 55.580 183.940 ;
        RECT 55.380 183.260 55.520 183.620 ;
        RECT 54.400 183.170 54.660 183.260 ;
        RECT 55.320 183.170 55.580 183.260 ;
        RECT 54.400 183.030 55.580 183.170 ;
        RECT 54.400 182.940 54.660 183.030 ;
        RECT 55.320 182.940 55.580 183.030 ;
        RECT 55.780 182.940 56.040 183.260 ;
        RECT 56.700 182.940 56.960 183.260 ;
        RECT 53.020 182.260 53.280 182.580 ;
        RECT 52.100 181.240 52.360 181.560 ;
        RECT 53.080 181.220 53.220 182.260 ;
        RECT 53.020 180.900 53.280 181.220 ;
        RECT 54.460 179.860 54.600 182.940 ;
        RECT 54.860 182.490 55.120 182.580 ;
        RECT 55.840 182.490 55.980 182.940 ;
        RECT 54.860 182.350 55.980 182.490 ;
        RECT 54.860 182.260 55.120 182.350 ;
        RECT 56.760 181.560 56.900 182.940 ;
        RECT 57.680 181.560 57.820 183.960 ;
        RECT 58.080 182.940 58.340 183.260 ;
        RECT 56.700 181.240 56.960 181.560 ;
        RECT 57.620 181.240 57.880 181.560 ;
        RECT 58.140 180.880 58.280 182.940 ;
        RECT 55.320 180.560 55.580 180.880 ;
        RECT 56.240 180.560 56.500 180.880 ;
        RECT 58.080 180.560 58.340 180.880 ;
        RECT 54.400 179.540 54.660 179.860 ;
        RECT 51.640 178.520 51.900 178.840 ;
        RECT 51.180 177.840 51.440 178.160 ;
        RECT 55.380 176.120 55.520 180.560 ;
        RECT 56.300 179.860 56.440 180.560 ;
        RECT 56.240 179.540 56.500 179.860 ;
        RECT 57.150 178.665 57.430 179.035 ;
        RECT 57.220 178.500 57.360 178.665 ;
        RECT 57.160 178.180 57.420 178.500 ;
        RECT 58.140 177.820 58.280 180.560 ;
        RECT 58.080 177.500 58.340 177.820 ;
        RECT 55.320 175.800 55.580 176.120 ;
        RECT 50.720 175.460 50.980 175.780 ;
        RECT 50.260 175.120 50.520 175.440 ;
        RECT 49.800 174.780 50.060 175.100 ;
        RECT 48.410 173.905 48.690 174.275 ;
        RECT 46.010 170.845 47.550 171.215 ;
        RECT 44.730 169.825 45.010 170.195 ;
        RECT 25.420 168.835 25.680 168.980 ;
        RECT 25.410 168.465 25.690 168.835 ;
        RECT 42.710 168.125 44.250 168.495 ;
        RECT 44.800 167.960 44.940 169.825 ;
        RECT 49.340 169.680 49.600 170.000 ;
        RECT 49.400 167.960 49.540 169.680 ;
        RECT 50.780 169.515 50.920 175.460 ;
        RECT 55.380 170.680 55.520 175.800 ;
        RECT 58.080 175.120 58.340 175.440 ;
        RECT 58.140 172.720 58.280 175.120 ;
        RECT 58.080 172.400 58.340 172.720 ;
        RECT 55.320 170.360 55.580 170.680 ;
        RECT 58.600 170.000 58.740 190.850 ;
        RECT 59.520 186.515 59.660 203.000 ;
        RECT 60.380 202.320 60.640 202.640 ;
        RECT 60.440 200.600 60.580 202.320 ;
        RECT 61.760 201.980 62.020 202.300 ;
        RECT 62.680 201.980 62.940 202.300 ;
        RECT 60.380 200.280 60.640 200.600 ;
        RECT 60.840 197.220 61.100 197.540 ;
        RECT 60.370 196.345 60.650 196.715 ;
        RECT 59.920 193.480 60.180 193.800 ;
        RECT 59.980 191.760 60.120 193.480 ;
        RECT 59.920 191.440 60.180 191.760 ;
        RECT 59.980 191.275 60.120 191.440 ;
        RECT 59.910 190.905 60.190 191.275 ;
        RECT 59.980 189.720 60.120 190.905 ;
        RECT 59.920 189.400 60.180 189.720 ;
        RECT 59.450 186.145 59.730 186.515 ;
        RECT 59.520 180.540 59.660 186.145 ;
        RECT 59.980 180.880 60.120 189.400 ;
        RECT 60.440 183.600 60.580 196.345 ;
        RECT 60.380 183.280 60.640 183.600 ;
        RECT 60.440 180.880 60.580 183.280 ;
        RECT 59.920 180.560 60.180 180.880 ;
        RECT 60.380 180.560 60.640 180.880 ;
        RECT 59.460 180.220 59.720 180.540 ;
        RECT 59.980 180.395 60.120 180.560 ;
        RECT 59.520 176.120 59.660 180.220 ;
        RECT 59.910 180.025 60.190 180.395 ;
        RECT 59.980 178.160 60.120 180.025 ;
        RECT 60.900 179.715 61.040 197.220 ;
        RECT 61.820 186.660 61.960 201.980 ;
        RECT 62.740 199.580 62.880 201.980 ;
        RECT 62.680 199.260 62.940 199.580 ;
        RECT 62.740 197.540 62.880 199.260 ;
        RECT 63.140 198.580 63.400 198.900 ;
        RECT 62.680 197.280 62.940 197.540 ;
        RECT 62.280 197.220 62.940 197.280 ;
        RECT 62.280 197.140 62.880 197.220 ;
        RECT 62.280 194.480 62.420 197.140 ;
        RECT 63.200 196.860 63.340 198.580 ;
        RECT 63.660 197.280 63.800 204.360 ;
        RECT 64.120 200.260 64.260 205.380 ;
        RECT 65.040 205.020 65.180 209.460 ;
        RECT 66.880 208.080 67.020 221.070 ;
        RECT 82.920 210.140 83.180 210.460 ;
        RECT 75.100 208.440 75.360 208.760 ;
        RECT 66.820 207.760 67.080 208.080 ;
        RECT 68.200 206.740 68.460 207.060 ;
        RECT 72.340 206.740 72.600 207.060 ;
        RECT 64.980 204.700 65.240 205.020 ;
        RECT 65.440 204.700 65.700 205.020 ;
        RECT 66.820 204.700 67.080 205.020 ;
        RECT 64.510 201.785 64.790 202.155 ;
        RECT 64.060 199.940 64.320 200.260 ;
        RECT 64.050 197.280 64.330 197.395 ;
        RECT 63.660 197.140 64.330 197.280 ;
        RECT 64.050 197.025 64.330 197.140 ;
        RECT 63.140 196.540 63.400 196.860 ;
        RECT 63.140 194.840 63.400 195.160 ;
        RECT 62.680 194.675 62.940 194.820 ;
        RECT 62.220 194.160 62.480 194.480 ;
        RECT 62.670 194.305 62.950 194.675 ;
        RECT 62.680 193.820 62.940 194.140 ;
        RECT 62.740 191.080 62.880 193.820 ;
        RECT 62.680 190.760 62.940 191.080 ;
        RECT 62.670 189.545 62.950 189.915 ;
        RECT 62.740 189.040 62.880 189.545 ;
        RECT 62.680 188.720 62.940 189.040 ;
        RECT 62.220 188.040 62.480 188.360 ;
        RECT 61.760 186.340 62.020 186.660 ;
        RECT 62.280 184.280 62.420 188.040 ;
        RECT 62.220 183.960 62.480 184.280 ;
        RECT 62.280 181.220 62.420 183.960 ;
        RECT 63.200 183.940 63.340 194.840 ;
        RECT 64.120 193.800 64.260 197.025 ;
        RECT 64.060 193.480 64.320 193.800 ;
        RECT 64.120 191.420 64.260 193.480 ;
        RECT 64.060 191.100 64.320 191.420 ;
        RECT 63.600 190.420 63.860 190.740 ;
        RECT 63.140 183.795 63.400 183.940 ;
        RECT 63.130 183.425 63.410 183.795 ;
        RECT 63.660 181.640 63.800 190.420 ;
        RECT 64.050 187.505 64.330 187.875 ;
        RECT 63.200 181.500 63.800 181.640 ;
        RECT 61.760 180.900 62.020 181.220 ;
        RECT 62.220 180.900 62.480 181.220 ;
        RECT 60.830 179.345 61.110 179.715 ;
        RECT 59.920 177.840 60.180 178.160 ;
        RECT 60.900 177.820 61.040 179.345 ;
        RECT 61.300 178.180 61.560 178.500 ;
        RECT 61.820 178.240 61.960 180.900 ;
        RECT 63.200 178.355 63.340 181.500 ;
        RECT 63.600 180.900 63.860 181.220 ;
        RECT 63.660 179.860 63.800 180.900 ;
        RECT 64.120 180.540 64.260 187.505 ;
        RECT 64.580 180.880 64.720 201.785 ;
        RECT 65.040 197.960 65.180 204.700 ;
        RECT 65.500 203.320 65.640 204.700 ;
        RECT 65.900 204.360 66.160 204.680 ;
        RECT 65.440 203.000 65.700 203.320 ;
        RECT 65.440 202.320 65.700 202.640 ;
        RECT 65.500 198.900 65.640 202.320 ;
        RECT 65.960 199.920 66.100 204.360 ;
        RECT 66.360 201.980 66.620 202.300 ;
        RECT 65.900 199.600 66.160 199.920 ;
        RECT 66.420 199.580 66.560 201.980 ;
        RECT 66.360 199.260 66.620 199.580 ;
        RECT 65.440 198.580 65.700 198.900 ;
        RECT 65.040 197.820 65.640 197.960 ;
        RECT 66.880 197.880 67.020 204.700 ;
        RECT 67.280 204.020 67.540 204.340 ;
        RECT 67.340 202.980 67.480 204.020 ;
        RECT 67.280 202.660 67.540 202.980 ;
        RECT 67.280 201.980 67.540 202.300 ;
        RECT 67.740 201.980 68.000 202.300 ;
        RECT 67.340 200.600 67.480 201.980 ;
        RECT 67.280 200.280 67.540 200.600 ;
        RECT 67.280 199.260 67.540 199.580 ;
        RECT 65.500 197.200 65.640 197.820 ;
        RECT 66.820 197.560 67.080 197.880 ;
        RECT 64.980 196.880 65.240 197.200 ;
        RECT 65.440 197.110 65.700 197.200 ;
        RECT 65.440 196.970 66.100 197.110 ;
        RECT 65.440 196.880 65.700 196.970 ;
        RECT 65.040 192.440 65.180 196.880 ;
        RECT 65.440 195.860 65.700 196.180 ;
        RECT 65.500 195.160 65.640 195.860 ;
        RECT 65.440 194.840 65.700 195.160 ;
        RECT 64.980 192.120 65.240 192.440 ;
        RECT 65.960 189.380 66.100 196.970 ;
        RECT 66.360 195.860 66.620 196.180 ;
        RECT 66.820 195.860 67.080 196.180 ;
        RECT 66.420 193.800 66.560 195.860 ;
        RECT 66.880 194.820 67.020 195.860 ;
        RECT 66.820 194.500 67.080 194.820 ;
        RECT 66.360 193.480 66.620 193.800 ;
        RECT 67.340 192.100 67.480 199.260 ;
        RECT 67.800 197.880 67.940 201.980 ;
        RECT 68.260 197.880 68.400 206.740 ;
        RECT 70.950 205.185 71.230 205.555 ;
        RECT 69.110 204.505 69.390 204.875 ;
        RECT 69.180 202.980 69.320 204.505 ;
        RECT 69.580 204.020 69.840 204.340 ;
        RECT 69.120 202.660 69.380 202.980 ;
        RECT 69.640 202.640 69.780 204.020 ;
        RECT 69.580 202.320 69.840 202.640 ;
        RECT 71.020 200.600 71.160 205.185 ;
        RECT 71.420 204.360 71.680 204.680 ;
        RECT 71.480 201.620 71.620 204.360 ;
        RECT 71.880 201.980 72.140 202.300 ;
        RECT 71.420 201.300 71.680 201.620 ;
        RECT 70.960 200.280 71.220 200.600 ;
        RECT 70.490 199.745 70.770 200.115 ;
        RECT 68.660 199.435 68.920 199.580 ;
        RECT 68.650 199.065 68.930 199.435 ;
        RECT 67.740 197.560 68.000 197.880 ;
        RECT 68.200 197.560 68.460 197.880 ;
        RECT 69.580 197.790 69.840 197.880 ;
        RECT 69.180 197.650 69.840 197.790 ;
        RECT 67.740 196.540 68.000 196.860 ;
        RECT 67.800 192.440 67.940 196.540 ;
        RECT 68.260 194.820 68.400 197.560 ;
        RECT 69.180 197.280 69.320 197.650 ;
        RECT 69.580 197.560 69.840 197.650 ;
        RECT 69.570 197.280 69.850 197.395 ;
        RECT 69.180 197.140 69.850 197.280 ;
        RECT 69.570 197.025 69.850 197.140 ;
        RECT 69.580 196.880 69.840 197.025 ;
        RECT 70.040 196.880 70.300 197.200 ;
        RECT 69.120 196.200 69.380 196.520 ;
        RECT 69.180 194.820 69.320 196.200 ;
        RECT 70.100 195.160 70.240 196.880 ;
        RECT 70.040 194.840 70.300 195.160 ;
        RECT 70.560 194.820 70.700 199.745 ;
        RECT 71.480 198.900 71.620 201.300 ;
        RECT 71.420 198.580 71.680 198.900 ;
        RECT 71.420 196.880 71.680 197.200 ;
        RECT 71.480 196.715 71.620 196.880 ;
        RECT 71.410 196.345 71.690 196.715 ;
        RECT 70.960 195.860 71.220 196.180 ;
        RECT 71.020 195.160 71.160 195.860 ;
        RECT 71.410 195.665 71.690 196.035 ;
        RECT 70.960 194.840 71.220 195.160 ;
        RECT 68.200 194.500 68.460 194.820 ;
        RECT 69.120 194.500 69.380 194.820 ;
        RECT 70.500 194.500 70.760 194.820 ;
        RECT 68.260 192.440 68.400 194.500 ;
        RECT 68.660 193.995 68.920 194.140 ;
        RECT 68.650 193.625 68.930 193.995 ;
        RECT 67.740 192.120 68.000 192.440 ;
        RECT 68.200 192.120 68.460 192.440 ;
        RECT 67.280 191.780 67.540 192.100 ;
        RECT 67.800 191.955 67.940 192.120 ;
        RECT 67.340 190.595 67.480 191.780 ;
        RECT 67.730 191.585 68.010 191.955 ;
        RECT 70.960 191.780 71.220 192.100 ;
        RECT 68.200 191.100 68.460 191.420 ;
        RECT 69.570 191.160 69.850 191.275 ;
        RECT 70.040 191.160 70.300 191.420 ;
        RECT 69.570 191.100 70.300 191.160 ;
        RECT 67.270 190.225 67.550 190.595 ;
        RECT 68.260 189.380 68.400 191.100 ;
        RECT 69.120 190.760 69.380 191.080 ;
        RECT 69.570 191.020 70.240 191.100 ;
        RECT 69.570 190.905 69.850 191.020 ;
        RECT 69.180 189.720 69.320 190.760 ;
        RECT 70.500 190.420 70.760 190.740 ;
        RECT 69.120 189.400 69.380 189.720 ;
        RECT 65.900 189.060 66.160 189.380 ;
        RECT 68.200 189.290 68.460 189.380 ;
        RECT 68.200 189.150 68.860 189.290 ;
        RECT 68.200 189.060 68.460 189.150 ;
        RECT 65.960 186.400 66.100 189.060 ;
        RECT 66.360 188.380 66.620 188.700 ;
        RECT 66.420 187.000 66.560 188.380 ;
        RECT 66.360 186.680 66.620 187.000 ;
        RECT 67.280 186.400 67.540 186.660 ;
        RECT 65.960 186.340 67.540 186.400 ;
        RECT 65.960 186.320 67.480 186.340 ;
        RECT 65.440 186.000 65.700 186.320 ;
        RECT 65.900 186.260 67.480 186.320 ;
        RECT 65.900 186.000 66.160 186.260 ;
        RECT 64.520 180.560 64.780 180.880 ;
        RECT 64.060 180.220 64.320 180.540 ;
        RECT 63.600 179.540 63.860 179.860 ;
        RECT 64.580 179.035 64.720 180.560 ;
        RECT 64.510 178.665 64.790 179.035 ;
        RECT 60.840 177.500 61.100 177.820 ;
        RECT 61.360 176.120 61.500 178.180 ;
        RECT 61.820 178.100 62.420 178.240 ;
        RECT 61.760 177.500 62.020 177.820 ;
        RECT 59.460 176.030 59.720 176.120 ;
        RECT 59.460 175.890 60.120 176.030 ;
        RECT 59.460 175.800 59.720 175.890 ;
        RECT 59.460 175.350 59.720 175.440 ;
        RECT 59.060 175.210 59.720 175.350 ;
        RECT 59.060 171.700 59.200 175.210 ;
        RECT 59.460 175.120 59.720 175.210 ;
        RECT 59.460 172.400 59.720 172.720 ;
        RECT 59.000 171.380 59.260 171.700 ;
        RECT 57.160 169.680 57.420 170.000 ;
        RECT 58.540 169.680 58.800 170.000 ;
        RECT 50.710 169.145 50.990 169.515 ;
        RECT 50.780 167.960 50.920 169.145 ;
        RECT 57.220 168.980 57.360 169.680 ;
        RECT 58.080 169.340 58.340 169.660 ;
        RECT 57.160 168.660 57.420 168.980 ;
        RECT 44.740 167.640 45.000 167.960 ;
        RECT 49.340 167.640 49.600 167.960 ;
        RECT 50.720 167.640 50.980 167.960 ;
        RECT 54.390 167.105 54.670 167.475 ;
        RECT 56.240 167.190 56.500 167.280 ;
        RECT 57.220 167.190 57.360 168.660 ;
        RECT 54.460 166.940 54.600 167.105 ;
        RECT 56.240 167.050 57.360 167.190 ;
        RECT 56.240 166.960 56.500 167.050 ;
        RECT 58.140 166.940 58.280 169.340 ;
        RECT 58.600 167.960 58.740 169.680 ;
        RECT 59.060 167.960 59.200 171.380 ;
        RECT 59.520 169.320 59.660 172.400 ;
        RECT 59.980 172.380 60.120 175.890 ;
        RECT 61.300 175.800 61.560 176.120 ;
        RECT 60.380 175.120 60.640 175.440 ;
        RECT 61.300 175.120 61.560 175.440 ;
        RECT 60.440 173.060 60.580 175.120 ;
        RECT 61.360 174.955 61.500 175.120 ;
        RECT 61.290 174.585 61.570 174.955 ;
        RECT 61.820 174.760 61.960 177.500 ;
        RECT 61.760 174.440 62.020 174.760 ;
        RECT 60.380 172.740 60.640 173.060 ;
        RECT 62.280 172.630 62.420 178.100 ;
        RECT 63.130 177.985 63.410 178.355 ;
        RECT 64.520 177.500 64.780 177.820 ;
        RECT 62.680 177.050 62.940 177.140 ;
        RECT 62.680 176.910 63.800 177.050 ;
        RECT 62.680 176.820 62.940 176.910 ;
        RECT 63.130 175.265 63.410 175.635 ;
        RECT 63.200 173.400 63.340 175.265 ;
        RECT 63.660 173.400 63.800 176.910 ;
        RECT 64.580 175.780 64.720 177.500 ;
        RECT 64.970 177.305 65.250 177.675 ;
        RECT 64.520 175.460 64.780 175.780 ;
        RECT 64.510 174.585 64.790 174.955 ;
        RECT 63.140 173.080 63.400 173.400 ;
        RECT 63.600 173.080 63.860 173.400 ;
        RECT 64.580 173.060 64.720 174.585 ;
        RECT 62.280 172.490 62.880 172.630 ;
        RECT 63.130 172.545 63.410 172.915 ;
        RECT 64.520 172.740 64.780 173.060 ;
        RECT 59.920 172.120 60.180 172.380 ;
        RECT 62.210 172.120 62.490 172.235 ;
        RECT 59.920 172.060 62.490 172.120 ;
        RECT 59.980 171.980 62.490 172.060 ;
        RECT 62.210 171.865 62.490 171.980 ;
        RECT 62.220 171.720 62.480 171.865 ;
        RECT 62.740 170.000 62.880 172.490 ;
        RECT 63.200 172.380 63.340 172.545 ;
        RECT 63.140 172.060 63.400 172.380 ;
        RECT 64.580 172.040 64.720 172.740 ;
        RECT 64.520 171.720 64.780 172.040 ;
        RECT 64.580 170.680 64.720 171.720 ;
        RECT 64.520 170.360 64.780 170.680 ;
        RECT 65.040 170.250 65.180 177.305 ;
        RECT 65.500 177.050 65.640 186.000 ;
        RECT 68.200 185.320 68.460 185.640 ;
        RECT 67.280 183.620 67.540 183.940 ;
        RECT 66.810 180.025 67.090 180.395 ;
        RECT 65.900 179.715 66.160 179.860 ;
        RECT 65.890 179.345 66.170 179.715 ;
        RECT 65.900 178.520 66.160 178.840 ;
        RECT 65.960 178.160 66.100 178.520 ;
        RECT 66.880 178.500 67.020 180.025 ;
        RECT 66.820 178.180 67.080 178.500 ;
        RECT 65.900 177.840 66.160 178.160 ;
        RECT 66.360 177.500 66.620 177.820 ;
        RECT 65.900 177.050 66.160 177.140 ;
        RECT 65.500 176.910 66.160 177.050 ;
        RECT 65.900 176.820 66.160 176.910 ;
        RECT 66.420 175.635 66.560 177.500 ;
        RECT 65.900 175.120 66.160 175.440 ;
        RECT 66.350 175.265 66.630 175.635 ;
        RECT 65.440 174.440 65.700 174.760 ;
        RECT 65.500 173.400 65.640 174.440 ;
        RECT 65.440 173.080 65.700 173.400 ;
        RECT 65.440 170.250 65.700 170.340 ;
        RECT 65.040 170.110 65.700 170.250 ;
        RECT 62.680 169.680 62.940 170.000 ;
        RECT 59.460 169.000 59.720 169.320 ;
        RECT 65.040 168.980 65.180 170.110 ;
        RECT 65.440 170.020 65.700 170.110 ;
        RECT 65.440 169.340 65.700 169.660 ;
        RECT 64.980 168.660 65.240 168.980 ;
        RECT 58.540 167.640 58.800 167.960 ;
        RECT 59.000 167.640 59.260 167.960 ;
        RECT 59.920 167.870 60.180 167.960 ;
        RECT 59.520 167.730 60.180 167.870 ;
        RECT 58.600 167.360 58.740 167.640 ;
        RECT 59.520 167.360 59.660 167.730 ;
        RECT 59.920 167.640 60.180 167.730 ;
        RECT 58.600 167.220 59.660 167.360 ;
        RECT 41.060 166.620 41.320 166.940 ;
        RECT 44.280 166.620 44.540 166.940 ;
        RECT 47.960 166.620 48.220 166.940 ;
        RECT 50.720 166.620 50.980 166.940 ;
        RECT 54.400 166.620 54.660 166.940 ;
        RECT 58.080 166.620 58.340 166.940 ;
        RECT 64.520 166.620 64.780 166.940 ;
        RECT 41.120 155.210 41.260 166.620 ;
        RECT 44.340 155.210 44.480 166.620 ;
        RECT 46.010 165.405 47.550 165.775 ;
        RECT 48.020 161.070 48.160 166.620 ;
        RECT 47.560 160.930 48.160 161.070 ;
        RECT 47.560 155.210 47.700 160.930 ;
        RECT 50.780 155.210 50.920 166.620 ;
        RECT 57.160 166.280 57.420 166.600 ;
        RECT 55.320 165.940 55.580 166.260 ;
        RECT 55.380 155.380 55.520 165.940 ;
        RECT 41.050 154.710 41.330 155.210 ;
        RECT 44.270 154.710 44.550 155.210 ;
        RECT 47.490 154.710 47.770 155.210 ;
        RECT 50.710 154.710 50.990 155.210 ;
        RECT 55.320 155.060 55.580 155.380 ;
        RECT 57.220 155.210 57.360 166.280 ;
        RECT 60.380 165.940 60.640 166.260 ;
        RECT 62.680 165.940 62.940 166.260 ;
        RECT 60.440 155.210 60.580 165.940 ;
        RECT 62.740 162.860 62.880 165.940 ;
        RECT 62.680 162.540 62.940 162.860 ;
        RECT 64.580 157.760 64.720 166.620 ;
        RECT 65.040 166.600 65.180 168.660 ;
        RECT 65.500 167.960 65.640 169.340 ;
        RECT 65.440 167.640 65.700 167.960 ;
        RECT 65.960 166.795 66.100 175.120 ;
        RECT 66.820 174.100 67.080 174.420 ;
        RECT 66.360 172.740 66.620 173.060 ;
        RECT 66.420 172.380 66.560 172.740 ;
        RECT 66.360 172.235 66.620 172.380 ;
        RECT 66.350 171.865 66.630 172.235 ;
        RECT 66.360 169.680 66.620 170.000 ;
        RECT 66.420 167.280 66.560 169.680 ;
        RECT 66.360 166.960 66.620 167.280 ;
        RECT 64.980 166.280 65.240 166.600 ;
        RECT 65.890 166.425 66.170 166.795 ;
        RECT 65.440 165.940 65.700 166.260 ;
        RECT 65.500 165.435 65.640 165.940 ;
        RECT 65.430 165.065 65.710 165.435 ;
        RECT 64.520 157.440 64.780 157.760 ;
        RECT 66.880 155.720 67.020 174.100 ;
        RECT 67.340 170.000 67.480 183.620 ;
        RECT 68.260 182.580 68.400 185.320 ;
        RECT 68.720 183.260 68.860 189.150 ;
        RECT 70.560 189.040 70.700 190.420 ;
        RECT 70.500 188.720 70.760 189.040 ;
        RECT 70.500 187.700 70.760 188.020 ;
        RECT 69.580 186.680 69.840 187.000 ;
        RECT 68.660 182.940 68.920 183.260 ;
        RECT 68.200 182.260 68.460 182.580 ;
        RECT 67.740 180.560 68.000 180.880 ;
        RECT 67.800 175.780 67.940 180.560 ;
        RECT 68.200 179.540 68.460 179.860 ;
        RECT 67.740 175.460 68.000 175.780 ;
        RECT 67.800 173.400 67.940 175.460 ;
        RECT 68.260 175.350 68.400 179.540 ;
        RECT 68.720 178.500 68.860 182.940 ;
        RECT 69.640 178.840 69.780 186.680 ;
        RECT 70.560 184.280 70.700 187.700 ;
        RECT 70.500 183.960 70.760 184.280 ;
        RECT 71.020 183.600 71.160 191.780 ;
        RECT 71.480 188.700 71.620 195.665 ;
        RECT 71.940 189.040 72.080 201.980 ;
        RECT 72.400 201.620 72.540 206.740 ;
        RECT 75.160 204.680 75.300 208.440 ;
        RECT 75.560 207.760 75.820 208.080 ;
        RECT 75.100 204.360 75.360 204.680 ;
        RECT 72.790 203.825 73.070 204.195 ;
        RECT 74.640 204.020 74.900 204.340 ;
        RECT 72.340 201.300 72.600 201.620 ;
        RECT 72.340 193.820 72.600 194.140 ;
        RECT 72.400 190.595 72.540 193.820 ;
        RECT 72.330 190.225 72.610 190.595 ;
        RECT 71.880 188.720 72.140 189.040 ;
        RECT 71.420 188.380 71.680 188.700 ;
        RECT 72.340 187.700 72.600 188.020 ;
        RECT 72.400 183.600 72.540 187.700 ;
        RECT 70.960 183.280 71.220 183.600 ;
        RECT 71.880 183.280 72.140 183.600 ;
        RECT 72.340 183.280 72.600 183.600 ;
        RECT 71.410 182.065 71.690 182.435 ;
        RECT 70.040 181.470 70.300 181.560 ;
        RECT 70.040 181.330 70.700 181.470 ;
        RECT 70.040 181.240 70.300 181.330 ;
        RECT 69.580 178.520 69.840 178.840 ;
        RECT 68.660 178.180 68.920 178.500 ;
        RECT 68.660 177.500 68.920 177.820 ;
        RECT 70.040 177.500 70.300 177.820 ;
        RECT 68.720 176.120 68.860 177.500 ;
        RECT 70.100 176.120 70.240 177.500 ;
        RECT 68.660 175.800 68.920 176.120 ;
        RECT 70.040 175.800 70.300 176.120 ;
        RECT 68.660 175.350 68.920 175.440 ;
        RECT 68.260 175.210 68.920 175.350 ;
        RECT 69.110 175.265 69.390 175.635 ;
        RECT 68.660 175.120 68.920 175.210 ;
        RECT 67.740 173.080 68.000 173.400 ;
        RECT 68.720 172.380 68.860 175.120 ;
        RECT 67.740 172.290 68.000 172.380 ;
        RECT 68.660 172.290 68.920 172.380 ;
        RECT 67.740 172.235 68.920 172.290 ;
        RECT 67.740 172.150 68.930 172.235 ;
        RECT 67.740 172.060 68.000 172.150 ;
        RECT 68.650 171.865 68.930 172.150 ;
        RECT 69.180 170.000 69.320 175.265 ;
        RECT 70.560 175.100 70.700 181.330 ;
        RECT 70.960 177.500 71.220 177.820 ;
        RECT 71.020 176.120 71.160 177.500 ;
        RECT 70.960 175.800 71.220 176.120 ;
        RECT 70.960 175.120 71.220 175.440 ;
        RECT 70.040 174.780 70.300 175.100 ;
        RECT 70.500 174.780 70.760 175.100 ;
        RECT 69.580 174.440 69.840 174.760 ;
        RECT 69.640 170.340 69.780 174.440 ;
        RECT 70.100 172.720 70.240 174.780 ;
        RECT 71.020 174.420 71.160 175.120 ;
        RECT 71.480 174.420 71.620 182.065 ;
        RECT 70.960 174.100 71.220 174.420 ;
        RECT 71.420 174.100 71.680 174.420 ;
        RECT 70.040 172.400 70.300 172.720 ;
        RECT 69.580 170.020 69.840 170.340 ;
        RECT 67.280 169.680 67.540 170.000 ;
        RECT 68.660 169.680 68.920 170.000 ;
        RECT 69.120 169.680 69.380 170.000 ;
        RECT 68.720 168.835 68.860 169.680 ;
        RECT 69.180 169.320 69.320 169.680 ;
        RECT 69.580 169.340 69.840 169.660 ;
        RECT 69.120 169.000 69.380 169.320 ;
        RECT 68.650 168.465 68.930 168.835 ;
        RECT 67.740 166.620 68.000 166.940 ;
        RECT 69.120 166.620 69.380 166.940 ;
        RECT 67.800 164.075 67.940 166.620 ;
        RECT 67.730 163.705 68.010 164.075 ;
        RECT 69.180 158.780 69.320 166.620 ;
        RECT 69.640 162.520 69.780 169.340 ;
        RECT 70.100 169.320 70.240 172.400 ;
        RECT 70.500 171.380 70.760 171.700 ;
        RECT 70.040 169.000 70.300 169.320 ;
        RECT 70.560 167.530 70.700 171.380 ;
        RECT 71.020 168.040 71.160 174.100 ;
        RECT 71.940 173.400 72.080 183.280 ;
        RECT 72.330 181.385 72.610 181.755 ;
        RECT 72.400 176.315 72.540 181.385 ;
        RECT 72.860 181.220 73.000 203.825 ;
        RECT 74.700 202.640 74.840 204.020 ;
        RECT 75.620 202.835 75.760 207.760 ;
        RECT 77.400 207.420 77.660 207.740 ;
        RECT 77.460 206.040 77.600 207.420 ;
        RECT 79.700 207.080 79.960 207.400 ;
        RECT 77.400 205.720 77.660 206.040 ;
        RECT 77.860 204.700 78.120 205.020 ;
        RECT 75.550 202.720 75.830 202.835 ;
        RECT 74.640 202.320 74.900 202.640 ;
        RECT 75.160 202.580 75.830 202.720 ;
        RECT 73.720 201.300 73.980 201.620 ;
        RECT 73.780 199.920 73.920 201.300 ;
        RECT 73.720 199.600 73.980 199.920 ;
        RECT 74.180 199.600 74.440 199.920 ;
        RECT 73.720 196.540 73.980 196.860 ;
        RECT 73.260 194.675 73.520 194.820 ;
        RECT 73.250 194.305 73.530 194.675 ;
        RECT 73.260 193.820 73.520 194.140 ;
        RECT 73.320 181.560 73.460 193.820 ;
        RECT 73.780 190.740 73.920 196.540 ;
        RECT 74.240 194.480 74.380 199.600 ;
        RECT 74.180 194.160 74.440 194.480 ;
        RECT 74.170 193.625 74.450 193.995 ;
        RECT 73.720 190.420 73.980 190.740 ;
        RECT 74.240 189.915 74.380 193.625 ;
        RECT 75.160 192.100 75.300 202.580 ;
        RECT 75.550 202.465 75.830 202.580 ;
        RECT 76.020 202.320 76.280 202.640 ;
        RECT 76.940 202.320 77.200 202.640 ;
        RECT 77.400 202.320 77.660 202.640 ;
        RECT 75.560 201.980 75.820 202.300 ;
        RECT 75.620 196.035 75.760 201.980 ;
        RECT 75.550 195.665 75.830 196.035 ;
        RECT 75.100 191.780 75.360 192.100 ;
        RECT 73.720 189.400 73.980 189.720 ;
        RECT 74.170 189.545 74.450 189.915 ;
        RECT 73.780 186.320 73.920 189.400 ;
        RECT 74.240 188.700 74.380 189.545 ;
        RECT 76.080 189.120 76.220 202.320 ;
        RECT 77.000 194.480 77.140 202.320 ;
        RECT 77.460 201.620 77.600 202.320 ;
        RECT 77.400 201.300 77.660 201.620 ;
        RECT 77.460 199.580 77.600 201.300 ;
        RECT 77.920 200.600 78.060 204.700 ;
        RECT 78.320 202.320 78.580 202.640 ;
        RECT 77.860 200.280 78.120 200.600 ;
        RECT 78.380 200.260 78.520 202.320 ;
        RECT 78.320 199.940 78.580 200.260 ;
        RECT 77.400 199.260 77.660 199.580 ;
        RECT 76.940 194.160 77.200 194.480 ;
        RECT 75.160 188.980 76.220 189.120 ;
        RECT 74.180 188.380 74.440 188.700 ;
        RECT 74.640 188.380 74.900 188.700 ;
        RECT 73.720 186.000 73.980 186.320 ;
        RECT 73.720 185.320 73.980 185.640 ;
        RECT 73.780 183.600 73.920 185.320 ;
        RECT 74.240 183.600 74.380 188.380 ;
        RECT 74.700 185.300 74.840 188.380 ;
        RECT 75.160 187.000 75.300 188.980 ;
        RECT 76.020 188.040 76.280 188.360 ;
        RECT 75.100 186.680 75.360 187.000 ;
        RECT 75.560 186.680 75.820 187.000 ;
        RECT 75.620 186.320 75.760 186.680 ;
        RECT 76.080 186.320 76.220 188.040 ;
        RECT 78.380 188.020 78.520 199.940 ;
        RECT 79.240 198.920 79.500 199.240 ;
        RECT 79.300 197.540 79.440 198.920 ;
        RECT 79.240 197.220 79.500 197.540 ;
        RECT 78.780 193.140 79.040 193.460 ;
        RECT 76.540 187.620 78.060 187.760 ;
        RECT 78.320 187.700 78.580 188.020 ;
        RECT 76.540 186.660 76.680 187.620 ;
        RECT 77.400 186.680 77.660 187.000 ;
        RECT 76.480 186.340 76.740 186.660 ;
        RECT 75.100 186.000 75.360 186.320 ;
        RECT 75.560 186.000 75.820 186.320 ;
        RECT 76.020 186.000 76.280 186.320 ;
        RECT 76.940 186.000 77.200 186.320 ;
        RECT 74.640 184.980 74.900 185.300 ;
        RECT 73.720 183.280 73.980 183.600 ;
        RECT 74.180 183.280 74.440 183.600 ;
        RECT 74.700 183.260 74.840 184.980 ;
        RECT 74.640 182.940 74.900 183.260 ;
        RECT 73.260 181.240 73.520 181.560 ;
        RECT 72.800 180.900 73.060 181.220 ;
        RECT 75.160 180.280 75.300 186.000 ;
        RECT 76.080 183.940 76.220 186.000 ;
        RECT 76.480 185.660 76.740 185.980 ;
        RECT 77.000 185.835 77.140 186.000 ;
        RECT 76.540 185.300 76.680 185.660 ;
        RECT 76.930 185.465 77.210 185.835 ;
        RECT 76.480 184.980 76.740 185.300 ;
        RECT 77.460 183.940 77.600 186.680 ;
        RECT 77.920 186.320 78.060 187.620 ;
        RECT 77.860 186.000 78.120 186.320 ;
        RECT 77.920 183.940 78.060 186.000 ;
        RECT 76.020 183.620 76.280 183.940 ;
        RECT 77.400 183.620 77.660 183.940 ;
        RECT 77.860 183.620 78.120 183.940 ;
        RECT 76.940 183.280 77.200 183.600 ;
        RECT 77.000 181.470 77.140 183.280 ;
        RECT 77.860 182.940 78.120 183.260 ;
        RECT 77.920 182.580 78.060 182.940 ;
        RECT 78.380 182.580 78.520 187.700 ;
        RECT 77.860 182.260 78.120 182.580 ;
        RECT 78.320 182.260 78.580 182.580 ;
        RECT 77.000 181.330 77.600 181.470 ;
        RECT 76.020 180.560 76.280 180.880 ;
        RECT 76.940 180.560 77.200 180.880 ;
        RECT 74.240 180.140 75.300 180.280 ;
        RECT 73.720 176.820 73.980 177.140 ;
        RECT 72.330 175.945 72.610 176.315 ;
        RECT 73.260 175.460 73.520 175.780 ;
        RECT 72.340 175.120 72.600 175.440 ;
        RECT 71.880 173.080 72.140 173.400 ;
        RECT 71.410 172.545 71.690 172.915 ;
        RECT 71.480 172.380 71.620 172.545 ;
        RECT 71.420 172.060 71.680 172.380 ;
        RECT 71.880 172.060 72.140 172.380 ;
        RECT 71.940 170.680 72.080 172.060 ;
        RECT 71.880 170.360 72.140 170.680 ;
        RECT 71.870 169.825 72.150 170.195 ;
        RECT 71.940 168.980 72.080 169.825 ;
        RECT 71.880 168.660 72.140 168.980 ;
        RECT 71.020 167.900 71.620 168.040 ;
        RECT 70.560 167.390 71.160 167.530 ;
        RECT 71.020 166.940 71.160 167.390 ;
        RECT 70.500 166.620 70.760 166.940 ;
        RECT 70.960 166.620 71.220 166.940 ;
        RECT 70.040 165.940 70.300 166.260 ;
        RECT 70.560 166.115 70.700 166.620 ;
        RECT 70.100 164.220 70.240 165.940 ;
        RECT 70.490 165.745 70.770 166.115 ;
        RECT 70.040 163.900 70.300 164.220 ;
        RECT 69.580 162.200 69.840 162.520 ;
        RECT 69.120 158.460 69.380 158.780 ;
        RECT 71.480 156.595 71.620 167.900 ;
        RECT 72.400 158.635 72.540 175.120 ;
        RECT 73.320 173.400 73.460 175.460 ;
        RECT 73.260 173.080 73.520 173.400 ;
        RECT 73.320 172.915 73.460 173.080 ;
        RECT 73.250 172.545 73.530 172.915 ;
        RECT 72.800 171.380 73.060 171.700 ;
        RECT 72.860 170.680 73.000 171.380 ;
        RECT 72.800 170.360 73.060 170.680 ;
        RECT 72.790 167.785 73.070 168.155 ;
        RECT 72.860 167.620 73.000 167.785 ;
        RECT 72.800 167.300 73.060 167.620 ;
        RECT 73.260 166.620 73.520 166.940 ;
        RECT 73.320 164.900 73.460 166.620 ;
        RECT 73.260 164.580 73.520 164.900 ;
        RECT 72.330 158.265 72.610 158.635 ;
        RECT 71.410 156.225 71.690 156.595 ;
        RECT 73.780 155.915 73.920 176.820 ;
        RECT 74.240 172.720 74.380 180.140 ;
        RECT 74.630 179.345 74.910 179.715 ;
        RECT 74.700 178.500 74.840 179.345 ;
        RECT 74.640 178.180 74.900 178.500 ;
        RECT 74.640 177.160 74.900 177.480 ;
        RECT 74.180 172.400 74.440 172.720 ;
        RECT 74.180 169.340 74.440 169.660 ;
        RECT 74.240 164.755 74.380 169.340 ;
        RECT 74.170 164.385 74.450 164.755 ;
        RECT 74.700 161.500 74.840 177.160 ;
        RECT 75.100 176.820 75.360 177.140 ;
        RECT 75.560 176.820 75.820 177.140 ;
        RECT 75.160 175.780 75.300 176.820 ;
        RECT 75.100 175.460 75.360 175.780 ;
        RECT 75.620 175.635 75.760 176.820 ;
        RECT 76.080 176.315 76.220 180.560 ;
        RECT 76.480 180.220 76.740 180.540 ;
        RECT 76.010 175.945 76.290 176.315 ;
        RECT 76.540 176.120 76.680 180.220 ;
        RECT 77.000 179.860 77.140 180.560 ;
        RECT 77.460 180.200 77.600 181.330 ;
        RECT 77.920 180.395 78.060 182.260 ;
        RECT 78.320 180.560 78.580 180.880 ;
        RECT 77.400 179.880 77.660 180.200 ;
        RECT 77.850 180.025 78.130 180.395 ;
        RECT 76.940 179.540 77.200 179.860 ;
        RECT 77.000 179.035 77.140 179.540 ;
        RECT 76.930 178.665 77.210 179.035 ;
        RECT 77.460 178.500 77.600 179.880 ;
        RECT 77.400 178.180 77.660 178.500 ;
        RECT 77.860 178.180 78.120 178.500 ;
        RECT 77.920 176.120 78.060 178.180 ;
        RECT 78.380 177.820 78.520 180.560 ;
        RECT 78.840 180.200 78.980 193.140 ;
        RECT 79.760 188.020 79.900 207.080 ;
        RECT 80.160 206.740 80.420 207.060 ;
        RECT 80.220 206.040 80.360 206.740 ;
        RECT 80.160 205.720 80.420 206.040 ;
        RECT 81.540 205.040 81.800 205.360 ;
        RECT 80.620 204.360 80.880 204.680 ;
        RECT 80.680 202.640 80.820 204.360 ;
        RECT 80.620 202.320 80.880 202.640 ;
        RECT 80.150 200.425 80.430 200.795 ;
        RECT 80.220 199.580 80.360 200.425 ;
        RECT 80.160 199.260 80.420 199.580 ;
        RECT 80.160 195.860 80.420 196.180 ;
        RECT 80.220 194.140 80.360 195.860 ;
        RECT 80.680 195.160 80.820 202.320 ;
        RECT 81.080 201.300 81.340 201.620 ;
        RECT 81.140 199.920 81.280 201.300 ;
        RECT 81.600 199.920 81.740 205.040 ;
        RECT 82.460 203.000 82.720 203.320 ;
        RECT 82.520 201.960 82.660 203.000 ;
        RECT 82.460 201.640 82.720 201.960 ;
        RECT 81.080 199.600 81.340 199.920 ;
        RECT 81.540 199.600 81.800 199.920 ;
        RECT 81.080 198.920 81.340 199.240 ;
        RECT 81.140 197.880 81.280 198.920 ;
        RECT 81.600 197.880 81.740 199.600 ;
        RECT 81.080 197.560 81.340 197.880 ;
        RECT 81.540 197.560 81.800 197.880 ;
        RECT 80.620 194.840 80.880 195.160 ;
        RECT 81.080 194.160 81.340 194.480 ;
        RECT 80.160 193.820 80.420 194.140 ;
        RECT 81.140 192.440 81.280 194.160 ;
        RECT 82.000 193.480 82.260 193.800 ;
        RECT 81.080 192.120 81.340 192.440 ;
        RECT 81.140 191.955 81.280 192.120 ;
        RECT 81.070 191.585 81.350 191.955 ;
        RECT 80.160 190.420 80.420 190.740 ;
        RECT 80.220 188.700 80.360 190.420 ;
        RECT 81.080 188.720 81.340 189.040 ;
        RECT 80.160 188.380 80.420 188.700 ;
        RECT 80.610 188.185 80.890 188.555 ;
        RECT 79.700 187.700 79.960 188.020 ;
        RECT 80.150 186.825 80.430 187.195 ;
        RECT 79.240 186.000 79.500 186.320 ;
        RECT 79.700 186.000 79.960 186.320 ;
        RECT 79.300 184.280 79.440 186.000 ;
        RECT 79.760 185.835 79.900 186.000 ;
        RECT 80.220 185.980 80.360 186.825 ;
        RECT 79.690 185.465 79.970 185.835 ;
        RECT 80.160 185.660 80.420 185.980 ;
        RECT 79.240 183.960 79.500 184.280 ;
        RECT 79.760 183.600 79.900 185.465 ;
        RECT 79.700 183.280 79.960 183.600 ;
        RECT 80.680 182.580 80.820 188.185 ;
        RECT 81.140 183.260 81.280 188.720 ;
        RECT 81.530 187.505 81.810 187.875 ;
        RECT 81.080 182.940 81.340 183.260 ;
        RECT 79.240 182.490 79.500 182.580 ;
        RECT 79.240 182.350 80.360 182.490 ;
        RECT 79.240 182.260 79.500 182.350 ;
        RECT 79.700 181.240 79.960 181.560 ;
        RECT 79.240 180.900 79.500 181.220 ;
        RECT 78.780 179.880 79.040 180.200 ;
        RECT 78.320 177.500 78.580 177.820 ;
        RECT 78.840 177.140 78.980 179.880 ;
        RECT 79.300 177.820 79.440 180.900 ;
        RECT 79.240 177.500 79.500 177.820 ;
        RECT 78.780 176.820 79.040 177.140 ;
        RECT 79.240 176.820 79.500 177.140 ;
        RECT 76.480 175.800 76.740 176.120 ;
        RECT 77.860 175.800 78.120 176.120 ;
        RECT 75.160 172.040 75.300 175.460 ;
        RECT 75.550 175.265 75.830 175.635 ;
        RECT 75.560 174.780 75.820 175.100 ;
        RECT 75.100 171.720 75.360 172.040 ;
        RECT 75.100 170.590 75.360 170.680 ;
        RECT 75.620 170.590 75.760 174.780 ;
        RECT 76.540 174.420 76.680 175.800 ;
        RECT 76.940 175.120 77.200 175.440 ;
        RECT 77.000 174.955 77.140 175.120 ;
        RECT 76.930 174.585 77.210 174.955 ;
        RECT 77.400 174.440 77.660 174.760 ;
        RECT 76.480 174.100 76.740 174.420 ;
        RECT 76.540 173.400 76.680 174.100 ;
        RECT 77.460 173.595 77.600 174.440 ;
        RECT 76.480 173.310 76.740 173.400 ;
        RECT 76.480 173.170 77.140 173.310 ;
        RECT 77.390 173.225 77.670 173.595 ;
        RECT 76.480 173.080 76.740 173.170 ;
        RECT 76.470 172.545 76.750 172.915 ;
        RECT 76.540 172.380 76.680 172.545 ;
        RECT 76.480 172.290 76.740 172.380 ;
        RECT 75.100 170.450 75.760 170.590 ;
        RECT 76.080 172.150 76.740 172.290 ;
        RECT 75.100 170.360 75.360 170.450 ;
        RECT 76.080 170.080 76.220 172.150 ;
        RECT 76.480 172.060 76.740 172.150 ;
        RECT 77.000 171.440 77.140 173.170 ;
        RECT 77.400 172.290 77.660 172.380 ;
        RECT 77.920 172.290 78.060 175.800 ;
        RECT 78.780 175.120 79.040 175.440 ;
        RECT 78.320 173.080 78.580 173.400 ;
        RECT 77.400 172.150 78.060 172.290 ;
        RECT 77.400 172.060 77.660 172.150 ;
        RECT 75.160 169.940 76.220 170.080 ;
        RECT 76.540 171.300 77.140 171.440 ;
        RECT 75.160 168.980 75.300 169.940 ;
        RECT 75.100 168.660 75.360 168.980 ;
        RECT 75.560 168.660 75.820 168.980 ;
        RECT 75.100 167.190 75.360 167.280 ;
        RECT 75.620 167.190 75.760 168.660 ;
        RECT 76.540 168.040 76.680 171.300 ;
        RECT 76.940 170.250 77.200 170.340 ;
        RECT 77.460 170.250 77.600 172.060 ;
        RECT 78.380 170.680 78.520 173.080 ;
        RECT 78.320 170.360 78.580 170.680 ;
        RECT 76.940 170.110 77.600 170.250 ;
        RECT 76.940 170.020 77.200 170.110 ;
        RECT 77.000 168.980 77.140 170.020 ;
        RECT 76.940 168.660 77.200 168.980 ;
        RECT 77.400 168.660 77.660 168.980 ;
        RECT 77.460 168.040 77.600 168.660 ;
        RECT 78.840 168.580 78.980 175.120 ;
        RECT 79.300 173.400 79.440 176.820 ;
        RECT 79.240 173.080 79.500 173.400 ;
        RECT 79.240 172.060 79.500 172.380 ;
        RECT 79.300 170.000 79.440 172.060 ;
        RECT 79.240 169.680 79.500 170.000 ;
        RECT 79.240 169.000 79.500 169.320 ;
        RECT 76.540 167.900 77.600 168.040 ;
        RECT 78.380 168.440 78.980 168.580 ;
        RECT 77.860 167.640 78.120 167.960 ;
        RECT 75.100 167.050 75.760 167.190 ;
        RECT 75.100 166.960 75.360 167.050 ;
        RECT 76.020 166.620 76.280 166.940 ;
        RECT 77.400 166.620 77.660 166.940 ;
        RECT 76.080 165.240 76.220 166.620 ;
        RECT 76.020 164.920 76.280 165.240 ;
        RECT 77.460 164.560 77.600 166.620 ;
        RECT 77.400 164.240 77.660 164.560 ;
        RECT 74.640 161.180 74.900 161.500 ;
        RECT 77.920 160.820 78.060 167.640 ;
        RECT 77.860 160.500 78.120 160.820 ;
        RECT 78.380 157.420 78.520 168.440 ;
        RECT 79.300 168.040 79.440 169.000 ;
        RECT 78.840 167.900 79.440 168.040 ;
        RECT 78.840 165.435 78.980 167.900 ;
        RECT 79.240 165.940 79.500 166.260 ;
        RECT 78.770 165.065 79.050 165.435 ;
        RECT 79.300 160.675 79.440 165.940 ;
        RECT 79.760 163.880 79.900 181.240 ;
        RECT 80.220 180.880 80.360 182.350 ;
        RECT 80.620 182.260 80.880 182.580 ;
        RECT 80.680 181.075 80.820 182.260 ;
        RECT 80.160 180.560 80.420 180.880 ;
        RECT 80.610 180.705 80.890 181.075 ;
        RECT 81.140 177.820 81.280 182.940 ;
        RECT 81.600 181.560 81.740 187.505 ;
        RECT 82.060 185.720 82.200 193.480 ;
        RECT 82.060 185.580 82.660 185.720 ;
        RECT 82.520 185.300 82.660 185.580 ;
        RECT 82.460 184.980 82.720 185.300 ;
        RECT 82.450 184.105 82.730 184.475 ;
        RECT 82.520 183.940 82.660 184.105 ;
        RECT 82.460 183.850 82.720 183.940 ;
        RECT 82.060 183.710 82.720 183.850 ;
        RECT 81.540 181.240 81.800 181.560 ;
        RECT 82.060 181.220 82.200 183.710 ;
        RECT 82.460 183.620 82.720 183.710 ;
        RECT 82.980 181.220 83.120 210.140 ;
        RECT 86.200 208.420 86.340 221.070 ;
        RECT 89.420 220.940 90.020 221.070 ;
        RECT 87.050 219.465 87.330 219.835 ;
        RECT 87.120 208.760 87.260 219.465 ;
        RECT 88.890 212.665 89.170 213.035 ;
        RECT 87.060 208.440 87.320 208.760 ;
        RECT 86.140 208.100 86.400 208.420 ;
        RECT 88.440 207.760 88.700 208.080 ;
        RECT 84.300 206.740 84.560 207.060 ;
        RECT 83.840 205.040 84.100 205.360 ;
        RECT 83.380 204.020 83.640 204.340 ;
        RECT 83.440 202.640 83.580 204.020 ;
        RECT 83.900 203.320 84.040 205.040 ;
        RECT 84.360 203.320 84.500 206.740 ;
        RECT 88.500 205.700 88.640 207.760 ;
        RECT 88.960 206.040 89.100 212.665 ;
        RECT 89.820 209.800 90.080 210.120 ;
        RECT 89.360 208.440 89.620 208.760 ;
        RECT 89.420 208.275 89.560 208.440 ;
        RECT 89.350 207.905 89.630 208.275 ;
        RECT 88.900 205.720 89.160 206.040 ;
        RECT 87.520 205.380 87.780 205.700 ;
        RECT 88.440 205.380 88.700 205.700 ;
        RECT 85.220 204.700 85.480 205.020 ;
        RECT 85.680 204.700 85.940 205.020 ;
        RECT 84.760 204.020 85.020 204.340 ;
        RECT 83.840 203.000 84.100 203.320 ;
        RECT 84.300 203.000 84.560 203.320 ;
        RECT 83.380 202.320 83.640 202.640 ;
        RECT 83.440 200.260 83.580 202.320 ;
        RECT 83.380 199.940 83.640 200.260 ;
        RECT 83.380 199.260 83.640 199.580 ;
        RECT 83.440 198.900 83.580 199.260 ;
        RECT 83.380 198.580 83.640 198.900 ;
        RECT 83.440 197.200 83.580 198.580 ;
        RECT 83.380 196.880 83.640 197.200 ;
        RECT 83.380 195.860 83.640 196.180 ;
        RECT 83.440 194.140 83.580 195.860 ;
        RECT 83.900 194.140 84.040 203.000 ;
        RECT 84.300 201.300 84.560 201.620 ;
        RECT 84.360 197.200 84.500 201.300 ;
        RECT 84.820 197.200 84.960 204.020 ;
        RECT 84.300 196.880 84.560 197.200 ;
        RECT 84.760 196.880 85.020 197.200 ;
        RECT 85.280 196.600 85.420 204.700 ;
        RECT 85.740 199.580 85.880 204.700 ;
        RECT 86.600 204.020 86.860 204.340 ;
        RECT 86.140 201.300 86.400 201.620 ;
        RECT 86.200 200.260 86.340 201.300 ;
        RECT 86.140 199.940 86.400 200.260 ;
        RECT 85.680 199.435 85.940 199.580 ;
        RECT 85.670 199.065 85.950 199.435 ;
        RECT 85.740 196.860 85.880 199.065 ;
        RECT 84.360 196.460 85.420 196.600 ;
        RECT 85.680 196.540 85.940 196.860 ;
        RECT 86.660 196.715 86.800 204.020 ;
        RECT 87.580 199.580 87.720 205.380 ;
        RECT 88.960 205.020 89.100 205.720 ;
        RECT 87.980 204.700 88.240 205.020 ;
        RECT 88.900 204.700 89.160 205.020 ;
        RECT 88.040 203.515 88.180 204.700 ;
        RECT 88.440 204.360 88.700 204.680 ;
        RECT 87.970 203.145 88.250 203.515 ;
        RECT 87.980 201.980 88.240 202.300 ;
        RECT 88.040 199.920 88.180 201.980 ;
        RECT 87.980 199.600 88.240 199.920 ;
        RECT 87.520 199.260 87.780 199.580 ;
        RECT 87.060 198.580 87.320 198.900 ;
        RECT 83.380 193.820 83.640 194.140 ;
        RECT 83.840 193.820 84.100 194.140 ;
        RECT 83.370 190.905 83.650 191.275 ;
        RECT 83.900 191.080 84.040 193.820 ;
        RECT 83.380 190.760 83.640 190.905 ;
        RECT 83.840 190.760 84.100 191.080 ;
        RECT 84.360 188.555 84.500 196.460 ;
        RECT 86.590 196.345 86.870 196.715 ;
        RECT 85.210 195.665 85.490 196.035 ;
        RECT 85.280 195.160 85.420 195.665 ;
        RECT 85.220 194.840 85.480 195.160 ;
        RECT 84.750 194.305 85.030 194.675 ;
        RECT 84.760 194.160 85.020 194.305 ;
        RECT 85.280 194.140 85.420 194.840 ;
        RECT 85.220 193.820 85.480 194.140 ;
        RECT 85.280 191.760 85.420 193.820 ;
        RECT 86.140 193.140 86.400 193.460 ;
        RECT 86.600 193.140 86.860 193.460 ;
        RECT 86.200 192.440 86.340 193.140 ;
        RECT 86.140 192.120 86.400 192.440 ;
        RECT 86.660 191.760 86.800 193.140 ;
        RECT 87.120 191.760 87.260 198.580 ;
        RECT 85.220 191.440 85.480 191.760 ;
        RECT 86.140 191.440 86.400 191.760 ;
        RECT 86.600 191.440 86.860 191.760 ;
        RECT 87.060 191.440 87.320 191.760 ;
        RECT 84.290 188.185 84.570 188.555 ;
        RECT 84.760 188.040 85.020 188.360 ;
        RECT 83.380 187.700 83.640 188.020 ;
        RECT 83.440 186.320 83.580 187.700 ;
        RECT 84.290 186.825 84.570 187.195 ;
        RECT 84.360 186.660 84.500 186.825 ;
        RECT 84.300 186.340 84.560 186.660 ;
        RECT 84.820 186.320 84.960 188.040 ;
        RECT 83.380 186.000 83.640 186.320 ;
        RECT 83.840 186.000 84.100 186.320 ;
        RECT 84.760 186.000 85.020 186.320 ;
        RECT 83.380 184.980 83.640 185.300 ;
        RECT 83.440 184.280 83.580 184.980 ;
        RECT 83.380 183.960 83.640 184.280 ;
        RECT 83.370 183.425 83.650 183.795 ;
        RECT 82.000 180.900 82.260 181.220 ;
        RECT 82.920 180.900 83.180 181.220 ;
        RECT 83.440 180.395 83.580 183.425 ;
        RECT 82.460 179.880 82.720 180.200 ;
        RECT 83.370 180.025 83.650 180.395 ;
        RECT 81.540 178.180 81.800 178.500 ;
        RECT 81.080 177.500 81.340 177.820 ;
        RECT 80.160 176.820 80.420 177.140 ;
        RECT 80.220 166.940 80.360 176.820 ;
        RECT 80.620 174.100 80.880 174.420 ;
        RECT 80.680 172.380 80.820 174.100 ;
        RECT 81.070 173.905 81.350 174.275 ;
        RECT 80.620 172.060 80.880 172.380 ;
        RECT 80.620 171.380 80.880 171.700 ;
        RECT 80.680 169.320 80.820 171.380 ;
        RECT 81.140 170.000 81.280 173.905 ;
        RECT 81.080 169.680 81.340 170.000 ;
        RECT 80.620 169.000 80.880 169.320 ;
        RECT 80.680 168.155 80.820 169.000 ;
        RECT 80.610 167.785 80.890 168.155 ;
        RECT 81.600 166.940 81.740 178.180 ;
        RECT 82.000 177.500 82.260 177.820 ;
        RECT 82.060 176.995 82.200 177.500 ;
        RECT 81.990 176.625 82.270 176.995 ;
        RECT 82.000 174.440 82.260 174.760 ;
        RECT 82.060 172.380 82.200 174.440 ;
        RECT 82.000 172.060 82.260 172.380 ;
        RECT 82.000 170.020 82.260 170.340 ;
        RECT 80.160 166.620 80.420 166.940 ;
        RECT 81.540 166.620 81.800 166.940 ;
        RECT 81.080 165.940 81.340 166.260 ;
        RECT 79.700 163.560 79.960 163.880 ;
        RECT 79.230 160.305 79.510 160.675 ;
        RECT 81.140 158.440 81.280 165.940 ;
        RECT 81.080 158.120 81.340 158.440 ;
        RECT 82.060 158.100 82.200 170.020 ;
        RECT 82.000 157.780 82.260 158.100 ;
        RECT 78.320 157.100 78.580 157.420 ;
        RECT 82.520 156.060 82.660 179.880 ;
        RECT 82.910 177.985 83.190 178.355 ;
        RECT 83.440 178.160 83.580 180.025 ;
        RECT 83.900 178.840 84.040 186.000 ;
        RECT 84.300 185.660 84.560 185.980 ;
        RECT 84.360 184.280 84.500 185.660 ;
        RECT 85.280 185.155 85.420 191.440 ;
        RECT 86.200 189.720 86.340 191.440 ;
        RECT 86.660 191.080 86.800 191.440 ;
        RECT 86.600 190.760 86.860 191.080 ;
        RECT 87.060 190.760 87.320 191.080 ;
        RECT 86.140 189.400 86.400 189.720 ;
        RECT 87.120 189.040 87.260 190.760 ;
        RECT 87.060 188.720 87.320 189.040 ;
        RECT 87.580 188.440 87.720 199.260 ;
        RECT 88.500 198.900 88.640 204.360 ;
        RECT 89.360 203.000 89.620 203.320 ;
        RECT 88.900 201.980 89.160 202.300 ;
        RECT 88.960 200.600 89.100 201.980 ;
        RECT 88.900 200.280 89.160 200.600 ;
        RECT 88.900 199.435 89.160 199.580 ;
        RECT 88.890 199.065 89.170 199.435 ;
        RECT 88.440 198.580 88.700 198.900 ;
        RECT 87.970 194.985 88.250 195.355 ;
        RECT 88.040 194.140 88.180 194.985 ;
        RECT 87.980 193.820 88.240 194.140 ;
        RECT 88.440 193.820 88.700 194.140 ;
        RECT 88.500 190.740 88.640 193.820 ;
        RECT 88.440 190.420 88.700 190.740 ;
        RECT 89.420 189.120 89.560 203.000 ;
        RECT 89.880 194.820 90.020 209.800 ;
        RECT 90.340 208.760 90.480 221.250 ;
        RECT 92.570 221.070 92.850 221.570 ;
        RECT 95.790 221.070 96.070 221.570 ;
        RECT 99.010 221.070 99.290 221.570 ;
        RECT 102.230 221.080 102.510 221.570 ;
        RECT 102.760 221.250 104.280 221.390 ;
        RECT 102.760 221.080 102.900 221.250 ;
        RECT 102.230 221.070 102.900 221.080 ;
        RECT 90.730 216.065 91.010 216.435 ;
        RECT 90.280 208.440 90.540 208.760 ;
        RECT 90.280 206.740 90.540 207.060 ;
        RECT 89.820 194.500 90.080 194.820 ;
        RECT 89.820 193.480 90.080 193.800 ;
        RECT 89.880 192.440 90.020 193.480 ;
        RECT 89.820 192.120 90.080 192.440 ;
        RECT 90.340 189.235 90.480 206.740 ;
        RECT 90.800 202.640 90.940 216.065 ;
        RECT 92.120 207.760 92.380 208.080 ;
        RECT 92.180 206.040 92.320 207.760 ;
        RECT 92.120 205.720 92.380 206.040 ;
        RECT 92.640 205.360 92.780 221.070 ;
        RECT 95.860 214.960 96.000 221.070 ;
        RECT 95.400 214.820 96.000 214.960 ;
        RECT 95.400 208.080 95.540 214.820 ;
        RECT 95.800 209.460 96.060 209.780 ;
        RECT 95.860 208.420 96.000 209.460 ;
        RECT 95.800 208.100 96.060 208.420 ;
        RECT 97.640 208.100 97.900 208.420 ;
        RECT 95.340 207.760 95.600 208.080 ;
        RECT 94.880 207.420 95.140 207.740 ;
        RECT 94.940 206.235 95.080 207.420 ;
        RECT 95.860 207.310 96.000 208.100 ;
        RECT 96.260 207.310 96.520 207.400 ;
        RECT 95.860 207.170 96.520 207.310 ;
        RECT 96.260 207.080 96.520 207.170 ;
        RECT 95.340 206.970 95.600 207.060 ;
        RECT 95.340 206.830 96.000 206.970 ;
        RECT 95.340 206.740 95.600 206.830 ;
        RECT 93.960 205.720 94.220 206.040 ;
        RECT 94.870 205.865 95.150 206.235 ;
        RECT 92.580 205.040 92.840 205.360 ;
        RECT 94.020 205.020 94.160 205.720 ;
        RECT 93.960 204.700 94.220 205.020 ;
        RECT 94.880 204.760 95.140 205.020 ;
        RECT 94.880 204.700 95.540 204.760 ;
        RECT 94.940 204.620 95.540 204.700 ;
        RECT 92.580 204.020 92.840 204.340 ;
        RECT 93.960 204.020 94.220 204.340 ;
        RECT 90.740 202.320 91.000 202.640 ;
        RECT 90.740 199.940 91.000 200.260 ;
        RECT 89.420 188.980 90.020 189.120 ;
        RECT 86.140 188.040 86.400 188.360 ;
        RECT 87.120 188.300 87.720 188.440 ;
        RECT 87.980 188.380 88.240 188.700 ;
        RECT 88.440 188.380 88.700 188.700 ;
        RECT 89.360 188.380 89.620 188.700 ;
        RECT 86.200 187.000 86.340 188.040 ;
        RECT 86.140 186.680 86.400 187.000 ;
        RECT 86.600 186.680 86.860 187.000 ;
        RECT 86.660 185.835 86.800 186.680 ;
        RECT 85.680 185.320 85.940 185.640 ;
        RECT 86.590 185.465 86.870 185.835 ;
        RECT 85.210 184.785 85.490 185.155 ;
        RECT 84.300 183.960 84.560 184.280 ;
        RECT 85.210 184.105 85.490 184.475 ;
        RECT 84.760 183.170 85.020 183.260 ;
        RECT 85.280 183.170 85.420 184.105 ;
        RECT 84.760 183.030 85.420 183.170 ;
        RECT 84.760 182.940 85.020 183.030 ;
        RECT 85.740 182.580 85.880 185.320 ;
        RECT 87.120 184.280 87.260 188.300 ;
        RECT 87.520 187.700 87.780 188.020 ;
        RECT 87.060 183.960 87.320 184.280 ;
        RECT 87.120 183.795 87.260 183.960 ;
        RECT 87.050 183.425 87.330 183.795 ;
        RECT 86.590 182.745 86.870 183.115 ;
        RECT 84.760 182.260 85.020 182.580 ;
        RECT 85.680 182.260 85.940 182.580 ;
        RECT 84.820 180.540 84.960 182.260 ;
        RECT 86.130 181.385 86.410 181.755 ;
        RECT 86.200 180.880 86.340 181.385 ;
        RECT 86.140 180.560 86.400 180.880 ;
        RECT 86.660 180.540 86.800 182.745 ;
        RECT 87.050 181.385 87.330 181.755 ;
        RECT 87.060 181.240 87.320 181.385 ;
        RECT 84.760 180.220 85.020 180.540 ;
        RECT 86.600 180.220 86.860 180.540 ;
        RECT 83.840 178.520 84.100 178.840 ;
        RECT 82.980 177.820 83.120 177.985 ;
        RECT 83.380 177.840 83.640 178.160 ;
        RECT 84.750 177.985 85.030 178.355 ;
        RECT 82.920 177.500 83.180 177.820 ;
        RECT 83.370 177.305 83.650 177.675 ;
        RECT 83.440 176.030 83.580 177.305 ;
        RECT 83.840 177.160 84.100 177.480 ;
        RECT 82.980 175.890 83.580 176.030 ;
        RECT 82.980 174.760 83.120 175.890 ;
        RECT 83.380 175.120 83.640 175.440 ;
        RECT 82.920 174.440 83.180 174.760 ;
        RECT 82.920 173.080 83.180 173.400 ;
        RECT 82.980 172.380 83.120 173.080 ;
        RECT 82.920 172.235 83.180 172.380 ;
        RECT 82.910 171.865 83.190 172.235 ;
        RECT 83.440 168.155 83.580 175.120 ;
        RECT 83.900 170.340 84.040 177.160 ;
        RECT 84.300 176.820 84.560 177.140 ;
        RECT 84.360 176.120 84.500 176.820 ;
        RECT 84.300 175.800 84.560 176.120 ;
        RECT 84.820 175.440 84.960 177.985 ;
        RECT 85.680 177.510 85.940 177.830 ;
        RECT 85.220 176.820 85.480 177.140 ;
        RECT 84.760 175.120 85.020 175.440 ;
        RECT 84.300 174.100 84.560 174.420 ;
        RECT 84.760 174.330 85.020 174.420 ;
        RECT 85.280 174.330 85.420 176.820 ;
        RECT 84.760 174.190 85.420 174.330 ;
        RECT 84.760 174.100 85.020 174.190 ;
        RECT 83.840 170.020 84.100 170.340 ;
        RECT 83.370 167.785 83.650 168.155 ;
        RECT 82.920 167.300 83.180 167.620 ;
        RECT 66.820 155.400 67.080 155.720 ;
        RECT 73.710 155.545 73.990 155.915 ;
        RECT 82.460 155.740 82.720 156.060 ;
        RECT 82.980 155.210 83.120 167.300 ;
        RECT 83.840 166.620 84.100 166.940 ;
        RECT 83.380 165.940 83.640 166.260 ;
        RECT 83.440 161.160 83.580 165.940 ;
        RECT 83.900 162.520 84.040 166.620 ;
        RECT 83.840 162.200 84.100 162.520 ;
        RECT 84.360 161.160 84.500 174.100 ;
        RECT 84.820 173.060 84.960 174.100 ;
        RECT 85.740 173.400 85.880 177.510 ;
        RECT 86.600 176.820 86.860 177.140 ;
        RECT 86.660 174.420 86.800 176.820 ;
        RECT 87.050 175.265 87.330 175.635 ;
        RECT 87.120 174.760 87.260 175.265 ;
        RECT 87.060 174.440 87.320 174.760 ;
        RECT 86.600 174.100 86.860 174.420 ;
        RECT 85.680 173.080 85.940 173.400 ;
        RECT 87.060 173.080 87.320 173.400 ;
        RECT 84.760 172.740 85.020 173.060 ;
        RECT 86.140 171.720 86.400 172.040 ;
        RECT 86.200 170.000 86.340 171.720 ;
        RECT 87.120 171.700 87.260 173.080 ;
        RECT 87.060 171.380 87.320 171.700 ;
        RECT 85.220 169.680 85.480 170.000 ;
        RECT 86.140 169.680 86.400 170.000 ;
        RECT 85.280 169.515 85.420 169.680 ;
        RECT 85.210 169.145 85.490 169.515 ;
        RECT 84.750 168.465 85.030 168.835 ;
        RECT 84.820 166.940 84.960 168.465 ;
        RECT 86.140 167.640 86.400 167.960 ;
        RECT 84.760 166.620 85.020 166.940 ;
        RECT 85.220 166.620 85.480 166.940 ;
        RECT 85.280 165.435 85.420 166.620 ;
        RECT 85.210 165.065 85.490 165.435 ;
        RECT 85.220 163.900 85.480 164.220 ;
        RECT 85.280 163.540 85.420 163.900 ;
        RECT 85.220 163.220 85.480 163.540 ;
        RECT 83.380 160.840 83.640 161.160 ;
        RECT 83.840 160.840 84.100 161.160 ;
        RECT 84.300 160.840 84.560 161.160 ;
        RECT 83.900 159.120 84.040 160.840 ;
        RECT 83.840 158.800 84.100 159.120 ;
        RECT 86.200 155.210 86.340 167.640 ;
        RECT 87.580 166.940 87.720 187.700 ;
        RECT 88.040 174.760 88.180 188.380 ;
        RECT 88.500 187.195 88.640 188.380 ;
        RECT 88.430 186.825 88.710 187.195 ;
        RECT 89.420 185.835 89.560 188.380 ;
        RECT 89.350 185.465 89.630 185.835 ;
        RECT 89.880 185.210 90.020 188.980 ;
        RECT 90.270 188.865 90.550 189.235 ;
        RECT 90.340 188.700 90.480 188.865 ;
        RECT 90.280 188.380 90.540 188.700 ;
        RECT 90.280 186.570 90.540 186.660 ;
        RECT 90.800 186.570 90.940 199.940 ;
        RECT 91.200 196.715 91.460 196.860 ;
        RECT 91.190 196.345 91.470 196.715 ;
        RECT 92.640 194.675 92.780 204.020 ;
        RECT 94.020 202.980 94.160 204.020 ;
        RECT 93.960 202.660 94.220 202.980 ;
        RECT 94.880 202.835 95.140 202.980 ;
        RECT 93.500 202.320 93.760 202.640 ;
        RECT 94.870 202.465 95.150 202.835 ;
        RECT 93.040 201.300 93.300 201.620 ;
        RECT 93.100 199.580 93.240 201.300 ;
        RECT 93.560 200.115 93.700 202.320 ;
        RECT 93.960 201.980 94.220 202.300 ;
        RECT 93.490 199.745 93.770 200.115 ;
        RECT 93.040 199.260 93.300 199.580 ;
        RECT 93.560 196.860 93.700 199.745 ;
        RECT 94.020 198.900 94.160 201.980 ;
        RECT 94.880 201.640 95.140 201.960 ;
        RECT 94.410 199.745 94.690 200.115 ;
        RECT 93.960 198.580 94.220 198.900 ;
        RECT 94.020 197.200 94.160 198.580 ;
        RECT 93.960 196.880 94.220 197.200 ;
        RECT 93.500 196.540 93.760 196.860 ;
        RECT 94.480 196.520 94.620 199.745 ;
        RECT 94.940 198.075 95.080 201.640 ;
        RECT 95.400 200.115 95.540 204.620 ;
        RECT 95.860 202.640 96.000 206.830 ;
        RECT 97.700 205.020 97.840 208.100 ;
        RECT 99.080 208.080 99.220 221.070 ;
        RECT 102.300 220.940 102.900 221.070 ;
        RECT 104.140 208.840 104.280 221.250 ;
        RECT 105.450 221.070 105.730 221.570 ;
        RECT 108.670 221.070 108.950 221.570 ;
        RECT 111.890 221.070 112.170 221.570 ;
        RECT 115.110 221.070 115.390 221.570 ;
        RECT 118.330 221.070 118.610 221.570 ;
        RECT 121.550 221.080 121.830 221.570 ;
        RECT 122.080 221.250 123.140 221.390 ;
        RECT 122.080 221.080 122.220 221.250 ;
        RECT 121.550 221.070 122.220 221.080 ;
        RECT 104.140 208.760 104.740 208.840 ;
        RECT 100.860 208.440 101.120 208.760 ;
        RECT 104.140 208.700 104.800 208.760 ;
        RECT 104.540 208.440 104.800 208.700 ;
        RECT 99.020 207.760 99.280 208.080 ;
        RECT 100.400 207.760 100.660 208.080 ;
        RECT 98.100 207.080 98.360 207.400 ;
        RECT 98.160 205.020 98.300 207.080 ;
        RECT 98.620 206.660 99.680 206.800 ;
        RECT 98.620 206.040 98.760 206.660 ;
        RECT 98.560 205.720 98.820 206.040 ;
        RECT 96.320 204.680 97.380 204.760 ;
        RECT 97.640 204.700 97.900 205.020 ;
        RECT 98.100 204.700 98.360 205.020 ;
        RECT 96.260 204.620 97.380 204.680 ;
        RECT 96.260 204.360 96.520 204.620 ;
        RECT 96.720 204.020 96.980 204.340 ;
        RECT 95.800 202.320 96.060 202.640 ;
        RECT 96.780 202.550 96.920 204.020 ;
        RECT 97.240 203.400 97.380 204.620 ;
        RECT 97.240 203.260 98.300 203.400 ;
        RECT 97.240 202.835 97.380 203.260 ;
        RECT 98.160 202.980 98.300 203.260 ;
        RECT 96.320 202.410 96.920 202.550 ;
        RECT 97.170 202.465 97.450 202.835 ;
        RECT 97.640 202.660 97.900 202.980 ;
        RECT 98.100 202.660 98.360 202.980 ;
        RECT 99.020 202.660 99.280 202.980 ;
        RECT 95.800 201.300 96.060 201.620 ;
        RECT 95.330 199.745 95.610 200.115 ;
        RECT 95.860 199.435 96.000 201.300 ;
        RECT 95.340 198.920 95.600 199.240 ;
        RECT 95.790 199.065 96.070 199.435 ;
        RECT 94.870 197.705 95.150 198.075 ;
        RECT 95.400 197.880 95.540 198.920 ;
        RECT 94.940 197.200 95.080 197.705 ;
        RECT 95.340 197.560 95.600 197.880 ;
        RECT 94.880 196.880 95.140 197.200 ;
        RECT 94.420 196.200 94.680 196.520 ;
        RECT 93.960 195.860 94.220 196.180 ;
        RECT 94.020 194.820 94.160 195.860 ;
        RECT 96.320 195.355 96.460 202.410 ;
        RECT 97.180 201.870 97.440 201.960 ;
        RECT 97.700 201.870 97.840 202.660 ;
        RECT 97.180 201.730 97.840 201.870 ;
        RECT 97.180 201.640 97.440 201.730 ;
        RECT 98.560 199.830 98.820 199.920 ;
        RECT 98.160 199.690 98.820 199.830 ;
        RECT 97.180 198.580 97.440 198.900 ;
        RECT 97.240 197.540 97.380 198.580 ;
        RECT 97.180 197.220 97.440 197.540 ;
        RECT 96.720 196.880 96.980 197.200 ;
        RECT 96.250 194.985 96.530 195.355 ;
        RECT 91.200 194.160 91.460 194.480 ;
        RECT 91.650 194.305 91.930 194.675 ;
        RECT 92.570 194.305 92.850 194.675 ;
        RECT 93.960 194.500 94.220 194.820 ;
        RECT 91.660 194.160 91.920 194.305 ;
        RECT 91.260 193.800 91.400 194.160 ;
        RECT 91.200 193.480 91.460 193.800 ;
        RECT 92.640 192.440 92.780 194.305 ;
        RECT 93.040 194.160 93.300 194.480 ;
        RECT 92.120 192.120 92.380 192.440 ;
        RECT 92.580 192.120 92.840 192.440 ;
        RECT 92.180 191.955 92.320 192.120 ;
        RECT 91.660 191.440 91.920 191.760 ;
        RECT 92.110 191.585 92.390 191.955 ;
        RECT 93.100 191.840 93.240 194.160 ;
        RECT 92.640 191.700 93.240 191.840 ;
        RECT 94.020 191.760 94.160 194.500 ;
        RECT 95.340 193.140 95.600 193.460 ;
        RECT 94.870 192.265 95.150 192.635 ;
        RECT 95.400 192.440 95.540 193.140 ;
        RECT 94.880 192.120 95.140 192.265 ;
        RECT 95.340 192.120 95.600 192.440 ;
        RECT 96.780 192.350 96.920 196.880 ;
        RECT 97.180 196.540 97.440 196.860 ;
        RECT 96.320 192.210 96.920 192.350 ;
        RECT 91.720 189.915 91.860 191.440 ;
        RECT 92.640 191.330 92.780 191.700 ;
        RECT 93.500 191.440 93.760 191.760 ;
        RECT 93.960 191.440 94.220 191.760 ;
        RECT 92.180 191.190 92.780 191.330 ;
        RECT 92.180 190.595 92.320 191.190 ;
        RECT 93.040 190.760 93.300 191.080 ;
        RECT 92.110 190.225 92.390 190.595 ;
        RECT 92.580 190.420 92.840 190.740 ;
        RECT 91.650 189.545 91.930 189.915 ;
        RECT 91.200 187.700 91.460 188.020 ;
        RECT 90.280 186.430 90.940 186.570 ;
        RECT 90.280 186.340 90.540 186.430 ;
        RECT 90.280 185.890 90.540 185.980 ;
        RECT 90.280 185.750 90.940 185.890 ;
        RECT 90.280 185.660 90.540 185.750 ;
        RECT 89.420 185.070 90.020 185.210 ;
        RECT 88.430 183.425 88.710 183.795 ;
        RECT 88.500 183.260 88.640 183.425 ;
        RECT 88.440 182.940 88.700 183.260 ;
        RECT 88.430 180.705 88.710 181.075 ;
        RECT 88.500 179.770 88.640 180.705 ;
        RECT 88.500 179.630 89.100 179.770 ;
        RECT 88.440 178.520 88.700 178.840 ;
        RECT 88.500 178.355 88.640 178.520 ;
        RECT 88.430 177.985 88.710 178.355 ;
        RECT 88.960 178.160 89.100 179.630 ;
        RECT 88.900 177.840 89.160 178.160 ;
        RECT 88.900 176.820 89.160 177.140 ;
        RECT 89.420 176.995 89.560 185.070 ;
        RECT 89.810 182.745 90.090 183.115 ;
        RECT 89.880 182.580 90.020 182.745 ;
        RECT 89.820 182.260 90.080 182.580 ;
        RECT 90.270 181.385 90.550 181.755 ;
        RECT 90.340 181.220 90.480 181.385 ;
        RECT 89.810 180.705 90.090 181.075 ;
        RECT 90.280 180.900 90.540 181.220 ;
        RECT 89.820 180.560 90.080 180.705 ;
        RECT 90.800 180.280 90.940 185.750 ;
        RECT 91.260 183.260 91.400 187.700 ;
        RECT 91.650 185.465 91.930 185.835 ;
        RECT 92.180 185.720 92.320 190.225 ;
        RECT 92.640 189.040 92.780 190.420 ;
        RECT 92.580 188.720 92.840 189.040 ;
        RECT 92.580 187.700 92.840 188.020 ;
        RECT 92.640 187.000 92.780 187.700 ;
        RECT 92.580 186.680 92.840 187.000 ;
        RECT 92.580 186.230 92.840 186.320 ;
        RECT 93.100 186.230 93.240 190.760 ;
        RECT 93.560 189.720 93.700 191.440 ;
        RECT 94.420 190.595 94.680 190.740 ;
        RECT 94.410 190.225 94.690 190.595 ;
        RECT 93.500 189.400 93.760 189.720 ;
        RECT 94.940 188.700 95.080 192.120 ;
        RECT 96.320 190.740 96.460 192.210 ;
        RECT 96.720 191.440 96.980 191.760 ;
        RECT 97.240 191.670 97.380 196.540 ;
        RECT 97.630 196.345 97.910 196.715 ;
        RECT 97.700 192.635 97.840 196.345 ;
        RECT 98.160 194.480 98.300 199.690 ;
        RECT 98.560 199.600 98.820 199.690 ;
        RECT 98.560 198.920 98.820 199.240 ;
        RECT 98.620 197.540 98.760 198.920 ;
        RECT 98.560 197.220 98.820 197.540 ;
        RECT 99.080 195.160 99.220 202.660 ;
        RECT 99.540 201.960 99.680 206.660 ;
        RECT 99.940 205.720 100.200 206.040 ;
        RECT 99.480 201.640 99.740 201.960 ;
        RECT 100.000 201.620 100.140 205.720 ;
        RECT 100.460 204.680 100.600 207.760 ;
        RECT 100.400 204.360 100.660 204.680 ;
        RECT 99.940 201.300 100.200 201.620 ;
        RECT 99.470 199.745 99.750 200.115 ;
        RECT 99.540 199.580 99.680 199.745 ;
        RECT 99.480 199.260 99.740 199.580 ;
        RECT 99.480 196.880 99.740 197.200 ;
        RECT 99.540 196.035 99.680 196.880 ;
        RECT 99.940 196.715 100.200 196.860 ;
        RECT 99.930 196.345 100.210 196.715 ;
        RECT 99.470 195.665 99.750 196.035 ;
        RECT 99.940 195.860 100.200 196.180 ;
        RECT 100.000 195.355 100.140 195.860 ;
        RECT 99.020 194.840 99.280 195.160 ;
        RECT 99.930 194.985 100.210 195.355 ;
        RECT 98.100 194.160 98.360 194.480 ;
        RECT 99.480 193.820 99.740 194.140 ;
        RECT 99.020 193.480 99.280 193.800 ;
        RECT 97.630 192.265 97.910 192.635 ;
        RECT 97.640 191.670 97.900 191.760 ;
        RECT 97.240 191.530 97.900 191.670 ;
        RECT 97.640 191.440 97.900 191.530 ;
        RECT 96.260 190.420 96.520 190.740 ;
        RECT 95.340 188.720 95.600 189.040 ;
        RECT 93.500 188.040 93.760 188.360 ;
        RECT 93.950 188.185 94.230 188.555 ;
        RECT 94.880 188.380 95.140 188.700 ;
        RECT 93.960 188.040 94.220 188.185 ;
        RECT 93.560 187.875 93.700 188.040 ;
        RECT 93.490 187.505 93.770 187.875 ;
        RECT 92.580 186.090 93.240 186.230 ;
        RECT 93.490 186.145 93.770 186.515 ;
        RECT 92.580 186.000 92.840 186.090 ;
        RECT 92.180 185.580 92.780 185.720 ;
        RECT 91.720 183.940 91.860 185.465 ;
        RECT 92.640 185.300 92.780 185.580 ;
        RECT 93.040 185.320 93.300 185.640 ;
        RECT 92.120 184.980 92.380 185.300 ;
        RECT 92.580 184.980 92.840 185.300 ;
        RECT 91.660 183.620 91.920 183.940 ;
        RECT 92.180 183.600 92.320 184.980 ;
        RECT 92.120 183.280 92.380 183.600 ;
        RECT 91.200 182.940 91.460 183.260 ;
        RECT 92.640 183.170 92.780 184.980 ;
        RECT 93.100 183.680 93.240 185.320 ;
        RECT 93.560 184.280 93.700 186.145 ;
        RECT 93.500 183.960 93.760 184.280 ;
        RECT 93.100 183.540 93.700 183.680 ;
        RECT 94.020 183.600 94.160 188.040 ;
        RECT 94.420 187.700 94.680 188.020 ;
        RECT 95.400 187.930 95.540 188.720 ;
        RECT 96.320 188.555 96.460 190.420 ;
        RECT 96.250 188.185 96.530 188.555 ;
        RECT 96.780 188.020 96.920 191.440 ;
        RECT 95.400 187.790 96.460 187.930 ;
        RECT 94.480 185.640 94.620 187.700 ;
        RECT 94.870 186.825 95.150 187.195 ;
        RECT 96.320 186.910 96.460 187.790 ;
        RECT 96.720 187.700 96.980 188.020 ;
        RECT 97.700 187.875 97.840 191.440 ;
        RECT 99.080 191.080 99.220 193.480 ;
        RECT 98.100 190.990 98.360 191.080 ;
        RECT 98.100 190.850 98.760 190.990 ;
        RECT 98.100 190.760 98.360 190.850 ;
        RECT 98.620 189.380 98.760 190.850 ;
        RECT 99.020 190.760 99.280 191.080 ;
        RECT 98.100 189.060 98.360 189.380 ;
        RECT 98.560 189.060 98.820 189.380 ;
        RECT 97.630 187.505 97.910 187.875 ;
        RECT 97.180 186.910 97.440 187.000 ;
        RECT 94.940 186.570 95.080 186.825 ;
        RECT 96.320 186.770 97.440 186.910 ;
        RECT 97.180 186.680 97.440 186.770 ;
        RECT 95.340 186.570 95.600 186.660 ;
        RECT 94.940 186.430 95.600 186.570 ;
        RECT 94.420 185.320 94.680 185.640 ;
        RECT 94.410 184.785 94.690 185.155 ;
        RECT 94.480 183.940 94.620 184.785 ;
        RECT 94.420 183.620 94.680 183.940 ;
        RECT 93.040 183.170 93.300 183.260 ;
        RECT 92.640 183.030 93.300 183.170 ;
        RECT 93.040 182.940 93.300 183.030 ;
        RECT 91.260 181.560 91.400 182.940 ;
        RECT 93.560 182.830 93.700 183.540 ;
        RECT 93.960 183.280 94.220 183.600 ;
        RECT 94.940 183.260 95.080 186.430 ;
        RECT 95.340 186.340 95.600 186.430 ;
        RECT 95.800 186.000 96.060 186.320 ;
        RECT 97.170 186.145 97.450 186.515 ;
        RECT 97.180 186.000 97.440 186.145 ;
        RECT 95.860 185.300 96.000 186.000 ;
        RECT 96.720 185.660 96.980 185.980 ;
        RECT 96.260 185.320 96.520 185.640 ;
        RECT 95.800 184.980 96.060 185.300 ;
        RECT 96.320 185.155 96.460 185.320 ;
        RECT 96.250 184.785 96.530 185.155 ;
        RECT 96.780 184.280 96.920 185.660 ;
        RECT 97.180 185.320 97.440 185.640 ;
        RECT 95.340 183.960 95.600 184.280 ;
        RECT 96.720 183.960 96.980 184.280 ;
        RECT 94.880 182.940 95.140 183.260 ;
        RECT 93.560 182.690 94.160 182.830 ;
        RECT 93.040 182.490 93.300 182.580 ;
        RECT 93.040 182.350 93.700 182.490 ;
        RECT 93.040 182.260 93.300 182.350 ;
        RECT 93.560 181.560 93.700 182.350 ;
        RECT 91.200 181.240 91.460 181.560 ;
        RECT 93.500 181.240 93.760 181.560 ;
        RECT 94.020 181.220 94.160 182.690 ;
        RECT 94.870 182.065 95.150 182.435 ;
        RECT 93.960 180.900 94.220 181.220 ;
        RECT 91.660 180.790 91.920 180.880 ;
        RECT 91.660 180.650 93.240 180.790 ;
        RECT 91.660 180.560 91.920 180.650 ;
        RECT 90.800 180.200 92.780 180.280 ;
        RECT 90.280 179.880 90.540 180.200 ;
        RECT 90.800 180.140 92.840 180.200 ;
        RECT 92.580 179.880 92.840 180.140 ;
        RECT 89.820 179.540 90.080 179.860 ;
        RECT 89.880 178.355 90.020 179.540 ;
        RECT 90.340 178.750 90.480 179.880 ;
        RECT 90.740 179.715 91.000 179.860 ;
        RECT 90.730 179.345 91.010 179.715 ;
        RECT 91.660 178.750 91.920 178.840 ;
        RECT 90.340 178.610 91.920 178.750 ;
        RECT 91.660 178.520 91.920 178.610 ;
        RECT 89.810 177.985 90.090 178.355 ;
        RECT 91.200 177.160 91.460 177.480 ;
        RECT 91.660 177.160 91.920 177.480 ;
        RECT 92.120 177.160 92.380 177.480 ;
        RECT 88.430 175.945 88.710 176.315 ;
        RECT 88.500 175.440 88.640 175.945 ;
        RECT 88.440 175.120 88.700 175.440 ;
        RECT 87.980 174.440 88.240 174.760 ;
        RECT 88.500 173.400 88.640 175.120 ;
        RECT 88.440 173.080 88.700 173.400 ;
        RECT 88.960 172.970 89.100 176.820 ;
        RECT 89.350 176.625 89.630 176.995 ;
        RECT 89.820 176.820 90.080 177.140 ;
        RECT 90.280 176.820 90.540 177.140 ;
        RECT 91.260 176.995 91.400 177.160 ;
        RECT 89.360 174.780 89.620 175.100 ;
        RECT 89.420 173.480 89.560 174.780 ;
        RECT 89.880 174.160 90.020 176.820 ;
        RECT 90.340 175.780 90.480 176.820 ;
        RECT 91.190 176.625 91.470 176.995 ;
        RECT 91.720 176.315 91.860 177.160 ;
        RECT 91.200 175.800 91.460 176.120 ;
        RECT 91.650 175.945 91.930 176.315 ;
        RECT 90.280 175.460 90.540 175.780 ;
        RECT 91.260 175.440 91.400 175.800 ;
        RECT 91.200 175.120 91.460 175.440 ;
        RECT 92.180 174.840 92.320 177.160 ;
        RECT 92.570 175.945 92.850 176.315 ;
        RECT 92.640 175.440 92.780 175.945 ;
        RECT 92.580 175.120 92.840 175.440 ;
        RECT 92.180 174.700 92.780 174.840 ;
        RECT 92.110 174.160 92.390 174.275 ;
        RECT 92.640 174.160 92.780 174.700 ;
        RECT 89.880 174.020 90.480 174.160 ;
        RECT 89.420 173.400 90.020 173.480 ;
        RECT 89.420 173.340 90.080 173.400 ;
        RECT 89.820 173.080 90.080 173.340 ;
        RECT 89.360 172.970 89.620 173.060 ;
        RECT 88.960 172.830 89.620 172.970 ;
        RECT 89.360 172.740 89.620 172.830 ;
        RECT 88.440 172.235 88.700 172.380 ;
        RECT 88.430 171.865 88.710 172.235 ;
        RECT 89.360 171.720 89.620 172.040 ;
        RECT 88.440 171.380 88.700 171.700 ;
        RECT 88.500 170.340 88.640 171.380 ;
        RECT 89.420 170.875 89.560 171.720 ;
        RECT 89.350 170.505 89.630 170.875 ;
        RECT 88.440 170.020 88.700 170.340 ;
        RECT 89.820 169.680 90.080 170.000 ;
        RECT 87.980 169.340 88.240 169.660 ;
        RECT 88.440 169.340 88.700 169.660 ;
        RECT 89.360 169.340 89.620 169.660 ;
        RECT 86.600 166.620 86.860 166.940 ;
        RECT 87.520 166.620 87.780 166.940 ;
        RECT 86.660 163.880 86.800 166.620 ;
        RECT 88.040 165.435 88.180 169.340 ;
        RECT 87.970 165.065 88.250 165.435 ;
        RECT 86.600 163.560 86.860 163.880 ;
        RECT 88.500 163.540 88.640 169.340 ;
        RECT 89.420 166.940 89.560 169.340 ;
        RECT 89.360 166.620 89.620 166.940 ;
        RECT 88.900 165.940 89.160 166.260 ;
        RECT 88.960 163.880 89.100 165.940 ;
        RECT 88.900 163.560 89.160 163.880 ;
        RECT 88.440 163.220 88.700 163.540 ;
        RECT 89.420 162.860 89.560 166.620 ;
        RECT 89.880 165.240 90.020 169.680 ;
        RECT 89.820 164.920 90.080 165.240 ;
        RECT 90.340 164.220 90.480 174.020 ;
        RECT 92.110 174.020 92.780 174.160 ;
        RECT 92.110 173.905 92.390 174.020 ;
        RECT 92.580 172.120 92.840 172.380 ;
        RECT 91.260 172.060 92.840 172.120 ;
        RECT 91.260 171.980 92.780 172.060 ;
        RECT 91.260 171.950 91.400 171.980 ;
        RECT 90.800 171.810 91.400 171.950 ;
        RECT 90.800 170.590 90.940 171.810 ;
        RECT 92.120 171.380 92.380 171.700 ;
        RECT 92.580 171.380 92.840 171.700 ;
        RECT 91.200 170.590 91.460 170.680 ;
        RECT 90.800 170.450 91.460 170.590 ;
        RECT 91.650 170.505 91.930 170.875 ;
        RECT 92.180 170.680 92.320 171.380 ;
        RECT 91.200 170.360 91.460 170.450 ;
        RECT 91.660 170.360 91.920 170.505 ;
        RECT 92.120 170.360 92.380 170.680 ;
        RECT 91.200 168.660 91.460 168.980 ;
        RECT 91.260 165.240 91.400 168.660 ;
        RECT 91.720 166.260 91.860 170.360 ;
        RECT 92.180 166.600 92.320 170.360 ;
        RECT 92.640 170.340 92.780 171.380 ;
        RECT 92.580 170.020 92.840 170.340 ;
        RECT 93.100 168.980 93.240 180.650 ;
        RECT 93.500 180.220 93.760 180.540 ;
        RECT 93.560 179.035 93.700 180.220 ;
        RECT 94.020 179.770 94.160 180.900 ;
        RECT 94.420 179.770 94.680 179.860 ;
        RECT 94.020 179.630 94.680 179.770 ;
        RECT 94.420 179.540 94.680 179.630 ;
        RECT 93.490 178.665 93.770 179.035 ;
        RECT 94.420 178.520 94.680 178.840 ;
        RECT 93.960 177.500 94.220 177.820 ;
        RECT 93.500 175.120 93.760 175.440 ;
        RECT 93.560 173.400 93.700 175.120 ;
        RECT 94.020 174.760 94.160 177.500 ;
        RECT 94.480 177.140 94.620 178.520 ;
        RECT 94.420 176.820 94.680 177.140 ;
        RECT 94.420 175.800 94.680 176.120 ;
        RECT 93.960 174.440 94.220 174.760 ;
        RECT 94.480 174.160 94.620 175.800 ;
        RECT 94.940 175.440 95.080 182.065 ;
        RECT 95.400 181.220 95.540 183.960 ;
        RECT 97.240 183.680 97.380 185.320 ;
        RECT 96.320 183.540 97.380 183.680 ;
        RECT 97.700 183.600 97.840 187.505 ;
        RECT 95.790 181.385 96.070 181.755 ;
        RECT 95.340 180.900 95.600 181.220 ;
        RECT 95.860 180.395 96.000 181.385 ;
        RECT 96.320 180.540 96.460 183.540 ;
        RECT 97.640 183.280 97.900 183.600 ;
        RECT 97.180 182.600 97.440 182.920 ;
        RECT 96.720 180.560 96.980 180.880 ;
        RECT 95.790 180.025 96.070 180.395 ;
        RECT 96.260 180.220 96.520 180.540 ;
        RECT 95.790 177.985 96.070 178.355 ;
        RECT 95.860 177.820 96.000 177.985 ;
        RECT 95.800 177.730 96.060 177.820 ;
        RECT 95.400 177.590 96.060 177.730 ;
        RECT 94.880 175.120 95.140 175.440 ;
        RECT 94.880 174.440 95.140 174.760 ;
        RECT 94.020 174.020 94.620 174.160 ;
        RECT 93.500 173.080 93.760 173.400 ;
        RECT 94.020 172.720 94.160 174.020 ;
        RECT 94.410 173.225 94.690 173.595 ;
        RECT 93.960 172.400 94.220 172.720 ;
        RECT 94.480 172.120 94.620 173.225 ;
        RECT 93.560 171.980 94.620 172.120 ;
        RECT 93.040 168.660 93.300 168.980 ;
        RECT 92.580 166.960 92.840 167.280 ;
        RECT 92.120 166.280 92.380 166.600 ;
        RECT 91.660 165.940 91.920 166.260 ;
        RECT 91.200 164.920 91.460 165.240 ;
        RECT 90.280 163.900 90.540 164.220 ;
        RECT 89.360 162.540 89.620 162.860 ;
        RECT 89.360 158.800 89.620 159.120 ;
        RECT 89.420 155.210 89.560 158.800 ;
        RECT 92.640 155.210 92.780 166.960 ;
        RECT 93.100 165.435 93.240 168.660 ;
        RECT 93.030 165.065 93.310 165.435 ;
        RECT 93.560 165.240 93.700 171.980 ;
        RECT 94.420 171.610 94.680 171.700 ;
        RECT 94.020 171.470 94.680 171.610 ;
        RECT 94.020 169.320 94.160 171.470 ;
        RECT 94.420 171.380 94.680 171.470 ;
        RECT 94.420 170.360 94.680 170.680 ;
        RECT 94.480 170.195 94.620 170.360 ;
        RECT 94.410 169.825 94.690 170.195 ;
        RECT 93.965 169.000 94.225 169.320 ;
        RECT 94.410 167.785 94.690 168.155 ;
        RECT 94.480 166.260 94.620 167.785 ;
        RECT 94.420 165.940 94.680 166.260 ;
        RECT 93.500 164.920 93.760 165.240 ;
        RECT 94.940 164.560 95.080 174.440 ;
        RECT 95.400 173.595 95.540 177.590 ;
        RECT 95.800 177.500 96.060 177.590 ;
        RECT 96.320 175.440 96.460 180.220 ;
        RECT 96.780 178.070 96.920 180.560 ;
        RECT 97.240 178.840 97.380 182.600 ;
        RECT 98.160 182.320 98.300 189.060 ;
        RECT 99.540 189.040 99.680 193.820 ;
        RECT 100.000 191.420 100.140 194.985 ;
        RECT 100.460 194.390 100.600 204.360 ;
        RECT 100.920 202.640 101.060 208.440 ;
        RECT 103.680 208.020 105.200 208.160 ;
        RECT 102.230 206.545 102.510 206.915 ;
        RECT 103.160 206.740 103.420 207.060 ;
        RECT 102.300 204.680 102.440 206.545 ;
        RECT 103.220 205.360 103.360 206.740 ;
        RECT 103.160 205.040 103.420 205.360 ;
        RECT 102.240 204.360 102.500 204.680 ;
        RECT 103.220 202.640 103.360 205.040 ;
        RECT 103.680 204.340 103.820 208.020 ;
        RECT 104.540 207.420 104.800 207.740 ;
        RECT 104.080 207.080 104.340 207.400 ;
        RECT 104.140 205.020 104.280 207.080 ;
        RECT 104.080 204.700 104.340 205.020 ;
        RECT 103.620 204.020 103.880 204.340 ;
        RECT 100.860 202.320 101.120 202.640 ;
        RECT 103.160 202.320 103.420 202.640 ;
        RECT 103.620 202.320 103.880 202.640 ;
        RECT 101.780 201.980 102.040 202.300 ;
        RECT 101.320 201.640 101.580 201.960 ;
        RECT 100.860 201.300 101.120 201.620 ;
        RECT 100.920 196.520 101.060 201.300 ;
        RECT 101.380 199.920 101.520 201.640 ;
        RECT 101.320 199.600 101.580 199.920 ;
        RECT 101.840 198.075 101.980 201.980 ;
        RECT 102.700 201.300 102.960 201.620 ;
        RECT 102.760 199.240 102.900 201.300 ;
        RECT 102.700 198.920 102.960 199.240 ;
        RECT 101.770 197.705 102.050 198.075 ;
        RECT 101.840 197.200 101.980 197.705 ;
        RECT 101.780 196.880 102.040 197.200 ;
        RECT 102.240 196.880 102.500 197.200 ;
        RECT 100.860 196.200 101.120 196.520 ;
        RECT 100.460 194.250 101.060 194.390 ;
        RECT 100.400 193.480 100.660 193.800 ;
        RECT 99.940 191.100 100.200 191.420 ;
        RECT 99.940 190.420 100.200 190.740 ;
        RECT 99.020 188.720 99.280 189.040 ;
        RECT 99.480 188.720 99.740 189.040 ;
        RECT 98.560 187.700 98.820 188.020 ;
        RECT 98.620 185.980 98.760 187.700 ;
        RECT 99.080 186.320 99.220 188.720 ;
        RECT 100.000 188.700 100.140 190.420 ;
        RECT 99.940 188.380 100.200 188.700 ;
        RECT 99.480 187.930 99.740 188.020 ;
        RECT 100.460 187.930 100.600 193.480 ;
        RECT 99.480 187.875 100.600 187.930 ;
        RECT 99.470 187.790 100.600 187.875 ;
        RECT 99.470 187.505 99.750 187.790 ;
        RECT 99.480 186.340 99.740 186.660 ;
        RECT 99.940 186.340 100.200 186.660 ;
        RECT 99.020 186.000 99.280 186.320 ;
        RECT 98.560 185.660 98.820 185.980 ;
        RECT 98.560 183.960 98.820 184.280 ;
        RECT 98.620 182.920 98.760 183.960 ;
        RECT 99.080 183.940 99.220 186.000 ;
        RECT 99.020 183.620 99.280 183.940 ;
        RECT 98.560 182.600 98.820 182.920 ;
        RECT 99.080 182.435 99.220 183.620 ;
        RECT 99.540 182.580 99.680 186.340 ;
        RECT 100.000 184.280 100.140 186.340 ;
        RECT 99.940 183.960 100.200 184.280 ;
        RECT 100.920 183.680 101.060 194.250 ;
        RECT 101.320 194.160 101.580 194.480 ;
        RECT 100.000 183.540 101.060 183.680 ;
        RECT 98.160 182.180 98.760 182.320 ;
        RECT 98.100 180.900 98.360 181.220 ;
        RECT 97.640 179.880 97.900 180.200 ;
        RECT 97.180 178.520 97.440 178.840 ;
        RECT 97.700 178.160 97.840 179.880 ;
        RECT 97.180 178.070 97.440 178.160 ;
        RECT 96.780 177.930 97.440 178.070 ;
        RECT 97.180 177.840 97.440 177.930 ;
        RECT 97.640 177.840 97.900 178.160 ;
        RECT 97.180 177.160 97.440 177.480 ;
        RECT 97.630 177.305 97.910 177.675 ;
        RECT 97.640 177.160 97.900 177.305 ;
        RECT 97.240 175.440 97.380 177.160 ;
        RECT 95.800 175.120 96.060 175.440 ;
        RECT 96.260 175.120 96.520 175.440 ;
        RECT 97.180 175.120 97.440 175.440 ;
        RECT 95.330 173.225 95.610 173.595 ;
        RECT 95.340 172.400 95.600 172.720 ;
        RECT 95.400 170.340 95.540 172.400 ;
        RECT 95.340 170.020 95.600 170.340 ;
        RECT 95.860 167.960 96.000 175.120 ;
        RECT 96.320 172.720 96.460 175.120 ;
        RECT 96.710 174.585 96.990 174.955 ;
        RECT 97.630 174.585 97.910 174.955 ;
        RECT 96.780 173.060 96.920 174.585 ;
        RECT 97.170 173.225 97.450 173.595 ;
        RECT 97.700 173.400 97.840 174.585 ;
        RECT 96.720 172.740 96.980 173.060 ;
        RECT 96.260 172.400 96.520 172.720 ;
        RECT 97.240 172.380 97.380 173.225 ;
        RECT 97.640 173.080 97.900 173.400 ;
        RECT 97.640 172.400 97.900 172.720 ;
        RECT 98.160 172.630 98.300 180.900 ;
        RECT 98.620 177.820 98.760 182.180 ;
        RECT 99.010 182.065 99.290 182.435 ;
        RECT 99.480 182.260 99.740 182.580 ;
        RECT 99.010 181.385 99.290 181.755 ;
        RECT 98.560 177.500 98.820 177.820 ;
        RECT 98.620 176.315 98.760 177.500 ;
        RECT 98.550 175.945 98.830 176.315 ;
        RECT 98.560 174.100 98.820 174.420 ;
        RECT 99.080 174.330 99.220 181.385 ;
        RECT 100.000 178.240 100.140 183.540 ;
        RECT 100.860 182.940 101.120 183.260 ;
        RECT 100.390 182.065 100.670 182.435 ;
        RECT 100.460 181.560 100.600 182.065 ;
        RECT 100.400 181.240 100.660 181.560 ;
        RECT 100.400 180.560 100.660 180.880 ;
        RECT 100.460 179.860 100.600 180.560 ;
        RECT 100.400 179.540 100.660 179.860 ;
        RECT 100.400 178.520 100.660 178.840 ;
        RECT 100.920 178.750 101.060 182.940 ;
        RECT 101.380 182.580 101.520 194.160 ;
        RECT 101.780 193.480 102.040 193.800 ;
        RECT 101.840 191.080 101.980 193.480 ;
        RECT 102.300 191.420 102.440 196.880 ;
        RECT 102.760 196.860 102.900 198.920 ;
        RECT 103.680 198.640 103.820 202.320 ;
        RECT 104.140 202.300 104.280 204.700 ;
        RECT 104.600 202.980 104.740 207.420 ;
        RECT 105.060 204.930 105.200 208.020 ;
        RECT 105.520 207.400 105.660 221.070 ;
        RECT 108.740 209.635 108.880 221.070 ;
        RECT 108.670 209.265 108.950 209.635 ;
        RECT 111.960 208.760 112.100 221.070 ;
        RECT 115.180 208.760 115.320 221.070 ;
        RECT 118.400 210.880 118.540 221.070 ;
        RECT 121.620 220.940 122.220 221.070 ;
        RECT 118.400 210.740 119.000 210.880 ;
        RECT 118.340 210.140 118.600 210.460 ;
        RECT 111.900 208.440 112.160 208.760 ;
        RECT 115.120 208.440 115.380 208.760 ;
        RECT 108.680 208.100 108.940 208.420 ;
        RECT 106.380 207.760 106.640 208.080 ;
        RECT 105.460 207.080 105.720 207.400 ;
        RECT 105.920 206.740 106.180 207.060 ;
        RECT 105.980 205.360 106.120 206.740 ;
        RECT 105.920 205.040 106.180 205.360 ;
        RECT 106.440 205.020 106.580 207.760 ;
        RECT 108.220 207.080 108.480 207.400 ;
        RECT 107.760 205.040 108.020 205.360 ;
        RECT 105.460 204.930 105.720 205.020 ;
        RECT 105.060 204.790 105.720 204.930 ;
        RECT 105.460 204.700 105.720 204.790 ;
        RECT 106.380 204.700 106.640 205.020 ;
        RECT 105.920 204.360 106.180 204.680 ;
        RECT 104.540 202.660 104.800 202.980 ;
        RECT 104.990 202.465 105.270 202.835 ;
        RECT 105.000 202.320 105.260 202.465 ;
        RECT 104.080 201.980 104.340 202.300 ;
        RECT 103.220 198.500 103.820 198.640 ;
        RECT 102.700 196.540 102.960 196.860 ;
        RECT 102.700 194.500 102.960 194.820 ;
        RECT 102.760 191.760 102.900 194.500 ;
        RECT 102.700 191.440 102.960 191.760 ;
        RECT 102.240 191.100 102.500 191.420 ;
        RECT 101.780 190.760 102.040 191.080 ;
        RECT 101.780 189.060 102.040 189.380 ;
        RECT 101.840 185.640 101.980 189.060 ;
        RECT 102.240 188.720 102.500 189.040 ;
        RECT 102.300 186.570 102.440 188.720 ;
        RECT 103.220 188.440 103.360 198.500 ;
        RECT 103.620 197.560 103.880 197.880 ;
        RECT 103.680 194.140 103.820 197.560 ;
        RECT 104.540 196.540 104.800 196.860 ;
        RECT 103.620 193.820 103.880 194.140 ;
        RECT 104.080 191.440 104.340 191.760 ;
        RECT 103.620 189.400 103.880 189.720 ;
        RECT 102.760 188.300 103.360 188.440 ;
        RECT 102.760 187.195 102.900 188.300 ;
        RECT 103.160 187.700 103.420 188.020 ;
        RECT 102.690 186.825 102.970 187.195 ;
        RECT 102.300 186.430 102.900 186.570 ;
        RECT 101.780 185.320 102.040 185.640 ;
        RECT 102.230 185.465 102.510 185.835 ;
        RECT 102.300 184.360 102.440 185.465 ;
        RECT 101.840 184.220 102.440 184.360 ;
        RECT 101.320 182.260 101.580 182.580 ;
        RECT 101.320 178.750 101.580 178.840 ;
        RECT 100.920 178.610 101.580 178.750 ;
        RECT 99.540 178.100 100.140 178.240 ;
        RECT 99.540 176.120 99.680 178.100 ;
        RECT 99.940 177.500 100.200 177.820 ;
        RECT 100.000 176.120 100.140 177.500 ;
        RECT 99.480 175.800 99.740 176.120 ;
        RECT 99.940 175.800 100.200 176.120 ;
        RECT 99.540 175.440 99.680 175.800 ;
        RECT 99.480 175.120 99.740 175.440 ;
        RECT 100.460 174.955 100.600 178.520 ;
        RECT 99.470 174.840 99.750 174.955 ;
        RECT 99.470 174.760 100.140 174.840 ;
        RECT 99.470 174.700 100.200 174.760 ;
        RECT 99.470 174.585 99.750 174.700 ;
        RECT 99.940 174.440 100.200 174.700 ;
        RECT 100.390 174.585 100.670 174.955 ;
        RECT 99.080 174.190 99.680 174.330 ;
        RECT 98.620 173.400 98.760 174.100 ;
        RECT 98.560 173.080 98.820 173.400 ;
        RECT 99.540 173.060 99.680 174.190 ;
        RECT 99.020 172.740 99.280 173.060 ;
        RECT 99.480 172.740 99.740 173.060 ;
        RECT 100.920 172.915 101.060 178.610 ;
        RECT 101.320 178.520 101.580 178.610 ;
        RECT 101.840 176.880 101.980 184.220 ;
        RECT 102.240 183.620 102.500 183.940 ;
        RECT 102.300 180.880 102.440 183.620 ;
        RECT 102.760 183.260 102.900 186.430 ;
        RECT 103.220 186.320 103.360 187.700 ;
        RECT 103.160 186.000 103.420 186.320 ;
        RECT 103.680 185.835 103.820 189.400 ;
        RECT 104.140 189.380 104.280 191.440 ;
        RECT 104.080 189.060 104.340 189.380 ;
        RECT 104.140 188.555 104.280 189.060 ;
        RECT 104.070 188.185 104.350 188.555 ;
        RECT 104.070 187.505 104.350 187.875 ;
        RECT 103.160 185.320 103.420 185.640 ;
        RECT 103.610 185.465 103.890 185.835 ;
        RECT 103.220 184.360 103.360 185.320 ;
        RECT 103.220 184.280 103.820 184.360 ;
        RECT 103.220 184.220 103.880 184.280 ;
        RECT 103.620 183.960 103.880 184.220 ;
        RECT 102.700 182.940 102.960 183.260 ;
        RECT 103.160 182.940 103.420 183.260 ;
        RECT 103.220 181.220 103.360 182.940 ;
        RECT 104.140 182.830 104.280 187.505 ;
        RECT 104.600 185.640 104.740 196.540 ;
        RECT 105.060 190.740 105.200 202.320 ;
        RECT 105.460 201.640 105.720 201.960 ;
        RECT 105.520 199.580 105.660 201.640 ;
        RECT 105.980 199.580 106.120 204.360 ;
        RECT 106.380 202.660 106.640 202.980 ;
        RECT 106.440 200.115 106.580 202.660 ;
        RECT 106.840 202.320 107.100 202.640 ;
        RECT 106.900 202.155 107.040 202.320 ;
        RECT 106.830 201.785 107.110 202.155 ;
        RECT 106.370 199.745 106.650 200.115 ;
        RECT 105.460 199.260 105.720 199.580 ;
        RECT 105.920 199.260 106.180 199.580 ;
        RECT 105.980 197.200 106.120 199.260 ;
        RECT 106.440 199.240 106.580 199.745 ;
        RECT 106.380 198.920 106.640 199.240 ;
        RECT 105.920 196.880 106.180 197.200 ;
        RECT 106.440 196.180 106.580 198.920 ;
        RECT 107.820 197.880 107.960 205.040 ;
        RECT 108.280 205.020 108.420 207.080 ;
        RECT 108.740 205.020 108.880 208.100 ;
        RECT 110.060 207.760 110.320 208.080 ;
        RECT 114.200 207.990 114.460 208.080 ;
        RECT 111.960 207.850 114.460 207.990 ;
        RECT 109.130 206.545 109.410 206.915 ;
        RECT 108.220 204.700 108.480 205.020 ;
        RECT 108.680 204.700 108.940 205.020 ;
        RECT 108.280 202.980 108.420 204.700 ;
        RECT 108.740 202.980 108.880 204.700 ;
        RECT 109.200 204.340 109.340 206.545 ;
        RECT 110.120 206.040 110.260 207.760 ;
        RECT 110.060 205.720 110.320 206.040 ;
        RECT 110.520 205.720 110.780 206.040 ;
        RECT 110.060 204.700 110.320 205.020 ;
        RECT 109.140 204.020 109.400 204.340 ;
        RECT 108.220 202.660 108.480 202.980 ;
        RECT 108.680 202.660 108.940 202.980 ;
        RECT 109.600 202.320 109.860 202.640 ;
        RECT 108.680 201.300 108.940 201.620 ;
        RECT 108.740 199.580 108.880 201.300 ;
        RECT 108.680 199.260 108.940 199.580 ;
        RECT 109.140 199.260 109.400 199.580 ;
        RECT 107.760 197.560 108.020 197.880 ;
        RECT 107.760 196.540 108.020 196.860 ;
        RECT 105.980 196.040 106.580 196.180 ;
        RECT 105.980 194.480 106.120 196.040 ;
        RECT 105.920 194.160 106.180 194.480 ;
        RECT 106.380 194.160 106.640 194.480 ;
        RECT 106.440 193.460 106.580 194.160 ;
        RECT 107.300 194.050 107.560 194.140 ;
        RECT 107.820 194.050 107.960 196.540 ;
        RECT 107.300 193.910 107.960 194.050 ;
        RECT 107.300 193.820 107.560 193.910 ;
        RECT 105.460 193.140 105.720 193.460 ;
        RECT 106.380 193.140 106.640 193.460 ;
        RECT 106.840 193.140 107.100 193.460 ;
        RECT 105.000 190.420 105.260 190.740 ;
        RECT 105.060 186.515 105.200 190.420 ;
        RECT 104.990 186.145 105.270 186.515 ;
        RECT 104.540 185.320 104.800 185.640 ;
        RECT 105.000 184.980 105.260 185.300 ;
        RECT 105.060 183.600 105.200 184.980 ;
        RECT 105.000 183.280 105.260 183.600 ;
        RECT 105.000 182.830 105.260 182.920 ;
        RECT 104.140 182.690 105.260 182.830 ;
        RECT 105.000 182.600 105.260 182.690 ;
        RECT 103.160 180.900 103.420 181.220 ;
        RECT 102.240 180.560 102.500 180.880 ;
        RECT 102.700 180.560 102.960 180.880 ;
        RECT 102.240 178.520 102.500 178.840 ;
        RECT 102.300 177.820 102.440 178.520 ;
        RECT 102.760 178.500 102.900 180.560 ;
        RECT 103.160 179.540 103.420 179.860 ;
        RECT 104.080 179.540 104.340 179.860 ;
        RECT 102.700 178.180 102.960 178.500 ;
        RECT 103.220 177.820 103.360 179.540 ;
        RECT 103.620 178.180 103.880 178.500 ;
        RECT 103.680 177.820 103.820 178.180 ;
        RECT 102.240 177.500 102.500 177.820 ;
        RECT 103.160 177.500 103.420 177.820 ;
        RECT 103.620 177.500 103.880 177.820 ;
        RECT 103.220 176.995 103.360 177.500 ;
        RECT 101.380 176.740 101.980 176.880 ;
        RECT 98.160 172.490 98.760 172.630 ;
        RECT 97.180 172.060 97.440 172.380 ;
        RECT 96.720 171.380 96.980 171.700 ;
        RECT 96.250 170.505 96.530 170.875 ;
        RECT 96.260 170.360 96.520 170.505 ;
        RECT 96.250 169.825 96.530 170.195 ;
        RECT 96.260 169.680 96.520 169.825 ;
        RECT 96.260 169.000 96.520 169.320 ;
        RECT 95.800 167.640 96.060 167.960 ;
        RECT 95.340 167.300 95.600 167.620 ;
        RECT 95.400 166.000 95.540 167.300 ;
        RECT 96.320 166.600 96.460 169.000 ;
        RECT 96.260 166.280 96.520 166.600 ;
        RECT 96.780 166.000 96.920 171.380 ;
        RECT 97.180 167.300 97.440 167.620 ;
        RECT 97.240 166.260 97.380 167.300 ;
        RECT 95.400 165.860 96.920 166.000 ;
        RECT 97.180 165.940 97.440 166.260 ;
        RECT 96.780 164.560 96.920 165.860 ;
        RECT 94.880 164.240 95.140 164.560 ;
        RECT 96.720 164.240 96.980 164.560 ;
        RECT 97.700 163.880 97.840 172.400 ;
        RECT 98.620 172.040 98.760 172.490 ;
        RECT 98.100 171.720 98.360 172.040 ;
        RECT 98.560 171.720 98.820 172.040 ;
        RECT 98.160 170.875 98.300 171.720 ;
        RECT 98.090 170.505 98.370 170.875 ;
        RECT 98.160 170.000 98.300 170.505 ;
        RECT 98.100 169.680 98.360 170.000 ;
        RECT 98.560 169.340 98.820 169.660 ;
        RECT 98.100 168.660 98.360 168.980 ;
        RECT 98.160 167.960 98.300 168.660 ;
        RECT 98.100 167.640 98.360 167.960 ;
        RECT 98.620 166.795 98.760 169.340 ;
        RECT 98.550 166.425 98.830 166.795 ;
        RECT 97.640 163.560 97.900 163.880 ;
        RECT 99.080 162.520 99.220 172.740 ;
        RECT 99.540 172.380 99.680 172.740 ;
        RECT 100.850 172.545 101.130 172.915 ;
        RECT 99.480 172.060 99.740 172.380 ;
        RECT 99.940 172.290 100.200 172.380 ;
        RECT 101.380 172.290 101.520 176.740 ;
        RECT 103.150 176.625 103.430 176.995 ;
        RECT 101.770 175.945 102.050 176.315 ;
        RECT 101.780 175.800 102.040 175.945 ;
        RECT 103.220 175.520 103.360 176.625 ;
        RECT 101.840 175.440 103.360 175.520 ;
        RECT 101.780 175.380 103.360 175.440 ;
        RECT 101.780 175.120 102.040 175.380 ;
        RECT 102.240 174.780 102.500 175.100 ;
        RECT 102.700 174.780 102.960 175.100 ;
        RECT 103.160 174.780 103.420 175.100 ;
        RECT 101.780 173.080 102.040 173.400 ;
        RECT 99.940 172.235 101.520 172.290 ;
        RECT 99.940 172.150 101.590 172.235 ;
        RECT 99.940 172.060 100.200 172.150 ;
        RECT 101.310 171.865 101.590 172.150 ;
        RECT 101.840 172.040 101.980 173.080 ;
        RECT 101.780 171.720 102.040 172.040 ;
        RECT 99.480 171.555 99.740 171.700 ;
        RECT 100.400 171.610 100.660 171.700 ;
        RECT 100.000 171.555 100.660 171.610 ;
        RECT 99.470 171.185 99.750 171.555 ;
        RECT 100.000 171.470 100.670 171.555 ;
        RECT 99.480 169.340 99.740 169.660 ;
        RECT 99.540 164.900 99.680 169.340 ;
        RECT 99.480 164.580 99.740 164.900 ;
        RECT 100.000 162.860 100.140 171.470 ;
        RECT 100.390 171.185 100.670 171.470 ;
        RECT 101.310 171.185 101.590 171.555 ;
        RECT 101.380 170.000 101.520 171.185 ;
        RECT 101.320 169.910 101.580 170.000 ;
        RECT 100.460 169.770 101.580 169.910 ;
        RECT 100.460 166.940 100.600 169.770 ;
        RECT 101.320 169.680 101.580 169.770 ;
        RECT 100.860 167.640 101.120 167.960 ;
        RECT 102.300 167.870 102.440 174.780 ;
        RECT 102.760 173.060 102.900 174.780 ;
        RECT 102.700 172.740 102.960 173.060 ;
        RECT 103.220 172.235 103.360 174.780 ;
        RECT 103.150 171.865 103.430 172.235 ;
        RECT 102.700 171.380 102.960 171.700 ;
        RECT 101.840 167.730 102.440 167.870 ;
        RECT 100.400 166.620 100.660 166.940 ;
        RECT 99.940 162.540 100.200 162.860 ;
        RECT 99.020 162.200 99.280 162.520 ;
        RECT 95.790 160.305 96.070 160.675 ;
        RECT 95.860 155.210 96.000 160.305 ;
        RECT 99.080 155.660 99.680 155.800 ;
        RECT 99.080 155.210 99.220 155.660 ;
        RECT 57.150 154.710 57.430 155.210 ;
        RECT 60.370 154.710 60.650 155.210 ;
        RECT 82.910 154.710 83.190 155.210 ;
        RECT 86.130 154.710 86.410 155.210 ;
        RECT 89.350 154.710 89.630 155.210 ;
        RECT 92.570 154.710 92.850 155.210 ;
        RECT 95.790 154.710 96.070 155.210 ;
        RECT 99.010 154.710 99.290 155.210 ;
        RECT 99.540 155.120 99.680 155.660 ;
        RECT 100.920 155.120 101.060 167.640 ;
        RECT 101.840 167.280 101.980 167.730 ;
        RECT 101.780 166.960 102.040 167.280 ;
        RECT 102.230 167.105 102.510 167.475 ;
        RECT 102.240 166.960 102.500 167.105 ;
        RECT 102.760 166.940 102.900 171.380 ;
        RECT 103.150 169.825 103.430 170.195 ;
        RECT 103.160 169.680 103.420 169.825 ;
        RECT 103.620 169.680 103.880 170.000 ;
        RECT 103.680 168.980 103.820 169.680 ;
        RECT 103.620 168.660 103.880 168.980 ;
        RECT 102.700 166.620 102.960 166.940 ;
        RECT 101.780 161.180 102.040 161.500 ;
        RECT 102.240 161.180 102.500 161.500 ;
        RECT 101.840 160.480 101.980 161.180 ;
        RECT 101.780 160.160 102.040 160.480 ;
        RECT 102.300 155.210 102.440 161.180 ;
        RECT 99.540 154.980 101.060 155.120 ;
        RECT 102.230 154.710 102.510 155.210 ;
        RECT 104.140 155.120 104.280 179.540 ;
        RECT 105.000 175.460 105.260 175.780 ;
        RECT 105.060 170.340 105.200 175.460 ;
        RECT 105.000 170.020 105.260 170.340 ;
        RECT 105.060 167.280 105.200 170.020 ;
        RECT 105.000 166.960 105.260 167.280 ;
        RECT 104.540 166.620 104.800 166.940 ;
        RECT 104.600 163.880 104.740 166.620 ;
        RECT 105.060 166.170 105.200 166.960 ;
        RECT 105.520 166.940 105.660 193.140 ;
        RECT 105.920 192.120 106.180 192.440 ;
        RECT 105.980 189.720 106.120 192.120 ;
        RECT 106.900 191.080 107.040 193.140 ;
        RECT 107.820 192.440 107.960 193.910 ;
        RECT 108.220 193.480 108.480 193.800 ;
        RECT 107.760 192.120 108.020 192.440 ;
        RECT 107.300 191.440 107.560 191.760 ;
        RECT 106.840 190.760 107.100 191.080 ;
        RECT 106.380 190.420 106.640 190.740 ;
        RECT 105.920 189.400 106.180 189.720 ;
        RECT 105.980 185.640 106.120 189.400 ;
        RECT 106.440 189.380 106.580 190.420 ;
        RECT 107.360 189.630 107.500 191.440 ;
        RECT 108.280 189.800 108.420 193.480 ;
        RECT 108.740 191.420 108.880 199.260 ;
        RECT 109.200 196.520 109.340 199.260 ;
        RECT 109.660 197.200 109.800 202.320 ;
        RECT 110.120 199.580 110.260 204.700 ;
        RECT 110.580 202.835 110.720 205.720 ;
        RECT 111.960 205.360 112.100 207.850 ;
        RECT 114.200 207.760 114.460 207.850 ;
        RECT 112.360 206.740 112.620 207.060 ;
        RECT 111.900 205.040 112.160 205.360 ;
        RECT 112.420 204.760 112.560 206.740 ;
        RECT 114.190 206.545 114.470 206.915 ;
        RECT 116.490 206.545 116.770 206.915 ;
        RECT 113.280 205.720 113.540 206.040 ;
        RECT 112.820 204.875 113.080 205.020 ;
        RECT 110.980 204.360 111.240 204.680 ;
        RECT 111.960 204.620 112.560 204.760 ;
        RECT 111.040 203.320 111.180 204.360 ;
        RECT 110.980 203.000 111.240 203.320 ;
        RECT 111.960 203.080 112.100 204.620 ;
        RECT 112.810 204.505 113.090 204.875 ;
        RECT 113.340 204.250 113.480 205.720 ;
        RECT 114.260 205.020 114.400 206.545 ;
        RECT 114.660 205.040 114.920 205.360 ;
        RECT 114.200 204.700 114.460 205.020 ;
        RECT 111.500 202.940 112.100 203.080 ;
        RECT 112.420 204.110 113.480 204.250 ;
        RECT 110.510 202.465 110.790 202.835 ;
        RECT 111.500 202.550 111.640 202.940 ;
        RECT 112.420 202.640 112.560 204.110 ;
        RECT 113.740 204.020 114.000 204.340 ;
        RECT 113.800 203.080 113.940 204.020 ;
        RECT 112.820 202.660 113.080 202.980 ;
        RECT 113.340 202.940 113.940 203.080 ;
        RECT 111.040 202.410 111.640 202.550 ;
        RECT 110.060 199.260 110.320 199.580 ;
        RECT 111.040 198.640 111.180 202.410 ;
        RECT 112.360 202.320 112.620 202.640 ;
        RECT 112.420 202.040 112.560 202.320 ;
        RECT 111.500 201.900 112.560 202.040 ;
        RECT 111.500 199.580 111.640 201.900 ;
        RECT 112.360 201.300 112.620 201.620 ;
        RECT 111.900 200.115 112.160 200.260 ;
        RECT 111.890 199.745 112.170 200.115 ;
        RECT 112.420 199.920 112.560 201.300 ;
        RECT 112.360 199.600 112.620 199.920 ;
        RECT 111.440 199.260 111.700 199.580 ;
        RECT 110.120 198.500 111.180 198.640 ;
        RECT 109.600 196.880 109.860 197.200 ;
        RECT 109.140 196.200 109.400 196.520 ;
        RECT 109.200 196.035 109.340 196.200 ;
        RECT 109.130 195.665 109.410 196.035 ;
        RECT 108.680 191.100 108.940 191.420 ;
        RECT 106.900 189.490 107.500 189.630 ;
        RECT 107.820 189.660 108.420 189.800 ;
        RECT 106.380 189.060 106.640 189.380 ;
        RECT 106.380 188.380 106.640 188.700 ;
        RECT 106.440 187.195 106.580 188.380 ;
        RECT 106.900 188.020 107.040 189.490 ;
        RECT 107.290 188.185 107.570 188.555 ;
        RECT 107.360 188.020 107.500 188.185 ;
        RECT 106.840 187.700 107.100 188.020 ;
        RECT 107.300 187.700 107.560 188.020 ;
        RECT 106.370 186.825 106.650 187.195 ;
        RECT 105.920 185.320 106.180 185.640 ;
        RECT 106.900 182.920 107.040 187.700 ;
        RECT 107.290 186.145 107.570 186.515 ;
        RECT 107.360 185.980 107.500 186.145 ;
        RECT 107.300 185.660 107.560 185.980 ;
        RECT 106.840 182.600 107.100 182.920 ;
        RECT 105.920 182.260 106.180 182.580 ;
        RECT 105.460 166.620 105.720 166.940 ;
        RECT 105.980 166.600 106.120 182.260 ;
        RECT 106.380 180.560 106.640 180.880 ;
        RECT 106.440 170.340 106.580 180.560 ;
        RECT 107.360 180.540 107.500 185.660 ;
        RECT 107.300 180.220 107.560 180.540 ;
        RECT 107.820 179.860 107.960 189.660 ;
        RECT 108.220 189.060 108.480 189.380 ;
        RECT 108.280 185.980 108.420 189.060 ;
        RECT 108.680 188.610 108.940 188.700 ;
        RECT 109.660 188.610 109.800 196.880 ;
        RECT 110.120 191.760 110.260 198.500 ;
        RECT 110.970 197.705 111.250 198.075 ;
        RECT 111.040 197.540 111.180 197.705 ;
        RECT 110.980 197.220 111.240 197.540 ;
        RECT 110.520 196.540 110.780 196.860 ;
        RECT 110.060 191.440 110.320 191.760 ;
        RECT 110.060 190.760 110.320 191.080 ;
        RECT 108.680 188.470 109.800 188.610 ;
        RECT 108.680 188.380 108.940 188.470 ;
        RECT 108.220 185.660 108.480 185.980 ;
        RECT 108.280 183.940 108.420 185.660 ;
        RECT 108.220 183.620 108.480 183.940 ;
        RECT 107.760 179.540 108.020 179.860 ;
        RECT 106.840 175.120 107.100 175.440 ;
        RECT 106.900 173.595 107.040 175.120 ;
        RECT 107.300 174.100 107.560 174.420 ;
        RECT 106.830 173.225 107.110 173.595 ;
        RECT 107.360 173.400 107.500 174.100 ;
        RECT 107.300 173.080 107.560 173.400 ;
        RECT 106.840 172.740 107.100 173.060 ;
        RECT 106.380 170.020 106.640 170.340 ;
        RECT 106.900 169.660 107.040 172.740 ;
        RECT 107.820 172.040 107.960 179.540 ;
        RECT 108.680 177.500 108.940 177.820 ;
        RECT 108.220 174.100 108.480 174.420 ;
        RECT 107.300 171.720 107.560 172.040 ;
        RECT 107.760 171.720 108.020 172.040 ;
        RECT 107.360 171.440 107.500 171.720 ;
        RECT 107.360 171.300 107.960 171.440 ;
        RECT 107.290 169.825 107.570 170.195 ;
        RECT 106.840 169.340 107.100 169.660 ;
        RECT 106.840 166.620 107.100 166.940 ;
        RECT 105.920 166.280 106.180 166.600 ;
        RECT 105.460 166.170 105.720 166.260 ;
        RECT 105.060 166.030 105.720 166.170 ;
        RECT 105.460 165.940 105.720 166.030 ;
        RECT 106.900 164.755 107.040 166.620 ;
        RECT 106.830 164.385 107.110 164.755 ;
        RECT 104.540 163.560 104.800 163.880 ;
        RECT 107.360 163.395 107.500 169.825 ;
        RECT 107.290 163.025 107.570 163.395 ;
        RECT 107.820 163.200 107.960 171.300 ;
        RECT 108.280 166.115 108.420 174.100 ;
        RECT 108.740 170.000 108.880 177.500 ;
        RECT 108.680 169.680 108.940 170.000 ;
        RECT 109.200 167.960 109.340 188.470 ;
        RECT 109.600 182.260 109.860 182.580 ;
        RECT 110.120 182.435 110.260 190.760 ;
        RECT 110.580 187.195 110.720 196.540 ;
        RECT 110.980 194.160 111.240 194.480 ;
        RECT 111.040 189.040 111.180 194.160 ;
        RECT 110.980 188.720 111.240 189.040 ;
        RECT 110.510 186.825 110.790 187.195 ;
        RECT 111.500 186.660 111.640 199.260 ;
        RECT 112.360 198.920 112.620 199.240 ;
        RECT 112.420 196.860 112.560 198.920 ;
        RECT 111.890 196.345 112.170 196.715 ;
        RECT 112.360 196.540 112.620 196.860 ;
        RECT 111.440 186.340 111.700 186.660 ;
        RECT 111.440 185.660 111.700 185.980 ;
        RECT 109.660 175.440 109.800 182.260 ;
        RECT 110.050 182.065 110.330 182.435 ;
        RECT 111.500 177.820 111.640 185.660 ;
        RECT 111.960 185.300 112.100 196.345 ;
        RECT 112.420 192.100 112.560 196.540 ;
        RECT 112.880 194.820 113.020 202.660 ;
        RECT 113.340 200.600 113.480 202.940 ;
        RECT 114.720 202.550 114.860 205.040 ;
        RECT 116.040 204.700 116.300 205.020 ;
        RECT 116.100 204.340 116.240 204.700 ;
        RECT 116.560 204.680 116.700 206.545 ;
        RECT 117.420 204.700 117.680 205.020 ;
        RECT 117.880 204.700 118.140 205.020 ;
        RECT 116.500 204.360 116.760 204.680 ;
        RECT 116.040 204.020 116.300 204.340 ;
        RECT 116.040 202.660 116.300 202.980 ;
        RECT 113.800 202.410 114.860 202.550 ;
        RECT 113.280 200.280 113.540 200.600 ;
        RECT 113.800 199.580 113.940 202.410 ;
        RECT 114.200 201.640 114.460 201.960 ;
        RECT 114.260 199.920 114.400 201.640 ;
        RECT 114.660 201.300 114.920 201.620 ;
        RECT 114.720 200.795 114.860 201.300 ;
        RECT 114.650 200.425 114.930 200.795 ;
        RECT 114.720 199.920 114.860 200.425 ;
        RECT 114.200 199.600 114.460 199.920 ;
        RECT 114.660 199.600 114.920 199.920 ;
        RECT 113.740 199.260 114.000 199.580 ;
        RECT 115.580 199.260 115.840 199.580 ;
        RECT 113.280 198.920 113.540 199.240 ;
        RECT 113.340 197.200 113.480 198.920 ;
        RECT 113.280 196.880 113.540 197.200 ;
        RECT 112.820 194.500 113.080 194.820 ;
        RECT 112.360 191.780 112.620 192.100 ;
        RECT 112.880 191.840 113.020 194.500 ;
        RECT 112.880 191.700 113.480 191.840 ;
        RECT 112.820 191.100 113.080 191.420 ;
        RECT 112.360 186.000 112.620 186.320 ;
        RECT 111.900 184.980 112.160 185.300 ;
        RECT 112.420 184.280 112.560 186.000 ;
        RECT 112.360 183.960 112.620 184.280 ;
        RECT 112.880 183.260 113.020 191.100 ;
        RECT 112.820 182.940 113.080 183.260 ;
        RECT 113.340 182.920 113.480 191.700 ;
        RECT 113.800 189.720 113.940 199.260 ;
        RECT 115.110 197.705 115.390 198.075 ;
        RECT 114.650 194.985 114.930 195.355 ;
        RECT 114.190 194.305 114.470 194.675 ;
        RECT 114.260 191.080 114.400 194.305 ;
        RECT 114.200 190.760 114.460 191.080 ;
        RECT 113.740 189.400 114.000 189.720 ;
        RECT 114.200 188.720 114.460 189.040 ;
        RECT 113.740 185.660 114.000 185.980 ;
        RECT 113.280 182.600 113.540 182.920 ;
        RECT 113.800 182.320 113.940 185.660 ;
        RECT 113.340 182.180 113.940 182.320 ;
        RECT 113.340 181.220 113.480 182.180 ;
        RECT 113.740 181.240 114.000 181.560 ;
        RECT 113.280 180.900 113.540 181.220 ;
        RECT 111.440 177.500 111.700 177.820 ;
        RECT 113.280 177.390 113.540 177.480 ;
        RECT 113.800 177.390 113.940 181.240 ;
        RECT 114.260 181.220 114.400 188.720 ;
        RECT 114.200 180.900 114.460 181.220 ;
        RECT 113.280 177.250 113.940 177.390 ;
        RECT 113.280 177.160 113.540 177.250 ;
        RECT 111.440 175.460 111.700 175.780 ;
        RECT 109.600 175.120 109.860 175.440 ;
        RECT 110.980 175.120 111.240 175.440 ;
        RECT 111.040 174.955 111.180 175.120 ;
        RECT 110.970 174.585 111.250 174.955 ;
        RECT 110.060 172.400 110.320 172.720 ;
        RECT 110.120 170.680 110.260 172.400 ;
        RECT 110.520 172.060 110.780 172.380 ;
        RECT 110.060 170.360 110.320 170.680 ;
        RECT 109.140 167.640 109.400 167.960 ;
        RECT 110.580 166.940 110.720 172.060 ;
        RECT 111.500 171.700 111.640 175.460 ;
        RECT 111.900 175.120 112.160 175.440 ;
        RECT 111.960 174.760 112.100 175.120 ;
        RECT 111.900 174.440 112.160 174.760 ;
        RECT 111.440 171.380 111.700 171.700 ;
        RECT 113.800 167.960 113.940 177.250 ;
        RECT 114.200 168.660 114.460 168.980 ;
        RECT 114.260 167.960 114.400 168.660 ;
        RECT 113.740 167.640 114.000 167.960 ;
        RECT 114.200 167.640 114.460 167.960 ;
        RECT 114.720 167.620 114.860 194.985 ;
        RECT 115.180 183.260 115.320 197.705 ;
        RECT 115.640 197.540 115.780 199.260 ;
        RECT 116.100 198.075 116.240 202.660 ;
        RECT 116.960 200.280 117.220 200.600 ;
        RECT 117.020 199.580 117.160 200.280 ;
        RECT 116.500 199.260 116.760 199.580 ;
        RECT 116.960 199.260 117.220 199.580 ;
        RECT 116.030 197.705 116.310 198.075 ;
        RECT 115.580 197.220 115.840 197.540 ;
        RECT 116.040 196.880 116.300 197.200 ;
        RECT 116.100 185.300 116.240 196.880 ;
        RECT 116.560 196.860 116.700 199.260 ;
        RECT 116.500 196.540 116.760 196.860 ;
        RECT 117.480 195.355 117.620 204.700 ;
        RECT 117.940 203.320 118.080 204.700 ;
        RECT 117.880 203.000 118.140 203.320 ;
        RECT 117.870 199.745 118.150 200.115 ;
        RECT 117.410 194.985 117.690 195.355 ;
        RECT 117.940 193.800 118.080 199.745 ;
        RECT 117.880 193.480 118.140 193.800 ;
        RECT 116.500 191.100 116.760 191.420 ;
        RECT 116.040 184.980 116.300 185.300 ;
        RECT 115.120 182.940 115.380 183.260 ;
        RECT 115.580 180.220 115.840 180.540 ;
        RECT 115.640 177.820 115.780 180.220 ;
        RECT 115.580 177.500 115.840 177.820 ;
        RECT 116.100 170.340 116.240 184.980 ;
        RECT 116.560 184.280 116.700 191.100 ;
        RECT 117.880 190.760 118.140 191.080 ;
        RECT 117.940 186.400 118.080 190.760 ;
        RECT 118.400 187.195 118.540 210.140 ;
        RECT 118.860 208.760 119.000 210.740 ;
        RECT 118.800 208.440 119.060 208.760 ;
        RECT 121.560 207.760 121.820 208.080 ;
        RECT 121.620 207.060 121.760 207.760 ;
        RECT 123.000 207.060 123.140 221.250 ;
        RECT 124.770 221.070 125.050 221.570 ;
        RECT 127.990 221.070 128.270 221.570 ;
        RECT 124.840 207.740 124.980 221.070 ;
        RECT 128.060 210.370 128.200 221.070 ;
        RECT 127.600 210.230 128.200 210.370 ;
        RECT 125.700 209.460 125.960 209.780 ;
        RECT 125.760 208.080 125.900 209.460 ;
        RECT 127.600 208.760 127.740 210.230 ;
        RECT 129.380 209.800 129.640 210.120 ;
        RECT 128.450 209.265 128.730 209.635 ;
        RECT 128.520 208.760 128.660 209.265 ;
        RECT 127.540 208.440 127.800 208.760 ;
        RECT 128.000 208.440 128.260 208.760 ;
        RECT 128.460 208.440 128.720 208.760 ;
        RECT 128.060 208.080 128.200 208.440 ;
        RECT 125.700 207.760 125.960 208.080 ;
        RECT 127.080 207.760 127.340 208.080 ;
        RECT 128.000 207.760 128.260 208.080 ;
        RECT 124.780 207.420 125.040 207.740 ;
        RECT 121.560 206.740 121.820 207.060 ;
        RECT 122.940 206.740 123.200 207.060 ;
        RECT 120.630 205.185 120.910 205.555 ;
        RECT 120.700 205.020 120.840 205.185 ;
        RECT 126.620 205.040 126.880 205.360 ;
        RECT 118.790 204.505 119.070 204.875 ;
        RECT 120.640 204.700 120.900 205.020 ;
        RECT 121.560 204.700 121.820 205.020 ;
        RECT 122.940 204.700 123.200 205.020 ;
        RECT 118.860 204.340 119.000 204.505 ;
        RECT 118.800 204.020 119.060 204.340 ;
        RECT 119.260 204.020 119.520 204.340 ;
        RECT 119.320 196.180 119.460 204.020 ;
        RECT 120.180 199.940 120.440 200.260 ;
        RECT 119.720 197.560 119.980 197.880 ;
        RECT 119.260 195.860 119.520 196.180 ;
        RECT 118.800 193.820 119.060 194.140 ;
        RECT 118.330 186.825 118.610 187.195 ;
        RECT 117.940 186.260 118.540 186.400 ;
        RECT 117.880 185.320 118.140 185.640 ;
        RECT 116.500 183.960 116.760 184.280 ;
        RECT 117.420 183.280 117.680 183.600 ;
        RECT 116.500 182.600 116.760 182.920 ;
        RECT 116.560 177.820 116.700 182.600 ;
        RECT 116.960 179.540 117.220 179.860 ;
        RECT 116.500 177.500 116.760 177.820 ;
        RECT 117.020 177.480 117.160 179.540 ;
        RECT 116.960 177.160 117.220 177.480 ;
        RECT 117.480 175.635 117.620 183.280 ;
        RECT 117.940 177.820 118.080 185.320 ;
        RECT 118.400 184.280 118.540 186.260 ;
        RECT 118.340 183.960 118.600 184.280 ;
        RECT 118.330 183.425 118.610 183.795 ;
        RECT 118.400 181.755 118.540 183.425 ;
        RECT 118.860 183.260 119.000 193.820 ;
        RECT 119.260 188.040 119.520 188.360 ;
        RECT 119.320 187.875 119.460 188.040 ;
        RECT 119.250 187.505 119.530 187.875 ;
        RECT 118.800 182.940 119.060 183.260 ;
        RECT 118.800 182.260 119.060 182.580 ;
        RECT 118.330 181.385 118.610 181.755 ;
        RECT 118.860 181.220 119.000 182.260 ;
        RECT 118.800 180.900 119.060 181.220 ;
        RECT 118.340 179.540 118.600 179.860 ;
        RECT 118.400 178.840 118.540 179.540 ;
        RECT 118.340 178.520 118.600 178.840 ;
        RECT 118.800 178.180 119.060 178.500 ;
        RECT 118.860 177.820 119.000 178.180 ;
        RECT 117.880 177.500 118.140 177.820 ;
        RECT 118.340 177.675 118.600 177.820 ;
        RECT 118.330 177.305 118.610 177.675 ;
        RECT 118.800 177.500 119.060 177.820 ;
        RECT 118.340 176.995 118.600 177.140 ;
        RECT 118.330 176.625 118.610 176.995 ;
        RECT 117.410 175.265 117.690 175.635 ;
        RECT 116.500 173.080 116.760 173.400 ;
        RECT 116.040 170.020 116.300 170.340 ;
        RECT 114.660 167.300 114.920 167.620 ;
        RECT 116.560 166.940 116.700 173.080 ;
        RECT 117.880 169.000 118.140 169.320 ;
        RECT 117.940 166.940 118.080 169.000 ;
        RECT 119.320 166.940 119.460 187.505 ;
        RECT 119.780 186.660 119.920 197.560 ;
        RECT 119.720 186.340 119.980 186.660 ;
        RECT 119.720 183.960 119.980 184.280 ;
        RECT 119.780 182.580 119.920 183.960 ;
        RECT 119.720 182.260 119.980 182.580 ;
        RECT 119.720 180.560 119.980 180.880 ;
        RECT 119.780 177.820 119.920 180.560 ;
        RECT 119.720 177.500 119.980 177.820 ;
        RECT 120.240 175.440 120.380 199.940 ;
        RECT 121.100 198.580 121.360 198.900 ;
        RECT 120.640 194.840 120.900 195.160 ;
        RECT 120.700 194.140 120.840 194.840 ;
        RECT 120.640 193.820 120.900 194.140 ;
        RECT 120.700 182.580 120.840 193.820 ;
        RECT 121.160 192.440 121.300 198.580 ;
        RECT 121.620 197.540 121.760 204.700 ;
        RECT 123.000 204.340 123.140 204.700 ;
        RECT 125.240 204.360 125.500 204.680 ;
        RECT 122.940 204.020 123.200 204.340 ;
        RECT 124.780 204.020 125.040 204.340 ;
        RECT 123.000 203.080 123.140 204.020 ;
        RECT 122.540 202.940 123.140 203.080 ;
        RECT 121.560 197.220 121.820 197.540 ;
        RECT 122.540 197.200 122.680 202.940 ;
        RECT 124.840 201.620 124.980 204.020 ;
        RECT 123.400 201.300 123.660 201.620 ;
        RECT 123.860 201.300 124.120 201.620 ;
        RECT 124.780 201.300 125.040 201.620 ;
        RECT 123.460 200.795 123.600 201.300 ;
        RECT 123.390 200.425 123.670 200.795 ;
        RECT 123.400 199.940 123.660 200.260 ;
        RECT 123.460 199.580 123.600 199.940 ;
        RECT 123.400 199.260 123.660 199.580 ;
        RECT 123.400 198.580 123.660 198.900 ;
        RECT 122.480 196.880 122.740 197.200 ;
        RECT 121.560 194.840 121.820 195.160 ;
        RECT 121.100 192.120 121.360 192.440 ;
        RECT 121.620 191.760 121.760 194.840 ;
        RECT 122.540 194.480 122.680 196.880 ;
        RECT 123.460 194.820 123.600 198.580 ;
        RECT 123.920 197.880 124.060 201.300 ;
        RECT 124.320 198.920 124.580 199.240 ;
        RECT 123.860 197.560 124.120 197.880 ;
        RECT 123.400 194.500 123.660 194.820 ;
        RECT 122.480 194.160 122.740 194.480 ;
        RECT 122.020 193.480 122.280 193.800 ;
        RECT 121.560 191.440 121.820 191.760 ;
        RECT 121.560 185.320 121.820 185.640 ;
        RECT 121.620 183.940 121.760 185.320 ;
        RECT 121.560 183.620 121.820 183.940 ;
        RECT 120.640 182.260 120.900 182.580 ;
        RECT 120.640 180.900 120.900 181.220 ;
        RECT 120.700 177.820 120.840 180.900 ;
        RECT 122.080 178.500 122.220 193.480 ;
        RECT 122.940 193.140 123.200 193.460 ;
        RECT 122.480 182.940 122.740 183.260 ;
        RECT 122.540 181.220 122.680 182.940 ;
        RECT 122.480 180.900 122.740 181.220 ;
        RECT 123.000 179.860 123.140 193.140 ;
        RECT 123.850 191.585 124.130 191.955 ;
        RECT 124.380 191.790 124.520 198.920 ;
        RECT 124.780 198.580 125.040 198.900 ;
        RECT 123.920 191.080 124.060 191.585 ;
        RECT 124.320 191.470 124.580 191.790 ;
        RECT 123.860 190.760 124.120 191.080 ;
        RECT 124.380 189.800 124.520 191.470 ;
        RECT 123.460 189.720 124.520 189.800 ;
        RECT 123.400 189.660 124.520 189.720 ;
        RECT 123.400 189.400 123.660 189.660 ;
        RECT 123.860 184.980 124.120 185.300 ;
        RECT 123.920 180.880 124.060 184.980 ;
        RECT 123.400 180.560 123.660 180.880 ;
        RECT 123.860 180.560 124.120 180.880 ;
        RECT 122.480 179.540 122.740 179.860 ;
        RECT 122.940 179.540 123.200 179.860 ;
        RECT 122.540 178.500 122.680 179.540 ;
        RECT 123.460 178.840 123.600 180.560 ;
        RECT 123.400 178.520 123.660 178.840 ;
        RECT 122.020 178.180 122.280 178.500 ;
        RECT 122.480 178.180 122.740 178.500 ;
        RECT 123.920 178.160 124.060 180.560 ;
        RECT 123.860 177.840 124.120 178.160 ;
        RECT 120.640 177.500 120.900 177.820 ;
        RECT 122.480 177.675 122.740 177.820 ;
        RECT 122.470 177.305 122.750 177.675 ;
        RECT 120.180 175.120 120.440 175.440 ;
        RECT 119.720 167.300 119.980 167.620 ;
        RECT 110.060 166.620 110.320 166.940 ;
        RECT 110.520 166.620 110.780 166.940 ;
        RECT 114.200 166.620 114.460 166.940 ;
        RECT 116.500 166.620 116.760 166.940 ;
        RECT 117.880 166.620 118.140 166.940 ;
        RECT 119.260 166.620 119.520 166.940 ;
        RECT 109.600 166.280 109.860 166.600 ;
        RECT 108.210 165.745 108.490 166.115 ;
        RECT 109.660 164.220 109.800 166.280 ;
        RECT 110.120 164.900 110.260 166.620 ;
        RECT 110.060 164.580 110.320 164.900 ;
        RECT 114.260 164.220 114.400 166.620 ;
        RECT 119.780 164.900 119.920 167.300 ;
        RECT 120.240 166.600 121.300 166.680 ;
        RECT 120.180 166.540 121.360 166.600 ;
        RECT 120.180 166.280 120.440 166.540 ;
        RECT 121.100 166.280 121.360 166.540 ;
        RECT 119.720 164.580 119.980 164.900 ;
        RECT 109.600 163.900 109.860 164.220 ;
        RECT 114.200 163.900 114.460 164.220 ;
        RECT 107.760 162.880 108.020 163.200 ;
        RECT 124.840 161.500 124.980 198.580 ;
        RECT 125.300 195.160 125.440 204.360 ;
        RECT 126.680 203.320 126.820 205.040 ;
        RECT 127.140 203.320 127.280 207.760 ;
        RECT 127.990 203.825 128.270 204.195 ;
        RECT 126.620 203.000 126.880 203.320 ;
        RECT 127.080 203.000 127.340 203.320 ;
        RECT 126.160 202.660 126.420 202.980 ;
        RECT 125.700 199.940 125.960 200.260 ;
        RECT 125.760 198.900 125.900 199.940 ;
        RECT 125.700 198.580 125.960 198.900 ;
        RECT 125.760 197.880 125.900 198.580 ;
        RECT 125.700 197.560 125.960 197.880 ;
        RECT 125.700 196.880 125.960 197.200 ;
        RECT 125.760 196.715 125.900 196.880 ;
        RECT 125.690 196.345 125.970 196.715 ;
        RECT 125.690 195.665 125.970 196.035 ;
        RECT 125.240 194.840 125.500 195.160 ;
        RECT 125.760 191.760 125.900 195.665 ;
        RECT 126.220 195.160 126.360 202.660 ;
        RECT 127.540 202.320 127.800 202.640 ;
        RECT 126.620 200.280 126.880 200.600 ;
        RECT 126.680 196.180 126.820 200.280 ;
        RECT 127.600 199.920 127.740 202.320 ;
        RECT 128.060 200.600 128.200 203.825 ;
        RECT 128.920 202.660 129.180 202.980 ;
        RECT 128.000 200.280 128.260 200.600 ;
        RECT 128.450 200.425 128.730 200.795 ;
        RECT 127.540 199.600 127.800 199.920 ;
        RECT 127.600 196.860 127.740 199.600 ;
        RECT 128.000 199.435 128.260 199.580 ;
        RECT 127.990 199.065 128.270 199.435 ;
        RECT 127.990 197.705 128.270 198.075 ;
        RECT 128.060 197.200 128.200 197.705 ;
        RECT 128.520 197.540 128.660 200.425 ;
        RECT 128.460 197.220 128.720 197.540 ;
        RECT 128.000 196.880 128.260 197.200 ;
        RECT 127.540 196.540 127.800 196.860 ;
        RECT 128.460 196.540 128.720 196.860 ;
        RECT 126.620 195.860 126.880 196.180 ;
        RECT 128.520 195.355 128.660 196.540 ;
        RECT 126.160 194.840 126.420 195.160 ;
        RECT 128.450 194.985 128.730 195.355 ;
        RECT 125.700 191.440 125.960 191.760 ;
        RECT 125.700 190.420 125.960 190.740 ;
        RECT 125.230 189.545 125.510 189.915 ;
        RECT 125.300 188.700 125.440 189.545 ;
        RECT 125.240 188.380 125.500 188.700 ;
        RECT 125.240 180.395 125.500 180.540 ;
        RECT 125.230 180.025 125.510 180.395 ;
        RECT 125.760 174.955 125.900 190.420 ;
        RECT 125.690 174.585 125.970 174.955 ;
        RECT 125.690 172.545 125.970 172.915 ;
        RECT 125.240 171.380 125.500 171.700 ;
        RECT 125.300 164.220 125.440 171.380 ;
        RECT 125.760 170.000 125.900 172.545 ;
        RECT 126.220 172.380 126.360 194.840 ;
        RECT 127.990 192.945 128.270 193.315 ;
        RECT 128.460 193.140 128.720 193.460 ;
        RECT 128.060 192.100 128.200 192.945 ;
        RECT 128.000 191.780 128.260 192.100 ;
        RECT 128.520 191.760 128.660 193.140 ;
        RECT 127.080 191.440 127.340 191.760 ;
        RECT 128.460 191.440 128.720 191.760 ;
        RECT 127.140 188.555 127.280 191.440 ;
        RECT 127.540 188.610 127.800 188.700 ;
        RECT 126.620 188.040 126.880 188.360 ;
        RECT 127.070 188.185 127.350 188.555 ;
        RECT 127.540 188.470 128.200 188.610 ;
        RECT 127.540 188.380 127.800 188.470 ;
        RECT 126.680 183.940 126.820 188.040 ;
        RECT 127.540 187.700 127.800 188.020 ;
        RECT 128.060 187.875 128.200 188.470 ;
        RECT 126.620 183.620 126.880 183.940 ;
        RECT 127.600 181.220 127.740 187.700 ;
        RECT 127.990 187.505 128.270 187.875 ;
        RECT 127.540 180.900 127.800 181.220 ;
        RECT 128.520 180.880 128.660 191.440 ;
        RECT 128.460 180.560 128.720 180.880 ;
        RECT 126.620 180.220 126.880 180.540 ;
        RECT 126.680 178.500 126.820 180.220 ;
        RECT 128.980 179.035 129.120 202.660 ;
        RECT 129.440 196.860 129.580 209.800 ;
        RECT 129.840 209.460 130.100 209.780 ;
        RECT 129.900 197.880 130.040 209.460 ;
        RECT 134.440 208.100 134.700 208.420 ;
        RECT 131.220 207.760 131.480 208.080 ;
        RECT 131.280 206.040 131.420 207.760 ;
        RECT 134.500 206.040 134.640 208.100 ;
        RECT 137.660 207.760 137.920 208.080 ;
        RECT 135.820 207.080 136.080 207.400 ;
        RECT 135.880 206.040 136.020 207.080 ;
        RECT 131.220 205.720 131.480 206.040 ;
        RECT 134.440 205.720 134.700 206.040 ;
        RECT 135.820 205.720 136.080 206.040 ;
        RECT 137.720 205.700 137.860 207.760 ;
        RECT 137.660 205.380 137.920 205.700 ;
        RECT 133.060 205.040 133.320 205.360 ;
        RECT 131.220 204.700 131.480 205.020 ;
        RECT 130.760 203.000 131.020 203.320 ;
        RECT 129.840 197.560 130.100 197.880 ;
        RECT 129.840 196.880 130.100 197.200 ;
        RECT 129.380 196.540 129.640 196.860 ;
        RECT 129.380 194.500 129.640 194.820 ;
        RECT 129.440 192.100 129.580 194.500 ;
        RECT 129.900 193.995 130.040 196.880 ;
        RECT 130.290 194.985 130.570 195.355 ;
        RECT 129.830 193.625 130.110 193.995 ;
        RECT 130.360 192.100 130.500 194.985 ;
        RECT 130.820 193.315 130.960 203.000 ;
        RECT 131.280 202.300 131.420 204.700 ;
        RECT 131.680 204.020 131.940 204.340 ;
        RECT 131.220 201.980 131.480 202.300 ;
        RECT 131.220 201.300 131.480 201.620 ;
        RECT 131.280 197.200 131.420 201.300 ;
        RECT 131.740 198.900 131.880 204.020 ;
        RECT 131.680 198.580 131.940 198.900 ;
        RECT 132.140 197.560 132.400 197.880 ;
        RECT 131.220 196.880 131.480 197.200 ;
        RECT 131.280 194.140 131.420 196.880 ;
        RECT 131.220 193.820 131.480 194.140 ;
        RECT 131.280 193.460 131.420 193.820 ;
        RECT 130.750 192.945 131.030 193.315 ;
        RECT 131.220 193.140 131.480 193.460 ;
        RECT 129.380 191.780 129.640 192.100 ;
        RECT 130.300 191.780 130.560 192.100 ;
        RECT 131.280 191.760 131.420 193.140 ;
        RECT 131.220 191.440 131.480 191.760 ;
        RECT 129.380 191.330 129.640 191.420 ;
        RECT 130.300 191.330 130.560 191.420 ;
        RECT 129.380 191.190 130.560 191.330 ;
        RECT 129.380 191.100 129.640 191.190 ;
        RECT 130.300 191.100 130.560 191.190 ;
        RECT 129.440 186.660 129.580 191.100 ;
        RECT 130.750 190.905 131.030 191.275 ;
        RECT 129.380 186.340 129.640 186.660 ;
        RECT 130.820 186.320 130.960 190.905 ;
        RECT 132.200 186.320 132.340 197.560 ;
        RECT 132.600 196.880 132.860 197.200 ;
        RECT 132.660 194.480 132.800 196.880 ;
        RECT 132.600 194.160 132.860 194.480 ;
        RECT 133.120 193.995 133.260 205.040 ;
        RECT 135.360 204.875 135.620 205.020 ;
        RECT 135.350 204.505 135.630 204.875 ;
        RECT 134.900 202.320 135.160 202.640 ;
        RECT 136.280 202.320 136.540 202.640 ;
        RECT 136.740 202.320 137.000 202.640 ;
        RECT 133.520 196.880 133.780 197.200 ;
        RECT 133.050 193.625 133.330 193.995 ;
        RECT 132.600 192.120 132.860 192.440 ;
        RECT 132.660 191.955 132.800 192.120 ;
        RECT 132.590 191.585 132.870 191.955 ;
        RECT 133.120 191.760 133.260 193.625 ;
        RECT 133.580 192.100 133.720 196.880 ;
        RECT 134.440 196.540 134.700 196.860 ;
        RECT 133.520 191.780 133.780 192.100 ;
        RECT 133.060 191.440 133.320 191.760 ;
        RECT 133.970 188.185 134.250 188.555 ;
        RECT 133.520 187.700 133.780 188.020 ;
        RECT 132.590 186.825 132.870 187.195 ;
        RECT 130.760 186.000 131.020 186.320 ;
        RECT 132.140 186.000 132.400 186.320 ;
        RECT 132.660 185.980 132.800 186.825 ;
        RECT 132.600 185.660 132.860 185.980 ;
        RECT 131.740 185.155 132.340 185.210 ;
        RECT 131.670 185.070 132.340 185.155 ;
        RECT 131.670 184.785 131.950 185.070 ;
        RECT 132.200 183.260 132.340 185.070 ;
        RECT 132.140 182.940 132.400 183.260 ;
        RECT 132.600 182.940 132.860 183.260 ;
        RECT 130.760 182.600 131.020 182.920 ;
        RECT 128.910 178.665 129.190 179.035 ;
        RECT 128.980 178.500 129.120 178.665 ;
        RECT 126.620 178.180 126.880 178.500 ;
        RECT 128.920 178.180 129.180 178.500 ;
        RECT 129.380 178.180 129.640 178.500 ;
        RECT 126.160 172.060 126.420 172.380 ;
        RECT 126.620 171.720 126.880 172.040 ;
        RECT 125.700 169.680 125.960 170.000 ;
        RECT 126.680 169.515 126.820 171.720 ;
        RECT 126.610 169.145 126.890 169.515 ;
        RECT 129.440 165.435 129.580 178.180 ;
        RECT 130.300 177.500 130.560 177.820 ;
        RECT 130.360 175.440 130.500 177.500 ;
        RECT 130.300 175.120 130.560 175.440 ;
        RECT 130.360 174.275 130.500 175.120 ;
        RECT 130.820 174.760 130.960 182.600 ;
        RECT 132.660 181.560 132.800 182.940 ;
        RECT 133.050 182.745 133.330 183.115 ;
        RECT 132.600 181.240 132.860 181.560 ;
        RECT 132.600 180.560 132.860 180.880 ;
        RECT 132.660 176.120 132.800 180.560 ;
        RECT 133.120 177.820 133.260 182.745 ;
        RECT 133.580 181.560 133.720 187.700 ;
        RECT 134.040 187.000 134.180 188.185 ;
        RECT 133.980 186.680 134.240 187.000 ;
        RECT 134.500 182.435 134.640 196.540 ;
        RECT 134.960 196.180 135.100 202.320 ;
        RECT 135.820 199.600 136.080 199.920 ;
        RECT 135.360 198.920 135.620 199.240 ;
        RECT 134.900 195.860 135.160 196.180 ;
        RECT 134.430 182.065 134.710 182.435 ;
        RECT 133.520 181.240 133.780 181.560 ;
        RECT 133.980 180.560 134.240 180.880 ;
        RECT 133.060 177.500 133.320 177.820 ;
        RECT 132.600 175.800 132.860 176.120 ;
        RECT 133.120 175.350 133.260 177.500 ;
        RECT 133.520 176.995 133.780 177.140 ;
        RECT 133.510 176.625 133.790 176.995 ;
        RECT 133.520 175.350 133.780 175.440 ;
        RECT 133.120 175.210 133.780 175.350 ;
        RECT 133.520 175.120 133.780 175.210 ;
        RECT 130.760 174.440 131.020 174.760 ;
        RECT 130.290 173.905 130.570 174.275 ;
        RECT 130.360 167.280 130.500 173.905 ;
        RECT 130.820 170.340 130.960 174.440 ;
        RECT 132.600 172.060 132.860 172.380 ;
        RECT 131.220 171.720 131.480 172.040 ;
        RECT 130.760 170.020 131.020 170.340 ;
        RECT 130.300 166.960 130.560 167.280 ;
        RECT 131.280 166.940 131.420 171.720 ;
        RECT 132.660 167.280 132.800 172.060 ;
        RECT 134.040 170.680 134.180 180.560 ;
        RECT 134.500 173.400 134.640 182.065 ;
        RECT 134.890 180.705 135.170 181.075 ;
        RECT 134.960 180.200 135.100 180.705 ;
        RECT 134.900 179.880 135.160 180.200 ;
        RECT 134.960 174.420 135.100 179.880 ;
        RECT 134.900 174.100 135.160 174.420 ;
        RECT 134.440 173.080 134.700 173.400 ;
        RECT 133.980 170.360 134.240 170.680 ;
        RECT 133.060 169.340 133.320 169.660 ;
        RECT 133.120 167.960 133.260 169.340 ;
        RECT 133.060 167.640 133.320 167.960 ;
        RECT 135.420 167.280 135.560 198.920 ;
        RECT 135.880 198.900 136.020 199.600 ;
        RECT 136.340 199.435 136.480 202.320 ;
        RECT 136.800 201.475 136.940 202.320 ;
        RECT 136.730 201.105 137.010 201.475 ;
        RECT 138.120 201.300 138.380 201.620 ;
        RECT 136.270 199.065 136.550 199.435 ;
        RECT 137.660 199.260 137.920 199.580 ;
        RECT 135.820 198.580 136.080 198.900 ;
        RECT 137.720 198.755 137.860 199.260 ;
        RECT 135.880 197.395 136.020 198.580 ;
        RECT 137.650 198.385 137.930 198.755 ;
        RECT 135.810 197.025 136.090 197.395 ;
        RECT 137.200 197.220 137.460 197.540 ;
        RECT 135.820 195.860 136.080 196.180 ;
        RECT 135.880 191.080 136.020 195.860 ;
        RECT 136.280 193.480 136.540 193.800 ;
        RECT 136.340 191.760 136.480 193.480 ;
        RECT 137.260 192.440 137.400 197.220 ;
        RECT 137.650 195.665 137.930 196.035 ;
        RECT 137.720 195.160 137.860 195.665 ;
        RECT 137.660 194.840 137.920 195.160 ;
        RECT 137.200 192.120 137.460 192.440 ;
        RECT 136.280 191.440 136.540 191.760 ;
        RECT 136.740 191.100 137.000 191.420 ;
        RECT 135.820 190.760 136.080 191.080 ;
        RECT 136.270 190.225 136.550 190.595 ;
        RECT 136.340 180.880 136.480 190.225 ;
        RECT 136.800 187.000 136.940 191.100 ;
        RECT 137.660 190.760 137.920 191.080 ;
        RECT 137.720 188.700 137.860 190.760 ;
        RECT 137.660 188.380 137.920 188.700 ;
        RECT 136.740 186.680 137.000 187.000 ;
        RECT 136.740 185.660 137.000 185.980 ;
        RECT 136.280 180.560 136.540 180.880 ;
        RECT 135.820 179.880 136.080 180.200 ;
        RECT 135.880 178.500 136.020 179.880 ;
        RECT 136.800 178.840 136.940 185.660 ;
        RECT 137.660 179.540 137.920 179.860 ;
        RECT 136.740 178.520 137.000 178.840 ;
        RECT 135.820 178.180 136.080 178.500 ;
        RECT 136.730 177.985 137.010 178.355 ;
        RECT 136.740 177.840 137.000 177.985 ;
        RECT 136.280 176.820 136.540 177.140 ;
        RECT 135.810 175.945 136.090 176.315 ;
        RECT 135.880 175.780 136.020 175.945 ;
        RECT 135.820 175.460 136.080 175.780 ;
        RECT 135.880 170.680 136.020 175.460 ;
        RECT 136.340 175.440 136.480 176.820 ;
        RECT 136.800 176.120 136.940 177.840 ;
        RECT 137.200 177.500 137.460 177.820 ;
        RECT 136.740 175.800 137.000 176.120 ;
        RECT 136.280 175.120 136.540 175.440 ;
        RECT 136.280 174.440 136.540 174.760 ;
        RECT 135.820 170.360 136.080 170.680 ;
        RECT 136.340 170.195 136.480 174.440 ;
        RECT 137.260 170.680 137.400 177.500 ;
        RECT 137.720 175.100 137.860 179.540 ;
        RECT 137.660 174.780 137.920 175.100 ;
        RECT 137.200 170.360 137.460 170.680 ;
        RECT 136.270 169.825 136.550 170.195 ;
        RECT 136.340 169.660 136.480 169.825 ;
        RECT 136.280 169.340 136.540 169.660 ;
        RECT 138.180 168.580 138.320 201.300 ;
        RECT 137.720 168.440 138.320 168.580 ;
        RECT 132.600 166.960 132.860 167.280 ;
        RECT 135.360 166.960 135.620 167.280 ;
        RECT 129.840 166.620 130.100 166.940 ;
        RECT 131.220 166.620 131.480 166.940 ;
        RECT 129.370 165.065 129.650 165.435 ;
        RECT 125.240 163.900 125.500 164.220 ;
        RECT 129.900 164.075 130.040 166.620 ;
        RECT 132.130 165.065 132.410 165.435 ;
        RECT 129.830 163.705 130.110 164.075 ;
        RECT 132.200 161.500 132.340 165.065 ;
        RECT 132.660 164.220 132.800 166.960 ;
        RECT 134.900 166.620 135.160 166.940 ;
        RECT 136.740 166.620 137.000 166.940 ;
        RECT 133.060 165.940 133.320 166.260 ;
        RECT 132.600 163.900 132.860 164.220 ;
        RECT 133.120 162.860 133.260 165.940 ;
        RECT 134.960 163.200 135.100 166.620 ;
        RECT 136.800 164.900 136.940 166.620 ;
        RECT 136.740 164.580 137.000 164.900 ;
        RECT 134.900 162.880 135.160 163.200 ;
        RECT 133.060 162.540 133.320 162.860 ;
        RECT 124.780 161.180 125.040 161.500 ;
        RECT 132.140 161.180 132.400 161.500 ;
        RECT 115.120 160.840 115.380 161.160 ;
        RECT 108.680 160.500 108.940 160.820 ;
        RECT 105.060 155.660 105.660 155.800 ;
        RECT 105.060 155.120 105.200 155.660 ;
        RECT 105.520 155.210 105.660 155.660 ;
        RECT 108.740 155.210 108.880 160.500 ;
        RECT 111.900 158.460 112.160 158.780 ;
        RECT 111.960 155.210 112.100 158.460 ;
        RECT 115.180 155.210 115.320 160.840 ;
        RECT 128.000 158.120 128.260 158.440 ;
        RECT 118.340 157.440 118.600 157.760 ;
        RECT 118.400 155.210 118.540 157.440 ;
        RECT 124.780 155.400 125.040 155.720 ;
        RECT 121.560 155.210 121.820 155.380 ;
        RECT 124.840 155.210 124.980 155.400 ;
        RECT 128.060 155.210 128.200 158.120 ;
        RECT 131.220 157.780 131.480 158.100 ;
        RECT 131.280 155.210 131.420 157.780 ;
        RECT 134.430 155.545 134.710 155.915 ;
        RECT 134.500 155.210 134.640 155.545 ;
        RECT 137.720 155.210 137.860 168.440 ;
        RECT 144.100 157.100 144.360 157.420 ;
        RECT 140.880 155.740 141.140 156.060 ;
        RECT 140.940 155.210 141.080 155.740 ;
        RECT 144.160 155.210 144.300 157.100 ;
        RECT 104.140 154.980 105.200 155.120 ;
        RECT 105.450 154.710 105.730 155.210 ;
        RECT 108.670 154.710 108.950 155.210 ;
        RECT 111.890 154.710 112.170 155.210 ;
        RECT 115.110 154.710 115.390 155.210 ;
        RECT 118.330 154.710 118.610 155.210 ;
        RECT 121.550 154.710 121.830 155.210 ;
        RECT 124.770 154.710 125.050 155.210 ;
        RECT 127.990 154.710 128.270 155.210 ;
        RECT 131.210 154.710 131.490 155.210 ;
        RECT 134.430 154.710 134.710 155.210 ;
        RECT 137.650 154.710 137.930 155.210 ;
        RECT 140.870 154.710 141.150 155.210 ;
        RECT 144.090 154.710 144.370 155.210 ;
      LAYER met3 ;
        RECT 87.025 219.800 87.355 219.815 ;
        RECT 144.930 219.800 145.430 219.950 ;
        RECT 87.025 219.500 145.430 219.800 ;
        RECT 87.025 219.485 87.355 219.500 ;
        RECT 144.930 219.350 145.430 219.500 ;
        RECT 90.705 216.400 91.035 216.415 ;
        RECT 144.930 216.400 145.430 216.550 ;
        RECT 90.705 216.100 145.430 216.400 ;
        RECT 90.705 216.085 91.035 216.100 ;
        RECT 144.930 215.950 145.430 216.100 ;
        RECT 88.865 213.000 89.195 213.015 ;
        RECT 144.930 213.000 145.430 213.150 ;
        RECT 88.865 212.700 145.430 213.000 ;
        RECT 88.865 212.685 89.195 212.700 ;
        RECT 144.930 212.550 145.430 212.700 ;
        RECT 21.640 209.600 22.140 209.750 ;
        RECT 27.225 209.600 27.555 209.615 ;
        RECT 21.640 209.300 27.555 209.600 ;
        RECT 21.640 209.150 22.140 209.300 ;
        RECT 27.225 209.285 27.555 209.300 ;
        RECT 108.645 209.600 108.975 209.615 ;
        RECT 128.425 209.600 128.755 209.615 ;
        RECT 144.930 209.600 145.430 209.750 ;
        RECT 108.645 209.300 128.755 209.600 ;
        RECT 108.645 209.285 108.975 209.300 ;
        RECT 128.425 209.285 128.755 209.300 ;
        RECT 131.890 209.300 145.430 209.600 ;
        RECT 45.990 208.945 47.570 209.275 ;
        RECT 89.325 208.240 89.655 208.255 ;
        RECT 131.890 208.240 132.190 209.300 ;
        RECT 144.930 209.150 145.430 209.300 ;
        RECT 89.325 207.940 132.190 208.240 ;
        RECT 89.325 207.925 89.655 207.940 ;
        RECT 102.205 206.880 102.535 206.895 ;
        RECT 109.105 206.880 109.435 206.895 ;
        RECT 114.165 206.880 114.495 206.895 ;
        RECT 116.465 206.880 116.795 206.895 ;
        RECT 102.205 206.580 116.795 206.880 ;
        RECT 102.205 206.565 102.535 206.580 ;
        RECT 109.105 206.565 109.435 206.580 ;
        RECT 114.165 206.565 114.495 206.580 ;
        RECT 116.465 206.565 116.795 206.580 ;
        RECT 21.640 206.200 22.140 206.350 ;
        RECT 42.690 206.225 44.270 206.555 ;
        RECT 25.385 206.200 25.715 206.215 ;
        RECT 21.640 205.900 25.715 206.200 ;
        RECT 21.640 205.750 22.140 205.900 ;
        RECT 25.385 205.885 25.715 205.900 ;
        RECT 94.845 206.200 95.175 206.215 ;
        RECT 144.930 206.200 145.430 206.350 ;
        RECT 94.845 205.900 145.430 206.200 ;
        RECT 94.845 205.885 95.175 205.900 ;
        RECT 144.930 205.750 145.430 205.900 ;
        RECT 70.925 205.520 71.255 205.535 ;
        RECT 120.605 205.520 120.935 205.535 ;
        RECT 70.925 205.220 120.935 205.520 ;
        RECT 70.925 205.205 71.255 205.220 ;
        RECT 120.605 205.205 120.935 205.220 ;
        RECT 69.085 204.840 69.415 204.855 ;
        RECT 112.785 204.840 113.115 204.855 ;
        RECT 69.085 204.540 113.115 204.840 ;
        RECT 69.085 204.525 69.415 204.540 ;
        RECT 112.785 204.525 113.115 204.540 ;
        RECT 118.765 204.840 119.095 204.855 ;
        RECT 135.325 204.840 135.655 204.855 ;
        RECT 118.765 204.540 135.655 204.840 ;
        RECT 118.765 204.525 119.095 204.540 ;
        RECT 135.325 204.525 135.655 204.540 ;
        RECT 72.765 204.160 73.095 204.175 ;
        RECT 127.965 204.160 128.295 204.175 ;
        RECT 72.765 203.860 128.295 204.160 ;
        RECT 72.765 203.845 73.095 203.860 ;
        RECT 127.965 203.845 128.295 203.860 ;
        RECT 45.990 203.505 47.570 203.835 ;
        RECT 87.945 203.480 88.275 203.495 ;
        RECT 87.945 203.180 132.190 203.480 ;
        RECT 87.945 203.165 88.275 203.180 ;
        RECT 21.640 202.800 22.140 202.950 ;
        RECT 25.385 202.800 25.715 202.815 ;
        RECT 21.640 202.500 25.715 202.800 ;
        RECT 21.640 202.350 22.140 202.500 ;
        RECT 25.385 202.485 25.715 202.500 ;
        RECT 75.525 202.800 75.855 202.815 ;
        RECT 93.670 202.800 94.050 202.810 ;
        RECT 75.525 202.500 94.050 202.800 ;
        RECT 75.525 202.485 75.855 202.500 ;
        RECT 93.670 202.490 94.050 202.500 ;
        RECT 94.845 202.800 95.175 202.815 ;
        RECT 97.145 202.800 97.475 202.815 ;
        RECT 94.845 202.500 97.475 202.800 ;
        RECT 94.845 202.485 95.175 202.500 ;
        RECT 97.145 202.485 97.475 202.500 ;
        RECT 104.965 202.800 105.295 202.815 ;
        RECT 110.485 202.800 110.815 202.815 ;
        RECT 104.965 202.500 110.815 202.800 ;
        RECT 131.890 202.800 132.190 203.180 ;
        RECT 144.930 202.800 145.430 202.950 ;
        RECT 131.890 202.500 145.430 202.800 ;
        RECT 104.965 202.485 105.295 202.500 ;
        RECT 110.485 202.485 110.815 202.500 ;
        RECT 144.930 202.350 145.430 202.500 ;
        RECT 64.485 202.120 64.815 202.135 ;
        RECT 106.805 202.120 107.135 202.135 ;
        RECT 64.485 201.820 107.135 202.120 ;
        RECT 64.485 201.805 64.815 201.820 ;
        RECT 106.805 201.805 107.135 201.820 ;
        RECT 71.590 201.440 71.970 201.450 ;
        RECT 136.705 201.440 137.035 201.455 ;
        RECT 71.590 201.140 137.035 201.440 ;
        RECT 71.590 201.130 71.970 201.140 ;
        RECT 136.705 201.125 137.035 201.140 ;
        RECT 42.690 200.785 44.270 201.115 ;
        RECT 80.125 200.760 80.455 200.775 ;
        RECT 114.625 200.760 114.955 200.775 ;
        RECT 80.125 200.460 114.955 200.760 ;
        RECT 80.125 200.445 80.455 200.460 ;
        RECT 114.625 200.445 114.955 200.460 ;
        RECT 123.365 200.760 123.695 200.775 ;
        RECT 128.425 200.760 128.755 200.775 ;
        RECT 123.365 200.460 128.755 200.760 ;
        RECT 123.365 200.445 123.695 200.460 ;
        RECT 128.425 200.445 128.755 200.460 ;
        RECT 70.465 200.080 70.795 200.095 ;
        RECT 93.465 200.080 93.795 200.095 ;
        RECT 70.465 199.780 93.795 200.080 ;
        RECT 70.465 199.765 70.795 199.780 ;
        RECT 93.465 199.765 93.795 199.780 ;
        RECT 94.385 200.080 94.715 200.095 ;
        RECT 95.305 200.080 95.635 200.095 ;
        RECT 99.445 200.080 99.775 200.095 ;
        RECT 106.345 200.080 106.675 200.095 ;
        RECT 94.385 199.780 106.675 200.080 ;
        RECT 94.385 199.765 94.715 199.780 ;
        RECT 95.305 199.765 95.635 199.780 ;
        RECT 99.445 199.765 99.775 199.780 ;
        RECT 106.345 199.765 106.675 199.780 ;
        RECT 111.865 200.080 112.195 200.095 ;
        RECT 117.845 200.080 118.175 200.095 ;
        RECT 111.865 199.780 118.175 200.080 ;
        RECT 111.865 199.765 112.195 199.780 ;
        RECT 117.845 199.765 118.175 199.780 ;
        RECT 68.625 199.410 68.955 199.415 ;
        RECT 68.625 199.400 69.210 199.410 ;
        RECT 68.400 199.100 69.210 199.400 ;
        RECT 68.625 199.090 69.210 199.100 ;
        RECT 85.645 199.400 85.975 199.415 ;
        RECT 88.865 199.400 89.195 199.415 ;
        RECT 95.765 199.400 96.095 199.415 ;
        RECT 85.645 199.100 96.095 199.400 ;
        RECT 68.625 199.085 68.955 199.090 ;
        RECT 85.645 199.085 85.975 199.100 ;
        RECT 88.865 199.085 89.195 199.100 ;
        RECT 95.765 199.085 96.095 199.100 ;
        RECT 96.430 199.400 96.810 199.410 ;
        RECT 127.965 199.400 128.295 199.415 ;
        RECT 96.430 199.100 128.295 199.400 ;
        RECT 96.430 199.090 96.810 199.100 ;
        RECT 127.965 199.085 128.295 199.100 ;
        RECT 136.245 199.400 136.575 199.415 ;
        RECT 144.930 199.400 145.430 199.550 ;
        RECT 136.245 199.100 145.430 199.400 ;
        RECT 136.245 199.085 136.575 199.100 ;
        RECT 144.930 198.950 145.430 199.100 ;
        RECT 87.230 198.720 87.610 198.730 ;
        RECT 137.625 198.720 137.955 198.735 ;
        RECT 87.230 198.420 137.955 198.720 ;
        RECT 87.230 198.410 87.610 198.420 ;
        RECT 137.625 198.405 137.955 198.420 ;
        RECT 45.990 198.065 47.570 198.395 ;
        RECT 94.845 198.040 95.175 198.055 ;
        RECT 101.745 198.040 102.075 198.055 ;
        RECT 94.845 197.740 102.075 198.040 ;
        RECT 94.845 197.725 95.175 197.740 ;
        RECT 101.745 197.725 102.075 197.740 ;
        RECT 110.945 198.040 111.275 198.055 ;
        RECT 115.085 198.040 115.415 198.055 ;
        RECT 110.945 197.740 115.415 198.040 ;
        RECT 110.945 197.725 111.275 197.740 ;
        RECT 115.085 197.725 115.415 197.740 ;
        RECT 116.005 198.040 116.335 198.055 ;
        RECT 127.965 198.040 128.295 198.055 ;
        RECT 116.005 197.740 128.295 198.040 ;
        RECT 116.005 197.725 116.335 197.740 ;
        RECT 127.965 197.725 128.295 197.740 ;
        RECT 64.025 197.360 64.355 197.375 ;
        RECT 69.545 197.360 69.875 197.375 ;
        RECT 135.785 197.360 136.115 197.375 ;
        RECT 64.025 197.060 69.875 197.360 ;
        RECT 64.025 197.045 64.355 197.060 ;
        RECT 69.545 197.045 69.875 197.060 ;
        RECT 98.310 197.060 136.115 197.360 ;
        RECT 47.925 196.680 48.255 196.695 ;
        RECT 60.345 196.680 60.675 196.695 ;
        RECT 71.385 196.680 71.715 196.695 ;
        RECT 47.925 196.380 71.715 196.680 ;
        RECT 47.925 196.365 48.255 196.380 ;
        RECT 60.345 196.365 60.675 196.380 ;
        RECT 71.385 196.365 71.715 196.380 ;
        RECT 83.550 196.680 83.930 196.690 ;
        RECT 86.565 196.680 86.895 196.695 ;
        RECT 83.550 196.380 86.895 196.680 ;
        RECT 83.550 196.370 83.930 196.380 ;
        RECT 86.565 196.365 86.895 196.380 ;
        RECT 91.165 196.680 91.495 196.695 ;
        RECT 97.605 196.680 97.935 196.695 ;
        RECT 91.165 196.380 97.935 196.680 ;
        RECT 91.165 196.365 91.495 196.380 ;
        RECT 97.605 196.365 97.935 196.380 ;
        RECT 71.385 196.000 71.715 196.015 ;
        RECT 75.525 196.000 75.855 196.015 ;
        RECT 85.185 196.000 85.515 196.015 ;
        RECT 71.385 195.700 85.515 196.000 ;
        RECT 71.385 195.685 71.715 195.700 ;
        RECT 75.525 195.685 75.855 195.700 ;
        RECT 85.185 195.685 85.515 195.700 ;
        RECT 89.990 196.000 90.370 196.010 ;
        RECT 98.310 196.000 98.610 197.060 ;
        RECT 135.785 197.045 136.115 197.060 ;
        RECT 99.190 196.680 99.570 196.690 ;
        RECT 99.905 196.680 100.235 196.695 ;
        RECT 99.190 196.380 100.235 196.680 ;
        RECT 99.190 196.370 99.570 196.380 ;
        RECT 99.905 196.365 100.235 196.380 ;
        RECT 111.865 196.680 112.195 196.695 ;
        RECT 125.665 196.680 125.995 196.695 ;
        RECT 111.865 196.380 125.995 196.680 ;
        RECT 111.865 196.365 112.195 196.380 ;
        RECT 125.665 196.365 125.995 196.380 ;
        RECT 89.990 195.700 98.610 196.000 ;
        RECT 99.445 196.000 99.775 196.015 ;
        RECT 101.950 196.000 102.330 196.010 ;
        RECT 99.445 195.700 102.330 196.000 ;
        RECT 89.990 195.690 90.370 195.700 ;
        RECT 99.445 195.685 99.775 195.700 ;
        RECT 101.950 195.690 102.330 195.700 ;
        RECT 109.105 196.000 109.435 196.015 ;
        RECT 125.665 196.000 125.995 196.015 ;
        RECT 109.105 195.700 125.995 196.000 ;
        RECT 109.105 195.685 109.435 195.700 ;
        RECT 125.665 195.685 125.995 195.700 ;
        RECT 137.625 196.000 137.955 196.015 ;
        RECT 144.930 196.000 145.430 196.150 ;
        RECT 137.625 195.700 145.430 196.000 ;
        RECT 137.625 195.685 137.955 195.700 ;
        RECT 42.690 195.345 44.270 195.675 ;
        RECT 144.930 195.550 145.430 195.700 ;
        RECT 87.945 195.320 88.275 195.335 ;
        RECT 69.790 195.020 88.275 195.320 ;
        RECT 62.645 194.640 62.975 194.655 ;
        RECT 69.790 194.640 70.090 195.020 ;
        RECT 87.945 195.005 88.275 195.020 ;
        RECT 95.510 195.320 95.890 195.330 ;
        RECT 96.225 195.320 96.555 195.335 ;
        RECT 95.510 195.020 96.555 195.320 ;
        RECT 95.510 195.010 95.890 195.020 ;
        RECT 96.225 195.005 96.555 195.020 ;
        RECT 97.350 195.320 97.730 195.330 ;
        RECT 99.905 195.320 100.235 195.335 ;
        RECT 97.350 195.020 100.235 195.320 ;
        RECT 97.350 195.010 97.730 195.020 ;
        RECT 99.905 195.005 100.235 195.020 ;
        RECT 114.625 195.320 114.955 195.335 ;
        RECT 117.385 195.320 117.715 195.335 ;
        RECT 128.425 195.320 128.755 195.335 ;
        RECT 130.265 195.320 130.595 195.335 ;
        RECT 114.625 195.020 130.595 195.320 ;
        RECT 114.625 195.005 114.955 195.020 ;
        RECT 117.385 195.005 117.715 195.020 ;
        RECT 128.425 195.005 128.755 195.020 ;
        RECT 130.265 195.005 130.595 195.020 ;
        RECT 62.645 194.340 70.090 194.640 ;
        RECT 62.645 194.325 62.975 194.340 ;
        RECT 73.225 194.325 73.555 194.655 ;
        RECT 84.725 194.640 85.055 194.655 ;
        RECT 91.625 194.640 91.955 194.655 ;
        RECT 84.725 194.340 91.955 194.640 ;
        RECT 84.725 194.325 85.055 194.340 ;
        RECT 91.625 194.325 91.955 194.340 ;
        RECT 92.545 194.640 92.875 194.655 ;
        RECT 114.165 194.640 114.495 194.655 ;
        RECT 92.545 194.340 114.495 194.640 ;
        RECT 92.545 194.325 92.875 194.340 ;
        RECT 114.165 194.325 114.495 194.340 ;
        RECT 68.625 193.960 68.955 193.975 ;
        RECT 73.240 193.960 73.540 194.325 ;
        RECT 68.625 193.660 73.540 193.960 ;
        RECT 74.145 193.960 74.475 193.975 ;
        RECT 129.805 193.960 130.135 193.975 ;
        RECT 133.025 193.960 133.355 193.975 ;
        RECT 74.145 193.660 133.355 193.960 ;
        RECT 68.625 193.645 68.955 193.660 ;
        RECT 74.145 193.645 74.475 193.660 ;
        RECT 129.805 193.645 130.135 193.660 ;
        RECT 133.025 193.645 133.355 193.660 ;
        RECT 127.965 193.280 128.295 193.295 ;
        RECT 130.725 193.280 131.055 193.295 ;
        RECT 83.590 192.980 131.055 193.280 ;
        RECT 21.640 192.600 22.140 192.750 ;
        RECT 45.990 192.625 47.570 192.955 ;
        RECT 25.385 192.600 25.715 192.615 ;
        RECT 21.640 192.300 25.715 192.600 ;
        RECT 21.640 192.150 22.140 192.300 ;
        RECT 25.385 192.285 25.715 192.300 ;
        RECT 48.385 192.600 48.715 192.615 ;
        RECT 83.590 192.600 83.890 192.980 ;
        RECT 127.965 192.965 128.295 192.980 ;
        RECT 130.725 192.965 131.055 192.980 ;
        RECT 94.845 192.600 95.175 192.615 ;
        RECT 48.385 192.300 83.890 192.600 ;
        RECT 91.180 192.300 95.175 192.600 ;
        RECT 48.385 192.285 48.715 192.300 ;
        RECT 49.765 191.920 50.095 191.935 ;
        RECT 67.705 191.920 68.035 191.935 ;
        RECT 49.765 191.620 68.035 191.920 ;
        RECT 49.765 191.605 50.095 191.620 ;
        RECT 67.705 191.605 68.035 191.620 ;
        RECT 81.045 191.920 81.375 191.935 ;
        RECT 91.180 191.920 91.480 192.300 ;
        RECT 94.845 192.285 95.175 192.300 ;
        RECT 97.605 192.600 97.935 192.615 ;
        RECT 144.930 192.600 145.430 192.750 ;
        RECT 97.605 192.300 145.430 192.600 ;
        RECT 97.605 192.285 97.935 192.300 ;
        RECT 144.930 192.150 145.430 192.300 ;
        RECT 81.045 191.620 91.480 191.920 ;
        RECT 92.085 191.920 92.415 191.935 ;
        RECT 98.270 191.920 98.650 191.930 ;
        RECT 92.085 191.620 98.650 191.920 ;
        RECT 81.045 191.605 81.375 191.620 ;
        RECT 92.085 191.605 92.415 191.620 ;
        RECT 98.270 191.610 98.650 191.620 ;
        RECT 123.825 191.920 124.155 191.935 ;
        RECT 132.565 191.920 132.895 191.935 ;
        RECT 123.825 191.620 132.895 191.920 ;
        RECT 123.825 191.605 124.155 191.620 ;
        RECT 132.565 191.605 132.895 191.620 ;
        RECT 29.985 191.240 30.315 191.255 ;
        RECT 59.885 191.240 60.215 191.255 ;
        RECT 29.985 190.940 60.215 191.240 ;
        RECT 29.985 190.925 30.315 190.940 ;
        RECT 59.885 190.925 60.215 190.940 ;
        RECT 68.830 191.240 69.210 191.250 ;
        RECT 69.545 191.240 69.875 191.255 ;
        RECT 68.830 190.940 69.875 191.240 ;
        RECT 68.830 190.930 69.210 190.940 ;
        RECT 69.545 190.925 69.875 190.940 ;
        RECT 83.345 191.240 83.675 191.255 ;
        RECT 130.725 191.240 131.055 191.255 ;
        RECT 83.345 190.940 131.055 191.240 ;
        RECT 83.345 190.925 83.675 190.940 ;
        RECT 130.725 190.925 131.055 190.940 ;
        RECT 67.245 190.560 67.575 190.575 ;
        RECT 72.305 190.560 72.635 190.575 ;
        RECT 92.085 190.560 92.415 190.575 ;
        RECT 67.245 190.260 92.415 190.560 ;
        RECT 67.245 190.245 67.575 190.260 ;
        RECT 72.305 190.245 72.635 190.260 ;
        RECT 92.085 190.245 92.415 190.260 ;
        RECT 94.385 190.560 94.715 190.575 ;
        RECT 136.245 190.560 136.575 190.575 ;
        RECT 94.385 190.260 136.575 190.560 ;
        RECT 94.385 190.245 94.715 190.260 ;
        RECT 136.245 190.245 136.575 190.260 ;
        RECT 42.690 189.905 44.270 190.235 ;
        RECT 55.285 189.880 55.615 189.895 ;
        RECT 62.645 189.880 62.975 189.895 ;
        RECT 74.145 189.880 74.475 189.895 ;
        RECT 55.285 189.580 74.475 189.880 ;
        RECT 55.285 189.565 55.615 189.580 ;
        RECT 62.645 189.565 62.975 189.580 ;
        RECT 74.145 189.565 74.475 189.580 ;
        RECT 91.625 189.880 91.955 189.895 ;
        RECT 103.790 189.880 104.170 189.890 ;
        RECT 91.625 189.580 104.170 189.880 ;
        RECT 91.625 189.565 91.955 189.580 ;
        RECT 103.790 189.570 104.170 189.580 ;
        RECT 125.205 189.880 125.535 189.895 ;
        RECT 125.205 189.580 131.960 189.880 ;
        RECT 125.205 189.565 125.535 189.580 ;
        RECT 21.640 189.200 22.140 189.350 ;
        RECT 25.385 189.200 25.715 189.215 ;
        RECT 21.640 188.900 25.715 189.200 ;
        RECT 21.640 188.750 22.140 188.900 ;
        RECT 25.385 188.885 25.715 188.900 ;
        RECT 90.245 189.200 90.575 189.215 ;
        RECT 131.660 189.200 131.960 189.580 ;
        RECT 144.930 189.200 145.430 189.350 ;
        RECT 90.245 188.900 128.050 189.200 ;
        RECT 131.660 188.900 145.430 189.200 ;
        RECT 90.245 188.885 90.575 188.900 ;
        RECT 53.905 188.520 54.235 188.535 ;
        RECT 57.585 188.520 57.915 188.535 ;
        RECT 53.905 188.220 57.915 188.520 ;
        RECT 53.905 188.205 54.235 188.220 ;
        RECT 57.585 188.205 57.915 188.220 ;
        RECT 80.585 188.520 80.915 188.535 ;
        RECT 84.265 188.520 84.595 188.535 ;
        RECT 91.830 188.520 92.210 188.530 ;
        RECT 80.585 188.220 92.210 188.520 ;
        RECT 80.585 188.205 80.915 188.220 ;
        RECT 84.265 188.205 84.595 188.220 ;
        RECT 91.830 188.210 92.210 188.220 ;
        RECT 93.925 188.520 94.255 188.535 ;
        RECT 96.225 188.520 96.555 188.535 ;
        RECT 93.925 188.220 96.555 188.520 ;
        RECT 93.925 188.205 94.255 188.220 ;
        RECT 96.225 188.205 96.555 188.220 ;
        RECT 100.110 188.520 100.490 188.530 ;
        RECT 104.045 188.520 104.375 188.535 ;
        RECT 100.110 188.220 104.375 188.520 ;
        RECT 100.110 188.210 100.490 188.220 ;
        RECT 104.045 188.205 104.375 188.220 ;
        RECT 107.265 188.520 107.595 188.535 ;
        RECT 127.045 188.520 127.375 188.535 ;
        RECT 107.265 188.220 127.375 188.520 ;
        RECT 127.750 188.520 128.050 188.900 ;
        RECT 144.930 188.750 145.430 188.900 ;
        RECT 133.945 188.520 134.275 188.535 ;
        RECT 127.750 188.220 134.275 188.520 ;
        RECT 107.265 188.205 107.595 188.220 ;
        RECT 127.045 188.205 127.375 188.220 ;
        RECT 133.945 188.205 134.275 188.220 ;
        RECT 48.385 187.840 48.715 187.855 ;
        RECT 64.025 187.840 64.355 187.855 ;
        RECT 81.505 187.840 81.835 187.855 ;
        RECT 93.465 187.840 93.795 187.855 ;
        RECT 97.605 187.840 97.935 187.855 ;
        RECT 48.385 187.540 97.935 187.840 ;
        RECT 48.385 187.525 48.715 187.540 ;
        RECT 64.025 187.525 64.355 187.540 ;
        RECT 81.505 187.525 81.835 187.540 ;
        RECT 93.465 187.525 93.795 187.540 ;
        RECT 97.605 187.525 97.935 187.540 ;
        RECT 99.445 187.840 99.775 187.855 ;
        RECT 104.045 187.840 104.375 187.855 ;
        RECT 99.445 187.540 104.375 187.840 ;
        RECT 99.445 187.525 99.775 187.540 ;
        RECT 104.045 187.525 104.375 187.540 ;
        RECT 119.225 187.840 119.555 187.855 ;
        RECT 127.965 187.840 128.295 187.855 ;
        RECT 119.225 187.540 128.295 187.840 ;
        RECT 119.225 187.525 119.555 187.540 ;
        RECT 127.965 187.525 128.295 187.540 ;
        RECT 45.990 187.185 47.570 187.515 ;
        RECT 80.125 187.160 80.455 187.175 ;
        RECT 84.265 187.160 84.595 187.175 ;
        RECT 88.405 187.170 88.735 187.175 ;
        RECT 80.125 186.860 84.595 187.160 ;
        RECT 80.125 186.845 80.455 186.860 ;
        RECT 84.265 186.845 84.595 186.860 ;
        RECT 88.150 187.160 88.735 187.170 ;
        RECT 93.670 187.160 94.050 187.170 ;
        RECT 94.845 187.160 95.175 187.175 ;
        RECT 102.665 187.160 102.995 187.175 ;
        RECT 88.150 186.860 88.960 187.160 ;
        RECT 93.670 186.860 102.995 187.160 ;
        RECT 88.150 186.850 88.735 186.860 ;
        RECT 93.670 186.850 94.050 186.860 ;
        RECT 88.405 186.845 88.735 186.850 ;
        RECT 94.845 186.845 95.175 186.860 ;
        RECT 102.665 186.845 102.995 186.860 ;
        RECT 106.345 187.160 106.675 187.175 ;
        RECT 110.485 187.160 110.815 187.175 ;
        RECT 106.345 186.860 110.815 187.160 ;
        RECT 106.345 186.845 106.675 186.860 ;
        RECT 110.485 186.845 110.815 186.860 ;
        RECT 118.305 187.160 118.635 187.175 ;
        RECT 132.565 187.160 132.895 187.175 ;
        RECT 118.305 186.860 132.895 187.160 ;
        RECT 118.305 186.845 118.635 186.860 ;
        RECT 132.565 186.845 132.895 186.860 ;
        RECT 59.425 186.480 59.755 186.495 ;
        RECT 93.465 186.480 93.795 186.495 ;
        RECT 97.145 186.480 97.475 186.495 ;
        RECT 59.425 186.180 91.250 186.480 ;
        RECT 59.425 186.165 59.755 186.180 ;
        RECT 21.640 185.800 22.140 185.950 ;
        RECT 24.465 185.800 24.795 185.815 ;
        RECT 21.640 185.500 24.795 185.800 ;
        RECT 21.640 185.350 22.140 185.500 ;
        RECT 24.465 185.485 24.795 185.500 ;
        RECT 76.905 185.800 77.235 185.815 ;
        RECT 79.665 185.800 79.995 185.815 ;
        RECT 86.565 185.800 86.895 185.815 ;
        RECT 89.325 185.810 89.655 185.815 ;
        RECT 76.905 185.500 79.995 185.800 ;
        RECT 76.905 185.485 77.235 185.500 ;
        RECT 79.665 185.485 79.995 185.500 ;
        RECT 82.670 185.500 86.895 185.800 ;
        RECT 42.690 184.465 44.270 184.795 ;
        RECT 82.670 184.455 82.970 185.500 ;
        RECT 86.565 185.485 86.895 185.500 ;
        RECT 89.070 185.800 89.655 185.810 ;
        RECT 89.070 185.500 89.880 185.800 ;
        RECT 89.070 185.490 89.655 185.500 ;
        RECT 89.325 185.485 89.655 185.490 ;
        RECT 85.185 185.120 85.515 185.135 ;
        RECT 86.310 185.120 86.690 185.130 ;
        RECT 85.185 184.820 86.690 185.120 ;
        RECT 90.950 185.120 91.250 186.180 ;
        RECT 93.465 186.180 97.475 186.480 ;
        RECT 93.465 186.165 93.795 186.180 ;
        RECT 97.145 186.165 97.475 186.180 ;
        RECT 104.965 186.480 105.295 186.495 ;
        RECT 107.265 186.480 107.595 186.495 ;
        RECT 104.965 186.180 107.595 186.480 ;
        RECT 104.965 186.165 105.295 186.180 ;
        RECT 107.265 186.165 107.595 186.180 ;
        RECT 91.625 185.800 91.955 185.815 ;
        RECT 102.205 185.800 102.535 185.815 ;
        RECT 91.625 185.500 102.535 185.800 ;
        RECT 91.625 185.485 91.955 185.500 ;
        RECT 102.205 185.485 102.535 185.500 ;
        RECT 103.585 185.800 103.915 185.815 ;
        RECT 144.930 185.800 145.430 185.950 ;
        RECT 103.585 185.500 145.430 185.800 ;
        RECT 103.585 185.485 103.915 185.500 ;
        RECT 144.930 185.350 145.430 185.500 ;
        RECT 94.385 185.120 94.715 185.135 ;
        RECT 90.950 184.820 94.715 185.120 ;
        RECT 85.185 184.805 85.515 184.820 ;
        RECT 86.310 184.810 86.690 184.820 ;
        RECT 94.385 184.805 94.715 184.820 ;
        RECT 96.225 185.120 96.555 185.135 ;
        RECT 131.645 185.120 131.975 185.135 ;
        RECT 96.225 184.820 131.975 185.120 ;
        RECT 96.225 184.805 96.555 184.820 ;
        RECT 131.645 184.805 131.975 184.820 ;
        RECT 82.425 184.140 82.970 184.455 ;
        RECT 85.185 184.440 85.515 184.455 ;
        RECT 124.950 184.440 125.330 184.450 ;
        RECT 85.185 184.140 125.330 184.440 ;
        RECT 82.425 184.125 82.755 184.140 ;
        RECT 85.185 184.125 85.515 184.140 ;
        RECT 124.950 184.130 125.330 184.140 ;
        RECT 47.005 183.760 47.335 183.775 ;
        RECT 63.105 183.760 63.435 183.775 ;
        RECT 47.005 183.460 63.435 183.760 ;
        RECT 47.005 183.445 47.335 183.460 ;
        RECT 63.105 183.445 63.435 183.460 ;
        RECT 83.345 183.760 83.675 183.775 ;
        RECT 87.025 183.760 87.355 183.775 ;
        RECT 83.345 183.460 87.355 183.760 ;
        RECT 83.345 183.445 83.675 183.460 ;
        RECT 87.025 183.445 87.355 183.460 ;
        RECT 88.405 183.760 88.735 183.775 ;
        RECT 118.305 183.760 118.635 183.775 ;
        RECT 88.405 183.460 118.635 183.760 ;
        RECT 88.405 183.445 88.735 183.460 ;
        RECT 118.305 183.445 118.635 183.460 ;
        RECT 86.565 183.080 86.895 183.095 ;
        RECT 89.785 183.080 90.115 183.095 ;
        RECT 133.025 183.080 133.355 183.095 ;
        RECT 86.565 182.780 89.410 183.080 ;
        RECT 86.565 182.765 86.895 182.780 ;
        RECT 21.640 182.400 22.140 182.550 ;
        RECT 25.385 182.400 25.715 182.415 ;
        RECT 21.640 182.100 25.715 182.400 ;
        RECT 21.640 181.950 22.140 182.100 ;
        RECT 25.385 182.085 25.715 182.100 ;
        RECT 71.385 182.400 71.715 182.415 ;
        RECT 88.150 182.400 88.530 182.410 ;
        RECT 71.385 182.100 88.530 182.400 ;
        RECT 89.110 182.400 89.410 182.780 ;
        RECT 89.785 182.780 133.355 183.080 ;
        RECT 89.785 182.765 90.115 182.780 ;
        RECT 133.025 182.765 133.355 182.780 ;
        RECT 92.750 182.400 93.130 182.410 ;
        RECT 89.110 182.100 93.130 182.400 ;
        RECT 71.385 182.085 71.715 182.100 ;
        RECT 88.150 182.090 88.530 182.100 ;
        RECT 92.750 182.090 93.130 182.100 ;
        RECT 94.845 182.400 95.175 182.415 ;
        RECT 98.985 182.400 99.315 182.415 ;
        RECT 94.845 182.100 99.315 182.400 ;
        RECT 94.845 182.085 95.175 182.100 ;
        RECT 98.985 182.085 99.315 182.100 ;
        RECT 100.365 182.400 100.695 182.415 ;
        RECT 110.025 182.400 110.355 182.415 ;
        RECT 134.405 182.400 134.735 182.415 ;
        RECT 144.930 182.400 145.430 182.550 ;
        RECT 100.365 182.100 134.735 182.400 ;
        RECT 100.365 182.085 100.695 182.100 ;
        RECT 110.025 182.085 110.355 182.100 ;
        RECT 134.405 182.085 134.735 182.100 ;
        RECT 138.790 182.100 145.430 182.400 ;
        RECT 45.990 181.745 47.570 182.075 ;
        RECT 72.305 181.720 72.635 181.735 ;
        RECT 85.390 181.720 85.770 181.730 ;
        RECT 86.105 181.720 86.435 181.735 ;
        RECT 87.025 181.730 87.355 181.735 ;
        RECT 87.025 181.720 87.610 181.730 ;
        RECT 72.305 181.420 81.820 181.720 ;
        RECT 72.305 181.405 72.635 181.420 ;
        RECT 50.225 181.040 50.555 181.055 ;
        RECT 80.585 181.040 80.915 181.055 ;
        RECT 50.225 180.740 80.915 181.040 ;
        RECT 81.520 181.040 81.820 181.420 ;
        RECT 85.390 181.420 86.435 181.720 ;
        RECT 86.800 181.420 87.610 181.720 ;
        RECT 85.390 181.410 85.770 181.420 ;
        RECT 86.105 181.405 86.435 181.420 ;
        RECT 87.025 181.410 87.610 181.420 ;
        RECT 90.245 181.720 90.575 181.735 ;
        RECT 95.765 181.720 96.095 181.735 ;
        RECT 90.245 181.420 96.095 181.720 ;
        RECT 87.025 181.405 87.355 181.410 ;
        RECT 90.245 181.405 90.575 181.420 ;
        RECT 95.765 181.405 96.095 181.420 ;
        RECT 98.270 181.720 98.650 181.730 ;
        RECT 98.985 181.720 99.315 181.735 ;
        RECT 98.270 181.420 99.315 181.720 ;
        RECT 98.270 181.410 98.650 181.420 ;
        RECT 98.985 181.405 99.315 181.420 ;
        RECT 118.305 181.720 118.635 181.735 ;
        RECT 138.790 181.720 139.090 182.100 ;
        RECT 144.930 181.950 145.430 182.100 ;
        RECT 118.305 181.420 139.090 181.720 ;
        RECT 118.305 181.405 118.635 181.420 ;
        RECT 88.405 181.040 88.735 181.055 ;
        RECT 81.520 180.740 88.735 181.040 ;
        RECT 50.225 180.725 50.555 180.740 ;
        RECT 80.585 180.725 80.915 180.740 ;
        RECT 88.405 180.725 88.735 180.740 ;
        RECT 89.785 181.040 90.115 181.055 ;
        RECT 134.865 181.040 135.195 181.055 ;
        RECT 89.785 180.740 135.195 181.040 ;
        RECT 89.785 180.725 90.115 180.740 ;
        RECT 134.865 180.725 135.195 180.740 ;
        RECT 59.885 180.360 60.215 180.375 ;
        RECT 66.785 180.360 67.115 180.375 ;
        RECT 59.885 180.060 67.115 180.360 ;
        RECT 59.885 180.045 60.215 180.060 ;
        RECT 66.785 180.045 67.115 180.060 ;
        RECT 77.825 180.360 78.155 180.375 ;
        RECT 83.345 180.360 83.675 180.375 ;
        RECT 77.825 180.060 83.675 180.360 ;
        RECT 77.825 180.045 78.155 180.060 ;
        RECT 83.345 180.045 83.675 180.060 ;
        RECT 95.765 180.360 96.095 180.375 ;
        RECT 125.205 180.360 125.535 180.375 ;
        RECT 95.765 180.060 125.535 180.360 ;
        RECT 95.765 180.045 96.095 180.060 ;
        RECT 125.205 180.045 125.535 180.060 ;
        RECT 60.805 179.680 61.135 179.695 ;
        RECT 65.865 179.680 66.195 179.695 ;
        RECT 60.805 179.380 66.195 179.680 ;
        RECT 60.805 179.365 61.135 179.380 ;
        RECT 65.865 179.365 66.195 179.380 ;
        RECT 74.605 179.680 74.935 179.695 ;
        RECT 90.705 179.690 91.035 179.695 ;
        RECT 84.470 179.680 84.850 179.690 ;
        RECT 89.990 179.680 90.370 179.690 ;
        RECT 74.605 179.380 90.370 179.680 ;
        RECT 74.605 179.365 74.935 179.380 ;
        RECT 84.470 179.370 84.850 179.380 ;
        RECT 89.990 179.370 90.370 179.380 ;
        RECT 90.705 179.680 91.290 179.690 ;
        RECT 90.705 179.380 91.490 179.680 ;
        RECT 91.870 179.380 130.810 179.680 ;
        RECT 90.705 179.370 91.290 179.380 ;
        RECT 90.705 179.365 91.035 179.370 ;
        RECT 21.640 179.000 22.140 179.150 ;
        RECT 42.690 179.025 44.270 179.355 ;
        RECT 25.385 179.000 25.715 179.015 ;
        RECT 21.640 178.700 25.715 179.000 ;
        RECT 21.640 178.550 22.140 178.700 ;
        RECT 25.385 178.685 25.715 178.700 ;
        RECT 57.125 179.000 57.455 179.015 ;
        RECT 64.485 179.000 64.815 179.015 ;
        RECT 57.125 178.700 64.815 179.000 ;
        RECT 57.125 178.685 57.455 178.700 ;
        RECT 64.485 178.685 64.815 178.700 ;
        RECT 76.905 179.000 77.235 179.015 ;
        RECT 91.870 179.000 92.170 179.380 ;
        RECT 76.905 178.700 92.170 179.000 ;
        RECT 93.465 179.000 93.795 179.015 ;
        RECT 128.885 179.000 129.215 179.015 ;
        RECT 93.465 178.700 129.215 179.000 ;
        RECT 130.510 179.000 130.810 179.380 ;
        RECT 144.930 179.000 145.430 179.150 ;
        RECT 130.510 178.700 145.430 179.000 ;
        RECT 76.905 178.685 77.235 178.700 ;
        RECT 93.465 178.685 93.795 178.700 ;
        RECT 128.885 178.685 129.215 178.700 ;
        RECT 144.930 178.550 145.430 178.700 ;
        RECT 63.105 178.005 63.435 178.335 ;
        RECT 82.885 178.320 83.215 178.335 ;
        RECT 83.550 178.320 83.930 178.330 ;
        RECT 82.885 178.020 83.930 178.320 ;
        RECT 82.885 178.005 83.215 178.020 ;
        RECT 83.550 178.010 83.930 178.020 ;
        RECT 84.725 178.320 85.055 178.335 ;
        RECT 88.405 178.320 88.735 178.335 ;
        RECT 84.725 178.020 88.735 178.320 ;
        RECT 84.725 178.005 85.055 178.020 ;
        RECT 88.405 178.005 88.735 178.020 ;
        RECT 89.785 178.320 90.115 178.335 ;
        RECT 94.590 178.320 94.970 178.330 ;
        RECT 89.785 178.020 94.970 178.320 ;
        RECT 89.785 178.005 90.115 178.020 ;
        RECT 94.590 178.010 94.970 178.020 ;
        RECT 95.765 178.320 96.095 178.335 ;
        RECT 100.110 178.320 100.490 178.330 ;
        RECT 136.705 178.320 137.035 178.335 ;
        RECT 95.765 178.020 100.490 178.320 ;
        RECT 95.765 178.005 96.095 178.020 ;
        RECT 100.110 178.010 100.490 178.020 ;
        RECT 101.070 178.020 137.035 178.320 ;
        RECT 63.120 177.640 63.420 178.005 ;
        RECT 64.945 177.640 65.275 177.655 ;
        RECT 63.120 177.340 65.275 177.640 ;
        RECT 64.945 177.325 65.275 177.340 ;
        RECT 83.345 177.640 83.675 177.655 ;
        RECT 97.605 177.640 97.935 177.655 ;
        RECT 101.070 177.640 101.370 178.020 ;
        RECT 136.705 178.005 137.035 178.020 ;
        RECT 83.345 177.340 101.370 177.640 ;
        RECT 118.305 177.640 118.635 177.655 ;
        RECT 122.445 177.640 122.775 177.655 ;
        RECT 118.305 177.340 122.775 177.640 ;
        RECT 83.345 177.325 83.675 177.340 ;
        RECT 97.605 177.325 97.935 177.340 ;
        RECT 118.305 177.325 118.635 177.340 ;
        RECT 122.445 177.325 122.775 177.340 ;
        RECT 81.965 176.960 82.295 176.975 ;
        RECT 89.325 176.960 89.655 176.975 ;
        RECT 89.990 176.960 90.370 176.970 ;
        RECT 81.965 176.660 90.370 176.960 ;
        RECT 81.965 176.645 82.295 176.660 ;
        RECT 89.325 176.645 89.655 176.660 ;
        RECT 89.990 176.650 90.370 176.660 ;
        RECT 91.165 176.960 91.495 176.975 ;
        RECT 103.125 176.960 103.455 176.975 ;
        RECT 91.165 176.660 103.455 176.960 ;
        RECT 91.165 176.645 91.495 176.660 ;
        RECT 103.125 176.645 103.455 176.660 ;
        RECT 118.305 176.960 118.635 176.975 ;
        RECT 133.485 176.960 133.815 176.975 ;
        RECT 118.305 176.660 133.815 176.960 ;
        RECT 118.305 176.645 118.635 176.660 ;
        RECT 133.485 176.645 133.815 176.660 ;
        RECT 45.990 176.305 47.570 176.635 ;
        RECT 49.765 176.280 50.095 176.295 ;
        RECT 72.305 176.280 72.635 176.295 ;
        RECT 49.765 175.980 72.635 176.280 ;
        RECT 49.765 175.965 50.095 175.980 ;
        RECT 72.305 175.965 72.635 175.980 ;
        RECT 75.985 176.280 76.315 176.295 ;
        RECT 87.230 176.280 87.610 176.290 ;
        RECT 75.985 175.980 87.610 176.280 ;
        RECT 75.985 175.965 76.315 175.980 ;
        RECT 87.230 175.970 87.610 175.980 ;
        RECT 88.405 176.280 88.735 176.295 ;
        RECT 91.625 176.280 91.955 176.295 ;
        RECT 88.405 175.980 91.955 176.280 ;
        RECT 88.405 175.965 88.735 175.980 ;
        RECT 91.625 175.965 91.955 175.980 ;
        RECT 92.545 176.280 92.875 176.295 ;
        RECT 96.430 176.280 96.810 176.290 ;
        RECT 92.545 175.980 96.810 176.280 ;
        RECT 92.545 175.965 92.875 175.980 ;
        RECT 96.430 175.970 96.810 175.980 ;
        RECT 98.525 176.280 98.855 176.295 ;
        RECT 101.745 176.280 102.075 176.295 ;
        RECT 135.785 176.280 136.115 176.295 ;
        RECT 98.525 175.980 102.075 176.280 ;
        RECT 98.525 175.965 98.855 175.980 ;
        RECT 101.745 175.965 102.075 175.980 ;
        RECT 102.680 175.980 136.115 176.280 ;
        RECT 63.105 175.600 63.435 175.615 ;
        RECT 66.325 175.600 66.655 175.615 ;
        RECT 63.105 175.300 66.655 175.600 ;
        RECT 63.105 175.285 63.435 175.300 ;
        RECT 66.325 175.285 66.655 175.300 ;
        RECT 69.085 175.600 69.415 175.615 ;
        RECT 75.525 175.600 75.855 175.615 ;
        RECT 69.085 175.300 75.855 175.600 ;
        RECT 69.085 175.285 69.415 175.300 ;
        RECT 75.525 175.285 75.855 175.300 ;
        RECT 87.025 175.600 87.355 175.615 ;
        RECT 93.670 175.600 94.050 175.610 ;
        RECT 102.680 175.600 102.980 175.980 ;
        RECT 135.785 175.965 136.115 175.980 ;
        RECT 117.385 175.600 117.715 175.615 ;
        RECT 87.025 175.300 94.050 175.600 ;
        RECT 87.025 175.285 87.355 175.300 ;
        RECT 93.670 175.290 94.050 175.300 ;
        RECT 95.550 175.300 102.980 175.600 ;
        RECT 103.600 175.300 117.715 175.600 ;
        RECT 61.265 174.920 61.595 174.935 ;
        RECT 64.485 174.920 64.815 174.935 ;
        RECT 61.265 174.620 64.815 174.920 ;
        RECT 66.340 174.920 66.640 175.285 ;
        RECT 76.905 174.920 77.235 174.935 ;
        RECT 66.340 174.620 77.235 174.920 ;
        RECT 61.265 174.605 61.595 174.620 ;
        RECT 64.485 174.605 64.815 174.620 ;
        RECT 76.905 174.605 77.235 174.620 ;
        RECT 93.670 174.920 94.050 174.930 ;
        RECT 95.550 174.920 95.850 175.300 ;
        RECT 96.685 174.930 97.015 174.935 ;
        RECT 93.670 174.620 95.850 174.920 ;
        RECT 96.430 174.920 97.015 174.930 ;
        RECT 97.605 174.920 97.935 174.935 ;
        RECT 99.445 174.920 99.775 174.935 ;
        RECT 96.430 174.620 97.240 174.920 ;
        RECT 97.605 174.620 99.775 174.920 ;
        RECT 93.670 174.610 94.050 174.620 ;
        RECT 96.430 174.610 97.015 174.620 ;
        RECT 96.685 174.605 97.015 174.610 ;
        RECT 97.605 174.605 97.935 174.620 ;
        RECT 99.445 174.605 99.775 174.620 ;
        RECT 100.365 174.920 100.695 174.935 ;
        RECT 103.600 174.920 103.900 175.300 ;
        RECT 117.385 175.285 117.715 175.300 ;
        RECT 124.950 175.600 125.330 175.610 ;
        RECT 144.930 175.600 145.430 175.750 ;
        RECT 124.950 175.300 145.430 175.600 ;
        RECT 124.950 175.290 125.330 175.300 ;
        RECT 144.930 175.150 145.430 175.300 ;
        RECT 100.365 174.620 103.900 174.920 ;
        RECT 110.945 174.920 111.275 174.935 ;
        RECT 125.665 174.920 125.995 174.935 ;
        RECT 110.945 174.620 125.995 174.920 ;
        RECT 100.365 174.605 100.695 174.620 ;
        RECT 110.945 174.605 111.275 174.620 ;
        RECT 125.665 174.605 125.995 174.620 ;
        RECT 48.385 174.240 48.715 174.255 ;
        RECT 81.045 174.240 81.375 174.255 ;
        RECT 92.085 174.240 92.415 174.255 ;
        RECT 48.385 173.940 92.415 174.240 ;
        RECT 48.385 173.925 48.715 173.940 ;
        RECT 81.045 173.925 81.375 173.940 ;
        RECT 92.085 173.925 92.415 173.940 ;
        RECT 92.750 174.240 93.130 174.250 ;
        RECT 130.265 174.240 130.595 174.255 ;
        RECT 92.750 173.940 130.595 174.240 ;
        RECT 92.750 173.930 93.130 173.940 ;
        RECT 130.265 173.925 130.595 173.940 ;
        RECT 42.690 173.585 44.270 173.915 ;
        RECT 77.365 173.560 77.695 173.575 ;
        RECT 89.070 173.560 89.450 173.570 ;
        RECT 77.365 173.260 89.450 173.560 ;
        RECT 77.365 173.245 77.695 173.260 ;
        RECT 89.070 173.250 89.450 173.260 ;
        RECT 89.990 173.560 90.370 173.570 ;
        RECT 93.670 173.560 94.050 173.570 ;
        RECT 89.990 173.260 94.050 173.560 ;
        RECT 89.990 173.250 90.370 173.260 ;
        RECT 93.670 173.250 94.050 173.260 ;
        RECT 94.385 173.560 94.715 173.575 ;
        RECT 95.305 173.560 95.635 173.575 ;
        RECT 94.385 173.260 95.635 173.560 ;
        RECT 94.385 173.245 94.715 173.260 ;
        RECT 95.305 173.245 95.635 173.260 ;
        RECT 97.145 173.560 97.475 173.575 ;
        RECT 106.805 173.560 107.135 173.575 ;
        RECT 97.145 173.260 107.135 173.560 ;
        RECT 97.145 173.245 97.475 173.260 ;
        RECT 106.805 173.245 107.135 173.260 ;
        RECT 63.105 172.880 63.435 172.895 ;
        RECT 71.385 172.880 71.715 172.895 ;
        RECT 63.105 172.580 71.715 172.880 ;
        RECT 63.105 172.565 63.435 172.580 ;
        RECT 71.385 172.565 71.715 172.580 ;
        RECT 73.225 172.880 73.555 172.895 ;
        RECT 76.445 172.880 76.775 172.895 ;
        RECT 100.825 172.880 101.155 172.895 ;
        RECT 125.665 172.880 125.995 172.895 ;
        RECT 73.225 172.580 76.775 172.880 ;
        RECT 73.225 172.565 73.555 172.580 ;
        RECT 76.445 172.565 76.775 172.580 ;
        RECT 77.150 172.580 101.155 172.880 ;
        RECT 62.185 172.200 62.515 172.215 ;
        RECT 66.325 172.200 66.655 172.215 ;
        RECT 62.185 171.900 66.655 172.200 ;
        RECT 62.185 171.885 62.515 171.900 ;
        RECT 66.325 171.885 66.655 171.900 ;
        RECT 68.625 172.200 68.955 172.215 ;
        RECT 77.150 172.200 77.450 172.580 ;
        RECT 100.825 172.565 101.155 172.580 ;
        RECT 103.140 172.580 125.995 172.880 ;
        RECT 103.140 172.215 103.440 172.580 ;
        RECT 125.665 172.565 125.995 172.580 ;
        RECT 68.625 171.900 77.450 172.200 ;
        RECT 82.885 172.200 83.215 172.215 ;
        RECT 88.405 172.200 88.735 172.215 ;
        RECT 82.885 171.900 88.735 172.200 ;
        RECT 68.625 171.885 68.955 171.900 ;
        RECT 82.885 171.885 83.215 171.900 ;
        RECT 88.405 171.885 88.735 171.900 ;
        RECT 89.070 172.200 89.450 172.210 ;
        RECT 101.285 172.200 101.615 172.215 ;
        RECT 103.125 172.200 103.455 172.215 ;
        RECT 89.070 171.900 100.680 172.200 ;
        RECT 89.070 171.890 89.450 171.900 ;
        RECT 100.380 171.535 100.680 171.900 ;
        RECT 101.285 171.900 103.455 172.200 ;
        RECT 101.285 171.885 101.615 171.900 ;
        RECT 103.125 171.885 103.455 171.900 ;
        RECT 103.790 172.200 104.170 172.210 ;
        RECT 144.930 172.200 145.430 172.350 ;
        RECT 103.790 171.900 145.430 172.200 ;
        RECT 103.790 171.890 104.170 171.900 ;
        RECT 144.930 171.750 145.430 171.900 ;
        RECT 88.150 171.520 88.530 171.530 ;
        RECT 99.445 171.520 99.775 171.535 ;
        RECT 88.150 171.220 99.775 171.520 ;
        RECT 88.150 171.210 88.530 171.220 ;
        RECT 99.445 171.205 99.775 171.220 ;
        RECT 100.365 171.205 100.695 171.535 ;
        RECT 101.285 171.520 101.615 171.535 ;
        RECT 101.950 171.520 102.330 171.530 ;
        RECT 101.285 171.220 102.330 171.520 ;
        RECT 101.285 171.205 101.615 171.220 ;
        RECT 101.950 171.210 102.330 171.220 ;
        RECT 45.990 170.865 47.570 171.195 ;
        RECT 86.310 170.840 86.690 170.850 ;
        RECT 89.325 170.840 89.655 170.855 ;
        RECT 48.630 170.540 85.730 170.840 ;
        RECT 44.705 170.160 45.035 170.175 ;
        RECT 48.630 170.160 48.930 170.540 ;
        RECT 71.845 170.170 72.175 170.175 ;
        RECT 71.590 170.160 72.175 170.170 ;
        RECT 44.705 169.860 48.930 170.160 ;
        RECT 71.390 169.860 72.175 170.160 ;
        RECT 85.430 170.160 85.730 170.540 ;
        RECT 86.310 170.540 89.655 170.840 ;
        RECT 86.310 170.530 86.690 170.540 ;
        RECT 89.325 170.525 89.655 170.540 ;
        RECT 91.625 170.840 91.955 170.855 ;
        RECT 96.225 170.840 96.555 170.855 ;
        RECT 91.625 170.540 96.555 170.840 ;
        RECT 91.625 170.525 91.955 170.540 ;
        RECT 96.225 170.525 96.555 170.540 ;
        RECT 98.065 170.840 98.395 170.855 ;
        RECT 99.190 170.840 99.570 170.850 ;
        RECT 98.065 170.540 99.570 170.840 ;
        RECT 98.065 170.525 98.395 170.540 ;
        RECT 99.190 170.530 99.570 170.540 ;
        RECT 94.385 170.160 94.715 170.175 ;
        RECT 85.430 169.860 94.715 170.160 ;
        RECT 44.705 169.845 45.035 169.860 ;
        RECT 71.590 169.850 72.175 169.860 ;
        RECT 71.845 169.845 72.175 169.850 ;
        RECT 94.385 169.845 94.715 169.860 ;
        RECT 95.510 170.160 95.890 170.170 ;
        RECT 96.225 170.160 96.555 170.175 ;
        RECT 103.125 170.160 103.455 170.175 ;
        RECT 95.510 169.860 103.455 170.160 ;
        RECT 95.510 169.850 95.890 169.860 ;
        RECT 96.225 169.845 96.555 169.860 ;
        RECT 103.125 169.845 103.455 169.860 ;
        RECT 107.265 170.160 107.595 170.175 ;
        RECT 136.245 170.160 136.575 170.175 ;
        RECT 107.265 169.860 136.575 170.160 ;
        RECT 107.265 169.845 107.595 169.860 ;
        RECT 136.245 169.845 136.575 169.860 ;
        RECT 50.685 169.480 51.015 169.495 ;
        RECT 85.185 169.480 85.515 169.495 ;
        RECT 50.685 169.180 85.515 169.480 ;
        RECT 50.685 169.165 51.015 169.180 ;
        RECT 85.185 169.165 85.515 169.180 ;
        RECT 87.230 169.480 87.610 169.490 ;
        RECT 90.910 169.480 91.290 169.490 ;
        RECT 126.585 169.480 126.915 169.495 ;
        RECT 87.230 169.180 89.410 169.480 ;
        RECT 87.230 169.170 87.610 169.180 ;
        RECT 21.640 168.800 22.140 168.950 ;
        RECT 25.385 168.800 25.715 168.815 ;
        RECT 21.640 168.500 25.715 168.800 ;
        RECT 21.640 168.350 22.140 168.500 ;
        RECT 25.385 168.485 25.715 168.500 ;
        RECT 68.625 168.800 68.955 168.815 ;
        RECT 84.725 168.800 85.055 168.815 ;
        RECT 68.625 168.500 85.055 168.800 ;
        RECT 89.110 168.800 89.410 169.180 ;
        RECT 90.910 169.180 126.915 169.480 ;
        RECT 90.910 169.170 91.290 169.180 ;
        RECT 126.585 169.165 126.915 169.180 ;
        RECT 144.930 168.800 145.430 168.950 ;
        RECT 89.110 168.500 97.690 168.800 ;
        RECT 68.625 168.485 68.955 168.500 ;
        RECT 84.725 168.485 85.055 168.500 ;
        RECT 42.690 168.145 44.270 168.475 ;
        RECT 72.765 168.120 73.095 168.135 ;
        RECT 80.585 168.120 80.915 168.135 ;
        RECT 72.765 167.820 80.915 168.120 ;
        RECT 72.765 167.805 73.095 167.820 ;
        RECT 80.585 167.805 80.915 167.820 ;
        RECT 83.345 168.120 83.675 168.135 ;
        RECT 94.385 168.120 94.715 168.135 ;
        RECT 83.345 167.820 94.715 168.120 ;
        RECT 97.390 168.120 97.690 168.500 ;
        RECT 132.350 168.500 145.430 168.800 ;
        RECT 132.350 168.120 132.650 168.500 ;
        RECT 144.930 168.350 145.430 168.500 ;
        RECT 97.390 167.820 132.650 168.120 ;
        RECT 83.345 167.805 83.675 167.820 ;
        RECT 94.385 167.805 94.715 167.820 ;
        RECT 54.365 167.440 54.695 167.455 ;
        RECT 102.205 167.440 102.535 167.455 ;
        RECT 54.365 167.140 102.535 167.440 ;
        RECT 54.365 167.125 54.695 167.140 ;
        RECT 102.205 167.125 102.535 167.140 ;
        RECT 65.865 166.760 66.195 166.775 ;
        RECT 98.525 166.760 98.855 166.775 ;
        RECT 65.865 166.460 98.855 166.760 ;
        RECT 65.865 166.445 66.195 166.460 ;
        RECT 98.525 166.445 98.855 166.460 ;
        RECT 70.465 166.080 70.795 166.095 ;
        RECT 108.185 166.080 108.515 166.095 ;
        RECT 70.465 165.780 108.515 166.080 ;
        RECT 70.465 165.765 70.795 165.780 ;
        RECT 108.185 165.765 108.515 165.780 ;
        RECT 45.990 165.425 47.570 165.755 ;
        RECT 65.405 165.400 65.735 165.415 ;
        RECT 78.745 165.400 79.075 165.415 ;
        RECT 65.405 165.100 79.075 165.400 ;
        RECT 65.405 165.085 65.735 165.100 ;
        RECT 78.745 165.085 79.075 165.100 ;
        RECT 84.470 165.400 84.850 165.410 ;
        RECT 85.185 165.400 85.515 165.415 ;
        RECT 84.470 165.100 85.515 165.400 ;
        RECT 84.470 165.090 84.850 165.100 ;
        RECT 85.185 165.085 85.515 165.100 ;
        RECT 87.945 165.400 88.275 165.415 ;
        RECT 93.005 165.400 93.335 165.415 ;
        RECT 87.945 165.100 93.335 165.400 ;
        RECT 87.945 165.085 88.275 165.100 ;
        RECT 93.005 165.085 93.335 165.100 ;
        RECT 97.350 165.400 97.730 165.410 ;
        RECT 129.345 165.400 129.675 165.415 ;
        RECT 97.350 165.100 129.675 165.400 ;
        RECT 97.350 165.090 97.730 165.100 ;
        RECT 129.345 165.085 129.675 165.100 ;
        RECT 132.105 165.400 132.435 165.415 ;
        RECT 144.930 165.400 145.430 165.550 ;
        RECT 132.105 165.100 145.430 165.400 ;
        RECT 132.105 165.085 132.435 165.100 ;
        RECT 144.930 164.950 145.430 165.100 ;
        RECT 74.145 164.720 74.475 164.735 ;
        RECT 90.910 164.720 91.290 164.730 ;
        RECT 74.145 164.420 91.290 164.720 ;
        RECT 74.145 164.405 74.475 164.420 ;
        RECT 90.910 164.410 91.290 164.420 ;
        RECT 91.830 164.720 92.210 164.730 ;
        RECT 106.805 164.720 107.135 164.735 ;
        RECT 91.830 164.420 107.135 164.720 ;
        RECT 91.830 164.410 92.210 164.420 ;
        RECT 106.805 164.405 107.135 164.420 ;
        RECT 67.705 164.040 68.035 164.055 ;
        RECT 129.805 164.040 130.135 164.055 ;
        RECT 67.705 163.740 130.135 164.040 ;
        RECT 67.705 163.725 68.035 163.740 ;
        RECT 129.805 163.725 130.135 163.740 ;
        RECT 83.550 163.360 83.930 163.370 ;
        RECT 107.265 163.360 107.595 163.375 ;
        RECT 83.550 163.060 107.595 163.360 ;
        RECT 83.550 163.050 83.930 163.060 ;
        RECT 107.265 163.045 107.595 163.060 ;
        RECT 85.390 162.000 85.770 162.010 ;
        RECT 144.930 162.000 145.430 162.150 ;
        RECT 85.390 161.700 145.430 162.000 ;
        RECT 85.390 161.690 85.770 161.700 ;
        RECT 144.930 161.550 145.430 161.700 ;
        RECT 79.205 160.640 79.535 160.655 ;
        RECT 95.765 160.640 96.095 160.655 ;
        RECT 79.205 160.340 96.095 160.640 ;
        RECT 79.205 160.325 79.535 160.340 ;
        RECT 95.765 160.325 96.095 160.340 ;
        RECT 72.305 158.600 72.635 158.615 ;
        RECT 144.930 158.600 145.430 158.750 ;
        RECT 72.305 158.300 145.430 158.600 ;
        RECT 72.305 158.285 72.635 158.300 ;
        RECT 144.930 158.150 145.430 158.300 ;
        RECT 71.385 156.560 71.715 156.575 ;
        RECT 71.385 156.260 135.410 156.560 ;
        RECT 71.385 156.245 71.715 156.260 ;
        RECT 73.685 155.880 74.015 155.895 ;
        RECT 134.405 155.880 134.735 155.895 ;
        RECT 73.685 155.580 134.735 155.880 ;
        RECT 73.685 155.565 74.015 155.580 ;
        RECT 134.405 155.565 134.735 155.580 ;
        RECT 135.110 155.200 135.410 156.260 ;
        RECT 144.930 155.200 145.430 155.350 ;
        RECT 135.110 154.900 145.430 155.200 ;
        RECT 144.930 154.750 145.430 154.900 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 42.680 165.350 44.280 209.350 ;
        RECT 45.980 165.350 47.580 209.350 ;
        RECT 93.695 202.485 94.025 202.815 ;
        RECT 71.615 201.125 71.945 201.455 ;
        RECT 68.855 199.085 69.185 199.415 ;
        RECT 68.870 191.255 69.170 199.085 ;
        RECT 68.855 190.925 69.185 191.255 ;
        RECT 71.630 170.175 71.930 201.125 ;
        RECT 87.255 198.405 87.585 198.735 ;
        RECT 83.575 196.365 83.905 196.695 ;
        RECT 83.590 178.335 83.890 196.365 ;
        RECT 86.335 184.805 86.665 185.135 ;
        RECT 85.415 181.405 85.745 181.735 ;
        RECT 84.495 179.365 84.825 179.695 ;
        RECT 83.575 178.005 83.905 178.335 ;
        RECT 71.615 169.845 71.945 170.175 ;
        RECT 83.590 163.375 83.890 178.005 ;
        RECT 84.510 165.415 84.810 179.365 ;
        RECT 84.495 165.085 84.825 165.415 ;
        RECT 83.575 163.045 83.905 163.375 ;
        RECT 85.430 162.015 85.730 181.405 ;
        RECT 86.350 170.855 86.650 184.805 ;
        RECT 87.270 181.735 87.570 198.405 ;
        RECT 90.015 195.685 90.345 196.015 ;
        RECT 88.175 186.845 88.505 187.175 ;
        RECT 88.190 182.415 88.490 186.845 ;
        RECT 89.095 185.485 89.425 185.815 ;
        RECT 88.175 182.085 88.505 182.415 ;
        RECT 87.255 181.405 87.585 181.735 ;
        RECT 87.255 175.965 87.585 176.295 ;
        RECT 86.335 170.525 86.665 170.855 ;
        RECT 87.270 169.495 87.570 175.965 ;
        RECT 88.190 171.535 88.490 182.085 ;
        RECT 89.110 173.575 89.410 185.485 ;
        RECT 90.030 179.695 90.330 195.685 ;
        RECT 91.855 188.205 92.185 188.535 ;
        RECT 90.015 179.365 90.345 179.695 ;
        RECT 90.935 179.365 91.265 179.695 ;
        RECT 90.015 176.645 90.345 176.975 ;
        RECT 90.030 173.575 90.330 176.645 ;
        RECT 89.095 173.245 89.425 173.575 ;
        RECT 90.015 173.245 90.345 173.575 ;
        RECT 89.110 172.215 89.410 173.245 ;
        RECT 89.095 171.885 89.425 172.215 ;
        RECT 88.175 171.205 88.505 171.535 ;
        RECT 90.950 169.495 91.250 179.365 ;
        RECT 87.255 169.165 87.585 169.495 ;
        RECT 90.935 169.165 91.265 169.495 ;
        RECT 90.950 164.735 91.250 169.165 ;
        RECT 91.870 164.735 92.170 188.205 ;
        RECT 93.710 187.175 94.010 202.485 ;
        RECT 96.455 199.085 96.785 199.415 ;
        RECT 95.535 195.005 95.865 195.335 ;
        RECT 93.695 186.845 94.025 187.175 ;
        RECT 92.775 182.085 93.105 182.415 ;
        RECT 92.790 174.255 93.090 182.085 ;
        RECT 93.710 175.615 94.010 186.845 ;
        RECT 94.615 178.005 94.945 178.335 ;
        RECT 93.695 175.285 94.025 175.615 ;
        RECT 93.695 174.605 94.025 174.935 ;
        RECT 92.775 173.925 93.105 174.255 ;
        RECT 93.710 173.575 94.010 174.605 ;
        RECT 93.695 173.245 94.025 173.575 ;
        RECT 94.630 168.660 94.930 178.005 ;
        RECT 95.550 170.175 95.850 195.005 ;
        RECT 96.470 176.295 96.770 199.085 ;
        RECT 99.215 196.365 99.545 196.695 ;
        RECT 97.375 195.005 97.705 195.335 ;
        RECT 96.455 175.965 96.785 176.295 ;
        RECT 96.455 174.920 96.785 174.935 ;
        RECT 97.390 174.920 97.690 195.005 ;
        RECT 98.295 191.605 98.625 191.935 ;
        RECT 98.310 181.735 98.610 191.605 ;
        RECT 98.295 181.405 98.625 181.735 ;
        RECT 96.455 174.620 97.690 174.920 ;
        RECT 96.455 174.605 96.785 174.620 ;
        RECT 99.230 170.855 99.530 196.365 ;
        RECT 101.975 195.685 102.305 196.015 ;
        RECT 100.135 188.205 100.465 188.535 ;
        RECT 100.150 178.335 100.450 188.205 ;
        RECT 100.135 178.005 100.465 178.335 ;
        RECT 101.990 171.535 102.290 195.685 ;
        RECT 103.815 189.565 104.145 189.895 ;
        RECT 103.830 172.215 104.130 189.565 ;
        RECT 124.975 184.125 125.305 184.455 ;
        RECT 124.990 175.615 125.290 184.125 ;
        RECT 124.975 175.285 125.305 175.615 ;
        RECT 103.815 171.885 104.145 172.215 ;
        RECT 101.975 171.205 102.305 171.535 ;
        RECT 99.215 170.525 99.545 170.855 ;
        RECT 95.535 169.845 95.865 170.175 ;
        RECT 94.630 168.360 97.690 168.660 ;
        RECT 97.390 165.415 97.690 168.360 ;
        RECT 97.375 165.085 97.705 165.415 ;
        RECT 90.935 164.405 91.265 164.735 ;
        RECT 91.855 164.405 92.185 164.735 ;
        RECT 85.415 161.685 85.745 162.015 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

