VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 54.135 151.435 54.305 151.625 ;
        RECT 56.435 151.435 56.605 151.625 ;
        RECT 56.895 151.435 57.065 151.625 ;
        RECT 60.115 151.435 60.285 151.625 ;
        RECT 61.955 151.435 62.125 151.625 ;
        RECT 62.415 151.455 62.585 151.625 ;
        RECT 62.420 151.435 62.585 151.455 ;
        RECT 66.550 151.435 66.720 151.625 ;
        RECT 69.310 151.435 69.480 151.625 ;
        RECT 69.775 151.455 69.945 151.625 ;
        RECT 69.805 151.435 69.945 151.455 ;
        RECT 72.535 151.435 72.705 151.625 ;
        RECT 75.730 151.435 75.900 151.625 ;
        RECT 80.365 151.480 80.525 151.590 ;
        RECT 90.015 151.435 90.185 151.625 ;
        RECT 90.480 151.435 90.650 151.625 ;
        RECT 95.990 151.435 96.160 151.625 ;
        RECT 105.195 151.435 105.365 151.625 ;
        RECT 107.495 151.435 107.665 151.625 ;
        RECT 107.955 151.435 108.125 151.625 ;
        RECT 117.155 151.435 117.325 151.625 ;
        RECT 118.995 151.455 119.165 151.625 ;
        RECT 118.995 151.435 119.195 151.455 ;
        RECT 123.585 151.435 123.755 151.625 ;
        RECT 124.975 151.435 125.145 151.625 ;
        RECT 53.995 150.625 55.365 151.435 ;
        RECT 55.385 150.525 56.735 151.435 ;
        RECT 56.755 150.755 58.585 151.435 ;
        RECT 57.240 150.525 58.585 150.755 ;
        RECT 58.595 150.755 60.425 151.435 ;
        RECT 60.435 150.755 62.265 151.435 ;
        RECT 62.420 150.755 64.255 151.435 ;
        RECT 58.595 150.525 59.940 150.755 ;
        RECT 60.435 150.525 61.780 150.755 ;
        RECT 63.325 150.525 64.255 150.755 ;
        RECT 64.675 150.525 66.865 151.435 ;
        RECT 66.885 150.565 67.315 151.350 ;
        RECT 67.435 150.525 69.625 151.435 ;
        RECT 69.805 150.615 72.375 151.435 ;
        RECT 72.395 150.755 75.605 151.435 ;
        RECT 70.785 150.525 72.375 150.615 ;
        RECT 74.470 150.525 75.605 150.755 ;
        RECT 75.670 150.525 79.745 151.435 ;
        RECT 79.765 150.565 80.195 151.350 ;
        RECT 81.220 150.755 90.325 151.435 ;
        RECT 90.335 150.755 92.610 151.435 ;
        RECT 91.240 150.525 92.610 150.755 ;
        RECT 92.645 150.565 93.075 151.350 ;
        RECT 93.385 150.525 96.305 151.435 ;
        RECT 96.400 150.755 105.505 151.435 ;
        RECT 105.525 150.565 105.955 151.350 ;
        RECT 105.975 150.525 107.790 151.435 ;
        RECT 107.815 150.755 116.920 151.435 ;
        RECT 117.025 150.525 118.375 151.435 ;
        RECT 118.405 150.565 118.835 151.350 ;
        RECT 118.995 150.755 122.525 151.435 ;
        RECT 119.700 150.525 122.525 150.755 ;
        RECT 122.535 150.655 123.905 151.435 ;
        RECT 123.915 150.625 125.285 151.435 ;
      LAYER nwell ;
        RECT 53.800 147.405 125.480 150.235 ;
      LAYER pwell ;
        RECT 56.495 147.025 57.445 147.115 ;
        RECT 53.995 146.205 55.365 147.015 ;
        RECT 56.495 146.205 58.425 147.025 ;
        RECT 58.595 146.885 59.940 147.115 ;
        RECT 61.575 147.025 62.525 147.115 ;
        RECT 58.595 146.205 60.425 146.885 ;
        RECT 60.595 146.205 62.525 147.025 ;
        RECT 65.020 146.915 66.405 147.115 ;
        RECT 62.735 146.235 66.405 146.915 ;
        RECT 66.885 146.290 67.315 147.075 ;
        RECT 54.135 145.995 54.305 146.205 ;
        RECT 58.275 146.185 58.425 146.205 ;
        RECT 55.525 146.050 55.685 146.160 ;
        RECT 56.895 145.995 57.065 146.185 ;
        RECT 57.350 145.995 57.520 146.185 ;
        RECT 58.275 146.015 58.445 146.185 ;
        RECT 58.730 145.995 58.900 146.185 ;
        RECT 60.115 146.015 60.285 146.205 ;
        RECT 60.595 146.185 60.745 146.205 ;
        RECT 60.575 146.015 60.745 146.185 ;
        RECT 61.950 145.995 62.120 146.185 ;
        RECT 62.875 146.015 63.045 146.235 ;
        RECT 65.035 146.205 66.405 146.235 ;
        RECT 67.795 146.205 71.465 147.115 ;
        RECT 71.475 146.885 73.065 147.115 ;
        RECT 71.475 146.205 75.145 146.885 ;
        RECT 75.240 146.205 84.345 146.885 ;
        RECT 84.355 146.205 88.455 147.115 ;
        RECT 88.495 146.205 92.165 147.115 ;
        RECT 92.645 146.290 93.075 147.075 ;
        RECT 96.515 146.885 100.445 147.115 ;
        RECT 110.500 146.885 113.325 147.115 ;
        RECT 114.180 146.885 117.005 147.115 ;
        RECT 93.095 146.205 95.835 146.885 ;
        RECT 96.030 146.205 100.445 146.885 ;
        RECT 100.455 146.205 109.560 146.885 ;
        RECT 109.795 146.205 113.325 146.885 ;
        RECT 113.475 146.205 117.005 146.885 ;
        RECT 117.025 146.205 118.375 147.115 ;
        RECT 118.405 146.290 118.835 147.075 ;
        RECT 119.700 146.885 122.525 147.115 ;
        RECT 118.995 146.205 122.525 146.885 ;
        RECT 122.535 146.205 123.905 146.985 ;
        RECT 123.915 146.205 125.285 147.015 ;
        RECT 53.995 145.185 55.365 145.995 ;
        RECT 55.375 145.315 57.205 145.995 ;
        RECT 55.375 145.085 56.720 145.315 ;
        RECT 57.235 145.085 58.585 145.995 ;
        RECT 58.615 145.085 59.965 145.995 ;
        RECT 60.430 145.765 62.120 145.995 ;
        RECT 62.275 145.965 63.670 145.995 ;
        RECT 64.715 145.965 64.885 146.185 ;
        RECT 65.175 146.015 65.345 146.185 ;
        RECT 66.550 146.045 66.670 146.155 ;
        RECT 67.470 146.045 67.590 146.155 ;
        RECT 67.940 146.015 68.110 146.205 ;
        RECT 65.205 145.995 65.345 146.015 ;
        RECT 70.235 145.995 70.405 146.185 ;
        RECT 74.830 146.015 75.000 146.205 ;
        RECT 79.435 145.995 79.605 146.185 ;
        RECT 80.365 146.040 80.525 146.150 ;
        RECT 81.275 145.995 81.445 146.185 ;
        RECT 84.035 146.015 84.205 146.205 ;
        RECT 84.500 146.015 84.670 146.205 ;
        RECT 91.850 146.015 92.020 146.205 ;
        RECT 92.310 146.045 92.430 146.155 ;
        RECT 93.235 146.015 93.405 146.205 ;
        RECT 96.030 146.185 96.140 146.205 ;
        RECT 100.595 146.185 100.765 146.205 ;
        RECT 109.795 146.185 109.995 146.205 ;
        RECT 113.475 146.185 113.675 146.205 ;
        RECT 95.970 146.015 96.140 146.185 ;
        RECT 99.215 145.995 99.385 146.185 ;
        RECT 100.590 146.015 100.765 146.185 ;
        RECT 100.590 145.995 100.760 146.015 ;
        RECT 101.060 145.995 101.230 146.185 ;
        RECT 104.745 146.040 104.905 146.150 ;
        RECT 109.335 146.015 109.505 146.185 ;
        RECT 109.305 145.995 109.505 146.015 ;
        RECT 109.795 145.995 109.965 146.185 ;
        RECT 113.475 146.015 113.645 146.185 ;
        RECT 118.075 146.015 118.245 146.205 ;
        RECT 118.995 146.185 119.195 146.205 ;
        RECT 118.995 146.015 119.165 146.185 ;
        RECT 119.915 145.995 120.085 146.185 ;
        RECT 123.130 145.995 123.300 146.185 ;
        RECT 123.595 146.155 123.765 146.205 ;
        RECT 123.590 146.045 123.765 146.155 ;
        RECT 123.595 146.015 123.765 146.045 ;
        RECT 124.975 145.995 125.145 146.205 ;
        RECT 60.430 145.085 62.265 145.765 ;
        RECT 62.275 145.285 65.010 145.965 ;
        RECT 62.275 145.085 63.685 145.285 ;
        RECT 65.205 145.175 67.775 145.995 ;
        RECT 67.805 145.315 70.545 145.995 ;
        RECT 70.640 145.315 79.745 145.995 ;
        RECT 66.185 145.085 67.775 145.175 ;
        RECT 79.765 145.125 80.195 145.910 ;
        RECT 81.135 145.315 90.240 145.995 ;
        RECT 90.420 145.315 99.525 145.995 ;
        RECT 99.555 145.085 100.905 145.995 ;
        RECT 100.915 145.085 104.515 145.995 ;
        RECT 105.525 145.125 105.955 145.910 ;
        RECT 105.975 145.315 109.505 145.995 ;
        RECT 105.975 145.085 108.800 145.315 ;
        RECT 109.665 145.085 111.015 145.995 ;
        RECT 111.120 145.315 120.225 145.995 ;
        RECT 120.235 145.085 123.445 145.995 ;
        RECT 123.915 145.185 125.285 145.995 ;
      LAYER nwell ;
        RECT 53.800 141.965 125.480 144.795 ;
      LAYER pwell ;
        RECT 53.995 140.765 55.365 141.575 ;
        RECT 56.780 141.445 58.125 141.675 ;
        RECT 56.295 140.765 58.125 141.445 ;
        RECT 58.135 141.445 59.480 141.675 ;
        RECT 58.135 140.765 59.965 141.445 ;
        RECT 60.915 140.765 62.265 141.675 ;
        RECT 63.415 141.585 64.365 141.675 ;
        RECT 62.435 140.765 64.365 141.585 ;
        RECT 64.575 140.765 66.865 141.675 ;
        RECT 66.885 140.850 67.315 141.635 ;
        RECT 67.335 140.765 68.705 141.545 ;
        RECT 68.725 140.765 71.455 141.675 ;
        RECT 71.475 140.765 74.215 141.445 ;
        RECT 74.320 140.765 83.425 141.445 ;
        RECT 83.520 140.765 92.625 141.445 ;
        RECT 92.645 140.850 93.075 141.635 ;
        RECT 93.095 140.765 97.225 141.675 ;
        RECT 97.255 140.765 98.605 141.675 ;
        RECT 98.615 140.765 107.720 141.445 ;
        RECT 107.815 140.765 116.920 141.445 ;
        RECT 117.015 140.765 118.385 141.545 ;
        RECT 118.405 140.850 118.835 141.635 ;
        RECT 118.865 140.995 122.065 141.675 ;
        RECT 122.560 141.445 123.905 141.675 ;
        RECT 118.865 140.765 121.920 140.995 ;
        RECT 122.075 140.765 123.905 141.445 ;
        RECT 123.915 140.765 125.285 141.575 ;
        RECT 54.135 140.555 54.305 140.765 ;
        RECT 55.525 140.610 55.685 140.720 ;
        RECT 56.435 140.575 56.605 140.765 ;
        RECT 56.895 140.555 57.065 140.745 ;
        RECT 57.350 140.605 57.470 140.715 ;
        RECT 58.275 140.595 58.445 140.745 ;
        RECT 53.995 139.745 55.365 140.555 ;
        RECT 55.375 139.875 57.205 140.555 ;
        RECT 55.375 139.645 56.720 139.875 ;
        RECT 57.675 139.645 58.565 140.595 ;
        RECT 58.745 140.555 58.915 140.745 ;
        RECT 59.655 140.575 59.825 140.765 ;
        RECT 60.120 140.555 60.290 140.745 ;
        RECT 61.030 140.575 61.200 140.765 ;
        RECT 62.435 140.745 62.585 140.765 ;
        RECT 62.415 140.575 62.585 140.745 ;
        RECT 63.795 140.555 63.965 140.745 ;
        RECT 66.550 140.575 66.720 140.765 ;
        RECT 68.395 140.575 68.565 140.765 ;
        RECT 68.395 140.555 68.560 140.575 ;
        RECT 68.855 140.555 69.025 140.745 ;
        RECT 71.155 140.575 71.325 140.765 ;
        RECT 71.615 140.575 71.785 140.765 ;
        RECT 74.835 140.555 75.005 140.745 ;
        RECT 76.220 140.555 76.390 140.745 ;
        RECT 76.680 140.555 76.850 140.745 ;
        RECT 58.595 139.775 59.965 140.555 ;
        RECT 59.975 139.645 63.645 140.555 ;
        RECT 63.655 139.645 66.405 140.555 ;
        RECT 66.725 139.875 68.560 140.555 ;
        RECT 66.725 139.645 67.655 139.875 ;
        RECT 68.715 139.645 71.925 140.555 ;
        RECT 71.935 139.645 75.145 140.555 ;
        RECT 75.155 139.645 76.505 140.555 ;
        RECT 76.535 139.645 79.455 140.555 ;
        RECT 79.765 139.685 80.195 140.470 ;
        RECT 80.360 140.325 80.530 140.745 ;
        RECT 83.115 140.575 83.285 140.765 ;
        RECT 84.960 140.555 85.130 140.745 ;
        RECT 88.635 140.555 88.805 140.745 ;
        RECT 92.315 140.575 92.485 140.765 ;
        RECT 96.910 140.575 97.080 140.765 ;
        RECT 98.290 140.575 98.460 140.765 ;
        RECT 98.755 140.575 98.925 140.765 ;
        RECT 101.510 140.555 101.680 140.745 ;
        RECT 101.980 140.575 102.150 140.745 ;
        RECT 105.190 140.605 105.310 140.715 ;
        RECT 102.005 140.555 102.150 140.575 ;
        RECT 106.115 140.555 106.285 140.745 ;
        RECT 107.955 140.575 108.125 140.765 ;
        RECT 115.320 140.555 115.490 140.745 ;
        RECT 117.155 140.575 117.325 140.765 ;
        RECT 119.000 140.555 119.170 140.745 ;
        RECT 121.750 140.575 121.920 140.765 ;
        RECT 122.215 140.575 122.385 140.765 ;
        RECT 123.585 140.555 123.755 140.745 ;
        RECT 124.975 140.555 125.145 140.765 ;
        RECT 81.640 140.325 84.800 140.555 ;
        RECT 80.255 139.875 84.800 140.325 ;
        RECT 80.255 139.645 81.630 139.875 ;
        RECT 83.420 139.645 84.800 139.875 ;
        RECT 84.815 139.645 88.470 140.555 ;
        RECT 88.495 139.875 97.600 140.555 ;
        RECT 97.695 139.645 101.825 140.555 ;
        RECT 102.005 139.645 105.045 140.555 ;
        RECT 105.525 139.685 105.955 140.470 ;
        RECT 105.975 139.875 115.080 140.555 ;
        RECT 115.175 139.645 118.720 140.555 ;
        RECT 118.855 139.645 122.400 140.555 ;
        RECT 122.535 139.775 123.905 140.555 ;
        RECT 123.915 139.745 125.285 140.555 ;
      LAYER nwell ;
        RECT 53.800 136.525 125.480 139.355 ;
      LAYER pwell ;
        RECT 55.845 136.145 57.435 136.235 ;
        RECT 53.995 135.325 55.365 136.135 ;
        RECT 55.845 135.325 58.415 136.145 ;
        RECT 59.645 136.005 60.575 136.235 ;
        RECT 54.135 135.115 54.305 135.325 ;
        RECT 58.275 135.305 58.415 135.325 ;
        RECT 58.740 135.325 60.575 136.005 ;
        RECT 60.895 135.325 64.565 136.235 ;
        RECT 65.495 135.325 66.865 136.105 ;
        RECT 66.885 135.410 67.315 136.195 ;
        RECT 67.335 135.325 68.685 136.235 ;
        RECT 68.715 135.325 70.545 136.235 ;
        RECT 70.705 135.325 74.360 136.235 ;
        RECT 75.155 135.325 78.365 136.235 ;
        RECT 78.460 135.325 87.565 136.005 ;
        RECT 87.575 135.325 91.705 136.235 ;
        RECT 92.645 135.410 93.075 136.195 ;
        RECT 93.180 135.325 102.285 136.005 ;
        RECT 102.295 135.325 105.505 136.235 ;
        RECT 105.515 135.325 109.185 136.235 ;
        RECT 109.280 135.325 118.385 136.005 ;
        RECT 118.405 135.410 118.835 136.195 ;
        RECT 119.700 136.005 122.525 136.235 ;
        RECT 118.995 135.325 122.525 136.005 ;
        RECT 122.545 135.325 123.895 136.235 ;
        RECT 123.915 135.325 125.285 136.135 ;
        RECT 58.740 135.305 58.905 135.325 ;
        RECT 55.510 135.165 55.630 135.275 ;
        RECT 56.895 135.115 57.065 135.305 ;
        RECT 57.365 135.115 57.535 135.305 ;
        RECT 58.275 135.135 58.445 135.305 ;
        RECT 58.735 135.135 58.905 135.305 ;
        RECT 59.655 135.115 59.825 135.305 ;
        RECT 61.035 135.115 61.205 135.305 ;
        RECT 61.490 135.165 61.610 135.275 ;
        RECT 61.955 135.115 62.125 135.305 ;
        RECT 64.250 135.135 64.420 135.325 ;
        RECT 64.725 135.170 64.885 135.280 ;
        RECT 66.555 135.135 66.725 135.325 ;
        RECT 67.010 135.165 67.130 135.275 ;
        RECT 66.555 135.115 66.720 135.135 ;
        RECT 67.485 135.115 67.655 135.305 ;
        RECT 68.400 135.135 68.570 135.325 ;
        RECT 68.860 135.135 69.030 135.325 ;
        RECT 70.705 135.305 70.865 135.325 ;
        RECT 70.235 135.115 70.405 135.305 ;
        RECT 70.695 135.135 70.865 135.305 ;
        RECT 73.455 135.135 73.625 135.305 ;
        RECT 73.455 135.115 73.605 135.135 ;
        RECT 73.915 135.115 74.085 135.305 ;
        RECT 74.830 135.165 74.950 135.275 ;
        RECT 75.295 135.135 75.465 135.325 ;
        RECT 79.430 135.115 79.600 135.305 ;
        RECT 83.115 135.115 83.285 135.305 ;
        RECT 83.575 135.115 83.745 135.305 ;
        RECT 87.255 135.135 87.425 135.325 ;
        RECT 87.720 135.135 87.890 135.325 ;
        RECT 91.865 135.170 92.025 135.280 ;
        RECT 95.535 135.115 95.705 135.305 ;
        RECT 95.990 135.165 96.110 135.275 ;
        RECT 101.975 135.135 102.145 135.325 ;
        RECT 105.190 135.305 105.360 135.325 ;
        RECT 105.190 135.135 105.365 135.305 ;
        RECT 105.660 135.135 105.830 135.325 ;
        RECT 105.195 135.115 105.365 135.135 ;
        RECT 106.115 135.115 106.285 135.305 ;
        RECT 109.330 135.165 109.450 135.275 ;
        RECT 109.800 135.115 109.970 135.305 ;
        RECT 113.945 135.160 114.105 135.270 ;
        RECT 118.075 135.135 118.245 135.325 ;
        RECT 118.995 135.305 119.195 135.325 ;
        RECT 118.995 135.135 119.165 135.305 ;
        RECT 122.675 135.135 122.845 135.325 ;
        RECT 123.595 135.115 123.765 135.305 ;
        RECT 124.975 135.115 125.145 135.325 ;
        RECT 53.995 134.305 55.365 135.115 ;
        RECT 55.375 134.435 57.205 135.115 ;
        RECT 55.375 134.205 56.720 134.435 ;
        RECT 57.215 134.335 58.585 135.115 ;
        RECT 58.595 134.335 59.965 135.115 ;
        RECT 59.985 134.205 61.335 135.115 ;
        RECT 61.825 134.205 64.555 135.115 ;
        RECT 64.885 134.435 66.720 135.115 ;
        RECT 64.885 134.205 65.815 134.435 ;
        RECT 67.335 134.335 68.705 135.115 ;
        RECT 68.715 134.205 70.530 135.115 ;
        RECT 71.675 134.295 73.605 135.115 ;
        RECT 73.775 134.435 76.525 135.115 ;
        RECT 71.675 134.205 72.625 134.295 ;
        RECT 75.595 134.205 76.525 134.435 ;
        RECT 76.535 134.205 79.745 135.115 ;
        RECT 79.765 134.245 80.195 135.030 ;
        RECT 80.215 134.205 83.425 135.115 ;
        RECT 83.435 134.205 86.645 135.115 ;
        RECT 86.740 134.435 95.845 135.115 ;
        RECT 96.400 134.435 105.505 135.115 ;
        RECT 105.975 135.085 107.815 135.115 ;
        RECT 105.525 134.245 105.955 135.030 ;
        RECT 105.975 134.435 109.140 135.085 ;
        RECT 106.460 134.405 109.140 134.435 ;
        RECT 106.460 134.205 107.815 134.405 ;
        RECT 109.655 134.205 113.785 135.115 ;
        RECT 114.800 134.435 123.905 135.115 ;
        RECT 123.915 134.305 125.285 135.115 ;
      LAYER nwell ;
        RECT 53.800 131.085 125.480 133.915 ;
      LAYER pwell ;
        RECT 53.995 129.885 55.365 130.695 ;
        RECT 56.295 129.885 57.665 130.665 ;
        RECT 57.675 129.885 59.045 130.665 ;
        RECT 59.055 129.885 60.425 130.665 ;
        RECT 62.865 130.565 63.795 130.795 ;
        RECT 61.960 129.885 63.795 130.565 ;
        RECT 64.115 130.565 65.460 130.795 ;
        RECT 64.115 129.885 65.945 130.565 ;
        RECT 66.885 129.970 67.315 130.755 ;
        RECT 68.255 130.565 69.185 130.795 ;
        RECT 68.255 129.885 72.155 130.565 ;
        RECT 72.855 129.885 74.225 130.665 ;
        RECT 74.235 129.885 76.050 130.795 ;
        RECT 76.160 129.885 85.265 130.565 ;
        RECT 85.275 129.885 88.930 130.795 ;
        RECT 88.955 129.885 92.625 130.795 ;
        RECT 92.645 129.970 93.075 130.755 ;
        RECT 93.105 129.885 95.845 130.565 ;
        RECT 95.855 129.885 99.930 130.795 ;
        RECT 99.995 129.885 109.100 130.565 ;
        RECT 109.280 129.885 118.385 130.565 ;
        RECT 118.405 129.970 118.835 130.755 ;
        RECT 118.855 129.885 121.895 130.795 ;
        RECT 122.075 129.885 123.905 130.795 ;
        RECT 123.915 129.885 125.285 130.695 ;
        RECT 54.135 129.675 54.305 129.885 ;
        RECT 57.355 129.865 57.525 129.885 ;
        RECT 55.525 129.730 55.685 129.840 ;
        RECT 56.895 129.675 57.065 129.865 ;
        RECT 57.350 129.695 57.525 129.865 ;
        RECT 58.735 129.695 58.905 129.885 ;
        RECT 60.115 129.695 60.285 129.885 ;
        RECT 61.960 129.865 62.125 129.885 ;
        RECT 60.575 129.695 60.745 129.865 ;
        RECT 57.350 129.675 57.520 129.695 ;
        RECT 61.495 129.675 61.665 129.865 ;
        RECT 61.955 129.695 62.125 129.865 ;
        RECT 62.880 129.675 63.050 129.865 ;
        RECT 65.635 129.695 65.805 129.885 ;
        RECT 66.105 129.730 66.265 129.840 ;
        RECT 66.560 129.675 66.730 129.865 ;
        RECT 67.485 129.730 67.645 129.840 ;
        RECT 67.935 129.675 68.105 129.865 ;
        RECT 68.670 129.695 68.840 129.885 ;
        RECT 69.590 129.675 69.760 129.865 ;
        RECT 72.530 129.725 72.650 129.835 ;
        RECT 72.995 129.695 73.165 129.885 ;
        RECT 73.730 129.675 73.900 129.865 ;
        RECT 75.755 129.695 75.925 129.885 ;
        RECT 77.590 129.725 77.710 129.835 ;
        RECT 78.055 129.675 78.225 129.865 ;
        RECT 80.360 129.675 80.530 129.865 ;
        RECT 84.955 129.695 85.125 129.885 ;
        RECT 85.420 129.695 85.590 129.885 ;
        RECT 85.880 129.675 86.050 129.865 ;
        RECT 86.310 129.675 86.480 129.865 ;
        RECT 92.310 129.695 92.480 129.885 ;
        RECT 93.240 129.675 93.410 129.865 ;
        RECT 95.535 129.695 95.705 129.885 ;
        RECT 95.995 129.675 96.165 129.865 ;
        RECT 99.700 129.695 99.870 129.885 ;
        RECT 100.135 129.695 100.305 129.885 ;
        RECT 105.195 129.675 105.365 129.865 ;
        RECT 106.105 129.675 106.275 129.865 ;
        RECT 112.555 129.695 112.725 129.865 ;
        RECT 118.075 129.695 118.245 129.885 ;
        RECT 121.750 129.865 121.895 129.885 ;
        RECT 123.590 129.865 123.760 129.885 ;
        RECT 121.750 129.695 121.925 129.865 ;
        RECT 123.590 129.695 123.765 129.865 ;
        RECT 112.555 129.675 112.695 129.695 ;
        RECT 121.755 129.675 121.925 129.695 ;
        RECT 123.595 129.675 123.765 129.695 ;
        RECT 124.975 129.675 125.145 129.885 ;
        RECT 53.995 128.865 55.365 129.675 ;
        RECT 55.375 128.995 57.205 129.675 ;
        RECT 55.375 128.765 56.720 128.995 ;
        RECT 57.235 128.765 58.585 129.675 ;
        RECT 58.725 128.765 61.725 129.675 ;
        RECT 62.735 128.995 66.405 129.675 ;
        RECT 62.735 128.765 63.660 128.995 ;
        RECT 66.415 128.765 67.765 129.675 ;
        RECT 67.805 128.765 69.155 129.675 ;
        RECT 69.175 128.995 73.075 129.675 ;
        RECT 73.315 128.995 77.215 129.675 ;
        RECT 77.915 128.995 79.745 129.675 ;
        RECT 69.175 128.765 70.105 128.995 ;
        RECT 73.315 128.765 74.245 128.995 ;
        RECT 78.400 128.765 79.745 128.995 ;
        RECT 79.765 128.805 80.195 129.590 ;
        RECT 80.215 128.765 84.515 129.675 ;
        RECT 84.815 128.765 86.165 129.675 ;
        RECT 86.250 128.765 90.325 129.675 ;
        RECT 90.335 128.765 93.535 129.675 ;
        RECT 93.565 128.995 96.305 129.675 ;
        RECT 96.400 128.995 105.505 129.675 ;
        RECT 105.525 128.805 105.955 129.590 ;
        RECT 105.975 128.995 110.105 129.675 ;
        RECT 105.975 128.765 107.345 128.995 ;
        RECT 110.125 128.855 112.695 129.675 ;
        RECT 112.960 128.995 122.065 129.675 ;
        RECT 122.075 128.995 123.905 129.675 ;
        RECT 123.915 128.865 125.285 129.675 ;
        RECT 110.125 128.765 111.715 128.855 ;
      LAYER nwell ;
        RECT 53.800 125.645 125.480 128.475 ;
      LAYER pwell ;
        RECT 53.995 124.445 55.365 125.255 ;
        RECT 55.375 124.445 56.745 125.225 ;
        RECT 57.235 124.445 58.585 125.355 ;
        RECT 58.725 124.445 61.725 125.355 ;
        RECT 62.275 125.125 63.200 125.355 ;
        RECT 62.275 124.445 65.945 125.125 ;
        RECT 66.885 124.530 67.315 125.315 ;
        RECT 67.335 124.445 68.705 125.225 ;
        RECT 68.715 125.125 69.645 125.355 ;
        RECT 68.715 124.445 72.615 125.125 ;
        RECT 72.855 124.445 74.225 125.225 ;
        RECT 74.695 124.445 76.065 125.225 ;
        RECT 77.005 124.445 79.735 125.355 ;
        RECT 80.215 124.445 84.290 125.355 ;
        RECT 85.275 124.445 88.485 125.355 ;
        RECT 88.495 124.445 90.310 125.355 ;
        RECT 90.435 124.445 92.625 125.355 ;
        RECT 92.645 124.530 93.075 125.315 ;
        RECT 93.180 124.445 102.285 125.125 ;
        RECT 102.305 124.445 105.045 125.125 ;
        RECT 105.055 124.445 114.160 125.125 ;
        RECT 114.255 124.445 117.910 125.355 ;
        RECT 118.405 124.530 118.835 125.315 ;
        RECT 118.855 124.675 122.055 125.355 ;
        RECT 119.000 124.445 122.055 124.675 ;
        RECT 122.075 124.445 123.425 125.355 ;
        RECT 123.915 124.445 125.285 125.255 ;
        RECT 54.135 124.235 54.305 124.445 ;
        RECT 55.525 124.255 55.695 124.445 ;
        RECT 57.350 124.425 57.520 124.445 ;
        RECT 56.890 124.285 57.010 124.395 ;
        RECT 57.350 124.255 57.525 124.425 ;
        RECT 57.355 124.235 57.525 124.255 ;
        RECT 58.725 124.235 58.895 124.425 ;
        RECT 59.195 124.235 59.365 124.425 ;
        RECT 61.040 124.235 61.210 124.425 ;
        RECT 61.495 124.255 61.665 124.445 ;
        RECT 61.950 124.285 62.070 124.395 ;
        RECT 62.420 124.255 62.590 124.445 ;
        RECT 63.325 124.235 63.495 124.425 ;
        RECT 63.805 124.235 63.975 124.425 ;
        RECT 65.185 124.235 65.355 124.425 ;
        RECT 66.105 124.290 66.265 124.400 ;
        RECT 66.555 124.235 66.725 124.425 ;
        RECT 68.385 124.255 68.555 124.445 ;
        RECT 68.845 124.235 69.015 124.425 ;
        RECT 69.130 124.255 69.300 124.445 ;
        RECT 69.325 124.280 69.485 124.390 ;
        RECT 70.230 124.235 70.400 124.425 ;
        RECT 71.615 124.235 71.785 124.425 ;
        RECT 72.995 124.255 73.165 124.445 ;
        RECT 74.370 124.285 74.490 124.395 ;
        RECT 75.745 124.255 75.915 124.445 ;
        RECT 76.225 124.290 76.385 124.400 ;
        RECT 77.135 124.235 77.305 124.425 ;
        RECT 79.435 124.255 79.605 124.445 ;
        RECT 84.060 124.425 84.230 124.445 ;
        RECT 85.415 124.425 85.585 124.445 ;
        RECT 79.890 124.285 80.010 124.395 ;
        RECT 82.655 124.235 82.825 124.425 ;
        RECT 84.025 124.255 84.230 124.425 ;
        RECT 84.505 124.290 84.665 124.400 ;
        RECT 85.405 124.255 85.585 124.425 ;
        RECT 84.025 124.235 84.195 124.255 ;
        RECT 85.405 124.235 85.575 124.255 ;
        RECT 85.885 124.235 86.055 124.425 ;
        RECT 88.165 124.235 88.335 124.425 ;
        RECT 89.545 124.235 89.715 124.425 ;
        RECT 90.015 124.235 90.185 124.445 ;
        RECT 92.310 124.255 92.480 124.445 ;
        RECT 96.915 124.255 97.085 124.425 ;
        RECT 96.915 124.235 97.075 124.255 ;
        RECT 100.135 124.235 100.305 124.425 ;
        RECT 100.605 124.280 100.765 124.390 ;
        RECT 101.975 124.255 102.145 124.445 ;
        RECT 104.735 124.255 104.905 124.445 ;
        RECT 105.195 124.395 105.365 124.445 ;
        RECT 105.190 124.285 105.365 124.395 ;
        RECT 105.195 124.255 105.365 124.285 ;
        RECT 104.705 124.235 104.905 124.255 ;
        RECT 112.090 124.235 112.260 124.425 ;
        RECT 112.560 124.235 112.730 124.425 ;
        RECT 114.400 124.255 114.570 124.445 ;
        RECT 118.070 124.285 118.190 124.395 ;
        RECT 119.000 124.255 119.170 124.445 ;
        RECT 122.220 124.255 122.390 124.445 ;
        RECT 123.595 124.395 123.765 124.425 ;
        RECT 123.590 124.285 123.765 124.395 ;
        RECT 123.595 124.235 123.765 124.285 ;
        RECT 124.975 124.235 125.145 124.445 ;
        RECT 53.995 123.425 55.365 124.235 ;
        RECT 56.295 123.455 57.665 124.235 ;
        RECT 57.675 123.455 59.045 124.235 ;
        RECT 59.055 123.555 60.885 124.235 ;
        RECT 60.895 123.325 62.245 124.235 ;
        RECT 62.275 123.455 63.645 124.235 ;
        RECT 63.655 123.455 65.025 124.235 ;
        RECT 65.035 123.455 66.405 124.235 ;
        RECT 66.425 123.325 67.775 124.235 ;
        RECT 67.795 123.455 69.165 124.235 ;
        RECT 70.115 123.325 71.465 124.235 ;
        RECT 71.475 123.425 76.985 124.235 ;
        RECT 76.995 123.425 79.745 124.235 ;
        RECT 79.765 123.365 80.195 124.150 ;
        RECT 80.245 123.325 82.965 124.235 ;
        RECT 82.975 123.455 84.345 124.235 ;
        RECT 84.355 123.455 85.725 124.235 ;
        RECT 85.735 123.455 87.105 124.235 ;
        RECT 87.115 123.455 88.485 124.235 ;
        RECT 88.495 123.455 89.865 124.235 ;
        RECT 89.875 123.325 93.085 124.235 ;
        RECT 93.420 123.325 97.075 124.235 ;
        RECT 97.235 123.325 100.445 124.235 ;
        RECT 101.375 123.555 104.905 124.235 ;
        RECT 101.375 123.325 104.200 123.555 ;
        RECT 105.525 123.365 105.955 124.150 ;
        RECT 106.335 123.325 112.405 124.235 ;
        RECT 112.560 124.005 114.250 124.235 ;
        RECT 112.415 123.325 114.250 124.005 ;
        RECT 114.800 123.555 123.905 124.235 ;
        RECT 123.915 123.425 125.285 124.235 ;
      LAYER nwell ;
        RECT 53.800 120.205 125.480 123.035 ;
      LAYER pwell ;
        RECT 53.995 119.005 55.365 119.815 ;
        RECT 57.345 119.685 58.275 119.915 ;
        RECT 56.440 119.005 58.275 119.685 ;
        RECT 58.595 119.685 59.960 119.915 ;
        RECT 63.635 119.685 64.565 119.915 ;
        RECT 58.595 119.005 61.805 119.685 ;
        RECT 61.815 119.005 64.565 119.685 ;
        RECT 65.035 119.005 66.850 119.915 ;
        RECT 66.885 119.090 67.315 119.875 ;
        RECT 68.255 119.005 71.175 119.915 ;
        RECT 71.475 119.005 73.305 119.915 ;
        RECT 73.330 119.005 76.985 119.915 ;
        RECT 76.995 119.005 80.665 119.915 ;
        RECT 80.675 119.685 81.595 119.915 ;
        RECT 80.675 119.005 84.260 119.685 ;
        RECT 84.815 119.005 86.645 119.915 ;
        RECT 86.655 119.685 87.585 119.915 ;
        RECT 91.235 119.685 92.165 119.915 ;
        RECT 86.655 119.005 89.405 119.685 ;
        RECT 89.415 119.005 92.165 119.685 ;
        RECT 92.645 119.090 93.075 119.875 ;
        RECT 93.095 119.005 96.305 119.915 ;
        RECT 97.235 119.005 99.985 119.915 ;
        RECT 100.480 119.685 101.825 119.915 ;
        RECT 99.995 119.005 101.825 119.685 ;
        RECT 101.835 119.005 105.310 119.915 ;
        RECT 105.525 119.005 106.875 119.915 ;
        RECT 106.895 119.005 116.000 119.685 ;
        RECT 116.095 119.005 118.305 119.915 ;
        RECT 118.405 119.090 118.835 119.875 ;
        RECT 118.855 119.005 122.065 119.915 ;
        RECT 122.560 119.685 123.905 119.915 ;
        RECT 122.075 119.005 123.905 119.685 ;
        RECT 123.915 119.005 125.285 119.815 ;
        RECT 54.135 118.795 54.305 119.005 ;
        RECT 56.440 118.985 56.605 119.005 ;
        RECT 61.490 118.985 61.660 119.005 ;
        RECT 55.525 118.795 55.695 118.985 ;
        RECT 56.435 118.815 56.605 118.985 ;
        RECT 56.905 118.840 57.065 118.950 ;
        RECT 57.820 118.795 57.990 118.985 ;
        RECT 61.490 118.815 61.665 118.985 ;
        RECT 61.955 118.815 62.125 119.005 ;
        RECT 61.495 118.795 61.665 118.815 ;
        RECT 62.875 118.795 63.045 118.985 ;
        RECT 63.335 118.795 63.505 118.985 ;
        RECT 64.715 118.955 64.885 118.985 ;
        RECT 64.710 118.845 64.885 118.955 ;
        RECT 64.715 118.795 64.885 118.845 ;
        RECT 66.555 118.815 66.725 119.005 ;
        RECT 67.485 118.850 67.645 118.960 ;
        RECT 68.400 118.815 68.570 119.005 ;
        RECT 69.310 118.795 69.480 118.985 ;
        RECT 70.695 118.795 70.865 118.985 ;
        RECT 71.620 118.815 71.790 119.005 ;
        RECT 76.215 118.795 76.385 118.985 ;
        RECT 76.670 118.815 76.840 119.005 ;
        RECT 77.140 118.815 77.310 119.005 ;
        RECT 80.355 118.795 80.525 118.985 ;
        RECT 80.820 118.815 80.990 119.005 ;
        RECT 83.575 118.795 83.745 118.985 ;
        RECT 84.490 118.845 84.610 118.955 ;
        RECT 85.410 118.845 85.530 118.955 ;
        RECT 86.330 118.815 86.500 119.005 ;
        RECT 86.800 118.795 86.970 118.985 ;
        RECT 88.175 118.795 88.345 118.985 ;
        RECT 89.095 118.815 89.265 119.005 ;
        RECT 89.555 118.985 89.725 119.005 ;
        RECT 89.545 118.815 89.725 118.985 ;
        RECT 89.545 118.795 89.715 118.815 ;
        RECT 90.940 118.795 91.110 118.985 ;
        RECT 92.305 118.795 92.475 118.985 ;
        RECT 93.235 118.815 93.405 119.005 ;
        RECT 95.995 118.815 96.165 118.985 ;
        RECT 96.465 118.850 96.625 118.960 ;
        RECT 95.965 118.795 96.165 118.815 ;
        RECT 97.380 118.795 97.550 119.005 ;
        RECT 97.840 118.795 98.010 118.985 ;
        RECT 100.135 118.815 100.305 119.005 ;
        RECT 100.590 118.845 100.710 118.955 ;
        RECT 101.060 118.795 101.230 118.985 ;
        RECT 101.980 118.815 102.150 119.005 ;
        RECT 104.745 118.840 104.905 118.950 ;
        RECT 105.655 118.815 105.825 119.005 ;
        RECT 107.035 118.815 107.205 119.005 ;
        RECT 108.875 118.795 109.045 118.985 ;
        RECT 109.330 118.845 109.450 118.955 ;
        RECT 109.800 118.795 109.970 118.985 ;
        RECT 113.025 118.840 113.185 118.950 ;
        RECT 113.935 118.795 114.105 118.985 ;
        RECT 116.240 118.815 116.410 119.005 ;
        RECT 119.000 118.815 119.170 119.005 ;
        RECT 122.215 118.815 122.385 119.005 ;
        RECT 123.145 118.840 123.305 118.950 ;
        RECT 124.975 118.795 125.145 119.005 ;
        RECT 53.995 117.985 55.365 118.795 ;
        RECT 55.375 118.015 56.745 118.795 ;
        RECT 57.820 118.565 59.510 118.795 ;
        RECT 57.675 117.885 59.510 118.565 ;
        RECT 59.975 118.115 61.805 118.795 ;
        RECT 59.975 117.885 61.320 118.115 ;
        RECT 61.815 118.015 63.185 118.795 ;
        RECT 63.195 118.015 64.565 118.795 ;
        RECT 64.575 117.985 68.245 118.795 ;
        RECT 69.195 117.885 70.545 118.795 ;
        RECT 70.555 117.985 76.065 118.795 ;
        RECT 76.075 117.985 79.745 118.795 ;
        RECT 79.765 117.925 80.195 118.710 ;
        RECT 80.215 118.115 83.425 118.795 ;
        RECT 82.290 117.885 83.425 118.115 ;
        RECT 83.450 117.885 85.265 118.795 ;
        RECT 85.735 117.885 87.085 118.795 ;
        RECT 87.115 118.015 88.485 118.795 ;
        RECT 88.495 118.015 89.865 118.795 ;
        RECT 89.875 117.885 91.225 118.795 ;
        RECT 91.255 118.015 92.625 118.795 ;
        RECT 92.635 118.115 96.165 118.795 ;
        RECT 92.635 117.885 95.460 118.115 ;
        RECT 96.315 117.885 97.665 118.795 ;
        RECT 97.695 117.885 100.445 118.795 ;
        RECT 100.915 118.115 104.500 118.795 ;
        RECT 100.915 117.885 101.835 118.115 ;
        RECT 105.525 117.925 105.955 118.710 ;
        RECT 105.975 117.885 109.185 118.795 ;
        RECT 109.800 118.565 112.855 118.795 ;
        RECT 109.655 117.885 112.855 118.565 ;
        RECT 113.795 118.115 122.900 118.795 ;
        RECT 123.915 117.985 125.285 118.795 ;
      LAYER nwell ;
        RECT 53.800 114.765 125.480 117.595 ;
      LAYER pwell ;
        RECT 53.995 113.565 55.365 114.375 ;
        RECT 56.295 113.565 59.505 114.475 ;
        RECT 59.515 113.565 65.025 114.375 ;
        RECT 65.035 113.565 66.865 114.375 ;
        RECT 66.885 113.650 67.315 114.435 ;
        RECT 67.345 113.565 70.075 114.475 ;
        RECT 70.095 113.565 73.765 114.375 ;
        RECT 74.235 113.565 75.585 114.475 ;
        RECT 75.615 113.565 81.125 114.375 ;
        RECT 81.135 113.565 86.645 114.375 ;
        RECT 87.590 113.565 89.405 114.475 ;
        RECT 90.350 113.565 92.165 114.475 ;
        RECT 92.645 113.650 93.075 114.435 ;
        RECT 93.555 113.565 94.925 114.345 ;
        RECT 94.945 113.565 96.295 114.475 ;
        RECT 96.335 113.565 97.685 114.475 ;
        RECT 97.695 113.565 100.905 114.475 ;
        RECT 101.375 113.565 102.745 114.345 ;
        RECT 102.775 113.565 104.125 114.475 ;
        RECT 104.145 113.565 105.495 114.475 ;
        RECT 105.615 113.565 107.805 114.475 ;
        RECT 108.080 113.565 111.015 114.475 ;
        RECT 111.045 113.565 113.980 114.475 ;
        RECT 114.725 113.795 117.925 114.475 ;
        RECT 114.725 113.565 117.780 113.795 ;
        RECT 118.405 113.650 118.835 114.435 ;
        RECT 118.865 113.795 122.065 114.475 ;
        RECT 122.560 114.245 123.905 114.475 ;
        RECT 118.865 113.565 121.920 113.795 ;
        RECT 122.075 113.565 123.905 114.245 ;
        RECT 123.915 113.565 125.285 114.375 ;
        RECT 54.135 113.355 54.305 113.565 ;
        RECT 55.515 113.355 55.685 113.545 ;
        RECT 56.435 113.375 56.605 113.565 ;
        RECT 57.350 113.405 57.470 113.515 ;
        RECT 58.090 113.355 58.260 113.545 ;
        RECT 59.655 113.375 59.825 113.565 ;
        RECT 61.955 113.355 62.125 113.545 ;
        RECT 65.175 113.375 65.345 113.565 ;
        RECT 66.095 113.355 66.265 113.545 ;
        RECT 68.395 113.375 68.565 113.545 ;
        RECT 69.775 113.375 69.945 113.565 ;
        RECT 70.235 113.375 70.405 113.565 ;
        RECT 68.395 113.355 68.560 113.375 ;
        RECT 71.615 113.355 71.785 113.545 ;
        RECT 72.085 113.400 72.245 113.510 ;
        RECT 73.270 113.355 73.440 113.545 ;
        RECT 73.910 113.405 74.030 113.515 ;
        RECT 75.300 113.375 75.470 113.565 ;
        RECT 75.755 113.375 75.925 113.565 ;
        RECT 77.135 113.355 77.305 113.545 ;
        RECT 81.275 113.375 81.445 113.565 ;
        RECT 81.735 113.355 81.905 113.545 ;
        RECT 82.190 113.405 82.310 113.515 ;
        RECT 82.655 113.355 82.825 113.545 ;
        RECT 85.415 113.355 85.585 113.545 ;
        RECT 86.805 113.410 86.965 113.520 ;
        RECT 87.715 113.375 87.885 113.565 ;
        RECT 88.175 113.355 88.345 113.545 ;
        RECT 89.565 113.410 89.725 113.520 ;
        RECT 90.025 113.400 90.185 113.510 ;
        RECT 90.475 113.375 90.645 113.565 ;
        RECT 90.935 113.355 91.105 113.545 ;
        RECT 92.310 113.405 92.430 113.515 ;
        RECT 92.785 113.400 92.945 113.510 ;
        RECT 93.230 113.405 93.350 113.515 ;
        RECT 94.605 113.355 94.775 113.565 ;
        RECT 95.075 113.375 95.245 113.565 ;
        RECT 96.450 113.375 96.620 113.565 ;
        RECT 98.295 113.375 98.465 113.545 ;
        RECT 98.265 113.355 98.465 113.375 ;
        RECT 98.755 113.355 98.925 113.545 ;
        RECT 100.595 113.375 100.765 113.565 ;
        RECT 101.055 113.515 101.225 113.545 ;
        RECT 101.050 113.405 101.225 113.515 ;
        RECT 101.055 113.355 101.225 113.405 ;
        RECT 101.525 113.355 101.695 113.545 ;
        RECT 102.425 113.375 102.595 113.565 ;
        RECT 103.810 113.545 103.980 113.565 ;
        RECT 103.805 113.375 103.980 113.545 ;
        RECT 103.805 113.355 103.975 113.375 ;
        RECT 104.275 113.355 104.445 113.565 ;
        RECT 106.110 113.405 106.230 113.515 ;
        RECT 106.585 113.355 106.755 113.545 ;
        RECT 107.490 113.375 107.660 113.565 ;
        RECT 108.080 113.545 108.125 113.565 ;
        RECT 113.935 113.545 113.980 113.565 ;
        RECT 107.955 113.375 108.125 113.545 ;
        RECT 108.875 113.355 109.045 113.545 ;
        RECT 112.555 113.355 112.725 113.545 ;
        RECT 113.015 113.355 113.185 113.545 ;
        RECT 113.935 113.375 114.105 113.545 ;
        RECT 114.390 113.405 114.510 113.515 ;
        RECT 114.855 113.355 115.025 113.545 ;
        RECT 117.610 113.375 117.780 113.565 ;
        RECT 118.070 113.405 118.190 113.515 ;
        RECT 121.750 113.375 121.920 113.565 ;
        RECT 122.215 113.375 122.385 113.565 ;
        RECT 124.975 113.355 125.145 113.565 ;
        RECT 53.995 112.545 55.365 113.355 ;
        RECT 55.375 112.545 57.205 113.355 ;
        RECT 57.675 112.675 61.575 113.355 ;
        RECT 57.675 112.445 58.605 112.675 ;
        RECT 61.815 112.545 64.565 113.355 ;
        RECT 64.575 112.445 66.390 113.355 ;
        RECT 66.725 112.675 68.560 113.355 ;
        RECT 66.725 112.445 67.655 112.675 ;
        RECT 68.715 112.445 71.925 113.355 ;
        RECT 72.855 112.675 76.755 113.355 ;
        RECT 72.855 112.445 73.785 112.675 ;
        RECT 76.995 112.545 79.745 113.355 ;
        RECT 79.765 112.485 80.195 113.270 ;
        RECT 80.215 112.445 82.030 113.355 ;
        RECT 82.525 112.445 85.255 113.355 ;
        RECT 85.275 112.545 88.025 113.355 ;
        RECT 88.050 112.445 89.865 113.355 ;
        RECT 90.810 112.445 92.625 113.355 ;
        RECT 93.555 112.575 94.925 113.355 ;
        RECT 94.935 112.675 98.465 113.355 ;
        RECT 94.935 112.445 97.760 112.675 ;
        RECT 98.615 112.575 99.985 113.355 ;
        RECT 99.995 112.575 101.365 113.355 ;
        RECT 101.375 112.575 102.745 113.355 ;
        RECT 102.755 112.575 104.125 113.355 ;
        RECT 104.135 112.575 105.505 113.355 ;
        RECT 105.525 112.485 105.955 113.270 ;
        RECT 106.435 112.575 107.805 113.355 ;
        RECT 107.825 112.445 109.175 113.355 ;
        RECT 109.335 112.445 112.785 113.355 ;
        RECT 112.875 112.675 114.705 113.355 ;
        RECT 114.715 112.675 123.820 113.355 ;
        RECT 113.360 112.445 114.705 112.675 ;
        RECT 123.915 112.545 125.285 113.355 ;
      LAYER nwell ;
        RECT 53.800 109.325 125.480 112.155 ;
      LAYER pwell ;
        RECT 53.995 108.125 55.365 108.935 ;
        RECT 55.375 108.125 57.205 108.935 ;
        RECT 57.215 108.805 58.145 109.035 ;
        RECT 57.215 108.125 61.115 108.805 ;
        RECT 61.355 108.125 64.105 108.935 ;
        RECT 64.115 108.125 65.930 109.035 ;
        RECT 66.885 108.210 67.315 108.995 ;
        RECT 67.645 108.805 68.575 109.035 ;
        RECT 67.645 108.125 69.480 108.805 ;
        RECT 69.635 108.125 71.450 109.035 ;
        RECT 72.395 108.805 73.325 109.035 ;
        RECT 72.395 108.125 76.295 108.805 ;
        RECT 76.545 108.125 77.895 109.035 ;
        RECT 77.915 108.125 79.265 109.035 ;
        RECT 80.215 108.125 82.030 109.035 ;
        RECT 82.065 108.125 83.415 109.035 ;
        RECT 83.435 108.125 84.805 108.935 ;
        RECT 84.815 108.125 86.165 109.035 ;
        RECT 86.195 108.125 91.705 108.935 ;
        RECT 92.645 108.210 93.075 108.995 ;
        RECT 93.095 108.835 94.040 109.035 ;
        RECT 95.375 108.835 96.305 109.035 ;
        RECT 93.095 108.355 96.305 108.835 ;
        RECT 93.095 108.155 96.165 108.355 ;
        RECT 93.095 108.125 94.040 108.155 ;
        RECT 54.135 107.915 54.305 108.125 ;
        RECT 55.515 107.915 55.685 108.125 ;
        RECT 57.630 107.935 57.800 108.125 ;
        RECT 61.495 107.935 61.665 108.125 ;
        RECT 61.680 107.915 61.850 108.105 ;
        RECT 65.175 107.915 65.345 108.105 ;
        RECT 65.635 107.915 65.805 108.125 ;
        RECT 69.315 108.105 69.480 108.125 ;
        RECT 66.105 107.970 66.265 108.080 ;
        RECT 69.315 107.935 69.485 108.105 ;
        RECT 71.155 107.915 71.325 108.125 ;
        RECT 71.625 107.970 71.785 108.080 ;
        RECT 72.810 107.935 72.980 108.125 ;
        RECT 76.675 107.915 76.845 108.125 ;
        RECT 78.980 107.935 79.150 108.125 ;
        RECT 79.445 108.075 79.605 108.080 ;
        RECT 79.430 107.970 79.605 108.075 ;
        RECT 79.430 107.965 79.550 107.970 ;
        RECT 80.355 107.915 80.525 108.105 ;
        RECT 81.735 107.935 81.905 108.125 ;
        RECT 82.195 107.935 82.365 108.125 ;
        RECT 83.575 108.105 83.745 108.125 ;
        RECT 83.110 107.965 83.230 108.075 ;
        RECT 83.575 107.935 83.750 108.105 ;
        RECT 85.880 107.935 86.050 108.125 ;
        RECT 86.335 107.935 86.505 108.125 ;
        RECT 83.580 107.915 83.750 107.935 ;
        RECT 87.255 107.915 87.425 108.105 ;
        RECT 89.100 107.915 89.270 108.105 ;
        RECT 91.865 107.970 92.025 108.080 ;
        RECT 95.530 107.915 95.700 108.105 ;
        RECT 95.995 107.935 96.165 108.155 ;
        RECT 96.315 108.125 98.145 108.935 ;
        RECT 98.615 108.125 101.825 109.035 ;
        RECT 101.850 108.125 105.505 109.035 ;
        RECT 105.515 108.125 107.330 109.035 ;
        RECT 108.405 108.125 111.405 109.035 ;
        RECT 113.320 108.805 114.690 109.035 ;
        RECT 112.415 108.125 114.690 108.805 ;
        RECT 114.725 108.125 117.465 108.805 ;
        RECT 118.405 108.210 118.835 108.995 ;
        RECT 118.935 108.125 121.145 109.035 ;
        RECT 121.155 108.125 123.895 108.805 ;
        RECT 123.915 108.125 125.285 108.935 ;
        RECT 96.455 107.935 96.625 108.125 ;
        RECT 98.290 107.965 98.410 108.075 ;
        RECT 98.745 107.935 98.915 108.125 ;
        RECT 96.000 107.915 96.165 107.935 ;
        RECT 99.220 107.915 99.390 108.105 ;
        RECT 99.675 107.915 99.845 108.105 ;
        RECT 102.435 107.915 102.605 108.105 ;
        RECT 104.285 107.915 104.455 108.105 ;
        RECT 105.190 107.935 105.360 108.125 ;
        RECT 106.125 107.960 106.285 108.070 ;
        RECT 107.035 107.915 107.205 108.125 ;
        RECT 107.505 107.970 107.665 108.080 ;
        RECT 108.415 107.915 108.585 108.105 ;
        RECT 109.795 107.915 109.965 108.105 ;
        RECT 111.175 107.935 111.345 108.125 ;
        RECT 111.645 107.970 111.805 108.080 ;
        RECT 112.560 107.935 112.730 108.125 ;
        RECT 53.995 107.105 55.365 107.915 ;
        RECT 55.375 107.105 58.125 107.915 ;
        RECT 58.365 107.235 62.265 107.915 ;
        RECT 61.335 107.005 62.265 107.235 ;
        RECT 62.275 107.005 65.485 107.915 ;
        RECT 65.495 107.105 71.005 107.915 ;
        RECT 71.015 107.105 76.525 107.915 ;
        RECT 76.535 107.105 79.285 107.915 ;
        RECT 79.765 107.045 80.195 107.830 ;
        RECT 80.215 107.105 82.965 107.915 ;
        RECT 83.435 107.235 87.105 107.915 ;
        RECT 83.435 107.005 84.360 107.235 ;
        RECT 87.115 107.105 88.945 107.915 ;
        RECT 88.955 107.005 91.875 107.915 ;
        RECT 92.370 107.005 95.845 107.915 ;
        RECT 96.000 107.235 97.835 107.915 ;
        RECT 96.905 107.005 97.835 107.235 ;
        RECT 98.155 107.005 99.505 107.915 ;
        RECT 99.535 107.105 102.285 107.915 ;
        RECT 102.310 107.005 104.125 107.915 ;
        RECT 104.135 107.135 105.505 107.915 ;
        RECT 105.525 107.045 105.955 107.830 ;
        RECT 106.895 107.135 108.265 107.915 ;
        RECT 108.275 107.135 109.645 107.915 ;
        RECT 109.735 107.005 113.185 107.915 ;
        RECT 113.470 107.885 113.640 108.105 ;
        RECT 115.785 107.960 115.945 108.070 ;
        RECT 116.695 107.915 116.865 108.105 ;
        RECT 117.155 107.935 117.325 108.125 ;
        RECT 117.625 107.970 117.785 108.080 ;
        RECT 120.830 107.935 121.000 108.125 ;
        RECT 121.295 107.935 121.465 108.125 ;
        RECT 114.670 107.885 115.625 107.915 ;
        RECT 113.345 107.205 115.625 107.885 ;
        RECT 116.555 107.235 119.305 107.915 ;
        RECT 114.670 107.005 115.625 107.205 ;
        RECT 118.375 107.005 119.305 107.235 ;
        RECT 119.315 107.885 120.710 107.915 ;
        RECT 121.755 107.885 121.925 108.105 ;
        RECT 122.215 107.915 122.385 108.105 ;
        RECT 124.975 107.915 125.145 108.125 ;
        RECT 119.315 107.205 122.050 107.885 ;
        RECT 122.075 107.235 123.905 107.915 ;
        RECT 119.315 107.005 120.725 107.205 ;
        RECT 122.560 107.005 123.905 107.235 ;
        RECT 123.915 107.105 125.285 107.915 ;
      LAYER nwell ;
        RECT 53.800 103.885 125.480 106.715 ;
      LAYER pwell ;
        RECT 53.995 102.685 55.365 103.495 ;
        RECT 55.375 102.685 58.125 103.495 ;
        RECT 61.335 103.365 62.265 103.595 ;
        RECT 58.365 102.685 62.265 103.365 ;
        RECT 62.275 102.685 65.025 103.495 ;
        RECT 65.495 102.685 66.845 103.595 ;
        RECT 66.885 102.770 67.315 103.555 ;
        RECT 67.335 102.685 70.545 103.595 ;
        RECT 71.015 103.365 71.945 103.595 ;
        RECT 71.015 102.685 74.915 103.365 ;
        RECT 75.155 102.685 76.505 103.595 ;
        RECT 76.535 102.685 79.285 103.495 ;
        RECT 79.295 102.685 82.505 103.595 ;
        RECT 82.515 102.685 88.025 103.495 ;
        RECT 88.035 102.685 91.705 103.495 ;
        RECT 92.645 102.770 93.075 103.555 ;
        RECT 93.095 103.395 94.040 103.595 ;
        RECT 95.375 103.395 96.305 103.595 ;
        RECT 93.095 102.915 96.305 103.395 ;
        RECT 93.095 102.715 96.165 102.915 ;
        RECT 93.095 102.685 94.040 102.715 ;
        RECT 54.135 102.475 54.305 102.685 ;
        RECT 55.515 102.495 55.685 102.685 ;
        RECT 56.895 102.475 57.065 102.665 ;
        RECT 57.355 102.475 57.525 102.665 ;
        RECT 60.115 102.475 60.285 102.665 ;
        RECT 60.575 102.475 60.745 102.665 ;
        RECT 61.680 102.495 61.850 102.685 ;
        RECT 62.415 102.495 62.585 102.685 ;
        RECT 65.170 102.525 65.290 102.635 ;
        RECT 66.090 102.525 66.210 102.635 ;
        RECT 66.560 102.495 66.730 102.685 ;
        RECT 67.475 102.475 67.645 102.665 ;
        RECT 67.935 102.495 68.105 102.665 ;
        RECT 70.235 102.495 70.405 102.685 ;
        RECT 70.690 102.525 70.810 102.635 ;
        RECT 67.965 102.475 68.105 102.495 ;
        RECT 70.970 102.475 71.140 102.665 ;
        RECT 71.430 102.495 71.600 102.685 ;
        RECT 74.835 102.475 75.005 102.665 ;
        RECT 76.220 102.495 76.390 102.685 ;
        RECT 76.675 102.495 76.845 102.685 ;
        RECT 78.985 102.520 79.145 102.630 ;
        RECT 79.425 102.495 79.595 102.685 ;
        RECT 82.655 102.495 82.825 102.685 ;
        RECT 84.035 102.495 84.205 102.665 ;
        RECT 76.680 102.475 76.845 102.495 ;
        RECT 84.035 102.475 84.195 102.495 ;
        RECT 87.710 102.475 87.880 102.665 ;
        RECT 88.175 102.475 88.345 102.685 ;
        RECT 91.395 102.475 91.565 102.665 ;
        RECT 91.865 102.530 92.025 102.640 ;
        RECT 95.995 102.495 96.165 102.715 ;
        RECT 96.315 102.685 101.825 103.495 ;
        RECT 101.835 102.685 105.505 103.495 ;
        RECT 105.515 102.685 106.885 103.495 ;
        RECT 96.455 102.495 96.625 102.685 ;
        RECT 96.920 102.475 97.090 102.665 ;
        RECT 101.975 102.495 102.145 102.685 ;
        RECT 103.815 102.475 103.985 102.665 ;
        RECT 104.275 102.475 104.445 102.665 ;
        RECT 105.655 102.495 105.825 102.685 ;
        RECT 106.115 102.475 106.285 102.665 ;
        RECT 106.895 102.645 107.785 103.595 ;
        RECT 109.185 103.365 110.105 103.595 ;
        RECT 107.815 102.685 110.105 103.365 ;
        RECT 110.135 102.685 111.485 103.595 ;
        RECT 111.955 102.685 113.325 103.465 ;
        RECT 114.670 103.395 115.625 103.595 ;
        RECT 113.345 102.715 115.625 103.395 ;
        RECT 107.495 102.495 107.665 102.645 ;
        RECT 107.955 102.495 108.125 102.685 ;
        RECT 109.335 102.475 109.505 102.665 ;
        RECT 111.170 102.495 111.340 102.685 ;
        RECT 111.635 102.635 111.805 102.665 ;
        RECT 111.630 102.525 111.805 102.635 ;
        RECT 111.635 102.475 111.805 102.525 ;
        RECT 112.105 102.495 112.275 102.685 ;
        RECT 113.470 102.495 113.640 102.715 ;
        RECT 114.670 102.685 115.625 102.715 ;
        RECT 116.175 102.685 118.385 103.595 ;
        RECT 118.405 102.770 118.835 103.555 ;
        RECT 118.865 102.685 120.215 103.595 ;
        RECT 120.315 102.685 123.900 103.595 ;
        RECT 123.915 102.685 125.285 103.495 ;
        RECT 113.945 102.520 114.105 102.630 ;
        RECT 114.855 102.475 115.025 102.665 ;
        RECT 115.770 102.525 115.890 102.635 ;
        RECT 118.070 102.495 118.240 102.685 ;
        RECT 118.995 102.495 119.165 102.685 ;
        RECT 123.590 102.495 123.760 102.685 ;
        RECT 124.975 102.475 125.145 102.685 ;
        RECT 53.995 101.665 55.365 102.475 ;
        RECT 55.375 101.795 57.205 102.475 ;
        RECT 57.215 101.795 59.045 102.475 ;
        RECT 55.375 101.565 56.720 101.795 ;
        RECT 59.055 101.695 60.425 102.475 ;
        RECT 60.435 101.665 65.945 102.475 ;
        RECT 66.425 101.565 67.775 102.475 ;
        RECT 67.965 101.655 70.535 102.475 ;
        RECT 68.945 101.565 70.535 101.655 ;
        RECT 70.555 101.795 74.455 102.475 ;
        RECT 70.555 101.565 71.485 101.795 ;
        RECT 74.695 101.665 76.525 102.475 ;
        RECT 76.680 101.795 78.515 102.475 ;
        RECT 77.585 101.565 78.515 101.795 ;
        RECT 79.765 101.605 80.195 102.390 ;
        RECT 80.540 101.565 84.195 102.475 ;
        RECT 84.355 101.565 88.025 102.475 ;
        RECT 88.035 101.565 91.245 102.475 ;
        RECT 91.255 101.665 96.765 102.475 ;
        RECT 96.775 101.565 101.165 102.475 ;
        RECT 101.385 101.565 104.115 102.475 ;
        RECT 104.135 101.665 105.505 102.475 ;
        RECT 105.525 101.605 105.955 102.390 ;
        RECT 105.975 101.565 109.185 102.475 ;
        RECT 109.195 101.795 111.485 102.475 ;
        RECT 111.495 101.795 113.785 102.475 ;
        RECT 114.715 101.795 123.820 102.475 ;
        RECT 110.565 101.565 111.485 101.795 ;
        RECT 112.865 101.565 113.785 101.795 ;
        RECT 123.915 101.665 125.285 102.475 ;
      LAYER nwell ;
        RECT 53.800 98.445 125.480 101.275 ;
      LAYER pwell ;
        RECT 53.995 97.245 55.365 98.055 ;
        RECT 56.295 97.245 58.125 98.155 ;
        RECT 59.980 97.925 61.345 98.155 ;
        RECT 58.135 97.245 61.345 97.925 ;
        RECT 61.355 97.245 63.185 98.155 ;
        RECT 63.195 97.245 66.865 98.055 ;
        RECT 66.885 97.330 67.315 98.115 ;
        RECT 67.335 97.925 68.680 98.155 ;
        RECT 74.915 98.065 75.865 98.155 ;
        RECT 67.335 97.245 69.165 97.925 ;
        RECT 69.175 97.245 72.845 98.055 ;
        RECT 73.935 97.245 75.865 98.065 ;
        RECT 76.075 97.245 81.585 98.055 ;
        RECT 81.595 97.245 83.425 98.055 ;
        RECT 83.435 97.245 86.185 98.155 ;
        RECT 86.195 97.245 88.025 98.055 ;
        RECT 89.880 97.925 91.245 98.155 ;
        RECT 88.035 97.245 91.245 97.925 ;
        RECT 91.255 97.245 92.625 98.055 ;
        RECT 92.645 97.330 93.075 98.115 ;
        RECT 93.525 97.245 96.305 98.155 ;
        RECT 96.315 97.245 98.145 98.055 ;
        RECT 98.615 97.245 100.430 98.155 ;
        RECT 102.720 97.955 103.665 98.155 ;
        RECT 100.915 97.275 103.665 97.955 ;
        RECT 54.135 97.035 54.305 97.245 ;
        RECT 55.490 97.200 55.660 97.225 ;
        RECT 55.490 97.090 55.685 97.200 ;
        RECT 55.490 97.055 55.660 97.090 ;
        RECT 56.440 97.055 56.610 97.245 ;
        RECT 58.280 97.055 58.450 97.245 ;
        RECT 60.125 97.080 60.285 97.190 ;
        RECT 55.550 97.035 55.660 97.055 ;
        RECT 61.035 97.035 61.205 97.225 ;
        RECT 62.870 97.055 63.040 97.245 ;
        RECT 63.335 97.055 63.505 97.245 ;
        RECT 64.715 97.035 64.885 97.225 ;
        RECT 68.855 97.055 69.025 97.245 ;
        RECT 69.315 97.035 69.485 97.245 ;
        RECT 73.935 97.225 74.085 97.245 ;
        RECT 73.005 97.090 73.165 97.200 ;
        RECT 73.915 97.055 74.085 97.225 ;
        RECT 75.295 97.035 75.465 97.225 ;
        RECT 75.755 97.035 75.925 97.225 ;
        RECT 76.215 97.055 76.385 97.245 ;
        RECT 79.430 97.085 79.550 97.195 ;
        RECT 80.345 97.035 80.515 97.225 ;
        RECT 81.735 97.055 81.905 97.245 ;
        RECT 83.575 97.035 83.745 97.245 ;
        RECT 86.335 97.035 86.505 97.245 ;
        RECT 88.180 97.055 88.350 97.245 ;
        RECT 89.090 97.035 89.260 97.225 ;
        RECT 89.555 97.035 89.725 97.225 ;
        RECT 91.395 97.055 91.565 97.245 ;
        RECT 95.075 97.035 95.245 97.225 ;
        RECT 95.995 97.055 96.165 97.245 ;
        RECT 96.455 97.055 96.625 97.245 ;
        RECT 98.290 97.085 98.410 97.195 ;
        RECT 98.755 97.035 98.925 97.225 ;
        RECT 100.135 97.055 100.305 97.245 ;
        RECT 101.060 97.225 101.230 97.275 ;
        RECT 102.720 97.245 103.665 97.275 ;
        RECT 103.675 97.245 106.425 98.055 ;
        RECT 108.265 97.925 109.185 98.155 ;
        RECT 106.895 97.245 109.185 97.925 ;
        RECT 109.215 97.245 110.565 98.155 ;
        RECT 110.575 97.245 114.245 98.055 ;
        RECT 115.175 97.245 116.545 98.025 ;
        RECT 116.555 97.245 118.385 97.925 ;
        RECT 118.405 97.330 118.835 98.115 ;
        RECT 119.800 97.925 121.140 98.155 ;
        RECT 119.315 97.245 123.905 97.925 ;
        RECT 123.915 97.245 125.285 98.055 ;
        RECT 100.590 97.085 100.710 97.195 ;
        RECT 101.055 97.055 101.230 97.225 ;
        RECT 101.055 97.035 101.225 97.055 ;
        RECT 101.515 97.035 101.685 97.225 ;
        RECT 103.815 97.055 103.985 97.245 ;
        RECT 105.190 97.085 105.310 97.195 ;
        RECT 106.570 97.085 106.690 97.195 ;
        RECT 107.035 97.055 107.205 97.245 ;
        RECT 108.415 97.035 108.585 97.225 ;
        RECT 110.250 97.055 110.420 97.245 ;
        RECT 110.715 97.055 110.885 97.245 ;
        RECT 110.715 97.035 110.865 97.055 ;
        RECT 111.175 97.035 111.345 97.225 ;
        RECT 114.405 97.090 114.565 97.200 ;
        RECT 115.325 97.055 115.495 97.245 ;
        RECT 116.705 97.080 116.865 97.190 ;
        RECT 118.075 97.055 118.245 97.245 ;
        RECT 118.525 97.035 118.695 97.225 ;
        RECT 119.005 97.195 119.175 97.225 ;
        RECT 118.990 97.085 119.175 97.195 ;
        RECT 119.005 97.035 119.175 97.085 ;
        RECT 119.460 97.055 119.630 97.245 ;
        RECT 121.755 97.035 121.925 97.225 ;
        RECT 122.215 97.035 122.385 97.225 ;
        RECT 124.975 97.035 125.145 97.245 ;
        RECT 53.995 96.225 55.365 97.035 ;
        RECT 55.550 96.355 59.965 97.035 ;
        RECT 60.895 96.355 64.565 97.035 ;
        RECT 64.575 96.805 66.145 97.035 ;
        RECT 68.235 96.995 69.155 97.035 ;
        RECT 68.235 96.805 69.165 96.995 ;
        RECT 64.575 96.445 69.165 96.805 ;
        RECT 64.575 96.355 69.155 96.445 ;
        RECT 56.035 96.125 59.965 96.355 ;
        RECT 63.635 96.125 64.565 96.355 ;
        RECT 66.155 96.125 69.155 96.355 ;
        RECT 69.175 96.225 71.925 97.035 ;
        RECT 72.075 96.125 75.525 97.035 ;
        RECT 75.615 96.225 79.285 97.035 ;
        RECT 79.765 96.165 80.195 96.950 ;
        RECT 80.215 96.125 83.425 97.035 ;
        RECT 83.445 96.125 86.175 97.035 ;
        RECT 86.195 96.225 88.025 97.035 ;
        RECT 88.055 96.125 89.405 97.035 ;
        RECT 89.415 96.225 94.925 97.035 ;
        RECT 94.935 96.225 98.605 97.035 ;
        RECT 98.615 96.225 99.985 97.035 ;
        RECT 100.005 96.125 101.355 97.035 ;
        RECT 101.375 96.225 105.045 97.035 ;
        RECT 105.525 96.165 105.955 96.950 ;
        RECT 105.985 96.125 108.715 97.035 ;
        RECT 108.935 96.215 110.865 97.035 ;
        RECT 111.035 96.225 116.545 97.035 ;
        RECT 117.475 96.255 118.845 97.035 ;
        RECT 118.855 96.255 120.225 97.035 ;
        RECT 120.235 96.355 122.065 97.035 ;
        RECT 122.075 96.355 123.905 97.035 ;
        RECT 108.935 96.125 109.885 96.215 ;
        RECT 120.235 96.125 121.580 96.355 ;
        RECT 122.560 96.125 123.905 96.355 ;
        RECT 123.915 96.225 125.285 97.035 ;
      LAYER nwell ;
        RECT 53.800 93.005 125.480 95.835 ;
      LAYER pwell ;
        RECT 55.385 92.625 56.975 92.715 ;
        RECT 53.995 91.805 55.365 92.615 ;
        RECT 55.385 91.805 57.955 92.625 ;
        RECT 59.955 92.485 60.885 92.715 ;
        RECT 58.135 91.805 60.885 92.485 ;
        RECT 60.895 91.805 62.725 92.615 ;
        RECT 63.195 92.515 64.125 92.715 ;
        RECT 65.455 92.515 66.405 92.715 ;
        RECT 63.195 92.035 66.405 92.515 ;
        RECT 63.340 91.835 66.405 92.035 ;
        RECT 66.885 91.890 67.315 92.675 ;
        RECT 67.335 92.515 68.265 92.715 ;
        RECT 69.595 92.515 70.545 92.715 ;
        RECT 67.335 92.035 70.545 92.515 ;
        RECT 54.135 91.595 54.305 91.805 ;
        RECT 57.815 91.785 57.955 91.805 ;
        RECT 56.895 91.595 57.065 91.785 ;
        RECT 57.355 91.595 57.525 91.785 ;
        RECT 57.815 91.615 57.985 91.785 ;
        RECT 58.275 91.615 58.445 91.805 ;
        RECT 59.655 91.595 59.825 91.785 ;
        RECT 60.115 91.595 60.285 91.785 ;
        RECT 61.035 91.615 61.205 91.805 ;
        RECT 62.870 91.645 62.990 91.755 ;
        RECT 63.340 91.615 63.510 91.835 ;
        RECT 65.470 91.805 66.405 91.835 ;
        RECT 67.480 91.835 70.545 92.035 ;
        RECT 65.635 91.595 65.805 91.785 ;
        RECT 66.550 91.645 66.670 91.755 ;
        RECT 67.480 91.615 67.650 91.835 ;
        RECT 69.610 91.805 70.545 91.835 ;
        RECT 71.485 91.805 75.605 92.715 ;
        RECT 75.615 91.805 77.445 92.485 ;
        RECT 77.475 91.805 78.825 92.715 ;
        RECT 80.435 92.625 81.385 92.715 ;
        RECT 79.455 91.805 81.385 92.625 ;
        RECT 81.595 92.035 83.430 92.715 ;
        RECT 81.740 91.805 83.430 92.035 ;
        RECT 83.895 91.805 85.725 92.615 ;
        RECT 86.195 91.805 89.865 92.715 ;
        RECT 90.360 92.485 91.705 92.715 ;
        RECT 89.875 91.805 91.705 92.485 ;
        RECT 92.645 91.890 93.075 92.675 ;
        RECT 93.095 91.805 96.305 92.715 ;
        RECT 96.355 92.485 97.730 92.715 ;
        RECT 99.520 92.485 100.900 92.715 ;
        RECT 96.355 92.035 100.900 92.485 ;
        RECT 70.705 91.650 70.865 91.760 ;
        RECT 71.155 91.595 71.325 91.785 ;
        RECT 72.995 91.595 73.165 91.785 ;
        RECT 73.455 91.615 73.625 91.805 ;
        RECT 74.835 91.595 75.005 91.785 ;
        RECT 75.295 91.615 75.465 91.805 ;
        RECT 77.135 91.615 77.305 91.805 ;
        RECT 78.510 91.785 78.680 91.805 ;
        RECT 79.455 91.785 79.605 91.805 ;
        RECT 78.510 91.615 78.685 91.785 ;
        RECT 78.970 91.645 79.090 91.755 ;
        RECT 79.435 91.615 79.605 91.785 ;
        RECT 78.515 91.595 78.685 91.615 ;
        RECT 80.355 91.595 80.525 91.785 ;
        RECT 81.740 91.615 81.910 91.805 ;
        RECT 84.035 91.615 84.205 91.805 ;
        RECT 85.870 91.645 85.990 91.755 ;
        RECT 86.335 91.595 86.505 91.805 ;
        RECT 90.015 91.615 90.185 91.805 ;
        RECT 91.855 91.615 92.025 91.785 ;
        RECT 91.855 91.595 92.020 91.615 ;
        RECT 92.320 91.595 92.490 91.785 ;
        RECT 93.235 91.615 93.405 91.805 ;
        RECT 93.695 91.595 93.865 91.785 ;
        RECT 96.460 91.615 96.630 92.035 ;
        RECT 97.740 91.805 100.900 92.035 ;
        RECT 100.915 91.805 102.265 92.715 ;
        RECT 102.295 91.805 103.665 92.615 ;
        RECT 103.685 91.805 106.415 92.715 ;
        RECT 106.435 91.805 108.250 92.715 ;
        RECT 108.275 91.805 113.785 92.615 ;
        RECT 113.795 91.805 117.465 92.615 ;
        RECT 118.405 91.890 118.835 92.675 ;
        RECT 118.855 91.805 120.685 92.615 ;
        RECT 120.695 91.805 122.065 92.585 ;
        RECT 122.075 91.805 123.905 92.485 ;
        RECT 123.915 91.805 125.285 92.615 ;
        RECT 96.910 91.595 97.080 91.785 ;
        RECT 98.295 91.595 98.465 91.785 ;
        RECT 101.980 91.615 102.150 91.805 ;
        RECT 102.435 91.615 102.605 91.805 ;
        RECT 105.195 91.595 105.365 91.785 ;
        RECT 106.115 91.595 106.285 91.805 ;
        RECT 107.955 91.615 108.125 91.805 ;
        RECT 108.415 91.615 108.585 91.805 ;
        RECT 111.635 91.595 111.805 91.785 ;
        RECT 113.935 91.615 114.105 91.805 ;
        RECT 117.155 91.595 117.325 91.785 ;
        RECT 117.625 91.650 117.785 91.760 ;
        RECT 118.995 91.615 119.165 91.805 ;
        RECT 120.845 91.615 121.015 91.805 ;
        RECT 122.215 91.615 122.385 91.805 ;
        RECT 123.595 91.595 123.765 91.785 ;
        RECT 124.975 91.595 125.145 91.805 ;
        RECT 53.995 90.785 55.365 91.595 ;
        RECT 55.375 90.915 57.205 91.595 ;
        RECT 55.375 90.685 56.720 90.915 ;
        RECT 57.225 90.685 58.575 91.595 ;
        RECT 58.595 90.815 59.965 91.595 ;
        RECT 59.975 90.785 65.485 91.595 ;
        RECT 65.495 90.785 71.005 91.595 ;
        RECT 71.030 90.685 72.845 91.595 ;
        RECT 72.855 90.915 74.685 91.595 ;
        RECT 73.340 90.685 74.685 90.915 ;
        RECT 74.695 90.785 78.365 91.595 ;
        RECT 78.375 90.785 79.745 91.595 ;
        RECT 79.765 90.725 80.195 91.510 ;
        RECT 80.215 90.785 85.725 91.595 ;
        RECT 86.195 90.685 89.865 91.595 ;
        RECT 90.185 90.915 92.020 91.595 ;
        RECT 90.185 90.685 91.115 90.915 ;
        RECT 92.175 90.685 93.525 91.595 ;
        RECT 93.555 90.685 96.765 91.595 ;
        RECT 96.795 90.685 98.145 91.595 ;
        RECT 98.155 90.785 103.665 91.595 ;
        RECT 103.675 90.685 105.490 91.595 ;
        RECT 105.525 90.725 105.955 91.510 ;
        RECT 105.975 90.785 111.485 91.595 ;
        RECT 111.495 90.785 117.005 91.595 ;
        RECT 117.015 90.785 122.525 91.595 ;
        RECT 122.535 90.815 123.905 91.595 ;
        RECT 123.915 90.785 125.285 91.595 ;
      LAYER nwell ;
        RECT 53.800 87.565 125.480 90.395 ;
      LAYER pwell ;
        RECT 53.995 86.365 55.365 87.175 ;
        RECT 55.375 86.365 60.885 87.175 ;
        RECT 60.895 86.365 66.405 87.175 ;
        RECT 66.885 86.450 67.315 87.235 ;
        RECT 67.335 86.365 69.165 87.175 ;
        RECT 69.655 86.365 71.005 87.275 ;
        RECT 71.015 86.365 74.675 87.275 ;
        RECT 74.865 86.365 78.365 87.275 ;
        RECT 78.375 86.365 81.125 87.175 ;
        RECT 81.145 86.595 84.345 87.275 ;
        RECT 81.145 86.365 84.200 86.595 ;
        RECT 84.355 86.365 89.865 87.175 ;
        RECT 89.875 86.365 92.625 87.175 ;
        RECT 92.645 86.450 93.075 87.235 ;
        RECT 93.590 87.045 94.965 87.275 ;
        RECT 96.735 87.045 97.685 87.275 ;
        RECT 98.180 87.045 99.525 87.275 ;
        RECT 100.020 87.045 103.630 87.275 ;
        RECT 93.590 86.595 97.685 87.045 ;
        RECT 54.135 86.155 54.305 86.365 ;
        RECT 55.515 86.155 55.685 86.365 ;
        RECT 61.035 86.155 61.205 86.365 ;
        RECT 66.555 86.315 66.725 86.345 ;
        RECT 66.550 86.205 66.725 86.315 ;
        RECT 66.555 86.155 66.725 86.205 ;
        RECT 67.475 86.175 67.645 86.365 ;
        RECT 69.310 86.205 69.430 86.315 ;
        RECT 69.770 86.175 69.940 86.365 ;
        RECT 73.450 86.155 73.620 86.345 ;
        RECT 74.390 86.175 74.560 86.365 ;
        RECT 74.865 86.345 75.000 86.365 ;
        RECT 74.830 86.175 75.000 86.345 ;
        RECT 75.755 86.175 75.925 86.345 ;
        RECT 76.225 86.200 76.385 86.310 ;
        RECT 75.755 86.155 75.905 86.175 ;
        RECT 77.140 86.155 77.310 86.345 ;
        RECT 78.515 86.175 78.685 86.365 ;
        RECT 79.430 86.205 79.550 86.315 ;
        RECT 81.735 86.155 81.905 86.345 ;
        RECT 82.195 86.155 82.365 86.345 ;
        RECT 83.575 86.155 83.745 86.345 ;
        RECT 84.030 86.175 84.200 86.365 ;
        RECT 84.495 86.175 84.665 86.365 ;
        RECT 89.095 86.155 89.265 86.345 ;
        RECT 90.015 86.175 90.185 86.365 ;
        RECT 93.230 86.205 93.350 86.315 ;
        RECT 93.695 86.175 93.865 86.595 ;
        RECT 94.975 86.365 97.685 86.595 ;
        RECT 97.695 86.365 99.525 87.045 ;
        RECT 99.535 86.365 103.630 87.045 ;
        RECT 103.675 86.365 109.185 87.175 ;
        RECT 109.195 86.365 114.705 87.175 ;
        RECT 114.715 86.365 118.385 87.175 ;
        RECT 118.405 86.450 118.835 87.235 ;
        RECT 118.855 86.365 121.605 87.175 ;
        RECT 122.075 86.365 123.905 87.045 ;
        RECT 123.915 86.365 125.285 87.175 ;
        RECT 94.615 86.155 94.785 86.345 ;
        RECT 97.835 86.175 98.005 86.365 ;
        RECT 98.290 86.205 98.410 86.315 ;
        RECT 99.680 86.175 99.850 86.365 ;
        RECT 102.430 86.155 102.600 86.345 ;
        RECT 102.895 86.155 103.065 86.345 ;
        RECT 103.815 86.175 103.985 86.365 ;
        RECT 106.115 86.155 106.285 86.345 ;
        RECT 109.335 86.175 109.505 86.365 ;
        RECT 111.635 86.155 111.805 86.345 ;
        RECT 114.855 86.175 115.025 86.365 ;
        RECT 117.155 86.155 117.325 86.345 ;
        RECT 118.995 86.175 119.165 86.365 ;
        RECT 121.750 86.205 121.870 86.315 ;
        RECT 123.595 86.175 123.765 86.365 ;
        RECT 124.975 86.155 125.145 86.365 ;
        RECT 53.995 85.345 55.365 86.155 ;
        RECT 55.375 85.345 60.885 86.155 ;
        RECT 60.895 85.345 66.405 86.155 ;
        RECT 66.415 85.345 71.925 86.155 ;
        RECT 71.935 85.245 73.765 86.155 ;
        RECT 73.975 85.335 75.905 86.155 ;
        RECT 76.995 85.475 79.270 86.155 ;
        RECT 73.975 85.245 74.925 85.335 ;
        RECT 77.900 85.245 79.270 85.475 ;
        RECT 79.765 85.285 80.195 86.070 ;
        RECT 80.215 85.475 82.045 86.155 ;
        RECT 82.055 85.375 83.425 86.155 ;
        RECT 83.435 85.345 88.945 86.155 ;
        RECT 88.955 85.345 94.465 86.155 ;
        RECT 94.475 85.345 98.145 86.155 ;
        RECT 98.650 85.475 102.745 86.155 ;
        RECT 98.650 85.245 102.260 85.475 ;
        RECT 102.755 85.345 105.505 86.155 ;
        RECT 105.525 85.285 105.955 86.070 ;
        RECT 105.975 85.345 111.485 86.155 ;
        RECT 111.495 85.345 117.005 86.155 ;
        RECT 117.015 85.345 122.525 86.155 ;
        RECT 123.915 85.345 125.285 86.155 ;
      LAYER nwell ;
        RECT 53.800 82.125 125.480 84.955 ;
      LAYER pwell ;
        RECT 53.995 80.925 55.365 81.735 ;
        RECT 55.375 80.925 60.885 81.735 ;
        RECT 63.195 80.925 66.865 81.735 ;
        RECT 66.885 81.010 67.315 81.795 ;
        RECT 67.335 80.925 71.005 81.735 ;
        RECT 71.475 80.925 72.845 81.705 ;
        RECT 72.855 80.925 74.685 81.735 ;
        RECT 75.180 81.605 76.525 81.835 ;
        RECT 74.695 80.925 76.525 81.605 ;
        RECT 76.535 80.925 77.885 81.835 ;
        RECT 77.915 80.925 79.285 81.705 ;
        RECT 79.765 81.010 80.195 81.795 ;
        RECT 81.135 80.925 82.965 81.605 ;
        RECT 82.975 80.925 84.345 81.735 ;
        RECT 84.840 81.605 86.185 81.835 ;
        RECT 84.355 80.925 86.185 81.605 ;
        RECT 86.195 80.925 91.705 81.735 ;
        RECT 92.645 81.010 93.075 81.795 ;
        RECT 93.095 80.925 98.605 81.735 ;
        RECT 98.615 80.925 104.125 81.735 ;
        RECT 104.135 80.925 105.505 81.735 ;
        RECT 105.525 81.010 105.955 81.795 ;
        RECT 105.975 80.925 111.485 81.735 ;
        RECT 111.495 80.925 117.005 81.735 ;
        RECT 117.015 80.925 118.385 81.735 ;
        RECT 118.405 81.010 118.835 81.795 ;
        RECT 118.855 80.925 122.525 81.735 ;
        RECT 122.535 80.925 123.905 81.735 ;
        RECT 123.915 80.925 125.285 81.735 ;
        RECT 54.135 80.735 54.305 80.925 ;
        RECT 55.515 80.735 55.685 80.925 ;
        RECT 61.045 80.770 61.205 80.880 ;
        RECT 62.875 80.735 63.045 80.905 ;
        RECT 63.335 80.735 63.505 80.925 ;
        RECT 67.475 80.735 67.645 80.925 ;
        RECT 71.150 80.765 71.270 80.875 ;
        RECT 72.535 80.735 72.705 80.925 ;
        RECT 72.995 80.735 73.165 80.925 ;
        RECT 74.835 80.735 75.005 80.925 ;
        RECT 77.600 80.735 77.770 80.925 ;
        RECT 78.065 80.735 78.235 80.925 ;
        RECT 79.430 80.765 79.550 80.875 ;
        RECT 80.365 80.770 80.525 80.880 ;
        RECT 81.275 80.735 81.445 80.925 ;
        RECT 83.115 80.735 83.285 80.925 ;
        RECT 84.495 80.735 84.665 80.925 ;
        RECT 86.335 80.735 86.505 80.925 ;
        RECT 91.865 80.770 92.025 80.880 ;
        RECT 93.235 80.735 93.405 80.925 ;
        RECT 98.755 80.735 98.925 80.925 ;
        RECT 104.275 80.735 104.445 80.925 ;
        RECT 106.115 80.735 106.285 80.925 ;
        RECT 111.635 80.735 111.805 80.925 ;
        RECT 117.155 80.735 117.325 80.925 ;
        RECT 118.995 80.735 119.165 80.925 ;
        RECT 122.675 80.735 122.845 80.925 ;
        RECT 124.975 80.735 125.145 80.925 ;
      LAYER li1 ;
        RECT 53.990 151.455 125.290 151.625 ;
        RECT 54.075 150.705 55.285 151.455 ;
        RECT 54.075 150.165 54.595 150.705 ;
        RECT 55.515 150.635 55.725 151.455 ;
        RECT 55.895 150.655 56.225 151.285 ;
        RECT 54.765 149.995 55.285 150.535 ;
        RECT 55.895 150.055 56.145 150.655 ;
        RECT 56.395 150.635 56.625 151.455 ;
        RECT 56.925 150.905 57.095 151.285 ;
        RECT 57.310 151.075 57.640 151.455 ;
        RECT 56.925 150.735 57.640 150.905 ;
        RECT 56.315 150.215 56.645 150.465 ;
        RECT 56.835 150.185 57.190 150.555 ;
        RECT 57.470 150.545 57.640 150.735 ;
        RECT 57.810 150.710 58.065 151.285 ;
        RECT 57.470 150.215 57.725 150.545 ;
        RECT 54.075 148.905 55.285 149.995 ;
        RECT 55.515 148.905 55.725 150.045 ;
        RECT 55.895 149.075 56.225 150.055 ;
        RECT 56.395 148.905 56.625 150.045 ;
        RECT 57.470 150.005 57.640 150.215 ;
        RECT 56.925 149.835 57.640 150.005 ;
        RECT 57.895 149.980 58.065 150.710 ;
        RECT 58.240 150.615 58.500 151.455 ;
        RECT 58.680 150.615 58.940 151.455 ;
        RECT 59.115 150.710 59.370 151.285 ;
        RECT 59.540 151.075 59.870 151.455 ;
        RECT 60.085 150.905 60.255 151.285 ;
        RECT 59.540 150.735 60.255 150.905 ;
        RECT 56.925 149.075 57.095 149.835 ;
        RECT 57.310 148.905 57.640 149.665 ;
        RECT 57.810 149.075 58.065 149.980 ;
        RECT 58.240 148.905 58.500 150.055 ;
        RECT 58.680 148.905 58.940 150.055 ;
        RECT 59.115 149.980 59.285 150.710 ;
        RECT 59.540 150.545 59.710 150.735 ;
        RECT 60.520 150.615 60.780 151.455 ;
        RECT 60.955 150.710 61.210 151.285 ;
        RECT 61.380 151.075 61.710 151.455 ;
        RECT 61.925 150.905 62.095 151.285 ;
        RECT 62.520 150.945 62.760 151.455 ;
        RECT 62.940 150.945 63.220 151.275 ;
        RECT 63.450 150.945 63.665 151.455 ;
        RECT 61.380 150.735 62.095 150.905 ;
        RECT 59.455 150.215 59.710 150.545 ;
        RECT 59.540 150.005 59.710 150.215 ;
        RECT 59.990 150.185 60.345 150.555 ;
        RECT 59.115 149.075 59.370 149.980 ;
        RECT 59.540 149.835 60.255 150.005 ;
        RECT 59.540 148.905 59.870 149.665 ;
        RECT 60.085 149.075 60.255 149.835 ;
        RECT 60.520 148.905 60.780 150.055 ;
        RECT 60.955 149.980 61.125 150.710 ;
        RECT 61.380 150.545 61.550 150.735 ;
        RECT 61.295 150.215 61.550 150.545 ;
        RECT 61.380 150.005 61.550 150.215 ;
        RECT 61.830 150.185 62.185 150.555 ;
        RECT 62.415 150.215 62.770 150.775 ;
        RECT 62.940 150.045 63.110 150.945 ;
        RECT 63.280 150.215 63.545 150.775 ;
        RECT 63.835 150.715 64.450 151.285 ;
        RECT 64.765 151.075 65.935 151.285 ;
        RECT 64.765 151.055 65.095 151.075 ;
        RECT 63.795 150.045 63.965 150.545 ;
        RECT 60.955 149.075 61.210 149.980 ;
        RECT 61.380 149.835 62.095 150.005 ;
        RECT 61.380 148.905 61.710 149.665 ;
        RECT 61.925 149.075 62.095 149.835 ;
        RECT 62.540 149.875 63.965 150.045 ;
        RECT 62.540 149.700 62.930 149.875 ;
        RECT 63.415 148.905 63.745 149.705 ;
        RECT 64.135 149.695 64.450 150.715 ;
        RECT 64.655 150.635 65.515 150.885 ;
        RECT 65.685 150.825 65.935 151.075 ;
        RECT 66.105 150.995 66.275 151.455 ;
        RECT 66.445 150.825 66.785 151.285 ;
        RECT 65.685 150.655 66.785 150.825 ;
        RECT 66.955 150.730 67.245 151.455 ;
        RECT 67.525 151.075 68.695 151.285 ;
        RECT 67.525 151.055 67.855 151.075 ;
        RECT 67.415 150.635 68.275 150.885 ;
        RECT 68.445 150.825 68.695 151.075 ;
        RECT 68.865 150.995 69.035 151.455 ;
        RECT 69.205 150.825 69.545 151.285 ;
        RECT 68.445 150.655 69.545 150.825 ;
        RECT 69.915 150.825 70.245 151.185 ;
        RECT 70.875 150.995 71.125 151.455 ;
        RECT 71.295 150.995 71.845 151.285 ;
        RECT 69.915 150.635 71.305 150.825 ;
        RECT 64.655 150.045 64.935 150.635 ;
        RECT 65.105 150.215 65.855 150.465 ;
        RECT 66.025 150.215 66.785 150.465 ;
        RECT 64.655 149.875 66.355 150.045 ;
        RECT 63.915 149.075 64.450 149.695 ;
        RECT 64.760 148.905 65.015 149.705 ;
        RECT 65.185 149.075 65.515 149.875 ;
        RECT 65.685 148.905 65.855 149.705 ;
        RECT 66.025 149.075 66.355 149.875 ;
        RECT 66.525 148.905 66.785 150.045 ;
        RECT 66.955 148.905 67.245 150.070 ;
        RECT 67.415 150.045 67.695 150.635 ;
        RECT 71.135 150.545 71.305 150.635 ;
        RECT 67.865 150.215 68.615 150.465 ;
        RECT 68.785 150.215 69.545 150.465 ;
        RECT 69.715 150.215 70.405 150.465 ;
        RECT 70.635 150.215 70.965 150.465 ;
        RECT 71.135 150.215 71.425 150.545 ;
        RECT 67.415 149.875 69.115 150.045 ;
        RECT 67.520 148.905 67.775 149.705 ;
        RECT 67.945 149.075 68.275 149.875 ;
        RECT 68.445 148.905 68.615 149.705 ;
        RECT 68.785 149.075 69.115 149.875 ;
        RECT 69.285 148.905 69.545 150.045 ;
        RECT 69.715 149.775 70.030 150.215 ;
        RECT 71.135 149.965 71.305 150.215 ;
        RECT 70.365 149.795 71.305 149.965 ;
        RECT 69.915 148.905 70.195 149.575 ;
        RECT 70.365 149.245 70.665 149.795 ;
        RECT 71.595 149.625 71.845 150.995 ;
        RECT 72.015 150.655 72.305 151.455 ;
        RECT 72.560 150.955 73.055 151.285 ;
        RECT 70.875 148.905 71.205 149.625 ;
        RECT 71.395 149.075 71.845 149.625 ;
        RECT 72.015 148.905 72.305 150.045 ;
        RECT 72.475 149.465 72.715 150.775 ;
        RECT 72.885 150.045 73.055 150.955 ;
        RECT 73.275 150.215 73.625 151.180 ;
        RECT 73.805 150.215 74.105 151.185 ;
        RECT 74.285 150.215 74.565 151.185 ;
        RECT 74.745 150.655 75.015 151.455 ;
        RECT 75.185 150.735 75.525 151.245 ;
        RECT 75.780 150.905 76.110 151.285 ;
        RECT 76.280 151.075 77.465 151.245 ;
        RECT 77.725 150.985 77.895 151.455 ;
        RECT 75.780 150.735 76.325 150.905 ;
        RECT 74.760 150.215 75.090 150.465 ;
        RECT 74.760 150.045 75.075 150.215 ;
        RECT 72.885 149.875 75.075 150.045 ;
        RECT 72.480 148.905 72.815 149.285 ;
        RECT 72.985 149.075 73.235 149.875 ;
        RECT 73.455 148.905 73.785 149.625 ;
        RECT 73.970 149.075 74.220 149.875 ;
        RECT 74.685 148.905 75.015 149.705 ;
        RECT 75.265 149.335 75.525 150.735 ;
        RECT 75.695 150.215 75.955 150.565 ;
        RECT 76.155 150.095 76.325 150.735 ;
        RECT 76.695 150.805 77.080 150.895 ;
        RECT 78.065 150.805 78.395 151.270 ;
        RECT 76.695 150.635 78.395 150.805 ;
        RECT 78.565 150.635 78.735 151.455 ;
        RECT 78.905 150.805 79.235 151.275 ;
        RECT 79.405 150.975 79.575 151.455 ;
        RECT 78.905 150.635 79.665 150.805 ;
        RECT 79.835 150.730 80.125 151.455 ;
        RECT 81.305 150.975 81.605 151.455 ;
        RECT 81.775 150.805 82.035 151.260 ;
        RECT 82.205 150.975 82.465 151.455 ;
        RECT 82.645 150.805 82.905 151.260 ;
        RECT 83.075 150.975 83.325 151.455 ;
        RECT 83.505 150.805 83.765 151.260 ;
        RECT 83.935 150.975 84.185 151.455 ;
        RECT 84.365 150.805 84.625 151.260 ;
        RECT 84.795 150.975 85.040 151.455 ;
        RECT 85.210 150.805 85.485 151.260 ;
        RECT 85.655 150.975 85.900 151.455 ;
        RECT 86.070 150.805 86.330 151.260 ;
        RECT 86.500 150.975 86.760 151.455 ;
        RECT 86.930 150.805 87.190 151.260 ;
        RECT 87.360 150.975 87.620 151.455 ;
        RECT 87.790 150.805 88.050 151.260 ;
        RECT 88.220 150.895 88.480 151.455 ;
        RECT 81.305 150.775 88.050 150.805 ;
        RECT 76.495 150.265 76.840 150.465 ;
        RECT 77.010 150.265 77.400 150.465 ;
        RECT 76.155 150.045 76.940 150.095 ;
        RECT 75.185 149.075 75.525 149.335 ;
        RECT 75.860 149.870 76.940 150.045 ;
        RECT 75.860 149.075 76.190 149.870 ;
        RECT 76.360 148.905 76.600 149.690 ;
        RECT 76.770 149.665 76.940 149.870 ;
        RECT 77.110 149.835 77.400 150.265 ;
        RECT 77.590 150.255 78.075 150.465 ;
        RECT 78.245 150.255 78.685 150.465 ;
        RECT 78.855 150.255 79.185 150.465 ;
        RECT 77.590 149.835 77.895 150.255 ;
        RECT 78.855 150.085 79.025 150.255 ;
        RECT 78.065 149.915 79.025 150.085 ;
        RECT 78.065 149.665 78.235 149.915 ;
        RECT 76.770 149.495 78.235 149.665 ;
        RECT 77.160 149.075 77.915 149.495 ;
        RECT 78.405 148.905 78.735 149.745 ;
        RECT 79.355 149.665 79.665 150.635 ;
        RECT 81.275 150.635 88.050 150.775 ;
        RECT 81.275 150.605 82.470 150.635 ;
        RECT 78.905 149.495 79.665 149.665 ;
        RECT 78.905 149.075 79.155 149.495 ;
        RECT 79.325 148.905 79.665 149.325 ;
        RECT 79.835 148.905 80.125 150.070 ;
        RECT 81.305 150.045 82.470 150.605 ;
        RECT 88.650 150.465 88.900 151.275 ;
        RECT 89.080 150.930 89.340 151.455 ;
        RECT 89.510 150.465 89.760 151.275 ;
        RECT 89.940 150.945 90.245 151.455 ;
        RECT 90.435 150.945 90.675 151.455 ;
        RECT 90.845 150.945 91.135 151.285 ;
        RECT 91.365 150.945 91.680 151.455 ;
        RECT 82.640 150.215 89.760 150.465 ;
        RECT 89.930 150.215 90.245 150.775 ;
        RECT 90.480 150.435 90.675 150.775 ;
        RECT 90.475 150.265 90.675 150.435 ;
        RECT 90.480 150.215 90.675 150.265 ;
        RECT 81.305 149.820 88.050 150.045 ;
        RECT 81.305 148.905 81.575 149.650 ;
        RECT 81.745 149.080 82.035 149.820 ;
        RECT 82.645 149.805 88.050 149.820 ;
        RECT 82.205 148.910 82.460 149.635 ;
        RECT 82.645 149.080 82.905 149.805 ;
        RECT 83.075 148.910 83.320 149.635 ;
        RECT 83.505 149.080 83.765 149.805 ;
        RECT 83.935 148.910 84.180 149.635 ;
        RECT 84.365 149.080 84.625 149.805 ;
        RECT 84.795 148.910 85.040 149.635 ;
        RECT 85.210 149.080 85.470 149.805 ;
        RECT 85.640 148.910 85.900 149.635 ;
        RECT 86.070 149.080 86.330 149.805 ;
        RECT 86.500 148.910 86.760 149.635 ;
        RECT 86.930 149.080 87.190 149.805 ;
        RECT 87.360 148.910 87.620 149.635 ;
        RECT 87.790 149.080 88.050 149.805 ;
        RECT 88.220 148.910 88.480 149.705 ;
        RECT 88.650 149.080 88.900 150.215 ;
        RECT 82.205 148.905 88.480 148.910 ;
        RECT 89.080 148.905 89.340 149.715 ;
        RECT 89.515 149.075 89.760 150.215 ;
        RECT 90.845 150.045 91.025 150.945 ;
        RECT 91.850 150.885 92.020 151.155 ;
        RECT 92.190 151.055 92.520 151.455 ;
        RECT 91.195 150.215 91.605 150.775 ;
        RECT 91.850 150.715 92.545 150.885 ;
        RECT 92.715 150.730 93.005 151.455 ;
        RECT 93.505 151.055 93.835 151.455 ;
        RECT 94.005 150.885 94.335 151.225 ;
        RECT 95.385 151.055 95.715 151.455 ;
        RECT 91.775 150.045 91.945 150.545 ;
        RECT 90.485 149.875 91.945 150.045 ;
        RECT 89.940 148.905 90.235 149.715 ;
        RECT 90.485 149.700 90.845 149.875 ;
        RECT 92.115 149.705 92.545 150.715 ;
        RECT 93.350 150.715 95.715 150.885 ;
        RECT 95.885 150.730 96.215 151.240 ;
        RECT 96.485 150.975 96.785 151.455 ;
        RECT 96.955 150.805 97.215 151.260 ;
        RECT 97.385 150.975 97.645 151.455 ;
        RECT 97.825 150.805 98.085 151.260 ;
        RECT 98.255 150.975 98.505 151.455 ;
        RECT 98.685 150.805 98.945 151.260 ;
        RECT 99.115 150.975 99.365 151.455 ;
        RECT 99.545 150.805 99.805 151.260 ;
        RECT 99.975 150.975 100.220 151.455 ;
        RECT 100.390 150.805 100.665 151.260 ;
        RECT 100.835 150.975 101.080 151.455 ;
        RECT 101.250 150.805 101.510 151.260 ;
        RECT 101.680 150.975 101.940 151.455 ;
        RECT 102.110 150.805 102.370 151.260 ;
        RECT 102.540 150.975 102.800 151.455 ;
        RECT 102.970 150.805 103.230 151.260 ;
        RECT 103.400 150.895 103.660 151.455 ;
        RECT 91.430 148.905 91.600 149.705 ;
        RECT 91.770 149.535 92.545 149.705 ;
        RECT 91.770 149.075 92.100 149.535 ;
        RECT 92.270 148.905 92.440 149.365 ;
        RECT 92.715 148.905 93.005 150.070 ;
        RECT 93.350 149.715 93.520 150.715 ;
        RECT 95.545 150.545 95.715 150.715 ;
        RECT 93.690 149.885 93.935 150.545 ;
        RECT 94.150 149.885 94.415 150.545 ;
        RECT 94.610 149.885 94.895 150.545 ;
        RECT 95.070 150.215 95.375 150.545 ;
        RECT 95.545 150.215 95.855 150.545 ;
        RECT 95.070 149.885 95.285 150.215 ;
        RECT 96.025 150.095 96.215 150.730 ;
        RECT 93.350 149.545 93.805 149.715 ;
        RECT 93.475 149.115 93.805 149.545 ;
        RECT 93.985 149.545 95.275 149.715 ;
        RECT 93.985 149.125 94.235 149.545 ;
        RECT 94.465 148.905 94.795 149.375 ;
        RECT 95.025 149.125 95.275 149.545 ;
        RECT 95.465 148.905 95.715 150.045 ;
        RECT 95.995 149.965 96.215 150.095 ;
        RECT 95.885 149.115 96.215 149.965 ;
        RECT 96.485 150.635 103.230 150.805 ;
        RECT 96.485 150.045 97.650 150.635 ;
        RECT 103.830 150.465 104.080 151.275 ;
        RECT 104.260 150.930 104.520 151.455 ;
        RECT 104.690 150.465 104.940 151.275 ;
        RECT 105.120 150.945 105.425 151.455 ;
        RECT 97.820 150.215 104.940 150.465 ;
        RECT 105.110 150.215 105.425 150.775 ;
        RECT 105.595 150.730 105.885 151.455 ;
        RECT 106.065 150.725 106.365 151.455 ;
        RECT 106.545 150.545 106.775 151.165 ;
        RECT 106.975 150.895 107.200 151.275 ;
        RECT 107.370 151.065 107.700 151.455 ;
        RECT 107.895 150.945 108.200 151.455 ;
        RECT 106.975 150.715 107.305 150.895 ;
        RECT 106.070 150.215 106.365 150.545 ;
        RECT 106.545 150.215 106.960 150.545 ;
        RECT 96.485 149.820 103.230 150.045 ;
        RECT 96.485 148.905 96.755 149.650 ;
        RECT 96.925 149.080 97.215 149.820 ;
        RECT 97.825 149.805 103.230 149.820 ;
        RECT 97.385 148.910 97.640 149.635 ;
        RECT 97.825 149.080 98.085 149.805 ;
        RECT 98.255 148.910 98.500 149.635 ;
        RECT 98.685 149.080 98.945 149.805 ;
        RECT 99.115 148.910 99.360 149.635 ;
        RECT 99.545 149.080 99.805 149.805 ;
        RECT 99.975 148.910 100.220 149.635 ;
        RECT 100.390 149.080 100.650 149.805 ;
        RECT 100.820 148.910 101.080 149.635 ;
        RECT 101.250 149.080 101.510 149.805 ;
        RECT 101.680 148.910 101.940 149.635 ;
        RECT 102.110 149.080 102.370 149.805 ;
        RECT 102.540 148.910 102.800 149.635 ;
        RECT 102.970 149.080 103.230 149.805 ;
        RECT 103.400 148.910 103.660 149.705 ;
        RECT 103.830 149.080 104.080 150.215 ;
        RECT 97.385 148.905 103.660 148.910 ;
        RECT 104.260 148.905 104.520 149.715 ;
        RECT 104.695 149.075 104.940 150.215 ;
        RECT 105.120 148.905 105.415 149.715 ;
        RECT 105.595 148.905 105.885 150.070 ;
        RECT 107.130 150.045 107.305 150.715 ;
        RECT 107.475 150.215 107.715 150.865 ;
        RECT 107.895 150.215 108.210 150.775 ;
        RECT 108.380 150.465 108.630 151.275 ;
        RECT 108.800 150.930 109.060 151.455 ;
        RECT 109.240 150.465 109.490 151.275 ;
        RECT 109.660 150.895 109.920 151.455 ;
        RECT 110.090 150.805 110.350 151.260 ;
        RECT 110.520 150.975 110.780 151.455 ;
        RECT 110.950 150.805 111.210 151.260 ;
        RECT 111.380 150.975 111.640 151.455 ;
        RECT 111.810 150.805 112.070 151.260 ;
        RECT 112.240 150.975 112.485 151.455 ;
        RECT 112.655 150.805 112.930 151.260 ;
        RECT 113.100 150.975 113.345 151.455 ;
        RECT 113.515 150.805 113.775 151.260 ;
        RECT 113.955 150.975 114.205 151.455 ;
        RECT 114.375 150.805 114.635 151.260 ;
        RECT 114.815 150.975 115.065 151.455 ;
        RECT 115.235 150.805 115.495 151.260 ;
        RECT 115.675 150.975 115.935 151.455 ;
        RECT 116.105 150.805 116.365 151.260 ;
        RECT 116.535 150.975 116.835 151.455 ;
        RECT 110.090 150.635 116.835 150.805 ;
        RECT 117.135 150.635 117.365 151.455 ;
        RECT 117.535 150.655 117.865 151.285 ;
        RECT 108.380 150.215 115.500 150.465 ;
        RECT 106.065 149.685 106.960 150.015 ;
        RECT 107.130 149.855 107.715 150.045 ;
        RECT 106.065 149.515 107.270 149.685 ;
        RECT 106.065 149.085 106.395 149.515 ;
        RECT 106.575 148.905 106.770 149.345 ;
        RECT 106.940 149.085 107.270 149.515 ;
        RECT 107.440 149.085 107.715 149.855 ;
        RECT 107.905 148.905 108.200 149.715 ;
        RECT 108.380 149.075 108.625 150.215 ;
        RECT 108.800 148.905 109.060 149.715 ;
        RECT 109.240 149.080 109.490 150.215 ;
        RECT 115.670 150.095 116.835 150.635 ;
        RECT 117.115 150.215 117.445 150.465 ;
        RECT 115.670 150.045 116.865 150.095 ;
        RECT 117.615 150.055 117.865 150.655 ;
        RECT 118.035 150.635 118.245 151.455 ;
        RECT 118.475 150.730 118.765 151.455 ;
        RECT 110.090 149.925 116.865 150.045 ;
        RECT 110.090 149.820 116.835 149.925 ;
        RECT 110.090 149.805 115.495 149.820 ;
        RECT 109.660 148.910 109.920 149.705 ;
        RECT 110.090 149.080 110.350 149.805 ;
        RECT 110.520 148.910 110.780 149.635 ;
        RECT 110.950 149.080 111.210 149.805 ;
        RECT 111.380 148.910 111.640 149.635 ;
        RECT 111.810 149.080 112.070 149.805 ;
        RECT 112.240 148.910 112.500 149.635 ;
        RECT 112.670 149.080 112.930 149.805 ;
        RECT 113.100 148.910 113.345 149.635 ;
        RECT 113.515 149.080 113.775 149.805 ;
        RECT 113.960 148.910 114.205 149.635 ;
        RECT 114.375 149.080 114.635 149.805 ;
        RECT 114.820 148.910 115.065 149.635 ;
        RECT 115.235 149.080 115.495 149.805 ;
        RECT 115.680 148.910 115.935 149.635 ;
        RECT 116.105 149.080 116.395 149.820 ;
        RECT 109.660 148.905 115.935 148.910 ;
        RECT 116.565 148.905 116.835 149.650 ;
        RECT 117.135 148.905 117.365 150.045 ;
        RECT 117.535 149.075 117.865 150.055 ;
        RECT 118.035 148.905 118.245 150.045 ;
        RECT 118.475 148.905 118.765 150.070 ;
        RECT 118.955 149.875 119.185 151.215 ;
        RECT 119.365 150.375 119.595 151.275 ;
        RECT 119.795 150.675 120.040 151.455 ;
        RECT 120.210 150.915 120.640 151.275 ;
        RECT 121.220 151.085 121.950 151.455 ;
        RECT 120.210 150.725 121.950 150.915 ;
        RECT 120.210 150.495 120.430 150.725 ;
        RECT 119.365 149.695 119.705 150.375 ;
        RECT 118.955 149.495 119.705 149.695 ;
        RECT 119.885 150.195 120.430 150.495 ;
        RECT 118.955 149.105 119.195 149.495 ;
        RECT 119.365 148.905 119.715 149.315 ;
        RECT 119.885 149.085 120.215 150.195 ;
        RECT 120.600 149.925 121.025 150.545 ;
        RECT 121.220 149.925 121.480 150.545 ;
        RECT 121.690 150.215 121.950 150.725 ;
        RECT 120.385 149.555 121.410 149.755 ;
        RECT 120.385 149.085 120.565 149.555 ;
        RECT 120.735 148.905 121.065 149.385 ;
        RECT 121.240 149.085 121.410 149.555 ;
        RECT 121.675 148.905 121.960 150.045 ;
        RECT 122.150 149.085 122.430 151.275 ;
        RECT 122.615 150.780 122.875 151.285 ;
        RECT 123.055 151.075 123.385 151.455 ;
        RECT 123.565 150.905 123.735 151.285 ;
        RECT 122.615 149.980 122.795 150.780 ;
        RECT 123.070 150.735 123.735 150.905 ;
        RECT 123.070 150.480 123.240 150.735 ;
        RECT 123.995 150.705 125.205 151.455 ;
        RECT 122.965 150.150 123.240 150.480 ;
        RECT 123.465 150.185 123.805 150.555 ;
        RECT 123.070 150.005 123.240 150.150 ;
        RECT 122.615 149.075 122.885 149.980 ;
        RECT 123.070 149.835 123.745 150.005 ;
        RECT 123.055 148.905 123.385 149.665 ;
        RECT 123.565 149.075 123.745 149.835 ;
        RECT 123.995 149.995 124.515 150.535 ;
        RECT 124.685 150.165 125.205 150.705 ;
        RECT 123.995 148.905 125.205 149.995 ;
        RECT 53.990 148.735 125.290 148.905 ;
        RECT 54.075 147.645 55.285 148.735 ;
        RECT 54.075 146.935 54.595 147.475 ;
        RECT 54.765 147.105 55.285 147.645 ;
        RECT 56.375 148.015 56.835 148.565 ;
        RECT 57.025 148.015 57.355 148.735 ;
        RECT 54.075 146.185 55.285 146.935 ;
        RECT 56.375 146.645 56.625 148.015 ;
        RECT 57.555 147.845 57.855 148.395 ;
        RECT 58.025 148.065 58.305 148.735 ;
        RECT 56.915 147.675 57.855 147.845 ;
        RECT 56.915 147.425 57.085 147.675 ;
        RECT 58.225 147.425 58.490 147.785 ;
        RECT 58.680 147.585 58.940 148.735 ;
        RECT 59.115 147.660 59.370 148.565 ;
        RECT 59.540 147.975 59.870 148.735 ;
        RECT 60.085 147.805 60.255 148.565 ;
        RECT 60.715 148.065 60.995 148.735 ;
        RECT 56.795 147.095 57.085 147.425 ;
        RECT 57.255 147.175 57.595 147.425 ;
        RECT 57.815 147.175 58.490 147.425 ;
        RECT 56.915 147.005 57.085 147.095 ;
        RECT 56.915 146.815 58.305 147.005 ;
        RECT 56.375 146.355 56.935 146.645 ;
        RECT 57.105 146.185 57.355 146.645 ;
        RECT 57.975 146.455 58.305 146.815 ;
        RECT 58.680 146.185 58.940 147.025 ;
        RECT 59.115 146.930 59.285 147.660 ;
        RECT 59.540 147.635 60.255 147.805 ;
        RECT 61.165 147.845 61.465 148.395 ;
        RECT 61.665 148.015 61.995 148.735 ;
        RECT 62.185 148.015 62.645 148.565 ;
        RECT 59.540 147.425 59.710 147.635 ;
        RECT 59.455 147.095 59.710 147.425 ;
        RECT 59.115 146.355 59.370 146.930 ;
        RECT 59.540 146.905 59.710 147.095 ;
        RECT 59.990 147.085 60.345 147.455 ;
        RECT 60.530 147.425 60.795 147.785 ;
        RECT 61.165 147.675 62.105 147.845 ;
        RECT 61.935 147.425 62.105 147.675 ;
        RECT 60.530 147.175 61.205 147.425 ;
        RECT 61.425 147.175 61.765 147.425 ;
        RECT 61.935 147.095 62.225 147.425 ;
        RECT 61.935 147.005 62.105 147.095 ;
        RECT 59.540 146.735 60.255 146.905 ;
        RECT 59.540 146.185 59.870 146.565 ;
        RECT 60.085 146.355 60.255 146.735 ;
        RECT 60.715 146.815 62.105 147.005 ;
        RECT 60.715 146.455 61.045 146.815 ;
        RECT 62.395 146.645 62.645 148.015 ;
        RECT 62.815 147.675 63.130 148.735 ;
        RECT 63.760 148.230 64.375 148.735 ;
        RECT 62.875 146.845 63.140 147.425 ;
        RECT 63.310 147.345 63.585 148.005 ;
        RECT 63.780 147.695 64.015 148.060 ;
        RECT 64.185 148.055 64.375 148.230 ;
        RECT 64.545 148.225 65.020 148.565 ;
        RECT 64.185 147.865 64.515 148.055 ;
        RECT 64.740 147.695 64.930 147.990 ;
        RECT 65.190 147.890 65.405 148.735 ;
        RECT 65.605 147.895 65.890 148.565 ;
        RECT 63.780 147.525 65.550 147.695 ;
        RECT 63.310 147.115 64.145 147.345 ;
        RECT 61.665 146.185 61.915 146.645 ;
        RECT 62.085 146.355 62.645 146.645 ;
        RECT 62.815 146.185 63.085 146.675 ;
        RECT 63.310 146.405 63.585 147.115 ;
        RECT 64.315 146.670 64.570 147.525 ;
        RECT 63.785 146.405 64.570 146.670 ;
        RECT 64.740 146.865 65.150 147.345 ;
        RECT 65.320 147.095 65.550 147.525 ;
        RECT 65.720 147.545 65.890 147.895 ;
        RECT 66.060 147.725 66.325 148.735 ;
        RECT 66.955 147.570 67.245 148.735 ;
        RECT 67.880 147.590 68.175 148.735 ;
        RECT 65.720 147.025 66.325 147.545 ;
        RECT 64.740 146.405 64.950 146.865 ;
        RECT 65.720 146.815 65.890 147.025 ;
        RECT 65.140 146.185 65.470 146.680 ;
        RECT 65.645 146.355 65.890 146.815 ;
        RECT 66.060 146.185 66.325 146.845 ;
        RECT 66.955 146.185 67.245 146.910 ;
        RECT 67.880 146.185 68.175 147.005 ;
        RECT 68.345 146.735 68.575 148.435 ;
        RECT 68.790 147.930 69.045 148.735 ;
        RECT 69.245 148.120 69.575 148.565 ;
        RECT 69.745 148.290 70.020 148.735 ;
        RECT 70.255 148.120 70.585 148.565 ;
        RECT 69.245 147.940 70.585 148.120 ;
        RECT 71.045 147.760 71.375 148.425 ;
        RECT 71.575 147.935 71.905 148.735 ;
        RECT 68.790 147.590 71.375 147.760 ;
        RECT 72.080 147.595 72.415 148.565 ;
        RECT 72.585 147.935 72.915 148.735 ;
        RECT 73.315 147.765 73.565 148.565 ;
        RECT 73.750 148.015 74.080 148.735 ;
        RECT 74.300 147.765 74.550 148.565 ;
        RECT 74.725 148.355 75.055 148.735 ;
        RECT 72.595 147.595 74.650 147.765 ;
        RECT 68.790 146.975 69.100 147.590 ;
        RECT 72.080 147.375 72.255 147.595 ;
        RECT 72.595 147.415 72.820 147.595 ;
        RECT 69.270 147.145 69.600 147.375 ;
        RECT 69.770 147.145 70.240 147.375 ;
        RECT 70.410 147.205 70.865 147.375 ;
        RECT 70.410 147.145 70.860 147.205 ;
        RECT 71.050 147.145 71.385 147.375 ;
        RECT 72.075 147.205 72.255 147.375 ;
        RECT 68.790 146.795 71.375 146.975 ;
        RECT 68.345 146.355 68.565 146.735 ;
        RECT 68.735 146.185 69.585 146.545 ;
        RECT 70.065 146.375 70.395 146.795 ;
        RECT 70.600 146.185 70.875 146.625 ;
        RECT 71.045 146.375 71.375 146.795 ;
        RECT 71.565 146.185 71.895 146.910 ;
        RECT 72.080 146.905 72.255 147.205 ;
        RECT 72.425 147.175 72.820 147.415 ;
        RECT 72.080 146.440 72.415 146.905 ;
        RECT 72.085 146.395 72.415 146.440 ;
        RECT 72.585 146.185 72.820 146.990 ;
        RECT 72.990 146.515 73.250 147.425 ;
        RECT 73.560 147.405 73.730 147.425 ;
        RECT 73.430 146.515 73.730 147.405 ;
        RECT 73.905 146.520 74.260 147.425 ;
        RECT 74.480 146.685 74.650 147.595 ;
        RECT 74.820 146.855 75.025 148.175 ;
        RECT 75.325 147.990 75.595 148.735 ;
        RECT 76.225 148.730 82.500 148.735 ;
        RECT 75.765 147.820 76.055 148.560 ;
        RECT 76.225 148.005 76.480 148.730 ;
        RECT 76.665 147.835 76.925 148.560 ;
        RECT 77.095 148.005 77.340 148.730 ;
        RECT 77.525 147.835 77.785 148.560 ;
        RECT 77.955 148.005 78.200 148.730 ;
        RECT 78.385 147.835 78.645 148.560 ;
        RECT 78.815 148.005 79.060 148.730 ;
        RECT 79.230 147.835 79.490 148.560 ;
        RECT 79.660 148.005 79.920 148.730 ;
        RECT 80.090 147.835 80.350 148.560 ;
        RECT 80.520 148.005 80.780 148.730 ;
        RECT 80.950 147.835 81.210 148.560 ;
        RECT 81.380 148.005 81.640 148.730 ;
        RECT 81.810 147.835 82.070 148.560 ;
        RECT 82.240 147.935 82.500 148.730 ;
        RECT 76.665 147.820 82.070 147.835 ;
        RECT 75.325 147.595 82.070 147.820 ;
        RECT 75.325 147.005 76.490 147.595 ;
        RECT 82.670 147.425 82.920 148.560 ;
        RECT 83.100 147.925 83.360 148.735 ;
        RECT 83.535 147.425 83.780 148.565 ;
        RECT 83.960 147.925 84.255 148.735 ;
        RECT 84.525 147.725 84.695 148.565 ;
        RECT 84.865 148.395 86.035 148.565 ;
        RECT 84.865 147.895 85.195 148.395 ;
        RECT 85.705 148.355 86.035 148.395 ;
        RECT 86.225 148.315 86.580 148.735 ;
        RECT 85.365 148.135 85.595 148.225 ;
        RECT 86.750 148.135 87.000 148.565 ;
        RECT 85.365 147.895 87.000 148.135 ;
        RECT 87.170 147.975 87.500 148.735 ;
        RECT 87.670 147.895 87.925 148.565 ;
        RECT 84.525 147.555 87.585 147.725 ;
        RECT 76.660 147.175 83.780 147.425 ;
        RECT 75.325 146.835 82.070 147.005 ;
        RECT 74.480 146.355 74.975 146.685 ;
        RECT 75.325 146.185 75.625 146.665 ;
        RECT 75.795 146.380 76.055 146.835 ;
        RECT 76.225 146.185 76.485 146.665 ;
        RECT 76.665 146.380 76.925 146.835 ;
        RECT 77.095 146.185 77.345 146.665 ;
        RECT 77.525 146.380 77.785 146.835 ;
        RECT 77.955 146.185 78.205 146.665 ;
        RECT 78.385 146.380 78.645 146.835 ;
        RECT 78.815 146.185 79.060 146.665 ;
        RECT 79.230 146.380 79.505 146.835 ;
        RECT 79.675 146.185 79.920 146.665 ;
        RECT 80.090 146.380 80.350 146.835 ;
        RECT 80.520 146.185 80.780 146.665 ;
        RECT 80.950 146.380 81.210 146.835 ;
        RECT 81.380 146.185 81.640 146.665 ;
        RECT 81.810 146.380 82.070 146.835 ;
        RECT 82.240 146.185 82.500 146.745 ;
        RECT 82.670 146.365 82.920 147.175 ;
        RECT 83.100 146.185 83.360 146.710 ;
        RECT 83.530 146.365 83.780 147.175 ;
        RECT 83.950 146.865 84.265 147.425 ;
        RECT 84.435 147.175 84.790 147.385 ;
        RECT 84.960 147.175 85.405 147.375 ;
        RECT 85.575 147.175 86.050 147.375 ;
        RECT 84.525 146.835 85.590 147.005 ;
        RECT 83.960 146.185 84.265 146.695 ;
        RECT 84.525 146.355 84.695 146.835 ;
        RECT 84.865 146.185 85.195 146.665 ;
        RECT 85.420 146.605 85.590 146.835 ;
        RECT 85.770 146.775 86.050 147.175 ;
        RECT 86.320 147.175 86.650 147.375 ;
        RECT 86.820 147.175 87.185 147.375 ;
        RECT 86.320 146.775 86.605 147.175 ;
        RECT 87.415 147.005 87.585 147.555 ;
        RECT 86.785 146.835 87.585 147.005 ;
        RECT 86.785 146.605 86.955 146.835 ;
        RECT 87.755 146.765 87.925 147.895 ;
        RECT 88.095 147.545 88.265 148.735 ;
        RECT 88.585 147.760 88.915 148.425 ;
        RECT 89.375 148.120 89.705 148.565 ;
        RECT 89.940 148.290 90.215 148.735 ;
        RECT 90.385 148.120 90.715 148.565 ;
        RECT 89.375 147.940 90.715 148.120 ;
        RECT 90.915 147.930 91.170 148.735 ;
        RECT 88.585 147.590 91.170 147.760 ;
        RECT 88.575 147.145 88.910 147.375 ;
        RECT 89.095 147.205 89.550 147.375 ;
        RECT 89.100 147.145 89.550 147.205 ;
        RECT 89.720 147.145 90.190 147.375 ;
        RECT 90.360 147.145 90.690 147.375 ;
        RECT 87.740 146.695 87.925 146.765 ;
        RECT 87.715 146.685 87.925 146.695 ;
        RECT 85.420 146.355 86.955 146.605 ;
        RECT 87.125 146.185 87.455 146.665 ;
        RECT 87.670 146.355 87.925 146.685 ;
        RECT 88.095 146.185 88.265 147.080 ;
        RECT 90.860 146.975 91.170 147.590 ;
        RECT 88.585 146.795 91.170 146.975 ;
        RECT 88.585 146.375 88.915 146.795 ;
        RECT 89.085 146.185 89.360 146.625 ;
        RECT 89.565 146.375 89.895 146.795 ;
        RECT 91.385 146.735 91.615 148.435 ;
        RECT 91.785 147.590 92.080 148.735 ;
        RECT 92.715 147.570 93.005 148.735 ;
        RECT 93.175 147.765 93.485 148.565 ;
        RECT 93.655 147.935 93.965 148.735 ;
        RECT 94.135 148.105 94.395 148.565 ;
        RECT 94.565 148.275 94.820 148.735 ;
        RECT 94.995 148.105 95.255 148.565 ;
        RECT 94.135 147.935 95.255 148.105 ;
        RECT 93.175 147.595 94.205 147.765 ;
        RECT 90.375 146.185 91.225 146.545 ;
        RECT 91.395 146.355 91.615 146.735 ;
        RECT 91.785 146.185 92.080 147.005 ;
        RECT 92.715 146.185 93.005 146.910 ;
        RECT 93.175 146.685 93.345 147.595 ;
        RECT 93.515 146.855 93.865 147.425 ;
        RECT 94.035 147.345 94.205 147.595 ;
        RECT 94.995 147.685 95.255 147.935 ;
        RECT 95.425 147.865 95.710 148.735 ;
        RECT 95.935 148.140 96.370 148.565 ;
        RECT 96.540 148.310 96.925 148.735 ;
        RECT 95.935 147.970 96.925 148.140 ;
        RECT 94.995 147.515 95.750 147.685 ;
        RECT 94.035 147.175 95.175 147.345 ;
        RECT 95.345 147.005 95.750 147.515 ;
        RECT 95.935 147.095 96.420 147.800 ;
        RECT 96.590 147.425 96.925 147.970 ;
        RECT 97.095 147.775 97.520 148.565 ;
        RECT 97.690 148.140 97.965 148.565 ;
        RECT 98.135 148.310 98.520 148.735 ;
        RECT 97.690 147.945 98.520 148.140 ;
        RECT 97.095 147.595 98.000 147.775 ;
        RECT 96.590 147.095 97.000 147.425 ;
        RECT 97.170 147.095 98.000 147.595 ;
        RECT 98.170 147.425 98.520 147.945 ;
        RECT 98.690 147.775 98.935 148.565 ;
        RECT 99.125 148.140 99.380 148.565 ;
        RECT 99.550 148.310 99.935 148.735 ;
        RECT 99.125 147.945 99.935 148.140 ;
        RECT 98.690 147.595 99.415 147.775 ;
        RECT 98.170 147.095 98.595 147.425 ;
        RECT 98.765 147.095 99.415 147.595 ;
        RECT 99.585 147.425 99.935 147.945 ;
        RECT 100.105 147.595 100.365 148.565 ;
        RECT 100.545 147.925 100.840 148.735 ;
        RECT 99.585 147.095 100.010 147.425 ;
        RECT 94.100 146.835 95.750 147.005 ;
        RECT 96.590 146.925 96.925 147.095 ;
        RECT 97.170 146.925 97.520 147.095 ;
        RECT 98.170 146.925 98.520 147.095 ;
        RECT 98.765 146.925 98.935 147.095 ;
        RECT 99.585 146.925 99.935 147.095 ;
        RECT 100.180 146.925 100.365 147.595 ;
        RECT 101.020 147.425 101.265 148.565 ;
        RECT 101.440 147.925 101.700 148.735 ;
        RECT 102.300 148.730 108.575 148.735 ;
        RECT 101.880 147.425 102.130 148.560 ;
        RECT 102.300 147.935 102.560 148.730 ;
        RECT 102.730 147.835 102.990 148.560 ;
        RECT 103.160 148.005 103.420 148.730 ;
        RECT 103.590 147.835 103.850 148.560 ;
        RECT 104.020 148.005 104.280 148.730 ;
        RECT 104.450 147.835 104.710 148.560 ;
        RECT 104.880 148.005 105.140 148.730 ;
        RECT 105.310 147.835 105.570 148.560 ;
        RECT 105.740 148.005 105.985 148.730 ;
        RECT 106.155 147.835 106.415 148.560 ;
        RECT 106.600 148.005 106.845 148.730 ;
        RECT 107.015 147.835 107.275 148.560 ;
        RECT 107.460 148.005 107.705 148.730 ;
        RECT 107.875 147.835 108.135 148.560 ;
        RECT 108.320 148.005 108.575 148.730 ;
        RECT 102.730 147.820 108.135 147.835 ;
        RECT 108.745 147.820 109.035 148.560 ;
        RECT 109.205 147.990 109.475 148.735 ;
        RECT 109.755 148.145 109.995 148.535 ;
        RECT 110.165 148.325 110.515 148.735 ;
        RECT 109.755 147.945 110.505 148.145 ;
        RECT 102.730 147.595 109.475 147.820 ;
        RECT 93.175 146.355 93.475 146.685 ;
        RECT 93.645 146.185 93.920 146.665 ;
        RECT 94.100 146.445 94.395 146.835 ;
        RECT 94.565 146.185 94.820 146.665 ;
        RECT 94.995 146.445 95.255 146.835 ;
        RECT 95.935 146.755 96.925 146.925 ;
        RECT 95.425 146.185 95.705 146.665 ;
        RECT 95.935 146.355 96.370 146.755 ;
        RECT 96.540 146.185 96.925 146.585 ;
        RECT 97.095 146.355 97.520 146.925 ;
        RECT 97.710 146.755 98.520 146.925 ;
        RECT 97.710 146.355 97.965 146.755 ;
        RECT 98.135 146.185 98.520 146.585 ;
        RECT 98.690 146.355 98.935 146.925 ;
        RECT 99.125 146.755 99.935 146.925 ;
        RECT 99.125 146.355 99.380 146.755 ;
        RECT 99.550 146.185 99.935 146.585 ;
        RECT 100.105 146.355 100.365 146.925 ;
        RECT 100.535 146.865 100.850 147.425 ;
        RECT 101.020 147.175 108.140 147.425 ;
        RECT 100.535 146.185 100.840 146.695 ;
        RECT 101.020 146.365 101.270 147.175 ;
        RECT 101.440 146.185 101.700 146.710 ;
        RECT 101.880 146.365 102.130 147.175 ;
        RECT 108.310 147.005 109.475 147.595 ;
        RECT 102.730 146.835 109.475 147.005 ;
        RECT 102.300 146.185 102.560 146.745 ;
        RECT 102.730 146.380 102.990 146.835 ;
        RECT 103.160 146.185 103.420 146.665 ;
        RECT 103.590 146.380 103.850 146.835 ;
        RECT 104.020 146.185 104.280 146.665 ;
        RECT 104.450 146.380 104.710 146.835 ;
        RECT 104.880 146.185 105.125 146.665 ;
        RECT 105.295 146.380 105.570 146.835 ;
        RECT 105.740 146.185 105.985 146.665 ;
        RECT 106.155 146.380 106.415 146.835 ;
        RECT 106.595 146.185 106.845 146.665 ;
        RECT 107.015 146.380 107.275 146.835 ;
        RECT 107.455 146.185 107.705 146.665 ;
        RECT 107.875 146.380 108.135 146.835 ;
        RECT 108.315 146.185 108.575 146.665 ;
        RECT 108.745 146.380 109.005 146.835 ;
        RECT 109.175 146.185 109.475 146.665 ;
        RECT 109.755 146.425 109.985 147.765 ;
        RECT 110.165 147.265 110.505 147.945 ;
        RECT 110.685 147.445 111.015 148.555 ;
        RECT 111.185 148.085 111.365 148.555 ;
        RECT 111.535 148.255 111.865 148.735 ;
        RECT 112.040 148.085 112.210 148.555 ;
        RECT 111.185 147.885 112.210 148.085 ;
        RECT 110.165 146.365 110.395 147.265 ;
        RECT 110.685 147.145 111.230 147.445 ;
        RECT 110.595 146.185 110.840 146.965 ;
        RECT 111.010 146.915 111.230 147.145 ;
        RECT 111.400 147.095 111.825 147.715 ;
        RECT 112.020 147.095 112.280 147.715 ;
        RECT 112.475 147.595 112.760 148.735 ;
        RECT 112.490 146.915 112.750 147.425 ;
        RECT 111.010 146.725 112.750 146.915 ;
        RECT 111.010 146.365 111.440 146.725 ;
        RECT 112.020 146.185 112.750 146.555 ;
        RECT 112.950 146.365 113.230 148.555 ;
        RECT 113.435 148.145 113.675 148.535 ;
        RECT 113.845 148.325 114.195 148.735 ;
        RECT 113.435 147.945 114.185 148.145 ;
        RECT 113.435 146.425 113.665 147.765 ;
        RECT 113.845 147.265 114.185 147.945 ;
        RECT 114.365 147.445 114.695 148.555 ;
        RECT 114.865 148.085 115.045 148.555 ;
        RECT 115.215 148.255 115.545 148.735 ;
        RECT 115.720 148.085 115.890 148.555 ;
        RECT 114.865 147.885 115.890 148.085 ;
        RECT 113.845 146.365 114.075 147.265 ;
        RECT 114.365 147.145 114.910 147.445 ;
        RECT 114.275 146.185 114.520 146.965 ;
        RECT 114.690 146.915 114.910 147.145 ;
        RECT 115.080 147.095 115.505 147.715 ;
        RECT 115.700 147.095 115.960 147.715 ;
        RECT 116.155 147.595 116.440 148.735 ;
        RECT 116.170 146.915 116.430 147.425 ;
        RECT 114.690 146.725 116.430 146.915 ;
        RECT 114.690 146.365 115.120 146.725 ;
        RECT 115.700 146.185 116.430 146.555 ;
        RECT 116.630 146.365 116.910 148.555 ;
        RECT 117.155 147.595 117.365 148.735 ;
        RECT 117.535 147.585 117.865 148.565 ;
        RECT 118.035 147.595 118.265 148.735 ;
        RECT 117.155 146.185 117.365 147.005 ;
        RECT 117.535 146.985 117.785 147.585 ;
        RECT 118.475 147.570 118.765 148.735 ;
        RECT 118.955 148.145 119.195 148.535 ;
        RECT 119.365 148.325 119.715 148.735 ;
        RECT 118.955 147.945 119.705 148.145 ;
        RECT 117.955 147.175 118.285 147.425 ;
        RECT 117.535 146.355 117.865 146.985 ;
        RECT 118.035 146.185 118.265 147.005 ;
        RECT 118.475 146.185 118.765 146.910 ;
        RECT 118.955 146.425 119.185 147.765 ;
        RECT 119.365 147.265 119.705 147.945 ;
        RECT 119.885 147.445 120.215 148.555 ;
        RECT 120.385 148.085 120.565 148.555 ;
        RECT 120.735 148.255 121.065 148.735 ;
        RECT 121.240 148.085 121.410 148.555 ;
        RECT 120.385 147.885 121.410 148.085 ;
        RECT 119.365 146.365 119.595 147.265 ;
        RECT 119.885 147.145 120.430 147.445 ;
        RECT 119.795 146.185 120.040 146.965 ;
        RECT 120.210 146.915 120.430 147.145 ;
        RECT 120.600 147.095 121.025 147.715 ;
        RECT 121.220 147.095 121.480 147.715 ;
        RECT 121.675 147.595 121.960 148.735 ;
        RECT 121.690 146.915 121.950 147.425 ;
        RECT 120.210 146.725 121.950 146.915 ;
        RECT 120.210 146.365 120.640 146.725 ;
        RECT 121.220 146.185 121.950 146.555 ;
        RECT 122.150 146.365 122.430 148.555 ;
        RECT 122.615 147.660 122.885 148.565 ;
        RECT 123.055 147.975 123.385 148.735 ;
        RECT 123.565 147.805 123.735 148.565 ;
        RECT 122.615 146.860 122.785 147.660 ;
        RECT 123.070 147.635 123.735 147.805 ;
        RECT 123.995 147.645 125.205 148.735 ;
        RECT 123.070 147.490 123.240 147.635 ;
        RECT 122.955 147.160 123.240 147.490 ;
        RECT 123.070 146.905 123.240 147.160 ;
        RECT 123.475 147.085 123.805 147.455 ;
        RECT 123.995 147.105 124.515 147.645 ;
        RECT 124.685 146.935 125.205 147.475 ;
        RECT 122.615 146.355 122.875 146.860 ;
        RECT 123.070 146.735 123.735 146.905 ;
        RECT 123.055 146.185 123.385 146.565 ;
        RECT 123.565 146.355 123.735 146.735 ;
        RECT 123.995 146.185 125.205 146.935 ;
        RECT 53.990 146.015 125.290 146.185 ;
        RECT 54.075 145.265 55.285 146.015 ;
        RECT 54.075 144.725 54.595 145.265 ;
        RECT 55.460 145.175 55.720 146.015 ;
        RECT 55.895 145.270 56.150 145.845 ;
        RECT 56.320 145.635 56.650 146.015 ;
        RECT 56.865 145.465 57.035 145.845 ;
        RECT 56.320 145.295 57.035 145.465 ;
        RECT 54.765 144.555 55.285 145.095 ;
        RECT 54.075 143.465 55.285 144.555 ;
        RECT 55.460 143.465 55.720 144.615 ;
        RECT 55.895 144.540 56.065 145.270 ;
        RECT 56.320 145.105 56.490 145.295 ;
        RECT 57.295 145.215 57.605 146.015 ;
        RECT 57.810 145.215 58.505 145.845 ;
        RECT 58.675 145.215 58.985 146.015 ;
        RECT 59.190 145.215 59.885 145.845 ;
        RECT 60.100 145.555 60.850 145.845 ;
        RECT 61.360 145.555 61.690 146.015 ;
        RECT 56.235 144.775 56.490 145.105 ;
        RECT 56.320 144.565 56.490 144.775 ;
        RECT 56.770 144.745 57.125 145.115 ;
        RECT 57.305 144.775 57.640 145.045 ;
        RECT 57.810 144.615 57.980 145.215 ;
        RECT 59.190 145.165 59.365 145.215 ;
        RECT 58.150 144.775 58.485 145.025 ;
        RECT 58.685 144.775 59.020 145.045 ;
        RECT 59.190 144.615 59.360 145.165 ;
        RECT 59.530 144.775 59.865 145.025 ;
        RECT 55.895 143.635 56.150 144.540 ;
        RECT 56.320 144.395 57.035 144.565 ;
        RECT 56.320 143.465 56.650 144.225 ;
        RECT 56.865 143.635 57.035 144.395 ;
        RECT 57.295 143.465 57.575 144.605 ;
        RECT 57.745 143.635 58.075 144.615 ;
        RECT 58.245 143.465 58.505 144.605 ;
        RECT 58.675 143.465 58.955 144.605 ;
        RECT 59.125 143.635 59.455 144.615 ;
        RECT 59.625 143.465 59.885 144.605 ;
        RECT 60.100 144.265 60.470 145.555 ;
        RECT 61.910 145.365 62.180 145.575 ;
        RECT 60.845 145.195 62.180 145.365 ;
        RECT 62.355 145.355 62.630 146.015 ;
        RECT 62.800 145.385 63.050 145.845 ;
        RECT 63.225 145.520 63.555 146.015 ;
        RECT 60.845 145.025 61.015 145.195 ;
        RECT 62.800 145.175 62.970 145.385 ;
        RECT 63.735 145.350 63.965 145.795 ;
        RECT 60.640 144.775 61.015 145.025 ;
        RECT 61.185 144.785 61.660 145.025 ;
        RECT 61.830 144.785 62.180 145.025 ;
        RECT 60.845 144.605 61.015 144.775 ;
        RECT 62.355 144.655 62.970 145.175 ;
        RECT 63.140 144.675 63.370 145.105 ;
        RECT 63.555 144.855 63.965 145.350 ;
        RECT 64.135 145.530 64.925 145.795 ;
        RECT 64.135 144.675 64.390 145.530 ;
        RECT 65.315 145.385 65.645 145.745 ;
        RECT 66.275 145.555 66.525 146.015 ;
        RECT 66.695 145.555 67.245 145.845 ;
        RECT 64.560 144.855 64.945 145.335 ;
        RECT 65.315 145.195 66.705 145.385 ;
        RECT 66.535 145.105 66.705 145.195 ;
        RECT 65.115 144.775 65.805 145.025 ;
        RECT 66.035 144.775 66.365 145.025 ;
        RECT 66.535 144.775 66.825 145.105 ;
        RECT 60.845 144.435 62.180 144.605 ;
        RECT 61.900 144.275 62.180 144.435 ;
        RECT 60.100 144.095 61.270 144.265 ;
        RECT 60.555 143.465 60.770 143.925 ;
        RECT 60.940 143.635 61.270 144.095 ;
        RECT 61.440 143.465 61.690 144.265 ;
        RECT 62.355 143.465 62.615 144.475 ;
        RECT 62.785 144.305 62.955 144.655 ;
        RECT 63.140 144.505 64.930 144.675 ;
        RECT 62.785 143.635 63.060 144.305 ;
        RECT 63.260 143.465 63.475 144.310 ;
        RECT 63.700 144.210 63.950 144.505 ;
        RECT 64.175 144.145 64.505 144.335 ;
        RECT 63.660 143.635 64.135 143.975 ;
        RECT 64.315 143.970 64.505 144.145 ;
        RECT 64.675 144.140 64.930 144.505 ;
        RECT 65.115 144.335 65.430 144.775 ;
        RECT 66.535 144.525 66.705 144.775 ;
        RECT 65.765 144.355 66.705 144.525 ;
        RECT 64.315 143.465 64.945 143.970 ;
        RECT 65.315 143.465 65.595 144.135 ;
        RECT 65.765 143.805 66.065 144.355 ;
        RECT 66.995 144.185 67.245 145.555 ;
        RECT 67.415 145.215 67.705 146.015 ;
        RECT 67.935 145.535 68.215 146.015 ;
        RECT 68.385 145.365 68.645 145.755 ;
        RECT 68.820 145.535 69.075 146.015 ;
        RECT 69.245 145.365 69.540 145.755 ;
        RECT 69.720 145.535 69.995 146.015 ;
        RECT 70.165 145.515 70.465 145.845 ;
        RECT 70.725 145.535 71.025 146.015 ;
        RECT 67.890 145.195 69.540 145.365 ;
        RECT 67.890 144.685 68.295 145.195 ;
        RECT 68.465 144.855 69.605 145.025 ;
        RECT 66.275 143.465 66.605 144.185 ;
        RECT 66.795 143.635 67.245 144.185 ;
        RECT 67.415 143.465 67.705 144.605 ;
        RECT 67.890 144.515 68.645 144.685 ;
        RECT 67.930 143.465 68.215 144.335 ;
        RECT 68.385 144.265 68.645 144.515 ;
        RECT 69.435 144.605 69.605 144.855 ;
        RECT 69.775 144.775 70.125 145.345 ;
        RECT 70.295 144.605 70.465 145.515 ;
        RECT 71.195 145.365 71.455 145.820 ;
        RECT 71.625 145.535 71.885 146.015 ;
        RECT 72.065 145.365 72.325 145.820 ;
        RECT 72.495 145.535 72.745 146.015 ;
        RECT 72.925 145.365 73.185 145.820 ;
        RECT 73.355 145.535 73.605 146.015 ;
        RECT 73.785 145.365 74.045 145.820 ;
        RECT 74.215 145.535 74.460 146.015 ;
        RECT 74.630 145.365 74.905 145.820 ;
        RECT 75.075 145.535 75.320 146.015 ;
        RECT 75.490 145.365 75.750 145.820 ;
        RECT 75.920 145.535 76.180 146.015 ;
        RECT 76.350 145.365 76.610 145.820 ;
        RECT 76.780 145.535 77.040 146.015 ;
        RECT 77.210 145.365 77.470 145.820 ;
        RECT 77.640 145.455 77.900 146.015 ;
        RECT 69.435 144.435 70.465 144.605 ;
        RECT 68.385 144.095 69.505 144.265 ;
        RECT 68.385 143.635 68.645 144.095 ;
        RECT 68.820 143.465 69.075 143.925 ;
        RECT 69.245 143.635 69.505 144.095 ;
        RECT 69.675 143.465 69.985 144.265 ;
        RECT 70.155 143.635 70.465 144.435 ;
        RECT 70.725 145.195 77.470 145.365 ;
        RECT 70.725 144.605 71.890 145.195 ;
        RECT 78.070 145.025 78.320 145.835 ;
        RECT 78.500 145.490 78.760 146.015 ;
        RECT 78.930 145.025 79.180 145.835 ;
        RECT 79.360 145.505 79.665 146.015 ;
        RECT 72.060 144.775 79.180 145.025 ;
        RECT 79.350 144.775 79.665 145.335 ;
        RECT 79.835 145.290 80.125 146.015 ;
        RECT 81.215 145.505 81.520 146.015 ;
        RECT 81.215 144.775 81.530 145.335 ;
        RECT 81.700 145.025 81.950 145.835 ;
        RECT 82.120 145.490 82.380 146.015 ;
        RECT 82.560 145.025 82.810 145.835 ;
        RECT 82.980 145.455 83.240 146.015 ;
        RECT 83.410 145.365 83.670 145.820 ;
        RECT 83.840 145.535 84.100 146.015 ;
        RECT 84.270 145.365 84.530 145.820 ;
        RECT 84.700 145.535 84.960 146.015 ;
        RECT 85.130 145.365 85.390 145.820 ;
        RECT 85.560 145.535 85.805 146.015 ;
        RECT 85.975 145.365 86.250 145.820 ;
        RECT 86.420 145.535 86.665 146.015 ;
        RECT 86.835 145.365 87.095 145.820 ;
        RECT 87.275 145.535 87.525 146.015 ;
        RECT 87.695 145.365 87.955 145.820 ;
        RECT 88.135 145.535 88.385 146.015 ;
        RECT 88.555 145.365 88.815 145.820 ;
        RECT 88.995 145.535 89.255 146.015 ;
        RECT 89.425 145.365 89.685 145.820 ;
        RECT 89.855 145.535 90.155 146.015 ;
        RECT 90.505 145.535 90.805 146.015 ;
        RECT 90.975 145.365 91.235 145.820 ;
        RECT 91.405 145.535 91.665 146.015 ;
        RECT 91.845 145.365 92.105 145.820 ;
        RECT 92.275 145.535 92.525 146.015 ;
        RECT 92.705 145.365 92.965 145.820 ;
        RECT 93.135 145.535 93.385 146.015 ;
        RECT 93.565 145.365 93.825 145.820 ;
        RECT 93.995 145.535 94.240 146.015 ;
        RECT 94.410 145.365 94.685 145.820 ;
        RECT 94.855 145.535 95.100 146.015 ;
        RECT 95.270 145.365 95.530 145.820 ;
        RECT 95.700 145.535 95.960 146.015 ;
        RECT 96.130 145.365 96.390 145.820 ;
        RECT 96.560 145.535 96.820 146.015 ;
        RECT 96.990 145.365 97.250 145.820 ;
        RECT 97.420 145.455 97.680 146.015 ;
        RECT 83.410 145.195 90.155 145.365 ;
        RECT 81.700 144.775 88.820 145.025 ;
        RECT 70.725 144.380 77.470 144.605 ;
        RECT 70.725 143.465 70.995 144.210 ;
        RECT 71.165 143.640 71.455 144.380 ;
        RECT 72.065 144.365 77.470 144.380 ;
        RECT 71.625 143.470 71.880 144.195 ;
        RECT 72.065 143.640 72.325 144.365 ;
        RECT 72.495 143.470 72.740 144.195 ;
        RECT 72.925 143.640 73.185 144.365 ;
        RECT 73.355 143.470 73.600 144.195 ;
        RECT 73.785 143.640 74.045 144.365 ;
        RECT 74.215 143.470 74.460 144.195 ;
        RECT 74.630 143.640 74.890 144.365 ;
        RECT 75.060 143.470 75.320 144.195 ;
        RECT 75.490 143.640 75.750 144.365 ;
        RECT 75.920 143.470 76.180 144.195 ;
        RECT 76.350 143.640 76.610 144.365 ;
        RECT 76.780 143.470 77.040 144.195 ;
        RECT 77.210 143.640 77.470 144.365 ;
        RECT 77.640 143.470 77.900 144.265 ;
        RECT 78.070 143.640 78.320 144.775 ;
        RECT 71.625 143.465 77.900 143.470 ;
        RECT 78.500 143.465 78.760 144.275 ;
        RECT 78.935 143.635 79.180 144.775 ;
        RECT 79.360 143.465 79.655 144.275 ;
        RECT 79.835 143.465 80.125 144.630 ;
        RECT 81.225 143.465 81.520 144.275 ;
        RECT 81.700 143.635 81.945 144.775 ;
        RECT 82.120 143.465 82.380 144.275 ;
        RECT 82.560 143.640 82.810 144.775 ;
        RECT 88.990 144.605 90.155 145.195 ;
        RECT 83.410 144.380 90.155 144.605 ;
        RECT 90.505 145.195 97.250 145.365 ;
        RECT 90.505 144.605 91.670 145.195 ;
        RECT 97.850 145.025 98.100 145.835 ;
        RECT 98.280 145.490 98.540 146.015 ;
        RECT 98.710 145.025 98.960 145.835 ;
        RECT 99.140 145.505 99.445 146.015 ;
        RECT 91.840 144.775 98.960 145.025 ;
        RECT 99.130 144.775 99.445 145.335 ;
        RECT 99.625 145.205 99.895 146.015 ;
        RECT 100.065 145.205 100.395 145.845 ;
        RECT 100.565 145.205 100.805 146.015 ;
        RECT 101.000 145.635 103.015 145.805 ;
        RECT 103.205 145.635 103.535 146.015 ;
        RECT 101.000 145.315 101.255 145.635 ;
        RECT 99.615 144.775 99.965 145.025 ;
        RECT 90.505 144.380 97.250 144.605 ;
        RECT 83.410 144.365 88.815 144.380 ;
        RECT 82.980 143.470 83.240 144.265 ;
        RECT 83.410 143.640 83.670 144.365 ;
        RECT 83.840 143.470 84.100 144.195 ;
        RECT 84.270 143.640 84.530 144.365 ;
        RECT 84.700 143.470 84.960 144.195 ;
        RECT 85.130 143.640 85.390 144.365 ;
        RECT 85.560 143.470 85.820 144.195 ;
        RECT 85.990 143.640 86.250 144.365 ;
        RECT 86.420 143.470 86.665 144.195 ;
        RECT 86.835 143.640 87.095 144.365 ;
        RECT 87.280 143.470 87.525 144.195 ;
        RECT 87.695 143.640 87.955 144.365 ;
        RECT 88.140 143.470 88.385 144.195 ;
        RECT 88.555 143.640 88.815 144.365 ;
        RECT 89.000 143.470 89.255 144.195 ;
        RECT 89.425 143.640 89.715 144.380 ;
        RECT 82.980 143.465 89.255 143.470 ;
        RECT 89.885 143.465 90.155 144.210 ;
        RECT 90.505 143.465 90.775 144.210 ;
        RECT 90.945 143.640 91.235 144.380 ;
        RECT 91.845 144.365 97.250 144.380 ;
        RECT 91.405 143.470 91.660 144.195 ;
        RECT 91.845 143.640 92.105 144.365 ;
        RECT 92.275 143.470 92.520 144.195 ;
        RECT 92.705 143.640 92.965 144.365 ;
        RECT 93.135 143.470 93.380 144.195 ;
        RECT 93.565 143.640 93.825 144.365 ;
        RECT 93.995 143.470 94.240 144.195 ;
        RECT 94.410 143.640 94.670 144.365 ;
        RECT 94.840 143.470 95.100 144.195 ;
        RECT 95.270 143.640 95.530 144.365 ;
        RECT 95.700 143.470 95.960 144.195 ;
        RECT 96.130 143.640 96.390 144.365 ;
        RECT 96.560 143.470 96.820 144.195 ;
        RECT 96.990 143.640 97.250 144.365 ;
        RECT 97.420 143.470 97.680 144.265 ;
        RECT 97.850 143.640 98.100 144.775 ;
        RECT 91.405 143.465 97.680 143.470 ;
        RECT 98.280 143.465 98.540 144.275 ;
        RECT 98.715 143.635 98.960 144.775 ;
        RECT 100.135 144.605 100.305 145.205 ;
        RECT 100.475 144.775 100.825 145.025 ;
        RECT 101.000 144.775 101.240 145.105 ;
        RECT 101.425 144.655 101.755 145.465 ;
        RECT 102.265 145.195 103.955 145.465 ;
        RECT 104.125 145.215 104.505 146.015 ;
        RECT 105.595 145.290 105.885 146.015 ;
        RECT 101.980 144.825 103.070 145.025 ;
        RECT 103.380 144.825 104.505 145.025 ;
        RECT 99.140 143.465 99.435 144.275 ;
        RECT 99.625 143.465 99.955 144.605 ;
        RECT 100.135 144.435 100.815 144.605 ;
        RECT 100.485 143.650 100.815 144.435 ;
        RECT 101.000 143.465 101.255 144.605 ;
        RECT 101.425 144.435 103.955 144.655 ;
        RECT 101.425 143.635 101.755 144.435 ;
        RECT 101.925 143.465 102.095 144.265 ;
        RECT 102.265 143.635 102.595 144.435 ;
        RECT 102.765 143.465 103.455 144.265 ;
        RECT 103.625 143.635 103.955 144.435 ;
        RECT 104.125 143.465 104.505 144.655 ;
        RECT 105.595 143.465 105.885 144.630 ;
        RECT 106.070 143.645 106.350 145.835 ;
        RECT 106.550 145.645 107.280 146.015 ;
        RECT 107.860 145.475 108.290 145.835 ;
        RECT 106.550 145.285 108.290 145.475 ;
        RECT 106.550 144.775 106.810 145.285 ;
        RECT 106.540 143.465 106.825 144.605 ;
        RECT 107.020 144.485 107.280 145.105 ;
        RECT 107.475 144.485 107.900 145.105 ;
        RECT 108.070 145.055 108.290 145.285 ;
        RECT 108.460 145.235 108.705 146.015 ;
        RECT 108.070 144.755 108.615 145.055 ;
        RECT 108.905 144.935 109.135 145.835 ;
        RECT 107.090 144.115 108.115 144.315 ;
        RECT 107.090 143.645 107.260 144.115 ;
        RECT 107.435 143.465 107.765 143.945 ;
        RECT 107.935 143.645 108.115 144.115 ;
        RECT 108.285 143.645 108.615 144.755 ;
        RECT 108.795 144.255 109.135 144.935 ;
        RECT 109.315 144.435 109.545 145.775 ;
        RECT 109.775 145.195 110.005 146.015 ;
        RECT 110.175 145.215 110.505 145.845 ;
        RECT 109.755 144.775 110.085 145.025 ;
        RECT 110.255 144.615 110.505 145.215 ;
        RECT 110.675 145.195 110.885 146.015 ;
        RECT 111.205 145.535 111.505 146.015 ;
        RECT 111.675 145.365 111.935 145.820 ;
        RECT 112.105 145.535 112.365 146.015 ;
        RECT 112.545 145.365 112.805 145.820 ;
        RECT 112.975 145.535 113.225 146.015 ;
        RECT 113.405 145.365 113.665 145.820 ;
        RECT 113.835 145.535 114.085 146.015 ;
        RECT 114.265 145.365 114.525 145.820 ;
        RECT 114.695 145.535 114.940 146.015 ;
        RECT 115.110 145.365 115.385 145.820 ;
        RECT 115.555 145.535 115.800 146.015 ;
        RECT 115.970 145.365 116.230 145.820 ;
        RECT 116.400 145.535 116.660 146.015 ;
        RECT 116.830 145.365 117.090 145.820 ;
        RECT 117.260 145.535 117.520 146.015 ;
        RECT 117.690 145.365 117.950 145.820 ;
        RECT 118.120 145.455 118.380 146.015 ;
        RECT 111.205 145.195 117.950 145.365 ;
        RECT 108.795 144.055 109.545 144.255 ;
        RECT 108.785 143.465 109.135 143.875 ;
        RECT 109.305 143.665 109.545 144.055 ;
        RECT 109.775 143.465 110.005 144.605 ;
        RECT 110.175 143.635 110.505 144.615 ;
        RECT 111.205 144.605 112.370 145.195 ;
        RECT 118.550 145.025 118.800 145.835 ;
        RECT 118.980 145.490 119.240 146.015 ;
        RECT 119.410 145.025 119.660 145.835 ;
        RECT 119.840 145.505 120.145 146.015 ;
        RECT 120.315 145.535 120.575 146.015 ;
        RECT 120.745 145.765 120.990 145.845 ;
        RECT 120.745 145.595 121.075 145.765 ;
        RECT 112.540 144.775 119.660 145.025 ;
        RECT 119.830 144.775 120.145 145.335 ;
        RECT 120.360 144.775 120.555 145.345 ;
        RECT 110.675 143.465 110.885 144.605 ;
        RECT 111.205 144.380 117.950 144.605 ;
        RECT 111.205 143.465 111.475 144.210 ;
        RECT 111.645 143.640 111.935 144.380 ;
        RECT 112.545 144.365 117.950 144.380 ;
        RECT 112.105 143.470 112.360 144.195 ;
        RECT 112.545 143.640 112.805 144.365 ;
        RECT 112.975 143.470 113.220 144.195 ;
        RECT 113.405 143.640 113.665 144.365 ;
        RECT 113.835 143.470 114.080 144.195 ;
        RECT 114.265 143.640 114.525 144.365 ;
        RECT 114.695 143.470 114.940 144.195 ;
        RECT 115.110 143.640 115.370 144.365 ;
        RECT 115.540 143.470 115.800 144.195 ;
        RECT 115.970 143.640 116.230 144.365 ;
        RECT 116.400 143.470 116.660 144.195 ;
        RECT 116.830 143.640 117.090 144.365 ;
        RECT 117.260 143.470 117.520 144.195 ;
        RECT 117.690 143.640 117.950 144.365 ;
        RECT 118.120 143.470 118.380 144.265 ;
        RECT 118.550 143.640 118.800 144.775 ;
        RECT 112.105 143.465 118.380 143.470 ;
        RECT 118.980 143.465 119.240 144.275 ;
        RECT 119.415 143.635 119.660 144.775 ;
        RECT 120.745 144.605 120.915 145.595 ;
        RECT 121.275 145.400 121.485 145.685 ;
        RECT 121.750 145.675 121.920 145.700 ;
        RECT 121.750 145.505 121.925 145.675 ;
        RECT 122.165 145.635 122.495 146.015 ;
        RECT 122.685 145.675 122.855 145.845 ;
        RECT 122.265 145.555 122.435 145.635 ;
        RECT 122.675 145.505 122.855 145.675 ;
        RECT 123.105 145.555 123.360 146.015 ;
        RECT 121.750 145.405 121.920 145.505 ;
        RECT 121.095 145.230 121.485 145.400 ;
        RECT 121.655 145.235 121.920 145.405 ;
        RECT 122.685 145.385 122.855 145.505 ;
        RECT 121.095 145.165 121.375 145.230 ;
        RECT 121.095 144.775 121.265 145.165 ;
        RECT 121.655 145.025 121.825 145.235 ;
        RECT 122.180 145.105 122.385 145.340 ;
        RECT 122.685 145.215 123.360 145.385 ;
        RECT 123.995 145.265 125.205 146.015 ;
        RECT 121.495 144.855 121.825 145.025 ;
        RECT 121.655 144.840 121.825 144.855 ;
        RECT 122.055 144.775 122.385 145.105 ;
        RECT 122.565 144.855 122.895 145.025 ;
        RECT 122.725 144.605 122.895 144.855 ;
        RECT 120.405 144.435 122.895 144.605 ;
        RECT 119.840 143.465 120.135 144.275 ;
        RECT 120.405 143.635 120.575 144.435 ;
        RECT 123.105 144.265 123.360 145.215 ;
        RECT 120.805 144.095 122.095 144.265 ;
        RECT 120.865 143.675 121.115 144.095 ;
        RECT 121.305 143.465 121.635 143.925 ;
        RECT 121.845 143.675 122.095 144.095 ;
        RECT 122.265 143.465 122.515 144.265 ;
        RECT 122.685 144.095 123.360 144.265 ;
        RECT 123.995 144.555 124.515 145.095 ;
        RECT 124.685 144.725 125.205 145.265 ;
        RECT 122.685 143.635 122.855 144.095 ;
        RECT 123.065 143.465 123.315 143.925 ;
        RECT 123.995 143.465 125.205 144.555 ;
        RECT 53.990 143.295 125.290 143.465 ;
        RECT 54.075 142.205 55.285 143.295 ;
        RECT 54.075 141.495 54.595 142.035 ;
        RECT 54.765 141.665 55.285 142.205 ;
        RECT 56.465 142.365 56.635 143.125 ;
        RECT 56.850 142.535 57.180 143.295 ;
        RECT 56.465 142.195 57.180 142.365 ;
        RECT 57.350 142.220 57.605 143.125 ;
        RECT 56.375 141.645 56.730 142.015 ;
        RECT 57.010 141.985 57.180 142.195 ;
        RECT 57.010 141.655 57.265 141.985 ;
        RECT 54.075 140.745 55.285 141.495 ;
        RECT 57.010 141.465 57.180 141.655 ;
        RECT 57.435 141.490 57.605 142.220 ;
        RECT 57.780 142.145 58.040 143.295 ;
        RECT 58.220 142.145 58.480 143.295 ;
        RECT 58.655 142.220 58.910 143.125 ;
        RECT 59.080 142.535 59.410 143.295 ;
        RECT 59.625 142.365 59.795 143.125 ;
        RECT 56.465 141.295 57.180 141.465 ;
        RECT 56.465 140.915 56.635 141.295 ;
        RECT 56.850 140.745 57.180 141.125 ;
        RECT 57.350 140.915 57.605 141.490 ;
        RECT 57.780 140.745 58.040 141.585 ;
        RECT 58.220 140.745 58.480 141.585 ;
        RECT 58.655 141.490 58.825 142.220 ;
        RECT 59.080 142.195 59.795 142.365 ;
        RECT 59.080 141.985 59.250 142.195 ;
        RECT 60.975 142.155 61.255 143.295 ;
        RECT 61.425 142.145 61.755 143.125 ;
        RECT 61.925 142.155 62.185 143.295 ;
        RECT 62.555 142.625 62.835 143.295 ;
        RECT 63.005 142.405 63.305 142.955 ;
        RECT 63.505 142.575 63.835 143.295 ;
        RECT 64.025 142.575 64.485 143.125 ;
        RECT 58.995 141.655 59.250 141.985 ;
        RECT 58.655 140.915 58.910 141.490 ;
        RECT 59.080 141.465 59.250 141.655 ;
        RECT 59.530 141.645 59.885 142.015 ;
        RECT 60.985 141.715 61.320 141.985 ;
        RECT 61.490 141.545 61.660 142.145 ;
        RECT 62.370 141.985 62.635 142.345 ;
        RECT 63.005 142.235 63.945 142.405 ;
        RECT 63.775 141.985 63.945 142.235 ;
        RECT 61.830 141.735 62.165 141.985 ;
        RECT 62.370 141.735 63.045 141.985 ;
        RECT 63.265 141.735 63.605 141.985 ;
        RECT 63.775 141.655 64.065 141.985 ;
        RECT 63.775 141.565 63.945 141.655 ;
        RECT 59.080 141.295 59.795 141.465 ;
        RECT 59.080 140.745 59.410 141.125 ;
        RECT 59.625 140.915 59.795 141.295 ;
        RECT 60.975 140.745 61.285 141.545 ;
        RECT 61.490 140.915 62.185 141.545 ;
        RECT 62.555 141.375 63.945 141.565 ;
        RECT 62.555 141.015 62.885 141.375 ;
        RECT 64.235 141.205 64.485 142.575 ;
        RECT 64.675 142.495 64.955 143.295 ;
        RECT 65.155 142.325 65.485 143.125 ;
        RECT 65.685 142.495 65.855 143.295 ;
        RECT 66.025 142.325 66.355 143.125 ;
        RECT 64.655 141.655 64.895 142.325 ;
        RECT 65.075 142.155 66.355 142.325 ;
        RECT 66.525 142.155 66.785 143.295 ;
        RECT 65.075 141.485 65.245 142.155 ;
        RECT 66.955 142.130 67.245 143.295 ;
        RECT 67.415 142.220 67.685 143.125 ;
        RECT 67.855 142.535 68.185 143.295 ;
        RECT 68.365 142.365 68.535 143.125 ;
        RECT 65.415 141.655 65.725 141.985 ;
        RECT 65.895 141.655 66.275 141.985 ;
        RECT 66.475 141.655 66.760 141.985 ;
        RECT 65.520 141.485 65.725 141.655 ;
        RECT 63.505 140.745 63.755 141.205 ;
        RECT 63.925 140.915 64.485 141.205 ;
        RECT 64.655 140.915 65.350 141.485 ;
        RECT 65.520 140.960 65.870 141.485 ;
        RECT 66.060 140.960 66.275 141.655 ;
        RECT 66.445 140.745 66.780 141.485 ;
        RECT 66.955 140.745 67.245 141.470 ;
        RECT 67.415 141.420 67.585 142.220 ;
        RECT 67.870 142.195 68.535 142.365 ;
        RECT 68.815 142.405 69.075 143.115 ;
        RECT 69.245 142.585 69.575 143.295 ;
        RECT 69.745 142.405 69.975 143.115 ;
        RECT 67.870 142.050 68.040 142.195 ;
        RECT 68.815 142.165 69.975 142.405 ;
        RECT 70.155 142.385 70.425 143.115 ;
        RECT 70.605 142.565 70.945 143.295 ;
        RECT 70.155 142.165 70.925 142.385 ;
        RECT 67.755 141.720 68.040 142.050 ;
        RECT 67.870 141.465 68.040 141.720 ;
        RECT 68.275 141.645 68.605 142.015 ;
        RECT 68.805 141.655 69.105 141.985 ;
        RECT 69.285 141.675 69.810 141.985 ;
        RECT 69.990 141.675 70.455 141.985 ;
        RECT 67.415 140.915 67.675 141.420 ;
        RECT 67.870 141.295 68.535 141.465 ;
        RECT 67.855 140.745 68.185 141.125 ;
        RECT 68.365 140.915 68.535 141.295 ;
        RECT 68.815 140.745 69.105 141.475 ;
        RECT 69.285 141.035 69.515 141.675 ;
        RECT 70.635 141.495 70.925 142.165 ;
        RECT 69.695 141.295 70.925 141.495 ;
        RECT 69.695 140.925 70.005 141.295 ;
        RECT 70.185 140.745 70.855 141.115 ;
        RECT 71.115 140.925 71.375 143.115 ;
        RECT 71.555 142.325 71.865 143.125 ;
        RECT 72.035 142.495 72.345 143.295 ;
        RECT 72.515 142.665 72.775 143.125 ;
        RECT 72.945 142.835 73.200 143.295 ;
        RECT 73.375 142.665 73.635 143.125 ;
        RECT 72.515 142.495 73.635 142.665 ;
        RECT 71.555 142.155 72.585 142.325 ;
        RECT 71.555 141.245 71.725 142.155 ;
        RECT 71.895 141.415 72.245 141.985 ;
        RECT 72.415 141.905 72.585 142.155 ;
        RECT 73.375 142.245 73.635 142.495 ;
        RECT 73.805 142.425 74.090 143.295 ;
        RECT 74.405 142.550 74.675 143.295 ;
        RECT 75.305 143.290 81.580 143.295 ;
        RECT 74.845 142.380 75.135 143.120 ;
        RECT 75.305 142.565 75.560 143.290 ;
        RECT 75.745 142.395 76.005 143.120 ;
        RECT 76.175 142.565 76.420 143.290 ;
        RECT 76.605 142.395 76.865 143.120 ;
        RECT 77.035 142.565 77.280 143.290 ;
        RECT 77.465 142.395 77.725 143.120 ;
        RECT 77.895 142.565 78.140 143.290 ;
        RECT 78.310 142.395 78.570 143.120 ;
        RECT 78.740 142.565 79.000 143.290 ;
        RECT 79.170 142.395 79.430 143.120 ;
        RECT 79.600 142.565 79.860 143.290 ;
        RECT 80.030 142.395 80.290 143.120 ;
        RECT 80.460 142.565 80.720 143.290 ;
        RECT 80.890 142.395 81.150 143.120 ;
        RECT 81.320 142.495 81.580 143.290 ;
        RECT 75.745 142.380 81.150 142.395 ;
        RECT 73.375 142.075 74.130 142.245 ;
        RECT 72.415 141.735 73.555 141.905 ;
        RECT 73.725 141.565 74.130 142.075 ;
        RECT 72.480 141.395 74.130 141.565 ;
        RECT 74.405 142.155 81.150 142.380 ;
        RECT 74.405 141.565 75.570 142.155 ;
        RECT 81.750 141.985 82.000 143.120 ;
        RECT 82.180 142.485 82.440 143.295 ;
        RECT 82.615 141.985 82.860 143.125 ;
        RECT 83.040 142.485 83.335 143.295 ;
        RECT 83.605 142.550 83.875 143.295 ;
        RECT 84.505 143.290 90.780 143.295 ;
        RECT 84.045 142.380 84.335 143.120 ;
        RECT 84.505 142.565 84.760 143.290 ;
        RECT 84.945 142.395 85.205 143.120 ;
        RECT 85.375 142.565 85.620 143.290 ;
        RECT 85.805 142.395 86.065 143.120 ;
        RECT 86.235 142.565 86.480 143.290 ;
        RECT 86.665 142.395 86.925 143.120 ;
        RECT 87.095 142.565 87.340 143.290 ;
        RECT 87.510 142.395 87.770 143.120 ;
        RECT 87.940 142.565 88.200 143.290 ;
        RECT 88.370 142.395 88.630 143.120 ;
        RECT 88.800 142.565 89.060 143.290 ;
        RECT 89.230 142.395 89.490 143.120 ;
        RECT 89.660 142.565 89.920 143.290 ;
        RECT 90.090 142.395 90.350 143.120 ;
        RECT 90.520 142.495 90.780 143.290 ;
        RECT 84.945 142.380 90.350 142.395 ;
        RECT 83.605 142.155 90.350 142.380 ;
        RECT 75.740 141.735 82.860 141.985 ;
        RECT 74.405 141.395 81.150 141.565 ;
        RECT 71.555 140.915 71.855 141.245 ;
        RECT 72.025 140.745 72.300 141.225 ;
        RECT 72.480 141.005 72.775 141.395 ;
        RECT 72.945 140.745 73.200 141.225 ;
        RECT 73.375 141.005 73.635 141.395 ;
        RECT 73.805 140.745 74.085 141.225 ;
        RECT 74.405 140.745 74.705 141.225 ;
        RECT 74.875 140.940 75.135 141.395 ;
        RECT 75.305 140.745 75.565 141.225 ;
        RECT 75.745 140.940 76.005 141.395 ;
        RECT 76.175 140.745 76.425 141.225 ;
        RECT 76.605 140.940 76.865 141.395 ;
        RECT 77.035 140.745 77.285 141.225 ;
        RECT 77.465 140.940 77.725 141.395 ;
        RECT 77.895 140.745 78.140 141.225 ;
        RECT 78.310 140.940 78.585 141.395 ;
        RECT 78.755 140.745 79.000 141.225 ;
        RECT 79.170 140.940 79.430 141.395 ;
        RECT 79.600 140.745 79.860 141.225 ;
        RECT 80.030 140.940 80.290 141.395 ;
        RECT 80.460 140.745 80.720 141.225 ;
        RECT 80.890 140.940 81.150 141.395 ;
        RECT 81.320 140.745 81.580 141.305 ;
        RECT 81.750 140.925 82.000 141.735 ;
        RECT 82.180 140.745 82.440 141.270 ;
        RECT 82.610 140.925 82.860 141.735 ;
        RECT 83.030 141.425 83.345 141.985 ;
        RECT 83.605 141.565 84.770 142.155 ;
        RECT 90.950 141.985 91.200 143.120 ;
        RECT 91.380 142.485 91.640 143.295 ;
        RECT 91.815 141.985 92.060 143.125 ;
        RECT 92.240 142.485 92.535 143.295 ;
        RECT 92.715 142.130 93.005 143.295 ;
        RECT 93.175 142.325 93.465 143.125 ;
        RECT 93.635 142.495 93.870 143.295 ;
        RECT 94.055 142.955 95.590 143.125 ;
        RECT 94.055 142.325 94.385 142.955 ;
        RECT 93.175 142.155 94.385 142.325 ;
        RECT 84.940 141.735 92.060 141.985 ;
        RECT 83.605 141.395 90.350 141.565 ;
        RECT 83.040 140.745 83.345 141.255 ;
        RECT 83.605 140.745 83.905 141.225 ;
        RECT 84.075 140.940 84.335 141.395 ;
        RECT 84.505 140.745 84.765 141.225 ;
        RECT 84.945 140.940 85.205 141.395 ;
        RECT 85.375 140.745 85.625 141.225 ;
        RECT 85.805 140.940 86.065 141.395 ;
        RECT 86.235 140.745 86.485 141.225 ;
        RECT 86.665 140.940 86.925 141.395 ;
        RECT 87.095 140.745 87.340 141.225 ;
        RECT 87.510 140.940 87.785 141.395 ;
        RECT 87.955 140.745 88.200 141.225 ;
        RECT 88.370 140.940 88.630 141.395 ;
        RECT 88.800 140.745 89.060 141.225 ;
        RECT 89.230 140.940 89.490 141.395 ;
        RECT 89.660 140.745 89.920 141.225 ;
        RECT 90.090 140.940 90.350 141.395 ;
        RECT 90.520 140.745 90.780 141.305 ;
        RECT 90.950 140.925 91.200 141.735 ;
        RECT 91.380 140.745 91.640 141.270 ;
        RECT 91.810 140.925 92.060 141.735 ;
        RECT 92.230 141.425 92.545 141.985 ;
        RECT 93.175 141.655 93.420 141.985 ;
        RECT 93.590 141.485 93.760 142.155 ;
        RECT 94.555 141.985 94.790 142.730 ;
        RECT 93.930 141.655 94.330 141.985 ;
        RECT 94.500 141.655 94.790 141.985 ;
        RECT 94.980 141.985 95.250 142.730 ;
        RECT 95.420 142.325 95.590 142.955 ;
        RECT 95.760 142.495 96.155 143.295 ;
        RECT 95.420 142.155 96.155 142.325 ;
        RECT 94.980 141.655 95.310 141.985 ;
        RECT 95.480 141.655 95.815 141.985 ;
        RECT 95.985 141.655 96.155 142.155 ;
        RECT 96.325 141.975 96.680 143.125 ;
        RECT 96.850 142.145 97.145 143.295 ;
        RECT 97.325 142.155 97.655 143.295 ;
        RECT 98.185 142.325 98.515 143.110 ;
        RECT 98.705 142.485 99.000 143.295 ;
        RECT 97.835 142.155 98.515 142.325 ;
        RECT 96.325 141.715 97.145 141.975 ;
        RECT 97.315 141.735 97.665 141.985 ;
        RECT 96.325 141.655 96.680 141.715 ;
        RECT 92.240 140.745 92.545 141.255 ;
        RECT 92.715 140.745 93.005 141.470 ;
        RECT 93.175 140.915 93.760 141.485 ;
        RECT 94.010 141.315 95.395 141.485 ;
        RECT 94.010 140.970 94.340 141.315 ;
        RECT 94.555 140.745 94.930 141.145 ;
        RECT 95.110 140.970 95.395 141.315 ;
        RECT 95.565 140.745 96.235 141.485 ;
        RECT 96.405 140.915 96.680 141.655 ;
        RECT 97.835 141.555 98.005 142.155 ;
        RECT 99.180 141.985 99.425 143.125 ;
        RECT 99.600 142.485 99.860 143.295 ;
        RECT 100.460 143.290 106.735 143.295 ;
        RECT 100.040 141.985 100.290 143.120 ;
        RECT 100.460 142.495 100.720 143.290 ;
        RECT 100.890 142.395 101.150 143.120 ;
        RECT 101.320 142.565 101.580 143.290 ;
        RECT 101.750 142.395 102.010 143.120 ;
        RECT 102.180 142.565 102.440 143.290 ;
        RECT 102.610 142.395 102.870 143.120 ;
        RECT 103.040 142.565 103.300 143.290 ;
        RECT 103.470 142.395 103.730 143.120 ;
        RECT 103.900 142.565 104.145 143.290 ;
        RECT 104.315 142.395 104.575 143.120 ;
        RECT 104.760 142.565 105.005 143.290 ;
        RECT 105.175 142.395 105.435 143.120 ;
        RECT 105.620 142.565 105.865 143.290 ;
        RECT 106.035 142.395 106.295 143.120 ;
        RECT 106.480 142.565 106.735 143.290 ;
        RECT 100.890 142.380 106.295 142.395 ;
        RECT 106.905 142.380 107.195 143.120 ;
        RECT 107.365 142.550 107.635 143.295 ;
        RECT 107.905 142.485 108.200 143.295 ;
        RECT 100.890 142.155 107.635 142.380 ;
        RECT 98.175 141.735 98.525 141.985 ;
        RECT 96.850 140.745 97.145 141.545 ;
        RECT 97.325 140.745 97.595 141.555 ;
        RECT 97.765 140.915 98.095 141.555 ;
        RECT 98.265 140.745 98.505 141.555 ;
        RECT 98.695 141.425 99.010 141.985 ;
        RECT 99.180 141.735 106.300 141.985 ;
        RECT 98.695 140.745 99.000 141.255 ;
        RECT 99.180 140.925 99.430 141.735 ;
        RECT 99.600 140.745 99.860 141.270 ;
        RECT 100.040 140.925 100.290 141.735 ;
        RECT 106.470 141.565 107.635 142.155 ;
        RECT 108.380 141.985 108.625 143.125 ;
        RECT 108.800 142.485 109.060 143.295 ;
        RECT 109.660 143.290 115.935 143.295 ;
        RECT 109.240 141.985 109.490 143.120 ;
        RECT 109.660 142.495 109.920 143.290 ;
        RECT 110.090 142.395 110.350 143.120 ;
        RECT 110.520 142.565 110.780 143.290 ;
        RECT 110.950 142.395 111.210 143.120 ;
        RECT 111.380 142.565 111.640 143.290 ;
        RECT 111.810 142.395 112.070 143.120 ;
        RECT 112.240 142.565 112.500 143.290 ;
        RECT 112.670 142.395 112.930 143.120 ;
        RECT 113.100 142.565 113.345 143.290 ;
        RECT 113.515 142.395 113.775 143.120 ;
        RECT 113.960 142.565 114.205 143.290 ;
        RECT 114.375 142.395 114.635 143.120 ;
        RECT 114.820 142.565 115.065 143.290 ;
        RECT 115.235 142.395 115.495 143.120 ;
        RECT 115.680 142.565 115.935 143.290 ;
        RECT 110.090 142.380 115.495 142.395 ;
        RECT 116.105 142.380 116.395 143.120 ;
        RECT 116.565 142.550 116.835 143.295 ;
        RECT 110.090 142.155 116.835 142.380 ;
        RECT 117.185 142.365 117.355 143.125 ;
        RECT 117.535 142.535 117.865 143.295 ;
        RECT 117.185 142.195 117.850 142.365 ;
        RECT 118.035 142.220 118.305 143.125 ;
        RECT 100.890 141.395 107.635 141.565 ;
        RECT 107.895 141.425 108.210 141.985 ;
        RECT 108.380 141.735 115.500 141.985 ;
        RECT 100.460 140.745 100.720 141.305 ;
        RECT 100.890 140.940 101.150 141.395 ;
        RECT 101.320 140.745 101.580 141.225 ;
        RECT 101.750 140.940 102.010 141.395 ;
        RECT 102.180 140.745 102.440 141.225 ;
        RECT 102.610 140.940 102.870 141.395 ;
        RECT 103.040 140.745 103.285 141.225 ;
        RECT 103.455 140.940 103.730 141.395 ;
        RECT 103.900 140.745 104.145 141.225 ;
        RECT 104.315 140.940 104.575 141.395 ;
        RECT 104.755 140.745 105.005 141.225 ;
        RECT 105.175 140.940 105.435 141.395 ;
        RECT 105.615 140.745 105.865 141.225 ;
        RECT 106.035 140.940 106.295 141.395 ;
        RECT 106.475 140.745 106.735 141.225 ;
        RECT 106.905 140.940 107.165 141.395 ;
        RECT 107.335 140.745 107.635 141.225 ;
        RECT 107.895 140.745 108.200 141.255 ;
        RECT 108.380 140.925 108.630 141.735 ;
        RECT 108.800 140.745 109.060 141.270 ;
        RECT 109.240 140.925 109.490 141.735 ;
        RECT 115.670 141.565 116.835 142.155 ;
        RECT 117.680 142.050 117.850 142.195 ;
        RECT 117.115 141.645 117.445 142.015 ;
        RECT 117.680 141.720 117.965 142.050 ;
        RECT 110.090 141.395 116.835 141.565 ;
        RECT 117.680 141.465 117.850 141.720 ;
        RECT 109.660 140.745 109.920 141.305 ;
        RECT 110.090 140.940 110.350 141.395 ;
        RECT 110.520 140.745 110.780 141.225 ;
        RECT 110.950 140.940 111.210 141.395 ;
        RECT 111.380 140.745 111.640 141.225 ;
        RECT 111.810 140.940 112.070 141.395 ;
        RECT 112.240 140.745 112.485 141.225 ;
        RECT 112.655 140.940 112.930 141.395 ;
        RECT 113.100 140.745 113.345 141.225 ;
        RECT 113.515 140.940 113.775 141.395 ;
        RECT 113.955 140.745 114.205 141.225 ;
        RECT 114.375 140.940 114.635 141.395 ;
        RECT 114.815 140.745 115.065 141.225 ;
        RECT 115.235 140.940 115.495 141.395 ;
        RECT 115.675 140.745 115.935 141.225 ;
        RECT 116.105 140.940 116.365 141.395 ;
        RECT 117.185 141.295 117.850 141.465 ;
        RECT 118.135 141.420 118.305 142.220 ;
        RECT 118.475 142.130 118.765 143.295 ;
        RECT 118.935 142.155 119.265 143.295 ;
        RECT 119.435 142.665 119.790 143.125 ;
        RECT 119.960 142.835 120.535 143.295 ;
        RECT 120.705 142.665 121.035 143.125 ;
        RECT 119.435 142.495 121.035 142.665 ;
        RECT 121.235 142.495 121.490 143.295 ;
        RECT 119.435 142.155 119.710 142.495 ;
        RECT 119.890 141.935 120.080 142.315 ;
        RECT 118.935 141.735 120.080 141.935 ;
        RECT 120.260 141.595 120.540 142.495 ;
        RECT 121.660 142.325 121.960 142.520 ;
        RECT 120.710 142.155 121.960 142.325 ;
        RECT 122.245 142.365 122.415 143.125 ;
        RECT 122.630 142.535 122.960 143.295 ;
        RECT 122.245 142.195 122.960 142.365 ;
        RECT 123.130 142.220 123.385 143.125 ;
        RECT 120.710 141.735 121.040 142.155 ;
        RECT 121.270 141.655 121.615 141.985 ;
        RECT 120.260 141.565 120.545 141.595 ;
        RECT 116.535 140.745 116.835 141.225 ;
        RECT 117.185 140.915 117.355 141.295 ;
        RECT 117.535 140.745 117.865 141.125 ;
        RECT 118.045 140.915 118.305 141.420 ;
        RECT 118.475 140.745 118.765 141.470 ;
        RECT 118.935 141.355 120.045 141.565 ;
        RECT 118.935 140.915 119.285 141.355 ;
        RECT 119.455 140.745 119.625 141.185 ;
        RECT 119.795 141.125 120.045 141.355 ;
        RECT 120.215 141.295 120.545 141.565 ;
        RECT 120.715 141.125 120.990 141.565 ;
        RECT 121.790 141.500 121.960 142.155 ;
        RECT 122.155 141.645 122.510 142.015 ;
        RECT 122.790 141.985 122.960 142.195 ;
        RECT 122.790 141.655 123.045 141.985 ;
        RECT 119.795 140.915 120.990 141.125 ;
        RECT 121.225 140.745 121.555 141.485 ;
        RECT 121.725 141.170 121.960 141.500 ;
        RECT 122.790 141.465 122.960 141.655 ;
        RECT 123.215 141.490 123.385 142.220 ;
        RECT 123.560 142.145 123.820 143.295 ;
        RECT 123.995 142.205 125.205 143.295 ;
        RECT 123.995 141.665 124.515 142.205 ;
        RECT 122.245 141.295 122.960 141.465 ;
        RECT 122.245 140.915 122.415 141.295 ;
        RECT 122.630 140.745 122.960 141.125 ;
        RECT 123.130 140.915 123.385 141.490 ;
        RECT 123.560 140.745 123.820 141.585 ;
        RECT 124.685 141.495 125.205 142.035 ;
        RECT 123.995 140.745 125.205 141.495 ;
        RECT 53.990 140.575 125.290 140.745 ;
        RECT 54.075 139.825 55.285 140.575 ;
        RECT 54.075 139.285 54.595 139.825 ;
        RECT 55.460 139.735 55.720 140.575 ;
        RECT 55.895 139.830 56.150 140.405 ;
        RECT 56.320 140.195 56.650 140.575 ;
        RECT 56.865 140.025 57.035 140.405 ;
        RECT 56.320 139.855 57.035 140.025 ;
        RECT 54.765 139.115 55.285 139.655 ;
        RECT 54.075 138.025 55.285 139.115 ;
        RECT 55.460 138.025 55.720 139.175 ;
        RECT 55.895 139.100 56.065 139.830 ;
        RECT 56.320 139.665 56.490 139.855 ;
        RECT 56.235 139.335 56.490 139.665 ;
        RECT 56.320 139.125 56.490 139.335 ;
        RECT 56.770 139.305 57.125 139.675 ;
        RECT 55.895 138.195 56.150 139.100 ;
        RECT 56.320 138.955 57.035 139.125 ;
        RECT 56.320 138.025 56.650 138.785 ;
        RECT 56.865 138.195 57.035 138.955 ;
        RECT 57.755 138.195 58.505 140.405 ;
        RECT 58.765 140.025 58.935 140.405 ;
        RECT 59.115 140.195 59.445 140.575 ;
        RECT 58.765 139.855 59.430 140.025 ;
        RECT 59.625 139.900 59.885 140.405 ;
        RECT 58.695 139.305 59.035 139.675 ;
        RECT 59.260 139.600 59.430 139.855 ;
        RECT 59.260 139.270 59.535 139.600 ;
        RECT 59.260 139.125 59.430 139.270 ;
        RECT 58.755 138.955 59.430 139.125 ;
        RECT 59.705 139.100 59.885 139.900 ;
        RECT 58.755 138.195 58.935 138.955 ;
        RECT 59.115 138.025 59.445 138.785 ;
        RECT 59.615 138.195 59.885 139.100 ;
        RECT 60.060 140.100 60.395 140.360 ;
        RECT 60.565 140.175 60.895 140.575 ;
        RECT 61.065 140.175 62.680 140.345 ;
        RECT 60.060 138.745 60.315 140.100 ;
        RECT 61.065 140.005 61.235 140.175 ;
        RECT 60.675 139.835 61.235 140.005 ;
        RECT 60.675 139.665 60.845 139.835 ;
        RECT 60.540 139.335 60.845 139.665 ;
        RECT 61.040 139.555 61.290 139.665 ;
        RECT 61.500 139.555 61.770 139.995 ;
        RECT 61.960 139.895 62.250 139.995 ;
        RECT 61.955 139.725 62.250 139.895 ;
        RECT 61.035 139.385 61.290 139.555 ;
        RECT 61.495 139.385 61.770 139.555 ;
        RECT 61.040 139.335 61.290 139.385 ;
        RECT 61.500 139.335 61.770 139.385 ;
        RECT 61.960 139.335 62.250 139.725 ;
        RECT 62.420 139.335 62.840 140.000 ;
        RECT 63.225 139.855 63.555 140.575 ;
        RECT 63.150 139.335 63.500 139.665 ;
        RECT 60.675 139.165 60.845 139.335 ;
        RECT 63.295 139.215 63.500 139.335 ;
        RECT 63.735 139.630 64.075 140.405 ;
        RECT 64.245 140.115 64.415 140.575 ;
        RECT 64.655 140.140 65.015 140.405 ;
        RECT 64.655 140.135 65.010 140.140 ;
        RECT 64.655 140.125 65.005 140.135 ;
        RECT 64.655 140.120 65.000 140.125 ;
        RECT 64.655 140.110 64.995 140.120 ;
        RECT 65.645 140.115 65.815 140.575 ;
        RECT 64.655 140.105 64.990 140.110 ;
        RECT 64.655 140.095 64.980 140.105 ;
        RECT 64.655 140.085 64.970 140.095 ;
        RECT 64.655 139.945 64.955 140.085 ;
        RECT 64.245 139.755 64.955 139.945 ;
        RECT 65.145 139.945 65.475 140.025 ;
        RECT 65.985 139.945 66.325 140.405 ;
        RECT 65.145 139.755 66.325 139.945 ;
        RECT 66.530 139.835 67.145 140.405 ;
        RECT 67.315 140.065 67.530 140.575 ;
        RECT 67.760 140.065 68.040 140.395 ;
        RECT 68.220 140.065 68.460 140.575 ;
        RECT 60.675 138.995 63.045 139.165 ;
        RECT 63.295 139.045 63.505 139.215 ;
        RECT 60.060 138.235 60.395 138.745 ;
        RECT 60.645 138.025 60.975 138.825 ;
        RECT 61.220 138.615 62.645 138.785 ;
        RECT 61.220 138.195 61.505 138.615 ;
        RECT 61.760 138.025 62.090 138.445 ;
        RECT 62.315 138.365 62.645 138.615 ;
        RECT 62.875 138.535 63.045 138.995 ;
        RECT 63.305 138.365 63.475 138.865 ;
        RECT 62.315 138.195 63.475 138.365 ;
        RECT 63.735 138.195 64.015 139.630 ;
        RECT 64.245 139.185 64.530 139.755 ;
        RECT 64.715 139.355 65.185 139.585 ;
        RECT 65.355 139.565 65.685 139.585 ;
        RECT 65.355 139.385 65.805 139.565 ;
        RECT 65.995 139.385 66.325 139.585 ;
        RECT 64.245 138.970 65.395 139.185 ;
        RECT 64.185 138.025 64.895 138.800 ;
        RECT 65.065 138.195 65.395 138.970 ;
        RECT 65.590 138.270 65.805 139.385 ;
        RECT 66.095 139.045 66.325 139.385 ;
        RECT 66.530 138.815 66.845 139.835 ;
        RECT 67.015 139.165 67.185 139.665 ;
        RECT 67.435 139.335 67.700 139.895 ;
        RECT 67.870 139.165 68.040 140.065 ;
        RECT 68.210 139.335 68.565 139.895 ;
        RECT 68.800 139.810 69.255 140.575 ;
        RECT 69.530 140.195 70.830 140.405 ;
        RECT 71.085 140.215 71.415 140.575 ;
        RECT 70.660 140.045 70.830 140.195 ;
        RECT 71.585 140.075 71.845 140.405 ;
        RECT 69.730 139.585 69.950 139.985 ;
        RECT 68.795 139.385 69.285 139.585 ;
        RECT 69.475 139.375 69.950 139.585 ;
        RECT 70.195 139.585 70.405 139.985 ;
        RECT 70.660 139.920 71.415 140.045 ;
        RECT 70.660 139.875 71.505 139.920 ;
        RECT 71.235 139.755 71.505 139.875 ;
        RECT 70.195 139.375 70.525 139.585 ;
        RECT 70.695 139.315 71.105 139.620 ;
        RECT 67.015 138.995 68.440 139.165 ;
        RECT 65.985 138.025 66.315 138.745 ;
        RECT 66.530 138.195 67.065 138.815 ;
        RECT 67.235 138.025 67.565 138.825 ;
        RECT 68.050 138.820 68.440 138.995 ;
        RECT 68.800 139.145 69.975 139.205 ;
        RECT 71.335 139.180 71.505 139.755 ;
        RECT 71.305 139.145 71.505 139.180 ;
        RECT 68.800 139.035 71.505 139.145 ;
        RECT 68.800 138.415 69.055 139.035 ;
        RECT 69.645 138.975 71.445 139.035 ;
        RECT 69.645 138.945 69.975 138.975 ;
        RECT 71.675 138.875 71.845 140.075 ;
        RECT 69.305 138.775 69.490 138.865 ;
        RECT 70.080 138.775 70.915 138.785 ;
        RECT 69.305 138.575 70.915 138.775 ;
        RECT 69.305 138.535 69.535 138.575 ;
        RECT 68.800 138.195 69.135 138.415 ;
        RECT 70.140 138.025 70.495 138.405 ;
        RECT 70.665 138.195 70.915 138.575 ;
        RECT 71.165 138.025 71.415 138.805 ;
        RECT 71.585 138.195 71.845 138.875 ;
        RECT 72.015 140.075 72.275 140.405 ;
        RECT 72.445 140.215 72.775 140.575 ;
        RECT 73.030 140.195 74.330 140.405 ;
        RECT 72.015 138.875 72.185 140.075 ;
        RECT 73.030 140.045 73.200 140.195 ;
        RECT 72.445 139.920 73.200 140.045 ;
        RECT 72.355 139.875 73.200 139.920 ;
        RECT 72.355 139.755 72.625 139.875 ;
        RECT 72.355 139.180 72.525 139.755 ;
        RECT 72.755 139.315 73.165 139.620 ;
        RECT 73.455 139.585 73.665 139.985 ;
        RECT 73.335 139.375 73.665 139.585 ;
        RECT 73.910 139.585 74.130 139.985 ;
        RECT 74.605 139.810 75.060 140.575 ;
        RECT 75.235 139.775 75.930 140.405 ;
        RECT 76.135 139.775 76.445 140.575 ;
        RECT 76.625 139.850 76.955 140.360 ;
        RECT 77.125 140.175 77.455 140.575 ;
        RECT 78.505 140.005 78.835 140.345 ;
        RECT 79.005 140.175 79.335 140.575 ;
        RECT 73.910 139.375 74.385 139.585 ;
        RECT 74.575 139.385 75.065 139.585 ;
        RECT 75.255 139.335 75.590 139.585 ;
        RECT 72.355 139.145 72.555 139.180 ;
        RECT 73.885 139.145 75.060 139.205 ;
        RECT 75.760 139.175 75.930 139.775 ;
        RECT 76.100 139.335 76.435 139.605 ;
        RECT 72.355 139.035 75.060 139.145 ;
        RECT 72.415 138.975 74.215 139.035 ;
        RECT 73.885 138.945 74.215 138.975 ;
        RECT 72.015 138.195 72.275 138.875 ;
        RECT 72.445 138.025 72.695 138.805 ;
        RECT 72.945 138.775 73.780 138.785 ;
        RECT 74.370 138.775 74.555 138.865 ;
        RECT 72.945 138.575 74.555 138.775 ;
        RECT 72.945 138.195 73.195 138.575 ;
        RECT 74.325 138.535 74.555 138.575 ;
        RECT 74.805 138.415 75.060 139.035 ;
        RECT 73.365 138.025 73.720 138.405 ;
        RECT 74.725 138.195 75.060 138.415 ;
        RECT 75.235 138.025 75.495 139.165 ;
        RECT 75.665 138.195 75.995 139.175 ;
        RECT 76.165 138.025 76.445 139.165 ;
        RECT 76.625 139.085 76.815 139.850 ;
        RECT 77.125 139.835 79.490 140.005 ;
        RECT 79.835 139.850 80.125 140.575 ;
        RECT 77.125 139.665 77.295 139.835 ;
        RECT 76.985 139.335 77.295 139.665 ;
        RECT 77.465 139.335 77.770 139.665 ;
        RECT 76.625 138.235 76.955 139.085 ;
        RECT 77.125 138.025 77.375 139.165 ;
        RECT 77.555 139.005 77.770 139.335 ;
        RECT 77.945 139.005 78.230 139.665 ;
        RECT 78.425 139.005 78.690 139.665 ;
        RECT 78.905 139.005 79.150 139.665 ;
        RECT 79.320 138.835 79.490 139.835 ;
        RECT 80.295 139.835 80.615 140.210 ;
        RECT 80.870 139.835 81.040 140.575 ;
        RECT 81.290 140.005 81.460 140.210 ;
        RECT 81.705 140.175 82.060 140.575 ;
        RECT 82.235 140.005 82.405 140.355 ;
        RECT 82.605 140.175 82.935 140.575 ;
        RECT 83.105 140.005 83.275 140.355 ;
        RECT 83.445 140.175 83.825 140.575 ;
        RECT 81.290 139.835 81.810 140.005 ;
        RECT 82.235 139.835 83.845 140.005 ;
        RECT 84.015 139.900 84.290 140.245 ;
        RECT 77.565 138.665 78.855 138.835 ;
        RECT 77.565 138.245 77.815 138.665 ;
        RECT 78.045 138.025 78.375 138.495 ;
        RECT 78.605 138.245 78.855 138.665 ;
        RECT 79.035 138.665 79.490 138.835 ;
        RECT 79.035 138.235 79.365 138.665 ;
        RECT 79.835 138.025 80.125 139.190 ;
        RECT 80.295 138.795 80.470 139.835 ;
        RECT 80.640 138.965 80.990 139.665 ;
        RECT 81.160 139.335 81.450 139.665 ;
        RECT 81.620 139.585 81.810 139.835 ;
        RECT 83.675 139.665 83.845 139.835 ;
        RECT 81.620 139.415 82.065 139.585 ;
        RECT 81.620 139.135 81.810 139.415 ;
        RECT 82.460 139.245 82.630 139.665 ;
        RECT 82.850 139.335 83.505 139.665 ;
        RECT 83.675 139.335 83.950 139.665 ;
        RECT 81.205 138.965 81.810 139.135 ;
        RECT 81.980 139.075 82.630 139.245 ;
        RECT 83.675 139.165 83.845 139.335 ;
        RECT 84.120 139.165 84.290 139.900 ;
        RECT 84.460 139.635 84.630 140.575 ;
        RECT 84.905 140.235 85.240 140.405 ;
        RECT 84.905 139.835 85.520 140.235 ;
        RECT 86.200 140.195 86.535 140.575 ;
        RECT 87.125 140.135 87.360 140.575 ;
        RECT 87.530 140.045 87.860 140.405 ;
        RECT 88.030 140.215 88.360 140.575 ;
        RECT 88.575 140.065 88.880 140.575 ;
        RECT 85.690 139.835 86.960 140.025 ;
        RECT 87.530 139.875 88.350 140.045 ;
        RECT 84.895 139.335 85.170 139.665 ;
        RECT 81.980 138.795 82.150 139.075 ;
        RECT 83.185 138.995 83.845 139.165 ;
        RECT 83.185 138.875 83.355 138.995 ;
        RECT 80.295 138.625 82.150 138.795 ;
        RECT 82.320 138.705 83.355 138.875 ;
        RECT 80.295 138.205 80.555 138.625 ;
        RECT 82.320 138.455 82.490 138.705 ;
        RECT 80.725 138.025 81.055 138.455 ;
        RECT 81.745 138.285 82.490 138.455 ;
        RECT 82.715 138.205 83.355 138.535 ;
        RECT 83.525 138.025 83.805 138.825 ;
        RECT 84.015 138.195 84.290 139.165 ;
        RECT 84.460 138.025 84.630 139.220 ;
        RECT 85.340 139.150 85.520 139.835 ;
        RECT 85.690 139.335 86.050 139.665 ;
        RECT 86.340 139.555 86.630 139.665 ;
        RECT 86.335 139.385 86.630 139.555 ;
        RECT 86.340 139.335 86.630 139.385 ;
        RECT 86.800 139.335 87.135 139.665 ;
        RECT 87.305 139.335 87.985 139.665 ;
        RECT 87.305 139.150 87.475 139.335 ;
        RECT 84.900 138.895 87.475 139.150 ;
        RECT 84.900 138.195 85.165 138.895 ;
        RECT 85.335 138.025 85.665 138.725 ;
        RECT 85.835 138.195 86.505 138.895 ;
        RECT 88.155 138.755 88.350 139.875 ;
        RECT 88.575 139.335 88.890 139.895 ;
        RECT 89.060 139.585 89.310 140.395 ;
        RECT 89.480 140.050 89.740 140.575 ;
        RECT 89.920 139.585 90.170 140.395 ;
        RECT 90.340 140.015 90.600 140.575 ;
        RECT 90.770 139.925 91.030 140.380 ;
        RECT 91.200 140.095 91.460 140.575 ;
        RECT 91.630 139.925 91.890 140.380 ;
        RECT 92.060 140.095 92.320 140.575 ;
        RECT 92.490 139.925 92.750 140.380 ;
        RECT 92.920 140.095 93.165 140.575 ;
        RECT 93.335 139.925 93.610 140.380 ;
        RECT 93.780 140.095 94.025 140.575 ;
        RECT 94.195 139.925 94.455 140.380 ;
        RECT 94.635 140.095 94.885 140.575 ;
        RECT 95.055 139.925 95.315 140.380 ;
        RECT 95.495 140.095 95.745 140.575 ;
        RECT 95.915 139.925 96.175 140.380 ;
        RECT 96.355 140.095 96.615 140.575 ;
        RECT 96.785 139.925 97.045 140.380 ;
        RECT 97.215 140.095 97.515 140.575 ;
        RECT 97.775 140.235 99.135 140.405 ;
        RECT 90.770 139.755 97.515 139.925 ;
        RECT 97.775 139.755 98.135 140.235 ;
        RECT 98.305 139.835 98.635 140.065 ;
        RECT 98.805 140.005 99.135 140.235 ;
        RECT 99.305 140.175 99.635 140.575 ;
        RECT 99.805 140.005 100.135 140.405 ;
        RECT 98.805 139.835 100.135 140.005 ;
        RECT 100.405 139.835 100.735 140.575 ;
        RECT 89.060 139.335 96.180 139.585 ;
        RECT 87.010 138.025 87.440 138.725 ;
        RECT 87.620 138.585 88.350 138.755 ;
        RECT 87.620 138.195 87.810 138.585 ;
        RECT 87.980 138.025 88.310 138.405 ;
        RECT 88.585 138.025 88.880 138.835 ;
        RECT 89.060 138.195 89.305 139.335 ;
        RECT 89.480 138.025 89.740 138.835 ;
        RECT 89.920 138.200 90.170 139.335 ;
        RECT 96.350 139.165 97.515 139.755 ;
        RECT 97.775 139.415 98.135 139.585 ;
        RECT 97.775 139.335 98.105 139.415 ;
        RECT 90.770 138.940 97.515 139.165 ;
        RECT 90.770 138.925 96.175 138.940 ;
        RECT 90.340 138.030 90.600 138.825 ;
        RECT 90.770 138.200 91.030 138.925 ;
        RECT 91.200 138.030 91.460 138.755 ;
        RECT 91.630 138.200 91.890 138.925 ;
        RECT 92.060 138.030 92.320 138.755 ;
        RECT 92.490 138.200 92.750 138.925 ;
        RECT 92.920 138.030 93.180 138.755 ;
        RECT 93.350 138.200 93.610 138.925 ;
        RECT 93.780 138.030 94.025 138.755 ;
        RECT 94.195 138.200 94.455 138.925 ;
        RECT 94.640 138.030 94.885 138.755 ;
        RECT 95.055 138.200 95.315 138.925 ;
        RECT 95.500 138.030 95.745 138.755 ;
        RECT 95.915 138.200 96.175 138.925 ;
        RECT 96.360 138.030 96.615 138.755 ;
        RECT 96.785 138.200 97.075 138.940 ;
        RECT 90.340 138.025 96.615 138.030 ;
        RECT 97.245 138.025 97.515 138.770 ;
        RECT 97.775 138.025 98.135 139.165 ;
        RECT 98.305 138.875 98.505 139.835 ;
        RECT 98.675 139.555 98.920 139.665 ;
        RECT 98.675 139.385 98.925 139.555 ;
        RECT 98.675 139.045 98.920 139.385 ;
        RECT 99.195 139.045 99.415 139.665 ;
        RECT 99.670 139.045 99.845 139.665 ;
        RECT 100.115 139.045 100.335 139.665 ;
        RECT 100.505 138.875 100.815 139.665 ;
        RECT 98.305 138.705 100.815 138.875 ;
        RECT 98.805 138.195 99.135 138.705 ;
        RECT 100.305 138.025 100.815 138.535 ;
        RECT 100.985 138.195 101.315 140.405 ;
        RECT 101.485 139.775 101.745 140.575 ;
        RECT 102.095 140.195 102.425 140.575 ;
        RECT 102.595 140.025 102.785 140.405 ;
        RECT 102.955 140.215 103.285 140.575 ;
        RECT 102.385 139.835 102.785 140.025 ;
        RECT 103.505 140.005 103.695 140.405 ;
        RECT 102.955 139.835 103.695 140.005 ;
        RECT 101.485 138.025 101.745 139.165 ;
        RECT 101.925 138.025 102.215 138.995 ;
        RECT 102.385 138.195 102.615 139.835 ;
        RECT 102.955 139.665 103.125 139.835 ;
        RECT 102.785 138.970 103.125 139.665 ;
        RECT 103.295 139.250 103.620 139.665 ;
        RECT 104.070 139.335 104.450 140.295 ;
        RECT 104.635 140.095 104.965 140.575 ;
        RECT 104.640 139.335 104.955 139.910 ;
        RECT 105.595 139.850 105.885 140.575 ;
        RECT 106.055 140.065 106.360 140.575 ;
        RECT 106.055 139.335 106.370 139.895 ;
        RECT 106.540 139.585 106.790 140.395 ;
        RECT 106.960 140.050 107.220 140.575 ;
        RECT 107.400 139.585 107.650 140.395 ;
        RECT 107.820 140.015 108.080 140.575 ;
        RECT 108.250 139.925 108.510 140.380 ;
        RECT 108.680 140.095 108.940 140.575 ;
        RECT 109.110 139.925 109.370 140.380 ;
        RECT 109.540 140.095 109.800 140.575 ;
        RECT 109.970 139.925 110.230 140.380 ;
        RECT 110.400 140.095 110.645 140.575 ;
        RECT 110.815 139.925 111.090 140.380 ;
        RECT 111.260 140.095 111.505 140.575 ;
        RECT 111.675 139.925 111.935 140.380 ;
        RECT 112.115 140.095 112.365 140.575 ;
        RECT 112.535 139.925 112.795 140.380 ;
        RECT 112.975 140.095 113.225 140.575 ;
        RECT 113.395 139.925 113.655 140.380 ;
        RECT 113.835 140.095 114.095 140.575 ;
        RECT 114.265 139.925 114.525 140.380 ;
        RECT 114.695 140.095 114.995 140.575 ;
        RECT 108.250 139.755 114.995 139.925 ;
        RECT 115.255 139.755 115.550 140.575 ;
        RECT 115.720 139.835 116.160 140.395 ;
        RECT 116.330 139.835 116.780 140.575 ;
        RECT 116.950 140.005 117.120 140.405 ;
        RECT 117.290 140.175 117.710 140.575 ;
        RECT 117.880 140.005 118.110 140.405 ;
        RECT 116.950 139.835 118.110 140.005 ;
        RECT 118.280 139.835 118.765 140.405 ;
        RECT 106.540 139.335 113.660 139.585 ;
        RECT 102.785 138.740 103.620 138.970 ;
        RECT 102.785 138.025 103.115 138.440 ;
        RECT 103.305 138.195 103.620 138.740 ;
        RECT 103.790 138.725 104.905 138.990 ;
        RECT 103.790 138.195 104.015 138.725 ;
        RECT 104.185 138.025 104.515 138.535 ;
        RECT 104.685 138.195 104.905 138.725 ;
        RECT 105.595 138.025 105.885 139.190 ;
        RECT 106.065 138.025 106.360 138.835 ;
        RECT 106.540 138.195 106.785 139.335 ;
        RECT 106.960 138.025 107.220 138.835 ;
        RECT 107.400 138.200 107.650 139.335 ;
        RECT 113.830 139.165 114.995 139.755 ;
        RECT 115.720 139.585 116.030 139.835 ;
        RECT 115.255 139.365 116.030 139.585 ;
        RECT 108.250 138.940 114.995 139.165 ;
        RECT 108.250 138.925 113.655 138.940 ;
        RECT 107.820 138.030 108.080 138.825 ;
        RECT 108.250 138.200 108.510 138.925 ;
        RECT 108.680 138.030 108.940 138.755 ;
        RECT 109.110 138.200 109.370 138.925 ;
        RECT 109.540 138.030 109.800 138.755 ;
        RECT 109.970 138.200 110.230 138.925 ;
        RECT 110.400 138.030 110.660 138.755 ;
        RECT 110.830 138.200 111.090 138.925 ;
        RECT 111.260 138.030 111.505 138.755 ;
        RECT 111.675 138.200 111.935 138.925 ;
        RECT 112.120 138.030 112.365 138.755 ;
        RECT 112.535 138.200 112.795 138.925 ;
        RECT 112.980 138.030 113.225 138.755 ;
        RECT 113.395 138.200 113.655 138.925 ;
        RECT 113.840 138.030 114.095 138.755 ;
        RECT 114.265 138.200 114.555 138.940 ;
        RECT 107.820 138.025 114.095 138.030 ;
        RECT 114.725 138.025 114.995 138.770 ;
        RECT 115.255 138.025 115.550 139.195 ;
        RECT 115.720 138.825 116.030 139.365 ;
        RECT 116.200 139.215 116.370 139.665 ;
        RECT 116.540 139.385 116.930 139.665 ;
        RECT 117.115 139.335 117.360 139.665 ;
        RECT 116.200 139.045 116.990 139.215 ;
        RECT 115.720 138.195 116.160 138.825 ;
        RECT 116.335 138.025 116.650 138.875 ;
        RECT 116.820 138.365 116.990 139.045 ;
        RECT 117.160 138.535 117.360 139.335 ;
        RECT 117.560 138.535 117.810 139.665 ;
        RECT 118.025 139.335 118.425 139.665 ;
        RECT 118.595 139.165 118.765 139.835 ;
        RECT 118.935 139.755 119.230 140.575 ;
        RECT 119.400 139.835 119.840 140.395 ;
        RECT 120.010 139.835 120.460 140.575 ;
        RECT 120.630 140.005 120.800 140.405 ;
        RECT 120.970 140.175 121.390 140.575 ;
        RECT 121.560 140.005 121.790 140.405 ;
        RECT 120.630 139.835 121.790 140.005 ;
        RECT 121.960 139.835 122.445 140.405 ;
        RECT 119.400 139.585 119.710 139.835 ;
        RECT 118.935 139.365 119.710 139.585 ;
        RECT 118.000 138.995 118.765 139.165 ;
        RECT 118.000 138.365 118.250 138.995 ;
        RECT 116.820 138.195 118.250 138.365 ;
        RECT 118.425 138.025 118.760 138.825 ;
        RECT 118.935 138.025 119.230 139.195 ;
        RECT 119.400 138.825 119.710 139.365 ;
        RECT 119.880 139.215 120.050 139.665 ;
        RECT 120.220 139.385 120.610 139.665 ;
        RECT 120.795 139.335 121.040 139.665 ;
        RECT 119.880 139.045 120.670 139.215 ;
        RECT 119.400 138.195 119.840 138.825 ;
        RECT 120.015 138.025 120.330 138.875 ;
        RECT 120.500 138.365 120.670 139.045 ;
        RECT 120.840 138.535 121.040 139.335 ;
        RECT 121.240 138.535 121.490 139.665 ;
        RECT 121.705 139.335 122.105 139.665 ;
        RECT 122.275 139.165 122.445 139.835 ;
        RECT 121.680 138.995 122.445 139.165 ;
        RECT 122.615 139.900 122.875 140.405 ;
        RECT 123.055 140.195 123.385 140.575 ;
        RECT 123.565 140.025 123.735 140.405 ;
        RECT 122.615 139.100 122.795 139.900 ;
        RECT 123.070 139.855 123.735 140.025 ;
        RECT 123.070 139.600 123.240 139.855 ;
        RECT 123.995 139.825 125.205 140.575 ;
        RECT 122.965 139.270 123.240 139.600 ;
        RECT 123.465 139.305 123.805 139.675 ;
        RECT 123.070 139.125 123.240 139.270 ;
        RECT 121.680 138.365 121.930 138.995 ;
        RECT 120.500 138.195 121.930 138.365 ;
        RECT 122.105 138.025 122.440 138.825 ;
        RECT 122.615 138.195 122.885 139.100 ;
        RECT 123.070 138.955 123.745 139.125 ;
        RECT 123.055 138.025 123.385 138.785 ;
        RECT 123.565 138.195 123.745 138.955 ;
        RECT 123.995 139.115 124.515 139.655 ;
        RECT 124.685 139.285 125.205 139.825 ;
        RECT 123.995 138.025 125.205 139.115 ;
        RECT 53.990 137.855 125.290 138.025 ;
        RECT 54.075 136.765 55.285 137.855 ;
        RECT 54.075 136.055 54.595 136.595 ;
        RECT 54.765 136.225 55.285 136.765 ;
        RECT 55.915 136.715 56.205 137.855 ;
        RECT 56.375 137.135 56.825 137.685 ;
        RECT 57.015 137.135 57.345 137.855 ;
        RECT 54.075 135.305 55.285 136.055 ;
        RECT 55.915 135.305 56.205 136.105 ;
        RECT 56.375 135.765 56.625 137.135 ;
        RECT 57.555 136.965 57.855 137.515 ;
        RECT 58.025 137.185 58.305 137.855 ;
        RECT 56.915 136.795 57.855 136.965 ;
        RECT 56.915 136.545 57.085 136.795 ;
        RECT 58.190 136.545 58.505 136.985 ;
        RECT 58.860 136.885 59.250 137.060 ;
        RECT 59.735 137.055 60.065 137.855 ;
        RECT 60.235 137.065 60.770 137.685 ;
        RECT 58.860 136.715 60.285 136.885 ;
        RECT 56.795 136.215 57.085 136.545 ;
        RECT 57.255 136.295 57.585 136.545 ;
        RECT 57.815 136.295 58.505 136.545 ;
        RECT 56.915 136.125 57.085 136.215 ;
        RECT 56.915 135.935 58.305 136.125 ;
        RECT 58.735 135.985 59.090 136.545 ;
        RECT 56.375 135.475 56.925 135.765 ;
        RECT 57.095 135.305 57.345 135.765 ;
        RECT 57.975 135.575 58.305 135.935 ;
        RECT 59.260 135.815 59.430 136.715 ;
        RECT 59.600 135.985 59.865 136.545 ;
        RECT 60.115 136.215 60.285 136.715 ;
        RECT 60.455 136.045 60.770 137.065 ;
        RECT 61.065 137.515 62.225 137.685 ;
        RECT 61.065 137.015 61.235 137.515 ;
        RECT 61.495 136.885 61.665 137.345 ;
        RECT 61.895 137.265 62.225 137.515 ;
        RECT 62.450 137.435 62.780 137.855 ;
        RECT 63.035 137.265 63.320 137.685 ;
        RECT 61.895 137.095 63.320 137.265 ;
        RECT 63.565 137.055 63.895 137.855 ;
        RECT 64.145 137.135 64.480 137.645 ;
        RECT 61.040 136.545 61.245 136.835 ;
        RECT 61.495 136.715 63.865 136.885 ;
        RECT 63.695 136.545 63.865 136.715 ;
        RECT 61.040 136.495 61.390 136.545 ;
        RECT 61.035 136.325 61.390 136.495 ;
        RECT 61.040 136.215 61.390 136.325 ;
        RECT 58.840 135.305 59.080 135.815 ;
        RECT 59.260 135.485 59.540 135.815 ;
        RECT 59.770 135.305 59.985 135.815 ;
        RECT 60.155 135.475 60.770 136.045 ;
        RECT 60.985 135.305 61.315 136.025 ;
        RECT 61.700 135.880 62.120 136.545 ;
        RECT 62.290 135.885 62.580 136.545 ;
        RECT 62.770 136.495 63.040 136.545 ;
        RECT 63.250 136.495 63.500 136.545 ;
        RECT 62.770 136.325 63.045 136.495 ;
        RECT 63.250 136.325 63.505 136.495 ;
        RECT 62.770 135.885 63.040 136.325 ;
        RECT 63.250 136.215 63.500 136.325 ;
        RECT 63.695 136.215 64.000 136.545 ;
        RECT 63.695 136.045 63.865 136.215 ;
        RECT 63.305 135.875 63.865 136.045 ;
        RECT 63.305 135.705 63.475 135.875 ;
        RECT 64.225 135.780 64.480 137.135 ;
        RECT 61.860 135.535 63.475 135.705 ;
        RECT 63.645 135.305 63.975 135.705 ;
        RECT 64.145 135.520 64.480 135.780 ;
        RECT 65.575 136.780 65.845 137.685 ;
        RECT 66.015 137.095 66.345 137.855 ;
        RECT 66.525 136.925 66.695 137.685 ;
        RECT 65.575 135.980 65.745 136.780 ;
        RECT 66.030 136.755 66.695 136.925 ;
        RECT 66.030 136.610 66.200 136.755 ;
        RECT 66.955 136.690 67.245 137.855 ;
        RECT 67.415 136.715 67.675 137.855 ;
        RECT 67.845 136.705 68.175 137.685 ;
        RECT 68.345 136.715 68.625 137.855 ;
        RECT 68.800 136.715 69.120 137.855 ;
        RECT 65.915 136.280 66.200 136.610 ;
        RECT 66.030 136.025 66.200 136.280 ;
        RECT 66.435 136.205 66.765 136.575 ;
        RECT 67.435 136.295 67.770 136.545 ;
        RECT 67.940 136.105 68.110 136.705 ;
        RECT 69.300 136.545 69.495 137.595 ;
        RECT 69.675 137.005 70.005 137.685 ;
        RECT 70.205 137.055 70.460 137.855 ;
        RECT 69.675 136.725 70.025 137.005 ;
        RECT 68.280 136.275 68.615 136.545 ;
        RECT 68.860 136.495 69.120 136.545 ;
        RECT 68.855 136.325 69.120 136.495 ;
        RECT 68.860 136.215 69.120 136.325 ;
        RECT 69.300 136.215 69.685 136.545 ;
        RECT 69.855 136.345 70.025 136.725 ;
        RECT 70.215 136.515 70.460 136.875 ;
        RECT 70.790 136.845 71.090 137.685 ;
        RECT 71.285 137.015 71.535 137.855 ;
        RECT 72.125 137.265 72.930 137.685 ;
        RECT 71.705 137.095 73.270 137.265 ;
        RECT 71.705 136.845 71.875 137.095 ;
        RECT 70.790 136.675 71.875 136.845 ;
        RECT 69.855 136.175 70.375 136.345 ;
        RECT 70.635 136.215 70.965 136.505 ;
        RECT 65.575 135.475 65.835 135.980 ;
        RECT 66.030 135.855 66.695 136.025 ;
        RECT 66.015 135.305 66.345 135.685 ;
        RECT 66.525 135.475 66.695 135.855 ;
        RECT 66.955 135.305 67.245 136.030 ;
        RECT 67.415 135.475 68.110 136.105 ;
        RECT 68.315 135.305 68.625 136.105 ;
        RECT 68.800 135.835 70.015 136.005 ;
        RECT 68.800 135.485 69.090 135.835 ;
        RECT 69.285 135.305 69.615 135.665 ;
        RECT 69.785 135.530 70.015 135.835 ;
        RECT 70.205 135.610 70.375 136.175 ;
        RECT 71.135 136.045 71.305 136.675 ;
        RECT 72.045 136.545 72.365 136.925 ;
        RECT 71.475 136.295 71.805 136.505 ;
        RECT 71.985 136.295 72.365 136.545 ;
        RECT 72.555 136.505 72.930 136.925 ;
        RECT 73.100 136.845 73.270 137.095 ;
        RECT 73.440 137.015 73.770 137.855 ;
        RECT 73.940 137.095 74.605 137.685 ;
        RECT 73.100 136.675 74.020 136.845 ;
        RECT 73.850 136.505 74.020 136.675 ;
        RECT 72.555 136.495 73.040 136.505 ;
        RECT 72.535 136.325 73.040 136.495 ;
        RECT 72.555 136.295 73.040 136.325 ;
        RECT 73.230 136.295 73.680 136.505 ;
        RECT 73.850 136.295 74.185 136.505 ;
        RECT 74.355 136.125 74.605 137.095 ;
        RECT 75.240 137.465 75.575 137.685 ;
        RECT 76.580 137.475 76.935 137.855 ;
        RECT 75.240 136.845 75.495 137.465 ;
        RECT 75.745 137.305 75.975 137.345 ;
        RECT 77.105 137.305 77.355 137.685 ;
        RECT 75.745 137.105 77.355 137.305 ;
        RECT 75.745 137.015 75.930 137.105 ;
        RECT 76.520 137.095 77.355 137.105 ;
        RECT 77.605 137.075 77.855 137.855 ;
        RECT 78.025 137.005 78.285 137.685 ;
        RECT 78.545 137.110 78.815 137.855 ;
        RECT 79.445 137.850 85.720 137.855 ;
        RECT 76.085 136.905 76.415 136.935 ;
        RECT 76.085 136.845 77.885 136.905 ;
        RECT 75.240 136.735 77.945 136.845 ;
        RECT 75.240 136.675 76.415 136.735 ;
        RECT 77.745 136.700 77.945 136.735 ;
        RECT 75.235 136.295 75.725 136.495 ;
        RECT 75.915 136.295 76.390 136.505 ;
        RECT 70.795 135.865 71.305 136.045 ;
        RECT 71.710 135.955 73.410 136.125 ;
        RECT 71.710 135.865 72.095 135.955 ;
        RECT 70.795 135.475 71.125 135.865 ;
        RECT 71.295 135.525 72.480 135.695 ;
        RECT 72.740 135.305 72.910 135.775 ;
        RECT 73.080 135.490 73.410 135.955 ;
        RECT 73.580 135.305 73.750 136.125 ;
        RECT 73.920 135.485 74.605 136.125 ;
        RECT 75.240 135.305 75.695 136.070 ;
        RECT 76.170 135.895 76.390 136.295 ;
        RECT 76.635 136.295 76.965 136.505 ;
        RECT 76.635 135.895 76.845 136.295 ;
        RECT 77.135 136.260 77.545 136.565 ;
        RECT 77.775 136.125 77.945 136.700 ;
        RECT 77.675 136.005 77.945 136.125 ;
        RECT 77.100 135.960 77.945 136.005 ;
        RECT 77.100 135.835 77.855 135.960 ;
        RECT 77.100 135.685 77.270 135.835 ;
        RECT 78.115 135.805 78.285 137.005 ;
        RECT 78.985 136.940 79.275 137.680 ;
        RECT 79.445 137.125 79.700 137.850 ;
        RECT 79.885 136.955 80.145 137.680 ;
        RECT 80.315 137.125 80.560 137.850 ;
        RECT 80.745 136.955 81.005 137.680 ;
        RECT 81.175 137.125 81.420 137.850 ;
        RECT 81.605 136.955 81.865 137.680 ;
        RECT 82.035 137.125 82.280 137.850 ;
        RECT 82.450 136.955 82.710 137.680 ;
        RECT 82.880 137.125 83.140 137.850 ;
        RECT 83.310 136.955 83.570 137.680 ;
        RECT 83.740 137.125 84.000 137.850 ;
        RECT 84.170 136.955 84.430 137.680 ;
        RECT 84.600 137.125 84.860 137.850 ;
        RECT 85.030 136.955 85.290 137.680 ;
        RECT 85.460 137.055 85.720 137.850 ;
        RECT 79.885 136.940 85.290 136.955 ;
        RECT 78.545 136.715 85.290 136.940 ;
        RECT 78.545 136.125 79.710 136.715 ;
        RECT 85.890 136.545 86.140 137.680 ;
        RECT 86.320 137.045 86.580 137.855 ;
        RECT 86.755 136.545 87.000 137.685 ;
        RECT 87.180 137.045 87.475 137.855 ;
        RECT 87.655 136.715 87.915 137.855 ;
        RECT 79.880 136.295 87.000 136.545 ;
        RECT 78.545 135.955 85.290 136.125 ;
        RECT 75.970 135.475 77.270 135.685 ;
        RECT 77.525 135.305 77.855 135.665 ;
        RECT 78.025 135.475 78.285 135.805 ;
        RECT 78.545 135.305 78.845 135.785 ;
        RECT 79.015 135.500 79.275 135.955 ;
        RECT 79.445 135.305 79.705 135.785 ;
        RECT 79.885 135.500 80.145 135.955 ;
        RECT 80.315 135.305 80.565 135.785 ;
        RECT 80.745 135.500 81.005 135.955 ;
        RECT 81.175 135.305 81.425 135.785 ;
        RECT 81.605 135.500 81.865 135.955 ;
        RECT 82.035 135.305 82.280 135.785 ;
        RECT 82.450 135.500 82.725 135.955 ;
        RECT 82.895 135.305 83.140 135.785 ;
        RECT 83.310 135.500 83.570 135.955 ;
        RECT 83.740 135.305 84.000 135.785 ;
        RECT 84.170 135.500 84.430 135.955 ;
        RECT 84.600 135.305 84.860 135.785 ;
        RECT 85.030 135.500 85.290 135.955 ;
        RECT 85.460 135.305 85.720 135.865 ;
        RECT 85.890 135.485 86.140 136.295 ;
        RECT 86.320 135.305 86.580 135.830 ;
        RECT 86.750 135.485 87.000 136.295 ;
        RECT 87.170 135.985 87.485 136.545 ;
        RECT 87.180 135.305 87.485 135.815 ;
        RECT 87.655 135.305 87.915 136.105 ;
        RECT 88.085 135.475 88.415 137.685 ;
        RECT 88.585 137.345 89.095 137.855 ;
        RECT 90.265 137.175 90.595 137.685 ;
        RECT 88.585 137.005 91.095 137.175 ;
        RECT 88.585 136.215 88.895 137.005 ;
        RECT 89.065 136.215 89.285 136.835 ;
        RECT 89.555 136.215 89.730 136.835 ;
        RECT 89.985 136.215 90.205 136.835 ;
        RECT 90.475 136.665 90.725 136.835 ;
        RECT 90.480 136.215 90.725 136.665 ;
        RECT 90.895 136.045 91.095 137.005 ;
        RECT 91.265 136.715 91.625 137.855 ;
        RECT 92.715 136.690 93.005 137.855 ;
        RECT 93.265 137.110 93.535 137.855 ;
        RECT 94.165 137.850 100.440 137.855 ;
        RECT 93.705 136.940 93.995 137.680 ;
        RECT 94.165 137.125 94.420 137.850 ;
        RECT 94.605 136.955 94.865 137.680 ;
        RECT 95.035 137.125 95.280 137.850 ;
        RECT 95.465 136.955 95.725 137.680 ;
        RECT 95.895 137.125 96.140 137.850 ;
        RECT 96.325 136.955 96.585 137.680 ;
        RECT 96.755 137.125 97.000 137.850 ;
        RECT 97.170 136.955 97.430 137.680 ;
        RECT 97.600 137.125 97.860 137.850 ;
        RECT 98.030 136.955 98.290 137.680 ;
        RECT 98.460 137.125 98.720 137.850 ;
        RECT 98.890 136.955 99.150 137.680 ;
        RECT 99.320 137.125 99.580 137.850 ;
        RECT 99.750 136.955 100.010 137.680 ;
        RECT 100.180 137.055 100.440 137.850 ;
        RECT 94.605 136.940 100.010 136.955 ;
        RECT 93.265 136.715 100.010 136.940 ;
        RECT 91.295 136.465 91.625 136.545 ;
        RECT 91.265 136.295 91.625 136.465 ;
        RECT 93.265 136.155 94.430 136.715 ;
        RECT 100.610 136.545 100.860 137.680 ;
        RECT 101.040 137.045 101.300 137.855 ;
        RECT 101.475 136.545 101.720 137.685 ;
        RECT 101.900 137.045 102.195 137.855 ;
        RECT 102.465 136.885 102.635 137.685 ;
        RECT 102.925 137.225 103.175 137.645 ;
        RECT 103.365 137.395 103.695 137.855 ;
        RECT 103.905 137.225 104.155 137.645 ;
        RECT 102.865 137.055 104.155 137.225 ;
        RECT 104.325 137.055 104.575 137.855 ;
        RECT 104.745 137.225 104.915 137.685 ;
        RECT 105.125 137.395 105.375 137.855 ;
        RECT 104.745 137.055 105.420 137.225 ;
        RECT 102.465 136.715 104.955 136.885 ;
        RECT 94.600 136.295 101.720 136.545 ;
        RECT 93.235 136.125 94.430 136.155 ;
        RECT 88.665 135.305 88.995 136.045 ;
        RECT 89.265 135.875 90.595 136.045 ;
        RECT 89.265 135.475 89.595 135.875 ;
        RECT 89.765 135.305 90.095 135.705 ;
        RECT 90.265 135.645 90.595 135.875 ;
        RECT 90.765 135.815 91.095 136.045 ;
        RECT 91.265 135.645 91.625 136.125 ;
        RECT 90.265 135.475 91.625 135.645 ;
        RECT 92.715 135.305 93.005 136.030 ;
        RECT 93.235 135.985 100.010 136.125 ;
        RECT 93.265 135.955 100.010 135.985 ;
        RECT 93.265 135.305 93.565 135.785 ;
        RECT 93.735 135.500 93.995 135.955 ;
        RECT 94.165 135.305 94.425 135.785 ;
        RECT 94.605 135.500 94.865 135.955 ;
        RECT 95.035 135.305 95.285 135.785 ;
        RECT 95.465 135.500 95.725 135.955 ;
        RECT 95.895 135.305 96.145 135.785 ;
        RECT 96.325 135.500 96.585 135.955 ;
        RECT 96.755 135.305 97.000 135.785 ;
        RECT 97.170 135.500 97.445 135.955 ;
        RECT 97.615 135.305 97.860 135.785 ;
        RECT 98.030 135.500 98.290 135.955 ;
        RECT 98.460 135.305 98.720 135.785 ;
        RECT 98.890 135.500 99.150 135.955 ;
        RECT 99.320 135.305 99.580 135.785 ;
        RECT 99.750 135.500 100.010 135.955 ;
        RECT 100.180 135.305 100.440 135.865 ;
        RECT 100.610 135.485 100.860 136.295 ;
        RECT 101.040 135.305 101.300 135.830 ;
        RECT 101.470 135.485 101.720 136.295 ;
        RECT 101.890 135.985 102.205 136.545 ;
        RECT 102.420 135.975 102.615 136.545 ;
        RECT 101.900 135.305 102.205 135.815 ;
        RECT 102.375 135.305 102.635 135.785 ;
        RECT 102.805 135.725 102.975 136.715 ;
        RECT 103.155 136.090 103.325 136.545 ;
        RECT 103.715 136.465 103.885 136.480 ;
        RECT 103.555 136.295 103.885 136.465 ;
        RECT 103.155 135.920 103.545 136.090 ;
        RECT 102.805 135.555 103.135 135.725 ;
        RECT 103.335 135.635 103.545 135.920 ;
        RECT 103.715 136.085 103.885 136.295 ;
        RECT 104.115 136.215 104.445 136.545 ;
        RECT 104.785 136.465 104.955 136.715 ;
        RECT 104.625 136.295 104.955 136.465 ;
        RECT 103.715 135.915 103.980 136.085 ;
        RECT 104.240 135.980 104.445 136.215 ;
        RECT 105.165 136.105 105.420 137.055 ;
        RECT 105.600 136.710 105.895 137.855 ;
        RECT 103.810 135.815 103.980 135.915 ;
        RECT 104.745 135.935 105.420 136.105 ;
        RECT 103.810 135.645 103.985 135.815 ;
        RECT 104.325 135.685 104.495 135.765 ;
        RECT 103.810 135.620 103.980 135.645 ;
        RECT 102.805 135.475 103.050 135.555 ;
        RECT 104.225 135.305 104.555 135.685 ;
        RECT 104.745 135.475 104.915 135.935 ;
        RECT 105.165 135.305 105.420 135.765 ;
        RECT 105.600 135.305 105.895 136.125 ;
        RECT 106.065 135.855 106.295 137.555 ;
        RECT 106.510 137.050 106.765 137.855 ;
        RECT 106.965 137.240 107.295 137.685 ;
        RECT 107.465 137.410 107.740 137.855 ;
        RECT 107.975 137.240 108.305 137.685 ;
        RECT 106.965 137.060 108.305 137.240 ;
        RECT 108.765 136.880 109.095 137.545 ;
        RECT 109.365 137.110 109.635 137.855 ;
        RECT 110.265 137.850 116.540 137.855 ;
        RECT 109.805 136.940 110.095 137.680 ;
        RECT 110.265 137.125 110.520 137.850 ;
        RECT 110.705 136.955 110.965 137.680 ;
        RECT 111.135 137.125 111.380 137.850 ;
        RECT 111.565 136.955 111.825 137.680 ;
        RECT 111.995 137.125 112.240 137.850 ;
        RECT 112.425 136.955 112.685 137.680 ;
        RECT 112.855 137.125 113.100 137.850 ;
        RECT 113.270 136.955 113.530 137.680 ;
        RECT 113.700 137.125 113.960 137.850 ;
        RECT 114.130 136.955 114.390 137.680 ;
        RECT 114.560 137.125 114.820 137.850 ;
        RECT 114.990 136.955 115.250 137.680 ;
        RECT 115.420 137.125 115.680 137.850 ;
        RECT 115.850 136.955 116.110 137.680 ;
        RECT 116.280 137.055 116.540 137.850 ;
        RECT 110.705 136.940 116.110 136.955 ;
        RECT 106.510 136.710 109.095 136.880 ;
        RECT 109.365 136.715 116.110 136.940 ;
        RECT 106.510 136.095 106.820 136.710 ;
        RECT 106.990 136.265 107.320 136.495 ;
        RECT 107.490 136.265 107.960 136.495 ;
        RECT 108.130 136.325 108.585 136.495 ;
        RECT 108.130 136.265 108.580 136.325 ;
        RECT 108.770 136.265 109.105 136.495 ;
        RECT 109.365 136.125 110.530 136.715 ;
        RECT 116.710 136.545 116.960 137.680 ;
        RECT 117.140 137.045 117.400 137.855 ;
        RECT 117.575 136.545 117.820 137.685 ;
        RECT 118.000 137.045 118.295 137.855 ;
        RECT 118.475 136.690 118.765 137.855 ;
        RECT 118.955 137.265 119.195 137.655 ;
        RECT 119.365 137.445 119.715 137.855 ;
        RECT 118.955 137.065 119.705 137.265 ;
        RECT 110.700 136.295 117.820 136.545 ;
        RECT 106.510 135.915 109.095 136.095 ;
        RECT 109.365 135.955 116.110 136.125 ;
        RECT 106.065 135.475 106.285 135.855 ;
        RECT 106.455 135.305 107.305 135.665 ;
        RECT 107.785 135.495 108.115 135.915 ;
        RECT 108.320 135.305 108.595 135.745 ;
        RECT 108.765 135.495 109.095 135.915 ;
        RECT 109.365 135.305 109.665 135.785 ;
        RECT 109.835 135.500 110.095 135.955 ;
        RECT 110.265 135.305 110.525 135.785 ;
        RECT 110.705 135.500 110.965 135.955 ;
        RECT 111.135 135.305 111.385 135.785 ;
        RECT 111.565 135.500 111.825 135.955 ;
        RECT 111.995 135.305 112.245 135.785 ;
        RECT 112.425 135.500 112.685 135.955 ;
        RECT 112.855 135.305 113.100 135.785 ;
        RECT 113.270 135.500 113.545 135.955 ;
        RECT 113.715 135.305 113.960 135.785 ;
        RECT 114.130 135.500 114.390 135.955 ;
        RECT 114.560 135.305 114.820 135.785 ;
        RECT 114.990 135.500 115.250 135.955 ;
        RECT 115.420 135.305 115.680 135.785 ;
        RECT 115.850 135.500 116.110 135.955 ;
        RECT 116.280 135.305 116.540 135.865 ;
        RECT 116.710 135.485 116.960 136.295 ;
        RECT 117.140 135.305 117.400 135.830 ;
        RECT 117.570 135.485 117.820 136.295 ;
        RECT 117.990 135.985 118.305 136.545 ;
        RECT 118.000 135.305 118.305 135.815 ;
        RECT 118.475 135.305 118.765 136.030 ;
        RECT 118.955 135.545 119.185 136.885 ;
        RECT 119.365 136.385 119.705 137.065 ;
        RECT 119.885 136.565 120.215 137.675 ;
        RECT 120.385 137.205 120.565 137.675 ;
        RECT 120.735 137.375 121.065 137.855 ;
        RECT 121.240 137.205 121.410 137.675 ;
        RECT 120.385 137.005 121.410 137.205 ;
        RECT 119.365 135.485 119.595 136.385 ;
        RECT 119.885 136.265 120.430 136.565 ;
        RECT 119.795 135.305 120.040 136.085 ;
        RECT 120.210 136.035 120.430 136.265 ;
        RECT 120.600 136.215 121.025 136.835 ;
        RECT 121.220 136.215 121.480 136.835 ;
        RECT 121.675 136.715 121.960 137.855 ;
        RECT 121.690 136.035 121.950 136.545 ;
        RECT 120.210 135.845 121.950 136.035 ;
        RECT 120.210 135.485 120.640 135.845 ;
        RECT 121.220 135.305 121.950 135.675 ;
        RECT 122.150 135.485 122.430 137.675 ;
        RECT 122.655 136.715 122.885 137.855 ;
        RECT 123.055 136.705 123.385 137.685 ;
        RECT 123.555 136.715 123.765 137.855 ;
        RECT 123.995 136.765 125.205 137.855 ;
        RECT 122.635 136.295 122.965 136.545 ;
        RECT 122.655 135.305 122.885 136.125 ;
        RECT 123.135 136.105 123.385 136.705 ;
        RECT 123.995 136.225 124.515 136.765 ;
        RECT 123.055 135.475 123.385 136.105 ;
        RECT 123.555 135.305 123.765 136.125 ;
        RECT 124.685 136.055 125.205 136.595 ;
        RECT 123.995 135.305 125.205 136.055 ;
        RECT 53.990 135.135 125.290 135.305 ;
        RECT 54.075 134.385 55.285 135.135 ;
        RECT 54.075 133.845 54.595 134.385 ;
        RECT 55.460 134.295 55.720 135.135 ;
        RECT 55.895 134.390 56.150 134.965 ;
        RECT 56.320 134.755 56.650 135.135 ;
        RECT 56.865 134.585 57.035 134.965 ;
        RECT 56.320 134.415 57.035 134.585 ;
        RECT 57.385 134.585 57.555 134.965 ;
        RECT 57.735 134.755 58.065 135.135 ;
        RECT 57.385 134.415 58.050 134.585 ;
        RECT 58.245 134.460 58.505 134.965 ;
        RECT 54.765 133.675 55.285 134.215 ;
        RECT 54.075 132.585 55.285 133.675 ;
        RECT 55.460 132.585 55.720 133.735 ;
        RECT 55.895 133.660 56.065 134.390 ;
        RECT 56.320 134.225 56.490 134.415 ;
        RECT 56.235 133.895 56.490 134.225 ;
        RECT 56.320 133.685 56.490 133.895 ;
        RECT 56.770 133.865 57.125 134.235 ;
        RECT 57.315 133.865 57.655 134.235 ;
        RECT 57.880 134.160 58.050 134.415 ;
        RECT 57.880 133.830 58.155 134.160 ;
        RECT 57.880 133.685 58.050 133.830 ;
        RECT 55.895 132.755 56.150 133.660 ;
        RECT 56.320 133.515 57.035 133.685 ;
        RECT 56.320 132.585 56.650 133.345 ;
        RECT 56.865 132.755 57.035 133.515 ;
        RECT 57.375 133.515 58.050 133.685 ;
        RECT 58.325 133.660 58.505 134.460 ;
        RECT 57.375 132.755 57.555 133.515 ;
        RECT 57.735 132.585 58.065 133.345 ;
        RECT 58.235 132.755 58.505 133.660 ;
        RECT 58.675 134.460 58.935 134.965 ;
        RECT 59.115 134.755 59.445 135.135 ;
        RECT 59.625 134.585 59.795 134.965 ;
        RECT 58.675 133.660 58.845 134.460 ;
        RECT 59.130 134.415 59.795 134.585 ;
        RECT 59.130 134.160 59.300 134.415 ;
        RECT 60.115 134.315 60.325 135.135 ;
        RECT 60.495 134.335 60.825 134.965 ;
        RECT 59.015 133.830 59.300 134.160 ;
        RECT 59.535 133.865 59.865 134.235 ;
        RECT 59.130 133.685 59.300 133.830 ;
        RECT 60.495 133.735 60.745 134.335 ;
        RECT 60.995 134.315 61.225 135.135 ;
        RECT 60.915 133.895 61.245 134.145 ;
        RECT 58.675 132.755 58.945 133.660 ;
        RECT 59.130 133.515 59.795 133.685 ;
        RECT 59.115 132.585 59.445 133.345 ;
        RECT 59.625 132.755 59.795 133.515 ;
        RECT 60.115 132.585 60.325 133.725 ;
        RECT 60.495 132.755 60.825 133.735 ;
        RECT 60.995 132.585 61.225 133.725 ;
        RECT 61.905 132.765 62.165 134.955 ;
        RECT 62.425 134.765 63.095 135.135 ;
        RECT 63.275 134.585 63.585 134.955 ;
        RECT 62.355 134.385 63.585 134.585 ;
        RECT 62.355 133.715 62.645 134.385 ;
        RECT 63.765 134.205 63.995 134.845 ;
        RECT 64.175 134.405 64.465 135.135 ;
        RECT 64.690 134.395 65.305 134.965 ;
        RECT 65.475 134.625 65.690 135.135 ;
        RECT 65.920 134.625 66.200 134.955 ;
        RECT 66.380 134.625 66.620 135.135 ;
        RECT 62.825 133.895 63.290 134.205 ;
        RECT 63.470 133.895 63.995 134.205 ;
        RECT 64.175 133.895 64.475 134.225 ;
        RECT 62.355 133.495 63.125 133.715 ;
        RECT 62.335 132.585 62.675 133.315 ;
        RECT 62.855 132.765 63.125 133.495 ;
        RECT 63.305 133.475 64.465 133.715 ;
        RECT 63.305 132.765 63.535 133.475 ;
        RECT 63.705 132.585 64.035 133.295 ;
        RECT 64.205 132.765 64.465 133.475 ;
        RECT 64.690 133.375 65.005 134.395 ;
        RECT 65.175 133.725 65.345 134.225 ;
        RECT 65.595 133.895 65.860 134.455 ;
        RECT 66.030 133.725 66.200 134.625 ;
        RECT 67.505 134.585 67.675 134.965 ;
        RECT 67.855 134.755 68.185 135.135 ;
        RECT 66.370 133.895 66.725 134.455 ;
        RECT 67.505 134.415 68.170 134.585 ;
        RECT 68.365 134.460 68.625 134.965 ;
        RECT 67.435 133.865 67.775 134.235 ;
        RECT 68.000 134.160 68.170 134.415 ;
        RECT 68.000 133.830 68.275 134.160 ;
        RECT 65.175 133.555 66.600 133.725 ;
        RECT 68.000 133.685 68.170 133.830 ;
        RECT 64.690 132.755 65.225 133.375 ;
        RECT 65.395 132.585 65.725 133.385 ;
        RECT 66.210 133.380 66.600 133.555 ;
        RECT 67.495 133.515 68.170 133.685 ;
        RECT 68.445 133.660 68.625 134.460 ;
        RECT 68.805 134.405 69.105 135.135 ;
        RECT 69.285 134.225 69.515 134.845 ;
        RECT 69.715 134.575 69.940 134.955 ;
        RECT 70.110 134.745 70.440 135.135 ;
        RECT 71.555 134.675 72.115 134.965 ;
        RECT 72.285 134.675 72.535 135.135 ;
        RECT 69.715 134.395 70.045 134.575 ;
        RECT 68.810 133.895 69.105 134.225 ;
        RECT 69.285 133.895 69.700 134.225 ;
        RECT 69.870 133.725 70.045 134.395 ;
        RECT 70.215 133.895 70.455 134.545 ;
        RECT 67.495 132.755 67.675 133.515 ;
        RECT 67.855 132.585 68.185 133.345 ;
        RECT 68.355 132.755 68.625 133.660 ;
        RECT 68.805 133.365 69.700 133.695 ;
        RECT 69.870 133.535 70.455 133.725 ;
        RECT 68.805 133.195 70.010 133.365 ;
        RECT 68.805 132.765 69.135 133.195 ;
        RECT 69.315 132.585 69.510 133.025 ;
        RECT 69.680 132.765 70.010 133.195 ;
        RECT 70.180 132.765 70.455 133.535 ;
        RECT 71.555 133.305 71.805 134.675 ;
        RECT 73.155 134.505 73.485 134.865 ;
        RECT 73.860 134.630 74.195 135.135 ;
        RECT 74.365 134.565 74.605 134.940 ;
        RECT 74.885 134.805 75.055 134.950 ;
        RECT 74.885 134.610 75.260 134.805 ;
        RECT 75.620 134.640 76.015 135.135 ;
        RECT 72.095 134.315 73.485 134.505 ;
        RECT 72.095 134.225 72.265 134.315 ;
        RECT 71.975 133.895 72.265 134.225 ;
        RECT 72.435 133.895 72.775 134.145 ;
        RECT 72.995 133.895 73.670 134.145 ;
        RECT 72.095 133.645 72.265 133.895 ;
        RECT 72.095 133.475 73.035 133.645 ;
        RECT 73.405 133.535 73.670 133.895 ;
        RECT 73.915 133.605 74.215 134.455 ;
        RECT 74.385 134.415 74.605 134.565 ;
        RECT 74.385 134.085 74.920 134.415 ;
        RECT 75.090 134.275 75.260 134.610 ;
        RECT 76.185 134.445 76.425 134.965 ;
        RECT 77.075 134.755 77.405 135.135 ;
        RECT 71.555 132.755 72.015 133.305 ;
        RECT 72.205 132.585 72.535 133.305 ;
        RECT 72.735 132.925 73.035 133.475 ;
        RECT 74.385 133.435 74.620 134.085 ;
        RECT 75.090 133.915 76.075 134.275 ;
        RECT 73.205 132.585 73.485 133.255 ;
        RECT 73.945 133.205 74.620 133.435 ;
        RECT 74.790 133.895 76.075 133.915 ;
        RECT 74.790 133.745 75.650 133.895 ;
        RECT 73.945 132.775 74.115 133.205 ;
        RECT 74.285 132.585 74.615 133.035 ;
        RECT 74.790 132.800 75.075 133.745 ;
        RECT 76.250 133.640 76.425 134.445 ;
        RECT 76.630 134.585 76.905 134.725 ;
        RECT 77.575 134.585 77.785 134.755 ;
        RECT 76.630 134.395 77.785 134.585 ;
        RECT 77.955 134.585 78.285 134.965 ;
        RECT 78.475 134.755 78.805 135.135 ;
        RECT 77.955 134.380 78.805 134.585 ;
        RECT 76.625 133.770 76.885 134.225 ;
        RECT 77.140 133.820 77.725 134.195 ;
        RECT 75.250 133.265 75.945 133.575 ;
        RECT 75.255 132.585 75.940 133.055 ;
        RECT 76.120 132.855 76.425 133.640 ;
        RECT 76.630 132.585 76.955 133.570 ;
        RECT 77.140 133.435 77.345 133.820 ;
        RECT 77.895 133.605 78.305 134.210 ;
        RECT 78.475 133.890 78.805 134.380 ;
        RECT 78.475 133.435 78.645 133.890 ;
        RECT 77.135 133.265 77.345 133.435 ;
        RECT 77.140 133.235 77.345 133.265 ;
        RECT 77.525 133.215 78.645 133.435 ;
        RECT 77.525 132.755 77.785 133.215 ;
        RECT 77.955 132.585 78.805 133.035 ;
        RECT 78.975 132.755 79.220 134.965 ;
        RECT 79.405 134.335 79.645 135.135 ;
        RECT 79.835 134.410 80.125 135.135 ;
        RECT 80.295 134.635 80.555 134.965 ;
        RECT 80.725 134.775 81.055 135.135 ;
        RECT 81.310 134.755 82.610 134.965 ;
        RECT 79.405 132.585 79.660 133.585 ;
        RECT 79.835 132.585 80.125 133.750 ;
        RECT 80.295 133.435 80.465 134.635 ;
        RECT 81.310 134.605 81.480 134.755 ;
        RECT 80.725 134.480 81.480 134.605 ;
        RECT 80.635 134.435 81.480 134.480 ;
        RECT 80.635 134.315 80.905 134.435 ;
        RECT 80.635 133.740 80.805 134.315 ;
        RECT 81.035 133.875 81.445 134.180 ;
        RECT 81.735 134.145 81.945 134.545 ;
        RECT 81.615 133.935 81.945 134.145 ;
        RECT 82.190 134.145 82.410 134.545 ;
        RECT 82.885 134.370 83.340 135.135 ;
        RECT 82.190 133.935 82.665 134.145 ;
        RECT 82.855 133.945 83.345 134.145 ;
        RECT 80.635 133.705 80.835 133.740 ;
        RECT 82.165 133.705 83.340 133.765 ;
        RECT 80.635 133.595 83.340 133.705 ;
        RECT 80.695 133.535 82.495 133.595 ;
        RECT 82.165 133.505 82.495 133.535 ;
        RECT 80.295 132.755 80.555 133.435 ;
        RECT 80.725 132.585 80.975 133.365 ;
        RECT 81.225 133.335 82.060 133.345 ;
        RECT 82.650 133.335 82.835 133.425 ;
        RECT 81.225 133.135 82.835 133.335 ;
        RECT 81.225 132.755 81.475 133.135 ;
        RECT 82.605 133.095 82.835 133.135 ;
        RECT 83.085 132.975 83.340 133.595 ;
        RECT 81.645 132.585 82.000 132.965 ;
        RECT 83.005 132.755 83.340 132.975 ;
        RECT 83.515 132.755 83.795 134.855 ;
        RECT 84.025 134.675 84.195 135.135 ;
        RECT 84.465 134.745 85.715 134.925 ;
        RECT 84.850 134.505 85.215 134.575 ;
        RECT 83.965 134.325 85.215 134.505 ;
        RECT 85.385 134.525 85.715 134.745 ;
        RECT 85.885 134.695 86.055 135.135 ;
        RECT 86.225 134.525 86.565 134.940 ;
        RECT 86.825 134.655 87.125 135.135 ;
        RECT 85.385 134.355 86.565 134.525 ;
        RECT 87.295 134.485 87.555 134.940 ;
        RECT 87.725 134.655 87.985 135.135 ;
        RECT 88.165 134.485 88.425 134.940 ;
        RECT 88.595 134.655 88.845 135.135 ;
        RECT 89.025 134.485 89.285 134.940 ;
        RECT 89.455 134.655 89.705 135.135 ;
        RECT 89.885 134.485 90.145 134.940 ;
        RECT 90.315 134.655 90.560 135.135 ;
        RECT 90.730 134.485 91.005 134.940 ;
        RECT 91.175 134.655 91.420 135.135 ;
        RECT 91.590 134.485 91.850 134.940 ;
        RECT 92.020 134.655 92.280 135.135 ;
        RECT 92.450 134.485 92.710 134.940 ;
        RECT 92.880 134.655 93.140 135.135 ;
        RECT 93.310 134.485 93.570 134.940 ;
        RECT 93.740 134.575 94.000 135.135 ;
        RECT 83.965 133.725 84.240 134.325 ;
        RECT 86.825 134.315 93.570 134.485 ;
        RECT 84.410 133.895 84.765 134.145 ;
        RECT 84.960 134.115 85.425 134.145 ;
        RECT 84.955 133.945 85.425 134.115 ;
        RECT 84.960 133.895 85.425 133.945 ;
        RECT 85.595 133.895 85.925 134.145 ;
        RECT 86.100 133.945 86.565 134.145 ;
        RECT 85.745 133.775 85.925 133.895 ;
        RECT 83.965 133.515 85.575 133.725 ;
        RECT 85.745 133.605 86.075 133.775 ;
        RECT 85.165 133.415 85.575 133.515 ;
        RECT 83.985 132.585 84.770 133.345 ;
        RECT 85.165 132.755 85.550 133.415 ;
        RECT 85.875 132.815 86.075 133.605 ;
        RECT 86.245 132.585 86.565 133.765 ;
        RECT 86.825 133.725 87.990 134.315 ;
        RECT 94.170 134.145 94.420 134.955 ;
        RECT 94.600 134.610 94.860 135.135 ;
        RECT 95.030 134.145 95.280 134.955 ;
        RECT 95.460 134.625 95.765 135.135 ;
        RECT 96.485 134.655 96.785 135.135 ;
        RECT 96.955 134.485 97.215 134.940 ;
        RECT 97.385 134.655 97.645 135.135 ;
        RECT 97.825 134.485 98.085 134.940 ;
        RECT 98.255 134.655 98.505 135.135 ;
        RECT 98.685 134.485 98.945 134.940 ;
        RECT 99.115 134.655 99.365 135.135 ;
        RECT 99.545 134.485 99.805 134.940 ;
        RECT 99.975 134.655 100.220 135.135 ;
        RECT 100.390 134.485 100.665 134.940 ;
        RECT 100.835 134.655 101.080 135.135 ;
        RECT 101.250 134.485 101.510 134.940 ;
        RECT 101.680 134.655 101.940 135.135 ;
        RECT 102.110 134.485 102.370 134.940 ;
        RECT 102.540 134.655 102.800 135.135 ;
        RECT 102.970 134.485 103.230 134.940 ;
        RECT 103.400 134.575 103.660 135.135 ;
        RECT 88.160 133.895 95.280 134.145 ;
        RECT 95.450 133.895 95.765 134.455 ;
        RECT 96.485 134.315 103.230 134.485 ;
        RECT 86.825 133.500 93.570 133.725 ;
        RECT 86.825 132.585 87.095 133.330 ;
        RECT 87.265 132.760 87.555 133.500 ;
        RECT 88.165 133.485 93.570 133.500 ;
        RECT 87.725 132.590 87.980 133.315 ;
        RECT 88.165 132.760 88.425 133.485 ;
        RECT 88.595 132.590 88.840 133.315 ;
        RECT 89.025 132.760 89.285 133.485 ;
        RECT 89.455 132.590 89.700 133.315 ;
        RECT 89.885 132.760 90.145 133.485 ;
        RECT 90.315 132.590 90.560 133.315 ;
        RECT 90.730 132.760 90.990 133.485 ;
        RECT 91.160 132.590 91.420 133.315 ;
        RECT 91.590 132.760 91.850 133.485 ;
        RECT 92.020 132.590 92.280 133.315 ;
        RECT 92.450 132.760 92.710 133.485 ;
        RECT 92.880 132.590 93.140 133.315 ;
        RECT 93.310 132.760 93.570 133.485 ;
        RECT 93.740 132.590 94.000 133.385 ;
        RECT 94.170 132.760 94.420 133.895 ;
        RECT 87.725 132.585 94.000 132.590 ;
        RECT 94.600 132.585 94.860 133.395 ;
        RECT 95.035 132.755 95.280 133.895 ;
        RECT 96.485 133.725 97.650 134.315 ;
        RECT 103.830 134.145 104.080 134.955 ;
        RECT 104.260 134.610 104.520 135.135 ;
        RECT 104.690 134.145 104.940 134.955 ;
        RECT 105.120 134.625 105.425 135.135 ;
        RECT 97.820 133.895 104.940 134.145 ;
        RECT 105.110 133.895 105.425 134.455 ;
        RECT 105.595 134.410 105.885 135.135 ;
        RECT 106.055 134.485 106.315 134.930 ;
        RECT 106.565 134.655 106.735 135.135 ;
        RECT 106.905 134.625 107.255 134.955 ;
        RECT 107.490 134.655 107.660 135.135 ;
        RECT 106.055 134.315 106.735 134.485 ;
        RECT 96.485 133.500 103.230 133.725 ;
        RECT 95.460 132.585 95.755 133.395 ;
        RECT 96.485 132.585 96.755 133.330 ;
        RECT 96.925 132.760 97.215 133.500 ;
        RECT 97.825 133.485 103.230 133.500 ;
        RECT 97.385 132.590 97.640 133.315 ;
        RECT 97.825 132.760 98.085 133.485 ;
        RECT 98.255 132.590 98.500 133.315 ;
        RECT 98.685 132.760 98.945 133.485 ;
        RECT 99.115 132.590 99.360 133.315 ;
        RECT 99.545 132.760 99.805 133.485 ;
        RECT 99.975 132.590 100.220 133.315 ;
        RECT 100.390 132.760 100.650 133.485 ;
        RECT 100.820 132.590 101.080 133.315 ;
        RECT 101.250 132.760 101.510 133.485 ;
        RECT 101.680 132.590 101.940 133.315 ;
        RECT 102.110 132.760 102.370 133.485 ;
        RECT 102.540 132.590 102.800 133.315 ;
        RECT 102.970 132.760 103.230 133.485 ;
        RECT 103.400 132.590 103.660 133.385 ;
        RECT 103.830 132.760 104.080 133.895 ;
        RECT 97.385 132.585 103.660 132.590 ;
        RECT 104.260 132.585 104.520 133.395 ;
        RECT 104.695 132.755 104.940 133.895 ;
        RECT 105.120 132.585 105.415 133.395 ;
        RECT 105.595 132.585 105.885 133.750 ;
        RECT 106.055 133.580 106.395 134.145 ;
        RECT 106.565 133.410 106.735 134.315 ;
        RECT 106.905 133.725 107.075 134.625 ;
        RECT 107.960 134.565 108.130 134.915 ;
        RECT 108.300 134.735 108.630 135.135 ;
        RECT 108.800 134.615 109.055 134.915 ;
        RECT 108.800 134.565 109.105 134.615 ;
        RECT 107.960 134.485 109.105 134.565 ;
        RECT 107.395 134.455 109.105 134.485 ;
        RECT 107.245 134.395 109.105 134.455 ;
        RECT 107.245 134.315 108.130 134.395 ;
        RECT 107.245 134.285 107.565 134.315 ;
        RECT 107.245 133.895 107.415 134.285 ;
        RECT 106.905 133.520 107.300 133.725 ;
        RECT 107.665 133.605 108.200 134.145 ;
        RECT 108.460 133.895 108.760 134.225 ;
        RECT 108.460 133.435 108.630 133.895 ;
        RECT 108.935 133.725 109.105 134.395 ;
        RECT 109.735 134.335 109.995 135.135 ;
        RECT 106.055 133.350 106.735 133.410 ;
        RECT 107.520 133.350 108.630 133.435 ;
        RECT 106.055 133.265 108.630 133.350 ;
        RECT 108.800 133.295 109.105 133.725 ;
        RECT 106.055 133.180 107.690 133.265 ;
        RECT 106.055 133.000 106.315 133.180 ;
        RECT 106.520 132.585 106.880 133.010 ;
        RECT 107.395 132.585 107.725 133.010 ;
        RECT 107.905 132.855 109.105 133.095 ;
        RECT 109.735 132.585 109.995 133.725 ;
        RECT 110.165 132.755 110.495 134.965 ;
        RECT 110.745 134.395 111.075 135.135 ;
        RECT 111.345 134.565 111.675 134.965 ;
        RECT 111.845 134.735 112.175 135.135 ;
        RECT 112.345 134.795 113.705 134.965 ;
        RECT 112.345 134.565 112.675 134.795 ;
        RECT 111.345 134.395 112.675 134.565 ;
        RECT 112.845 134.395 113.175 134.625 ;
        RECT 110.665 133.435 110.975 134.225 ;
        RECT 111.145 133.605 111.365 134.225 ;
        RECT 111.635 133.605 111.810 134.225 ;
        RECT 112.065 133.605 112.285 134.225 ;
        RECT 112.560 134.115 112.805 134.225 ;
        RECT 112.555 133.945 112.805 134.115 ;
        RECT 112.560 133.605 112.805 133.945 ;
        RECT 112.975 133.435 113.175 134.395 ;
        RECT 113.345 134.315 113.705 134.795 ;
        RECT 114.885 134.655 115.185 135.135 ;
        RECT 115.355 134.485 115.615 134.940 ;
        RECT 115.785 134.655 116.045 135.135 ;
        RECT 116.225 134.485 116.485 134.940 ;
        RECT 116.655 134.655 116.905 135.135 ;
        RECT 117.085 134.485 117.345 134.940 ;
        RECT 117.515 134.655 117.765 135.135 ;
        RECT 117.945 134.485 118.205 134.940 ;
        RECT 118.375 134.655 118.620 135.135 ;
        RECT 118.790 134.485 119.065 134.940 ;
        RECT 119.235 134.655 119.480 135.135 ;
        RECT 119.650 134.485 119.910 134.940 ;
        RECT 120.080 134.655 120.340 135.135 ;
        RECT 120.510 134.485 120.770 134.940 ;
        RECT 120.940 134.655 121.200 135.135 ;
        RECT 121.370 134.485 121.630 134.940 ;
        RECT 121.800 134.575 122.060 135.135 ;
        RECT 114.885 134.315 121.630 134.485 ;
        RECT 113.345 133.975 113.705 134.145 ;
        RECT 113.375 133.895 113.705 133.975 ;
        RECT 114.885 133.725 116.050 134.315 ;
        RECT 122.230 134.145 122.480 134.955 ;
        RECT 122.660 134.610 122.920 135.135 ;
        RECT 123.090 134.145 123.340 134.955 ;
        RECT 123.520 134.625 123.825 135.135 ;
        RECT 116.220 133.895 123.340 134.145 ;
        RECT 123.510 133.895 123.825 134.455 ;
        RECT 123.995 134.385 125.205 135.135 ;
        RECT 110.665 133.265 113.175 133.435 ;
        RECT 110.665 132.585 111.175 133.095 ;
        RECT 112.345 132.755 112.675 133.265 ;
        RECT 113.345 132.585 113.705 133.725 ;
        RECT 114.885 133.500 121.630 133.725 ;
        RECT 114.885 132.585 115.155 133.330 ;
        RECT 115.325 132.760 115.615 133.500 ;
        RECT 116.225 133.485 121.630 133.500 ;
        RECT 115.785 132.590 116.040 133.315 ;
        RECT 116.225 132.760 116.485 133.485 ;
        RECT 116.655 132.590 116.900 133.315 ;
        RECT 117.085 132.760 117.345 133.485 ;
        RECT 117.515 132.590 117.760 133.315 ;
        RECT 117.945 132.760 118.205 133.485 ;
        RECT 118.375 132.590 118.620 133.315 ;
        RECT 118.790 132.760 119.050 133.485 ;
        RECT 119.220 132.590 119.480 133.315 ;
        RECT 119.650 132.760 119.910 133.485 ;
        RECT 120.080 132.590 120.340 133.315 ;
        RECT 120.510 132.760 120.770 133.485 ;
        RECT 120.940 132.590 121.200 133.315 ;
        RECT 121.370 132.760 121.630 133.485 ;
        RECT 121.800 132.590 122.060 133.385 ;
        RECT 122.230 132.760 122.480 133.895 ;
        RECT 115.785 132.585 122.060 132.590 ;
        RECT 122.660 132.585 122.920 133.395 ;
        RECT 123.095 132.755 123.340 133.895 ;
        RECT 123.995 133.675 124.515 134.215 ;
        RECT 124.685 133.845 125.205 134.385 ;
        RECT 123.520 132.585 123.815 133.395 ;
        RECT 123.995 132.585 125.205 133.675 ;
        RECT 53.990 132.415 125.290 132.585 ;
        RECT 54.075 131.325 55.285 132.415 ;
        RECT 54.075 130.615 54.595 131.155 ;
        RECT 54.765 130.785 55.285 131.325 ;
        RECT 56.375 131.340 56.645 132.245 ;
        RECT 56.815 131.655 57.145 132.415 ;
        RECT 57.325 131.485 57.495 132.245 ;
        RECT 54.075 129.865 55.285 130.615 ;
        RECT 56.375 130.540 56.545 131.340 ;
        RECT 56.830 131.315 57.495 131.485 ;
        RECT 57.755 131.340 58.025 132.245 ;
        RECT 58.195 131.655 58.525 132.415 ;
        RECT 58.705 131.485 58.875 132.245 ;
        RECT 56.830 131.170 57.000 131.315 ;
        RECT 56.715 130.840 57.000 131.170 ;
        RECT 56.830 130.585 57.000 130.840 ;
        RECT 57.235 130.765 57.565 131.135 ;
        RECT 56.375 130.035 56.635 130.540 ;
        RECT 56.830 130.415 57.495 130.585 ;
        RECT 56.815 129.865 57.145 130.245 ;
        RECT 57.325 130.035 57.495 130.415 ;
        RECT 57.755 130.540 57.925 131.340 ;
        RECT 58.210 131.315 58.875 131.485 ;
        RECT 59.135 131.340 59.405 132.245 ;
        RECT 59.575 131.655 59.905 132.415 ;
        RECT 60.085 131.485 60.255 132.245 ;
        RECT 60.705 131.690 61.035 132.415 ;
        RECT 58.210 131.170 58.380 131.315 ;
        RECT 58.095 130.840 58.380 131.170 ;
        RECT 58.210 130.585 58.380 130.840 ;
        RECT 58.615 130.765 58.945 131.135 ;
        RECT 57.755 130.035 58.015 130.540 ;
        RECT 58.210 130.415 58.875 130.585 ;
        RECT 58.195 129.865 58.525 130.245 ;
        RECT 58.705 130.035 58.875 130.415 ;
        RECT 59.135 130.540 59.305 131.340 ;
        RECT 59.590 131.315 60.255 131.485 ;
        RECT 59.590 131.170 59.760 131.315 ;
        RECT 59.475 130.840 59.760 131.170 ;
        RECT 59.590 130.585 59.760 130.840 ;
        RECT 59.995 130.765 60.325 131.135 ;
        RECT 59.135 130.035 59.395 130.540 ;
        RECT 59.590 130.415 60.255 130.585 ;
        RECT 59.575 129.865 59.905 130.245 ;
        RECT 60.085 130.035 60.255 130.415 ;
        RECT 60.515 130.035 61.035 131.520 ;
        RECT 61.205 130.695 61.725 132.245 ;
        RECT 62.080 131.445 62.470 131.620 ;
        RECT 62.955 131.615 63.285 132.415 ;
        RECT 63.455 131.625 63.990 132.245 ;
        RECT 62.080 131.275 63.505 131.445 ;
        RECT 61.955 130.545 62.310 131.105 ;
        RECT 61.205 129.865 61.545 130.525 ;
        RECT 62.480 130.375 62.650 131.275 ;
        RECT 62.820 130.545 63.085 131.105 ;
        RECT 63.335 130.775 63.505 131.275 ;
        RECT 63.675 130.605 63.990 131.625 ;
        RECT 64.200 131.265 64.460 132.415 ;
        RECT 64.635 131.340 64.890 132.245 ;
        RECT 65.060 131.655 65.390 132.415 ;
        RECT 65.605 131.485 65.775 132.245 ;
        RECT 62.060 129.865 62.300 130.375 ;
        RECT 62.480 130.045 62.760 130.375 ;
        RECT 62.990 129.865 63.205 130.375 ;
        RECT 63.375 130.035 63.990 130.605 ;
        RECT 64.200 129.865 64.460 130.705 ;
        RECT 64.635 130.610 64.805 131.340 ;
        RECT 65.060 131.315 65.775 131.485 ;
        RECT 65.060 131.105 65.230 131.315 ;
        RECT 66.955 131.250 67.245 132.415 ;
        RECT 68.340 131.275 68.675 132.245 ;
        RECT 68.845 131.275 69.015 132.415 ;
        RECT 69.185 132.075 71.215 132.245 ;
        RECT 64.975 130.775 65.230 131.105 ;
        RECT 64.635 130.035 64.890 130.610 ;
        RECT 65.060 130.585 65.230 130.775 ;
        RECT 65.510 130.765 65.865 131.135 ;
        RECT 68.340 130.605 68.510 131.275 ;
        RECT 69.185 131.105 69.355 132.075 ;
        RECT 68.680 130.775 68.935 131.105 ;
        RECT 69.160 130.775 69.355 131.105 ;
        RECT 69.525 131.735 70.650 131.905 ;
        RECT 68.765 130.605 68.935 130.775 ;
        RECT 69.525 130.605 69.695 131.735 ;
        RECT 65.060 130.415 65.775 130.585 ;
        RECT 65.060 129.865 65.390 130.245 ;
        RECT 65.605 130.035 65.775 130.415 ;
        RECT 66.955 129.865 67.245 130.590 ;
        RECT 68.340 130.035 68.595 130.605 ;
        RECT 68.765 130.435 69.695 130.605 ;
        RECT 69.865 131.395 70.875 131.565 ;
        RECT 69.865 130.595 70.035 131.395 ;
        RECT 69.520 130.400 69.695 130.435 ;
        RECT 68.765 129.865 69.095 130.265 ;
        RECT 69.520 130.035 70.050 130.400 ;
        RECT 70.240 130.375 70.515 131.195 ;
        RECT 70.235 130.205 70.515 130.375 ;
        RECT 70.240 130.035 70.515 130.205 ;
        RECT 70.685 130.035 70.875 131.395 ;
        RECT 71.045 131.410 71.215 132.075 ;
        RECT 71.385 131.655 71.555 132.415 ;
        RECT 71.790 131.655 72.305 132.065 ;
        RECT 71.045 131.220 71.795 131.410 ;
        RECT 71.965 130.845 72.305 131.655 ;
        RECT 73.025 131.485 73.195 132.245 ;
        RECT 73.375 131.655 73.705 132.415 ;
        RECT 73.025 131.315 73.690 131.485 ;
        RECT 73.875 131.340 74.145 132.245 ;
        RECT 73.520 131.170 73.690 131.315 ;
        RECT 71.075 130.675 72.305 130.845 ;
        RECT 72.955 130.765 73.285 131.135 ;
        RECT 73.520 130.840 73.805 131.170 ;
        RECT 71.055 129.865 71.565 130.400 ;
        RECT 71.785 130.070 72.030 130.675 ;
        RECT 73.520 130.585 73.690 130.840 ;
        RECT 73.025 130.415 73.690 130.585 ;
        RECT 73.975 130.540 74.145 131.340 ;
        RECT 74.325 131.805 74.655 132.235 ;
        RECT 74.835 131.975 75.030 132.415 ;
        RECT 75.200 131.805 75.530 132.235 ;
        RECT 74.325 131.635 75.530 131.805 ;
        RECT 74.325 131.305 75.220 131.635 ;
        RECT 75.700 131.465 75.975 132.235 ;
        RECT 76.245 131.670 76.515 132.415 ;
        RECT 77.145 132.410 83.420 132.415 ;
        RECT 76.685 131.500 76.975 132.240 ;
        RECT 77.145 131.685 77.400 132.410 ;
        RECT 77.585 131.515 77.845 132.240 ;
        RECT 78.015 131.685 78.260 132.410 ;
        RECT 78.445 131.515 78.705 132.240 ;
        RECT 78.875 131.685 79.120 132.410 ;
        RECT 79.305 131.515 79.565 132.240 ;
        RECT 79.735 131.685 79.980 132.410 ;
        RECT 80.150 131.515 80.410 132.240 ;
        RECT 80.580 131.685 80.840 132.410 ;
        RECT 81.010 131.515 81.270 132.240 ;
        RECT 81.440 131.685 81.700 132.410 ;
        RECT 81.870 131.515 82.130 132.240 ;
        RECT 82.300 131.685 82.560 132.410 ;
        RECT 82.730 131.515 82.990 132.240 ;
        RECT 83.160 131.615 83.420 132.410 ;
        RECT 77.585 131.500 82.990 131.515 ;
        RECT 75.390 131.275 75.975 131.465 ;
        RECT 76.245 131.275 82.990 131.500 ;
        RECT 74.330 130.775 74.625 131.105 ;
        RECT 74.805 130.775 75.220 131.105 ;
        RECT 73.025 130.035 73.195 130.415 ;
        RECT 73.375 129.865 73.705 130.245 ;
        RECT 73.885 130.035 74.145 130.540 ;
        RECT 74.325 129.865 74.625 130.595 ;
        RECT 74.805 130.155 75.035 130.775 ;
        RECT 75.390 130.605 75.565 131.275 ;
        RECT 75.235 130.425 75.565 130.605 ;
        RECT 75.735 130.455 75.975 131.105 ;
        RECT 76.245 130.685 77.410 131.275 ;
        RECT 83.590 131.105 83.840 132.240 ;
        RECT 84.020 131.605 84.280 132.415 ;
        RECT 84.455 131.105 84.700 132.245 ;
        RECT 84.880 131.605 85.175 132.415 ;
        RECT 85.360 131.545 85.625 132.245 ;
        RECT 85.795 131.715 86.125 132.415 ;
        RECT 86.295 131.545 86.965 132.245 ;
        RECT 87.470 131.715 87.900 132.415 ;
        RECT 88.080 131.855 88.270 132.245 ;
        RECT 88.440 132.035 88.770 132.415 ;
        RECT 89.125 132.075 90.285 132.245 ;
        RECT 88.080 131.685 88.810 131.855 ;
        RECT 85.360 131.290 87.935 131.545 ;
        RECT 77.580 130.855 84.700 131.105 ;
        RECT 76.245 130.515 82.990 130.685 ;
        RECT 75.235 130.045 75.460 130.425 ;
        RECT 75.630 129.865 75.960 130.255 ;
        RECT 76.245 129.865 76.545 130.345 ;
        RECT 76.715 130.060 76.975 130.515 ;
        RECT 77.145 129.865 77.405 130.345 ;
        RECT 77.585 130.060 77.845 130.515 ;
        RECT 78.015 129.865 78.265 130.345 ;
        RECT 78.445 130.060 78.705 130.515 ;
        RECT 78.875 129.865 79.125 130.345 ;
        RECT 79.305 130.060 79.565 130.515 ;
        RECT 79.735 129.865 79.980 130.345 ;
        RECT 80.150 130.060 80.425 130.515 ;
        RECT 80.595 129.865 80.840 130.345 ;
        RECT 81.010 130.060 81.270 130.515 ;
        RECT 81.440 129.865 81.700 130.345 ;
        RECT 81.870 130.060 82.130 130.515 ;
        RECT 82.300 129.865 82.560 130.345 ;
        RECT 82.730 130.060 82.990 130.515 ;
        RECT 83.160 129.865 83.420 130.425 ;
        RECT 83.590 130.045 83.840 130.855 ;
        RECT 84.020 129.865 84.280 130.390 ;
        RECT 84.450 130.045 84.700 130.855 ;
        RECT 84.870 130.545 85.185 131.105 ;
        RECT 85.355 130.775 85.630 131.105 ;
        RECT 85.800 130.605 85.980 131.290 ;
        RECT 87.765 131.105 87.935 131.290 ;
        RECT 86.150 130.775 86.510 131.105 ;
        RECT 86.800 131.055 87.090 131.105 ;
        RECT 86.795 130.885 87.090 131.055 ;
        RECT 86.800 130.775 87.090 130.885 ;
        RECT 87.260 130.775 87.595 131.105 ;
        RECT 87.765 130.775 88.445 131.105 ;
        RECT 84.880 129.865 85.185 130.375 ;
        RECT 85.365 130.205 85.980 130.605 ;
        RECT 86.150 130.415 87.420 130.605 ;
        RECT 88.615 130.565 88.810 131.685 ;
        RECT 89.125 131.575 89.295 132.075 ;
        RECT 89.555 131.445 89.725 131.905 ;
        RECT 89.955 131.825 90.285 132.075 ;
        RECT 90.510 131.995 90.840 132.415 ;
        RECT 91.095 131.825 91.380 132.245 ;
        RECT 89.955 131.655 91.380 131.825 ;
        RECT 91.625 131.615 91.955 132.415 ;
        RECT 92.205 131.695 92.540 132.205 ;
        RECT 89.100 131.105 89.305 131.395 ;
        RECT 89.555 131.275 91.925 131.445 ;
        RECT 91.755 131.105 91.925 131.275 ;
        RECT 89.100 131.055 89.450 131.105 ;
        RECT 89.095 130.885 89.450 131.055 ;
        RECT 89.100 130.775 89.450 130.885 ;
        RECT 87.990 130.395 88.810 130.565 ;
        RECT 85.365 130.035 85.700 130.205 ;
        RECT 86.660 129.865 86.995 130.245 ;
        RECT 87.585 129.865 87.820 130.305 ;
        RECT 87.990 130.035 88.320 130.395 ;
        RECT 88.490 129.865 88.820 130.225 ;
        RECT 89.045 129.865 89.375 130.585 ;
        RECT 89.760 130.440 90.180 131.105 ;
        RECT 90.350 130.715 90.640 131.105 ;
        RECT 90.830 131.055 91.100 131.105 ;
        RECT 91.310 131.055 91.560 131.105 ;
        RECT 90.830 130.885 91.105 131.055 ;
        RECT 91.310 130.885 91.565 131.055 ;
        RECT 90.350 130.545 90.645 130.715 ;
        RECT 90.350 130.445 90.640 130.545 ;
        RECT 90.830 130.445 91.100 130.885 ;
        RECT 91.310 130.775 91.560 130.885 ;
        RECT 91.755 130.775 92.060 131.105 ;
        RECT 91.755 130.605 91.925 130.775 ;
        RECT 91.365 130.435 91.925 130.605 ;
        RECT 91.365 130.265 91.535 130.435 ;
        RECT 92.285 130.340 92.540 131.695 ;
        RECT 92.715 131.250 93.005 132.415 ;
        RECT 93.230 131.545 93.515 132.415 ;
        RECT 93.685 131.785 93.945 132.245 ;
        RECT 94.120 131.955 94.375 132.415 ;
        RECT 94.545 131.785 94.805 132.245 ;
        RECT 93.685 131.615 94.805 131.785 ;
        RECT 94.975 131.615 95.285 132.415 ;
        RECT 93.685 131.365 93.945 131.615 ;
        RECT 95.455 131.445 95.765 132.245 ;
        RECT 95.935 131.995 96.275 132.415 ;
        RECT 96.445 131.825 96.695 132.245 ;
        RECT 93.190 131.195 93.945 131.365 ;
        RECT 94.735 131.275 95.765 131.445 ;
        RECT 93.190 130.685 93.595 131.195 ;
        RECT 94.735 131.025 94.905 131.275 ;
        RECT 93.765 130.855 94.905 131.025 ;
        RECT 89.920 130.095 91.535 130.265 ;
        RECT 91.705 129.865 92.035 130.265 ;
        RECT 92.205 130.080 92.540 130.340 ;
        RECT 92.715 129.865 93.005 130.590 ;
        RECT 93.190 130.515 94.840 130.685 ;
        RECT 95.075 130.535 95.425 131.105 ;
        RECT 93.235 129.865 93.515 130.345 ;
        RECT 93.685 130.125 93.945 130.515 ;
        RECT 94.120 129.865 94.375 130.345 ;
        RECT 94.545 130.125 94.840 130.515 ;
        RECT 95.595 130.365 95.765 131.275 ;
        RECT 95.935 131.655 96.695 131.825 ;
        RECT 95.935 130.685 96.245 131.655 ;
        RECT 96.865 131.575 97.195 132.415 ;
        RECT 97.685 131.825 98.440 132.245 ;
        RECT 97.365 131.655 98.830 131.825 ;
        RECT 97.365 131.405 97.535 131.655 ;
        RECT 96.575 131.235 97.535 131.405 ;
        RECT 96.575 131.065 96.745 131.235 ;
        RECT 97.705 131.065 98.010 131.485 ;
        RECT 96.415 130.855 96.745 131.065 ;
        RECT 96.915 130.855 97.355 131.065 ;
        RECT 97.525 130.855 98.010 131.065 ;
        RECT 98.200 131.055 98.490 131.485 ;
        RECT 98.660 131.450 98.830 131.655 ;
        RECT 99.000 131.630 99.240 132.415 ;
        RECT 99.410 131.450 99.740 132.245 ;
        RECT 100.085 131.605 100.380 132.415 ;
        RECT 98.660 131.275 99.740 131.450 ;
        RECT 98.660 131.225 99.445 131.275 ;
        RECT 98.200 130.855 98.590 131.055 ;
        RECT 98.760 130.855 99.105 131.055 ;
        RECT 95.935 130.515 96.695 130.685 ;
        RECT 95.020 129.865 95.295 130.345 ;
        RECT 95.465 130.035 95.765 130.365 ;
        RECT 96.025 129.865 96.195 130.345 ;
        RECT 96.365 130.045 96.695 130.515 ;
        RECT 96.865 129.865 97.035 130.685 ;
        RECT 97.205 130.515 98.905 130.685 ;
        RECT 97.205 130.050 97.535 130.515 ;
        RECT 98.520 130.425 98.905 130.515 ;
        RECT 99.275 130.585 99.445 131.225 ;
        RECT 100.560 131.105 100.805 132.245 ;
        RECT 100.980 131.605 101.240 132.415 ;
        RECT 101.840 132.410 108.115 132.415 ;
        RECT 101.420 131.105 101.670 132.240 ;
        RECT 101.840 131.615 102.100 132.410 ;
        RECT 102.270 131.515 102.530 132.240 ;
        RECT 102.700 131.685 102.960 132.410 ;
        RECT 103.130 131.515 103.390 132.240 ;
        RECT 103.560 131.685 103.820 132.410 ;
        RECT 103.990 131.515 104.250 132.240 ;
        RECT 104.420 131.685 104.680 132.410 ;
        RECT 104.850 131.515 105.110 132.240 ;
        RECT 105.280 131.685 105.525 132.410 ;
        RECT 105.695 131.515 105.955 132.240 ;
        RECT 106.140 131.685 106.385 132.410 ;
        RECT 106.555 131.515 106.815 132.240 ;
        RECT 107.000 131.685 107.245 132.410 ;
        RECT 107.415 131.515 107.675 132.240 ;
        RECT 107.860 131.685 108.115 132.410 ;
        RECT 102.270 131.500 107.675 131.515 ;
        RECT 108.285 131.500 108.575 132.240 ;
        RECT 108.745 131.670 109.015 132.415 ;
        RECT 109.365 131.670 109.635 132.415 ;
        RECT 110.265 132.410 116.540 132.415 ;
        RECT 109.805 131.500 110.095 132.240 ;
        RECT 110.265 131.685 110.520 132.410 ;
        RECT 110.705 131.515 110.965 132.240 ;
        RECT 111.135 131.685 111.380 132.410 ;
        RECT 111.565 131.515 111.825 132.240 ;
        RECT 111.995 131.685 112.240 132.410 ;
        RECT 112.425 131.515 112.685 132.240 ;
        RECT 112.855 131.685 113.100 132.410 ;
        RECT 113.270 131.515 113.530 132.240 ;
        RECT 113.700 131.685 113.960 132.410 ;
        RECT 114.130 131.515 114.390 132.240 ;
        RECT 114.560 131.685 114.820 132.410 ;
        RECT 114.990 131.515 115.250 132.240 ;
        RECT 115.420 131.685 115.680 132.410 ;
        RECT 115.850 131.515 116.110 132.240 ;
        RECT 116.280 131.615 116.540 132.410 ;
        RECT 110.705 131.500 116.110 131.515 ;
        RECT 102.270 131.275 109.015 131.500 ;
        RECT 99.645 130.755 99.905 131.105 ;
        RECT 99.275 130.415 99.820 130.585 ;
        RECT 100.075 130.545 100.390 131.105 ;
        RECT 100.560 130.855 107.680 131.105 ;
        RECT 107.850 131.055 109.015 131.275 ;
        RECT 109.365 131.275 116.110 131.500 ;
        RECT 107.850 130.885 109.045 131.055 ;
        RECT 97.705 129.865 97.875 130.335 ;
        RECT 98.135 130.075 99.320 130.245 ;
        RECT 99.490 130.035 99.820 130.415 ;
        RECT 100.075 129.865 100.380 130.375 ;
        RECT 100.560 130.045 100.810 130.855 ;
        RECT 100.980 129.865 101.240 130.390 ;
        RECT 101.420 130.045 101.670 130.855 ;
        RECT 107.850 130.685 109.015 130.885 ;
        RECT 102.270 130.515 109.015 130.685 ;
        RECT 109.365 130.685 110.530 131.275 ;
        RECT 116.710 131.105 116.960 132.240 ;
        RECT 117.140 131.605 117.400 132.415 ;
        RECT 117.575 131.105 117.820 132.245 ;
        RECT 118.000 131.605 118.295 132.415 ;
        RECT 118.475 131.250 118.765 132.415 ;
        RECT 118.995 131.715 119.215 132.245 ;
        RECT 119.385 131.905 119.715 132.415 ;
        RECT 119.885 131.715 120.110 132.245 ;
        RECT 118.995 131.450 120.110 131.715 ;
        RECT 120.280 131.700 120.595 132.245 ;
        RECT 120.785 132.000 121.115 132.415 ;
        RECT 120.280 131.470 121.115 131.700 ;
        RECT 110.700 130.855 117.820 131.105 ;
        RECT 109.365 130.515 116.110 130.685 ;
        RECT 101.840 129.865 102.100 130.425 ;
        RECT 102.270 130.060 102.530 130.515 ;
        RECT 102.700 129.865 102.960 130.345 ;
        RECT 103.130 130.060 103.390 130.515 ;
        RECT 103.560 129.865 103.820 130.345 ;
        RECT 103.990 130.060 104.250 130.515 ;
        RECT 104.420 129.865 104.665 130.345 ;
        RECT 104.835 130.060 105.110 130.515 ;
        RECT 105.280 129.865 105.525 130.345 ;
        RECT 105.695 130.060 105.955 130.515 ;
        RECT 106.135 129.865 106.385 130.345 ;
        RECT 106.555 130.060 106.815 130.515 ;
        RECT 106.995 129.865 107.245 130.345 ;
        RECT 107.415 130.060 107.675 130.515 ;
        RECT 107.855 129.865 108.115 130.345 ;
        RECT 108.285 130.060 108.545 130.515 ;
        RECT 108.715 129.865 109.015 130.345 ;
        RECT 109.365 129.865 109.665 130.345 ;
        RECT 109.835 130.060 110.095 130.515 ;
        RECT 110.265 129.865 110.525 130.345 ;
        RECT 110.705 130.060 110.965 130.515 ;
        RECT 111.135 129.865 111.385 130.345 ;
        RECT 111.565 130.060 111.825 130.515 ;
        RECT 111.995 129.865 112.245 130.345 ;
        RECT 112.425 130.060 112.685 130.515 ;
        RECT 112.855 129.865 113.100 130.345 ;
        RECT 113.270 130.060 113.545 130.515 ;
        RECT 113.715 129.865 113.960 130.345 ;
        RECT 114.130 130.060 114.390 130.515 ;
        RECT 114.560 129.865 114.820 130.345 ;
        RECT 114.990 130.060 115.250 130.515 ;
        RECT 115.420 129.865 115.680 130.345 ;
        RECT 115.850 130.060 116.110 130.515 ;
        RECT 116.280 129.865 116.540 130.425 ;
        RECT 116.710 130.045 116.960 130.855 ;
        RECT 117.140 129.865 117.400 130.390 ;
        RECT 117.570 130.045 117.820 130.855 ;
        RECT 117.990 130.545 118.305 131.105 ;
        RECT 118.000 129.865 118.305 130.375 ;
        RECT 118.475 129.865 118.765 130.590 ;
        RECT 118.945 130.530 119.260 131.105 ;
        RECT 118.935 129.865 119.265 130.345 ;
        RECT 119.450 130.145 119.830 131.105 ;
        RECT 120.280 130.775 120.605 131.190 ;
        RECT 120.775 130.775 121.115 131.470 ;
        RECT 120.775 130.605 120.945 130.775 ;
        RECT 121.285 130.605 121.515 132.245 ;
        RECT 121.685 131.445 121.975 132.415 ;
        RECT 122.160 131.615 122.415 132.415 ;
        RECT 122.615 131.565 122.945 132.245 ;
        RECT 122.160 131.075 122.405 131.435 ;
        RECT 122.595 131.285 122.945 131.565 ;
        RECT 122.595 130.905 122.765 131.285 ;
        RECT 123.125 131.105 123.320 132.155 ;
        RECT 123.500 131.275 123.820 132.415 ;
        RECT 123.995 131.325 125.205 132.415 ;
        RECT 120.205 130.435 120.945 130.605 ;
        RECT 120.205 130.035 120.395 130.435 ;
        RECT 121.115 130.415 121.515 130.605 ;
        RECT 122.245 130.735 122.765 130.905 ;
        RECT 122.935 130.775 123.320 131.105 ;
        RECT 123.500 131.055 123.760 131.105 ;
        RECT 123.500 130.885 123.765 131.055 ;
        RECT 123.500 130.775 123.760 130.885 ;
        RECT 123.995 130.785 124.515 131.325 ;
        RECT 120.615 129.865 120.945 130.225 ;
        RECT 121.115 130.035 121.305 130.415 ;
        RECT 121.475 129.865 121.805 130.245 ;
        RECT 122.245 130.170 122.415 130.735 ;
        RECT 124.685 130.615 125.205 131.155 ;
        RECT 122.605 130.395 123.820 130.565 ;
        RECT 122.605 130.090 122.835 130.395 ;
        RECT 123.005 129.865 123.335 130.225 ;
        RECT 123.530 130.045 123.820 130.395 ;
        RECT 123.995 129.865 125.205 130.615 ;
        RECT 53.990 129.695 125.290 129.865 ;
        RECT 54.075 128.945 55.285 129.695 ;
        RECT 54.075 128.405 54.595 128.945 ;
        RECT 55.460 128.855 55.720 129.695 ;
        RECT 55.895 128.950 56.150 129.525 ;
        RECT 56.320 129.315 56.650 129.695 ;
        RECT 56.865 129.145 57.035 129.525 ;
        RECT 56.320 128.975 57.035 129.145 ;
        RECT 54.765 128.235 55.285 128.775 ;
        RECT 54.075 127.145 55.285 128.235 ;
        RECT 55.460 127.145 55.720 128.295 ;
        RECT 55.895 128.220 56.065 128.950 ;
        RECT 56.320 128.785 56.490 128.975 ;
        RECT 57.295 128.895 57.605 129.695 ;
        RECT 57.810 128.895 58.505 129.525 ;
        RECT 58.675 128.955 59.165 129.525 ;
        RECT 59.335 129.125 59.565 129.525 ;
        RECT 59.735 129.295 60.155 129.695 ;
        RECT 60.325 129.125 60.495 129.525 ;
        RECT 59.335 128.955 60.495 129.125 ;
        RECT 60.665 128.955 61.115 129.695 ;
        RECT 61.285 128.955 61.725 129.515 ;
        RECT 57.810 128.845 57.985 128.895 ;
        RECT 56.235 128.455 56.490 128.785 ;
        RECT 56.320 128.245 56.490 128.455 ;
        RECT 56.770 128.425 57.125 128.795 ;
        RECT 57.305 128.455 57.640 128.725 ;
        RECT 57.810 128.295 57.980 128.845 ;
        RECT 58.150 128.455 58.485 128.705 ;
        RECT 55.895 127.315 56.150 128.220 ;
        RECT 56.320 128.075 57.035 128.245 ;
        RECT 56.320 127.145 56.650 127.905 ;
        RECT 56.865 127.315 57.035 128.075 ;
        RECT 57.295 127.145 57.575 128.285 ;
        RECT 57.745 127.315 58.075 128.295 ;
        RECT 58.675 128.285 58.845 128.955 ;
        RECT 59.015 128.455 59.420 128.785 ;
        RECT 58.245 127.145 58.505 128.285 ;
        RECT 58.675 128.115 59.445 128.285 ;
        RECT 58.685 127.145 59.015 127.945 ;
        RECT 59.195 127.485 59.445 128.115 ;
        RECT 59.635 127.655 59.885 128.785 ;
        RECT 60.085 128.455 60.330 128.785 ;
        RECT 60.515 128.505 60.905 128.785 ;
        RECT 60.085 127.655 60.285 128.455 ;
        RECT 61.075 128.335 61.245 128.785 ;
        RECT 60.455 128.165 61.245 128.335 ;
        RECT 60.455 127.485 60.625 128.165 ;
        RECT 59.195 127.315 60.625 127.485 ;
        RECT 60.795 127.145 61.110 127.995 ;
        RECT 61.415 127.945 61.725 128.955 ;
        RECT 61.285 127.315 61.725 127.945 ;
        RECT 62.815 128.955 63.155 129.525 ;
        RECT 63.350 129.030 63.520 129.695 ;
        RECT 63.800 129.355 64.020 129.400 ;
        RECT 63.795 129.185 64.020 129.355 ;
        RECT 64.190 129.215 64.635 129.385 ;
        RECT 63.800 129.045 64.020 129.185 ;
        RECT 62.815 127.985 62.990 128.955 ;
        RECT 63.800 128.875 64.295 129.045 ;
        RECT 63.160 128.335 63.330 128.785 ;
        RECT 63.500 128.505 63.950 128.705 ;
        RECT 64.120 128.680 64.295 128.875 ;
        RECT 64.465 128.425 64.635 129.215 ;
        RECT 64.805 129.090 65.055 129.460 ;
        RECT 64.885 128.705 65.055 129.090 ;
        RECT 65.225 129.055 65.475 129.460 ;
        RECT 65.645 129.225 65.815 129.695 ;
        RECT 65.985 129.055 66.325 129.460 ;
        RECT 65.225 128.875 66.325 129.055 ;
        RECT 66.515 128.885 66.755 129.695 ;
        RECT 66.925 128.885 67.255 129.525 ;
        RECT 67.425 128.885 67.695 129.695 ;
        RECT 64.885 128.535 65.080 128.705 ;
        RECT 63.160 128.165 63.555 128.335 ;
        RECT 64.465 128.285 64.740 128.425 ;
        RECT 62.815 127.315 63.075 127.985 ;
        RECT 63.385 127.895 63.555 128.165 ;
        RECT 63.725 128.065 64.740 128.285 ;
        RECT 64.910 128.285 65.080 128.535 ;
        RECT 65.250 128.455 65.810 128.705 ;
        RECT 64.910 127.895 65.465 128.285 ;
        RECT 63.385 127.725 65.465 127.895 ;
        RECT 63.245 127.145 63.575 127.545 ;
        RECT 64.445 127.145 64.845 127.545 ;
        RECT 65.135 127.490 65.465 127.725 ;
        RECT 65.635 127.355 65.810 128.455 ;
        RECT 65.980 128.135 66.325 128.705 ;
        RECT 66.495 128.455 66.845 128.705 ;
        RECT 67.015 128.285 67.185 128.885 ;
        RECT 67.915 128.875 68.145 129.695 ;
        RECT 68.315 128.895 68.645 129.525 ;
        RECT 67.355 128.455 67.705 128.705 ;
        RECT 67.895 128.455 68.225 128.705 ;
        RECT 68.395 128.295 68.645 128.895 ;
        RECT 68.815 128.875 69.025 129.695 ;
        RECT 69.260 128.955 69.515 129.525 ;
        RECT 69.685 129.295 70.015 129.695 ;
        RECT 70.440 129.160 70.970 129.525 ;
        RECT 70.440 129.125 70.615 129.160 ;
        RECT 69.685 128.955 70.615 129.125 ;
        RECT 71.160 129.015 71.435 129.525 ;
        RECT 66.505 128.115 67.185 128.285 ;
        RECT 65.980 127.145 66.325 127.965 ;
        RECT 66.505 127.330 66.835 128.115 ;
        RECT 67.365 127.145 67.695 128.285 ;
        RECT 67.915 127.145 68.145 128.285 ;
        RECT 68.315 127.315 68.645 128.295 ;
        RECT 69.260 128.285 69.430 128.955 ;
        RECT 69.685 128.785 69.855 128.955 ;
        RECT 69.600 128.455 69.855 128.785 ;
        RECT 70.080 128.455 70.275 128.785 ;
        RECT 68.815 127.145 69.025 128.285 ;
        RECT 69.260 127.315 69.595 128.285 ;
        RECT 69.765 127.145 69.935 128.285 ;
        RECT 70.105 127.485 70.275 128.455 ;
        RECT 70.445 127.825 70.615 128.955 ;
        RECT 70.785 128.165 70.955 128.965 ;
        RECT 71.155 128.845 71.435 129.015 ;
        RECT 71.160 128.365 71.435 128.845 ;
        RECT 71.605 128.165 71.795 129.525 ;
        RECT 71.975 129.160 72.485 129.695 ;
        RECT 72.705 128.885 72.950 129.490 ;
        RECT 73.400 128.955 73.655 129.525 ;
        RECT 73.825 129.295 74.155 129.695 ;
        RECT 74.580 129.160 75.110 129.525 ;
        RECT 74.580 129.125 74.755 129.160 ;
        RECT 73.825 128.955 74.755 129.125 ;
        RECT 71.995 128.715 73.225 128.885 ;
        RECT 70.785 127.995 71.795 128.165 ;
        RECT 71.965 128.150 72.715 128.340 ;
        RECT 70.445 127.655 71.570 127.825 ;
        RECT 71.965 127.485 72.135 128.150 ;
        RECT 72.885 127.905 73.225 128.715 ;
        RECT 70.105 127.315 72.135 127.485 ;
        RECT 72.305 127.145 72.475 127.905 ;
        RECT 72.710 127.495 73.225 127.905 ;
        RECT 73.400 128.285 73.570 128.955 ;
        RECT 73.825 128.785 73.995 128.955 ;
        RECT 73.740 128.455 73.995 128.785 ;
        RECT 74.220 128.455 74.415 128.785 ;
        RECT 73.400 127.315 73.735 128.285 ;
        RECT 73.905 127.145 74.075 128.285 ;
        RECT 74.245 127.485 74.415 128.455 ;
        RECT 74.585 127.825 74.755 128.955 ;
        RECT 74.925 128.165 75.095 128.965 ;
        RECT 75.300 128.675 75.575 129.525 ;
        RECT 75.295 128.505 75.575 128.675 ;
        RECT 75.300 128.365 75.575 128.505 ;
        RECT 75.745 128.165 75.935 129.525 ;
        RECT 76.115 129.160 76.625 129.695 ;
        RECT 76.845 128.885 77.090 129.490 ;
        RECT 78.085 129.145 78.255 129.525 ;
        RECT 78.470 129.315 78.800 129.695 ;
        RECT 78.085 128.975 78.800 129.145 ;
        RECT 76.135 128.715 77.365 128.885 ;
        RECT 74.925 127.995 75.935 128.165 ;
        RECT 76.105 128.150 76.855 128.340 ;
        RECT 74.585 127.655 75.710 127.825 ;
        RECT 76.105 127.485 76.275 128.150 ;
        RECT 77.025 127.905 77.365 128.715 ;
        RECT 77.995 128.425 78.350 128.795 ;
        RECT 78.630 128.785 78.800 128.975 ;
        RECT 78.970 128.950 79.225 129.525 ;
        RECT 78.630 128.455 78.885 128.785 ;
        RECT 78.630 128.245 78.800 128.455 ;
        RECT 74.245 127.315 76.275 127.485 ;
        RECT 76.445 127.145 76.615 127.905 ;
        RECT 76.850 127.495 77.365 127.905 ;
        RECT 78.085 128.075 78.800 128.245 ;
        RECT 79.055 128.220 79.225 128.950 ;
        RECT 79.400 128.855 79.660 129.695 ;
        RECT 79.835 128.970 80.125 129.695 ;
        RECT 80.345 128.895 80.555 129.695 ;
        RECT 78.085 127.315 78.255 128.075 ;
        RECT 78.470 127.145 78.800 127.905 ;
        RECT 78.970 127.315 79.225 128.220 ;
        RECT 79.400 127.145 79.660 128.295 ;
        RECT 79.835 127.145 80.125 128.310 ;
        RECT 80.345 127.145 80.555 128.285 ;
        RECT 80.725 127.315 81.065 129.525 ;
        RECT 81.245 129.235 81.495 129.695 ;
        RECT 81.685 129.065 82.015 129.525 ;
        RECT 82.215 129.355 82.600 129.525 ;
        RECT 82.195 129.185 82.600 129.355 ;
        RECT 81.240 128.895 82.015 129.065 ;
        RECT 81.240 127.995 81.515 128.895 ;
        RECT 81.715 128.165 82.045 128.705 ;
        RECT 82.215 128.165 82.600 129.185 ;
        RECT 83.075 129.155 83.405 129.525 ;
        RECT 83.595 129.325 83.925 129.695 ;
        RECT 84.095 129.155 84.425 129.525 ;
        RECT 83.075 128.955 84.425 129.155 ;
        RECT 84.895 128.895 85.590 129.525 ;
        RECT 85.795 128.895 86.105 129.695 ;
        RECT 86.360 129.145 86.690 129.525 ;
        RECT 86.860 129.315 88.045 129.485 ;
        RECT 88.305 129.225 88.475 129.695 ;
        RECT 86.360 128.975 86.905 129.145 ;
        RECT 82.890 128.165 83.310 128.705 ;
        RECT 83.510 128.455 83.870 128.785 ;
        RECT 84.040 128.465 84.725 128.775 ;
        RECT 81.240 127.755 83.405 127.995 ;
        RECT 81.245 127.145 81.865 127.585 ;
        RECT 82.070 127.315 82.350 127.755 ;
        RECT 82.535 127.145 82.865 127.525 ;
        RECT 83.075 127.315 83.405 127.755 ;
        RECT 83.580 127.655 83.870 128.455 ;
        RECT 83.575 127.485 83.870 127.655 ;
        RECT 83.580 127.410 83.870 127.485 ;
        RECT 84.095 127.145 84.350 128.285 ;
        RECT 84.520 127.425 84.725 128.465 ;
        RECT 84.915 128.455 85.250 128.705 ;
        RECT 85.420 128.295 85.590 128.895 ;
        RECT 85.760 128.455 86.095 128.725 ;
        RECT 86.275 128.455 86.535 128.805 ;
        RECT 86.735 128.335 86.905 128.975 ;
        RECT 87.275 129.045 87.660 129.135 ;
        RECT 88.645 129.045 88.975 129.510 ;
        RECT 87.275 128.875 88.975 129.045 ;
        RECT 89.145 128.875 89.315 129.695 ;
        RECT 89.485 129.045 89.815 129.515 ;
        RECT 89.985 129.215 90.155 129.695 ;
        RECT 90.425 129.355 91.615 129.525 ;
        RECT 90.425 129.185 90.735 129.355 ;
        RECT 89.485 128.875 90.245 129.045 ;
        RECT 87.075 128.505 87.420 128.705 ;
        RECT 87.590 128.505 87.980 128.705 ;
        RECT 84.895 127.145 85.155 128.285 ;
        RECT 85.325 127.315 85.655 128.295 ;
        RECT 86.735 128.285 87.520 128.335 ;
        RECT 85.825 127.145 86.105 128.285 ;
        RECT 86.440 128.110 87.520 128.285 ;
        RECT 86.440 127.315 86.770 128.110 ;
        RECT 86.940 127.145 87.180 127.930 ;
        RECT 87.350 127.905 87.520 128.110 ;
        RECT 87.690 128.075 87.980 128.505 ;
        RECT 88.170 128.495 88.655 128.705 ;
        RECT 88.825 128.495 89.265 128.705 ;
        RECT 89.435 128.495 89.765 128.705 ;
        RECT 88.170 128.075 88.475 128.495 ;
        RECT 89.435 128.325 89.605 128.495 ;
        RECT 88.645 128.155 89.605 128.325 ;
        RECT 88.645 127.905 88.815 128.155 ;
        RECT 87.350 127.735 88.815 127.905 ;
        RECT 87.740 127.315 88.495 127.735 ;
        RECT 88.985 127.145 89.315 127.985 ;
        RECT 89.935 127.905 90.245 128.875 ;
        RECT 90.420 128.380 90.735 129.015 ;
        RECT 89.485 127.735 90.245 127.905 ;
        RECT 89.485 127.315 89.735 127.735 ;
        RECT 89.905 127.145 90.245 127.565 ;
        RECT 90.425 127.145 90.735 128.210 ;
        RECT 90.905 127.995 91.115 129.185 ;
        RECT 91.285 129.065 91.615 129.355 ;
        RECT 91.855 129.235 92.025 129.695 ;
        RECT 92.255 129.065 92.585 129.525 ;
        RECT 92.765 129.235 92.935 129.695 ;
        RECT 93.115 129.065 93.445 129.525 ;
        RECT 93.695 129.215 93.975 129.695 ;
        RECT 91.285 128.895 93.445 129.065 ;
        RECT 94.145 129.045 94.405 129.435 ;
        RECT 94.580 129.215 94.835 129.695 ;
        RECT 95.005 129.045 95.300 129.435 ;
        RECT 95.480 129.215 95.755 129.695 ;
        RECT 95.925 129.195 96.225 129.525 ;
        RECT 96.485 129.215 96.785 129.695 ;
        RECT 93.650 128.875 95.300 129.045 ;
        RECT 91.455 128.335 91.950 128.705 ;
        RECT 92.130 128.505 92.930 128.705 ;
        RECT 93.100 128.335 93.430 128.725 ;
        RECT 91.395 128.165 93.430 128.335 ;
        RECT 93.650 128.365 94.055 128.875 ;
        RECT 94.225 128.535 95.365 128.705 ;
        RECT 93.650 128.195 94.405 128.365 ;
        RECT 90.905 127.815 92.555 127.995 ;
        RECT 90.905 127.315 91.140 127.815 ;
        RECT 92.255 127.655 92.555 127.815 ;
        RECT 91.310 127.145 91.640 127.605 ;
        RECT 91.835 127.485 92.025 127.645 ;
        RECT 92.725 127.485 92.945 127.995 ;
        RECT 91.835 127.315 92.945 127.485 ;
        RECT 93.115 127.145 93.445 127.995 ;
        RECT 93.690 127.145 93.975 128.015 ;
        RECT 94.145 127.945 94.405 128.195 ;
        RECT 95.195 128.285 95.365 128.535 ;
        RECT 95.535 128.455 95.885 129.025 ;
        RECT 96.055 128.285 96.225 129.195 ;
        RECT 96.955 129.045 97.215 129.500 ;
        RECT 97.385 129.215 97.645 129.695 ;
        RECT 97.825 129.045 98.085 129.500 ;
        RECT 98.255 129.215 98.505 129.695 ;
        RECT 98.685 129.045 98.945 129.500 ;
        RECT 99.115 129.215 99.365 129.695 ;
        RECT 99.545 129.045 99.805 129.500 ;
        RECT 99.975 129.215 100.220 129.695 ;
        RECT 100.390 129.045 100.665 129.500 ;
        RECT 100.835 129.215 101.080 129.695 ;
        RECT 101.250 129.045 101.510 129.500 ;
        RECT 101.680 129.215 101.940 129.695 ;
        RECT 102.110 129.045 102.370 129.500 ;
        RECT 102.540 129.215 102.800 129.695 ;
        RECT 102.970 129.045 103.230 129.500 ;
        RECT 103.400 129.135 103.660 129.695 ;
        RECT 95.195 128.115 96.225 128.285 ;
        RECT 94.145 127.775 95.265 127.945 ;
        RECT 94.145 127.315 94.405 127.775 ;
        RECT 94.580 127.145 94.835 127.605 ;
        RECT 95.005 127.315 95.265 127.775 ;
        RECT 95.435 127.145 95.745 127.945 ;
        RECT 95.915 127.315 96.225 128.115 ;
        RECT 96.485 128.875 103.230 129.045 ;
        RECT 96.485 128.285 97.650 128.875 ;
        RECT 103.830 128.705 104.080 129.515 ;
        RECT 104.260 129.170 104.520 129.695 ;
        RECT 104.690 128.705 104.940 129.515 ;
        RECT 105.120 129.185 105.425 129.695 ;
        RECT 97.820 128.455 104.940 128.705 ;
        RECT 105.110 128.455 105.425 129.015 ;
        RECT 105.595 128.970 105.885 129.695 ;
        RECT 106.080 128.870 106.335 129.695 ;
        RECT 106.505 128.955 106.840 129.525 ;
        RECT 107.035 129.030 107.205 129.695 ;
        RECT 107.485 129.045 107.705 129.400 ;
        RECT 107.875 129.215 108.335 129.385 ;
        RECT 107.485 129.010 107.990 129.045 ;
        RECT 96.485 128.060 103.230 128.285 ;
        RECT 96.485 127.145 96.755 127.890 ;
        RECT 96.925 127.320 97.215 128.060 ;
        RECT 97.825 128.045 103.230 128.060 ;
        RECT 97.385 127.150 97.640 127.875 ;
        RECT 97.825 127.320 98.085 128.045 ;
        RECT 98.255 127.150 98.500 127.875 ;
        RECT 98.685 127.320 98.945 128.045 ;
        RECT 99.115 127.150 99.360 127.875 ;
        RECT 99.545 127.320 99.805 128.045 ;
        RECT 99.975 127.150 100.220 127.875 ;
        RECT 100.390 127.320 100.650 128.045 ;
        RECT 100.820 127.150 101.080 127.875 ;
        RECT 101.250 127.320 101.510 128.045 ;
        RECT 101.680 127.150 101.940 127.875 ;
        RECT 102.110 127.320 102.370 128.045 ;
        RECT 102.540 127.150 102.800 127.875 ;
        RECT 102.970 127.320 103.230 128.045 ;
        RECT 103.400 127.150 103.660 127.945 ;
        RECT 103.830 127.320 104.080 128.455 ;
        RECT 97.385 127.145 103.660 127.150 ;
        RECT 104.260 127.145 104.520 127.955 ;
        RECT 104.695 127.315 104.940 128.455 ;
        RECT 105.120 127.145 105.415 127.955 ;
        RECT 105.595 127.145 105.885 128.310 ;
        RECT 106.080 127.145 106.335 128.370 ;
        RECT 106.505 127.995 106.675 128.955 ;
        RECT 107.485 128.875 107.995 129.010 ;
        RECT 106.845 128.335 107.015 128.785 ;
        RECT 107.185 128.505 107.655 128.705 ;
        RECT 107.825 128.680 107.995 128.875 ;
        RECT 108.165 128.425 108.335 129.215 ;
        RECT 108.505 129.090 108.750 129.460 ;
        RECT 108.580 128.705 108.750 129.090 ;
        RECT 108.925 129.055 109.155 129.460 ;
        RECT 109.345 129.225 109.515 129.695 ;
        RECT 109.685 129.055 110.015 129.460 ;
        RECT 108.925 128.875 110.015 129.055 ;
        RECT 110.195 128.895 110.485 129.695 ;
        RECT 110.655 129.235 111.205 129.525 ;
        RECT 111.375 129.235 111.625 129.695 ;
        RECT 108.580 128.535 108.770 128.705 ;
        RECT 106.845 128.165 107.240 128.335 ;
        RECT 108.165 128.285 108.430 128.425 ;
        RECT 106.505 127.985 106.745 127.995 ;
        RECT 106.505 127.315 106.760 127.985 ;
        RECT 107.070 127.895 107.240 128.165 ;
        RECT 107.410 128.065 108.430 128.285 ;
        RECT 108.600 128.285 108.770 128.535 ;
        RECT 108.940 128.455 109.495 128.705 ;
        RECT 108.600 127.895 109.155 128.285 ;
        RECT 107.070 127.725 109.155 127.895 ;
        RECT 106.930 127.145 107.260 127.545 ;
        RECT 108.130 127.145 108.535 127.545 ;
        RECT 108.805 127.355 109.155 127.725 ;
        RECT 109.325 127.655 109.495 128.455 ;
        RECT 109.670 128.135 110.015 128.705 ;
        RECT 109.325 127.485 109.505 127.655 ;
        RECT 109.325 127.355 109.495 127.485 ;
        RECT 109.700 127.145 110.015 127.965 ;
        RECT 110.195 127.145 110.485 128.285 ;
        RECT 110.655 127.865 110.905 129.235 ;
        RECT 112.255 129.065 112.585 129.425 ;
        RECT 113.045 129.215 113.345 129.695 ;
        RECT 111.195 128.875 112.585 129.065 ;
        RECT 113.515 129.045 113.775 129.500 ;
        RECT 113.945 129.215 114.205 129.695 ;
        RECT 114.385 129.045 114.645 129.500 ;
        RECT 114.815 129.215 115.065 129.695 ;
        RECT 115.245 129.045 115.505 129.500 ;
        RECT 115.675 129.215 115.925 129.695 ;
        RECT 116.105 129.045 116.365 129.500 ;
        RECT 116.535 129.215 116.780 129.695 ;
        RECT 116.950 129.045 117.225 129.500 ;
        RECT 117.395 129.215 117.640 129.695 ;
        RECT 117.810 129.045 118.070 129.500 ;
        RECT 118.240 129.215 118.500 129.695 ;
        RECT 118.670 129.045 118.930 129.500 ;
        RECT 119.100 129.215 119.360 129.695 ;
        RECT 119.530 129.045 119.790 129.500 ;
        RECT 119.960 129.135 120.220 129.695 ;
        RECT 113.045 128.875 119.790 129.045 ;
        RECT 111.195 128.785 111.365 128.875 ;
        RECT 111.075 128.455 111.365 128.785 ;
        RECT 111.535 128.455 111.865 128.705 ;
        RECT 112.095 128.455 112.785 128.705 ;
        RECT 111.195 128.205 111.365 128.455 ;
        RECT 111.195 128.035 112.135 128.205 ;
        RECT 110.655 127.315 111.105 127.865 ;
        RECT 111.295 127.145 111.625 127.865 ;
        RECT 111.835 127.485 112.135 128.035 ;
        RECT 112.470 128.015 112.785 128.455 ;
        RECT 113.045 128.285 114.210 128.875 ;
        RECT 120.390 128.705 120.640 129.515 ;
        RECT 120.820 129.170 121.080 129.695 ;
        RECT 121.250 128.705 121.500 129.515 ;
        RECT 121.680 129.185 121.985 129.695 ;
        RECT 122.160 129.295 122.495 129.695 ;
        RECT 122.665 129.125 122.870 129.525 ;
        RECT 123.080 129.215 123.355 129.695 ;
        RECT 123.565 129.195 123.825 129.525 ;
        RECT 114.380 128.455 121.500 128.705 ;
        RECT 121.670 128.455 121.985 129.015 ;
        RECT 122.185 128.955 122.870 129.125 ;
        RECT 113.045 128.060 119.790 128.285 ;
        RECT 112.305 127.145 112.585 127.815 ;
        RECT 113.045 127.145 113.315 127.890 ;
        RECT 113.485 127.320 113.775 128.060 ;
        RECT 114.385 128.045 119.790 128.060 ;
        RECT 113.945 127.150 114.200 127.875 ;
        RECT 114.385 127.320 114.645 128.045 ;
        RECT 114.815 127.150 115.060 127.875 ;
        RECT 115.245 127.320 115.505 128.045 ;
        RECT 115.675 127.150 115.920 127.875 ;
        RECT 116.105 127.320 116.365 128.045 ;
        RECT 116.535 127.150 116.780 127.875 ;
        RECT 116.950 127.320 117.210 128.045 ;
        RECT 117.380 127.150 117.640 127.875 ;
        RECT 117.810 127.320 118.070 128.045 ;
        RECT 118.240 127.150 118.500 127.875 ;
        RECT 118.670 127.320 118.930 128.045 ;
        RECT 119.100 127.150 119.360 127.875 ;
        RECT 119.530 127.320 119.790 128.045 ;
        RECT 119.960 127.150 120.220 127.945 ;
        RECT 120.390 127.320 120.640 128.455 ;
        RECT 113.945 127.145 120.220 127.150 ;
        RECT 120.820 127.145 121.080 127.955 ;
        RECT 121.255 127.315 121.500 128.455 ;
        RECT 121.680 127.145 121.975 127.955 ;
        RECT 122.185 127.925 122.525 128.955 ;
        RECT 122.695 128.285 122.945 128.785 ;
        RECT 123.125 128.455 123.485 129.035 ;
        RECT 123.655 128.285 123.825 129.195 ;
        RECT 123.995 128.945 125.205 129.695 ;
        RECT 122.695 128.115 123.825 128.285 ;
        RECT 122.185 127.750 122.850 127.925 ;
        RECT 122.160 127.145 122.495 127.570 ;
        RECT 122.665 127.345 122.850 127.750 ;
        RECT 123.055 127.145 123.385 127.925 ;
        RECT 123.555 127.345 123.825 128.115 ;
        RECT 123.995 128.235 124.515 128.775 ;
        RECT 124.685 128.405 125.205 128.945 ;
        RECT 123.995 127.145 125.205 128.235 ;
        RECT 53.990 126.975 125.290 127.145 ;
        RECT 54.075 125.885 55.285 126.975 ;
        RECT 54.075 125.175 54.595 125.715 ;
        RECT 54.765 125.345 55.285 125.885 ;
        RECT 55.535 126.045 55.715 126.805 ;
        RECT 55.895 126.215 56.225 126.975 ;
        RECT 55.535 125.875 56.210 126.045 ;
        RECT 56.395 125.900 56.665 126.805 ;
        RECT 56.040 125.730 56.210 125.875 ;
        RECT 55.475 125.325 55.815 125.695 ;
        RECT 56.040 125.400 56.315 125.730 ;
        RECT 54.075 124.425 55.285 125.175 ;
        RECT 56.040 125.145 56.210 125.400 ;
        RECT 55.545 124.975 56.210 125.145 ;
        RECT 56.485 125.100 56.665 125.900 ;
        RECT 57.295 125.835 57.575 126.975 ;
        RECT 57.745 125.825 58.075 126.805 ;
        RECT 58.245 125.835 58.505 126.975 ;
        RECT 58.685 126.175 59.015 126.975 ;
        RECT 59.195 126.635 60.625 126.805 ;
        RECT 59.195 126.005 59.445 126.635 ;
        RECT 58.675 125.835 59.445 126.005 ;
        RECT 57.810 125.785 57.985 125.825 ;
        RECT 57.305 125.395 57.640 125.665 ;
        RECT 57.810 125.225 57.980 125.785 ;
        RECT 58.150 125.415 58.485 125.665 ;
        RECT 55.545 124.595 55.715 124.975 ;
        RECT 55.895 124.425 56.225 124.805 ;
        RECT 56.405 124.595 56.665 125.100 ;
        RECT 57.295 124.425 57.605 125.225 ;
        RECT 57.810 124.595 58.505 125.225 ;
        RECT 58.675 125.165 58.845 125.835 ;
        RECT 59.015 125.335 59.420 125.665 ;
        RECT 59.635 125.335 59.885 126.465 ;
        RECT 60.085 125.665 60.285 126.465 ;
        RECT 60.455 125.955 60.625 126.635 ;
        RECT 60.795 126.125 61.110 126.975 ;
        RECT 61.285 126.175 61.725 126.805 ;
        RECT 60.455 125.785 61.245 125.955 ;
        RECT 60.085 125.335 60.330 125.665 ;
        RECT 60.515 125.335 60.905 125.615 ;
        RECT 61.075 125.335 61.245 125.785 ;
        RECT 61.415 125.165 61.725 126.175 ;
        RECT 58.675 124.595 59.165 125.165 ;
        RECT 59.335 124.995 60.495 125.165 ;
        RECT 59.335 124.595 59.565 124.995 ;
        RECT 59.735 124.425 60.155 124.825 ;
        RECT 60.325 124.595 60.495 124.995 ;
        RECT 60.665 124.425 61.115 125.165 ;
        RECT 61.285 124.605 61.725 125.165 ;
        RECT 62.355 126.135 62.615 126.805 ;
        RECT 62.785 126.575 63.115 126.975 ;
        RECT 63.985 126.575 64.385 126.975 ;
        RECT 64.675 126.395 65.005 126.630 ;
        RECT 62.925 126.225 65.005 126.395 ;
        RECT 62.355 126.125 62.585 126.135 ;
        RECT 62.355 125.165 62.530 126.125 ;
        RECT 62.925 125.955 63.095 126.225 ;
        RECT 62.700 125.785 63.095 125.955 ;
        RECT 63.265 125.835 64.280 126.055 ;
        RECT 62.700 125.335 62.870 125.785 ;
        RECT 64.005 125.695 64.280 125.835 ;
        RECT 64.450 125.835 65.005 126.225 ;
        RECT 63.040 125.415 63.490 125.615 ;
        RECT 63.660 125.245 63.835 125.440 ;
        RECT 62.355 124.595 62.695 125.165 ;
        RECT 62.890 124.425 63.060 125.090 ;
        RECT 63.340 125.075 63.835 125.245 ;
        RECT 63.340 124.935 63.560 125.075 ;
        RECT 63.335 124.765 63.560 124.935 ;
        RECT 64.005 124.905 64.175 125.695 ;
        RECT 64.450 125.585 64.620 125.835 ;
        RECT 65.175 125.665 65.350 126.765 ;
        RECT 65.520 126.155 65.865 126.975 ;
        RECT 64.425 125.415 64.620 125.585 ;
        RECT 64.790 125.415 65.350 125.665 ;
        RECT 65.520 125.415 65.865 125.985 ;
        RECT 66.955 125.810 67.245 126.975 ;
        RECT 67.415 125.900 67.685 126.805 ;
        RECT 67.855 126.215 68.185 126.975 ;
        RECT 68.365 126.045 68.545 126.805 ;
        RECT 64.425 125.030 64.595 125.415 ;
        RECT 63.340 124.720 63.560 124.765 ;
        RECT 63.730 124.735 64.175 124.905 ;
        RECT 64.345 124.660 64.595 125.030 ;
        RECT 64.765 125.065 65.865 125.245 ;
        RECT 64.765 124.660 65.015 125.065 ;
        RECT 65.185 124.425 65.355 124.895 ;
        RECT 65.525 124.660 65.865 125.065 ;
        RECT 66.955 124.425 67.245 125.150 ;
        RECT 67.415 125.100 67.595 125.900 ;
        RECT 67.870 125.875 68.545 126.045 ;
        RECT 67.870 125.730 68.040 125.875 ;
        RECT 67.765 125.400 68.040 125.730 ;
        RECT 68.800 125.835 69.135 126.805 ;
        RECT 69.305 125.835 69.475 126.975 ;
        RECT 69.645 126.635 71.675 126.805 ;
        RECT 67.870 125.145 68.040 125.400 ;
        RECT 68.265 125.325 68.605 125.695 ;
        RECT 68.800 125.165 68.970 125.835 ;
        RECT 69.645 125.665 69.815 126.635 ;
        RECT 69.140 125.335 69.395 125.665 ;
        RECT 69.620 125.335 69.815 125.665 ;
        RECT 69.985 126.295 71.110 126.465 ;
        RECT 69.225 125.165 69.395 125.335 ;
        RECT 69.985 125.165 70.155 126.295 ;
        RECT 67.415 124.595 67.675 125.100 ;
        RECT 67.870 124.975 68.535 125.145 ;
        RECT 67.855 124.425 68.185 124.805 ;
        RECT 68.365 124.595 68.535 124.975 ;
        RECT 68.800 124.595 69.055 125.165 ;
        RECT 69.225 124.995 70.155 125.165 ;
        RECT 70.325 125.955 71.335 126.125 ;
        RECT 70.325 125.155 70.495 125.955 ;
        RECT 70.700 125.275 70.975 125.755 ;
        RECT 70.695 125.105 70.975 125.275 ;
        RECT 69.980 124.960 70.155 124.995 ;
        RECT 69.225 124.425 69.555 124.825 ;
        RECT 69.980 124.595 70.510 124.960 ;
        RECT 70.700 124.595 70.975 125.105 ;
        RECT 71.145 124.595 71.335 125.955 ;
        RECT 71.505 125.970 71.675 126.635 ;
        RECT 71.845 126.215 72.015 126.975 ;
        RECT 72.250 126.215 72.765 126.625 ;
        RECT 71.505 125.780 72.255 125.970 ;
        RECT 72.425 125.405 72.765 126.215 ;
        RECT 73.025 126.045 73.195 126.805 ;
        RECT 73.375 126.215 73.705 126.975 ;
        RECT 73.025 125.875 73.690 126.045 ;
        RECT 73.875 125.900 74.145 126.805 ;
        RECT 73.520 125.730 73.690 125.875 ;
        RECT 71.535 125.235 72.765 125.405 ;
        RECT 72.955 125.325 73.285 125.695 ;
        RECT 73.520 125.400 73.805 125.730 ;
        RECT 71.515 124.425 72.025 124.960 ;
        RECT 72.245 124.630 72.490 125.235 ;
        RECT 73.520 125.145 73.690 125.400 ;
        RECT 73.025 124.975 73.690 125.145 ;
        RECT 73.975 125.100 74.145 125.900 ;
        RECT 73.025 124.595 73.195 124.975 ;
        RECT 73.375 124.425 73.705 124.805 ;
        RECT 73.885 124.595 74.145 125.100 ;
        RECT 74.775 125.900 75.045 126.805 ;
        RECT 75.215 126.215 75.545 126.975 ;
        RECT 75.725 126.045 75.905 126.805 ;
        RECT 74.775 125.100 74.955 125.900 ;
        RECT 75.230 125.875 75.905 126.045 ;
        RECT 77.095 126.085 77.355 126.795 ;
        RECT 77.525 126.265 77.855 126.975 ;
        RECT 78.025 126.085 78.255 126.795 ;
        RECT 75.230 125.730 75.400 125.875 ;
        RECT 77.095 125.845 78.255 126.085 ;
        RECT 78.435 126.065 78.705 126.795 ;
        RECT 78.885 126.245 79.225 126.975 ;
        RECT 78.435 125.845 79.205 126.065 ;
        RECT 75.125 125.400 75.400 125.730 ;
        RECT 75.230 125.145 75.400 125.400 ;
        RECT 75.625 125.325 75.965 125.695 ;
        RECT 77.085 125.335 77.385 125.665 ;
        RECT 77.565 125.355 78.090 125.665 ;
        RECT 78.270 125.355 78.735 125.665 ;
        RECT 74.775 124.595 75.035 125.100 ;
        RECT 75.230 124.975 75.895 125.145 ;
        RECT 75.215 124.425 75.545 124.805 ;
        RECT 75.725 124.595 75.895 124.975 ;
        RECT 77.095 124.425 77.385 125.155 ;
        RECT 77.565 124.715 77.795 125.355 ;
        RECT 78.915 125.175 79.205 125.845 ;
        RECT 77.975 124.975 79.205 125.175 ;
        RECT 77.975 124.605 78.285 124.975 ;
        RECT 78.465 124.425 79.135 124.795 ;
        RECT 79.395 124.605 79.655 126.795 ;
        RECT 80.295 126.555 80.635 126.975 ;
        RECT 80.805 126.385 81.055 126.805 ;
        RECT 80.295 126.215 81.055 126.385 ;
        RECT 80.295 125.245 80.605 126.215 ;
        RECT 81.225 126.135 81.555 126.975 ;
        RECT 82.045 126.385 82.800 126.805 ;
        RECT 81.725 126.215 83.190 126.385 ;
        RECT 81.725 125.965 81.895 126.215 ;
        RECT 80.935 125.795 81.895 125.965 ;
        RECT 80.935 125.625 81.105 125.795 ;
        RECT 82.065 125.625 82.370 126.045 ;
        RECT 80.775 125.415 81.105 125.625 ;
        RECT 81.275 125.415 81.715 125.625 ;
        RECT 81.885 125.415 82.370 125.625 ;
        RECT 82.560 125.615 82.850 126.045 ;
        RECT 83.020 126.010 83.190 126.215 ;
        RECT 83.360 126.190 83.600 126.975 ;
        RECT 83.770 126.010 84.100 126.805 ;
        RECT 83.020 125.835 84.100 126.010 ;
        RECT 83.020 125.785 83.805 125.835 ;
        RECT 82.560 125.415 82.950 125.615 ;
        RECT 83.120 125.415 83.465 125.615 ;
        RECT 80.295 125.075 81.055 125.245 ;
        RECT 80.385 124.425 80.555 124.905 ;
        RECT 80.725 124.605 81.055 125.075 ;
        RECT 81.225 124.425 81.395 125.245 ;
        RECT 81.565 125.075 83.265 125.245 ;
        RECT 81.565 124.610 81.895 125.075 ;
        RECT 82.880 124.985 83.265 125.075 ;
        RECT 83.635 125.145 83.805 125.785 ;
        RECT 84.005 125.315 84.265 125.665 ;
        RECT 83.635 124.975 84.180 125.145 ;
        RECT 82.065 124.425 82.235 124.895 ;
        RECT 82.495 124.635 83.680 124.805 ;
        RECT 83.850 124.595 84.180 124.975 ;
        RECT 85.355 124.705 85.635 126.805 ;
        RECT 85.825 126.215 86.610 126.975 ;
        RECT 87.005 126.145 87.390 126.805 ;
        RECT 87.005 126.045 87.415 126.145 ;
        RECT 85.805 125.835 87.415 126.045 ;
        RECT 87.715 125.955 87.915 126.745 ;
        RECT 85.805 125.235 86.080 125.835 ;
        RECT 87.585 125.785 87.915 125.955 ;
        RECT 88.085 125.795 88.405 126.975 ;
        RECT 88.585 126.365 88.915 126.795 ;
        RECT 89.095 126.535 89.290 126.975 ;
        RECT 89.460 126.365 89.790 126.795 ;
        RECT 88.585 126.195 89.790 126.365 ;
        RECT 88.585 125.865 89.480 126.195 ;
        RECT 89.960 126.025 90.235 126.795 ;
        RECT 90.520 126.175 90.775 126.975 ;
        RECT 89.650 125.835 90.235 126.025 ;
        RECT 90.945 126.005 91.275 126.805 ;
        RECT 91.445 126.175 91.615 126.975 ;
        RECT 91.785 126.005 92.115 126.805 ;
        RECT 90.415 125.835 92.115 126.005 ;
        RECT 92.285 125.835 92.545 126.975 ;
        RECT 87.585 125.665 87.765 125.785 ;
        RECT 86.250 125.415 86.605 125.665 ;
        RECT 86.800 125.615 87.265 125.665 ;
        RECT 86.795 125.445 87.265 125.615 ;
        RECT 86.800 125.415 87.265 125.445 ;
        RECT 87.435 125.415 87.765 125.665 ;
        RECT 87.940 125.415 88.405 125.615 ;
        RECT 88.590 125.335 88.885 125.665 ;
        RECT 89.065 125.335 89.480 125.665 ;
        RECT 85.805 125.055 87.055 125.235 ;
        RECT 86.690 124.985 87.055 125.055 ;
        RECT 87.225 125.035 88.405 125.205 ;
        RECT 85.865 124.425 86.035 124.885 ;
        RECT 87.225 124.815 87.555 125.035 ;
        RECT 86.305 124.635 87.555 124.815 ;
        RECT 87.725 124.425 87.895 124.865 ;
        RECT 88.065 124.620 88.405 125.035 ;
        RECT 88.585 124.425 88.885 125.155 ;
        RECT 89.065 124.715 89.295 125.335 ;
        RECT 89.650 125.165 89.825 125.835 ;
        RECT 89.495 124.985 89.825 125.165 ;
        RECT 89.995 125.015 90.235 125.665 ;
        RECT 90.415 125.245 90.695 125.835 ;
        RECT 92.715 125.810 93.005 126.975 ;
        RECT 93.265 126.230 93.535 126.975 ;
        RECT 94.165 126.970 100.440 126.975 ;
        RECT 93.705 126.060 93.995 126.800 ;
        RECT 94.165 126.245 94.420 126.970 ;
        RECT 94.605 126.075 94.865 126.800 ;
        RECT 95.035 126.245 95.280 126.970 ;
        RECT 95.465 126.075 95.725 126.800 ;
        RECT 95.895 126.245 96.140 126.970 ;
        RECT 96.325 126.075 96.585 126.800 ;
        RECT 96.755 126.245 97.000 126.970 ;
        RECT 97.170 126.075 97.430 126.800 ;
        RECT 97.600 126.245 97.860 126.970 ;
        RECT 98.030 126.075 98.290 126.800 ;
        RECT 98.460 126.245 98.720 126.970 ;
        RECT 98.890 126.075 99.150 126.800 ;
        RECT 99.320 126.245 99.580 126.970 ;
        RECT 99.750 126.075 100.010 126.800 ;
        RECT 100.180 126.175 100.440 126.970 ;
        RECT 94.605 126.060 100.010 126.075 ;
        RECT 93.265 125.835 100.010 126.060 ;
        RECT 90.865 125.415 91.615 125.665 ;
        RECT 91.785 125.415 92.545 125.665 ;
        RECT 93.265 125.245 94.430 125.835 ;
        RECT 100.610 125.665 100.860 126.800 ;
        RECT 101.040 126.165 101.300 126.975 ;
        RECT 101.475 125.665 101.720 126.805 ;
        RECT 101.900 126.165 102.195 126.975 ;
        RECT 102.430 126.105 102.715 126.975 ;
        RECT 102.885 126.345 103.145 126.805 ;
        RECT 103.320 126.515 103.575 126.975 ;
        RECT 103.745 126.345 104.005 126.805 ;
        RECT 102.885 126.175 104.005 126.345 ;
        RECT 104.175 126.175 104.485 126.975 ;
        RECT 102.885 125.925 103.145 126.175 ;
        RECT 104.655 126.005 104.965 126.805 ;
        RECT 105.145 126.165 105.440 126.975 ;
        RECT 102.390 125.755 103.145 125.925 ;
        RECT 103.935 125.835 104.965 126.005 ;
        RECT 94.600 125.415 101.720 125.665 ;
        RECT 90.415 124.995 91.275 125.245 ;
        RECT 91.445 125.055 92.545 125.225 ;
        RECT 89.495 124.605 89.720 124.985 ;
        RECT 89.890 124.425 90.220 124.815 ;
        RECT 90.525 124.805 90.855 124.825 ;
        RECT 91.445 124.805 91.695 125.055 ;
        RECT 90.525 124.595 91.695 124.805 ;
        RECT 91.865 124.425 92.035 124.885 ;
        RECT 92.205 124.595 92.545 125.055 ;
        RECT 92.715 124.425 93.005 125.150 ;
        RECT 93.265 125.075 100.010 125.245 ;
        RECT 93.265 124.425 93.565 124.905 ;
        RECT 93.735 124.620 93.995 125.075 ;
        RECT 94.165 124.425 94.425 124.905 ;
        RECT 94.605 124.620 94.865 125.075 ;
        RECT 95.035 124.425 95.285 124.905 ;
        RECT 95.465 124.620 95.725 125.075 ;
        RECT 95.895 124.425 96.145 124.905 ;
        RECT 96.325 124.620 96.585 125.075 ;
        RECT 96.755 124.425 97.000 124.905 ;
        RECT 97.170 124.620 97.445 125.075 ;
        RECT 97.615 124.425 97.860 124.905 ;
        RECT 98.030 124.620 98.290 125.075 ;
        RECT 98.460 124.425 98.720 124.905 ;
        RECT 98.890 124.620 99.150 125.075 ;
        RECT 99.320 124.425 99.580 124.905 ;
        RECT 99.750 124.620 100.010 125.075 ;
        RECT 100.180 124.425 100.440 124.985 ;
        RECT 100.610 124.605 100.860 125.415 ;
        RECT 101.040 124.425 101.300 124.950 ;
        RECT 101.470 124.605 101.720 125.415 ;
        RECT 101.890 125.105 102.205 125.665 ;
        RECT 102.390 125.245 102.795 125.755 ;
        RECT 103.935 125.585 104.105 125.835 ;
        RECT 102.965 125.415 104.105 125.585 ;
        RECT 102.390 125.075 104.040 125.245 ;
        RECT 104.275 125.095 104.625 125.665 ;
        RECT 101.900 124.425 102.205 124.935 ;
        RECT 102.435 124.425 102.715 124.905 ;
        RECT 102.885 124.685 103.145 125.075 ;
        RECT 103.320 124.425 103.575 124.905 ;
        RECT 103.745 124.685 104.040 125.075 ;
        RECT 104.795 124.925 104.965 125.835 ;
        RECT 105.620 125.665 105.865 126.805 ;
        RECT 106.040 126.165 106.300 126.975 ;
        RECT 106.900 126.970 113.175 126.975 ;
        RECT 106.480 125.665 106.730 126.800 ;
        RECT 106.900 126.175 107.160 126.970 ;
        RECT 107.330 126.075 107.590 126.800 ;
        RECT 107.760 126.245 108.020 126.970 ;
        RECT 108.190 126.075 108.450 126.800 ;
        RECT 108.620 126.245 108.880 126.970 ;
        RECT 109.050 126.075 109.310 126.800 ;
        RECT 109.480 126.245 109.740 126.970 ;
        RECT 109.910 126.075 110.170 126.800 ;
        RECT 110.340 126.245 110.585 126.970 ;
        RECT 110.755 126.075 111.015 126.800 ;
        RECT 111.200 126.245 111.445 126.970 ;
        RECT 111.615 126.075 111.875 126.800 ;
        RECT 112.060 126.245 112.305 126.970 ;
        RECT 112.475 126.075 112.735 126.800 ;
        RECT 112.920 126.245 113.175 126.970 ;
        RECT 107.330 126.060 112.735 126.075 ;
        RECT 113.345 126.060 113.635 126.800 ;
        RECT 113.805 126.230 114.075 126.975 ;
        RECT 114.340 126.105 114.605 126.805 ;
        RECT 114.775 126.275 115.105 126.975 ;
        RECT 115.275 126.105 115.945 126.805 ;
        RECT 116.450 126.275 116.880 126.975 ;
        RECT 117.060 126.415 117.250 126.805 ;
        RECT 117.420 126.595 117.750 126.975 ;
        RECT 117.060 126.245 117.790 126.415 ;
        RECT 107.330 125.835 114.075 126.060 ;
        RECT 114.340 125.850 116.915 126.105 ;
        RECT 105.135 125.105 105.450 125.665 ;
        RECT 105.620 125.415 112.740 125.665 ;
        RECT 104.220 124.425 104.495 124.905 ;
        RECT 104.665 124.595 104.965 124.925 ;
        RECT 105.135 124.425 105.440 124.935 ;
        RECT 105.620 124.605 105.870 125.415 ;
        RECT 106.040 124.425 106.300 124.950 ;
        RECT 106.480 124.605 106.730 125.415 ;
        RECT 112.910 125.245 114.075 125.835 ;
        RECT 114.335 125.335 114.610 125.665 ;
        RECT 107.330 125.075 114.075 125.245 ;
        RECT 114.780 125.165 114.960 125.850 ;
        RECT 116.745 125.665 116.915 125.850 ;
        RECT 115.130 125.335 115.490 125.665 ;
        RECT 115.780 125.615 116.070 125.665 ;
        RECT 115.775 125.445 116.070 125.615 ;
        RECT 115.780 125.335 116.070 125.445 ;
        RECT 116.240 125.335 116.575 125.665 ;
        RECT 116.745 125.335 117.425 125.665 ;
        RECT 106.900 124.425 107.160 124.985 ;
        RECT 107.330 124.620 107.590 125.075 ;
        RECT 107.760 124.425 108.020 124.905 ;
        RECT 108.190 124.620 108.450 125.075 ;
        RECT 108.620 124.425 108.880 124.905 ;
        RECT 109.050 124.620 109.310 125.075 ;
        RECT 109.480 124.425 109.725 124.905 ;
        RECT 109.895 124.620 110.170 125.075 ;
        RECT 110.340 124.425 110.585 124.905 ;
        RECT 110.755 124.620 111.015 125.075 ;
        RECT 111.195 124.425 111.445 124.905 ;
        RECT 111.615 124.620 111.875 125.075 ;
        RECT 112.055 124.425 112.305 124.905 ;
        RECT 112.475 124.620 112.735 125.075 ;
        RECT 112.915 124.425 113.175 124.905 ;
        RECT 113.345 124.620 113.605 125.075 ;
        RECT 113.775 124.425 114.075 124.905 ;
        RECT 114.345 124.765 114.960 125.165 ;
        RECT 115.130 124.975 116.400 125.165 ;
        RECT 117.595 125.125 117.790 126.245 ;
        RECT 118.475 125.810 118.765 126.975 ;
        RECT 118.960 126.005 119.260 126.200 ;
        RECT 119.430 126.175 119.685 126.975 ;
        RECT 119.885 126.345 120.215 126.805 ;
        RECT 120.385 126.515 120.960 126.975 ;
        RECT 121.130 126.345 121.485 126.805 ;
        RECT 119.885 126.175 121.485 126.345 ;
        RECT 118.960 125.835 120.210 126.005 ;
        RECT 118.960 125.180 119.130 125.835 ;
        RECT 119.305 125.335 119.650 125.665 ;
        RECT 119.880 125.415 120.210 125.835 ;
        RECT 120.380 125.245 120.660 126.175 ;
        RECT 120.840 125.615 121.030 125.995 ;
        RECT 121.210 125.835 121.485 126.175 ;
        RECT 121.655 125.835 121.985 126.975 ;
        RECT 122.165 126.005 122.495 126.790 ;
        RECT 122.165 125.835 122.845 126.005 ;
        RECT 123.025 125.835 123.355 126.975 ;
        RECT 123.995 125.885 125.205 126.975 ;
        RECT 120.840 125.415 121.985 125.615 ;
        RECT 122.155 125.415 122.505 125.665 ;
        RECT 116.970 124.955 117.790 125.125 ;
        RECT 114.345 124.595 114.680 124.765 ;
        RECT 115.640 124.425 115.975 124.805 ;
        RECT 116.565 124.425 116.800 124.865 ;
        RECT 116.970 124.595 117.300 124.955 ;
        RECT 117.470 124.425 117.800 124.785 ;
        RECT 118.475 124.425 118.765 125.150 ;
        RECT 118.960 124.850 119.195 125.180 ;
        RECT 119.365 124.425 119.695 125.165 ;
        RECT 119.930 124.805 120.205 125.245 ;
        RECT 120.380 125.145 120.705 125.245 ;
        RECT 120.375 124.975 120.705 125.145 ;
        RECT 120.875 125.035 121.985 125.245 ;
        RECT 122.675 125.235 122.845 125.835 ;
        RECT 123.015 125.415 123.365 125.665 ;
        RECT 123.995 125.345 124.515 125.885 ;
        RECT 120.875 124.805 121.125 125.035 ;
        RECT 119.930 124.595 121.125 124.805 ;
        RECT 121.295 124.425 121.465 124.865 ;
        RECT 121.635 124.595 121.985 125.035 ;
        RECT 122.175 124.425 122.415 125.235 ;
        RECT 122.585 124.595 122.915 125.235 ;
        RECT 123.085 124.425 123.355 125.235 ;
        RECT 124.685 125.175 125.205 125.715 ;
        RECT 123.995 124.425 125.205 125.175 ;
        RECT 53.990 124.255 125.290 124.425 ;
        RECT 54.075 123.505 55.285 124.255 ;
        RECT 56.375 123.580 56.635 124.085 ;
        RECT 56.815 123.875 57.145 124.255 ;
        RECT 57.325 123.705 57.495 124.085 ;
        RECT 54.075 122.965 54.595 123.505 ;
        RECT 54.765 122.795 55.285 123.335 ;
        RECT 54.075 121.705 55.285 122.795 ;
        RECT 56.375 122.780 56.545 123.580 ;
        RECT 56.830 123.535 57.495 123.705 ;
        RECT 57.755 123.580 58.015 124.085 ;
        RECT 58.195 123.875 58.525 124.255 ;
        RECT 58.705 123.705 58.875 124.085 ;
        RECT 56.830 123.280 57.000 123.535 ;
        RECT 56.715 122.950 57.000 123.280 ;
        RECT 57.235 122.985 57.565 123.355 ;
        RECT 56.830 122.805 57.000 122.950 ;
        RECT 56.375 121.875 56.645 122.780 ;
        RECT 56.830 122.635 57.495 122.805 ;
        RECT 56.815 121.705 57.145 122.465 ;
        RECT 57.325 121.875 57.495 122.635 ;
        RECT 57.755 122.780 57.935 123.580 ;
        RECT 58.210 123.535 58.875 123.705 ;
        RECT 59.135 123.755 59.395 124.085 ;
        RECT 59.605 123.775 59.880 124.255 ;
        RECT 58.210 123.280 58.380 123.535 ;
        RECT 58.105 122.950 58.380 123.280 ;
        RECT 58.605 122.985 58.945 123.355 ;
        RECT 58.210 122.805 58.380 122.950 ;
        RECT 59.135 122.845 59.305 123.755 ;
        RECT 60.090 123.685 60.295 124.085 ;
        RECT 60.465 123.855 60.800 124.255 ;
        RECT 59.475 123.015 59.835 123.595 ;
        RECT 60.090 123.515 60.775 123.685 ;
        RECT 60.015 122.845 60.265 123.345 ;
        RECT 57.755 121.875 58.025 122.780 ;
        RECT 58.210 122.635 58.885 122.805 ;
        RECT 58.195 121.705 58.525 122.465 ;
        RECT 58.705 121.875 58.885 122.635 ;
        RECT 59.135 122.675 60.265 122.845 ;
        RECT 59.135 121.905 59.405 122.675 ;
        RECT 60.435 122.485 60.775 123.515 ;
        RECT 60.995 123.445 61.235 124.255 ;
        RECT 61.405 123.445 61.735 124.085 ;
        RECT 61.905 123.445 62.175 124.255 ;
        RECT 62.355 123.580 62.615 124.085 ;
        RECT 62.795 123.875 63.125 124.255 ;
        RECT 63.305 123.705 63.475 124.085 ;
        RECT 60.975 123.015 61.325 123.265 ;
        RECT 61.495 122.845 61.665 123.445 ;
        RECT 61.835 123.015 62.185 123.265 ;
        RECT 59.575 121.705 59.905 122.485 ;
        RECT 60.110 122.310 60.775 122.485 ;
        RECT 60.985 122.675 61.665 122.845 ;
        RECT 60.110 121.905 60.295 122.310 ;
        RECT 60.465 121.705 60.800 122.130 ;
        RECT 60.985 121.890 61.315 122.675 ;
        RECT 61.845 121.705 62.175 122.845 ;
        RECT 62.355 122.780 62.535 123.580 ;
        RECT 62.810 123.535 63.475 123.705 ;
        RECT 63.825 123.705 63.995 124.085 ;
        RECT 64.175 123.875 64.505 124.255 ;
        RECT 63.825 123.535 64.490 123.705 ;
        RECT 64.685 123.580 64.945 124.085 ;
        RECT 62.810 123.280 62.980 123.535 ;
        RECT 62.705 122.950 62.980 123.280 ;
        RECT 63.205 122.985 63.545 123.355 ;
        RECT 63.755 122.985 64.095 123.355 ;
        RECT 64.320 123.280 64.490 123.535 ;
        RECT 62.810 122.805 62.980 122.950 ;
        RECT 64.320 122.950 64.595 123.280 ;
        RECT 64.320 122.805 64.490 122.950 ;
        RECT 62.355 121.875 62.625 122.780 ;
        RECT 62.810 122.635 63.485 122.805 ;
        RECT 62.795 121.705 63.125 122.465 ;
        RECT 63.305 121.875 63.485 122.635 ;
        RECT 63.815 122.635 64.490 122.805 ;
        RECT 64.765 122.780 64.945 123.580 ;
        RECT 65.205 123.705 65.375 124.085 ;
        RECT 65.555 123.875 65.885 124.255 ;
        RECT 65.205 123.535 65.870 123.705 ;
        RECT 66.065 123.580 66.325 124.085 ;
        RECT 65.135 122.985 65.475 123.355 ;
        RECT 65.700 123.280 65.870 123.535 ;
        RECT 65.700 122.950 65.975 123.280 ;
        RECT 65.700 122.805 65.870 122.950 ;
        RECT 63.815 121.875 63.995 122.635 ;
        RECT 64.175 121.705 64.505 122.465 ;
        RECT 64.675 121.875 64.945 122.780 ;
        RECT 65.195 122.635 65.870 122.805 ;
        RECT 66.145 122.780 66.325 123.580 ;
        RECT 66.535 123.435 66.765 124.255 ;
        RECT 66.935 123.455 67.265 124.085 ;
        RECT 66.515 123.015 66.845 123.265 ;
        RECT 67.015 122.855 67.265 123.455 ;
        RECT 67.435 123.435 67.645 124.255 ;
        RECT 67.875 123.580 68.135 124.085 ;
        RECT 68.315 123.875 68.645 124.255 ;
        RECT 68.825 123.705 68.995 124.085 ;
        RECT 65.195 121.875 65.375 122.635 ;
        RECT 65.555 121.705 65.885 122.465 ;
        RECT 66.055 121.875 66.325 122.780 ;
        RECT 66.535 121.705 66.765 122.845 ;
        RECT 66.935 121.875 67.265 122.855 ;
        RECT 67.435 121.705 67.645 122.845 ;
        RECT 67.875 122.780 68.055 123.580 ;
        RECT 68.330 123.535 68.995 123.705 ;
        RECT 68.330 123.280 68.500 123.535 ;
        RECT 70.175 123.455 70.485 124.255 ;
        RECT 70.690 123.455 71.385 124.085 ;
        RECT 71.555 123.710 76.900 124.255 ;
        RECT 68.225 122.950 68.500 123.280 ;
        RECT 68.725 122.985 69.065 123.355 ;
        RECT 70.185 123.015 70.520 123.285 ;
        RECT 68.330 122.805 68.500 122.950 ;
        RECT 70.690 122.855 70.860 123.455 ;
        RECT 71.030 123.015 71.365 123.265 ;
        RECT 73.140 122.880 73.480 123.710 ;
        RECT 77.075 123.485 79.665 124.255 ;
        RECT 79.835 123.530 80.125 124.255 ;
        RECT 80.295 123.495 81.005 124.085 ;
        RECT 81.515 123.725 81.845 124.085 ;
        RECT 82.045 123.895 82.375 124.255 ;
        RECT 82.545 123.725 82.875 124.085 ;
        RECT 81.515 123.515 82.875 123.725 ;
        RECT 83.055 123.580 83.315 124.085 ;
        RECT 83.495 123.875 83.825 124.255 ;
        RECT 84.005 123.705 84.175 124.085 ;
        RECT 67.875 121.875 68.145 122.780 ;
        RECT 68.330 122.635 69.005 122.805 ;
        RECT 68.315 121.705 68.645 122.465 ;
        RECT 68.825 121.875 69.005 122.635 ;
        RECT 70.175 121.705 70.455 122.845 ;
        RECT 70.625 121.875 70.955 122.855 ;
        RECT 71.125 121.705 71.385 122.845 ;
        RECT 74.960 122.140 75.310 123.390 ;
        RECT 77.075 122.965 78.285 123.485 ;
        RECT 78.455 122.795 79.665 123.315 ;
        RECT 71.555 121.705 76.900 122.140 ;
        RECT 77.075 121.705 79.665 122.795 ;
        RECT 79.835 121.705 80.125 122.870 ;
        RECT 80.295 122.525 80.500 123.495 ;
        RECT 80.670 122.725 81.000 123.265 ;
        RECT 81.175 123.015 81.670 123.345 ;
        RECT 81.990 123.015 82.365 123.345 ;
        RECT 82.575 123.015 82.885 123.345 ;
        RECT 81.175 122.725 81.500 123.015 ;
        RECT 81.695 122.525 82.025 122.745 ;
        RECT 80.295 122.295 82.025 122.525 ;
        RECT 80.295 121.875 80.995 122.295 ;
        RECT 81.195 121.705 81.525 122.065 ;
        RECT 81.695 121.895 82.025 122.295 ;
        RECT 82.195 122.045 82.365 123.015 ;
        RECT 83.055 122.780 83.235 123.580 ;
        RECT 83.510 123.535 84.175 123.705 ;
        RECT 84.435 123.580 84.695 124.085 ;
        RECT 84.875 123.875 85.205 124.255 ;
        RECT 85.385 123.705 85.555 124.085 ;
        RECT 83.510 123.280 83.680 123.535 ;
        RECT 83.405 122.950 83.680 123.280 ;
        RECT 83.905 122.985 84.245 123.355 ;
        RECT 83.510 122.805 83.680 122.950 ;
        RECT 82.545 121.705 82.875 122.765 ;
        RECT 83.055 121.875 83.325 122.780 ;
        RECT 83.510 122.635 84.185 122.805 ;
        RECT 83.495 121.705 83.825 122.465 ;
        RECT 84.005 121.875 84.185 122.635 ;
        RECT 84.435 122.780 84.615 123.580 ;
        RECT 84.890 123.535 85.555 123.705 ;
        RECT 85.905 123.705 86.075 124.085 ;
        RECT 86.255 123.875 86.585 124.255 ;
        RECT 85.905 123.535 86.570 123.705 ;
        RECT 86.765 123.580 87.025 124.085 ;
        RECT 84.890 123.280 85.060 123.535 ;
        RECT 84.785 122.950 85.060 123.280 ;
        RECT 85.285 122.985 85.625 123.355 ;
        RECT 85.835 122.985 86.175 123.355 ;
        RECT 86.400 123.280 86.570 123.535 ;
        RECT 84.890 122.805 85.060 122.950 ;
        RECT 86.400 122.950 86.675 123.280 ;
        RECT 86.400 122.805 86.570 122.950 ;
        RECT 84.435 121.875 84.705 122.780 ;
        RECT 84.890 122.635 85.565 122.805 ;
        RECT 84.875 121.705 85.205 122.465 ;
        RECT 85.385 121.875 85.565 122.635 ;
        RECT 85.895 122.635 86.570 122.805 ;
        RECT 86.845 122.780 87.025 123.580 ;
        RECT 85.895 121.875 86.075 122.635 ;
        RECT 86.255 121.705 86.585 122.465 ;
        RECT 86.755 121.875 87.025 122.780 ;
        RECT 87.195 123.580 87.455 124.085 ;
        RECT 87.635 123.875 87.965 124.255 ;
        RECT 88.145 123.705 88.315 124.085 ;
        RECT 87.195 122.780 87.375 123.580 ;
        RECT 87.650 123.535 88.315 123.705 ;
        RECT 88.575 123.580 88.835 124.085 ;
        RECT 89.015 123.875 89.345 124.255 ;
        RECT 89.525 123.705 89.695 124.085 ;
        RECT 87.650 123.280 87.820 123.535 ;
        RECT 87.545 122.950 87.820 123.280 ;
        RECT 88.045 122.985 88.385 123.355 ;
        RECT 87.650 122.805 87.820 122.950 ;
        RECT 87.195 121.875 87.465 122.780 ;
        RECT 87.650 122.635 88.325 122.805 ;
        RECT 87.635 121.705 87.965 122.465 ;
        RECT 88.145 121.875 88.325 122.635 ;
        RECT 88.575 122.780 88.755 123.580 ;
        RECT 89.030 123.535 89.695 123.705 ;
        RECT 89.030 123.280 89.200 123.535 ;
        RECT 89.960 123.490 90.415 124.255 ;
        RECT 90.690 123.875 91.990 124.085 ;
        RECT 92.245 123.895 92.575 124.255 ;
        RECT 91.820 123.725 91.990 123.875 ;
        RECT 92.745 123.755 93.005 124.085 ;
        RECT 88.925 122.950 89.200 123.280 ;
        RECT 89.425 122.985 89.765 123.355 ;
        RECT 90.890 123.265 91.110 123.665 ;
        RECT 89.955 123.065 90.445 123.265 ;
        RECT 90.635 123.055 91.110 123.265 ;
        RECT 91.355 123.265 91.565 123.665 ;
        RECT 91.820 123.600 92.575 123.725 ;
        RECT 91.820 123.555 92.665 123.600 ;
        RECT 92.395 123.435 92.665 123.555 ;
        RECT 91.355 123.055 91.685 123.265 ;
        RECT 91.855 122.995 92.265 123.300 ;
        RECT 89.030 122.805 89.200 122.950 ;
        RECT 89.960 122.825 91.135 122.885 ;
        RECT 92.495 122.860 92.665 123.435 ;
        RECT 92.465 122.825 92.665 122.860 ;
        RECT 88.575 121.875 88.845 122.780 ;
        RECT 89.030 122.635 89.705 122.805 ;
        RECT 89.015 121.705 89.345 122.465 ;
        RECT 89.525 121.875 89.705 122.635 ;
        RECT 89.960 122.715 92.665 122.825 ;
        RECT 89.960 122.095 90.215 122.715 ;
        RECT 90.805 122.655 92.605 122.715 ;
        RECT 90.805 122.625 91.135 122.655 ;
        RECT 92.835 122.555 93.005 123.755 ;
        RECT 90.465 122.455 90.650 122.545 ;
        RECT 91.240 122.455 92.075 122.465 ;
        RECT 90.465 122.255 92.075 122.455 ;
        RECT 90.465 122.215 90.695 122.255 ;
        RECT 89.960 121.875 90.295 122.095 ;
        RECT 91.300 121.705 91.655 122.085 ;
        RECT 91.825 121.875 92.075 122.255 ;
        RECT 92.325 121.705 92.575 122.485 ;
        RECT 92.745 121.875 93.005 122.555 ;
        RECT 93.175 123.435 93.860 124.075 ;
        RECT 94.030 123.435 94.200 124.255 ;
        RECT 94.370 123.605 94.700 124.070 ;
        RECT 94.870 123.785 95.040 124.255 ;
        RECT 95.300 123.865 96.485 124.035 ;
        RECT 96.655 123.695 96.985 124.085 ;
        RECT 95.685 123.605 96.070 123.695 ;
        RECT 94.370 123.435 96.070 123.605 ;
        RECT 96.475 123.515 96.985 123.695 ;
        RECT 97.315 123.755 97.575 124.085 ;
        RECT 97.745 123.895 98.075 124.255 ;
        RECT 98.330 123.875 99.630 124.085 ;
        RECT 93.175 122.465 93.425 123.435 ;
        RECT 93.595 123.055 93.930 123.265 ;
        RECT 94.100 123.055 94.550 123.265 ;
        RECT 94.740 123.055 95.225 123.265 ;
        RECT 93.760 122.885 93.930 123.055 ;
        RECT 94.850 122.895 95.225 123.055 ;
        RECT 95.415 123.015 95.795 123.265 ;
        RECT 95.975 123.055 96.305 123.265 ;
        RECT 93.760 122.715 94.680 122.885 ;
        RECT 93.175 121.875 93.840 122.465 ;
        RECT 94.010 121.705 94.340 122.545 ;
        RECT 94.510 122.465 94.680 122.715 ;
        RECT 94.850 122.725 95.245 122.895 ;
        RECT 94.850 122.635 95.225 122.725 ;
        RECT 95.415 122.635 95.735 123.015 ;
        RECT 96.475 122.885 96.645 123.515 ;
        RECT 96.815 123.055 97.145 123.345 ;
        RECT 95.905 122.715 96.990 122.885 ;
        RECT 95.905 122.465 96.075 122.715 ;
        RECT 94.510 122.295 96.075 122.465 ;
        RECT 94.850 121.875 95.655 122.295 ;
        RECT 96.245 121.705 96.495 122.545 ;
        RECT 96.690 121.875 96.990 122.715 ;
        RECT 97.315 122.555 97.485 123.755 ;
        RECT 98.330 123.725 98.500 123.875 ;
        RECT 97.745 123.600 98.500 123.725 ;
        RECT 97.655 123.555 98.500 123.600 ;
        RECT 97.655 123.435 97.925 123.555 ;
        RECT 97.655 122.860 97.825 123.435 ;
        RECT 98.055 122.995 98.465 123.300 ;
        RECT 98.755 123.265 98.965 123.665 ;
        RECT 98.635 123.055 98.965 123.265 ;
        RECT 99.210 123.265 99.430 123.665 ;
        RECT 99.905 123.490 100.360 124.255 ;
        RECT 99.210 123.055 99.685 123.265 ;
        RECT 99.875 123.065 100.365 123.265 ;
        RECT 97.655 122.825 97.855 122.860 ;
        RECT 99.185 122.825 100.360 122.885 ;
        RECT 97.655 122.715 100.360 122.825 ;
        RECT 97.715 122.655 99.515 122.715 ;
        RECT 99.185 122.625 99.515 122.655 ;
        RECT 97.315 121.875 97.575 122.555 ;
        RECT 97.745 121.705 97.995 122.485 ;
        RECT 98.245 122.455 99.080 122.465 ;
        RECT 99.670 122.455 99.855 122.545 ;
        RECT 98.245 122.255 99.855 122.455 ;
        RECT 98.245 121.875 98.495 122.255 ;
        RECT 99.625 122.215 99.855 122.255 ;
        RECT 100.105 122.095 100.360 122.715 ;
        RECT 98.665 121.705 99.020 122.085 ;
        RECT 100.025 121.875 100.360 122.095 ;
        RECT 101.470 121.885 101.750 124.075 ;
        RECT 101.950 123.885 102.680 124.255 ;
        RECT 103.260 123.715 103.690 124.075 ;
        RECT 101.950 123.525 103.690 123.715 ;
        RECT 101.950 123.015 102.210 123.525 ;
        RECT 101.940 121.705 102.225 122.845 ;
        RECT 102.420 122.725 102.680 123.345 ;
        RECT 102.875 122.725 103.300 123.345 ;
        RECT 103.470 123.295 103.690 123.525 ;
        RECT 103.860 123.475 104.105 124.255 ;
        RECT 103.470 122.995 104.015 123.295 ;
        RECT 104.305 123.175 104.535 124.075 ;
        RECT 102.490 122.355 103.515 122.555 ;
        RECT 102.490 121.885 102.660 122.355 ;
        RECT 102.835 121.705 103.165 122.185 ;
        RECT 103.335 121.885 103.515 122.355 ;
        RECT 103.685 121.885 104.015 122.995 ;
        RECT 104.195 122.495 104.535 123.175 ;
        RECT 104.715 122.675 104.945 124.015 ;
        RECT 105.595 123.530 105.885 124.255 ;
        RECT 106.505 123.775 106.675 124.255 ;
        RECT 106.845 123.605 107.175 124.080 ;
        RECT 107.345 123.775 107.515 124.255 ;
        RECT 107.685 123.605 108.015 124.080 ;
        RECT 108.185 123.775 108.355 124.255 ;
        RECT 108.525 123.605 108.855 124.080 ;
        RECT 109.025 123.775 109.195 124.255 ;
        RECT 109.365 123.605 109.695 124.080 ;
        RECT 109.865 123.775 110.035 124.255 ;
        RECT 110.205 123.605 110.535 124.080 ;
        RECT 110.705 123.775 110.875 124.255 ;
        RECT 111.045 123.605 111.375 124.080 ;
        RECT 106.055 123.435 109.695 123.605 ;
        RECT 109.865 123.435 111.375 123.605 ;
        RECT 111.565 123.435 111.895 124.080 ;
        RECT 112.065 123.435 112.235 124.255 ;
        RECT 112.500 123.605 112.770 123.815 ;
        RECT 112.990 123.795 113.320 124.255 ;
        RECT 113.830 123.795 114.580 124.085 ;
        RECT 112.500 123.435 113.835 123.605 ;
        RECT 106.055 122.895 106.440 123.435 ;
        RECT 109.865 123.265 110.035 123.435 ;
        RECT 111.565 123.265 111.735 123.435 ;
        RECT 113.665 123.265 113.835 123.435 ;
        RECT 106.650 123.065 110.035 123.265 ;
        RECT 110.205 123.065 111.735 123.265 ;
        RECT 111.905 123.065 112.325 123.265 ;
        RECT 109.865 122.895 110.035 123.065 ;
        RECT 104.195 122.295 104.945 122.495 ;
        RECT 104.185 121.705 104.535 122.115 ;
        RECT 104.705 121.905 104.945 122.295 ;
        RECT 105.595 121.705 105.885 122.870 ;
        RECT 106.055 122.725 109.695 122.895 ;
        RECT 109.865 122.725 111.375 122.895 ;
        RECT 106.505 121.705 106.675 122.505 ;
        RECT 106.845 121.875 107.175 122.725 ;
        RECT 107.345 121.705 107.515 122.505 ;
        RECT 107.685 121.875 108.015 122.725 ;
        RECT 108.185 121.705 108.355 122.505 ;
        RECT 108.525 121.875 108.855 122.725 ;
        RECT 109.025 121.705 109.195 122.505 ;
        RECT 109.365 121.875 109.695 122.725 ;
        RECT 109.865 121.705 110.035 122.555 ;
        RECT 110.205 121.875 110.535 122.725 ;
        RECT 110.705 121.705 110.875 122.555 ;
        RECT 111.045 121.875 111.375 122.725 ;
        RECT 111.565 122.795 111.735 123.065 ;
        RECT 112.500 123.025 112.850 123.265 ;
        RECT 113.020 123.025 113.495 123.265 ;
        RECT 113.665 123.015 114.040 123.265 ;
        RECT 111.565 121.875 111.895 122.795 ;
        RECT 112.065 121.705 112.235 122.895 ;
        RECT 113.665 122.845 113.835 123.015 ;
        RECT 112.500 122.675 113.835 122.845 ;
        RECT 112.500 122.515 112.780 122.675 ;
        RECT 114.210 122.505 114.580 123.795 ;
        RECT 114.885 123.775 115.185 124.255 ;
        RECT 115.355 123.605 115.615 124.060 ;
        RECT 115.785 123.775 116.045 124.255 ;
        RECT 116.225 123.605 116.485 124.060 ;
        RECT 116.655 123.775 116.905 124.255 ;
        RECT 117.085 123.605 117.345 124.060 ;
        RECT 117.515 123.775 117.765 124.255 ;
        RECT 117.945 123.605 118.205 124.060 ;
        RECT 118.375 123.775 118.620 124.255 ;
        RECT 118.790 123.605 119.065 124.060 ;
        RECT 119.235 123.775 119.480 124.255 ;
        RECT 119.650 123.605 119.910 124.060 ;
        RECT 120.080 123.775 120.340 124.255 ;
        RECT 120.510 123.605 120.770 124.060 ;
        RECT 120.940 123.775 121.200 124.255 ;
        RECT 121.370 123.605 121.630 124.060 ;
        RECT 121.800 123.695 122.060 124.255 ;
        RECT 114.885 123.435 121.630 123.605 ;
        RECT 114.885 122.845 116.050 123.435 ;
        RECT 122.230 123.265 122.480 124.075 ;
        RECT 122.660 123.730 122.920 124.255 ;
        RECT 123.090 123.265 123.340 124.075 ;
        RECT 123.520 123.745 123.825 124.255 ;
        RECT 116.220 123.015 123.340 123.265 ;
        RECT 123.510 123.015 123.825 123.575 ;
        RECT 123.995 123.505 125.205 124.255 ;
        RECT 114.885 122.620 121.630 122.845 ;
        RECT 112.990 121.705 113.240 122.505 ;
        RECT 113.410 122.335 114.580 122.505 ;
        RECT 113.410 121.875 113.740 122.335 ;
        RECT 113.910 121.705 114.125 122.165 ;
        RECT 114.885 121.705 115.155 122.450 ;
        RECT 115.325 121.880 115.615 122.620 ;
        RECT 116.225 122.605 121.630 122.620 ;
        RECT 115.785 121.710 116.040 122.435 ;
        RECT 116.225 121.880 116.485 122.605 ;
        RECT 116.655 121.710 116.900 122.435 ;
        RECT 117.085 121.880 117.345 122.605 ;
        RECT 117.515 121.710 117.760 122.435 ;
        RECT 117.945 121.880 118.205 122.605 ;
        RECT 118.375 121.710 118.620 122.435 ;
        RECT 118.790 121.880 119.050 122.605 ;
        RECT 119.220 121.710 119.480 122.435 ;
        RECT 119.650 121.880 119.910 122.605 ;
        RECT 120.080 121.710 120.340 122.435 ;
        RECT 120.510 121.880 120.770 122.605 ;
        RECT 120.940 121.710 121.200 122.435 ;
        RECT 121.370 121.880 121.630 122.605 ;
        RECT 121.800 121.710 122.060 122.505 ;
        RECT 122.230 121.880 122.480 123.015 ;
        RECT 115.785 121.705 122.060 121.710 ;
        RECT 122.660 121.705 122.920 122.515 ;
        RECT 123.095 121.875 123.340 123.015 ;
        RECT 123.995 122.795 124.515 123.335 ;
        RECT 124.685 122.965 125.205 123.505 ;
        RECT 123.520 121.705 123.815 122.515 ;
        RECT 123.995 121.705 125.205 122.795 ;
        RECT 53.990 121.535 125.290 121.705 ;
        RECT 54.075 120.445 55.285 121.535 ;
        RECT 54.075 119.735 54.595 120.275 ;
        RECT 54.765 119.905 55.285 120.445 ;
        RECT 56.560 120.565 56.950 120.740 ;
        RECT 57.435 120.735 57.765 121.535 ;
        RECT 57.935 120.745 58.470 121.365 ;
        RECT 56.560 120.395 57.985 120.565 ;
        RECT 54.075 118.985 55.285 119.735 ;
        RECT 56.435 119.665 56.790 120.225 ;
        RECT 56.960 119.495 57.130 120.395 ;
        RECT 57.300 119.665 57.565 120.225 ;
        RECT 57.815 119.895 57.985 120.395 ;
        RECT 58.155 119.725 58.470 120.745 ;
        RECT 58.675 120.580 58.945 121.535 ;
        RECT 56.540 118.985 56.780 119.495 ;
        RECT 56.960 119.165 57.240 119.495 ;
        RECT 57.470 118.985 57.685 119.495 ;
        RECT 57.855 119.155 58.470 119.725 ;
        RECT 59.130 120.480 59.435 121.265 ;
        RECT 59.615 121.065 60.300 121.535 ;
        RECT 59.610 120.545 60.305 120.855 ;
        RECT 59.130 119.675 59.305 120.480 ;
        RECT 60.480 120.375 60.765 121.320 ;
        RECT 60.965 121.085 61.295 121.535 ;
        RECT 61.465 120.915 61.635 121.345 ;
        RECT 59.905 120.225 60.765 120.375 ;
        RECT 59.475 120.205 60.765 120.225 ;
        RECT 60.955 120.685 61.635 120.915 ;
        RECT 61.985 120.915 62.155 121.345 ;
        RECT 62.325 121.085 62.655 121.535 ;
        RECT 61.985 120.685 62.660 120.915 ;
        RECT 59.475 119.845 60.465 120.205 ;
        RECT 60.955 120.035 61.190 120.685 ;
        RECT 58.675 118.985 58.945 119.620 ;
        RECT 59.130 119.155 59.365 119.675 ;
        RECT 60.295 119.510 60.465 119.845 ;
        RECT 60.635 119.705 61.190 120.035 ;
        RECT 60.975 119.555 61.190 119.705 ;
        RECT 61.360 120.345 61.665 120.515 ;
        RECT 61.360 119.665 61.660 120.345 ;
        RECT 61.955 119.665 62.255 120.515 ;
        RECT 62.425 120.035 62.660 120.685 ;
        RECT 62.830 120.375 63.115 121.320 ;
        RECT 63.295 121.065 63.980 121.535 ;
        RECT 63.290 120.545 63.985 120.855 ;
        RECT 64.160 120.480 64.465 121.265 ;
        RECT 62.830 120.225 63.690 120.375 ;
        RECT 62.830 120.205 64.115 120.225 ;
        RECT 62.425 119.705 62.960 120.035 ;
        RECT 63.130 119.845 64.115 120.205 ;
        RECT 62.425 119.555 62.645 119.705 ;
        RECT 59.535 118.985 59.935 119.480 ;
        RECT 60.295 119.315 60.695 119.510 ;
        RECT 60.525 119.170 60.695 119.315 ;
        RECT 60.975 119.180 61.215 119.555 ;
        RECT 61.385 118.985 61.715 119.490 ;
        RECT 61.900 118.985 62.235 119.490 ;
        RECT 62.405 119.180 62.645 119.555 ;
        RECT 63.130 119.510 63.300 119.845 ;
        RECT 64.290 119.675 64.465 120.480 ;
        RECT 65.125 120.925 65.455 121.355 ;
        RECT 65.635 121.095 65.830 121.535 ;
        RECT 66.000 120.925 66.330 121.355 ;
        RECT 65.125 120.755 66.330 120.925 ;
        RECT 65.125 120.425 66.020 120.755 ;
        RECT 66.500 120.585 66.775 121.355 ;
        RECT 66.190 120.395 66.775 120.585 ;
        RECT 65.130 119.895 65.425 120.225 ;
        RECT 65.605 119.895 66.020 120.225 ;
        RECT 62.925 119.315 63.300 119.510 ;
        RECT 62.925 119.170 63.095 119.315 ;
        RECT 63.660 118.985 64.055 119.480 ;
        RECT 64.225 119.155 64.465 119.675 ;
        RECT 65.125 118.985 65.425 119.715 ;
        RECT 65.605 119.275 65.835 119.895 ;
        RECT 66.190 119.725 66.365 120.395 ;
        RECT 66.955 120.370 67.245 121.535 ;
        RECT 68.345 120.475 68.675 121.325 ;
        RECT 68.345 120.345 68.565 120.475 ;
        RECT 68.845 120.395 69.095 121.535 ;
        RECT 69.285 120.895 69.535 121.315 ;
        RECT 69.765 121.065 70.095 121.535 ;
        RECT 70.325 120.895 70.575 121.315 ;
        RECT 69.285 120.725 70.575 120.895 ;
        RECT 70.755 120.895 71.085 121.325 ;
        RECT 70.755 120.725 71.210 120.895 ;
        RECT 66.035 119.545 66.365 119.725 ;
        RECT 66.535 119.575 66.775 120.225 ;
        RECT 68.345 119.710 68.535 120.345 ;
        RECT 69.275 120.225 69.490 120.555 ;
        RECT 68.705 119.895 69.015 120.225 ;
        RECT 69.185 119.895 69.490 120.225 ;
        RECT 69.665 119.895 69.950 120.555 ;
        RECT 70.145 119.895 70.410 120.555 ;
        RECT 70.625 119.895 70.870 120.555 ;
        RECT 68.845 119.725 69.015 119.895 ;
        RECT 71.040 119.725 71.210 120.725 ;
        RECT 71.560 120.395 71.880 121.535 ;
        RECT 72.060 120.225 72.255 121.275 ;
        RECT 72.435 120.685 72.765 121.365 ;
        RECT 72.965 120.735 73.220 121.535 ;
        RECT 73.415 120.695 73.670 121.365 ;
        RECT 73.840 120.775 74.170 121.535 ;
        RECT 74.340 120.935 74.590 121.365 ;
        RECT 74.760 121.115 75.115 121.535 ;
        RECT 75.305 121.195 76.475 121.365 ;
        RECT 75.305 121.155 75.635 121.195 ;
        RECT 75.745 120.935 75.975 121.025 ;
        RECT 74.340 120.695 75.975 120.935 ;
        RECT 76.145 120.695 76.475 121.195 ;
        RECT 73.415 120.685 73.625 120.695 ;
        RECT 72.435 120.405 72.785 120.685 ;
        RECT 71.620 120.175 71.880 120.225 ;
        RECT 71.615 120.005 71.880 120.175 ;
        RECT 71.620 119.895 71.880 120.005 ;
        RECT 72.060 119.895 72.445 120.225 ;
        RECT 72.615 120.025 72.785 120.405 ;
        RECT 72.975 120.195 73.220 120.555 ;
        RECT 72.615 119.855 73.135 120.025 ;
        RECT 66.035 119.165 66.260 119.545 ;
        RECT 66.430 118.985 66.760 119.375 ;
        RECT 66.955 118.985 67.245 119.710 ;
        RECT 68.345 119.200 68.675 119.710 ;
        RECT 68.845 119.555 71.210 119.725 ;
        RECT 68.845 118.985 69.175 119.385 ;
        RECT 70.225 119.215 70.555 119.555 ;
        RECT 71.560 119.515 72.775 119.685 ;
        RECT 70.725 118.985 71.055 119.385 ;
        RECT 71.560 119.165 71.850 119.515 ;
        RECT 72.045 118.985 72.375 119.345 ;
        RECT 72.545 119.210 72.775 119.515 ;
        RECT 72.965 119.290 73.135 119.855 ;
        RECT 73.415 119.565 73.585 120.685 ;
        RECT 76.645 120.525 76.815 121.365 ;
        RECT 73.755 120.355 76.815 120.525 ;
        RECT 77.080 120.815 77.415 121.325 ;
        RECT 73.755 119.805 73.925 120.355 ;
        RECT 74.155 119.975 74.520 120.175 ;
        RECT 74.690 119.975 75.020 120.175 ;
        RECT 73.755 119.635 74.555 119.805 ;
        RECT 73.415 119.485 73.600 119.565 ;
        RECT 73.415 119.155 73.670 119.485 ;
        RECT 73.885 118.985 74.215 119.465 ;
        RECT 74.385 119.405 74.555 119.635 ;
        RECT 74.735 119.575 75.020 119.975 ;
        RECT 75.290 119.975 75.765 120.175 ;
        RECT 75.935 119.975 76.380 120.175 ;
        RECT 76.550 119.975 76.900 120.185 ;
        RECT 75.290 119.575 75.570 119.975 ;
        RECT 75.750 119.635 76.815 119.805 ;
        RECT 75.750 119.405 75.920 119.635 ;
        RECT 74.385 119.155 75.920 119.405 ;
        RECT 76.145 118.985 76.475 119.465 ;
        RECT 76.645 119.155 76.815 119.635 ;
        RECT 77.080 119.460 77.335 120.815 ;
        RECT 77.665 120.735 77.995 121.535 ;
        RECT 78.240 120.945 78.525 121.365 ;
        RECT 78.780 121.115 79.110 121.535 ;
        RECT 79.335 121.195 80.495 121.365 ;
        RECT 79.335 120.945 79.665 121.195 ;
        RECT 78.240 120.775 79.665 120.945 ;
        RECT 79.895 120.565 80.065 121.025 ;
        RECT 80.325 120.695 80.495 121.195 ;
        RECT 77.695 120.395 80.065 120.565 ;
        RECT 77.695 120.225 77.865 120.395 ;
        RECT 80.315 120.345 80.525 120.515 ;
        RECT 80.755 120.425 81.015 121.365 ;
        RECT 81.185 121.135 81.515 121.535 ;
        RECT 82.660 121.270 82.915 121.365 ;
        RECT 81.775 121.100 82.915 121.270 ;
        RECT 83.085 121.155 83.415 121.325 ;
        RECT 81.775 120.875 81.945 121.100 ;
        RECT 81.185 120.705 81.945 120.875 ;
        RECT 82.660 120.965 82.915 121.100 ;
        RECT 80.315 120.225 80.520 120.345 ;
        RECT 77.560 119.895 77.865 120.225 ;
        RECT 78.060 120.175 78.310 120.225 ;
        RECT 78.055 120.005 78.310 120.175 ;
        RECT 78.060 119.895 78.310 120.005 ;
        RECT 77.695 119.725 77.865 119.895 ;
        RECT 78.520 119.835 78.790 120.225 ;
        RECT 78.980 120.175 79.270 120.225 ;
        RECT 78.975 120.005 79.270 120.175 ;
        RECT 77.695 119.555 78.255 119.725 ;
        RECT 78.515 119.665 78.790 119.835 ;
        RECT 78.520 119.565 78.790 119.665 ;
        RECT 78.980 119.565 79.270 120.005 ;
        RECT 79.440 119.560 79.860 120.225 ;
        RECT 80.170 119.895 80.520 120.225 ;
        RECT 80.755 119.710 80.930 120.425 ;
        RECT 81.185 120.225 81.355 120.705 ;
        RECT 82.210 120.615 82.380 120.805 ;
        RECT 82.660 120.795 83.070 120.965 ;
        RECT 81.100 119.895 81.355 120.225 ;
        RECT 81.580 119.895 81.910 120.515 ;
        RECT 82.210 120.445 82.730 120.615 ;
        RECT 82.080 119.895 82.370 120.275 ;
        RECT 82.560 119.725 82.730 120.445 ;
        RECT 77.080 119.200 77.415 119.460 ;
        RECT 78.085 119.385 78.255 119.555 ;
        RECT 77.585 118.985 77.915 119.385 ;
        RECT 78.085 119.215 79.700 119.385 ;
        RECT 80.245 118.985 80.575 119.705 ;
        RECT 80.755 119.155 81.015 119.710 ;
        RECT 81.850 119.555 82.730 119.725 ;
        RECT 82.900 119.770 83.070 120.795 ;
        RECT 83.245 120.905 83.415 121.155 ;
        RECT 83.585 121.075 83.835 121.535 ;
        RECT 84.005 120.905 84.185 121.365 ;
        RECT 83.245 120.735 84.185 120.905 ;
        RECT 84.900 120.735 85.155 121.535 ;
        RECT 85.355 120.685 85.685 121.365 ;
        RECT 83.270 120.255 83.750 120.555 ;
        RECT 82.900 119.600 83.250 119.770 ;
        RECT 83.490 119.665 83.750 120.255 ;
        RECT 83.950 119.665 84.210 120.555 ;
        RECT 84.900 120.195 85.145 120.555 ;
        RECT 85.335 120.405 85.685 120.685 ;
        RECT 85.335 120.025 85.505 120.405 ;
        RECT 85.865 120.225 86.060 121.275 ;
        RECT 86.240 120.395 86.560 121.535 ;
        RECT 86.755 120.480 87.060 121.265 ;
        RECT 87.240 121.065 87.925 121.535 ;
        RECT 87.235 120.545 87.930 120.855 ;
        RECT 84.985 119.855 85.505 120.025 ;
        RECT 85.675 119.895 86.060 120.225 ;
        RECT 86.240 120.175 86.500 120.225 ;
        RECT 86.240 120.005 86.505 120.175 ;
        RECT 86.240 119.895 86.500 120.005 ;
        RECT 84.985 119.835 85.155 119.855 ;
        RECT 84.955 119.665 85.155 119.835 ;
        RECT 81.185 118.985 81.615 119.430 ;
        RECT 81.850 119.155 82.020 119.555 ;
        RECT 82.190 118.985 82.910 119.385 ;
        RECT 83.080 119.155 83.250 119.600 ;
        RECT 83.825 118.985 84.225 119.495 ;
        RECT 84.985 119.290 85.155 119.665 ;
        RECT 85.345 119.515 86.560 119.685 ;
        RECT 85.345 119.210 85.575 119.515 ;
        RECT 85.745 118.985 86.075 119.345 ;
        RECT 86.270 119.165 86.560 119.515 ;
        RECT 86.755 119.675 86.930 120.480 ;
        RECT 88.105 120.375 88.390 121.320 ;
        RECT 88.565 121.085 88.895 121.535 ;
        RECT 89.065 120.915 89.235 121.345 ;
        RECT 87.530 120.225 88.390 120.375 ;
        RECT 87.105 120.205 88.390 120.225 ;
        RECT 88.560 120.685 89.235 120.915 ;
        RECT 89.585 120.915 89.755 121.345 ;
        RECT 89.925 121.085 90.255 121.535 ;
        RECT 89.585 120.685 90.260 120.915 ;
        RECT 87.105 119.845 88.090 120.205 ;
        RECT 88.560 120.035 88.795 120.685 ;
        RECT 86.755 119.155 86.995 119.675 ;
        RECT 87.920 119.510 88.090 119.845 ;
        RECT 88.260 119.705 88.795 120.035 ;
        RECT 88.575 119.555 88.795 119.705 ;
        RECT 88.965 119.665 89.265 120.515 ;
        RECT 89.555 119.665 89.855 120.515 ;
        RECT 90.025 120.035 90.260 120.685 ;
        RECT 90.430 120.375 90.715 121.320 ;
        RECT 90.895 121.065 91.580 121.535 ;
        RECT 90.890 120.545 91.585 120.855 ;
        RECT 91.760 120.480 92.065 121.265 ;
        RECT 90.430 120.225 91.290 120.375 ;
        RECT 90.430 120.205 91.715 120.225 ;
        RECT 90.025 119.705 90.560 120.035 ;
        RECT 90.730 119.845 91.715 120.205 ;
        RECT 90.025 119.555 90.245 119.705 ;
        RECT 87.165 118.985 87.560 119.480 ;
        RECT 87.920 119.315 88.295 119.510 ;
        RECT 88.125 119.170 88.295 119.315 ;
        RECT 88.575 119.180 88.815 119.555 ;
        RECT 88.985 118.985 89.320 119.490 ;
        RECT 89.500 118.985 89.835 119.490 ;
        RECT 90.005 119.180 90.245 119.555 ;
        RECT 90.730 119.510 90.900 119.845 ;
        RECT 91.890 119.675 92.065 120.480 ;
        RECT 92.715 120.370 93.005 121.535 ;
        RECT 93.180 121.145 93.515 121.365 ;
        RECT 94.520 121.155 94.875 121.535 ;
        RECT 93.180 120.525 93.435 121.145 ;
        RECT 93.685 120.985 93.915 121.025 ;
        RECT 95.045 120.985 95.295 121.365 ;
        RECT 93.685 120.785 95.295 120.985 ;
        RECT 93.685 120.695 93.870 120.785 ;
        RECT 94.460 120.775 95.295 120.785 ;
        RECT 95.545 120.755 95.795 121.535 ;
        RECT 95.965 120.685 96.225 121.365 ;
        RECT 94.025 120.585 94.355 120.615 ;
        RECT 94.025 120.525 95.825 120.585 ;
        RECT 93.180 120.415 95.885 120.525 ;
        RECT 93.180 120.355 94.355 120.415 ;
        RECT 95.685 120.380 95.885 120.415 ;
        RECT 93.175 119.975 93.665 120.175 ;
        RECT 93.855 119.975 94.330 120.185 ;
        RECT 90.525 119.315 90.900 119.510 ;
        RECT 90.525 119.170 90.695 119.315 ;
        RECT 91.260 118.985 91.655 119.480 ;
        RECT 91.825 119.155 92.065 119.675 ;
        RECT 92.715 118.985 93.005 119.710 ;
        RECT 93.180 118.985 93.635 119.750 ;
        RECT 94.110 119.575 94.330 119.975 ;
        RECT 94.575 119.975 94.905 120.185 ;
        RECT 94.575 119.575 94.785 119.975 ;
        RECT 95.075 119.940 95.485 120.245 ;
        RECT 95.715 119.805 95.885 120.380 ;
        RECT 95.615 119.685 95.885 119.805 ;
        RECT 95.040 119.640 95.885 119.685 ;
        RECT 95.040 119.515 95.795 119.640 ;
        RECT 95.040 119.365 95.210 119.515 ;
        RECT 96.055 119.485 96.225 120.685 ;
        RECT 97.325 121.195 98.495 121.365 ;
        RECT 97.325 120.525 97.655 121.195 ;
        RECT 98.165 121.155 98.495 121.195 ;
        RECT 98.665 121.155 99.040 121.535 ;
        RECT 97.825 120.985 98.055 121.025 ;
        RECT 97.825 120.935 98.440 120.985 ;
        RECT 99.185 120.935 99.355 121.065 ;
        RECT 97.825 120.735 99.355 120.935 ;
        RECT 99.590 120.755 99.855 121.535 ;
        RECT 97.825 120.695 98.705 120.735 ;
        RECT 100.165 120.605 100.335 121.365 ;
        RECT 100.550 120.775 100.880 121.535 ;
        RECT 98.845 120.525 99.905 120.565 ;
        RECT 97.325 120.395 99.905 120.525 ;
        RECT 100.165 120.435 100.880 120.605 ;
        RECT 101.050 120.460 101.305 121.365 ;
        RECT 97.325 120.345 99.070 120.395 ;
        RECT 97.355 119.665 97.805 120.175 ;
        RECT 97.995 119.975 98.470 120.175 ;
        RECT 98.220 119.575 98.470 119.975 ;
        RECT 98.720 119.975 99.070 120.175 ;
        RECT 98.720 119.575 98.930 119.975 ;
        RECT 99.240 119.895 99.565 120.225 ;
        RECT 99.735 119.725 99.905 120.395 ;
        RECT 100.075 119.885 100.430 120.255 ;
        RECT 100.710 120.225 100.880 120.435 ;
        RECT 100.710 119.895 100.965 120.225 ;
        RECT 99.175 119.555 99.905 119.725 ;
        RECT 100.710 119.705 100.880 119.895 ;
        RECT 101.135 119.730 101.305 120.460 ;
        RECT 101.480 120.385 101.740 121.535 ;
        RECT 101.915 120.395 102.255 121.365 ;
        RECT 102.425 120.395 102.595 121.535 ;
        RECT 102.865 120.735 103.115 121.535 ;
        RECT 103.760 120.565 104.090 121.365 ;
        RECT 104.390 120.735 104.720 121.535 ;
        RECT 104.890 120.565 105.220 121.365 ;
        RECT 102.785 120.395 105.220 120.565 ;
        RECT 105.635 120.395 105.865 121.535 ;
        RECT 93.910 119.155 95.210 119.365 ;
        RECT 95.465 118.985 95.795 119.345 ;
        RECT 95.965 119.155 96.225 119.485 ;
        RECT 97.325 118.985 97.775 119.495 ;
        RECT 99.175 119.405 99.355 119.555 ;
        RECT 98.050 119.155 99.355 119.405 ;
        RECT 100.165 119.535 100.880 119.705 ;
        RECT 99.535 118.985 99.865 119.385 ;
        RECT 100.165 119.155 100.335 119.535 ;
        RECT 100.550 118.985 100.880 119.365 ;
        RECT 101.050 119.155 101.305 119.730 ;
        RECT 101.480 118.985 101.740 119.825 ;
        RECT 101.915 119.785 102.090 120.395 ;
        RECT 102.785 120.145 102.955 120.395 ;
        RECT 102.260 119.975 102.955 120.145 ;
        RECT 103.130 119.975 103.550 120.175 ;
        RECT 103.720 119.975 104.050 120.175 ;
        RECT 104.220 119.975 104.550 120.175 ;
        RECT 101.915 119.155 102.255 119.785 ;
        RECT 102.425 118.985 102.675 119.785 ;
        RECT 102.865 119.635 104.090 119.805 ;
        RECT 102.865 119.155 103.195 119.635 ;
        RECT 103.365 118.985 103.590 119.445 ;
        RECT 103.760 119.155 104.090 119.635 ;
        RECT 104.720 119.765 104.890 120.395 ;
        RECT 106.035 120.385 106.365 121.365 ;
        RECT 106.535 120.395 106.745 121.535 ;
        RECT 106.985 120.725 107.280 121.535 ;
        RECT 105.075 119.975 105.425 120.225 ;
        RECT 105.615 119.975 105.945 120.225 ;
        RECT 104.720 119.155 105.220 119.765 ;
        RECT 105.635 118.985 105.865 119.805 ;
        RECT 106.115 119.785 106.365 120.385 ;
        RECT 107.460 120.225 107.705 121.365 ;
        RECT 107.880 120.725 108.140 121.535 ;
        RECT 108.740 121.530 115.015 121.535 ;
        RECT 108.320 120.225 108.570 121.360 ;
        RECT 108.740 120.735 109.000 121.530 ;
        RECT 109.170 120.635 109.430 121.360 ;
        RECT 109.600 120.805 109.860 121.530 ;
        RECT 110.030 120.635 110.290 121.360 ;
        RECT 110.460 120.805 110.720 121.530 ;
        RECT 110.890 120.635 111.150 121.360 ;
        RECT 111.320 120.805 111.580 121.530 ;
        RECT 111.750 120.635 112.010 121.360 ;
        RECT 112.180 120.805 112.425 121.530 ;
        RECT 112.595 120.635 112.855 121.360 ;
        RECT 113.040 120.805 113.285 121.530 ;
        RECT 113.455 120.635 113.715 121.360 ;
        RECT 113.900 120.805 114.145 121.530 ;
        RECT 114.315 120.635 114.575 121.360 ;
        RECT 114.760 120.805 115.015 121.530 ;
        RECT 109.170 120.620 114.575 120.635 ;
        RECT 115.185 120.620 115.475 121.360 ;
        RECT 115.645 120.790 115.915 121.535 ;
        RECT 109.170 120.395 115.915 120.620 ;
        RECT 106.035 119.155 106.365 119.785 ;
        RECT 106.535 118.985 106.745 119.805 ;
        RECT 106.975 119.665 107.290 120.225 ;
        RECT 107.460 119.975 114.580 120.225 ;
        RECT 106.975 118.985 107.280 119.495 ;
        RECT 107.460 119.165 107.710 119.975 ;
        RECT 107.880 118.985 108.140 119.510 ;
        RECT 108.320 119.165 108.570 119.975 ;
        RECT 114.750 119.805 115.915 120.395 ;
        RECT 116.180 120.565 116.455 121.365 ;
        RECT 116.625 120.735 116.955 121.535 ;
        RECT 117.125 121.195 118.265 121.365 ;
        RECT 117.125 120.565 117.295 121.195 ;
        RECT 116.180 120.355 117.295 120.565 ;
        RECT 117.465 120.565 117.795 121.025 ;
        RECT 117.965 120.735 118.265 121.195 ;
        RECT 117.465 120.345 118.225 120.565 ;
        RECT 118.475 120.370 118.765 121.535 ;
        RECT 118.940 120.535 119.195 121.535 ;
        RECT 116.180 119.975 116.900 120.175 ;
        RECT 117.070 119.975 117.840 120.175 ;
        RECT 118.010 119.805 118.225 120.345 ;
        RECT 109.170 119.635 115.915 119.805 ;
        RECT 108.740 118.985 109.000 119.545 ;
        RECT 109.170 119.180 109.430 119.635 ;
        RECT 109.600 118.985 109.860 119.465 ;
        RECT 110.030 119.180 110.290 119.635 ;
        RECT 110.460 118.985 110.720 119.465 ;
        RECT 110.890 119.180 111.150 119.635 ;
        RECT 111.320 118.985 111.565 119.465 ;
        RECT 111.735 119.180 112.010 119.635 ;
        RECT 112.180 118.985 112.425 119.465 ;
        RECT 112.595 119.180 112.855 119.635 ;
        RECT 113.035 118.985 113.285 119.465 ;
        RECT 113.455 119.180 113.715 119.635 ;
        RECT 113.895 118.985 114.145 119.465 ;
        RECT 114.315 119.180 114.575 119.635 ;
        RECT 114.755 118.985 115.015 119.465 ;
        RECT 115.185 119.180 115.445 119.635 ;
        RECT 115.615 118.985 115.915 119.465 ;
        RECT 116.180 118.985 116.455 119.805 ;
        RECT 116.625 119.635 118.225 119.805 ;
        RECT 116.625 119.625 117.795 119.635 ;
        RECT 116.625 119.155 116.955 119.625 ;
        RECT 117.125 118.985 117.295 119.455 ;
        RECT 117.465 119.155 117.795 119.625 ;
        RECT 117.965 118.985 118.255 119.455 ;
        RECT 118.475 118.985 118.765 119.710 ;
        RECT 118.955 118.985 119.195 119.785 ;
        RECT 119.380 119.155 119.625 121.365 ;
        RECT 119.795 121.085 120.645 121.535 ;
        RECT 120.815 120.905 121.075 121.365 ;
        RECT 119.955 120.685 121.075 120.905 ;
        RECT 121.255 120.855 121.460 120.885 ;
        RECT 121.255 120.685 121.465 120.855 ;
        RECT 119.955 120.230 120.125 120.685 ;
        RECT 119.795 119.740 120.125 120.230 ;
        RECT 120.295 119.910 120.705 120.515 ;
        RECT 121.255 120.300 121.460 120.685 ;
        RECT 121.645 120.550 121.970 121.535 ;
        RECT 122.245 120.605 122.415 121.365 ;
        RECT 122.630 120.775 122.960 121.535 ;
        RECT 122.245 120.435 122.960 120.605 ;
        RECT 123.130 120.460 123.385 121.365 ;
        RECT 120.875 119.925 121.460 120.300 ;
        RECT 121.715 119.895 121.975 120.350 ;
        RECT 122.155 119.885 122.510 120.255 ;
        RECT 122.790 120.225 122.960 120.435 ;
        RECT 122.790 119.895 123.045 120.225 ;
        RECT 119.795 119.535 120.645 119.740 ;
        RECT 119.795 118.985 120.125 119.365 ;
        RECT 120.315 119.155 120.645 119.535 ;
        RECT 120.815 119.535 121.970 119.725 ;
        RECT 122.790 119.705 122.960 119.895 ;
        RECT 123.215 119.730 123.385 120.460 ;
        RECT 123.560 120.385 123.820 121.535 ;
        RECT 123.995 120.445 125.205 121.535 ;
        RECT 123.995 119.905 124.515 120.445 ;
        RECT 120.815 119.365 121.025 119.535 ;
        RECT 121.695 119.395 121.970 119.535 ;
        RECT 122.245 119.535 122.960 119.705 ;
        RECT 121.195 118.985 121.525 119.365 ;
        RECT 122.245 119.155 122.415 119.535 ;
        RECT 122.630 118.985 122.960 119.365 ;
        RECT 123.130 119.155 123.385 119.730 ;
        RECT 123.560 118.985 123.820 119.825 ;
        RECT 124.685 119.735 125.205 120.275 ;
        RECT 123.995 118.985 125.205 119.735 ;
        RECT 53.990 118.815 125.290 118.985 ;
        RECT 54.075 118.065 55.285 118.815 ;
        RECT 55.545 118.265 55.715 118.645 ;
        RECT 55.895 118.435 56.225 118.815 ;
        RECT 55.545 118.095 56.210 118.265 ;
        RECT 56.405 118.140 56.665 118.645 ;
        RECT 54.075 117.525 54.595 118.065 ;
        RECT 54.765 117.355 55.285 117.895 ;
        RECT 55.475 117.545 55.815 117.915 ;
        RECT 56.040 117.840 56.210 118.095 ;
        RECT 56.040 117.510 56.315 117.840 ;
        RECT 56.040 117.365 56.210 117.510 ;
        RECT 54.075 116.265 55.285 117.355 ;
        RECT 55.535 117.195 56.210 117.365 ;
        RECT 56.485 117.340 56.665 118.140 ;
        RECT 57.760 118.165 58.030 118.375 ;
        RECT 58.250 118.355 58.580 118.815 ;
        RECT 59.090 118.355 59.840 118.645 ;
        RECT 57.760 117.995 59.095 118.165 ;
        RECT 58.925 117.825 59.095 117.995 ;
        RECT 57.760 117.585 58.110 117.825 ;
        RECT 58.280 117.585 58.755 117.825 ;
        RECT 58.925 117.575 59.300 117.825 ;
        RECT 58.925 117.405 59.095 117.575 ;
        RECT 55.535 116.435 55.715 117.195 ;
        RECT 55.895 116.265 56.225 117.025 ;
        RECT 56.395 116.435 56.665 117.340 ;
        RECT 57.760 117.235 59.095 117.405 ;
        RECT 57.760 117.075 58.040 117.235 ;
        RECT 59.470 117.065 59.840 118.355 ;
        RECT 60.060 117.975 60.320 118.815 ;
        RECT 60.495 118.070 60.750 118.645 ;
        RECT 60.920 118.435 61.250 118.815 ;
        RECT 61.465 118.265 61.635 118.645 ;
        RECT 60.920 118.095 61.635 118.265 ;
        RECT 61.895 118.140 62.155 118.645 ;
        RECT 62.335 118.435 62.665 118.815 ;
        RECT 62.845 118.265 63.015 118.645 ;
        RECT 58.250 116.265 58.500 117.065 ;
        RECT 58.670 116.895 59.840 117.065 ;
        RECT 58.670 116.435 59.000 116.895 ;
        RECT 59.170 116.265 59.385 116.725 ;
        RECT 60.060 116.265 60.320 117.415 ;
        RECT 60.495 117.340 60.665 118.070 ;
        RECT 60.920 117.905 61.090 118.095 ;
        RECT 60.835 117.575 61.090 117.905 ;
        RECT 60.920 117.365 61.090 117.575 ;
        RECT 61.370 117.545 61.725 117.915 ;
        RECT 60.495 116.435 60.750 117.340 ;
        RECT 60.920 117.195 61.635 117.365 ;
        RECT 60.920 116.265 61.250 117.025 ;
        RECT 61.465 116.435 61.635 117.195 ;
        RECT 61.895 117.340 62.065 118.140 ;
        RECT 62.350 118.095 63.015 118.265 ;
        RECT 63.365 118.265 63.535 118.645 ;
        RECT 63.715 118.435 64.045 118.815 ;
        RECT 63.365 118.095 64.030 118.265 ;
        RECT 64.225 118.140 64.485 118.645 ;
        RECT 62.350 117.840 62.520 118.095 ;
        RECT 62.235 117.510 62.520 117.840 ;
        RECT 62.755 117.545 63.085 117.915 ;
        RECT 63.295 117.545 63.625 117.915 ;
        RECT 63.860 117.840 64.030 118.095 ;
        RECT 62.350 117.365 62.520 117.510 ;
        RECT 63.860 117.510 64.145 117.840 ;
        RECT 63.860 117.365 64.030 117.510 ;
        RECT 61.895 116.435 62.165 117.340 ;
        RECT 62.350 117.195 63.015 117.365 ;
        RECT 62.335 116.265 62.665 117.025 ;
        RECT 62.845 116.435 63.015 117.195 ;
        RECT 63.365 117.195 64.030 117.365 ;
        RECT 64.315 117.340 64.485 118.140 ;
        RECT 64.655 118.045 68.165 118.815 ;
        RECT 64.655 117.525 66.305 118.045 ;
        RECT 69.255 118.015 69.565 118.815 ;
        RECT 69.770 118.015 70.465 118.645 ;
        RECT 70.635 118.270 75.980 118.815 ;
        RECT 69.770 117.965 69.945 118.015 ;
        RECT 66.475 117.355 68.165 117.875 ;
        RECT 69.265 117.575 69.600 117.845 ;
        RECT 69.770 117.415 69.940 117.965 ;
        RECT 70.110 117.575 70.445 117.825 ;
        RECT 72.220 117.440 72.560 118.270 ;
        RECT 76.155 118.045 79.665 118.815 ;
        RECT 79.835 118.090 80.125 118.815 ;
        RECT 80.380 118.315 80.875 118.645 ;
        RECT 63.365 116.435 63.535 117.195 ;
        RECT 63.715 116.265 64.045 117.025 ;
        RECT 64.215 116.435 64.485 117.340 ;
        RECT 64.655 116.265 68.165 117.355 ;
        RECT 69.255 116.265 69.535 117.405 ;
        RECT 69.705 116.435 70.035 117.415 ;
        RECT 70.205 116.265 70.465 117.405 ;
        RECT 74.040 116.700 74.390 117.950 ;
        RECT 76.155 117.525 77.805 118.045 ;
        RECT 77.975 117.355 79.665 117.875 ;
        RECT 70.635 116.265 75.980 116.700 ;
        RECT 76.155 116.265 79.665 117.355 ;
        RECT 79.835 116.265 80.125 117.430 ;
        RECT 80.295 116.825 80.535 118.135 ;
        RECT 80.705 117.405 80.875 118.315 ;
        RECT 81.095 117.575 81.445 118.540 ;
        RECT 81.625 117.575 81.925 118.545 ;
        RECT 82.105 117.575 82.385 118.545 ;
        RECT 82.565 118.015 82.835 118.815 ;
        RECT 83.005 118.095 83.345 118.605 ;
        RECT 83.540 118.425 83.870 118.815 ;
        RECT 84.040 118.255 84.265 118.635 ;
        RECT 82.580 117.575 82.910 117.825 ;
        RECT 82.580 117.405 82.895 117.575 ;
        RECT 80.705 117.235 82.895 117.405 ;
        RECT 80.300 116.265 80.635 116.645 ;
        RECT 80.805 116.435 81.055 117.235 ;
        RECT 81.275 116.265 81.605 116.985 ;
        RECT 81.790 116.435 82.040 117.235 ;
        RECT 82.505 116.265 82.835 117.065 ;
        RECT 83.085 116.695 83.345 118.095 ;
        RECT 83.525 117.575 83.765 118.225 ;
        RECT 83.935 118.075 84.265 118.255 ;
        RECT 83.935 117.405 84.110 118.075 ;
        RECT 84.465 117.905 84.695 118.525 ;
        RECT 84.875 118.085 85.175 118.815 ;
        RECT 85.815 118.015 86.510 118.645 ;
        RECT 86.715 118.015 87.025 118.815 ;
        RECT 87.195 118.140 87.455 118.645 ;
        RECT 87.635 118.435 87.965 118.815 ;
        RECT 88.145 118.265 88.315 118.645 ;
        RECT 84.280 117.575 84.695 117.905 ;
        RECT 84.875 117.575 85.170 117.905 ;
        RECT 85.835 117.575 86.170 117.825 ;
        RECT 86.340 117.415 86.510 118.015 ;
        RECT 86.680 117.575 87.015 117.845 ;
        RECT 83.005 116.435 83.345 116.695 ;
        RECT 83.525 117.215 84.110 117.405 ;
        RECT 83.525 116.445 83.800 117.215 ;
        RECT 84.280 117.045 85.175 117.375 ;
        RECT 83.970 116.875 85.175 117.045 ;
        RECT 83.970 116.445 84.300 116.875 ;
        RECT 84.470 116.265 84.665 116.705 ;
        RECT 84.845 116.445 85.175 116.875 ;
        RECT 85.815 116.265 86.075 117.405 ;
        RECT 86.245 116.435 86.575 117.415 ;
        RECT 86.745 116.265 87.025 117.405 ;
        RECT 87.195 117.340 87.365 118.140 ;
        RECT 87.650 118.095 88.315 118.265 ;
        RECT 88.575 118.140 88.835 118.645 ;
        RECT 89.015 118.435 89.345 118.815 ;
        RECT 89.525 118.265 89.695 118.645 ;
        RECT 87.650 117.840 87.820 118.095 ;
        RECT 87.535 117.510 87.820 117.840 ;
        RECT 88.055 117.545 88.385 117.915 ;
        RECT 87.650 117.365 87.820 117.510 ;
        RECT 87.195 116.435 87.465 117.340 ;
        RECT 87.650 117.195 88.315 117.365 ;
        RECT 87.635 116.265 87.965 117.025 ;
        RECT 88.145 116.435 88.315 117.195 ;
        RECT 88.575 117.340 88.755 118.140 ;
        RECT 89.030 118.095 89.695 118.265 ;
        RECT 89.030 117.840 89.200 118.095 ;
        RECT 89.955 118.015 90.650 118.645 ;
        RECT 90.855 118.015 91.165 118.815 ;
        RECT 91.335 118.140 91.595 118.645 ;
        RECT 91.775 118.435 92.105 118.815 ;
        RECT 92.285 118.265 92.455 118.645 ;
        RECT 88.925 117.510 89.200 117.840 ;
        RECT 89.425 117.545 89.765 117.915 ;
        RECT 89.975 117.575 90.310 117.825 ;
        RECT 89.030 117.365 89.200 117.510 ;
        RECT 90.480 117.455 90.650 118.015 ;
        RECT 90.820 117.575 91.155 117.845 ;
        RECT 90.475 117.415 90.650 117.455 ;
        RECT 88.575 116.435 88.845 117.340 ;
        RECT 89.030 117.195 89.705 117.365 ;
        RECT 89.015 116.265 89.345 117.025 ;
        RECT 89.525 116.435 89.705 117.195 ;
        RECT 89.955 116.265 90.215 117.405 ;
        RECT 90.385 116.435 90.715 117.415 ;
        RECT 90.885 116.265 91.165 117.405 ;
        RECT 91.335 117.340 91.515 118.140 ;
        RECT 91.790 118.095 92.455 118.265 ;
        RECT 91.790 117.840 91.960 118.095 ;
        RECT 91.685 117.510 91.960 117.840 ;
        RECT 92.185 117.545 92.525 117.915 ;
        RECT 91.790 117.365 91.960 117.510 ;
        RECT 91.335 116.435 91.605 117.340 ;
        RECT 91.790 117.195 92.465 117.365 ;
        RECT 91.775 116.265 92.105 117.025 ;
        RECT 92.285 116.435 92.465 117.195 ;
        RECT 92.730 116.445 93.010 118.635 ;
        RECT 93.210 118.445 93.940 118.815 ;
        RECT 94.520 118.275 94.950 118.635 ;
        RECT 93.210 118.085 94.950 118.275 ;
        RECT 93.210 117.575 93.470 118.085 ;
        RECT 93.200 116.265 93.485 117.405 ;
        RECT 93.680 117.285 93.940 117.905 ;
        RECT 94.135 117.285 94.560 117.905 ;
        RECT 94.730 117.855 94.950 118.085 ;
        RECT 95.120 118.035 95.365 118.815 ;
        RECT 94.730 117.555 95.275 117.855 ;
        RECT 95.565 117.735 95.795 118.635 ;
        RECT 93.750 116.915 94.775 117.115 ;
        RECT 93.750 116.445 93.920 116.915 ;
        RECT 94.095 116.265 94.425 116.745 ;
        RECT 94.595 116.445 94.775 116.915 ;
        RECT 94.945 116.445 95.275 117.555 ;
        RECT 95.455 117.055 95.795 117.735 ;
        RECT 95.975 117.235 96.205 118.575 ;
        RECT 96.395 118.015 97.090 118.645 ;
        RECT 97.295 118.015 97.605 118.815 ;
        RECT 97.785 118.305 98.235 118.815 ;
        RECT 98.510 118.395 99.815 118.645 ;
        RECT 99.995 118.415 100.325 118.815 ;
        RECT 99.635 118.245 99.815 118.395 ;
        RECT 96.415 117.575 96.750 117.825 ;
        RECT 96.920 117.415 97.090 118.015 ;
        RECT 97.260 117.575 97.595 117.845 ;
        RECT 97.815 117.625 98.265 118.135 ;
        RECT 98.680 117.825 98.930 118.225 ;
        RECT 98.455 117.625 98.930 117.825 ;
        RECT 99.180 117.825 99.390 118.225 ;
        RECT 99.635 118.075 100.365 118.245 ;
        RECT 99.180 117.625 99.530 117.825 ;
        RECT 99.700 117.575 100.025 117.905 ;
        RECT 95.455 116.855 96.205 117.055 ;
        RECT 95.445 116.265 95.795 116.675 ;
        RECT 95.965 116.465 96.205 116.855 ;
        RECT 96.395 116.265 96.655 117.405 ;
        RECT 96.825 116.435 97.155 117.415 ;
        RECT 97.785 117.405 99.530 117.455 ;
        RECT 100.195 117.405 100.365 118.075 ;
        RECT 97.325 116.265 97.605 117.405 ;
        RECT 97.785 117.275 100.365 117.405 ;
        RECT 97.785 116.605 98.115 117.275 ;
        RECT 99.305 117.235 100.365 117.275 ;
        RECT 100.995 118.090 101.255 118.645 ;
        RECT 101.425 118.370 101.855 118.815 ;
        RECT 102.090 118.245 102.260 118.645 ;
        RECT 102.430 118.415 103.150 118.815 ;
        RECT 100.995 117.375 101.170 118.090 ;
        RECT 102.090 118.075 102.970 118.245 ;
        RECT 103.320 118.200 103.490 118.645 ;
        RECT 104.065 118.305 104.465 118.815 ;
        RECT 101.340 117.575 101.595 117.905 ;
        RECT 98.285 117.065 99.165 117.105 ;
        RECT 98.285 116.865 99.815 117.065 ;
        RECT 98.285 116.815 98.900 116.865 ;
        RECT 98.285 116.775 98.515 116.815 ;
        RECT 99.645 116.735 99.815 116.865 ;
        RECT 98.625 116.605 98.955 116.645 ;
        RECT 97.785 116.435 98.955 116.605 ;
        RECT 99.125 116.265 99.500 116.645 ;
        RECT 100.050 116.265 100.315 117.045 ;
        RECT 100.995 116.435 101.255 117.375 ;
        RECT 101.425 117.095 101.595 117.575 ;
        RECT 101.820 117.285 102.150 117.905 ;
        RECT 102.320 117.525 102.610 117.905 ;
        RECT 102.800 117.355 102.970 118.075 ;
        RECT 102.450 117.185 102.970 117.355 ;
        RECT 103.140 118.030 103.490 118.200 ;
        RECT 101.425 116.925 102.185 117.095 ;
        RECT 102.450 116.995 102.620 117.185 ;
        RECT 103.140 117.005 103.310 118.030 ;
        RECT 103.730 117.545 103.990 118.135 ;
        RECT 103.510 117.245 103.990 117.545 ;
        RECT 104.190 117.245 104.450 118.135 ;
        RECT 105.595 118.090 105.885 118.815 ;
        RECT 106.055 118.315 106.315 118.645 ;
        RECT 106.485 118.455 106.815 118.815 ;
        RECT 107.070 118.435 108.370 118.645 ;
        RECT 102.015 116.700 102.185 116.925 ;
        RECT 102.900 116.835 103.310 117.005 ;
        RECT 103.485 116.895 104.425 117.065 ;
        RECT 102.900 116.700 103.155 116.835 ;
        RECT 101.425 116.265 101.755 116.665 ;
        RECT 102.015 116.530 103.155 116.700 ;
        RECT 103.485 116.645 103.655 116.895 ;
        RECT 102.900 116.435 103.155 116.530 ;
        RECT 103.325 116.475 103.655 116.645 ;
        RECT 103.825 116.265 104.075 116.725 ;
        RECT 104.245 116.435 104.425 116.895 ;
        RECT 105.595 116.265 105.885 117.430 ;
        RECT 106.055 117.115 106.225 118.315 ;
        RECT 107.070 118.285 107.240 118.435 ;
        RECT 106.485 118.160 107.240 118.285 ;
        RECT 106.395 118.115 107.240 118.160 ;
        RECT 106.395 117.995 106.665 118.115 ;
        RECT 106.395 117.420 106.565 117.995 ;
        RECT 106.795 117.555 107.205 117.860 ;
        RECT 107.495 117.825 107.705 118.225 ;
        RECT 107.375 117.615 107.705 117.825 ;
        RECT 107.950 117.825 108.170 118.225 ;
        RECT 108.645 118.050 109.100 118.815 ;
        RECT 109.760 118.060 109.995 118.390 ;
        RECT 110.165 118.075 110.495 118.815 ;
        RECT 110.730 118.435 111.925 118.645 ;
        RECT 107.950 117.615 108.425 117.825 ;
        RECT 108.615 117.625 109.105 117.825 ;
        RECT 106.395 117.385 106.595 117.420 ;
        RECT 107.925 117.385 109.100 117.445 ;
        RECT 106.395 117.275 109.100 117.385 ;
        RECT 106.455 117.215 108.255 117.275 ;
        RECT 107.925 117.185 108.255 117.215 ;
        RECT 106.055 116.435 106.315 117.115 ;
        RECT 106.485 116.265 106.735 117.045 ;
        RECT 106.985 117.015 107.820 117.025 ;
        RECT 108.410 117.015 108.595 117.105 ;
        RECT 106.985 116.815 108.595 117.015 ;
        RECT 106.985 116.435 107.235 116.815 ;
        RECT 108.365 116.775 108.595 116.815 ;
        RECT 108.845 116.655 109.100 117.275 ;
        RECT 109.760 117.405 109.930 118.060 ;
        RECT 110.730 117.995 111.005 118.435 ;
        RECT 111.175 118.095 111.505 118.265 ;
        RECT 111.180 117.995 111.505 118.095 ;
        RECT 111.675 118.205 111.925 118.435 ;
        RECT 112.095 118.375 112.265 118.815 ;
        RECT 112.435 118.205 112.785 118.645 ;
        RECT 113.875 118.305 114.180 118.815 ;
        RECT 111.675 117.995 112.785 118.205 ;
        RECT 110.105 117.575 110.450 117.905 ;
        RECT 110.680 117.405 111.010 117.825 ;
        RECT 109.760 117.235 111.010 117.405 ;
        RECT 109.760 117.040 110.060 117.235 ;
        RECT 111.180 117.065 111.460 117.995 ;
        RECT 111.640 117.625 112.785 117.825 ;
        RECT 111.640 117.455 111.830 117.625 ;
        RECT 113.875 117.575 114.190 118.135 ;
        RECT 114.360 117.825 114.610 118.635 ;
        RECT 114.780 118.290 115.040 118.815 ;
        RECT 115.220 117.825 115.470 118.635 ;
        RECT 115.640 118.255 115.900 118.815 ;
        RECT 116.070 118.165 116.330 118.620 ;
        RECT 116.500 118.335 116.760 118.815 ;
        RECT 116.930 118.165 117.190 118.620 ;
        RECT 117.360 118.335 117.620 118.815 ;
        RECT 117.790 118.165 118.050 118.620 ;
        RECT 118.220 118.335 118.465 118.815 ;
        RECT 118.635 118.165 118.910 118.620 ;
        RECT 119.080 118.335 119.325 118.815 ;
        RECT 119.495 118.165 119.755 118.620 ;
        RECT 119.935 118.335 120.185 118.815 ;
        RECT 120.355 118.165 120.615 118.620 ;
        RECT 120.795 118.335 121.045 118.815 ;
        RECT 121.215 118.165 121.475 118.620 ;
        RECT 121.655 118.335 121.915 118.815 ;
        RECT 122.085 118.165 122.345 118.620 ;
        RECT 122.515 118.335 122.815 118.815 ;
        RECT 116.070 117.995 122.815 118.165 ;
        RECT 123.995 118.065 125.205 118.815 ;
        RECT 114.360 117.575 121.480 117.825 ;
        RECT 111.635 117.285 111.830 117.455 ;
        RECT 112.095 117.405 112.265 117.455 ;
        RECT 111.640 117.245 111.830 117.285 ;
        RECT 112.010 117.065 112.285 117.405 ;
        RECT 107.405 116.265 107.760 116.645 ;
        RECT 108.765 116.435 109.100 116.655 ;
        RECT 110.230 116.265 110.485 117.065 ;
        RECT 110.685 116.895 112.285 117.065 ;
        RECT 110.685 116.435 111.015 116.895 ;
        RECT 111.185 116.265 111.760 116.725 ;
        RECT 111.930 116.435 112.285 116.895 ;
        RECT 112.455 116.265 112.785 117.405 ;
        RECT 113.885 116.265 114.180 117.075 ;
        RECT 114.360 116.435 114.605 117.575 ;
        RECT 114.780 116.265 115.040 117.075 ;
        RECT 115.220 116.440 115.470 117.575 ;
        RECT 121.650 117.405 122.815 117.995 ;
        RECT 116.070 117.180 122.815 117.405 ;
        RECT 123.995 117.355 124.515 117.895 ;
        RECT 124.685 117.525 125.205 118.065 ;
        RECT 116.070 117.165 121.475 117.180 ;
        RECT 115.640 116.270 115.900 117.065 ;
        RECT 116.070 116.440 116.330 117.165 ;
        RECT 116.500 116.270 116.760 116.995 ;
        RECT 116.930 116.440 117.190 117.165 ;
        RECT 117.360 116.270 117.620 116.995 ;
        RECT 117.790 116.440 118.050 117.165 ;
        RECT 118.220 116.270 118.480 116.995 ;
        RECT 118.650 116.440 118.910 117.165 ;
        RECT 119.080 116.270 119.325 116.995 ;
        RECT 119.495 116.440 119.755 117.165 ;
        RECT 119.940 116.270 120.185 116.995 ;
        RECT 120.355 116.440 120.615 117.165 ;
        RECT 120.800 116.270 121.045 116.995 ;
        RECT 121.215 116.440 121.475 117.165 ;
        RECT 121.660 116.270 121.915 116.995 ;
        RECT 122.085 116.440 122.375 117.180 ;
        RECT 115.640 116.265 121.915 116.270 ;
        RECT 122.545 116.265 122.815 117.010 ;
        RECT 123.995 116.265 125.205 117.355 ;
        RECT 53.990 116.095 125.290 116.265 ;
        RECT 54.075 115.005 55.285 116.095 ;
        RECT 54.075 114.295 54.595 114.835 ;
        RECT 54.765 114.465 55.285 115.005 ;
        RECT 54.075 113.545 55.285 114.295 ;
        RECT 56.375 113.825 56.655 115.925 ;
        RECT 56.845 115.335 57.630 116.095 ;
        RECT 58.025 115.265 58.410 115.925 ;
        RECT 58.025 115.165 58.435 115.265 ;
        RECT 56.825 114.955 58.435 115.165 ;
        RECT 58.735 115.075 58.935 115.865 ;
        RECT 56.825 114.355 57.100 114.955 ;
        RECT 58.605 114.905 58.935 115.075 ;
        RECT 59.105 114.915 59.425 116.095 ;
        RECT 59.595 115.660 64.940 116.095 ;
        RECT 58.605 114.785 58.785 114.905 ;
        RECT 57.270 114.535 57.625 114.785 ;
        RECT 57.820 114.735 58.285 114.785 ;
        RECT 57.815 114.565 58.285 114.735 ;
        RECT 57.820 114.535 58.285 114.565 ;
        RECT 58.455 114.535 58.785 114.785 ;
        RECT 58.960 114.535 59.425 114.735 ;
        RECT 56.825 114.175 58.075 114.355 ;
        RECT 57.710 114.105 58.075 114.175 ;
        RECT 58.245 114.155 59.425 114.325 ;
        RECT 56.885 113.545 57.055 114.005 ;
        RECT 58.245 113.935 58.575 114.155 ;
        RECT 57.325 113.755 58.575 113.935 ;
        RECT 58.745 113.545 58.915 113.985 ;
        RECT 59.085 113.740 59.425 114.155 ;
        RECT 61.180 114.090 61.520 114.920 ;
        RECT 63.000 114.410 63.350 115.660 ;
        RECT 65.115 115.005 66.785 116.095 ;
        RECT 65.115 114.315 65.865 114.835 ;
        RECT 66.035 114.485 66.785 115.005 ;
        RECT 66.955 114.930 67.245 116.095 ;
        RECT 67.435 115.205 67.695 115.915 ;
        RECT 67.865 115.385 68.195 116.095 ;
        RECT 68.365 115.205 68.595 115.915 ;
        RECT 67.435 114.965 68.595 115.205 ;
        RECT 68.775 115.185 69.045 115.915 ;
        RECT 69.225 115.365 69.565 116.095 ;
        RECT 68.775 114.965 69.545 115.185 ;
        RECT 67.425 114.455 67.725 114.785 ;
        RECT 67.905 114.475 68.430 114.785 ;
        RECT 68.610 114.475 69.075 114.785 ;
        RECT 59.595 113.545 64.940 114.090 ;
        RECT 65.115 113.545 66.785 114.315 ;
        RECT 66.955 113.545 67.245 114.270 ;
        RECT 67.435 113.545 67.725 114.275 ;
        RECT 67.905 113.835 68.135 114.475 ;
        RECT 69.255 114.295 69.545 114.965 ;
        RECT 68.315 114.095 69.545 114.295 ;
        RECT 68.315 113.725 68.625 114.095 ;
        RECT 68.805 113.545 69.475 113.915 ;
        RECT 69.735 113.725 69.995 115.915 ;
        RECT 70.175 115.005 73.685 116.095 ;
        RECT 70.175 114.315 71.825 114.835 ;
        RECT 71.995 114.485 73.685 115.005 ;
        RECT 74.315 114.955 74.575 116.095 ;
        RECT 74.745 114.945 75.075 115.925 ;
        RECT 75.245 114.955 75.525 116.095 ;
        RECT 75.695 115.660 81.040 116.095 ;
        RECT 81.215 115.660 86.560 116.095 ;
        RECT 74.335 114.535 74.670 114.785 ;
        RECT 74.840 114.345 75.010 114.945 ;
        RECT 75.180 114.515 75.515 114.785 ;
        RECT 70.175 113.545 73.685 114.315 ;
        RECT 74.315 113.715 75.010 114.345 ;
        RECT 75.215 113.545 75.525 114.345 ;
        RECT 77.280 114.090 77.620 114.920 ;
        RECT 79.100 114.410 79.450 115.660 ;
        RECT 82.800 114.090 83.140 114.920 ;
        RECT 84.620 114.410 84.970 115.660 ;
        RECT 87.665 115.145 87.940 115.915 ;
        RECT 88.110 115.485 88.440 115.915 ;
        RECT 88.610 115.655 88.805 116.095 ;
        RECT 88.985 115.485 89.315 115.915 ;
        RECT 88.110 115.315 89.315 115.485 ;
        RECT 87.665 114.955 88.250 115.145 ;
        RECT 88.420 114.985 89.315 115.315 ;
        RECT 90.425 115.145 90.700 115.915 ;
        RECT 90.870 115.485 91.200 115.915 ;
        RECT 91.370 115.655 91.565 116.095 ;
        RECT 91.745 115.485 92.075 115.915 ;
        RECT 90.870 115.315 92.075 115.485 ;
        RECT 90.425 114.955 91.010 115.145 ;
        RECT 91.180 114.985 92.075 115.315 ;
        RECT 87.665 114.135 87.905 114.785 ;
        RECT 88.075 114.285 88.250 114.955 ;
        RECT 88.420 114.455 88.835 114.785 ;
        RECT 89.015 114.455 89.310 114.785 ;
        RECT 88.075 114.105 88.405 114.285 ;
        RECT 75.695 113.545 81.040 114.090 ;
        RECT 81.215 113.545 86.560 114.090 ;
        RECT 87.680 113.545 88.010 113.935 ;
        RECT 88.180 113.725 88.405 114.105 ;
        RECT 88.605 113.835 88.835 114.455 ;
        RECT 89.015 113.545 89.315 114.275 ;
        RECT 90.425 114.135 90.665 114.785 ;
        RECT 90.835 114.285 91.010 114.955 ;
        RECT 92.715 114.930 93.005 116.095 ;
        RECT 93.635 115.020 93.905 115.925 ;
        RECT 94.075 115.335 94.405 116.095 ;
        RECT 94.585 115.165 94.765 115.925 ;
        RECT 91.180 114.455 91.595 114.785 ;
        RECT 91.775 114.455 92.070 114.785 ;
        RECT 90.835 114.105 91.165 114.285 ;
        RECT 90.440 113.545 90.770 113.935 ;
        RECT 90.940 113.725 91.165 114.105 ;
        RECT 91.365 113.835 91.595 114.455 ;
        RECT 91.775 113.545 92.075 114.275 ;
        RECT 92.715 113.545 93.005 114.270 ;
        RECT 93.635 114.220 93.815 115.020 ;
        RECT 94.090 114.995 94.765 115.165 ;
        RECT 94.090 114.850 94.260 114.995 ;
        RECT 95.055 114.955 95.285 116.095 ;
        RECT 95.455 114.945 95.785 115.925 ;
        RECT 95.955 114.955 96.165 116.095 ;
        RECT 96.395 114.955 96.675 116.095 ;
        RECT 96.845 114.945 97.175 115.925 ;
        RECT 97.345 114.955 97.605 116.095 ;
        RECT 97.775 115.245 98.035 115.925 ;
        RECT 98.205 115.315 98.455 116.095 ;
        RECT 98.705 115.545 98.955 115.925 ;
        RECT 99.125 115.715 99.480 116.095 ;
        RECT 100.485 115.705 100.820 115.925 ;
        RECT 100.085 115.545 100.315 115.585 ;
        RECT 98.705 115.345 100.315 115.545 ;
        RECT 98.705 115.335 99.540 115.345 ;
        RECT 100.130 115.255 100.315 115.345 ;
        RECT 93.985 114.520 94.260 114.850 ;
        RECT 94.090 114.265 94.260 114.520 ;
        RECT 94.485 114.445 94.825 114.815 ;
        RECT 95.035 114.535 95.365 114.785 ;
        RECT 93.635 113.715 93.895 114.220 ;
        RECT 94.090 114.095 94.755 114.265 ;
        RECT 94.075 113.545 94.405 113.925 ;
        RECT 94.585 113.715 94.755 114.095 ;
        RECT 95.055 113.545 95.285 114.365 ;
        RECT 95.535 114.345 95.785 114.945 ;
        RECT 96.405 114.515 96.740 114.785 ;
        RECT 95.455 113.715 95.785 114.345 ;
        RECT 95.955 113.545 96.165 114.365 ;
        RECT 96.910 114.345 97.080 114.945 ;
        RECT 97.250 114.535 97.585 114.785 ;
        RECT 96.395 113.545 96.705 114.345 ;
        RECT 96.910 113.715 97.605 114.345 ;
        RECT 97.775 114.045 97.945 115.245 ;
        RECT 99.645 115.145 99.975 115.175 ;
        RECT 98.175 115.085 99.975 115.145 ;
        RECT 100.565 115.085 100.820 115.705 ;
        RECT 98.115 114.975 100.820 115.085 ;
        RECT 98.115 114.940 98.315 114.975 ;
        RECT 98.115 114.365 98.285 114.940 ;
        RECT 99.645 114.915 100.820 114.975 ;
        RECT 101.455 115.020 101.725 115.925 ;
        RECT 101.895 115.335 102.225 116.095 ;
        RECT 102.405 115.165 102.585 115.925 ;
        RECT 98.515 114.500 98.925 114.805 ;
        RECT 99.095 114.535 99.425 114.745 ;
        RECT 98.115 114.245 98.385 114.365 ;
        RECT 98.115 114.200 98.960 114.245 ;
        RECT 98.205 114.075 98.960 114.200 ;
        RECT 99.215 114.135 99.425 114.535 ;
        RECT 99.670 114.535 100.145 114.745 ;
        RECT 100.335 114.535 100.825 114.735 ;
        RECT 99.670 114.135 99.890 114.535 ;
        RECT 97.775 113.715 98.035 114.045 ;
        RECT 98.790 113.925 98.960 114.075 ;
        RECT 98.205 113.545 98.535 113.905 ;
        RECT 98.790 113.715 100.090 113.925 ;
        RECT 100.365 113.545 100.820 114.310 ;
        RECT 101.455 114.220 101.635 115.020 ;
        RECT 101.910 114.995 102.585 115.165 ;
        RECT 101.910 114.850 102.080 114.995 ;
        RECT 102.845 114.955 103.175 116.095 ;
        RECT 103.705 115.125 104.035 115.910 ;
        RECT 103.355 114.955 104.035 115.125 ;
        RECT 104.255 114.955 104.485 116.095 ;
        RECT 101.805 114.520 102.080 114.850 ;
        RECT 101.910 114.265 102.080 114.520 ;
        RECT 102.305 114.445 102.645 114.815 ;
        RECT 102.835 114.535 103.185 114.785 ;
        RECT 103.355 114.355 103.525 114.955 ;
        RECT 104.655 114.945 104.985 115.925 ;
        RECT 105.155 114.955 105.365 116.095 ;
        RECT 105.700 115.295 105.955 116.095 ;
        RECT 106.125 115.125 106.455 115.925 ;
        RECT 106.625 115.295 106.795 116.095 ;
        RECT 106.965 115.125 107.295 115.925 ;
        RECT 105.595 114.955 107.295 115.125 ;
        RECT 107.465 114.955 107.725 116.095 ;
        RECT 108.100 115.655 108.430 116.095 ;
        RECT 108.600 115.485 108.835 115.925 ;
        RECT 109.020 115.715 109.350 116.095 ;
        RECT 109.560 115.485 109.905 115.925 ;
        RECT 107.895 115.245 109.905 115.485 ;
        RECT 103.695 114.535 104.045 114.785 ;
        RECT 104.235 114.535 104.565 114.785 ;
        RECT 101.455 113.715 101.715 114.220 ;
        RECT 101.910 114.095 102.575 114.265 ;
        RECT 101.895 113.545 102.225 113.925 ;
        RECT 102.405 113.715 102.575 114.095 ;
        RECT 102.845 113.545 103.115 114.355 ;
        RECT 103.285 113.715 103.615 114.355 ;
        RECT 103.785 113.545 104.025 114.355 ;
        RECT 104.255 113.545 104.485 114.365 ;
        RECT 104.735 114.345 104.985 114.945 ;
        RECT 105.595 114.365 105.875 114.955 ;
        RECT 106.045 114.535 106.795 114.785 ;
        RECT 106.965 114.535 107.725 114.785 ;
        RECT 104.655 113.715 104.985 114.345 ;
        RECT 105.155 113.545 105.365 114.365 ;
        RECT 105.595 114.115 106.455 114.365 ;
        RECT 107.895 114.345 108.125 115.245 ;
        RECT 110.080 115.075 110.425 115.830 ;
        RECT 110.595 115.255 110.925 116.095 ;
        RECT 111.135 115.255 111.465 116.095 ;
        RECT 111.635 115.075 111.980 115.830 ;
        RECT 112.155 115.485 112.500 115.925 ;
        RECT 112.710 115.715 113.040 116.095 ;
        RECT 113.225 115.485 113.460 115.925 ;
        RECT 113.630 115.655 113.960 116.095 ;
        RECT 112.155 115.245 114.165 115.485 ;
        RECT 108.295 114.535 108.625 115.075 ;
        RECT 106.625 114.175 107.725 114.345 ;
        RECT 105.705 113.925 106.035 113.945 ;
        RECT 106.625 113.925 106.875 114.175 ;
        RECT 105.705 113.715 106.875 113.925 ;
        RECT 107.045 113.545 107.215 114.005 ;
        RECT 107.385 113.715 107.725 114.175 ;
        RECT 107.895 113.715 108.500 114.345 ;
        RECT 108.835 113.715 109.165 115.075 ;
        RECT 109.335 114.455 109.625 115.075 ;
        RECT 109.795 114.455 110.425 115.075 ;
        RECT 110.595 114.465 110.925 115.075 ;
        RECT 111.135 114.465 111.465 115.075 ;
        RECT 111.635 114.455 112.265 115.075 ;
        RECT 112.435 114.455 112.725 115.075 ;
        RECT 109.560 114.085 110.925 114.285 ;
        RECT 109.560 113.715 109.905 114.085 ;
        RECT 110.095 113.545 110.425 113.915 ;
        RECT 110.595 113.715 110.925 114.085 ;
        RECT 111.135 114.085 112.500 114.285 ;
        RECT 111.135 113.715 111.465 114.085 ;
        RECT 111.635 113.545 111.965 113.915 ;
        RECT 112.155 113.715 112.500 114.085 ;
        RECT 112.895 113.715 113.225 115.075 ;
        RECT 113.435 114.535 113.765 115.075 ;
        RECT 113.935 114.345 114.165 115.245 ;
        RECT 114.795 114.955 115.125 116.095 ;
        RECT 115.295 115.465 115.650 115.925 ;
        RECT 115.820 115.635 116.395 116.095 ;
        RECT 116.565 115.465 116.895 115.925 ;
        RECT 115.295 115.295 116.895 115.465 ;
        RECT 117.095 115.295 117.350 116.095 ;
        RECT 115.295 114.955 115.570 115.295 ;
        RECT 115.750 114.735 115.940 115.115 ;
        RECT 114.795 114.535 115.940 114.735 ;
        RECT 116.120 114.365 116.400 115.295 ;
        RECT 117.520 115.125 117.820 115.320 ;
        RECT 116.570 114.955 117.820 115.125 ;
        RECT 116.570 114.535 116.900 114.955 ;
        RECT 117.130 114.455 117.475 114.785 ;
        RECT 113.560 113.715 114.165 114.345 ;
        RECT 114.795 114.155 115.905 114.365 ;
        RECT 114.795 113.715 115.145 114.155 ;
        RECT 115.315 113.545 115.485 113.985 ;
        RECT 115.655 113.925 115.905 114.155 ;
        RECT 116.075 114.265 116.400 114.365 ;
        RECT 116.075 114.095 116.405 114.265 ;
        RECT 116.575 113.925 116.850 114.365 ;
        RECT 117.650 114.300 117.820 114.955 ;
        RECT 118.475 114.930 118.765 116.095 ;
        RECT 118.935 114.955 119.265 116.095 ;
        RECT 119.435 115.465 119.790 115.925 ;
        RECT 119.960 115.635 120.535 116.095 ;
        RECT 120.705 115.465 121.035 115.925 ;
        RECT 119.435 115.295 121.035 115.465 ;
        RECT 121.235 115.295 121.490 116.095 ;
        RECT 119.435 114.955 119.710 115.295 ;
        RECT 119.890 114.735 120.080 115.115 ;
        RECT 118.935 114.565 120.085 114.735 ;
        RECT 118.935 114.535 120.080 114.565 ;
        RECT 120.260 114.365 120.540 115.295 ;
        RECT 121.660 115.125 121.960 115.320 ;
        RECT 120.710 114.955 121.960 115.125 ;
        RECT 122.245 115.165 122.415 115.925 ;
        RECT 122.630 115.335 122.960 116.095 ;
        RECT 122.245 114.995 122.960 115.165 ;
        RECT 123.130 115.020 123.385 115.925 ;
        RECT 120.710 114.535 121.040 114.955 ;
        RECT 121.270 114.455 121.615 114.785 ;
        RECT 115.655 113.715 116.850 113.925 ;
        RECT 117.085 113.545 117.415 114.285 ;
        RECT 117.585 113.970 117.820 114.300 ;
        RECT 118.475 113.545 118.765 114.270 ;
        RECT 118.935 114.155 120.045 114.365 ;
        RECT 118.935 113.715 119.285 114.155 ;
        RECT 119.455 113.545 119.625 113.985 ;
        RECT 119.795 113.925 120.045 114.155 ;
        RECT 120.215 114.265 120.540 114.365 ;
        RECT 120.215 114.095 120.545 114.265 ;
        RECT 120.715 113.925 120.990 114.365 ;
        RECT 121.790 114.300 121.960 114.955 ;
        RECT 122.155 114.445 122.510 114.815 ;
        RECT 122.790 114.785 122.960 114.995 ;
        RECT 122.790 114.455 123.045 114.785 ;
        RECT 119.795 113.715 120.990 113.925 ;
        RECT 121.225 113.545 121.555 114.285 ;
        RECT 121.725 113.970 121.960 114.300 ;
        RECT 122.790 114.265 122.960 114.455 ;
        RECT 123.215 114.290 123.385 115.020 ;
        RECT 123.560 114.945 123.820 116.095 ;
        RECT 123.995 115.005 125.205 116.095 ;
        RECT 123.995 114.465 124.515 115.005 ;
        RECT 122.245 114.095 122.960 114.265 ;
        RECT 122.245 113.715 122.415 114.095 ;
        RECT 122.630 113.545 122.960 113.925 ;
        RECT 123.130 113.715 123.385 114.290 ;
        RECT 123.560 113.545 123.820 114.385 ;
        RECT 124.685 114.295 125.205 114.835 ;
        RECT 123.995 113.545 125.205 114.295 ;
        RECT 53.990 113.375 125.290 113.545 ;
        RECT 54.075 112.625 55.285 113.375 ;
        RECT 54.075 112.085 54.595 112.625 ;
        RECT 55.455 112.605 57.125 113.375 ;
        RECT 57.760 112.635 58.015 113.205 ;
        RECT 58.185 112.975 58.515 113.375 ;
        RECT 58.940 112.840 59.470 113.205 ;
        RECT 59.660 113.035 59.935 113.205 ;
        RECT 59.655 112.865 59.935 113.035 ;
        RECT 58.940 112.805 59.115 112.840 ;
        RECT 58.185 112.635 59.115 112.805 ;
        RECT 54.765 111.915 55.285 112.455 ;
        RECT 55.455 112.085 56.205 112.605 ;
        RECT 56.375 111.915 57.125 112.435 ;
        RECT 54.075 110.825 55.285 111.915 ;
        RECT 55.455 110.825 57.125 111.915 ;
        RECT 57.760 111.965 57.930 112.635 ;
        RECT 58.185 112.465 58.355 112.635 ;
        RECT 58.100 112.135 58.355 112.465 ;
        RECT 58.580 112.135 58.775 112.465 ;
        RECT 57.760 110.995 58.095 111.965 ;
        RECT 58.265 110.825 58.435 111.965 ;
        RECT 58.605 111.165 58.775 112.135 ;
        RECT 58.945 111.505 59.115 112.635 ;
        RECT 59.285 111.845 59.455 112.645 ;
        RECT 59.660 112.045 59.935 112.865 ;
        RECT 60.105 111.845 60.295 113.205 ;
        RECT 60.475 112.840 60.985 113.375 ;
        RECT 61.205 112.565 61.450 113.170 ;
        RECT 61.895 112.605 64.485 113.375 ;
        RECT 64.665 112.645 64.965 113.375 ;
        RECT 60.495 112.395 61.725 112.565 ;
        RECT 59.285 111.675 60.295 111.845 ;
        RECT 60.465 111.830 61.215 112.020 ;
        RECT 58.945 111.335 60.070 111.505 ;
        RECT 60.465 111.165 60.635 111.830 ;
        RECT 61.385 111.585 61.725 112.395 ;
        RECT 61.895 112.085 63.105 112.605 ;
        RECT 65.145 112.465 65.375 113.085 ;
        RECT 65.575 112.815 65.800 113.195 ;
        RECT 65.970 112.985 66.300 113.375 ;
        RECT 65.575 112.635 65.905 112.815 ;
        RECT 63.275 111.915 64.485 112.435 ;
        RECT 64.670 112.135 64.965 112.465 ;
        RECT 65.145 112.135 65.560 112.465 ;
        RECT 65.730 111.965 65.905 112.635 ;
        RECT 66.075 112.135 66.315 112.785 ;
        RECT 66.530 112.635 67.145 113.205 ;
        RECT 67.315 112.865 67.530 113.375 ;
        RECT 67.760 112.865 68.040 113.195 ;
        RECT 68.220 112.865 68.460 113.375 ;
        RECT 58.605 110.995 60.635 111.165 ;
        RECT 60.805 110.825 60.975 111.585 ;
        RECT 61.210 111.175 61.725 111.585 ;
        RECT 61.895 110.825 64.485 111.915 ;
        RECT 64.665 111.605 65.560 111.935 ;
        RECT 65.730 111.775 66.315 111.965 ;
        RECT 64.665 111.435 65.870 111.605 ;
        RECT 64.665 111.005 64.995 111.435 ;
        RECT 65.175 110.825 65.370 111.265 ;
        RECT 65.540 111.005 65.870 111.435 ;
        RECT 66.040 111.005 66.315 111.775 ;
        RECT 66.530 111.615 66.845 112.635 ;
        RECT 67.015 111.965 67.185 112.465 ;
        RECT 67.435 112.135 67.700 112.695 ;
        RECT 67.870 111.965 68.040 112.865 ;
        RECT 68.795 112.765 69.135 113.180 ;
        RECT 69.305 112.935 69.475 113.375 ;
        RECT 69.645 112.985 70.895 113.165 ;
        RECT 69.645 112.765 69.975 112.985 ;
        RECT 71.165 112.915 71.335 113.375 ;
        RECT 68.210 112.135 68.565 112.695 ;
        RECT 68.795 112.595 69.975 112.765 ;
        RECT 70.145 112.745 70.510 112.815 ;
        RECT 70.145 112.565 71.395 112.745 ;
        RECT 68.795 112.185 69.260 112.385 ;
        RECT 69.435 112.135 69.765 112.385 ;
        RECT 69.935 112.355 70.400 112.385 ;
        RECT 69.935 112.185 70.405 112.355 ;
        RECT 69.935 112.135 70.400 112.185 ;
        RECT 70.595 112.135 70.950 112.385 ;
        RECT 69.435 112.015 69.615 112.135 ;
        RECT 67.015 111.795 68.440 111.965 ;
        RECT 66.530 110.995 67.065 111.615 ;
        RECT 67.235 110.825 67.565 111.625 ;
        RECT 68.050 111.620 68.440 111.795 ;
        RECT 68.795 110.825 69.115 112.005 ;
        RECT 69.285 111.845 69.615 112.015 ;
        RECT 71.120 111.965 71.395 112.565 ;
        RECT 69.285 111.055 69.485 111.845 ;
        RECT 69.785 111.755 71.395 111.965 ;
        RECT 69.785 111.655 70.195 111.755 ;
        RECT 69.810 110.995 70.195 111.655 ;
        RECT 70.590 110.825 71.375 111.585 ;
        RECT 71.565 110.995 71.845 113.095 ;
        RECT 72.940 112.635 73.195 113.205 ;
        RECT 73.365 112.975 73.695 113.375 ;
        RECT 74.120 112.840 74.650 113.205 ;
        RECT 74.120 112.805 74.295 112.840 ;
        RECT 73.365 112.635 74.295 112.805 ;
        RECT 72.940 111.965 73.110 112.635 ;
        RECT 73.365 112.465 73.535 112.635 ;
        RECT 73.280 112.135 73.535 112.465 ;
        RECT 73.760 112.135 73.955 112.465 ;
        RECT 72.940 110.995 73.275 111.965 ;
        RECT 73.445 110.825 73.615 111.965 ;
        RECT 73.785 111.165 73.955 112.135 ;
        RECT 74.125 111.505 74.295 112.635 ;
        RECT 74.465 111.845 74.635 112.645 ;
        RECT 74.840 112.355 75.115 113.205 ;
        RECT 74.835 112.185 75.115 112.355 ;
        RECT 74.840 112.045 75.115 112.185 ;
        RECT 75.285 111.845 75.475 113.205 ;
        RECT 75.655 112.840 76.165 113.375 ;
        RECT 76.385 112.565 76.630 113.170 ;
        RECT 77.075 112.605 79.665 113.375 ;
        RECT 79.835 112.650 80.125 113.375 ;
        RECT 80.305 112.645 80.605 113.375 ;
        RECT 75.675 112.395 76.905 112.565 ;
        RECT 74.465 111.675 75.475 111.845 ;
        RECT 75.645 111.830 76.395 112.020 ;
        RECT 74.125 111.335 75.250 111.505 ;
        RECT 75.645 111.165 75.815 111.830 ;
        RECT 76.565 111.585 76.905 112.395 ;
        RECT 77.075 112.085 78.285 112.605 ;
        RECT 80.785 112.465 81.015 113.085 ;
        RECT 81.215 112.815 81.440 113.195 ;
        RECT 81.610 112.985 81.940 113.375 ;
        RECT 81.215 112.635 81.545 112.815 ;
        RECT 78.455 111.915 79.665 112.435 ;
        RECT 80.310 112.135 80.605 112.465 ;
        RECT 80.785 112.135 81.200 112.465 ;
        RECT 73.785 110.995 75.815 111.165 ;
        RECT 75.985 110.825 76.155 111.585 ;
        RECT 76.390 111.175 76.905 111.585 ;
        RECT 77.075 110.825 79.665 111.915 ;
        RECT 79.835 110.825 80.125 111.990 ;
        RECT 81.370 111.965 81.545 112.635 ;
        RECT 81.715 112.135 81.955 112.785 ;
        RECT 80.305 111.605 81.200 111.935 ;
        RECT 81.370 111.775 81.955 111.965 ;
        RECT 80.305 111.435 81.510 111.605 ;
        RECT 80.305 111.005 80.635 111.435 ;
        RECT 80.815 110.825 81.010 111.265 ;
        RECT 81.180 111.005 81.510 111.435 ;
        RECT 81.680 111.005 81.955 111.775 ;
        RECT 82.605 111.005 82.865 113.195 ;
        RECT 83.125 113.005 83.795 113.375 ;
        RECT 83.975 112.825 84.285 113.195 ;
        RECT 83.055 112.625 84.285 112.825 ;
        RECT 83.055 111.955 83.345 112.625 ;
        RECT 84.465 112.445 84.695 113.085 ;
        RECT 84.875 112.645 85.165 113.375 ;
        RECT 85.355 112.605 87.945 113.375 ;
        RECT 88.140 112.985 88.470 113.375 ;
        RECT 88.640 112.815 88.865 113.195 ;
        RECT 83.525 112.135 83.990 112.445 ;
        RECT 84.170 112.135 84.695 112.445 ;
        RECT 84.875 112.135 85.175 112.465 ;
        RECT 85.355 112.085 86.565 112.605 ;
        RECT 83.055 111.735 83.825 111.955 ;
        RECT 83.035 110.825 83.375 111.555 ;
        RECT 83.555 111.005 83.825 111.735 ;
        RECT 84.005 111.715 85.165 111.955 ;
        RECT 86.735 111.915 87.945 112.435 ;
        RECT 88.125 112.135 88.365 112.785 ;
        RECT 88.535 112.635 88.865 112.815 ;
        RECT 88.535 111.965 88.710 112.635 ;
        RECT 89.065 112.465 89.295 113.085 ;
        RECT 89.475 112.645 89.775 113.375 ;
        RECT 90.900 112.985 91.230 113.375 ;
        RECT 91.400 112.815 91.625 113.195 ;
        RECT 88.880 112.135 89.295 112.465 ;
        RECT 89.475 112.135 89.770 112.465 ;
        RECT 90.885 112.135 91.125 112.785 ;
        RECT 91.295 112.635 91.625 112.815 ;
        RECT 91.295 111.965 91.470 112.635 ;
        RECT 91.825 112.465 92.055 113.085 ;
        RECT 92.235 112.645 92.535 113.375 ;
        RECT 93.635 112.700 93.895 113.205 ;
        RECT 94.075 112.995 94.405 113.375 ;
        RECT 94.585 112.825 94.755 113.205 ;
        RECT 91.640 112.135 92.055 112.465 ;
        RECT 92.235 112.135 92.530 112.465 ;
        RECT 84.005 111.005 84.235 111.715 ;
        RECT 84.405 110.825 84.735 111.535 ;
        RECT 84.905 111.005 85.165 111.715 ;
        RECT 85.355 110.825 87.945 111.915 ;
        RECT 88.125 111.775 88.710 111.965 ;
        RECT 88.125 111.005 88.400 111.775 ;
        RECT 88.880 111.605 89.775 111.935 ;
        RECT 88.570 111.435 89.775 111.605 ;
        RECT 88.570 111.005 88.900 111.435 ;
        RECT 89.070 110.825 89.265 111.265 ;
        RECT 89.445 111.005 89.775 111.435 ;
        RECT 90.885 111.775 91.470 111.965 ;
        RECT 90.885 111.005 91.160 111.775 ;
        RECT 91.640 111.605 92.535 111.935 ;
        RECT 91.330 111.435 92.535 111.605 ;
        RECT 91.330 111.005 91.660 111.435 ;
        RECT 91.830 110.825 92.025 111.265 ;
        RECT 92.205 111.005 92.535 111.435 ;
        RECT 93.635 111.900 93.815 112.700 ;
        RECT 94.090 112.655 94.755 112.825 ;
        RECT 94.090 112.400 94.260 112.655 ;
        RECT 93.985 112.070 94.260 112.400 ;
        RECT 94.485 112.105 94.825 112.475 ;
        RECT 94.090 111.925 94.260 112.070 ;
        RECT 93.635 110.995 93.905 111.900 ;
        RECT 94.090 111.755 94.765 111.925 ;
        RECT 94.075 110.825 94.405 111.585 ;
        RECT 94.585 110.995 94.765 111.755 ;
        RECT 95.030 111.005 95.310 113.195 ;
        RECT 95.510 113.005 96.240 113.375 ;
        RECT 96.820 112.835 97.250 113.195 ;
        RECT 95.510 112.645 97.250 112.835 ;
        RECT 95.510 112.135 95.770 112.645 ;
        RECT 95.500 110.825 95.785 111.965 ;
        RECT 95.980 111.845 96.240 112.465 ;
        RECT 96.435 111.845 96.860 112.465 ;
        RECT 97.030 112.415 97.250 112.645 ;
        RECT 97.420 112.595 97.665 113.375 ;
        RECT 97.030 112.115 97.575 112.415 ;
        RECT 97.865 112.295 98.095 113.195 ;
        RECT 96.050 111.475 97.075 111.675 ;
        RECT 96.050 111.005 96.220 111.475 ;
        RECT 96.395 110.825 96.725 111.305 ;
        RECT 96.895 111.005 97.075 111.475 ;
        RECT 97.245 111.005 97.575 112.115 ;
        RECT 97.755 111.615 98.095 112.295 ;
        RECT 98.275 111.795 98.505 113.135 ;
        RECT 98.785 112.825 98.955 113.205 ;
        RECT 99.135 112.995 99.465 113.375 ;
        RECT 98.785 112.655 99.450 112.825 ;
        RECT 99.645 112.700 99.905 113.205 ;
        RECT 98.715 112.105 99.045 112.475 ;
        RECT 99.280 112.400 99.450 112.655 ;
        RECT 99.280 112.070 99.565 112.400 ;
        RECT 99.280 111.925 99.450 112.070 ;
        RECT 98.785 111.755 99.450 111.925 ;
        RECT 99.735 111.900 99.905 112.700 ;
        RECT 97.755 111.415 98.505 111.615 ;
        RECT 97.745 110.825 98.095 111.235 ;
        RECT 98.265 111.025 98.505 111.415 ;
        RECT 98.785 110.995 98.955 111.755 ;
        RECT 99.135 110.825 99.465 111.585 ;
        RECT 99.635 110.995 99.905 111.900 ;
        RECT 100.075 112.700 100.335 113.205 ;
        RECT 100.515 112.995 100.845 113.375 ;
        RECT 101.025 112.825 101.195 113.205 ;
        RECT 100.075 111.900 100.245 112.700 ;
        RECT 100.530 112.655 101.195 112.825 ;
        RECT 101.545 112.825 101.715 113.205 ;
        RECT 101.895 112.995 102.225 113.375 ;
        RECT 101.545 112.655 102.210 112.825 ;
        RECT 102.405 112.700 102.665 113.205 ;
        RECT 100.530 112.400 100.700 112.655 ;
        RECT 100.415 112.070 100.700 112.400 ;
        RECT 100.935 112.105 101.265 112.475 ;
        RECT 101.475 112.105 101.815 112.475 ;
        RECT 102.040 112.400 102.210 112.655 ;
        RECT 100.530 111.925 100.700 112.070 ;
        RECT 102.040 112.070 102.315 112.400 ;
        RECT 102.040 111.925 102.210 112.070 ;
        RECT 100.075 110.995 100.345 111.900 ;
        RECT 100.530 111.755 101.195 111.925 ;
        RECT 100.515 110.825 100.845 111.585 ;
        RECT 101.025 110.995 101.195 111.755 ;
        RECT 101.535 111.755 102.210 111.925 ;
        RECT 102.485 111.900 102.665 112.700 ;
        RECT 101.535 110.995 101.715 111.755 ;
        RECT 101.895 110.825 102.225 111.585 ;
        RECT 102.395 110.995 102.665 111.900 ;
        RECT 102.835 112.700 103.095 113.205 ;
        RECT 103.275 112.995 103.605 113.375 ;
        RECT 103.785 112.825 103.955 113.205 ;
        RECT 102.835 111.900 103.015 112.700 ;
        RECT 103.290 112.655 103.955 112.825 ;
        RECT 104.305 112.825 104.475 113.205 ;
        RECT 104.655 112.995 104.985 113.375 ;
        RECT 104.305 112.655 104.970 112.825 ;
        RECT 105.165 112.700 105.425 113.205 ;
        RECT 103.290 112.400 103.460 112.655 ;
        RECT 103.185 112.070 103.460 112.400 ;
        RECT 103.685 112.105 104.025 112.475 ;
        RECT 104.235 112.105 104.565 112.475 ;
        RECT 104.800 112.400 104.970 112.655 ;
        RECT 103.290 111.925 103.460 112.070 ;
        RECT 104.800 112.070 105.085 112.400 ;
        RECT 104.800 111.925 104.970 112.070 ;
        RECT 102.835 110.995 103.105 111.900 ;
        RECT 103.290 111.755 103.965 111.925 ;
        RECT 103.275 110.825 103.605 111.585 ;
        RECT 103.785 110.995 103.965 111.755 ;
        RECT 104.305 111.755 104.970 111.925 ;
        RECT 105.255 111.900 105.425 112.700 ;
        RECT 105.595 112.650 105.885 113.375 ;
        RECT 106.605 112.825 106.775 113.205 ;
        RECT 106.955 112.995 107.285 113.375 ;
        RECT 106.605 112.655 107.270 112.825 ;
        RECT 107.465 112.700 107.725 113.205 ;
        RECT 106.535 112.105 106.875 112.475 ;
        RECT 107.100 112.400 107.270 112.655 ;
        RECT 107.100 112.070 107.375 112.400 ;
        RECT 104.305 110.995 104.475 111.755 ;
        RECT 104.655 110.825 104.985 111.585 ;
        RECT 105.155 110.995 105.425 111.900 ;
        RECT 105.595 110.825 105.885 111.990 ;
        RECT 107.100 111.925 107.270 112.070 ;
        RECT 106.595 111.755 107.270 111.925 ;
        RECT 107.545 111.900 107.725 112.700 ;
        RECT 107.955 112.555 108.165 113.375 ;
        RECT 108.335 112.575 108.665 113.205 ;
        RECT 108.335 111.975 108.585 112.575 ;
        RECT 108.835 112.555 109.065 113.375 ;
        RECT 109.430 112.725 109.760 113.190 ;
        RECT 109.930 112.905 110.100 113.375 ;
        RECT 110.270 112.725 110.600 113.205 ;
        RECT 109.430 112.555 110.600 112.725 ;
        RECT 108.755 112.135 109.085 112.385 ;
        RECT 109.275 112.175 109.920 112.385 ;
        RECT 110.090 112.175 110.660 112.385 ;
        RECT 110.830 112.005 111.000 113.205 ;
        RECT 111.540 112.805 111.710 113.010 ;
        RECT 106.595 110.995 106.775 111.755 ;
        RECT 106.955 110.825 107.285 111.585 ;
        RECT 107.455 110.995 107.725 111.900 ;
        RECT 107.955 110.825 108.165 111.965 ;
        RECT 108.335 110.995 108.665 111.975 ;
        RECT 108.835 110.825 109.065 111.965 ;
        RECT 109.490 110.825 109.820 111.925 ;
        RECT 110.295 111.595 111.000 112.005 ;
        RECT 111.170 112.635 111.710 112.805 ;
        RECT 111.990 112.635 112.160 113.375 ;
        RECT 112.425 112.635 112.785 113.010 ;
        RECT 113.045 112.825 113.215 113.205 ;
        RECT 113.430 112.995 113.760 113.375 ;
        RECT 113.045 112.655 113.760 112.825 ;
        RECT 111.170 111.935 111.340 112.635 ;
        RECT 111.510 112.135 111.840 112.465 ;
        RECT 112.010 112.135 112.360 112.465 ;
        RECT 111.170 111.765 111.795 111.935 ;
        RECT 112.010 111.595 112.275 112.135 ;
        RECT 112.530 111.980 112.785 112.635 ;
        RECT 112.955 112.105 113.310 112.475 ;
        RECT 113.590 112.465 113.760 112.655 ;
        RECT 113.930 112.630 114.185 113.205 ;
        RECT 113.590 112.135 113.845 112.465 ;
        RECT 110.295 111.425 112.275 111.595 ;
        RECT 110.295 110.995 110.620 111.425 ;
        RECT 110.790 110.825 111.120 111.245 ;
        RECT 111.865 110.825 112.275 111.255 ;
        RECT 112.445 110.995 112.785 111.980 ;
        RECT 113.590 111.925 113.760 112.135 ;
        RECT 113.045 111.755 113.760 111.925 ;
        RECT 114.015 111.900 114.185 112.630 ;
        RECT 114.360 112.535 114.620 113.375 ;
        RECT 114.795 112.865 115.100 113.375 ;
        RECT 114.795 112.135 115.110 112.695 ;
        RECT 115.280 112.385 115.530 113.195 ;
        RECT 115.700 112.850 115.960 113.375 ;
        RECT 116.140 112.385 116.390 113.195 ;
        RECT 116.560 112.815 116.820 113.375 ;
        RECT 116.990 112.725 117.250 113.180 ;
        RECT 117.420 112.895 117.680 113.375 ;
        RECT 117.850 112.725 118.110 113.180 ;
        RECT 118.280 112.895 118.540 113.375 ;
        RECT 118.710 112.725 118.970 113.180 ;
        RECT 119.140 112.895 119.385 113.375 ;
        RECT 119.555 112.725 119.830 113.180 ;
        RECT 120.000 112.895 120.245 113.375 ;
        RECT 120.415 112.725 120.675 113.180 ;
        RECT 120.855 112.895 121.105 113.375 ;
        RECT 121.275 112.725 121.535 113.180 ;
        RECT 121.715 112.895 121.965 113.375 ;
        RECT 122.135 112.725 122.395 113.180 ;
        RECT 122.575 112.895 122.835 113.375 ;
        RECT 123.005 112.725 123.265 113.180 ;
        RECT 123.435 112.895 123.735 113.375 ;
        RECT 116.990 112.555 123.735 112.725 ;
        RECT 123.995 112.625 125.205 113.375 ;
        RECT 115.280 112.135 122.400 112.385 ;
        RECT 113.045 110.995 113.215 111.755 ;
        RECT 113.430 110.825 113.760 111.585 ;
        RECT 113.930 110.995 114.185 111.900 ;
        RECT 114.360 110.825 114.620 111.975 ;
        RECT 114.805 110.825 115.100 111.635 ;
        RECT 115.280 110.995 115.525 112.135 ;
        RECT 115.700 110.825 115.960 111.635 ;
        RECT 116.140 111.000 116.390 112.135 ;
        RECT 122.570 111.965 123.735 112.555 ;
        RECT 116.990 111.740 123.735 111.965 ;
        RECT 123.995 111.915 124.515 112.455 ;
        RECT 124.685 112.085 125.205 112.625 ;
        RECT 116.990 111.725 122.395 111.740 ;
        RECT 116.560 110.830 116.820 111.625 ;
        RECT 116.990 111.000 117.250 111.725 ;
        RECT 117.420 110.830 117.680 111.555 ;
        RECT 117.850 111.000 118.110 111.725 ;
        RECT 118.280 110.830 118.540 111.555 ;
        RECT 118.710 111.000 118.970 111.725 ;
        RECT 119.140 110.830 119.400 111.555 ;
        RECT 119.570 111.000 119.830 111.725 ;
        RECT 120.000 110.830 120.245 111.555 ;
        RECT 120.415 111.000 120.675 111.725 ;
        RECT 120.860 110.830 121.105 111.555 ;
        RECT 121.275 111.000 121.535 111.725 ;
        RECT 121.720 110.830 121.965 111.555 ;
        RECT 122.135 111.000 122.395 111.725 ;
        RECT 122.580 110.830 122.835 111.555 ;
        RECT 123.005 111.000 123.295 111.740 ;
        RECT 116.560 110.825 122.835 110.830 ;
        RECT 123.465 110.825 123.735 111.570 ;
        RECT 123.995 110.825 125.205 111.915 ;
        RECT 53.990 110.655 125.290 110.825 ;
        RECT 54.075 109.565 55.285 110.655 ;
        RECT 55.455 109.565 57.125 110.655 ;
        RECT 54.075 108.855 54.595 109.395 ;
        RECT 54.765 109.025 55.285 109.565 ;
        RECT 55.455 108.875 56.205 109.395 ;
        RECT 56.375 109.045 57.125 109.565 ;
        RECT 57.300 109.515 57.635 110.485 ;
        RECT 57.805 109.515 57.975 110.655 ;
        RECT 58.145 110.315 60.175 110.485 ;
        RECT 54.075 108.105 55.285 108.855 ;
        RECT 55.455 108.105 57.125 108.875 ;
        RECT 57.300 108.845 57.470 109.515 ;
        RECT 58.145 109.345 58.315 110.315 ;
        RECT 57.640 109.015 57.895 109.345 ;
        RECT 58.120 109.015 58.315 109.345 ;
        RECT 58.485 109.975 59.610 110.145 ;
        RECT 57.725 108.845 57.895 109.015 ;
        RECT 58.485 108.845 58.655 109.975 ;
        RECT 57.300 108.275 57.555 108.845 ;
        RECT 57.725 108.675 58.655 108.845 ;
        RECT 58.825 109.635 59.835 109.805 ;
        RECT 58.825 108.835 58.995 109.635 ;
        RECT 58.480 108.640 58.655 108.675 ;
        RECT 57.725 108.105 58.055 108.505 ;
        RECT 58.480 108.275 59.010 108.640 ;
        RECT 59.200 108.615 59.475 109.435 ;
        RECT 59.195 108.445 59.475 108.615 ;
        RECT 59.200 108.275 59.475 108.445 ;
        RECT 59.645 108.275 59.835 109.635 ;
        RECT 60.005 109.650 60.175 110.315 ;
        RECT 60.345 109.895 60.515 110.655 ;
        RECT 60.750 109.895 61.265 110.305 ;
        RECT 60.005 109.460 60.755 109.650 ;
        RECT 60.925 109.085 61.265 109.895 ;
        RECT 61.435 109.565 64.025 110.655 ;
        RECT 60.035 108.915 61.265 109.085 ;
        RECT 60.015 108.105 60.525 108.640 ;
        RECT 60.745 108.310 60.990 108.915 ;
        RECT 61.435 108.875 62.645 109.395 ;
        RECT 62.815 109.045 64.025 109.565 ;
        RECT 64.205 110.045 64.535 110.475 ;
        RECT 64.715 110.215 64.910 110.655 ;
        RECT 65.080 110.045 65.410 110.475 ;
        RECT 64.205 109.875 65.410 110.045 ;
        RECT 64.205 109.545 65.100 109.875 ;
        RECT 65.580 109.705 65.855 110.475 ;
        RECT 65.270 109.515 65.855 109.705 ;
        RECT 64.210 109.015 64.505 109.345 ;
        RECT 64.685 109.015 65.100 109.345 ;
        RECT 61.435 108.105 64.025 108.875 ;
        RECT 64.205 108.105 64.505 108.835 ;
        RECT 64.685 108.395 64.915 109.015 ;
        RECT 65.270 108.845 65.445 109.515 ;
        RECT 66.955 109.490 67.245 110.655 ;
        RECT 67.450 109.865 67.985 110.485 ;
        RECT 65.115 108.665 65.445 108.845 ;
        RECT 65.615 108.695 65.855 109.345 ;
        RECT 67.450 108.845 67.765 109.865 ;
        RECT 68.155 109.855 68.485 110.655 ;
        RECT 69.725 110.045 70.055 110.475 ;
        RECT 70.235 110.215 70.430 110.655 ;
        RECT 70.600 110.045 70.930 110.475 ;
        RECT 69.725 109.875 70.930 110.045 ;
        RECT 68.970 109.685 69.360 109.860 ;
        RECT 67.935 109.515 69.360 109.685 ;
        RECT 69.725 109.545 70.620 109.875 ;
        RECT 71.100 109.705 71.375 110.475 ;
        RECT 70.790 109.515 71.375 109.705 ;
        RECT 72.480 109.515 72.815 110.485 ;
        RECT 72.985 109.515 73.155 110.655 ;
        RECT 73.325 110.315 75.355 110.485 ;
        RECT 67.935 109.015 68.105 109.515 ;
        RECT 65.115 108.285 65.340 108.665 ;
        RECT 65.510 108.105 65.840 108.495 ;
        RECT 66.955 108.105 67.245 108.830 ;
        RECT 67.450 108.275 68.065 108.845 ;
        RECT 68.355 108.785 68.620 109.345 ;
        RECT 68.790 108.615 68.960 109.515 ;
        RECT 69.130 108.785 69.485 109.345 ;
        RECT 69.730 109.015 70.025 109.345 ;
        RECT 70.205 109.015 70.620 109.345 ;
        RECT 68.235 108.105 68.450 108.615 ;
        RECT 68.680 108.285 68.960 108.615 ;
        RECT 69.140 108.105 69.380 108.615 ;
        RECT 69.725 108.105 70.025 108.835 ;
        RECT 70.205 108.395 70.435 109.015 ;
        RECT 70.790 108.845 70.965 109.515 ;
        RECT 70.635 108.665 70.965 108.845 ;
        RECT 71.135 108.695 71.375 109.345 ;
        RECT 72.480 108.845 72.650 109.515 ;
        RECT 73.325 109.345 73.495 110.315 ;
        RECT 72.820 109.015 73.075 109.345 ;
        RECT 73.300 109.015 73.495 109.345 ;
        RECT 73.665 109.975 74.790 110.145 ;
        RECT 72.905 108.845 73.075 109.015 ;
        RECT 73.665 108.845 73.835 109.975 ;
        RECT 70.635 108.285 70.860 108.665 ;
        RECT 71.030 108.105 71.360 108.495 ;
        RECT 72.480 108.275 72.735 108.845 ;
        RECT 72.905 108.675 73.835 108.845 ;
        RECT 74.005 109.635 75.015 109.805 ;
        RECT 74.005 108.835 74.175 109.635 ;
        RECT 73.660 108.640 73.835 108.675 ;
        RECT 72.905 108.105 73.235 108.505 ;
        RECT 73.660 108.275 74.190 108.640 ;
        RECT 74.380 108.615 74.655 109.435 ;
        RECT 74.375 108.445 74.655 108.615 ;
        RECT 74.380 108.275 74.655 108.445 ;
        RECT 74.825 108.275 75.015 109.635 ;
        RECT 75.185 109.650 75.355 110.315 ;
        RECT 75.525 109.895 75.695 110.655 ;
        RECT 75.930 109.895 76.445 110.305 ;
        RECT 75.185 109.460 75.935 109.650 ;
        RECT 76.105 109.085 76.445 109.895 ;
        RECT 76.655 109.515 76.885 110.655 ;
        RECT 77.055 109.505 77.385 110.485 ;
        RECT 77.555 109.515 77.765 110.655 ;
        RECT 77.995 109.515 78.255 110.655 ;
        RECT 78.425 109.505 78.755 110.485 ;
        RECT 78.925 109.515 79.205 110.655 ;
        RECT 80.305 110.045 80.635 110.475 ;
        RECT 80.815 110.215 81.010 110.655 ;
        RECT 81.180 110.045 81.510 110.475 ;
        RECT 80.305 109.875 81.510 110.045 ;
        RECT 80.305 109.545 81.200 109.875 ;
        RECT 81.680 109.705 81.955 110.475 ;
        RECT 81.370 109.515 81.955 109.705 ;
        RECT 82.175 109.515 82.405 110.655 ;
        RECT 76.635 109.095 76.965 109.345 ;
        RECT 75.215 108.915 76.445 109.085 ;
        RECT 75.195 108.105 75.705 108.640 ;
        RECT 75.925 108.310 76.170 108.915 ;
        RECT 76.655 108.105 76.885 108.925 ;
        RECT 77.135 108.905 77.385 109.505 ;
        RECT 78.015 109.095 78.350 109.345 ;
        RECT 77.055 108.275 77.385 108.905 ;
        RECT 77.555 108.105 77.765 108.925 ;
        RECT 78.520 108.905 78.690 109.505 ;
        RECT 78.860 109.075 79.195 109.345 ;
        RECT 80.310 109.015 80.605 109.345 ;
        RECT 80.785 109.015 81.200 109.345 ;
        RECT 77.995 108.275 78.690 108.905 ;
        RECT 78.895 108.105 79.205 108.905 ;
        RECT 80.305 108.105 80.605 108.835 ;
        RECT 80.785 108.395 81.015 109.015 ;
        RECT 81.370 108.845 81.545 109.515 ;
        RECT 82.575 109.505 82.905 110.485 ;
        RECT 83.075 109.515 83.285 110.655 ;
        RECT 83.515 109.565 84.725 110.655 ;
        RECT 81.215 108.665 81.545 108.845 ;
        RECT 81.715 108.695 81.955 109.345 ;
        RECT 82.155 109.095 82.485 109.345 ;
        RECT 81.215 108.285 81.440 108.665 ;
        RECT 81.610 108.105 81.940 108.495 ;
        RECT 82.175 108.105 82.405 108.925 ;
        RECT 82.655 108.905 82.905 109.505 ;
        RECT 82.575 108.275 82.905 108.905 ;
        RECT 83.075 108.105 83.285 108.925 ;
        RECT 83.515 108.855 84.035 109.395 ;
        RECT 84.205 109.025 84.725 109.565 ;
        RECT 84.895 109.515 85.155 110.655 ;
        RECT 85.325 109.505 85.655 110.485 ;
        RECT 85.825 109.515 86.105 110.655 ;
        RECT 86.275 110.220 91.620 110.655 ;
        RECT 84.915 109.095 85.250 109.345 ;
        RECT 85.420 108.905 85.590 109.505 ;
        RECT 85.760 109.075 86.095 109.345 ;
        RECT 83.515 108.105 84.725 108.855 ;
        RECT 84.895 108.275 85.590 108.905 ;
        RECT 85.795 108.105 86.105 108.905 ;
        RECT 87.860 108.650 88.200 109.480 ;
        RECT 89.680 108.970 90.030 110.220 ;
        RECT 92.715 109.490 93.005 110.655 ;
        RECT 93.175 109.515 93.450 110.485 ;
        RECT 93.660 109.855 93.940 110.655 ;
        RECT 94.110 110.145 95.725 110.475 ;
        RECT 94.110 109.805 95.285 109.975 ;
        RECT 94.110 109.685 94.280 109.805 ;
        RECT 93.620 109.515 94.280 109.685 ;
        RECT 86.275 108.105 91.620 108.650 ;
        RECT 92.715 108.105 93.005 108.830 ;
        RECT 93.175 108.780 93.345 109.515 ;
        RECT 93.620 109.345 93.790 109.515 ;
        RECT 94.540 109.345 94.785 109.635 ;
        RECT 94.955 109.515 95.285 109.805 ;
        RECT 95.545 109.345 95.715 109.905 ;
        RECT 95.965 109.515 96.225 110.655 ;
        RECT 96.395 109.565 98.065 110.655 ;
        RECT 93.515 109.015 93.790 109.345 ;
        RECT 93.960 109.015 94.785 109.345 ;
        RECT 95.000 109.015 95.715 109.345 ;
        RECT 95.885 109.095 96.220 109.345 ;
        RECT 93.620 108.845 93.790 109.015 ;
        RECT 95.465 108.925 95.715 109.015 ;
        RECT 93.175 108.435 93.450 108.780 ;
        RECT 93.620 108.675 95.285 108.845 ;
        RECT 93.640 108.105 94.015 108.505 ;
        RECT 94.185 108.325 94.355 108.675 ;
        RECT 94.525 108.105 94.855 108.505 ;
        RECT 95.025 108.275 95.285 108.675 ;
        RECT 95.465 108.505 95.795 108.925 ;
        RECT 95.965 108.105 96.225 108.925 ;
        RECT 96.395 108.875 97.145 109.395 ;
        RECT 97.315 109.045 98.065 109.565 ;
        RECT 98.700 109.705 98.965 110.475 ;
        RECT 99.135 109.935 99.465 110.655 ;
        RECT 99.655 110.115 99.915 110.475 ;
        RECT 100.085 110.285 100.415 110.655 ;
        RECT 100.585 110.115 100.845 110.475 ;
        RECT 99.655 109.885 100.845 110.115 ;
        RECT 101.415 109.705 101.705 110.475 ;
        RECT 96.395 108.105 98.065 108.875 ;
        RECT 98.700 108.285 99.035 109.705 ;
        RECT 99.210 109.525 101.705 109.705 ;
        RECT 101.935 109.815 102.190 110.485 ;
        RECT 102.360 109.895 102.690 110.655 ;
        RECT 102.860 110.055 103.110 110.485 ;
        RECT 103.280 110.235 103.635 110.655 ;
        RECT 103.825 110.315 104.995 110.485 ;
        RECT 103.825 110.275 104.155 110.315 ;
        RECT 104.265 110.055 104.495 110.145 ;
        RECT 102.860 109.815 104.495 110.055 ;
        RECT 104.665 109.815 104.995 110.315 ;
        RECT 101.935 109.805 102.145 109.815 ;
        RECT 99.210 108.835 99.435 109.525 ;
        RECT 99.635 109.015 99.915 109.345 ;
        RECT 100.095 109.015 100.670 109.345 ;
        RECT 100.850 109.015 101.285 109.345 ;
        RECT 101.465 109.015 101.735 109.345 ;
        RECT 99.210 108.645 101.695 108.835 ;
        RECT 99.215 108.105 99.960 108.475 ;
        RECT 100.525 108.285 100.780 108.645 ;
        RECT 100.960 108.105 101.290 108.475 ;
        RECT 101.470 108.285 101.695 108.645 ;
        RECT 101.935 108.685 102.105 109.805 ;
        RECT 105.165 109.645 105.335 110.485 ;
        RECT 102.275 109.475 105.335 109.645 ;
        RECT 105.605 110.045 105.935 110.475 ;
        RECT 106.115 110.215 106.310 110.655 ;
        RECT 106.480 110.045 106.810 110.475 ;
        RECT 105.605 109.875 106.810 110.045 ;
        RECT 105.605 109.545 106.500 109.875 ;
        RECT 106.980 109.705 107.255 110.475 ;
        RECT 108.365 109.855 108.695 110.655 ;
        RECT 108.875 110.315 110.305 110.485 ;
        RECT 106.670 109.515 107.255 109.705 ;
        RECT 108.875 109.685 109.125 110.315 ;
        RECT 108.355 109.515 109.125 109.685 ;
        RECT 102.275 108.925 102.445 109.475 ;
        RECT 102.675 109.095 103.040 109.295 ;
        RECT 103.210 109.095 103.540 109.295 ;
        RECT 102.275 108.755 103.075 108.925 ;
        RECT 101.935 108.605 102.120 108.685 ;
        RECT 101.935 108.275 102.190 108.605 ;
        RECT 102.405 108.105 102.735 108.585 ;
        RECT 102.905 108.525 103.075 108.755 ;
        RECT 103.255 108.695 103.540 109.095 ;
        RECT 103.810 109.095 104.285 109.295 ;
        RECT 104.455 109.095 104.900 109.295 ;
        RECT 105.070 109.095 105.420 109.305 ;
        RECT 103.810 108.695 104.090 109.095 ;
        RECT 105.610 109.015 105.905 109.345 ;
        RECT 106.085 109.015 106.500 109.345 ;
        RECT 104.270 108.755 105.335 108.925 ;
        RECT 104.270 108.525 104.440 108.755 ;
        RECT 102.905 108.275 104.440 108.525 ;
        RECT 104.665 108.105 104.995 108.585 ;
        RECT 105.165 108.275 105.335 108.755 ;
        RECT 105.605 108.105 105.905 108.835 ;
        RECT 106.085 108.395 106.315 109.015 ;
        RECT 106.670 108.845 106.845 109.515 ;
        RECT 106.515 108.665 106.845 108.845 ;
        RECT 107.015 108.695 107.255 109.345 ;
        RECT 108.355 108.845 108.525 109.515 ;
        RECT 108.695 109.015 109.100 109.345 ;
        RECT 109.315 109.015 109.565 110.145 ;
        RECT 109.765 109.345 109.965 110.145 ;
        RECT 110.135 109.635 110.305 110.315 ;
        RECT 110.475 109.805 110.790 110.655 ;
        RECT 110.965 109.855 111.405 110.485 ;
        RECT 110.135 109.465 110.925 109.635 ;
        RECT 109.765 109.015 110.010 109.345 ;
        RECT 110.195 109.015 110.585 109.295 ;
        RECT 110.755 109.015 110.925 109.465 ;
        RECT 111.095 108.845 111.405 109.855 ;
        RECT 112.565 109.685 112.925 109.860 ;
        RECT 113.510 109.855 113.680 110.655 ;
        RECT 113.850 110.025 114.180 110.485 ;
        RECT 114.350 110.195 114.520 110.655 ;
        RECT 113.850 109.855 114.625 110.025 ;
        RECT 112.565 109.515 114.025 109.685 ;
        RECT 112.560 109.295 112.755 109.345 ;
        RECT 112.555 109.125 112.755 109.295 ;
        RECT 106.515 108.285 106.740 108.665 ;
        RECT 106.910 108.105 107.240 108.495 ;
        RECT 108.355 108.275 108.845 108.845 ;
        RECT 109.015 108.675 110.175 108.845 ;
        RECT 109.015 108.275 109.245 108.675 ;
        RECT 109.415 108.105 109.835 108.505 ;
        RECT 110.005 108.275 110.175 108.675 ;
        RECT 110.345 108.105 110.795 108.845 ;
        RECT 110.965 108.285 111.405 108.845 ;
        RECT 112.560 108.785 112.755 109.125 ;
        RECT 112.925 108.615 113.105 109.515 ;
        RECT 113.275 108.785 113.685 109.345 ;
        RECT 113.855 109.015 114.025 109.515 ;
        RECT 114.195 108.845 114.625 109.855 ;
        RECT 114.850 109.785 115.135 110.655 ;
        RECT 115.305 110.025 115.565 110.485 ;
        RECT 115.740 110.195 115.995 110.655 ;
        RECT 116.165 110.025 116.425 110.485 ;
        RECT 115.305 109.855 116.425 110.025 ;
        RECT 116.595 109.855 116.905 110.655 ;
        RECT 115.305 109.605 115.565 109.855 ;
        RECT 117.075 109.685 117.385 110.485 ;
        RECT 113.930 108.675 114.625 108.845 ;
        RECT 114.810 109.435 115.565 109.605 ;
        RECT 116.355 109.515 117.385 109.685 ;
        RECT 114.810 108.925 115.215 109.435 ;
        RECT 116.355 109.265 116.525 109.515 ;
        RECT 115.385 109.095 116.525 109.265 ;
        RECT 114.810 108.755 116.460 108.925 ;
        RECT 116.695 108.775 117.045 109.345 ;
        RECT 112.515 108.105 112.755 108.615 ;
        RECT 112.925 108.275 113.215 108.615 ;
        RECT 113.445 108.105 113.760 108.615 ;
        RECT 113.930 108.405 114.100 108.675 ;
        RECT 114.270 108.105 114.600 108.505 ;
        RECT 114.855 108.105 115.135 108.585 ;
        RECT 115.305 108.365 115.565 108.755 ;
        RECT 115.740 108.105 115.995 108.585 ;
        RECT 116.165 108.365 116.460 108.755 ;
        RECT 117.215 108.605 117.385 109.515 ;
        RECT 118.475 109.490 118.765 110.655 ;
        RECT 118.975 110.315 120.115 110.485 ;
        RECT 118.975 109.855 119.275 110.315 ;
        RECT 119.445 109.685 119.775 110.145 ;
        RECT 119.015 109.635 119.775 109.685 ;
        RECT 118.995 109.465 119.775 109.635 ;
        RECT 119.945 109.685 120.115 110.315 ;
        RECT 120.285 109.855 120.615 110.655 ;
        RECT 120.785 109.685 121.060 110.485 ;
        RECT 119.945 109.475 121.060 109.685 ;
        RECT 121.235 109.685 121.545 110.485 ;
        RECT 121.715 109.855 122.025 110.655 ;
        RECT 122.195 110.025 122.455 110.485 ;
        RECT 122.625 110.195 122.880 110.655 ;
        RECT 123.055 110.025 123.315 110.485 ;
        RECT 122.195 109.855 123.315 110.025 ;
        RECT 121.235 109.515 122.265 109.685 ;
        RECT 119.015 108.925 119.230 109.465 ;
        RECT 119.400 109.095 120.170 109.295 ;
        RECT 120.340 109.095 121.060 109.295 ;
        RECT 116.640 108.105 116.915 108.585 ;
        RECT 117.085 108.275 117.385 108.605 ;
        RECT 118.475 108.105 118.765 108.830 ;
        RECT 119.015 108.755 120.615 108.925 ;
        RECT 119.445 108.745 120.615 108.755 ;
        RECT 118.985 108.105 119.275 108.575 ;
        RECT 119.445 108.275 119.775 108.745 ;
        RECT 119.945 108.105 120.115 108.575 ;
        RECT 120.285 108.275 120.615 108.745 ;
        RECT 120.785 108.105 121.060 108.925 ;
        RECT 121.235 108.605 121.405 109.515 ;
        RECT 121.575 108.775 121.925 109.345 ;
        RECT 122.095 109.265 122.265 109.515 ;
        RECT 123.055 109.605 123.315 109.855 ;
        RECT 123.485 109.785 123.770 110.655 ;
        RECT 123.055 109.435 123.810 109.605 ;
        RECT 122.095 109.095 123.235 109.265 ;
        RECT 123.405 108.925 123.810 109.435 ;
        RECT 123.995 109.565 125.205 110.655 ;
        RECT 123.995 109.025 124.515 109.565 ;
        RECT 122.160 108.755 123.810 108.925 ;
        RECT 124.685 108.855 125.205 109.395 ;
        RECT 121.235 108.275 121.535 108.605 ;
        RECT 121.705 108.105 121.980 108.585 ;
        RECT 122.160 108.365 122.455 108.755 ;
        RECT 122.625 108.105 122.880 108.585 ;
        RECT 123.055 108.365 123.315 108.755 ;
        RECT 123.485 108.105 123.765 108.585 ;
        RECT 123.995 108.105 125.205 108.855 ;
        RECT 53.990 107.935 125.290 108.105 ;
        RECT 54.075 107.185 55.285 107.935 ;
        RECT 54.075 106.645 54.595 107.185 ;
        RECT 55.455 107.165 58.045 107.935 ;
        RECT 54.765 106.475 55.285 107.015 ;
        RECT 55.455 106.645 56.665 107.165 ;
        RECT 58.490 107.125 58.735 107.730 ;
        RECT 58.955 107.400 59.465 107.935 ;
        RECT 56.835 106.475 58.045 106.995 ;
        RECT 54.075 105.385 55.285 106.475 ;
        RECT 55.455 105.385 58.045 106.475 ;
        RECT 58.215 106.955 59.445 107.125 ;
        RECT 58.215 106.145 58.555 106.955 ;
        RECT 58.725 106.390 59.475 106.580 ;
        RECT 58.215 105.735 58.730 106.145 ;
        RECT 58.965 105.385 59.135 106.145 ;
        RECT 59.305 105.725 59.475 106.390 ;
        RECT 59.645 106.405 59.835 107.765 ;
        RECT 60.005 106.915 60.280 107.765 ;
        RECT 60.470 107.400 61.000 107.765 ;
        RECT 61.425 107.535 61.755 107.935 ;
        RECT 60.825 107.365 61.000 107.400 ;
        RECT 60.005 106.745 60.285 106.915 ;
        RECT 60.005 106.605 60.280 106.745 ;
        RECT 60.485 106.405 60.655 107.205 ;
        RECT 59.645 106.235 60.655 106.405 ;
        RECT 60.825 107.195 61.755 107.365 ;
        RECT 61.925 107.195 62.180 107.765 ;
        RECT 60.825 106.065 60.995 107.195 ;
        RECT 61.585 107.025 61.755 107.195 ;
        RECT 59.870 105.895 60.995 106.065 ;
        RECT 61.165 106.695 61.360 107.025 ;
        RECT 61.585 106.695 61.840 107.025 ;
        RECT 61.165 105.725 61.335 106.695 ;
        RECT 62.010 106.525 62.180 107.195 ;
        RECT 62.355 107.325 62.695 107.740 ;
        RECT 62.865 107.495 63.035 107.935 ;
        RECT 63.205 107.545 64.455 107.725 ;
        RECT 63.205 107.325 63.535 107.545 ;
        RECT 64.725 107.475 64.895 107.935 ;
        RECT 62.355 107.155 63.535 107.325 ;
        RECT 63.705 107.305 64.070 107.375 ;
        RECT 63.705 107.125 64.955 107.305 ;
        RECT 62.355 106.745 62.820 106.945 ;
        RECT 62.995 106.695 63.325 106.945 ;
        RECT 63.495 106.915 63.960 106.945 ;
        RECT 63.495 106.745 63.965 106.915 ;
        RECT 63.495 106.695 63.960 106.745 ;
        RECT 64.155 106.695 64.510 106.945 ;
        RECT 62.995 106.575 63.175 106.695 ;
        RECT 59.305 105.555 61.335 105.725 ;
        RECT 61.505 105.385 61.675 106.525 ;
        RECT 61.845 105.555 62.180 106.525 ;
        RECT 62.355 105.385 62.675 106.565 ;
        RECT 62.845 106.405 63.175 106.575 ;
        RECT 64.680 106.525 64.955 107.125 ;
        RECT 62.845 105.615 63.045 106.405 ;
        RECT 63.345 106.315 64.955 106.525 ;
        RECT 63.345 106.215 63.755 106.315 ;
        RECT 63.370 105.555 63.755 106.215 ;
        RECT 64.150 105.385 64.935 106.145 ;
        RECT 65.125 105.555 65.405 107.655 ;
        RECT 65.575 107.390 70.920 107.935 ;
        RECT 71.095 107.390 76.440 107.935 ;
        RECT 67.160 106.560 67.500 107.390 ;
        RECT 68.980 105.820 69.330 107.070 ;
        RECT 72.680 106.560 73.020 107.390 ;
        RECT 76.615 107.165 79.205 107.935 ;
        RECT 79.835 107.210 80.125 107.935 ;
        RECT 80.295 107.165 82.885 107.935 ;
        RECT 83.515 107.195 83.855 107.765 ;
        RECT 84.050 107.270 84.220 107.935 ;
        RECT 84.500 107.595 84.720 107.640 ;
        RECT 84.495 107.425 84.720 107.595 ;
        RECT 84.890 107.455 85.335 107.625 ;
        RECT 84.500 107.285 84.720 107.425 ;
        RECT 74.500 105.820 74.850 107.070 ;
        RECT 76.615 106.645 77.825 107.165 ;
        RECT 77.995 106.475 79.205 106.995 ;
        RECT 80.295 106.645 81.505 107.165 ;
        RECT 65.575 105.385 70.920 105.820 ;
        RECT 71.095 105.385 76.440 105.820 ;
        RECT 76.615 105.385 79.205 106.475 ;
        RECT 79.835 105.385 80.125 106.550 ;
        RECT 81.675 106.475 82.885 106.995 ;
        RECT 80.295 105.385 82.885 106.475 ;
        RECT 83.515 106.225 83.690 107.195 ;
        RECT 84.500 107.115 84.995 107.285 ;
        RECT 83.860 106.575 84.030 107.025 ;
        RECT 84.200 106.745 84.650 106.945 ;
        RECT 84.820 106.920 84.995 107.115 ;
        RECT 85.165 106.665 85.335 107.455 ;
        RECT 85.505 107.330 85.755 107.700 ;
        RECT 85.585 106.945 85.755 107.330 ;
        RECT 85.925 107.295 86.175 107.700 ;
        RECT 86.345 107.465 86.515 107.935 ;
        RECT 86.685 107.295 87.025 107.700 ;
        RECT 85.925 107.115 87.025 107.295 ;
        RECT 87.195 107.165 88.865 107.935 ;
        RECT 89.045 107.210 89.375 107.720 ;
        RECT 89.545 107.535 89.875 107.935 ;
        RECT 90.925 107.365 91.255 107.705 ;
        RECT 91.425 107.535 91.755 107.935 ;
        RECT 85.585 106.775 85.780 106.945 ;
        RECT 83.860 106.405 84.255 106.575 ;
        RECT 85.165 106.525 85.440 106.665 ;
        RECT 83.515 105.555 83.775 106.225 ;
        RECT 84.085 106.135 84.255 106.405 ;
        RECT 84.425 106.305 85.440 106.525 ;
        RECT 85.610 106.525 85.780 106.775 ;
        RECT 85.950 106.695 86.510 106.945 ;
        RECT 85.610 106.135 86.165 106.525 ;
        RECT 84.085 105.965 86.165 106.135 ;
        RECT 83.945 105.385 84.275 105.785 ;
        RECT 85.145 105.385 85.545 105.785 ;
        RECT 85.835 105.730 86.165 105.965 ;
        RECT 86.335 105.595 86.510 106.695 ;
        RECT 86.680 106.375 87.025 106.945 ;
        RECT 87.195 106.645 87.945 107.165 ;
        RECT 88.115 106.475 88.865 106.995 ;
        RECT 86.680 105.385 87.025 106.205 ;
        RECT 87.195 105.385 88.865 106.475 ;
        RECT 89.045 106.445 89.235 107.210 ;
        RECT 89.545 107.195 91.910 107.365 ;
        RECT 89.545 107.025 89.715 107.195 ;
        RECT 89.405 106.695 89.715 107.025 ;
        RECT 89.885 106.695 90.190 107.025 ;
        RECT 89.045 105.595 89.375 106.445 ;
        RECT 89.545 105.385 89.795 106.525 ;
        RECT 89.975 106.365 90.190 106.695 ;
        RECT 90.365 106.365 90.650 107.025 ;
        RECT 90.845 106.365 91.110 107.025 ;
        RECT 91.325 106.365 91.570 107.025 ;
        RECT 91.740 106.195 91.910 107.195 ;
        RECT 92.460 107.155 92.960 107.765 ;
        RECT 92.255 106.695 92.605 106.945 ;
        RECT 92.790 106.525 92.960 107.155 ;
        RECT 93.590 107.285 93.920 107.765 ;
        RECT 94.090 107.475 94.315 107.935 ;
        RECT 94.485 107.285 94.815 107.765 ;
        RECT 93.590 107.115 94.815 107.285 ;
        RECT 95.005 107.135 95.255 107.935 ;
        RECT 95.425 107.135 95.765 107.765 ;
        RECT 96.100 107.425 96.340 107.935 ;
        RECT 96.520 107.425 96.800 107.755 ;
        RECT 97.030 107.425 97.245 107.935 ;
        RECT 93.130 106.745 93.460 106.945 ;
        RECT 93.630 106.745 93.960 106.945 ;
        RECT 94.130 106.745 94.550 106.945 ;
        RECT 94.725 106.775 95.420 106.945 ;
        RECT 94.725 106.525 94.895 106.775 ;
        RECT 95.590 106.525 95.765 107.135 ;
        RECT 95.995 106.695 96.350 107.255 ;
        RECT 96.520 106.525 96.690 107.425 ;
        RECT 96.860 106.695 97.125 107.255 ;
        RECT 97.415 107.195 98.030 107.765 ;
        RECT 97.375 106.525 97.545 107.025 ;
        RECT 89.985 106.025 91.275 106.195 ;
        RECT 89.985 105.605 90.235 106.025 ;
        RECT 90.465 105.385 90.795 105.855 ;
        RECT 91.025 105.605 91.275 106.025 ;
        RECT 91.455 106.025 91.910 106.195 ;
        RECT 92.460 106.355 94.895 106.525 ;
        RECT 91.455 105.595 91.785 106.025 ;
        RECT 92.460 105.555 92.790 106.355 ;
        RECT 92.960 105.385 93.290 106.185 ;
        RECT 93.590 105.555 93.920 106.355 ;
        RECT 94.565 105.385 94.815 106.185 ;
        RECT 95.085 105.385 95.255 106.525 ;
        RECT 95.425 105.555 95.765 106.525 ;
        RECT 96.120 106.355 97.545 106.525 ;
        RECT 96.120 106.180 96.510 106.355 ;
        RECT 96.995 105.385 97.325 106.185 ;
        RECT 97.715 106.175 98.030 107.195 ;
        RECT 98.235 107.135 98.930 107.765 ;
        RECT 99.135 107.135 99.445 107.935 ;
        RECT 99.615 107.165 102.205 107.935 ;
        RECT 102.400 107.545 102.730 107.935 ;
        RECT 102.900 107.375 103.125 107.755 ;
        RECT 98.255 106.695 98.590 106.945 ;
        RECT 98.760 106.575 98.930 107.135 ;
        RECT 99.100 106.695 99.435 106.965 ;
        RECT 99.615 106.645 100.825 107.165 ;
        RECT 98.755 106.535 98.930 106.575 ;
        RECT 97.495 105.555 98.030 106.175 ;
        RECT 98.235 105.385 98.495 106.525 ;
        RECT 98.665 105.555 98.995 106.535 ;
        RECT 99.165 105.385 99.445 106.525 ;
        RECT 100.995 106.475 102.205 106.995 ;
        RECT 102.385 106.695 102.625 107.345 ;
        RECT 102.795 107.195 103.125 107.375 ;
        RECT 102.795 106.525 102.970 107.195 ;
        RECT 103.325 107.025 103.555 107.645 ;
        RECT 103.735 107.205 104.035 107.935 ;
        RECT 104.305 107.385 104.475 107.765 ;
        RECT 104.655 107.555 104.985 107.935 ;
        RECT 104.305 107.215 104.970 107.385 ;
        RECT 105.165 107.260 105.425 107.765 ;
        RECT 103.140 106.695 103.555 107.025 ;
        RECT 103.735 106.695 104.030 107.025 ;
        RECT 104.235 106.665 104.575 107.035 ;
        RECT 104.800 106.960 104.970 107.215 ;
        RECT 99.615 105.385 102.205 106.475 ;
        RECT 102.385 106.335 102.970 106.525 ;
        RECT 104.800 106.630 105.075 106.960 ;
        RECT 102.385 105.565 102.660 106.335 ;
        RECT 103.140 106.165 104.035 106.495 ;
        RECT 104.800 106.485 104.970 106.630 ;
        RECT 102.830 105.995 104.035 106.165 ;
        RECT 102.830 105.565 103.160 105.995 ;
        RECT 103.330 105.385 103.525 105.825 ;
        RECT 103.705 105.565 104.035 105.995 ;
        RECT 104.295 106.315 104.970 106.485 ;
        RECT 105.245 106.460 105.425 107.260 ;
        RECT 105.595 107.210 105.885 107.935 ;
        RECT 107.065 107.385 107.235 107.765 ;
        RECT 107.415 107.555 107.745 107.935 ;
        RECT 107.065 107.215 107.730 107.385 ;
        RECT 107.925 107.260 108.185 107.765 ;
        RECT 106.995 106.665 107.325 107.035 ;
        RECT 107.560 106.960 107.730 107.215 ;
        RECT 107.560 106.630 107.845 106.960 ;
        RECT 104.295 105.555 104.475 106.315 ;
        RECT 104.655 105.385 104.985 106.145 ;
        RECT 105.155 105.555 105.425 106.460 ;
        RECT 105.595 105.385 105.885 106.550 ;
        RECT 107.560 106.485 107.730 106.630 ;
        RECT 107.065 106.315 107.730 106.485 ;
        RECT 108.015 106.460 108.185 107.260 ;
        RECT 108.445 107.385 108.615 107.765 ;
        RECT 108.795 107.555 109.125 107.935 ;
        RECT 108.445 107.215 109.110 107.385 ;
        RECT 109.305 107.260 109.565 107.765 ;
        RECT 108.375 106.665 108.705 107.035 ;
        RECT 108.940 106.960 109.110 107.215 ;
        RECT 108.940 106.630 109.225 106.960 ;
        RECT 108.940 106.485 109.110 106.630 ;
        RECT 107.065 105.555 107.235 106.315 ;
        RECT 107.415 105.385 107.745 106.145 ;
        RECT 107.915 105.555 108.185 106.460 ;
        RECT 108.445 106.315 109.110 106.485 ;
        RECT 109.395 106.460 109.565 107.260 ;
        RECT 108.445 105.555 108.615 106.315 ;
        RECT 108.795 105.385 109.125 106.145 ;
        RECT 109.295 105.555 109.565 106.460 ;
        RECT 109.735 107.195 110.095 107.570 ;
        RECT 110.360 107.195 110.530 107.935 ;
        RECT 110.810 107.365 110.980 107.570 ;
        RECT 110.810 107.195 111.350 107.365 ;
        RECT 109.735 106.540 109.990 107.195 ;
        RECT 110.160 106.695 110.510 107.025 ;
        RECT 110.680 106.695 111.010 107.025 ;
        RECT 109.735 105.555 110.075 106.540 ;
        RECT 110.245 106.155 110.510 106.695 ;
        RECT 111.180 106.495 111.350 107.195 ;
        RECT 110.725 106.325 111.350 106.495 ;
        RECT 111.520 106.565 111.690 107.765 ;
        RECT 111.920 107.285 112.250 107.765 ;
        RECT 112.420 107.465 112.590 107.935 ;
        RECT 112.760 107.285 113.090 107.750 ;
        RECT 111.920 107.115 113.090 107.285 ;
        RECT 113.430 107.365 113.685 107.715 ;
        RECT 113.855 107.535 114.185 107.935 ;
        RECT 114.355 107.365 114.525 107.715 ;
        RECT 114.695 107.535 115.075 107.935 ;
        RECT 113.430 107.195 115.095 107.365 ;
        RECT 115.265 107.260 115.540 107.605 ;
        RECT 116.640 107.430 116.975 107.935 ;
        RECT 117.145 107.365 117.385 107.740 ;
        RECT 117.665 107.605 117.835 107.750 ;
        RECT 117.665 107.410 118.040 107.605 ;
        RECT 118.400 107.440 118.795 107.935 ;
        RECT 114.925 107.025 115.095 107.195 ;
        RECT 111.860 106.735 112.430 106.945 ;
        RECT 112.600 106.735 113.245 106.945 ;
        RECT 113.415 106.695 113.760 107.025 ;
        RECT 113.930 106.695 114.755 107.025 ;
        RECT 114.925 106.695 115.200 107.025 ;
        RECT 111.520 106.155 112.225 106.565 ;
        RECT 110.245 105.985 112.225 106.155 ;
        RECT 110.245 105.385 110.655 105.815 ;
        RECT 111.400 105.385 111.730 105.805 ;
        RECT 111.900 105.555 112.225 105.985 ;
        RECT 112.700 105.385 113.030 106.485 ;
        RECT 113.435 106.235 113.760 106.525 ;
        RECT 113.930 106.405 114.125 106.695 ;
        RECT 114.925 106.525 115.095 106.695 ;
        RECT 115.370 106.525 115.540 107.260 ;
        RECT 114.435 106.355 115.095 106.525 ;
        RECT 114.435 106.235 114.605 106.355 ;
        RECT 113.435 106.065 114.605 106.235 ;
        RECT 113.415 105.605 114.605 105.895 ;
        RECT 114.775 105.385 115.055 106.185 ;
        RECT 115.265 105.555 115.540 106.525 ;
        RECT 116.695 106.405 116.995 107.255 ;
        RECT 117.165 107.215 117.385 107.365 ;
        RECT 117.165 106.885 117.700 107.215 ;
        RECT 117.870 107.075 118.040 107.410 ;
        RECT 118.965 107.245 119.205 107.765 ;
        RECT 119.395 107.275 119.670 107.935 ;
        RECT 119.840 107.305 120.090 107.765 ;
        RECT 120.265 107.440 120.595 107.935 ;
        RECT 117.165 106.235 117.400 106.885 ;
        RECT 117.870 106.715 118.855 107.075 ;
        RECT 116.725 106.005 117.400 106.235 ;
        RECT 117.570 106.695 118.855 106.715 ;
        RECT 117.570 106.545 118.430 106.695 ;
        RECT 116.725 105.575 116.895 106.005 ;
        RECT 117.065 105.385 117.395 105.835 ;
        RECT 117.570 105.600 117.855 106.545 ;
        RECT 119.030 106.440 119.205 107.245 ;
        RECT 119.840 107.095 120.010 107.305 ;
        RECT 120.775 107.270 121.005 107.715 ;
        RECT 119.395 106.575 120.010 107.095 ;
        RECT 120.180 106.595 120.410 107.025 ;
        RECT 120.595 106.775 121.005 107.270 ;
        RECT 121.175 107.450 121.965 107.715 ;
        RECT 121.175 106.595 121.430 107.450 ;
        RECT 122.245 107.385 122.415 107.765 ;
        RECT 122.630 107.555 122.960 107.935 ;
        RECT 121.600 106.775 121.985 107.255 ;
        RECT 122.245 107.215 122.960 107.385 ;
        RECT 122.155 106.665 122.510 107.035 ;
        RECT 122.790 107.025 122.960 107.215 ;
        RECT 123.130 107.190 123.385 107.765 ;
        RECT 122.790 106.695 123.045 107.025 ;
        RECT 118.030 106.065 118.725 106.375 ;
        RECT 118.035 105.385 118.720 105.855 ;
        RECT 118.900 105.655 119.205 106.440 ;
        RECT 119.395 105.385 119.655 106.395 ;
        RECT 119.825 106.225 119.995 106.575 ;
        RECT 120.180 106.425 121.970 106.595 ;
        RECT 122.790 106.485 122.960 106.695 ;
        RECT 119.825 105.555 120.100 106.225 ;
        RECT 120.300 105.385 120.515 106.230 ;
        RECT 120.740 106.130 120.990 106.425 ;
        RECT 121.215 106.065 121.545 106.255 ;
        RECT 120.700 105.555 121.175 105.895 ;
        RECT 121.355 105.890 121.545 106.065 ;
        RECT 121.715 106.060 121.970 106.425 ;
        RECT 122.245 106.315 122.960 106.485 ;
        RECT 123.215 106.460 123.385 107.190 ;
        RECT 123.560 107.095 123.820 107.935 ;
        RECT 123.995 107.185 125.205 107.935 ;
        RECT 121.355 105.385 121.985 105.890 ;
        RECT 122.245 105.555 122.415 106.315 ;
        RECT 122.630 105.385 122.960 106.145 ;
        RECT 123.130 105.555 123.385 106.460 ;
        RECT 123.560 105.385 123.820 106.535 ;
        RECT 123.995 106.475 124.515 107.015 ;
        RECT 124.685 106.645 125.205 107.185 ;
        RECT 123.995 105.385 125.205 106.475 ;
        RECT 53.990 105.215 125.290 105.385 ;
        RECT 54.075 104.125 55.285 105.215 ;
        RECT 55.455 104.125 58.045 105.215 ;
        RECT 54.075 103.415 54.595 103.955 ;
        RECT 54.765 103.585 55.285 104.125 ;
        RECT 55.455 103.435 56.665 103.955 ;
        RECT 56.835 103.605 58.045 104.125 ;
        RECT 58.215 104.455 58.730 104.865 ;
        RECT 58.965 104.455 59.135 105.215 ;
        RECT 59.305 104.875 61.335 105.045 ;
        RECT 58.215 103.645 58.555 104.455 ;
        RECT 59.305 104.210 59.475 104.875 ;
        RECT 59.870 104.535 60.995 104.705 ;
        RECT 58.725 104.020 59.475 104.210 ;
        RECT 59.645 104.195 60.655 104.365 ;
        RECT 58.215 103.475 59.445 103.645 ;
        RECT 54.075 102.665 55.285 103.415 ;
        RECT 55.455 102.665 58.045 103.435 ;
        RECT 58.490 102.870 58.735 103.475 ;
        RECT 58.955 102.665 59.465 103.200 ;
        RECT 59.645 102.835 59.835 104.195 ;
        RECT 60.005 103.855 60.280 103.995 ;
        RECT 60.005 103.685 60.285 103.855 ;
        RECT 60.005 102.835 60.280 103.685 ;
        RECT 60.485 103.395 60.655 104.195 ;
        RECT 60.825 103.405 60.995 104.535 ;
        RECT 61.165 103.905 61.335 104.875 ;
        RECT 61.505 104.075 61.675 105.215 ;
        RECT 61.845 104.075 62.180 105.045 ;
        RECT 62.355 104.125 64.945 105.215 ;
        RECT 61.165 103.575 61.360 103.905 ;
        RECT 61.585 103.575 61.840 103.905 ;
        RECT 61.585 103.405 61.755 103.575 ;
        RECT 62.010 103.405 62.180 104.075 ;
        RECT 60.825 103.235 61.755 103.405 ;
        RECT 60.825 103.200 61.000 103.235 ;
        RECT 60.470 102.835 61.000 103.200 ;
        RECT 61.425 102.665 61.755 103.065 ;
        RECT 61.925 102.835 62.180 103.405 ;
        RECT 62.355 103.435 63.565 103.955 ;
        RECT 63.735 103.605 64.945 104.125 ;
        RECT 65.575 104.075 65.835 105.215 ;
        RECT 66.005 104.065 66.335 105.045 ;
        RECT 66.505 104.075 66.785 105.215 ;
        RECT 65.595 103.655 65.930 103.905 ;
        RECT 66.100 103.465 66.270 104.065 ;
        RECT 66.955 104.050 67.245 105.215 ;
        RECT 67.415 104.035 67.735 105.215 ;
        RECT 67.905 104.195 68.105 104.985 ;
        RECT 68.430 104.385 68.815 105.045 ;
        RECT 69.210 104.455 69.995 105.215 ;
        RECT 68.405 104.285 68.815 104.385 ;
        RECT 67.905 104.025 68.235 104.195 ;
        RECT 68.405 104.075 70.015 104.285 ;
        RECT 68.055 103.905 68.235 104.025 ;
        RECT 66.440 103.635 66.775 103.905 ;
        RECT 67.415 103.655 67.880 103.855 ;
        RECT 68.055 103.655 68.385 103.905 ;
        RECT 68.555 103.855 69.020 103.905 ;
        RECT 68.555 103.685 69.025 103.855 ;
        RECT 68.555 103.655 69.020 103.685 ;
        RECT 69.215 103.655 69.570 103.905 ;
        RECT 69.740 103.475 70.015 104.075 ;
        RECT 62.355 102.665 64.945 103.435 ;
        RECT 65.575 102.835 66.270 103.465 ;
        RECT 66.475 102.665 66.785 103.465 ;
        RECT 66.955 102.665 67.245 103.390 ;
        RECT 67.415 103.275 68.595 103.445 ;
        RECT 67.415 102.860 67.755 103.275 ;
        RECT 67.925 102.665 68.095 103.105 ;
        RECT 68.265 103.055 68.595 103.275 ;
        RECT 68.765 103.295 70.015 103.475 ;
        RECT 68.765 103.225 69.130 103.295 ;
        RECT 68.265 102.875 69.515 103.055 ;
        RECT 69.785 102.665 69.955 103.125 ;
        RECT 70.185 102.945 70.465 105.045 ;
        RECT 71.100 104.075 71.435 105.045 ;
        RECT 71.605 104.075 71.775 105.215 ;
        RECT 71.945 104.875 73.975 105.045 ;
        RECT 71.100 103.405 71.270 104.075 ;
        RECT 71.945 103.905 72.115 104.875 ;
        RECT 71.440 103.575 71.695 103.905 ;
        RECT 71.920 103.575 72.115 103.905 ;
        RECT 72.285 104.535 73.410 104.705 ;
        RECT 71.525 103.405 71.695 103.575 ;
        RECT 72.285 103.405 72.455 104.535 ;
        RECT 71.100 102.835 71.355 103.405 ;
        RECT 71.525 103.235 72.455 103.405 ;
        RECT 72.625 104.195 73.635 104.365 ;
        RECT 72.625 103.395 72.795 104.195 ;
        RECT 72.280 103.200 72.455 103.235 ;
        RECT 71.525 102.665 71.855 103.065 ;
        RECT 72.280 102.835 72.810 103.200 ;
        RECT 73.000 103.175 73.275 103.995 ;
        RECT 72.995 103.005 73.275 103.175 ;
        RECT 73.000 102.835 73.275 103.005 ;
        RECT 73.445 102.835 73.635 104.195 ;
        RECT 73.805 104.210 73.975 104.875 ;
        RECT 74.145 104.455 74.315 105.215 ;
        RECT 74.550 104.455 75.065 104.865 ;
        RECT 73.805 104.020 74.555 104.210 ;
        RECT 74.725 103.645 75.065 104.455 ;
        RECT 75.235 104.075 75.495 105.215 ;
        RECT 75.665 104.065 75.995 105.045 ;
        RECT 76.165 104.075 76.445 105.215 ;
        RECT 76.615 104.125 79.205 105.215 ;
        RECT 75.255 103.655 75.590 103.905 ;
        RECT 73.835 103.475 75.065 103.645 ;
        RECT 73.815 102.665 74.325 103.200 ;
        RECT 74.545 102.870 74.790 103.475 ;
        RECT 75.760 103.465 75.930 104.065 ;
        RECT 76.100 103.635 76.435 103.905 ;
        RECT 75.235 102.835 75.930 103.465 ;
        RECT 76.135 102.665 76.445 103.465 ;
        RECT 76.615 103.435 77.825 103.955 ;
        RECT 77.995 103.605 79.205 104.125 ;
        RECT 79.380 104.265 79.645 105.035 ;
        RECT 79.815 104.495 80.145 105.215 ;
        RECT 80.335 104.675 80.595 105.035 ;
        RECT 80.765 104.845 81.095 105.215 ;
        RECT 81.265 104.675 81.525 105.035 ;
        RECT 80.335 104.445 81.525 104.675 ;
        RECT 82.095 104.265 82.385 105.035 ;
        RECT 82.595 104.780 87.940 105.215 ;
        RECT 76.615 102.665 79.205 103.435 ;
        RECT 79.380 102.845 79.715 104.265 ;
        RECT 79.890 104.085 82.385 104.265 ;
        RECT 79.890 103.395 80.115 104.085 ;
        RECT 80.315 103.575 80.595 103.905 ;
        RECT 80.775 103.575 81.350 103.905 ;
        RECT 81.530 103.575 81.965 103.905 ;
        RECT 82.145 103.575 82.415 103.905 ;
        RECT 79.890 103.205 82.375 103.395 ;
        RECT 84.180 103.210 84.520 104.040 ;
        RECT 86.000 103.530 86.350 104.780 ;
        RECT 88.115 104.125 91.625 105.215 ;
        RECT 88.115 103.435 89.765 103.955 ;
        RECT 89.935 103.605 91.625 104.125 ;
        RECT 92.715 104.050 93.005 105.215 ;
        RECT 93.175 104.075 93.450 105.045 ;
        RECT 93.660 104.415 93.940 105.215 ;
        RECT 94.110 104.705 95.725 105.035 ;
        RECT 94.110 104.365 95.285 104.535 ;
        RECT 94.110 104.245 94.280 104.365 ;
        RECT 93.620 104.075 94.280 104.245 ;
        RECT 79.895 102.665 80.640 103.035 ;
        RECT 81.205 102.845 81.460 103.205 ;
        RECT 81.640 102.665 81.970 103.035 ;
        RECT 82.150 102.845 82.375 103.205 ;
        RECT 82.595 102.665 87.940 103.210 ;
        RECT 88.115 102.665 91.625 103.435 ;
        RECT 92.715 102.665 93.005 103.390 ;
        RECT 93.175 103.340 93.345 104.075 ;
        RECT 93.620 103.905 93.790 104.075 ;
        RECT 94.540 103.905 94.785 104.195 ;
        RECT 94.955 104.075 95.285 104.365 ;
        RECT 95.545 103.905 95.715 104.465 ;
        RECT 95.965 104.075 96.225 105.215 ;
        RECT 96.395 104.780 101.740 105.215 ;
        RECT 93.515 103.575 93.790 103.905 ;
        RECT 93.960 103.575 94.785 103.905 ;
        RECT 95.000 103.575 95.715 103.905 ;
        RECT 95.885 103.655 96.220 103.905 ;
        RECT 93.620 103.405 93.790 103.575 ;
        RECT 95.465 103.485 95.715 103.575 ;
        RECT 93.175 102.995 93.450 103.340 ;
        RECT 93.620 103.235 95.285 103.405 ;
        RECT 93.640 102.665 94.015 103.065 ;
        RECT 94.185 102.885 94.355 103.235 ;
        RECT 94.525 102.665 94.855 103.065 ;
        RECT 95.025 102.835 95.285 103.235 ;
        RECT 95.465 103.065 95.795 103.485 ;
        RECT 95.965 102.665 96.225 103.485 ;
        RECT 97.980 103.210 98.320 104.040 ;
        RECT 99.800 103.530 100.150 104.780 ;
        RECT 101.915 104.125 105.425 105.215 ;
        RECT 105.595 104.125 106.805 105.215 ;
        RECT 101.915 103.435 103.565 103.955 ;
        RECT 103.735 103.605 105.425 104.125 ;
        RECT 96.395 102.665 101.740 103.210 ;
        RECT 101.915 102.665 105.425 103.435 ;
        RECT 105.595 103.415 106.115 103.955 ;
        RECT 106.285 103.585 106.805 104.125 ;
        RECT 105.595 102.665 106.805 103.415 ;
        RECT 106.975 102.835 107.725 105.045 ;
        RECT 107.895 104.660 108.500 105.215 ;
        RECT 108.675 104.705 109.155 105.045 ;
        RECT 109.325 104.670 109.580 105.215 ;
        RECT 107.895 104.560 108.510 104.660 ;
        RECT 108.325 104.535 108.510 104.560 ;
        RECT 107.895 103.940 108.155 104.390 ;
        RECT 108.325 104.290 108.655 104.535 ;
        RECT 108.825 104.215 109.580 104.465 ;
        RECT 109.750 104.345 110.025 105.045 ;
        RECT 108.810 104.180 109.580 104.215 ;
        RECT 108.795 104.170 109.580 104.180 ;
        RECT 108.790 104.155 109.685 104.170 ;
        RECT 108.770 104.140 109.685 104.155 ;
        RECT 108.750 104.130 109.685 104.140 ;
        RECT 108.725 104.120 109.685 104.130 ;
        RECT 108.655 104.090 109.685 104.120 ;
        RECT 108.635 104.060 109.685 104.090 ;
        RECT 108.615 104.030 109.685 104.060 ;
        RECT 108.585 104.005 109.685 104.030 ;
        RECT 108.550 103.970 109.685 104.005 ;
        RECT 108.520 103.965 109.685 103.970 ;
        RECT 108.520 103.960 108.910 103.965 ;
        RECT 108.520 103.950 108.885 103.960 ;
        RECT 108.520 103.945 108.870 103.950 ;
        RECT 108.520 103.940 108.855 103.945 ;
        RECT 107.895 103.935 108.855 103.940 ;
        RECT 107.895 103.925 108.845 103.935 ;
        RECT 107.895 103.920 108.835 103.925 ;
        RECT 107.895 103.910 108.825 103.920 ;
        RECT 107.895 103.900 108.820 103.910 ;
        RECT 107.895 103.895 108.815 103.900 ;
        RECT 107.895 103.880 108.805 103.895 ;
        RECT 107.895 103.865 108.800 103.880 ;
        RECT 107.895 103.840 108.790 103.865 ;
        RECT 107.895 103.770 108.785 103.840 ;
        RECT 107.895 103.215 108.445 103.600 ;
        RECT 108.615 103.045 108.785 103.770 ;
        RECT 107.895 102.875 108.785 103.045 ;
        RECT 108.955 103.370 109.285 103.795 ;
        RECT 109.455 103.570 109.685 103.965 ;
        RECT 108.955 102.885 109.175 103.370 ;
        RECT 109.855 103.315 110.025 104.345 ;
        RECT 110.205 104.075 110.535 105.215 ;
        RECT 111.065 104.245 111.395 105.030 ;
        RECT 110.715 104.075 111.395 104.245 ;
        RECT 112.115 104.285 112.295 105.045 ;
        RECT 112.475 104.455 112.805 105.215 ;
        RECT 112.115 104.115 112.790 104.285 ;
        RECT 112.975 104.140 113.245 105.045 ;
        RECT 113.415 104.705 114.605 104.995 ;
        RECT 110.195 103.655 110.545 103.905 ;
        RECT 110.715 103.475 110.885 104.075 ;
        RECT 112.620 103.970 112.790 104.115 ;
        RECT 111.055 103.655 111.405 103.905 ;
        RECT 112.055 103.565 112.395 103.935 ;
        RECT 112.620 103.640 112.895 103.970 ;
        RECT 109.345 102.665 109.595 103.205 ;
        RECT 109.765 102.835 110.025 103.315 ;
        RECT 110.205 102.665 110.475 103.475 ;
        RECT 110.645 102.835 110.975 103.475 ;
        RECT 111.145 102.665 111.385 103.475 ;
        RECT 112.620 103.385 112.790 103.640 ;
        RECT 112.125 103.215 112.790 103.385 ;
        RECT 113.065 103.340 113.245 104.140 ;
        RECT 113.435 104.365 114.605 104.535 ;
        RECT 114.775 104.415 115.055 105.215 ;
        RECT 113.435 104.075 113.760 104.365 ;
        RECT 114.435 104.245 114.605 104.365 ;
        RECT 113.930 103.905 114.125 104.195 ;
        RECT 114.435 104.075 115.095 104.245 ;
        RECT 115.265 104.075 115.540 105.045 ;
        RECT 116.215 104.875 117.355 105.045 ;
        RECT 116.215 104.415 116.515 104.875 ;
        RECT 116.685 104.245 117.015 104.705 ;
        RECT 116.255 104.195 117.015 104.245 ;
        RECT 114.925 103.905 115.095 104.075 ;
        RECT 113.415 103.575 113.760 103.905 ;
        RECT 113.930 103.575 114.755 103.905 ;
        RECT 114.925 103.575 115.200 103.905 ;
        RECT 114.925 103.405 115.095 103.575 ;
        RECT 112.125 102.835 112.295 103.215 ;
        RECT 112.475 102.665 112.805 103.045 ;
        RECT 112.985 102.835 113.245 103.340 ;
        RECT 113.430 103.235 115.095 103.405 ;
        RECT 115.370 103.340 115.540 104.075 ;
        RECT 116.235 104.025 117.015 104.195 ;
        RECT 117.185 104.245 117.355 104.875 ;
        RECT 117.525 104.415 117.855 105.215 ;
        RECT 118.025 104.245 118.300 105.045 ;
        RECT 117.185 104.035 118.300 104.245 ;
        RECT 118.475 104.050 118.765 105.215 ;
        RECT 118.975 104.075 119.205 105.215 ;
        RECT 119.375 104.065 119.705 105.045 ;
        RECT 119.875 104.075 120.085 105.215 ;
        RECT 120.445 104.875 122.495 105.045 ;
        RECT 120.445 104.375 120.695 104.875 ;
        RECT 120.865 104.205 121.075 104.705 ;
        RECT 121.285 104.375 121.495 104.875 ;
        RECT 121.825 104.205 122.075 104.705 ;
        RECT 122.245 104.375 122.495 104.875 ;
        RECT 122.665 104.205 122.915 105.045 ;
        RECT 123.085 104.375 123.335 105.215 ;
        RECT 123.505 104.205 123.760 105.045 ;
        RECT 113.430 102.885 113.685 103.235 ;
        RECT 113.855 102.665 114.185 103.065 ;
        RECT 114.355 102.885 114.525 103.235 ;
        RECT 114.695 102.665 115.075 103.065 ;
        RECT 115.265 102.995 115.540 103.340 ;
        RECT 116.255 103.485 116.470 104.025 ;
        RECT 116.640 103.655 117.410 103.855 ;
        RECT 117.580 103.655 118.300 103.855 ;
        RECT 118.955 103.655 119.285 103.905 ;
        RECT 116.255 103.315 117.855 103.485 ;
        RECT 116.685 103.305 117.855 103.315 ;
        RECT 116.225 102.665 116.515 103.135 ;
        RECT 116.685 102.835 117.015 103.305 ;
        RECT 117.185 102.665 117.355 103.135 ;
        RECT 117.525 102.835 117.855 103.305 ;
        RECT 118.025 102.665 118.300 103.485 ;
        RECT 118.475 102.665 118.765 103.390 ;
        RECT 118.975 102.665 119.205 103.485 ;
        RECT 119.455 103.465 119.705 104.065 ;
        RECT 120.315 104.035 121.075 104.205 ;
        RECT 120.315 103.485 120.775 104.035 ;
        RECT 121.270 103.865 121.535 104.205 ;
        RECT 121.825 104.035 123.760 104.205 ;
        RECT 123.995 104.125 125.205 105.215 ;
        RECT 120.945 103.655 121.535 103.865 ;
        RECT 121.725 103.655 122.775 103.865 ;
        RECT 122.945 103.655 123.775 103.865 ;
        RECT 123.995 103.585 124.515 104.125 ;
        RECT 119.375 102.835 119.705 103.465 ;
        RECT 119.875 102.665 120.085 103.485 ;
        RECT 120.315 103.305 123.375 103.485 ;
        RECT 120.365 102.665 120.655 103.135 ;
        RECT 120.825 102.835 121.155 103.305 ;
        RECT 121.325 102.665 122.035 103.135 ;
        RECT 122.205 102.835 122.535 103.305 ;
        RECT 122.705 102.665 122.875 103.135 ;
        RECT 123.045 102.835 123.375 103.305 ;
        RECT 123.545 102.665 123.820 103.485 ;
        RECT 124.685 103.415 125.205 103.955 ;
        RECT 123.995 102.665 125.205 103.415 ;
        RECT 53.990 102.495 125.290 102.665 ;
        RECT 54.075 101.745 55.285 102.495 ;
        RECT 54.075 101.205 54.595 101.745 ;
        RECT 55.460 101.655 55.720 102.495 ;
        RECT 55.895 101.750 56.150 102.325 ;
        RECT 56.320 102.115 56.650 102.495 ;
        RECT 56.865 101.945 57.035 102.325 ;
        RECT 56.320 101.775 57.035 101.945 ;
        RECT 57.295 101.995 57.555 102.325 ;
        RECT 57.765 102.015 58.040 102.495 ;
        RECT 54.765 101.035 55.285 101.575 ;
        RECT 54.075 99.945 55.285 101.035 ;
        RECT 55.460 99.945 55.720 101.095 ;
        RECT 55.895 101.020 56.065 101.750 ;
        RECT 56.320 101.585 56.490 101.775 ;
        RECT 56.235 101.255 56.490 101.585 ;
        RECT 56.320 101.045 56.490 101.255 ;
        RECT 56.770 101.225 57.125 101.595 ;
        RECT 57.295 101.085 57.465 101.995 ;
        RECT 58.250 101.925 58.455 102.325 ;
        RECT 58.625 102.095 58.960 102.495 ;
        RECT 57.635 101.255 57.995 101.835 ;
        RECT 58.250 101.755 58.935 101.925 ;
        RECT 58.175 101.085 58.425 101.585 ;
        RECT 55.895 100.115 56.150 101.020 ;
        RECT 56.320 100.875 57.035 101.045 ;
        RECT 56.320 99.945 56.650 100.705 ;
        RECT 56.865 100.115 57.035 100.875 ;
        RECT 57.295 100.915 58.425 101.085 ;
        RECT 57.295 100.145 57.565 100.915 ;
        RECT 58.595 100.725 58.935 101.755 ;
        RECT 57.735 99.945 58.065 100.725 ;
        RECT 58.270 100.550 58.935 100.725 ;
        RECT 59.135 101.820 59.395 102.325 ;
        RECT 59.575 102.115 59.905 102.495 ;
        RECT 60.085 101.945 60.255 102.325 ;
        RECT 60.515 101.950 65.860 102.495 ;
        RECT 59.135 101.020 59.305 101.820 ;
        RECT 59.590 101.775 60.255 101.945 ;
        RECT 59.590 101.520 59.760 101.775 ;
        RECT 59.475 101.190 59.760 101.520 ;
        RECT 59.995 101.225 60.325 101.595 ;
        RECT 59.590 101.045 59.760 101.190 ;
        RECT 62.100 101.120 62.440 101.950 ;
        RECT 66.555 101.675 66.765 102.495 ;
        RECT 66.935 101.695 67.265 102.325 ;
        RECT 58.270 100.145 58.455 100.550 ;
        RECT 58.625 99.945 58.960 100.370 ;
        RECT 59.135 100.115 59.405 101.020 ;
        RECT 59.590 100.875 60.255 101.045 ;
        RECT 59.575 99.945 59.905 100.705 ;
        RECT 60.085 100.115 60.255 100.875 ;
        RECT 63.920 100.380 64.270 101.630 ;
        RECT 66.935 101.095 67.185 101.695 ;
        RECT 67.435 101.675 67.665 102.495 ;
        RECT 68.075 101.865 68.405 102.225 ;
        RECT 69.035 102.035 69.285 102.495 ;
        RECT 69.455 102.035 70.005 102.325 ;
        RECT 68.075 101.675 69.465 101.865 ;
        RECT 69.295 101.585 69.465 101.675 ;
        RECT 67.355 101.255 67.685 101.505 ;
        RECT 67.875 101.255 68.565 101.505 ;
        RECT 68.795 101.255 69.125 101.505 ;
        RECT 69.295 101.255 69.585 101.585 ;
        RECT 60.515 99.945 65.860 100.380 ;
        RECT 66.555 99.945 66.765 101.085 ;
        RECT 66.935 100.115 67.265 101.095 ;
        RECT 67.435 99.945 67.665 101.085 ;
        RECT 67.875 100.815 68.190 101.255 ;
        RECT 69.295 101.005 69.465 101.255 ;
        RECT 68.525 100.835 69.465 101.005 ;
        RECT 68.075 99.945 68.355 100.615 ;
        RECT 68.525 100.285 68.825 100.835 ;
        RECT 69.755 100.665 70.005 102.035 ;
        RECT 70.175 101.695 70.465 102.495 ;
        RECT 70.640 101.755 70.895 102.325 ;
        RECT 71.065 102.095 71.395 102.495 ;
        RECT 71.820 101.960 72.350 102.325 ;
        RECT 71.820 101.925 71.995 101.960 ;
        RECT 71.065 101.755 71.995 101.925 ;
        RECT 70.640 101.085 70.810 101.755 ;
        RECT 71.065 101.585 71.235 101.755 ;
        RECT 70.980 101.255 71.235 101.585 ;
        RECT 71.460 101.255 71.655 101.585 ;
        RECT 69.035 99.945 69.365 100.665 ;
        RECT 69.555 100.115 70.005 100.665 ;
        RECT 70.175 99.945 70.465 101.085 ;
        RECT 70.640 100.115 70.975 101.085 ;
        RECT 71.145 99.945 71.315 101.085 ;
        RECT 71.485 100.285 71.655 101.255 ;
        RECT 71.825 100.625 71.995 101.755 ;
        RECT 72.165 100.965 72.335 101.765 ;
        RECT 72.540 101.475 72.815 102.325 ;
        RECT 72.535 101.305 72.815 101.475 ;
        RECT 72.540 101.165 72.815 101.305 ;
        RECT 72.985 100.965 73.175 102.325 ;
        RECT 73.355 101.960 73.865 102.495 ;
        RECT 74.085 101.685 74.330 102.290 ;
        RECT 74.775 101.725 76.445 102.495 ;
        RECT 76.780 101.985 77.020 102.495 ;
        RECT 77.200 101.985 77.480 102.315 ;
        RECT 77.710 101.985 77.925 102.495 ;
        RECT 73.375 101.515 74.605 101.685 ;
        RECT 72.165 100.795 73.175 100.965 ;
        RECT 73.345 100.950 74.095 101.140 ;
        RECT 71.825 100.455 72.950 100.625 ;
        RECT 73.345 100.285 73.515 100.950 ;
        RECT 74.265 100.705 74.605 101.515 ;
        RECT 74.775 101.205 75.525 101.725 ;
        RECT 75.695 101.035 76.445 101.555 ;
        RECT 76.675 101.255 77.030 101.815 ;
        RECT 77.200 101.085 77.370 101.985 ;
        RECT 77.540 101.255 77.805 101.815 ;
        RECT 78.095 101.755 78.710 102.325 ;
        RECT 79.835 101.770 80.125 102.495 ;
        RECT 78.055 101.085 78.225 101.585 ;
        RECT 71.485 100.115 73.515 100.285 ;
        RECT 73.685 99.945 73.855 100.705 ;
        RECT 74.090 100.295 74.605 100.705 ;
        RECT 74.775 99.945 76.445 101.035 ;
        RECT 76.800 100.915 78.225 101.085 ;
        RECT 76.800 100.740 77.190 100.915 ;
        RECT 77.675 99.945 78.005 100.745 ;
        RECT 78.395 100.735 78.710 101.755 ;
        RECT 80.295 101.675 80.980 102.315 ;
        RECT 81.150 101.675 81.320 102.495 ;
        RECT 81.490 101.845 81.820 102.310 ;
        RECT 81.990 102.025 82.160 102.495 ;
        RECT 82.420 102.105 83.605 102.275 ;
        RECT 83.775 101.935 84.105 102.325 ;
        RECT 82.805 101.845 83.190 101.935 ;
        RECT 81.490 101.675 83.190 101.845 ;
        RECT 83.595 101.755 84.105 101.935 ;
        RECT 84.445 101.775 84.775 102.495 ;
        RECT 85.320 102.095 86.935 102.265 ;
        RECT 87.105 102.095 87.435 102.495 ;
        RECT 86.765 101.925 86.935 102.095 ;
        RECT 87.605 102.020 87.940 102.280 ;
        RECT 78.175 100.115 78.710 100.735 ;
        RECT 79.835 99.945 80.125 101.110 ;
        RECT 80.295 100.705 80.545 101.675 ;
        RECT 80.715 101.295 81.050 101.505 ;
        RECT 81.220 101.295 81.670 101.505 ;
        RECT 81.860 101.295 82.345 101.505 ;
        RECT 80.880 101.125 81.050 101.295 ;
        RECT 81.970 101.135 82.345 101.295 ;
        RECT 82.535 101.255 82.915 101.505 ;
        RECT 83.095 101.295 83.425 101.505 ;
        RECT 80.880 100.955 81.800 101.125 ;
        RECT 80.295 100.115 80.960 100.705 ;
        RECT 81.130 99.945 81.460 100.785 ;
        RECT 81.630 100.705 81.800 100.955 ;
        RECT 81.970 100.965 82.365 101.135 ;
        RECT 81.970 100.875 82.345 100.965 ;
        RECT 82.535 100.875 82.855 101.255 ;
        RECT 83.595 101.125 83.765 101.755 ;
        RECT 83.935 101.295 84.265 101.585 ;
        RECT 84.500 101.475 84.850 101.585 ;
        RECT 84.495 101.305 84.850 101.475 ;
        RECT 84.500 101.255 84.850 101.305 ;
        RECT 85.160 101.255 85.580 101.920 ;
        RECT 85.750 101.815 86.040 101.915 ;
        RECT 86.230 101.815 86.500 101.915 ;
        RECT 85.750 101.645 86.045 101.815 ;
        RECT 86.230 101.645 86.505 101.815 ;
        RECT 86.765 101.755 87.325 101.925 ;
        RECT 85.750 101.255 86.040 101.645 ;
        RECT 86.230 101.255 86.500 101.645 ;
        RECT 87.155 101.585 87.325 101.755 ;
        RECT 86.710 101.475 86.960 101.585 ;
        RECT 86.710 101.305 86.965 101.475 ;
        RECT 86.710 101.255 86.960 101.305 ;
        RECT 87.155 101.255 87.460 101.585 ;
        RECT 83.025 100.955 84.110 101.125 ;
        RECT 84.500 100.965 84.705 101.255 ;
        RECT 87.155 101.085 87.325 101.255 ;
        RECT 83.025 100.705 83.195 100.955 ;
        RECT 81.630 100.535 83.195 100.705 ;
        RECT 81.970 100.115 82.775 100.535 ;
        RECT 83.365 99.945 83.615 100.785 ;
        RECT 83.810 100.115 84.110 100.955 ;
        RECT 84.955 100.915 87.325 101.085 ;
        RECT 84.525 100.285 84.695 100.785 ;
        RECT 84.955 100.455 85.125 100.915 ;
        RECT 85.355 100.535 86.780 100.705 ;
        RECT 85.355 100.285 85.685 100.535 ;
        RECT 84.525 100.115 85.685 100.285 ;
        RECT 85.910 99.945 86.240 100.365 ;
        RECT 86.495 100.115 86.780 100.535 ;
        RECT 87.025 99.945 87.355 100.745 ;
        RECT 87.685 100.665 87.940 102.020 ;
        RECT 88.120 101.730 88.575 102.495 ;
        RECT 88.850 102.115 90.150 102.325 ;
        RECT 90.405 102.135 90.735 102.495 ;
        RECT 89.980 101.965 90.150 102.115 ;
        RECT 90.905 101.995 91.165 102.325 ;
        RECT 90.935 101.985 91.165 101.995 ;
        RECT 89.050 101.505 89.270 101.905 ;
        RECT 88.115 101.305 88.605 101.505 ;
        RECT 88.795 101.295 89.270 101.505 ;
        RECT 89.515 101.505 89.725 101.905 ;
        RECT 89.980 101.840 90.735 101.965 ;
        RECT 89.980 101.795 90.825 101.840 ;
        RECT 90.555 101.675 90.825 101.795 ;
        RECT 89.515 101.295 89.845 101.505 ;
        RECT 90.015 101.235 90.425 101.540 ;
        RECT 87.605 100.155 87.940 100.665 ;
        RECT 88.120 101.065 89.295 101.125 ;
        RECT 90.655 101.100 90.825 101.675 ;
        RECT 90.625 101.065 90.825 101.100 ;
        RECT 88.120 100.955 90.825 101.065 ;
        RECT 88.120 100.335 88.375 100.955 ;
        RECT 88.965 100.895 90.765 100.955 ;
        RECT 88.965 100.865 89.295 100.895 ;
        RECT 90.995 100.795 91.165 101.985 ;
        RECT 91.335 101.950 96.680 102.495 ;
        RECT 92.920 101.120 93.260 101.950 ;
        RECT 96.865 101.900 97.115 102.325 ;
        RECT 97.285 102.070 97.615 102.495 ;
        RECT 97.785 102.075 98.875 102.325 ;
        RECT 99.065 102.075 100.155 102.325 ;
        RECT 97.785 101.900 97.955 102.075 ;
        RECT 96.865 101.730 97.955 101.900 ;
        RECT 98.125 101.735 99.815 101.905 ;
        RECT 99.985 101.900 100.155 102.075 ;
        RECT 100.325 102.070 100.655 102.495 ;
        RECT 100.825 101.900 101.145 102.325 ;
        RECT 88.625 100.695 88.810 100.785 ;
        RECT 89.400 100.695 90.235 100.705 ;
        RECT 88.625 100.495 90.235 100.695 ;
        RECT 88.625 100.455 88.855 100.495 ;
        RECT 88.120 100.115 88.455 100.335 ;
        RECT 89.460 99.945 89.815 100.325 ;
        RECT 89.985 100.115 90.235 100.495 ;
        RECT 90.485 99.945 90.735 100.725 ;
        RECT 90.905 100.115 91.165 100.795 ;
        RECT 94.740 100.380 95.090 101.630 ;
        RECT 96.920 101.475 97.550 101.505 ;
        RECT 97.840 101.475 98.470 101.505 ;
        RECT 96.915 101.305 97.550 101.475 ;
        RECT 97.835 101.305 98.470 101.475 ;
        RECT 98.640 101.095 98.930 101.735 ;
        RECT 99.985 101.730 101.145 101.900 ;
        RECT 101.475 101.765 101.765 102.495 ;
        RECT 99.215 101.305 99.870 101.505 ;
        RECT 100.160 101.475 101.270 101.505 ;
        RECT 100.135 101.305 101.270 101.475 ;
        RECT 101.465 101.255 101.765 101.585 ;
        RECT 101.945 101.565 102.175 102.205 ;
        RECT 102.355 101.945 102.665 102.315 ;
        RECT 102.845 102.125 103.515 102.495 ;
        RECT 102.355 101.745 103.585 101.945 ;
        RECT 101.945 101.255 102.470 101.565 ;
        RECT 102.650 101.255 103.115 101.565 ;
        RECT 96.865 100.925 98.930 101.095 ;
        RECT 91.335 99.945 96.680 100.380 ;
        RECT 96.865 100.115 97.115 100.925 ;
        RECT 97.285 100.285 97.535 100.755 ;
        RECT 97.705 100.455 98.035 100.925 ;
        RECT 98.205 100.285 98.375 100.755 ;
        RECT 98.545 100.455 98.930 100.925 ;
        RECT 99.145 100.925 101.075 101.095 ;
        RECT 103.295 101.075 103.585 101.745 ;
        RECT 99.145 100.285 99.395 100.925 ;
        RECT 97.285 100.115 99.395 100.285 ;
        RECT 99.565 99.945 99.735 100.755 ;
        RECT 99.905 100.115 100.235 100.925 ;
        RECT 100.405 99.945 100.575 100.755 ;
        RECT 100.745 100.115 101.075 100.925 ;
        RECT 101.475 100.835 102.635 101.075 ;
        RECT 101.475 100.125 101.735 100.835 ;
        RECT 101.905 99.945 102.235 100.655 ;
        RECT 102.405 100.125 102.635 100.835 ;
        RECT 102.815 100.855 103.585 101.075 ;
        RECT 102.815 100.125 103.085 100.855 ;
        RECT 103.265 99.945 103.605 100.675 ;
        RECT 103.775 100.125 104.035 102.315 ;
        RECT 104.215 101.745 105.425 102.495 ;
        RECT 105.595 101.770 105.885 102.495 ;
        RECT 104.215 101.205 104.735 101.745 ;
        RECT 104.905 101.035 105.425 101.575 ;
        RECT 104.215 99.945 105.425 101.035 ;
        RECT 105.595 99.945 105.885 101.110 ;
        RECT 106.055 100.115 106.335 102.215 ;
        RECT 106.565 102.035 106.735 102.495 ;
        RECT 107.005 102.105 108.255 102.285 ;
        RECT 107.390 101.865 107.755 101.935 ;
        RECT 106.505 101.685 107.755 101.865 ;
        RECT 107.925 101.885 108.255 102.105 ;
        RECT 108.425 102.055 108.595 102.495 ;
        RECT 108.765 101.885 109.105 102.300 ;
        RECT 109.275 102.115 110.165 102.285 ;
        RECT 107.925 101.715 109.105 101.885 ;
        RECT 106.505 101.085 106.780 101.685 ;
        RECT 109.275 101.560 109.825 101.945 ;
        RECT 106.950 101.255 107.305 101.505 ;
        RECT 107.500 101.475 107.965 101.505 ;
        RECT 107.495 101.305 107.965 101.475 ;
        RECT 107.500 101.255 107.965 101.305 ;
        RECT 108.135 101.255 108.465 101.505 ;
        RECT 108.640 101.305 109.105 101.505 ;
        RECT 109.995 101.390 110.165 102.115 ;
        RECT 109.275 101.320 110.165 101.390 ;
        RECT 110.335 101.790 110.555 102.275 ;
        RECT 110.725 101.955 110.975 102.495 ;
        RECT 111.145 101.845 111.405 102.325 ;
        RECT 111.575 102.115 112.465 102.285 ;
        RECT 110.335 101.365 110.665 101.790 ;
        RECT 108.285 101.135 108.465 101.255 ;
        RECT 109.275 101.295 110.170 101.320 ;
        RECT 109.275 101.280 110.180 101.295 ;
        RECT 109.275 101.265 110.185 101.280 ;
        RECT 109.275 101.260 110.195 101.265 ;
        RECT 109.275 101.250 110.200 101.260 ;
        RECT 109.275 101.240 110.205 101.250 ;
        RECT 109.275 101.235 110.215 101.240 ;
        RECT 109.275 101.225 110.225 101.235 ;
        RECT 109.275 101.220 110.235 101.225 ;
        RECT 106.505 100.875 108.115 101.085 ;
        RECT 108.285 100.965 108.615 101.135 ;
        RECT 107.705 100.775 108.115 100.875 ;
        RECT 106.525 99.945 107.310 100.705 ;
        RECT 107.705 100.115 108.090 100.775 ;
        RECT 108.415 100.175 108.615 100.965 ;
        RECT 108.785 99.945 109.105 101.125 ;
        RECT 109.275 100.770 109.535 101.220 ;
        RECT 109.900 101.215 110.235 101.220 ;
        RECT 109.900 101.210 110.250 101.215 ;
        RECT 109.900 101.200 110.265 101.210 ;
        RECT 109.900 101.195 110.290 101.200 ;
        RECT 110.835 101.195 111.065 101.590 ;
        RECT 109.900 101.190 111.065 101.195 ;
        RECT 109.930 101.155 111.065 101.190 ;
        RECT 109.965 101.130 111.065 101.155 ;
        RECT 109.995 101.100 111.065 101.130 ;
        RECT 110.015 101.070 111.065 101.100 ;
        RECT 110.035 101.040 111.065 101.070 ;
        RECT 110.105 101.030 111.065 101.040 ;
        RECT 110.130 101.020 111.065 101.030 ;
        RECT 110.150 101.005 111.065 101.020 ;
        RECT 110.170 100.990 111.065 101.005 ;
        RECT 110.175 100.980 110.960 100.990 ;
        RECT 110.190 100.945 110.960 100.980 ;
        RECT 109.705 100.625 110.035 100.870 ;
        RECT 110.205 100.695 110.960 100.945 ;
        RECT 111.235 100.815 111.405 101.845 ;
        RECT 111.575 101.560 112.125 101.945 ;
        RECT 112.295 101.390 112.465 102.115 ;
        RECT 109.705 100.600 109.890 100.625 ;
        RECT 109.275 100.500 109.890 100.600 ;
        RECT 109.275 99.945 109.880 100.500 ;
        RECT 110.055 100.115 110.535 100.455 ;
        RECT 110.705 99.945 110.960 100.490 ;
        RECT 111.130 100.115 111.405 100.815 ;
        RECT 111.575 101.320 112.465 101.390 ;
        RECT 112.635 101.790 112.855 102.275 ;
        RECT 113.025 101.955 113.275 102.495 ;
        RECT 113.445 101.845 113.705 102.325 ;
        RECT 114.795 101.985 115.100 102.495 ;
        RECT 112.635 101.365 112.965 101.790 ;
        RECT 111.575 101.295 112.470 101.320 ;
        RECT 111.575 101.280 112.480 101.295 ;
        RECT 111.575 101.265 112.485 101.280 ;
        RECT 111.575 101.260 112.495 101.265 ;
        RECT 111.575 101.250 112.500 101.260 ;
        RECT 111.575 101.240 112.505 101.250 ;
        RECT 111.575 101.235 112.515 101.240 ;
        RECT 111.575 101.225 112.525 101.235 ;
        RECT 111.575 101.220 112.535 101.225 ;
        RECT 111.575 100.770 111.835 101.220 ;
        RECT 112.200 101.215 112.535 101.220 ;
        RECT 112.200 101.210 112.550 101.215 ;
        RECT 112.200 101.200 112.565 101.210 ;
        RECT 112.200 101.195 112.590 101.200 ;
        RECT 113.135 101.195 113.365 101.590 ;
        RECT 112.200 101.190 113.365 101.195 ;
        RECT 112.230 101.155 113.365 101.190 ;
        RECT 112.265 101.130 113.365 101.155 ;
        RECT 112.295 101.100 113.365 101.130 ;
        RECT 112.315 101.070 113.365 101.100 ;
        RECT 112.335 101.040 113.365 101.070 ;
        RECT 112.405 101.030 113.365 101.040 ;
        RECT 112.430 101.020 113.365 101.030 ;
        RECT 112.450 101.005 113.365 101.020 ;
        RECT 112.470 100.990 113.365 101.005 ;
        RECT 112.475 100.980 113.260 100.990 ;
        RECT 112.490 100.945 113.260 100.980 ;
        RECT 112.005 100.625 112.335 100.870 ;
        RECT 112.505 100.695 113.260 100.945 ;
        RECT 113.535 100.815 113.705 101.845 ;
        RECT 114.795 101.255 115.110 101.815 ;
        RECT 115.280 101.505 115.530 102.315 ;
        RECT 115.700 101.970 115.960 102.495 ;
        RECT 116.140 101.505 116.390 102.315 ;
        RECT 116.560 101.935 116.820 102.495 ;
        RECT 116.990 101.845 117.250 102.300 ;
        RECT 117.420 102.015 117.680 102.495 ;
        RECT 117.850 101.845 118.110 102.300 ;
        RECT 118.280 102.015 118.540 102.495 ;
        RECT 118.710 101.845 118.970 102.300 ;
        RECT 119.140 102.015 119.385 102.495 ;
        RECT 119.555 101.845 119.830 102.300 ;
        RECT 120.000 102.015 120.245 102.495 ;
        RECT 120.415 101.845 120.675 102.300 ;
        RECT 120.855 102.015 121.105 102.495 ;
        RECT 121.275 101.845 121.535 102.300 ;
        RECT 121.715 102.015 121.965 102.495 ;
        RECT 122.135 101.845 122.395 102.300 ;
        RECT 122.575 102.015 122.835 102.495 ;
        RECT 123.005 101.845 123.265 102.300 ;
        RECT 123.435 102.015 123.735 102.495 ;
        RECT 116.990 101.675 123.735 101.845 ;
        RECT 123.995 101.745 125.205 102.495 ;
        RECT 115.280 101.255 122.400 101.505 ;
        RECT 112.005 100.600 112.190 100.625 ;
        RECT 111.575 100.500 112.190 100.600 ;
        RECT 111.575 99.945 112.180 100.500 ;
        RECT 112.355 100.115 112.835 100.455 ;
        RECT 113.005 99.945 113.260 100.490 ;
        RECT 113.430 100.115 113.705 100.815 ;
        RECT 114.805 99.945 115.100 100.755 ;
        RECT 115.280 100.115 115.525 101.255 ;
        RECT 115.700 99.945 115.960 100.755 ;
        RECT 116.140 100.120 116.390 101.255 ;
        RECT 122.570 101.085 123.735 101.675 ;
        RECT 116.990 100.860 123.735 101.085 ;
        RECT 123.995 101.035 124.515 101.575 ;
        RECT 124.685 101.205 125.205 101.745 ;
        RECT 116.990 100.845 122.395 100.860 ;
        RECT 116.560 99.950 116.820 100.745 ;
        RECT 116.990 100.120 117.250 100.845 ;
        RECT 117.420 99.950 117.680 100.675 ;
        RECT 117.850 100.120 118.110 100.845 ;
        RECT 118.280 99.950 118.540 100.675 ;
        RECT 118.710 100.120 118.970 100.845 ;
        RECT 119.140 99.950 119.400 100.675 ;
        RECT 119.570 100.120 119.830 100.845 ;
        RECT 120.000 99.950 120.245 100.675 ;
        RECT 120.415 100.120 120.675 100.845 ;
        RECT 120.860 99.950 121.105 100.675 ;
        RECT 121.275 100.120 121.535 100.845 ;
        RECT 121.720 99.950 121.965 100.675 ;
        RECT 122.135 100.120 122.395 100.845 ;
        RECT 122.580 99.950 122.835 100.675 ;
        RECT 123.005 100.120 123.295 100.860 ;
        RECT 116.560 99.945 122.835 99.950 ;
        RECT 123.465 99.945 123.735 100.690 ;
        RECT 123.995 99.945 125.205 101.035 ;
        RECT 53.990 99.775 125.290 99.945 ;
        RECT 54.075 98.685 55.285 99.775 ;
        RECT 54.075 97.975 54.595 98.515 ;
        RECT 54.765 98.145 55.285 98.685 ;
        RECT 56.380 98.635 56.700 99.775 ;
        RECT 56.880 98.465 57.075 99.515 ;
        RECT 57.255 98.925 57.585 99.605 ;
        RECT 57.785 98.975 58.040 99.775 ;
        RECT 58.305 99.155 58.475 99.585 ;
        RECT 58.645 99.325 58.975 99.775 ;
        RECT 58.305 98.925 58.985 99.155 ;
        RECT 57.255 98.645 57.605 98.925 ;
        RECT 56.440 98.415 56.700 98.465 ;
        RECT 56.435 98.245 56.700 98.415 ;
        RECT 56.440 98.135 56.700 98.245 ;
        RECT 56.880 98.135 57.265 98.465 ;
        RECT 57.435 98.265 57.605 98.645 ;
        RECT 57.795 98.435 58.040 98.795 ;
        RECT 57.435 98.095 57.955 98.265 ;
        RECT 54.075 97.225 55.285 97.975 ;
        RECT 56.380 97.755 57.595 97.925 ;
        RECT 56.380 97.405 56.670 97.755 ;
        RECT 56.865 97.225 57.195 97.585 ;
        RECT 57.365 97.450 57.595 97.755 ;
        RECT 57.785 97.530 57.955 98.095 ;
        RECT 58.280 98.075 58.580 98.755 ;
        RECT 58.275 97.905 58.580 98.075 ;
        RECT 58.750 98.275 58.985 98.925 ;
        RECT 59.175 98.615 59.460 99.560 ;
        RECT 59.640 99.305 60.325 99.775 ;
        RECT 59.635 98.785 60.330 99.095 ;
        RECT 60.505 98.720 60.810 99.505 ;
        RECT 60.995 98.820 61.265 99.775 ;
        RECT 61.440 98.975 61.695 99.775 ;
        RECT 61.895 98.925 62.225 99.605 ;
        RECT 59.175 98.465 60.035 98.615 ;
        RECT 59.175 98.445 60.465 98.465 ;
        RECT 58.750 97.945 59.305 98.275 ;
        RECT 59.475 98.085 60.465 98.445 ;
        RECT 58.750 97.795 58.965 97.945 ;
        RECT 58.225 97.225 58.555 97.730 ;
        RECT 58.725 97.420 58.965 97.795 ;
        RECT 59.475 97.750 59.645 98.085 ;
        RECT 60.635 97.915 60.810 98.720 ;
        RECT 61.440 98.435 61.685 98.795 ;
        RECT 61.875 98.645 62.225 98.925 ;
        RECT 61.875 98.265 62.045 98.645 ;
        RECT 62.405 98.465 62.600 99.515 ;
        RECT 62.780 98.635 63.100 99.775 ;
        RECT 63.275 98.685 66.785 99.775 ;
        RECT 59.245 97.555 59.645 97.750 ;
        RECT 59.245 97.410 59.415 97.555 ;
        RECT 60.005 97.225 60.405 97.720 ;
        RECT 60.575 97.395 60.810 97.915 ;
        RECT 61.525 98.095 62.045 98.265 ;
        RECT 62.215 98.135 62.600 98.465 ;
        RECT 62.780 98.415 63.040 98.465 ;
        RECT 62.780 98.245 63.045 98.415 ;
        RECT 62.780 98.135 63.040 98.245 ;
        RECT 60.995 97.225 61.265 97.860 ;
        RECT 61.525 97.530 61.695 98.095 ;
        RECT 63.275 97.995 64.925 98.515 ;
        RECT 65.095 98.165 66.785 98.685 ;
        RECT 66.955 98.610 67.245 99.775 ;
        RECT 67.420 98.625 67.680 99.775 ;
        RECT 67.855 98.700 68.110 99.605 ;
        RECT 68.280 99.015 68.610 99.775 ;
        RECT 68.825 98.845 68.995 99.605 ;
        RECT 61.885 97.755 63.100 97.925 ;
        RECT 61.885 97.450 62.115 97.755 ;
        RECT 62.285 97.225 62.615 97.585 ;
        RECT 62.810 97.405 63.100 97.755 ;
        RECT 63.275 97.225 66.785 97.995 ;
        RECT 66.955 97.225 67.245 97.950 ;
        RECT 67.420 97.225 67.680 98.065 ;
        RECT 67.855 97.970 68.025 98.700 ;
        RECT 68.280 98.675 68.995 98.845 ;
        RECT 69.255 98.685 72.765 99.775 ;
        RECT 74.055 99.105 74.335 99.775 ;
        RECT 74.505 98.885 74.805 99.435 ;
        RECT 75.005 99.055 75.335 99.775 ;
        RECT 75.525 99.055 75.985 99.605 ;
        RECT 76.155 99.340 81.500 99.775 ;
        RECT 68.280 98.465 68.450 98.675 ;
        RECT 68.195 98.135 68.450 98.465 ;
        RECT 67.855 97.395 68.110 97.970 ;
        RECT 68.280 97.945 68.450 98.135 ;
        RECT 68.730 98.125 69.085 98.495 ;
        RECT 69.255 97.995 70.905 98.515 ;
        RECT 71.075 98.165 72.765 98.685 ;
        RECT 73.870 98.465 74.135 98.825 ;
        RECT 74.505 98.715 75.445 98.885 ;
        RECT 75.275 98.465 75.445 98.715 ;
        RECT 73.870 98.215 74.545 98.465 ;
        RECT 74.765 98.215 75.105 98.465 ;
        RECT 75.275 98.135 75.565 98.465 ;
        RECT 75.275 98.045 75.445 98.135 ;
        RECT 68.280 97.775 68.995 97.945 ;
        RECT 68.280 97.225 68.610 97.605 ;
        RECT 68.825 97.395 68.995 97.775 ;
        RECT 69.255 97.225 72.765 97.995 ;
        RECT 74.055 97.855 75.445 98.045 ;
        RECT 74.055 97.495 74.385 97.855 ;
        RECT 75.735 97.685 75.985 99.055 ;
        RECT 77.740 97.770 78.080 98.600 ;
        RECT 79.560 98.090 79.910 99.340 ;
        RECT 81.675 98.685 83.345 99.775 ;
        RECT 81.675 97.995 82.425 98.515 ;
        RECT 82.595 98.165 83.345 98.685 ;
        RECT 83.515 98.170 83.795 99.605 ;
        RECT 83.965 99.000 84.675 99.775 ;
        RECT 84.845 98.830 85.175 99.605 ;
        RECT 84.025 98.615 85.175 98.830 ;
        RECT 75.005 97.225 75.255 97.685 ;
        RECT 75.425 97.395 75.985 97.685 ;
        RECT 76.155 97.225 81.500 97.770 ;
        RECT 81.675 97.225 83.345 97.995 ;
        RECT 83.515 97.395 83.855 98.170 ;
        RECT 84.025 98.045 84.310 98.615 ;
        RECT 84.495 98.215 84.965 98.445 ;
        RECT 85.370 98.415 85.585 99.530 ;
        RECT 85.765 99.055 86.095 99.775 ;
        RECT 85.875 98.415 86.105 98.755 ;
        RECT 86.275 98.685 87.945 99.775 ;
        RECT 88.205 99.155 88.375 99.585 ;
        RECT 88.545 99.325 88.875 99.775 ;
        RECT 88.205 98.925 88.885 99.155 ;
        RECT 85.135 98.235 85.585 98.415 ;
        RECT 85.135 98.215 85.465 98.235 ;
        RECT 85.775 98.215 86.105 98.415 ;
        RECT 84.025 97.855 84.735 98.045 ;
        RECT 84.435 97.715 84.735 97.855 ;
        RECT 84.925 97.855 86.105 98.045 ;
        RECT 84.925 97.775 85.255 97.855 ;
        RECT 84.435 97.705 84.750 97.715 ;
        RECT 84.435 97.695 84.760 97.705 ;
        RECT 84.435 97.690 84.770 97.695 ;
        RECT 84.025 97.225 84.195 97.685 ;
        RECT 84.435 97.680 84.775 97.690 ;
        RECT 84.435 97.675 84.780 97.680 ;
        RECT 84.435 97.665 84.785 97.675 ;
        RECT 84.435 97.660 84.790 97.665 ;
        RECT 84.435 97.395 84.795 97.660 ;
        RECT 85.425 97.225 85.595 97.685 ;
        RECT 85.765 97.395 86.105 97.855 ;
        RECT 86.275 97.995 87.025 98.515 ;
        RECT 87.195 98.165 87.945 98.685 ;
        RECT 88.180 98.415 88.480 98.755 ;
        RECT 88.175 98.245 88.480 98.415 ;
        RECT 86.275 97.225 87.945 97.995 ;
        RECT 88.180 97.905 88.480 98.245 ;
        RECT 88.650 98.275 88.885 98.925 ;
        RECT 89.075 98.615 89.360 99.560 ;
        RECT 89.540 99.305 90.225 99.775 ;
        RECT 89.535 98.785 90.230 99.095 ;
        RECT 90.405 98.720 90.710 99.505 ;
        RECT 90.895 98.820 91.165 99.775 ;
        RECT 89.075 98.465 89.935 98.615 ;
        RECT 89.075 98.445 90.365 98.465 ;
        RECT 88.650 97.945 89.205 98.275 ;
        RECT 89.375 98.085 90.365 98.445 ;
        RECT 88.650 97.795 88.865 97.945 ;
        RECT 88.125 97.225 88.455 97.730 ;
        RECT 88.625 97.420 88.865 97.795 ;
        RECT 89.375 97.750 89.545 98.085 ;
        RECT 90.535 97.915 90.710 98.720 ;
        RECT 91.335 98.685 92.545 99.775 ;
        RECT 89.145 97.555 89.545 97.750 ;
        RECT 89.145 97.410 89.315 97.555 ;
        RECT 89.905 97.225 90.305 97.720 ;
        RECT 90.475 97.395 90.710 97.915 ;
        RECT 91.335 97.975 91.855 98.515 ;
        RECT 92.025 98.145 92.545 98.685 ;
        RECT 92.715 98.610 93.005 99.775 ;
        RECT 93.615 98.635 93.955 99.775 ;
        RECT 94.125 99.095 94.295 99.605 ;
        RECT 94.505 99.275 94.755 99.775 ;
        RECT 94.965 99.395 96.225 99.605 ;
        RECT 94.965 99.095 95.215 99.395 ;
        RECT 94.125 98.925 95.215 99.095 ;
        RECT 95.445 98.925 95.795 99.225 ;
        RECT 95.965 98.975 96.225 99.395 ;
        RECT 94.125 98.885 94.295 98.925 ;
        RECT 95.055 98.565 95.455 98.755 ;
        RECT 93.560 98.155 93.975 98.465 ;
        RECT 94.145 98.135 94.505 98.465 ;
        RECT 94.715 98.215 95.080 98.395 ;
        RECT 90.895 97.225 91.165 97.860 ;
        RECT 91.335 97.225 92.545 97.975 ;
        RECT 92.715 97.225 93.005 97.950 ;
        RECT 93.615 97.225 93.955 97.945 ;
        RECT 94.145 97.555 94.345 98.135 ;
        RECT 94.715 97.905 94.905 98.215 ;
        RECT 95.285 98.135 95.455 98.565 ;
        RECT 95.625 97.945 95.795 98.925 ;
        RECT 96.395 98.685 98.065 99.775 ;
        RECT 95.965 98.135 96.225 98.465 ;
        RECT 94.605 97.485 94.905 97.905 ;
        RECT 95.145 97.775 95.795 97.945 ;
        RECT 96.395 97.995 97.145 98.515 ;
        RECT 97.315 98.165 98.065 98.685 ;
        RECT 98.705 99.165 99.035 99.595 ;
        RECT 99.215 99.335 99.410 99.775 ;
        RECT 99.580 99.165 99.910 99.595 ;
        RECT 98.705 98.995 99.910 99.165 ;
        RECT 98.705 98.665 99.600 98.995 ;
        RECT 100.080 98.825 100.355 99.595 ;
        RECT 101.000 99.265 102.655 99.555 ;
        RECT 99.770 98.635 100.355 98.825 ;
        RECT 101.000 98.925 102.590 99.095 ;
        RECT 102.825 98.975 103.105 99.775 ;
        RECT 101.000 98.635 101.320 98.925 ;
        RECT 102.420 98.805 102.590 98.925 ;
        RECT 98.710 98.135 99.005 98.465 ;
        RECT 99.185 98.135 99.600 98.465 ;
        RECT 95.145 97.735 95.395 97.775 ;
        RECT 95.075 97.565 95.395 97.735 ;
        RECT 95.145 97.435 95.395 97.565 ;
        RECT 95.885 97.225 96.215 97.605 ;
        RECT 96.395 97.225 98.065 97.995 ;
        RECT 98.705 97.225 99.005 97.955 ;
        RECT 99.185 97.515 99.415 98.135 ;
        RECT 99.770 97.965 99.945 98.635 ;
        RECT 101.515 98.585 102.230 98.755 ;
        RECT 102.420 98.635 103.145 98.805 ;
        RECT 103.315 98.635 103.585 99.605 ;
        RECT 103.755 98.685 106.345 99.775 ;
        RECT 106.975 99.220 107.580 99.775 ;
        RECT 107.755 99.265 108.235 99.605 ;
        RECT 108.405 99.230 108.660 99.775 ;
        RECT 106.975 99.120 107.590 99.220 ;
        RECT 107.405 99.095 107.590 99.120 ;
        RECT 99.615 97.785 99.945 97.965 ;
        RECT 100.115 97.815 100.355 98.465 ;
        RECT 101.000 97.895 101.350 98.465 ;
        RECT 101.520 98.135 102.230 98.585 ;
        RECT 102.975 98.465 103.145 98.635 ;
        RECT 102.400 98.135 102.805 98.465 ;
        RECT 102.975 98.135 103.245 98.465 ;
        RECT 102.975 97.965 103.145 98.135 ;
        RECT 101.535 97.795 103.145 97.965 ;
        RECT 103.415 97.900 103.585 98.635 ;
        RECT 99.615 97.405 99.840 97.785 ;
        RECT 100.010 97.225 100.340 97.615 ;
        RECT 101.005 97.225 101.335 97.725 ;
        RECT 101.535 97.445 101.705 97.795 ;
        RECT 101.905 97.225 102.235 97.625 ;
        RECT 102.405 97.445 102.575 97.795 ;
        RECT 102.745 97.225 103.125 97.625 ;
        RECT 103.315 97.555 103.585 97.900 ;
        RECT 103.755 97.995 104.965 98.515 ;
        RECT 105.135 98.165 106.345 98.685 ;
        RECT 106.975 98.500 107.235 98.950 ;
        RECT 107.405 98.850 107.735 99.095 ;
        RECT 107.905 98.775 108.660 99.025 ;
        RECT 108.830 98.905 109.105 99.605 ;
        RECT 107.890 98.740 108.660 98.775 ;
        RECT 107.875 98.730 108.660 98.740 ;
        RECT 107.870 98.715 108.765 98.730 ;
        RECT 107.850 98.700 108.765 98.715 ;
        RECT 107.830 98.690 108.765 98.700 ;
        RECT 107.805 98.680 108.765 98.690 ;
        RECT 107.735 98.650 108.765 98.680 ;
        RECT 107.715 98.620 108.765 98.650 ;
        RECT 107.695 98.590 108.765 98.620 ;
        RECT 107.665 98.565 108.765 98.590 ;
        RECT 107.630 98.530 108.765 98.565 ;
        RECT 107.600 98.525 108.765 98.530 ;
        RECT 107.600 98.520 107.990 98.525 ;
        RECT 107.600 98.510 107.965 98.520 ;
        RECT 107.600 98.505 107.950 98.510 ;
        RECT 107.600 98.500 107.935 98.505 ;
        RECT 106.975 98.495 107.935 98.500 ;
        RECT 106.975 98.485 107.925 98.495 ;
        RECT 106.975 98.480 107.915 98.485 ;
        RECT 106.975 98.470 107.905 98.480 ;
        RECT 106.975 98.460 107.900 98.470 ;
        RECT 106.975 98.455 107.895 98.460 ;
        RECT 106.975 98.440 107.885 98.455 ;
        RECT 106.975 98.425 107.880 98.440 ;
        RECT 106.975 98.400 107.870 98.425 ;
        RECT 106.975 98.330 107.865 98.400 ;
        RECT 103.755 97.225 106.345 97.995 ;
        RECT 106.975 97.775 107.525 98.160 ;
        RECT 107.695 97.605 107.865 98.330 ;
        RECT 106.975 97.435 107.865 97.605 ;
        RECT 108.035 97.930 108.365 98.355 ;
        RECT 108.535 98.130 108.765 98.525 ;
        RECT 108.035 97.445 108.255 97.930 ;
        RECT 108.935 97.875 109.105 98.905 ;
        RECT 109.285 98.635 109.615 99.775 ;
        RECT 110.145 98.805 110.475 99.590 ;
        RECT 109.795 98.635 110.475 98.805 ;
        RECT 110.655 98.685 114.165 99.775 ;
        RECT 109.275 98.215 109.625 98.465 ;
        RECT 109.795 98.035 109.965 98.635 ;
        RECT 110.135 98.215 110.485 98.465 ;
        RECT 108.425 97.225 108.675 97.765 ;
        RECT 108.845 97.395 109.105 97.875 ;
        RECT 109.285 97.225 109.555 98.035 ;
        RECT 109.725 97.395 110.055 98.035 ;
        RECT 110.225 97.225 110.465 98.035 ;
        RECT 110.655 97.995 112.305 98.515 ;
        RECT 112.475 98.165 114.165 98.685 ;
        RECT 115.335 98.845 115.515 99.605 ;
        RECT 115.695 99.015 116.025 99.775 ;
        RECT 115.335 98.675 116.010 98.845 ;
        RECT 116.195 98.700 116.465 99.605 ;
        RECT 116.640 99.350 116.975 99.775 ;
        RECT 117.145 99.170 117.330 99.575 ;
        RECT 115.840 98.530 116.010 98.675 ;
        RECT 115.275 98.125 115.615 98.495 ;
        RECT 115.840 98.200 116.115 98.530 ;
        RECT 110.655 97.225 114.165 97.995 ;
        RECT 115.840 97.945 116.010 98.200 ;
        RECT 115.345 97.775 116.010 97.945 ;
        RECT 116.285 97.900 116.465 98.700 ;
        RECT 115.345 97.395 115.515 97.775 ;
        RECT 115.695 97.225 116.025 97.605 ;
        RECT 116.205 97.395 116.465 97.900 ;
        RECT 116.665 98.995 117.330 99.170 ;
        RECT 117.535 98.995 117.865 99.775 ;
        RECT 116.665 97.965 117.005 98.995 ;
        RECT 118.035 98.805 118.305 99.575 ;
        RECT 117.175 98.635 118.305 98.805 ;
        RECT 117.175 98.135 117.425 98.635 ;
        RECT 116.665 97.795 117.350 97.965 ;
        RECT 117.605 97.885 117.965 98.465 ;
        RECT 116.640 97.225 116.975 97.625 ;
        RECT 117.145 97.395 117.350 97.795 ;
        RECT 118.135 97.725 118.305 98.635 ;
        RECT 118.475 98.610 118.765 99.775 ;
        RECT 119.485 99.195 119.655 99.605 ;
        RECT 119.825 99.395 120.155 99.775 ;
        RECT 120.800 99.395 121.470 99.775 ;
        RECT 121.705 99.225 121.875 99.605 ;
        RECT 122.045 99.395 122.385 99.775 ;
        RECT 122.555 99.225 122.725 99.605 ;
        RECT 123.065 99.395 123.395 99.775 ;
        RECT 123.565 99.225 123.825 99.605 ;
        RECT 119.485 99.025 121.235 99.195 ;
        RECT 119.460 98.415 119.640 98.775 ;
        RECT 119.455 98.245 119.640 98.415 ;
        RECT 119.460 98.135 119.640 98.245 ;
        RECT 117.560 97.225 117.835 97.705 ;
        RECT 118.045 97.395 118.305 97.725 ;
        RECT 118.475 97.225 118.765 97.950 ;
        RECT 119.810 97.945 119.980 99.025 ;
        RECT 120.300 98.685 120.630 98.855 ;
        RECT 119.485 97.775 119.980 97.945 ;
        RECT 119.485 97.395 119.655 97.775 ;
        RECT 119.825 97.225 120.155 97.605 ;
        RECT 120.325 97.395 120.550 98.685 ;
        RECT 121.065 98.465 121.235 99.025 ;
        RECT 121.545 99.055 122.725 99.225 ;
        RECT 122.895 99.055 123.825 99.225 ;
        RECT 120.725 97.945 120.895 98.465 ;
        RECT 121.065 98.135 121.375 98.465 ;
        RECT 121.545 97.945 121.715 99.055 ;
        RECT 122.895 98.885 123.065 99.055 ;
        RECT 121.885 98.715 123.065 98.885 ;
        RECT 121.885 98.540 122.055 98.715 ;
        RECT 122.215 98.245 122.485 98.415 ;
        RECT 120.725 97.775 121.715 97.945 ;
        RECT 120.720 97.225 121.050 97.605 ;
        RECT 121.320 97.395 121.490 97.775 ;
        RECT 122.220 97.560 122.485 98.245 ;
        RECT 122.660 97.565 122.965 98.545 ;
        RECT 123.135 97.905 123.485 98.445 ;
        RECT 123.655 97.725 123.825 99.055 ;
        RECT 123.995 98.685 125.205 99.775 ;
        RECT 123.995 98.145 124.515 98.685 ;
        RECT 124.685 97.975 125.205 98.515 ;
        RECT 123.145 97.225 123.395 97.725 ;
        RECT 123.565 97.395 123.825 97.725 ;
        RECT 123.995 97.225 125.205 97.975 ;
        RECT 53.990 97.055 125.290 97.225 ;
        RECT 54.075 96.305 55.285 97.055 ;
        RECT 55.455 96.485 55.890 96.885 ;
        RECT 56.060 96.655 56.445 97.055 ;
        RECT 55.455 96.315 56.445 96.485 ;
        RECT 56.615 96.315 57.040 96.885 ;
        RECT 57.230 96.485 57.485 96.885 ;
        RECT 57.655 96.655 58.040 97.055 ;
        RECT 57.230 96.315 58.040 96.485 ;
        RECT 58.210 96.315 58.455 96.885 ;
        RECT 58.645 96.485 58.900 96.885 ;
        RECT 59.070 96.655 59.455 97.055 ;
        RECT 58.645 96.315 59.455 96.485 ;
        RECT 59.625 96.315 59.885 96.885 ;
        RECT 61.060 96.485 61.235 96.885 ;
        RECT 61.405 96.675 61.735 97.055 ;
        RECT 61.980 96.555 62.210 96.885 ;
        RECT 61.060 96.315 61.690 96.485 ;
        RECT 54.075 95.765 54.595 96.305 ;
        RECT 56.110 96.145 56.445 96.315 ;
        RECT 56.690 96.145 57.040 96.315 ;
        RECT 57.690 96.145 58.040 96.315 ;
        RECT 58.285 96.145 58.455 96.315 ;
        RECT 59.105 96.145 59.455 96.315 ;
        RECT 54.765 95.595 55.285 96.135 ;
        RECT 54.075 94.505 55.285 95.595 ;
        RECT 55.455 95.440 55.940 96.145 ;
        RECT 56.110 95.815 56.520 96.145 ;
        RECT 56.110 95.270 56.445 95.815 ;
        RECT 56.690 95.645 57.520 96.145 ;
        RECT 55.455 95.100 56.445 95.270 ;
        RECT 56.615 95.465 57.520 95.645 ;
        RECT 57.690 95.815 58.115 96.145 ;
        RECT 55.455 94.675 55.890 95.100 ;
        RECT 56.060 94.505 56.445 94.930 ;
        RECT 56.615 94.675 57.040 95.465 ;
        RECT 57.690 95.295 58.040 95.815 ;
        RECT 58.285 95.645 58.935 96.145 ;
        RECT 57.210 95.100 58.040 95.295 ;
        RECT 58.210 95.465 58.935 95.645 ;
        RECT 59.105 95.815 59.530 96.145 ;
        RECT 57.210 94.675 57.485 95.100 ;
        RECT 57.655 94.505 58.040 94.930 ;
        RECT 58.210 94.675 58.455 95.465 ;
        RECT 59.105 95.295 59.455 95.815 ;
        RECT 59.700 95.645 59.885 96.315 ;
        RECT 61.520 96.145 61.690 96.315 ;
        RECT 58.645 95.100 59.455 95.295 ;
        RECT 58.645 94.675 58.900 95.100 ;
        RECT 59.070 94.505 59.455 94.930 ;
        RECT 59.625 94.675 59.885 95.645 ;
        RECT 60.975 95.465 61.340 96.145 ;
        RECT 61.520 95.815 61.870 96.145 ;
        RECT 61.520 95.295 61.690 95.815 ;
        RECT 61.060 95.125 61.690 95.295 ;
        RECT 62.040 95.265 62.210 96.555 ;
        RECT 62.410 95.445 62.690 96.720 ;
        RECT 62.915 95.695 63.185 96.720 ;
        RECT 63.645 96.675 63.975 97.055 ;
        RECT 64.145 96.800 64.480 96.845 ;
        RECT 62.875 95.525 63.185 95.695 ;
        RECT 62.915 95.445 63.185 95.525 ;
        RECT 63.375 95.445 63.715 96.475 ;
        RECT 64.145 96.335 64.485 96.800 ;
        RECT 63.885 95.815 64.145 96.145 ;
        RECT 63.885 95.265 64.055 95.815 ;
        RECT 64.315 95.645 64.485 96.335 ;
        RECT 61.060 94.675 61.235 95.125 ;
        RECT 62.040 95.095 64.055 95.265 ;
        RECT 61.405 94.505 61.735 94.945 ;
        RECT 62.040 94.675 62.210 95.095 ;
        RECT 62.445 94.505 63.115 94.915 ;
        RECT 63.330 94.675 63.500 95.095 ;
        RECT 63.700 94.505 64.030 94.915 ;
        RECT 64.225 94.675 64.485 95.645 ;
        RECT 64.655 96.555 64.915 96.885 ;
        RECT 65.225 96.675 65.555 97.055 ;
        RECT 65.735 96.715 67.215 96.885 ;
        RECT 64.655 95.855 64.825 96.555 ;
        RECT 65.735 96.385 66.135 96.715 ;
        RECT 65.175 96.195 65.385 96.375 ;
        RECT 65.175 96.025 65.795 96.195 ;
        RECT 65.965 95.905 66.135 96.385 ;
        RECT 66.325 96.215 66.875 96.545 ;
        RECT 64.655 95.685 65.785 95.855 ;
        RECT 65.965 95.735 66.535 95.905 ;
        RECT 64.655 95.005 64.825 95.685 ;
        RECT 65.615 95.565 65.785 95.685 ;
        RECT 64.995 95.185 65.345 95.515 ;
        RECT 65.615 95.395 66.195 95.565 ;
        RECT 66.365 95.225 66.535 95.735 ;
        RECT 65.795 95.055 66.535 95.225 ;
        RECT 66.705 95.225 66.875 96.215 ;
        RECT 67.045 95.815 67.215 96.715 ;
        RECT 67.465 96.145 67.650 96.725 ;
        RECT 67.920 96.145 68.115 96.720 ;
        RECT 68.325 96.675 68.655 97.055 ;
        RECT 67.465 95.815 67.695 96.145 ;
        RECT 67.920 95.815 68.175 96.145 ;
        RECT 67.465 95.505 67.650 95.815 ;
        RECT 67.920 95.505 68.115 95.815 ;
        RECT 68.485 95.225 68.655 96.145 ;
        RECT 66.705 95.055 68.655 95.225 ;
        RECT 64.655 94.675 64.915 95.005 ;
        RECT 65.225 94.505 65.555 94.885 ;
        RECT 65.795 94.675 65.985 95.055 ;
        RECT 66.235 94.505 66.565 94.885 ;
        RECT 66.775 94.675 66.945 95.055 ;
        RECT 67.140 94.505 67.470 94.885 ;
        RECT 67.730 94.675 67.900 95.055 ;
        RECT 68.325 94.505 68.655 94.885 ;
        RECT 68.825 94.675 69.085 96.885 ;
        RECT 69.255 96.285 71.845 97.055 ;
        RECT 72.170 96.405 72.500 96.870 ;
        RECT 72.670 96.585 72.840 97.055 ;
        RECT 73.010 96.405 73.340 96.885 ;
        RECT 69.255 95.765 70.465 96.285 ;
        RECT 72.170 96.235 73.340 96.405 ;
        RECT 70.635 95.595 71.845 96.115 ;
        RECT 72.015 95.855 72.660 96.065 ;
        RECT 72.830 95.855 73.400 96.065 ;
        RECT 73.570 95.685 73.740 96.885 ;
        RECT 74.280 96.485 74.450 96.690 ;
        RECT 69.255 94.505 71.845 95.595 ;
        RECT 72.230 94.505 72.560 95.605 ;
        RECT 73.035 95.275 73.740 95.685 ;
        RECT 73.910 96.315 74.450 96.485 ;
        RECT 74.730 96.315 74.900 97.055 ;
        RECT 75.165 96.315 75.525 96.690 ;
        RECT 73.910 95.615 74.080 96.315 ;
        RECT 74.250 95.815 74.580 96.145 ;
        RECT 74.750 95.815 75.100 96.145 ;
        RECT 73.910 95.445 74.535 95.615 ;
        RECT 74.750 95.275 75.015 95.815 ;
        RECT 75.270 95.660 75.525 96.315 ;
        RECT 75.695 96.285 79.205 97.055 ;
        RECT 79.835 96.330 80.125 97.055 ;
        RECT 75.695 95.765 77.345 96.285 ;
        RECT 73.035 95.105 75.015 95.275 ;
        RECT 73.035 94.675 73.360 95.105 ;
        RECT 73.530 94.505 73.860 94.925 ;
        RECT 74.605 94.505 75.015 94.935 ;
        RECT 75.185 94.675 75.525 95.660 ;
        RECT 77.515 95.595 79.205 96.115 ;
        RECT 75.695 94.505 79.205 95.595 ;
        RECT 79.835 94.505 80.125 95.670 ;
        RECT 80.300 95.455 80.635 96.875 ;
        RECT 80.815 96.685 81.560 97.055 ;
        RECT 82.125 96.515 82.380 96.875 ;
        RECT 82.560 96.685 82.890 97.055 ;
        RECT 83.070 96.515 83.295 96.875 ;
        RECT 80.810 96.325 83.295 96.515 ;
        RECT 80.810 95.635 81.035 96.325 ;
        RECT 81.235 95.815 81.515 96.145 ;
        RECT 81.695 95.815 82.270 96.145 ;
        RECT 82.450 95.815 82.885 96.145 ;
        RECT 83.065 95.815 83.335 96.145 ;
        RECT 80.810 95.455 83.305 95.635 ;
        RECT 80.300 94.685 80.565 95.455 ;
        RECT 80.735 94.505 81.065 95.225 ;
        RECT 81.255 95.045 82.445 95.275 ;
        RECT 81.255 94.685 81.515 95.045 ;
        RECT 81.685 94.505 82.015 94.875 ;
        RECT 82.185 94.685 82.445 95.045 ;
        RECT 83.015 94.685 83.305 95.455 ;
        RECT 83.525 94.685 83.785 96.875 ;
        RECT 84.045 96.685 84.715 97.055 ;
        RECT 84.895 96.505 85.205 96.875 ;
        RECT 83.975 96.305 85.205 96.505 ;
        RECT 83.975 95.635 84.265 96.305 ;
        RECT 85.385 96.125 85.615 96.765 ;
        RECT 85.795 96.325 86.085 97.055 ;
        RECT 86.275 96.285 87.945 97.055 ;
        RECT 84.445 95.815 84.910 96.125 ;
        RECT 85.090 95.815 85.615 96.125 ;
        RECT 85.795 95.815 86.095 96.145 ;
        RECT 86.275 95.765 87.025 96.285 ;
        RECT 88.125 96.245 88.395 97.055 ;
        RECT 88.565 96.245 88.895 96.885 ;
        RECT 89.065 96.245 89.305 97.055 ;
        RECT 89.495 96.510 94.840 97.055 ;
        RECT 83.975 95.415 84.745 95.635 ;
        RECT 83.955 94.505 84.295 95.235 ;
        RECT 84.475 94.685 84.745 95.415 ;
        RECT 84.925 95.395 86.085 95.635 ;
        RECT 87.195 95.595 87.945 96.115 ;
        RECT 88.115 95.815 88.465 96.065 ;
        RECT 88.635 95.645 88.805 96.245 ;
        RECT 88.975 95.815 89.325 96.065 ;
        RECT 91.080 95.680 91.420 96.510 ;
        RECT 95.015 96.285 98.525 97.055 ;
        RECT 98.695 96.305 99.905 97.055 ;
        RECT 84.925 94.685 85.155 95.395 ;
        RECT 85.325 94.505 85.655 95.215 ;
        RECT 85.825 94.685 86.085 95.395 ;
        RECT 86.275 94.505 87.945 95.595 ;
        RECT 88.125 94.505 88.455 95.645 ;
        RECT 88.635 95.475 89.315 95.645 ;
        RECT 88.985 94.690 89.315 95.475 ;
        RECT 92.900 94.940 93.250 96.190 ;
        RECT 95.015 95.765 96.665 96.285 ;
        RECT 96.835 95.595 98.525 96.115 ;
        RECT 98.695 95.765 99.215 96.305 ;
        RECT 100.135 96.235 100.345 97.055 ;
        RECT 100.515 96.255 100.845 96.885 ;
        RECT 99.385 95.595 99.905 96.135 ;
        RECT 100.515 95.655 100.765 96.255 ;
        RECT 101.015 96.235 101.245 97.055 ;
        RECT 101.455 96.285 104.965 97.055 ;
        RECT 105.595 96.330 105.885 97.055 ;
        RECT 106.075 96.325 106.365 97.055 ;
        RECT 100.935 95.815 101.265 96.065 ;
        RECT 101.455 95.765 103.105 96.285 ;
        RECT 89.495 94.505 94.840 94.940 ;
        RECT 95.015 94.505 98.525 95.595 ;
        RECT 98.695 94.505 99.905 95.595 ;
        RECT 100.135 94.505 100.345 95.645 ;
        RECT 100.515 94.675 100.845 95.655 ;
        RECT 101.015 94.505 101.245 95.645 ;
        RECT 103.275 95.595 104.965 96.115 ;
        RECT 106.065 95.815 106.365 96.145 ;
        RECT 106.545 96.125 106.775 96.765 ;
        RECT 106.955 96.505 107.265 96.875 ;
        RECT 107.445 96.685 108.115 97.055 ;
        RECT 106.955 96.305 108.185 96.505 ;
        RECT 106.545 95.815 107.070 96.125 ;
        RECT 107.250 95.815 107.715 96.125 ;
        RECT 101.455 94.505 104.965 95.595 ;
        RECT 105.595 94.505 105.885 95.670 ;
        RECT 107.895 95.635 108.185 96.305 ;
        RECT 106.075 95.395 107.235 95.635 ;
        RECT 106.075 94.685 106.335 95.395 ;
        RECT 106.505 94.505 106.835 95.215 ;
        RECT 107.005 94.685 107.235 95.395 ;
        RECT 107.415 95.415 108.185 95.635 ;
        RECT 107.415 94.685 107.685 95.415 ;
        RECT 107.865 94.505 108.205 95.235 ;
        RECT 108.375 94.685 108.635 96.875 ;
        RECT 108.815 96.595 109.375 96.885 ;
        RECT 109.545 96.595 109.795 97.055 ;
        RECT 108.815 95.225 109.065 96.595 ;
        RECT 110.415 96.425 110.745 96.785 ;
        RECT 111.115 96.510 116.460 97.055 ;
        RECT 109.355 96.235 110.745 96.425 ;
        RECT 109.355 96.145 109.525 96.235 ;
        RECT 109.235 95.815 109.525 96.145 ;
        RECT 109.695 95.815 110.035 96.065 ;
        RECT 110.255 95.815 110.930 96.065 ;
        RECT 109.355 95.565 109.525 95.815 ;
        RECT 109.355 95.395 110.295 95.565 ;
        RECT 110.665 95.455 110.930 95.815 ;
        RECT 112.700 95.680 113.040 96.510 ;
        RECT 117.555 96.380 117.815 96.885 ;
        RECT 117.995 96.675 118.325 97.055 ;
        RECT 118.505 96.505 118.675 96.885 ;
        RECT 108.815 94.675 109.275 95.225 ;
        RECT 109.465 94.505 109.795 95.225 ;
        RECT 109.995 94.845 110.295 95.395 ;
        RECT 110.465 94.505 110.745 95.175 ;
        RECT 114.520 94.940 114.870 96.190 ;
        RECT 117.555 95.580 117.735 96.380 ;
        RECT 118.010 96.335 118.675 96.505 ;
        RECT 119.025 96.505 119.195 96.885 ;
        RECT 119.375 96.675 119.705 97.055 ;
        RECT 119.025 96.335 119.690 96.505 ;
        RECT 119.885 96.380 120.145 96.885 ;
        RECT 118.010 96.080 118.180 96.335 ;
        RECT 117.905 95.750 118.180 96.080 ;
        RECT 118.405 95.785 118.745 96.155 ;
        RECT 118.955 95.785 119.295 96.155 ;
        RECT 119.520 96.080 119.690 96.335 ;
        RECT 118.010 95.605 118.180 95.750 ;
        RECT 119.520 95.750 119.795 96.080 ;
        RECT 119.520 95.605 119.690 95.750 ;
        RECT 111.115 94.505 116.460 94.940 ;
        RECT 117.555 94.675 117.825 95.580 ;
        RECT 118.010 95.435 118.685 95.605 ;
        RECT 117.995 94.505 118.325 95.265 ;
        RECT 118.505 94.675 118.685 95.435 ;
        RECT 119.015 95.435 119.690 95.605 ;
        RECT 119.965 95.580 120.145 96.380 ;
        RECT 120.320 96.215 120.580 97.055 ;
        RECT 120.755 96.310 121.010 96.885 ;
        RECT 121.180 96.675 121.510 97.055 ;
        RECT 121.725 96.505 121.895 96.885 ;
        RECT 121.180 96.335 121.895 96.505 ;
        RECT 122.245 96.505 122.415 96.885 ;
        RECT 122.630 96.675 122.960 97.055 ;
        RECT 122.245 96.335 122.960 96.505 ;
        RECT 119.015 94.675 119.195 95.435 ;
        RECT 119.375 94.505 119.705 95.265 ;
        RECT 119.875 94.675 120.145 95.580 ;
        RECT 120.320 94.505 120.580 95.655 ;
        RECT 120.755 95.580 120.925 96.310 ;
        RECT 121.180 96.145 121.350 96.335 ;
        RECT 121.095 95.815 121.350 96.145 ;
        RECT 121.180 95.605 121.350 95.815 ;
        RECT 121.630 95.785 121.985 96.155 ;
        RECT 122.155 95.785 122.510 96.155 ;
        RECT 122.790 96.145 122.960 96.335 ;
        RECT 123.130 96.310 123.385 96.885 ;
        RECT 122.790 95.815 123.045 96.145 ;
        RECT 122.790 95.605 122.960 95.815 ;
        RECT 120.755 94.675 121.010 95.580 ;
        RECT 121.180 95.435 121.895 95.605 ;
        RECT 121.180 94.505 121.510 95.265 ;
        RECT 121.725 94.675 121.895 95.435 ;
        RECT 122.245 95.435 122.960 95.605 ;
        RECT 123.215 95.580 123.385 96.310 ;
        RECT 123.560 96.215 123.820 97.055 ;
        RECT 123.995 96.305 125.205 97.055 ;
        RECT 122.245 94.675 122.415 95.435 ;
        RECT 122.630 94.505 122.960 95.265 ;
        RECT 123.130 94.675 123.385 95.580 ;
        RECT 123.560 94.505 123.820 95.655 ;
        RECT 123.995 95.595 124.515 96.135 ;
        RECT 124.685 95.765 125.205 96.305 ;
        RECT 123.995 94.505 125.205 95.595 ;
        RECT 53.990 94.335 125.290 94.505 ;
        RECT 54.075 93.245 55.285 94.335 ;
        RECT 54.075 92.535 54.595 93.075 ;
        RECT 54.765 92.705 55.285 93.245 ;
        RECT 55.455 93.195 55.745 94.335 ;
        RECT 55.915 93.615 56.365 94.165 ;
        RECT 56.555 93.615 56.885 94.335 ;
        RECT 54.075 91.785 55.285 92.535 ;
        RECT 55.455 91.785 55.745 92.585 ;
        RECT 55.915 92.245 56.165 93.615 ;
        RECT 57.095 93.445 57.395 93.995 ;
        RECT 57.565 93.665 57.845 94.335 ;
        RECT 58.305 93.715 58.475 94.145 ;
        RECT 58.645 93.885 58.975 94.335 ;
        RECT 58.305 93.485 58.980 93.715 ;
        RECT 56.455 93.275 57.395 93.445 ;
        RECT 56.455 93.025 56.625 93.275 ;
        RECT 57.730 93.025 58.045 93.465 ;
        RECT 56.335 92.695 56.625 93.025 ;
        RECT 56.795 92.775 57.125 93.025 ;
        RECT 57.355 92.775 58.045 93.025 ;
        RECT 56.455 92.605 56.625 92.695 ;
        RECT 56.455 92.415 57.845 92.605 ;
        RECT 58.275 92.465 58.575 93.315 ;
        RECT 58.745 92.835 58.980 93.485 ;
        RECT 59.150 93.175 59.435 94.120 ;
        RECT 59.615 93.865 60.300 94.335 ;
        RECT 59.610 93.345 60.305 93.655 ;
        RECT 60.480 93.280 60.785 94.065 ;
        RECT 59.150 93.025 60.010 93.175 ;
        RECT 59.150 93.005 60.435 93.025 ;
        RECT 58.745 92.505 59.280 92.835 ;
        RECT 59.450 92.645 60.435 93.005 ;
        RECT 55.915 91.955 56.465 92.245 ;
        RECT 56.635 91.785 56.885 92.245 ;
        RECT 57.515 92.055 57.845 92.415 ;
        RECT 58.745 92.355 58.965 92.505 ;
        RECT 58.220 91.785 58.555 92.290 ;
        RECT 58.725 91.980 58.965 92.355 ;
        RECT 59.450 92.310 59.620 92.645 ;
        RECT 60.610 92.475 60.785 93.280 ;
        RECT 60.975 93.245 62.645 94.335 ;
        RECT 63.275 93.825 63.535 94.335 ;
        RECT 59.245 92.115 59.620 92.310 ;
        RECT 59.245 91.970 59.415 92.115 ;
        RECT 59.980 91.785 60.375 92.280 ;
        RECT 60.545 91.955 60.785 92.475 ;
        RECT 60.975 92.555 61.725 93.075 ;
        RECT 61.895 92.725 62.645 93.245 ;
        RECT 63.275 92.775 63.615 93.655 ;
        RECT 63.785 92.945 63.955 94.165 ;
        RECT 64.195 93.830 64.810 94.335 ;
        RECT 64.195 93.295 64.445 93.660 ;
        RECT 64.615 93.655 64.810 93.830 ;
        RECT 64.980 93.825 65.455 94.165 ;
        RECT 65.625 93.790 65.840 94.335 ;
        RECT 64.615 93.465 64.945 93.655 ;
        RECT 65.165 93.295 65.880 93.590 ;
        RECT 66.050 93.465 66.325 94.165 ;
        RECT 64.195 93.125 65.985 93.295 ;
        RECT 63.785 92.695 64.580 92.945 ;
        RECT 63.785 92.605 64.035 92.695 ;
        RECT 60.975 91.785 62.645 92.555 ;
        RECT 63.275 91.785 63.535 92.605 ;
        RECT 63.705 92.185 64.035 92.605 ;
        RECT 64.750 92.270 65.005 93.125 ;
        RECT 64.215 92.005 65.005 92.270 ;
        RECT 65.175 92.425 65.585 92.945 ;
        RECT 65.755 92.695 65.985 93.125 ;
        RECT 66.155 92.435 66.325 93.465 ;
        RECT 66.955 93.170 67.245 94.335 ;
        RECT 67.415 93.825 67.675 94.335 ;
        RECT 67.415 92.775 67.755 93.655 ;
        RECT 67.925 92.945 68.095 94.165 ;
        RECT 68.335 93.830 68.950 94.335 ;
        RECT 68.335 93.295 68.585 93.660 ;
        RECT 68.755 93.655 68.950 93.830 ;
        RECT 69.120 93.825 69.595 94.165 ;
        RECT 69.765 93.790 69.980 94.335 ;
        RECT 68.755 93.465 69.085 93.655 ;
        RECT 69.305 93.295 70.020 93.590 ;
        RECT 70.190 93.465 70.465 94.165 ;
        RECT 68.335 93.125 70.125 93.295 ;
        RECT 67.925 92.695 68.720 92.945 ;
        RECT 67.925 92.605 68.175 92.695 ;
        RECT 65.175 92.005 65.375 92.425 ;
        RECT 65.565 91.785 65.895 92.245 ;
        RECT 66.065 91.955 66.325 92.435 ;
        RECT 66.955 91.785 67.245 92.510 ;
        RECT 67.415 91.785 67.675 92.605 ;
        RECT 67.845 92.185 68.175 92.605 ;
        RECT 68.890 92.270 69.145 93.125 ;
        RECT 68.355 92.005 69.145 92.270 ;
        RECT 69.315 92.425 69.725 92.945 ;
        RECT 69.895 92.695 70.125 93.125 ;
        RECT 70.295 92.435 70.465 93.465 ;
        RECT 71.620 93.365 71.890 94.160 ;
        RECT 72.070 93.535 72.285 94.335 ;
        RECT 72.465 93.365 72.750 94.160 ;
        RECT 71.620 93.195 72.750 93.365 ;
        RECT 71.600 92.725 72.100 92.990 ;
        RECT 72.320 92.695 72.705 93.025 ;
        RECT 72.930 92.695 73.210 94.165 ;
        RECT 73.390 92.750 73.720 94.165 ;
        RECT 73.890 92.990 74.095 94.165 ;
        RECT 74.265 93.345 74.475 94.160 ;
        RECT 74.715 93.515 75.045 94.335 ;
        RECT 74.265 93.165 74.915 93.345 ;
        RECT 75.220 93.320 75.475 94.160 ;
        RECT 75.700 93.910 76.035 94.335 ;
        RECT 76.205 93.730 76.390 94.135 ;
        RECT 73.890 92.750 74.320 92.990 ;
        RECT 72.320 92.545 72.625 92.695 ;
        RECT 69.315 92.005 69.515 92.425 ;
        RECT 69.705 91.785 70.035 92.245 ;
        RECT 70.205 91.955 70.465 92.435 ;
        RECT 71.655 91.785 71.895 92.460 ;
        RECT 72.070 91.985 72.625 92.545 ;
        RECT 74.695 92.525 74.915 93.165 ;
        RECT 72.805 92.355 74.915 92.525 ;
        RECT 72.805 91.960 73.010 92.355 ;
        RECT 73.695 92.350 74.915 92.355 ;
        RECT 73.180 91.785 73.525 92.185 ;
        RECT 73.695 91.960 74.025 92.350 ;
        RECT 74.300 91.785 74.975 92.170 ;
        RECT 75.145 91.955 75.475 93.320 ;
        RECT 75.725 93.555 76.390 93.730 ;
        RECT 76.595 93.555 76.925 94.335 ;
        RECT 75.725 92.525 76.065 93.555 ;
        RECT 77.095 93.365 77.365 94.135 ;
        RECT 76.235 93.195 77.365 93.365 ;
        RECT 77.545 93.195 77.875 94.335 ;
        RECT 78.405 93.365 78.735 94.150 ;
        RECT 79.575 93.665 79.855 94.335 ;
        RECT 80.025 93.445 80.325 93.995 ;
        RECT 80.525 93.615 80.855 94.335 ;
        RECT 81.045 93.615 81.505 94.165 ;
        RECT 78.055 93.195 78.735 93.365 ;
        RECT 76.235 92.695 76.485 93.195 ;
        RECT 75.725 92.355 76.410 92.525 ;
        RECT 76.665 92.445 77.025 93.025 ;
        RECT 75.700 91.785 76.035 92.185 ;
        RECT 76.205 91.955 76.410 92.355 ;
        RECT 77.195 92.285 77.365 93.195 ;
        RECT 77.535 92.775 77.885 93.025 ;
        RECT 78.055 92.595 78.225 93.195 ;
        RECT 79.390 93.025 79.655 93.385 ;
        RECT 80.025 93.275 80.965 93.445 ;
        RECT 80.795 93.025 80.965 93.275 ;
        RECT 78.395 92.775 78.745 93.025 ;
        RECT 79.390 92.775 80.065 93.025 ;
        RECT 80.285 92.775 80.625 93.025 ;
        RECT 80.795 92.695 81.085 93.025 ;
        RECT 80.795 92.605 80.965 92.695 ;
        RECT 76.620 91.785 76.895 92.265 ;
        RECT 77.105 91.955 77.365 92.285 ;
        RECT 77.545 91.785 77.815 92.595 ;
        RECT 77.985 91.955 78.315 92.595 ;
        RECT 78.485 91.785 78.725 92.595 ;
        RECT 79.575 92.415 80.965 92.605 ;
        RECT 79.575 92.055 79.905 92.415 ;
        RECT 81.255 92.245 81.505 93.615 ;
        RECT 82.170 93.535 82.420 94.335 ;
        RECT 82.590 93.705 82.920 94.165 ;
        RECT 83.090 93.875 83.305 94.335 ;
        RECT 82.590 93.535 83.760 93.705 ;
        RECT 81.680 93.365 81.960 93.525 ;
        RECT 81.680 93.195 83.015 93.365 ;
        RECT 82.845 93.025 83.015 93.195 ;
        RECT 81.680 92.775 82.030 93.015 ;
        RECT 82.200 92.775 82.675 93.015 ;
        RECT 82.845 92.775 83.220 93.025 ;
        RECT 82.845 92.605 83.015 92.775 ;
        RECT 80.525 91.785 80.775 92.245 ;
        RECT 80.945 91.955 81.505 92.245 ;
        RECT 81.680 92.435 83.015 92.605 ;
        RECT 81.680 92.225 81.950 92.435 ;
        RECT 83.390 92.245 83.760 93.535 ;
        RECT 83.975 93.245 85.645 94.335 ;
        RECT 82.170 91.785 82.500 92.245 ;
        RECT 83.010 91.955 83.760 92.245 ;
        RECT 83.975 92.555 84.725 93.075 ;
        RECT 84.895 92.725 85.645 93.245 ;
        RECT 86.275 93.485 86.615 94.125 ;
        RECT 86.785 93.875 87.030 94.335 ;
        RECT 87.205 93.705 87.455 94.165 ;
        RECT 87.645 93.955 88.315 94.335 ;
        RECT 88.515 93.705 88.765 94.165 ;
        RECT 87.205 93.535 88.765 93.705 ;
        RECT 83.975 91.785 85.645 92.555 ;
        RECT 86.275 92.370 86.445 93.485 ;
        RECT 89.525 93.365 89.695 94.165 ;
        RECT 86.755 93.195 89.695 93.365 ;
        RECT 90.045 93.405 90.215 94.165 ;
        RECT 90.430 93.575 90.760 94.335 ;
        RECT 90.045 93.235 90.760 93.405 ;
        RECT 90.930 93.260 91.185 94.165 ;
        RECT 86.755 93.025 86.925 93.195 ;
        RECT 86.615 92.695 86.925 93.025 ;
        RECT 87.095 92.695 87.430 93.025 ;
        RECT 86.755 92.525 86.925 92.695 ;
        RECT 86.275 91.955 86.585 92.370 ;
        RECT 86.755 92.355 87.450 92.525 ;
        RECT 87.700 92.450 87.895 93.025 ;
        RECT 88.155 92.695 88.500 93.025 ;
        RECT 88.810 92.695 89.285 93.025 ;
        RECT 89.540 92.695 89.725 93.025 ;
        RECT 88.155 92.465 88.345 92.695 ;
        RECT 89.955 92.685 90.310 93.055 ;
        RECT 90.590 93.025 90.760 93.235 ;
        RECT 90.590 92.695 90.845 93.025 ;
        RECT 86.780 91.785 87.110 92.165 ;
        RECT 87.280 92.125 87.450 92.355 ;
        RECT 88.515 92.355 89.695 92.525 ;
        RECT 90.590 92.505 90.760 92.695 ;
        RECT 91.015 92.530 91.185 93.260 ;
        RECT 91.360 93.185 91.620 94.335 ;
        RECT 92.715 93.170 93.005 94.335 ;
        RECT 88.515 92.125 88.685 92.355 ;
        RECT 87.280 91.955 88.685 92.125 ;
        RECT 88.955 91.785 89.285 92.185 ;
        RECT 89.525 91.955 89.695 92.355 ;
        RECT 90.045 92.335 90.760 92.505 ;
        RECT 90.045 91.955 90.215 92.335 ;
        RECT 90.430 91.785 90.760 92.165 ;
        RECT 90.930 91.955 91.185 92.530 ;
        RECT 91.360 91.785 91.620 92.625 ;
        RECT 92.715 91.785 93.005 92.510 ;
        RECT 93.175 92.065 93.455 94.165 ;
        RECT 93.645 93.575 94.430 94.335 ;
        RECT 94.825 93.505 95.210 94.165 ;
        RECT 94.825 93.405 95.235 93.505 ;
        RECT 93.625 93.195 95.235 93.405 ;
        RECT 95.535 93.315 95.735 94.105 ;
        RECT 93.625 92.595 93.900 93.195 ;
        RECT 95.405 93.145 95.735 93.315 ;
        RECT 95.905 93.155 96.225 94.335 ;
        RECT 96.395 93.735 96.655 94.155 ;
        RECT 96.825 93.905 97.155 94.335 ;
        RECT 97.845 93.905 98.590 94.075 ;
        RECT 96.395 93.565 98.250 93.735 ;
        RECT 95.405 93.025 95.585 93.145 ;
        RECT 94.070 92.775 94.425 93.025 ;
        RECT 94.620 92.975 95.085 93.025 ;
        RECT 94.615 92.805 95.085 92.975 ;
        RECT 94.620 92.775 95.085 92.805 ;
        RECT 95.255 92.775 95.585 93.025 ;
        RECT 95.760 92.775 96.225 92.975 ;
        RECT 93.625 92.415 94.875 92.595 ;
        RECT 94.510 92.345 94.875 92.415 ;
        RECT 95.045 92.395 96.225 92.565 ;
        RECT 93.685 91.785 93.855 92.245 ;
        RECT 95.045 92.175 95.375 92.395 ;
        RECT 94.125 91.995 95.375 92.175 ;
        RECT 95.545 91.785 95.715 92.225 ;
        RECT 95.885 91.980 96.225 92.395 ;
        RECT 96.395 92.525 96.570 93.565 ;
        RECT 96.740 92.695 97.090 93.395 ;
        RECT 97.305 93.225 97.910 93.395 ;
        RECT 97.260 92.695 97.550 93.025 ;
        RECT 97.720 92.945 97.910 93.225 ;
        RECT 98.080 93.285 98.250 93.565 ;
        RECT 98.420 93.655 98.590 93.905 ;
        RECT 98.815 93.825 99.455 94.155 ;
        RECT 98.420 93.485 99.455 93.655 ;
        RECT 99.625 93.535 99.905 94.335 ;
        RECT 99.285 93.365 99.455 93.485 ;
        RECT 98.080 93.115 98.730 93.285 ;
        RECT 99.285 93.195 99.945 93.365 ;
        RECT 100.115 93.195 100.390 94.165 ;
        RECT 97.720 92.775 98.165 92.945 ;
        RECT 97.720 92.525 97.910 92.775 ;
        RECT 98.560 92.695 98.730 93.115 ;
        RECT 99.775 93.025 99.945 93.195 ;
        RECT 98.950 92.695 99.605 93.025 ;
        RECT 99.775 92.695 100.050 93.025 ;
        RECT 99.775 92.525 99.945 92.695 ;
        RECT 96.395 92.150 96.715 92.525 ;
        RECT 96.970 91.785 97.140 92.525 ;
        RECT 97.390 92.355 97.910 92.525 ;
        RECT 98.335 92.355 99.945 92.525 ;
        RECT 100.220 92.460 100.390 93.195 ;
        RECT 100.560 93.140 100.730 94.335 ;
        RECT 100.995 93.195 101.255 94.335 ;
        RECT 101.425 93.185 101.755 94.165 ;
        RECT 101.925 93.195 102.205 94.335 ;
        RECT 102.375 93.245 103.585 94.335 ;
        RECT 101.015 92.775 101.350 93.025 ;
        RECT 97.390 92.150 97.560 92.355 ;
        RECT 97.805 91.785 98.160 92.185 ;
        RECT 98.335 92.005 98.505 92.355 ;
        RECT 98.705 91.785 99.035 92.185 ;
        RECT 99.205 92.005 99.375 92.355 ;
        RECT 99.545 91.785 99.925 92.185 ;
        RECT 100.115 92.115 100.390 92.460 ;
        RECT 100.560 91.785 100.730 92.725 ;
        RECT 101.520 92.585 101.690 93.185 ;
        RECT 101.860 92.755 102.195 93.025 ;
        RECT 100.995 91.955 101.690 92.585 ;
        RECT 101.895 91.785 102.205 92.585 ;
        RECT 102.375 92.535 102.895 93.075 ;
        RECT 103.065 92.705 103.585 93.245 ;
        RECT 103.775 93.445 104.035 94.155 ;
        RECT 104.205 93.625 104.535 94.335 ;
        RECT 104.705 93.445 104.935 94.155 ;
        RECT 103.775 93.205 104.935 93.445 ;
        RECT 105.115 93.425 105.385 94.155 ;
        RECT 105.565 93.605 105.905 94.335 ;
        RECT 105.115 93.205 105.885 93.425 ;
        RECT 103.765 92.695 104.065 93.025 ;
        RECT 104.245 92.715 104.770 93.025 ;
        RECT 104.950 92.715 105.415 93.025 ;
        RECT 102.375 91.785 103.585 92.535 ;
        RECT 103.775 91.785 104.065 92.515 ;
        RECT 104.245 92.075 104.475 92.715 ;
        RECT 105.595 92.535 105.885 93.205 ;
        RECT 104.655 92.335 105.885 92.535 ;
        RECT 104.655 91.965 104.965 92.335 ;
        RECT 105.145 91.785 105.815 92.155 ;
        RECT 106.075 91.965 106.335 94.155 ;
        RECT 106.525 93.725 106.855 94.155 ;
        RECT 107.035 93.895 107.230 94.335 ;
        RECT 107.400 93.725 107.730 94.155 ;
        RECT 106.525 93.555 107.730 93.725 ;
        RECT 106.525 93.225 107.420 93.555 ;
        RECT 107.900 93.385 108.175 94.155 ;
        RECT 108.355 93.900 113.700 94.335 ;
        RECT 107.590 93.195 108.175 93.385 ;
        RECT 106.530 92.695 106.825 93.025 ;
        RECT 107.005 92.695 107.420 93.025 ;
        RECT 106.525 91.785 106.825 92.515 ;
        RECT 107.005 92.075 107.235 92.695 ;
        RECT 107.590 92.525 107.765 93.195 ;
        RECT 107.435 92.345 107.765 92.525 ;
        RECT 107.935 92.375 108.175 93.025 ;
        RECT 107.435 91.965 107.660 92.345 ;
        RECT 109.940 92.330 110.280 93.160 ;
        RECT 111.760 92.650 112.110 93.900 ;
        RECT 113.875 93.245 117.385 94.335 ;
        RECT 113.875 92.555 115.525 93.075 ;
        RECT 115.695 92.725 117.385 93.245 ;
        RECT 118.475 93.170 118.765 94.335 ;
        RECT 118.935 93.245 120.605 94.335 ;
        RECT 118.935 92.555 119.685 93.075 ;
        RECT 119.855 92.725 120.605 93.245 ;
        RECT 120.855 93.405 121.035 94.165 ;
        RECT 121.215 93.575 121.545 94.335 ;
        RECT 120.855 93.235 121.530 93.405 ;
        RECT 121.715 93.260 121.985 94.165 ;
        RECT 121.360 93.090 121.530 93.235 ;
        RECT 120.795 92.685 121.135 93.055 ;
        RECT 121.360 92.760 121.635 93.090 ;
        RECT 107.830 91.785 108.160 92.175 ;
        RECT 108.355 91.785 113.700 92.330 ;
        RECT 113.875 91.785 117.385 92.555 ;
        RECT 118.475 91.785 118.765 92.510 ;
        RECT 118.935 91.785 120.605 92.555 ;
        RECT 121.360 92.505 121.530 92.760 ;
        RECT 120.865 92.335 121.530 92.505 ;
        RECT 121.805 92.460 121.985 93.260 ;
        RECT 120.865 91.955 121.035 92.335 ;
        RECT 121.215 91.785 121.545 92.165 ;
        RECT 121.725 91.955 121.985 92.460 ;
        RECT 122.155 93.365 122.425 94.135 ;
        RECT 122.595 93.555 122.925 94.335 ;
        RECT 123.130 93.730 123.315 94.135 ;
        RECT 123.485 93.910 123.820 94.335 ;
        RECT 123.130 93.555 123.795 93.730 ;
        RECT 122.155 93.195 123.285 93.365 ;
        RECT 122.155 92.285 122.325 93.195 ;
        RECT 122.495 92.445 122.855 93.025 ;
        RECT 123.035 92.695 123.285 93.195 ;
        RECT 123.455 92.525 123.795 93.555 ;
        RECT 123.995 93.245 125.205 94.335 ;
        RECT 123.995 92.705 124.515 93.245 ;
        RECT 124.685 92.535 125.205 93.075 ;
        RECT 123.110 92.355 123.795 92.525 ;
        RECT 122.155 91.955 122.415 92.285 ;
        RECT 122.625 91.785 122.900 92.265 ;
        RECT 123.110 91.955 123.315 92.355 ;
        RECT 123.485 91.785 123.820 92.185 ;
        RECT 123.995 91.785 125.205 92.535 ;
        RECT 53.990 91.615 125.290 91.785 ;
        RECT 54.075 90.865 55.285 91.615 ;
        RECT 54.075 90.325 54.595 90.865 ;
        RECT 55.460 90.775 55.720 91.615 ;
        RECT 55.895 90.870 56.150 91.445 ;
        RECT 56.320 91.235 56.650 91.615 ;
        RECT 56.865 91.065 57.035 91.445 ;
        RECT 56.320 90.895 57.035 91.065 ;
        RECT 54.765 90.155 55.285 90.695 ;
        RECT 54.075 89.065 55.285 90.155 ;
        RECT 55.460 89.065 55.720 90.215 ;
        RECT 55.895 90.140 56.065 90.870 ;
        RECT 56.320 90.705 56.490 90.895 ;
        RECT 57.335 90.795 57.565 91.615 ;
        RECT 57.735 90.815 58.065 91.445 ;
        RECT 56.235 90.375 56.490 90.705 ;
        RECT 56.320 90.165 56.490 90.375 ;
        RECT 56.770 90.345 57.125 90.715 ;
        RECT 57.315 90.375 57.645 90.625 ;
        RECT 57.815 90.215 58.065 90.815 ;
        RECT 58.235 90.795 58.445 91.615 ;
        RECT 58.675 90.940 58.935 91.445 ;
        RECT 59.115 91.235 59.445 91.615 ;
        RECT 59.625 91.065 59.795 91.445 ;
        RECT 60.055 91.070 65.400 91.615 ;
        RECT 65.575 91.070 70.920 91.615 ;
        RECT 71.120 91.225 71.450 91.615 ;
        RECT 55.895 89.235 56.150 90.140 ;
        RECT 56.320 89.995 57.035 90.165 ;
        RECT 56.320 89.065 56.650 89.825 ;
        RECT 56.865 89.235 57.035 89.995 ;
        RECT 57.335 89.065 57.565 90.205 ;
        RECT 57.735 89.235 58.065 90.215 ;
        RECT 58.235 89.065 58.445 90.205 ;
        RECT 58.675 90.140 58.845 90.940 ;
        RECT 59.130 90.895 59.795 91.065 ;
        RECT 59.130 90.640 59.300 90.895 ;
        RECT 59.015 90.310 59.300 90.640 ;
        RECT 59.535 90.345 59.865 90.715 ;
        RECT 59.130 90.165 59.300 90.310 ;
        RECT 61.640 90.240 61.980 91.070 ;
        RECT 58.675 89.235 58.945 90.140 ;
        RECT 59.130 89.995 59.795 90.165 ;
        RECT 59.115 89.065 59.445 89.825 ;
        RECT 59.625 89.235 59.795 89.995 ;
        RECT 63.460 89.500 63.810 90.750 ;
        RECT 67.160 90.240 67.500 91.070 ;
        RECT 71.620 91.055 71.845 91.435 ;
        RECT 68.980 89.500 69.330 90.750 ;
        RECT 71.105 90.375 71.345 91.025 ;
        RECT 71.515 90.875 71.845 91.055 ;
        RECT 71.515 90.205 71.690 90.875 ;
        RECT 72.045 90.705 72.275 91.325 ;
        RECT 72.455 90.885 72.755 91.615 ;
        RECT 73.025 91.065 73.195 91.445 ;
        RECT 73.410 91.235 73.740 91.615 ;
        RECT 73.025 90.895 73.740 91.065 ;
        RECT 71.860 90.375 72.275 90.705 ;
        RECT 72.455 90.375 72.750 90.705 ;
        RECT 72.935 90.345 73.290 90.715 ;
        RECT 73.570 90.705 73.740 90.895 ;
        RECT 73.910 90.870 74.165 91.445 ;
        RECT 73.570 90.375 73.825 90.705 ;
        RECT 71.105 90.015 71.690 90.205 ;
        RECT 60.055 89.065 65.400 89.500 ;
        RECT 65.575 89.065 70.920 89.500 ;
        RECT 71.105 89.245 71.380 90.015 ;
        RECT 71.860 89.845 72.755 90.175 ;
        RECT 73.570 90.165 73.740 90.375 ;
        RECT 71.550 89.675 72.755 89.845 ;
        RECT 71.550 89.245 71.880 89.675 ;
        RECT 72.050 89.065 72.245 89.505 ;
        RECT 72.425 89.245 72.755 89.675 ;
        RECT 73.025 89.995 73.740 90.165 ;
        RECT 73.995 90.140 74.165 90.870 ;
        RECT 74.340 90.775 74.600 91.615 ;
        RECT 74.775 90.845 78.285 91.615 ;
        RECT 78.455 90.865 79.665 91.615 ;
        RECT 79.835 90.890 80.125 91.615 ;
        RECT 80.295 91.070 85.640 91.615 ;
        RECT 74.775 90.325 76.425 90.845 ;
        RECT 73.025 89.235 73.195 89.995 ;
        RECT 73.410 89.065 73.740 89.825 ;
        RECT 73.910 89.235 74.165 90.140 ;
        RECT 74.340 89.065 74.600 90.215 ;
        RECT 76.595 90.155 78.285 90.675 ;
        RECT 78.455 90.325 78.975 90.865 ;
        RECT 79.145 90.155 79.665 90.695 ;
        RECT 81.880 90.240 82.220 91.070 ;
        RECT 86.275 91.030 86.585 91.445 ;
        RECT 86.780 91.235 87.110 91.615 ;
        RECT 87.280 91.275 88.685 91.445 ;
        RECT 87.280 91.045 87.450 91.275 ;
        RECT 74.775 89.065 78.285 90.155 ;
        RECT 78.455 89.065 79.665 90.155 ;
        RECT 79.835 89.065 80.125 90.230 ;
        RECT 83.700 89.500 84.050 90.750 ;
        RECT 86.275 89.915 86.445 91.030 ;
        RECT 86.755 90.875 87.450 91.045 ;
        RECT 88.515 91.045 88.685 91.275 ;
        RECT 88.955 91.215 89.285 91.615 ;
        RECT 89.525 91.045 89.695 91.445 ;
        RECT 86.755 90.705 86.925 90.875 ;
        RECT 86.615 90.375 86.925 90.705 ;
        RECT 87.095 90.375 87.430 90.705 ;
        RECT 87.700 90.375 87.895 90.950 ;
        RECT 88.155 90.705 88.345 90.935 ;
        RECT 88.515 90.875 89.695 91.045 ;
        RECT 89.990 90.875 90.605 91.445 ;
        RECT 90.775 91.105 90.990 91.615 ;
        RECT 91.220 91.105 91.500 91.435 ;
        RECT 91.680 91.105 91.920 91.615 ;
        RECT 88.155 90.375 88.500 90.705 ;
        RECT 88.810 90.375 89.285 90.705 ;
        RECT 89.540 90.375 89.725 90.705 ;
        RECT 86.755 90.205 86.925 90.375 ;
        RECT 86.755 90.035 89.695 90.205 ;
        RECT 80.295 89.065 85.640 89.500 ;
        RECT 86.275 89.275 86.615 89.915 ;
        RECT 87.205 89.695 88.765 89.865 ;
        RECT 86.785 89.065 87.030 89.525 ;
        RECT 87.205 89.235 87.455 89.695 ;
        RECT 87.645 89.065 88.315 89.445 ;
        RECT 88.515 89.235 88.765 89.695 ;
        RECT 89.525 89.235 89.695 90.035 ;
        RECT 89.990 89.855 90.305 90.875 ;
        RECT 90.475 90.205 90.645 90.705 ;
        RECT 90.895 90.375 91.160 90.935 ;
        RECT 91.330 90.205 91.500 91.105 ;
        RECT 91.670 90.375 92.025 90.935 ;
        RECT 92.275 90.805 92.515 91.615 ;
        RECT 92.685 90.805 93.015 91.445 ;
        RECT 93.185 90.805 93.455 91.615 ;
        RECT 92.255 90.375 92.605 90.625 ;
        RECT 92.775 90.205 92.945 90.805 ;
        RECT 93.115 90.375 93.465 90.625 ;
        RECT 90.475 90.035 91.900 90.205 ;
        RECT 89.990 89.235 90.525 89.855 ;
        RECT 90.695 89.065 91.025 89.865 ;
        RECT 91.510 89.860 91.900 90.035 ;
        RECT 92.265 90.035 92.945 90.205 ;
        RECT 92.265 89.250 92.595 90.035 ;
        RECT 93.125 89.065 93.455 90.205 ;
        RECT 93.635 89.235 93.915 91.335 ;
        RECT 94.145 91.155 94.315 91.615 ;
        RECT 94.585 91.225 95.835 91.405 ;
        RECT 94.970 90.985 95.335 91.055 ;
        RECT 94.085 90.805 95.335 90.985 ;
        RECT 95.505 91.005 95.835 91.225 ;
        RECT 96.005 91.175 96.175 91.615 ;
        RECT 96.345 91.005 96.685 91.420 ;
        RECT 95.505 90.835 96.685 91.005 ;
        RECT 96.855 90.815 97.165 91.615 ;
        RECT 97.370 90.815 98.065 91.445 ;
        RECT 98.235 91.070 103.580 91.615 ;
        RECT 94.085 90.205 94.360 90.805 ;
        RECT 94.530 90.375 94.885 90.625 ;
        RECT 95.080 90.595 95.545 90.625 ;
        RECT 95.075 90.425 95.545 90.595 ;
        RECT 95.080 90.375 95.545 90.425 ;
        RECT 95.715 90.375 96.045 90.625 ;
        RECT 96.220 90.425 96.685 90.625 ;
        RECT 96.865 90.375 97.200 90.645 ;
        RECT 95.865 90.255 96.045 90.375 ;
        RECT 94.085 89.995 95.695 90.205 ;
        RECT 95.865 90.085 96.195 90.255 ;
        RECT 95.285 89.895 95.695 89.995 ;
        RECT 94.105 89.065 94.890 89.825 ;
        RECT 95.285 89.235 95.670 89.895 ;
        RECT 95.995 89.295 96.195 90.085 ;
        RECT 96.365 89.065 96.685 90.245 ;
        RECT 97.370 90.215 97.540 90.815 ;
        RECT 97.710 90.375 98.045 90.625 ;
        RECT 99.820 90.240 100.160 91.070 ;
        RECT 103.765 90.885 104.065 91.615 ;
        RECT 96.855 89.065 97.135 90.205 ;
        RECT 97.305 89.235 97.635 90.215 ;
        RECT 97.805 89.065 98.065 90.205 ;
        RECT 101.640 89.500 101.990 90.750 ;
        RECT 104.245 90.705 104.475 91.325 ;
        RECT 104.675 91.055 104.900 91.435 ;
        RECT 105.070 91.225 105.400 91.615 ;
        RECT 104.675 90.875 105.005 91.055 ;
        RECT 103.770 90.375 104.065 90.705 ;
        RECT 104.245 90.375 104.660 90.705 ;
        RECT 104.830 90.205 105.005 90.875 ;
        RECT 105.175 90.375 105.415 91.025 ;
        RECT 105.595 90.890 105.885 91.615 ;
        RECT 106.055 91.070 111.400 91.615 ;
        RECT 111.575 91.070 116.920 91.615 ;
        RECT 117.095 91.070 122.440 91.615 ;
        RECT 107.640 90.240 107.980 91.070 ;
        RECT 103.765 89.845 104.660 90.175 ;
        RECT 104.830 90.015 105.415 90.205 ;
        RECT 103.765 89.675 104.970 89.845 ;
        RECT 98.235 89.065 103.580 89.500 ;
        RECT 103.765 89.245 104.095 89.675 ;
        RECT 104.275 89.065 104.470 89.505 ;
        RECT 104.640 89.245 104.970 89.675 ;
        RECT 105.140 89.245 105.415 90.015 ;
        RECT 105.595 89.065 105.885 90.230 ;
        RECT 109.460 89.500 109.810 90.750 ;
        RECT 113.160 90.240 113.500 91.070 ;
        RECT 114.980 89.500 115.330 90.750 ;
        RECT 118.680 90.240 119.020 91.070 ;
        RECT 122.615 90.940 122.875 91.445 ;
        RECT 123.055 91.235 123.385 91.615 ;
        RECT 123.565 91.065 123.735 91.445 ;
        RECT 120.500 89.500 120.850 90.750 ;
        RECT 122.615 90.140 122.785 90.940 ;
        RECT 123.070 90.895 123.735 91.065 ;
        RECT 123.070 90.640 123.240 90.895 ;
        RECT 123.995 90.865 125.205 91.615 ;
        RECT 122.955 90.310 123.240 90.640 ;
        RECT 123.475 90.345 123.805 90.715 ;
        RECT 123.070 90.165 123.240 90.310 ;
        RECT 106.055 89.065 111.400 89.500 ;
        RECT 111.575 89.065 116.920 89.500 ;
        RECT 117.095 89.065 122.440 89.500 ;
        RECT 122.615 89.235 122.885 90.140 ;
        RECT 123.070 89.995 123.735 90.165 ;
        RECT 123.055 89.065 123.385 89.825 ;
        RECT 123.565 89.235 123.735 89.995 ;
        RECT 123.995 90.155 124.515 90.695 ;
        RECT 124.685 90.325 125.205 90.865 ;
        RECT 123.995 89.065 125.205 90.155 ;
        RECT 53.990 88.895 125.290 89.065 ;
        RECT 54.075 87.805 55.285 88.895 ;
        RECT 55.455 88.460 60.800 88.895 ;
        RECT 60.975 88.460 66.320 88.895 ;
        RECT 54.075 87.095 54.595 87.635 ;
        RECT 54.765 87.265 55.285 87.805 ;
        RECT 54.075 86.345 55.285 87.095 ;
        RECT 57.040 86.890 57.380 87.720 ;
        RECT 58.860 87.210 59.210 88.460 ;
        RECT 62.560 86.890 62.900 87.720 ;
        RECT 64.380 87.210 64.730 88.460 ;
        RECT 66.955 87.730 67.245 88.895 ;
        RECT 67.415 87.805 69.085 88.895 ;
        RECT 67.415 87.115 68.165 87.635 ;
        RECT 68.335 87.285 69.085 87.805 ;
        RECT 69.715 87.755 69.995 88.895 ;
        RECT 70.165 87.745 70.495 88.725 ;
        RECT 70.665 87.755 70.925 88.895 ;
        RECT 71.100 88.055 71.420 88.895 ;
        RECT 71.590 87.875 71.790 88.665 ;
        RECT 72.115 87.965 72.500 88.725 ;
        RECT 72.895 88.135 73.695 88.895 ;
        RECT 70.230 87.705 70.405 87.745 ;
        RECT 69.725 87.315 70.060 87.585 ;
        RECT 70.230 87.145 70.400 87.705 ;
        RECT 70.570 87.335 70.905 87.585 ;
        RECT 71.100 87.535 71.420 87.875 ;
        RECT 71.590 87.705 71.945 87.875 ;
        RECT 72.115 87.755 73.715 87.965 ;
        RECT 71.765 87.585 71.945 87.705 ;
        RECT 71.100 87.335 71.595 87.535 ;
        RECT 71.765 87.335 72.095 87.585 ;
        RECT 72.265 87.335 72.730 87.585 ;
        RECT 72.900 87.335 73.255 87.585 ;
        RECT 73.435 87.155 73.715 87.755 ;
        RECT 55.455 86.345 60.800 86.890 ;
        RECT 60.975 86.345 66.320 86.890 ;
        RECT 66.955 86.345 67.245 87.070 ;
        RECT 67.415 86.345 69.085 87.115 ;
        RECT 69.715 86.345 70.025 87.145 ;
        RECT 70.230 86.515 70.925 87.145 ;
        RECT 71.100 87.085 72.130 87.125 ;
        RECT 71.100 86.955 72.300 87.085 ;
        RECT 71.100 86.540 71.435 86.955 ;
        RECT 71.605 86.345 71.775 86.785 ;
        RECT 71.960 86.735 72.300 86.955 ;
        RECT 72.475 86.975 73.715 87.155 ;
        RECT 72.475 86.905 72.840 86.975 ;
        RECT 71.960 86.555 73.225 86.735 ;
        RECT 73.485 86.345 73.665 86.805 ;
        RECT 73.885 86.625 74.100 88.725 ;
        RECT 74.325 87.705 74.575 88.895 ;
        RECT 74.775 87.755 75.160 88.715 ;
        RECT 75.375 88.095 75.665 88.895 ;
        RECT 75.835 88.555 77.200 88.725 ;
        RECT 75.835 87.925 76.005 88.555 ;
        RECT 75.330 87.755 76.005 87.925 ;
        RECT 74.335 86.345 74.505 87.145 ;
        RECT 74.775 87.085 74.950 87.755 ;
        RECT 75.330 87.585 75.500 87.755 ;
        RECT 76.175 87.585 76.500 88.385 ;
        RECT 76.870 88.345 77.200 88.555 ;
        RECT 76.870 88.095 77.825 88.345 ;
        RECT 75.135 87.335 75.500 87.585 ;
        RECT 75.695 87.335 75.945 87.585 ;
        RECT 75.135 87.255 75.325 87.335 ;
        RECT 75.695 87.255 75.865 87.335 ;
        RECT 76.155 87.255 76.500 87.585 ;
        RECT 76.670 87.255 76.945 87.920 ;
        RECT 77.130 87.255 77.485 87.920 ;
        RECT 77.655 87.085 77.825 88.095 ;
        RECT 77.995 87.755 78.285 88.895 ;
        RECT 78.455 87.805 81.045 88.895 ;
        RECT 78.010 87.255 78.285 87.585 ;
        RECT 74.775 86.515 75.285 87.085 ;
        RECT 75.830 86.915 77.230 87.085 ;
        RECT 75.455 86.345 75.625 86.905 ;
        RECT 75.830 86.515 76.160 86.915 ;
        RECT 76.335 86.345 76.665 86.745 ;
        RECT 76.900 86.725 77.230 86.915 ;
        RECT 77.400 86.895 77.825 87.085 ;
        RECT 78.455 87.115 79.665 87.635 ;
        RECT 79.835 87.285 81.045 87.805 ;
        RECT 81.215 87.755 81.545 88.895 ;
        RECT 81.715 88.265 82.070 88.725 ;
        RECT 82.240 88.435 82.815 88.895 ;
        RECT 82.985 88.265 83.315 88.725 ;
        RECT 81.715 88.095 83.315 88.265 ;
        RECT 83.515 88.095 83.770 88.895 ;
        RECT 84.435 88.460 89.780 88.895 ;
        RECT 81.715 87.755 81.990 88.095 ;
        RECT 82.170 87.535 82.360 87.915 ;
        RECT 81.215 87.335 82.360 87.535 ;
        RECT 82.540 87.165 82.820 88.095 ;
        RECT 83.940 87.925 84.240 88.120 ;
        RECT 82.990 87.755 84.240 87.925 ;
        RECT 82.990 87.335 83.320 87.755 ;
        RECT 83.550 87.255 83.895 87.585 ;
        RECT 77.995 86.725 78.285 86.995 ;
        RECT 76.900 86.515 78.285 86.725 ;
        RECT 78.455 86.345 81.045 87.115 ;
        RECT 81.215 86.955 82.325 87.165 ;
        RECT 81.215 86.515 81.565 86.955 ;
        RECT 81.735 86.345 81.905 86.785 ;
        RECT 82.075 86.725 82.325 86.955 ;
        RECT 82.495 87.065 82.820 87.165 ;
        RECT 82.495 86.895 82.825 87.065 ;
        RECT 82.995 86.725 83.270 87.165 ;
        RECT 84.070 87.100 84.240 87.755 ;
        RECT 82.075 86.515 83.270 86.725 ;
        RECT 83.505 86.345 83.835 87.085 ;
        RECT 84.005 86.770 84.240 87.100 ;
        RECT 86.020 86.890 86.360 87.720 ;
        RECT 87.840 87.210 88.190 88.460 ;
        RECT 89.955 87.805 92.545 88.895 ;
        RECT 89.955 87.115 91.165 87.635 ;
        RECT 91.335 87.285 92.545 87.805 ;
        RECT 92.715 87.730 93.005 88.895 ;
        RECT 93.635 88.295 93.895 88.715 ;
        RECT 94.065 88.465 94.395 88.895 ;
        RECT 95.060 88.465 95.805 88.635 ;
        RECT 96.030 88.555 96.670 88.715 ;
        RECT 93.635 88.125 95.465 88.295 ;
        RECT 84.435 86.345 89.780 86.890 ;
        RECT 89.955 86.345 92.545 87.115 ;
        RECT 93.635 87.085 93.805 88.125 ;
        RECT 93.975 87.255 94.325 87.955 ;
        RECT 94.540 87.785 95.125 87.955 ;
        RECT 94.495 87.255 94.785 87.585 ;
        RECT 94.955 87.505 95.125 87.785 ;
        RECT 95.295 87.845 95.465 88.125 ;
        RECT 95.635 88.215 95.805 88.465 ;
        RECT 95.995 88.385 96.670 88.555 ;
        RECT 95.635 88.045 96.670 88.215 ;
        RECT 96.840 88.095 97.120 88.895 ;
        RECT 96.500 87.925 96.670 88.045 ;
        RECT 95.295 87.675 95.945 87.845 ;
        RECT 96.500 87.755 97.160 87.925 ;
        RECT 97.330 87.755 97.605 88.725 ;
        RECT 97.865 87.965 98.035 88.725 ;
        RECT 98.250 88.135 98.580 88.895 ;
        RECT 97.865 87.795 98.580 87.965 ;
        RECT 98.750 87.820 99.005 88.725 ;
        RECT 94.955 87.335 95.380 87.505 ;
        RECT 94.955 87.085 95.125 87.335 ;
        RECT 95.775 87.255 95.945 87.675 ;
        RECT 96.990 87.585 97.160 87.755 ;
        RECT 96.165 87.255 96.820 87.585 ;
        RECT 96.990 87.255 97.265 87.585 ;
        RECT 96.990 87.085 97.160 87.255 ;
        RECT 92.715 86.345 93.005 87.070 ;
        RECT 93.635 86.710 93.950 87.085 ;
        RECT 94.205 86.345 94.375 87.085 ;
        RECT 94.625 86.915 95.125 87.085 ;
        RECT 95.565 86.915 97.160 87.085 ;
        RECT 97.435 87.020 97.605 87.755 ;
        RECT 97.775 87.245 98.130 87.615 ;
        RECT 98.410 87.585 98.580 87.795 ;
        RECT 98.410 87.255 98.665 87.585 ;
        RECT 98.410 87.065 98.580 87.255 ;
        RECT 98.835 87.090 99.005 87.820 ;
        RECT 99.180 87.745 99.440 88.895 ;
        RECT 99.620 88.325 99.940 88.725 ;
        RECT 99.620 87.875 99.790 88.325 ;
        RECT 100.110 88.095 100.420 88.895 ;
        RECT 100.590 88.265 100.920 88.725 ;
        RECT 101.090 88.435 101.260 88.895 ;
        RECT 101.430 88.265 101.760 88.725 ;
        RECT 101.930 88.435 102.180 88.895 ;
        RECT 102.370 88.435 102.620 88.895 ;
        RECT 100.590 88.215 101.760 88.265 ;
        RECT 102.790 88.265 103.040 88.725 ;
        RECT 103.290 88.435 103.580 88.895 ;
        RECT 103.755 88.460 109.100 88.895 ;
        RECT 109.275 88.460 114.620 88.895 ;
        RECT 102.790 88.215 103.580 88.265 ;
        RECT 100.590 88.045 103.580 88.215 ;
        RECT 99.620 87.705 103.180 87.875 ;
        RECT 94.625 86.710 94.795 86.915 ;
        RECT 95.020 86.345 95.395 86.745 ;
        RECT 95.565 86.565 95.735 86.915 ;
        RECT 95.920 86.345 96.250 86.745 ;
        RECT 96.420 86.565 96.590 86.915 ;
        RECT 96.760 86.345 97.140 86.745 ;
        RECT 97.330 86.675 97.605 87.020 ;
        RECT 97.865 86.895 98.580 87.065 ;
        RECT 97.865 86.515 98.035 86.895 ;
        RECT 98.250 86.345 98.580 86.725 ;
        RECT 98.750 86.515 99.005 87.090 ;
        RECT 99.180 86.345 99.440 87.185 ;
        RECT 99.620 86.915 99.790 87.705 ;
        RECT 99.960 87.335 100.310 87.535 ;
        RECT 100.590 87.335 101.270 87.535 ;
        RECT 101.480 87.335 102.670 87.535 ;
        RECT 102.850 87.335 103.180 87.705 ;
        RECT 103.380 87.165 103.580 88.045 ;
        RECT 99.620 86.515 99.940 86.915 ;
        RECT 100.110 86.345 100.420 87.165 ;
        RECT 100.590 86.975 102.280 87.165 ;
        RECT 100.590 86.515 100.920 86.975 ;
        RECT 101.530 86.895 102.280 86.975 ;
        RECT 101.090 86.345 101.340 86.805 ;
        RECT 102.450 86.725 102.620 87.165 ;
        RECT 102.790 86.895 103.580 87.165 ;
        RECT 105.340 86.890 105.680 87.720 ;
        RECT 107.160 87.210 107.510 88.460 ;
        RECT 110.860 86.890 111.200 87.720 ;
        RECT 112.680 87.210 113.030 88.460 ;
        RECT 114.795 87.805 118.305 88.895 ;
        RECT 114.795 87.115 116.445 87.635 ;
        RECT 116.615 87.285 118.305 87.805 ;
        RECT 118.475 87.730 118.765 88.895 ;
        RECT 118.935 87.805 121.525 88.895 ;
        RECT 122.160 88.470 122.495 88.895 ;
        RECT 122.665 88.290 122.850 88.695 ;
        RECT 118.935 87.115 120.145 87.635 ;
        RECT 120.315 87.285 121.525 87.805 ;
        RECT 122.185 88.115 122.850 88.290 ;
        RECT 123.055 88.115 123.385 88.895 ;
        RECT 101.530 86.515 103.580 86.725 ;
        RECT 103.755 86.345 109.100 86.890 ;
        RECT 109.275 86.345 114.620 86.890 ;
        RECT 114.795 86.345 118.305 87.115 ;
        RECT 118.475 86.345 118.765 87.070 ;
        RECT 118.935 86.345 121.525 87.115 ;
        RECT 122.185 87.085 122.525 88.115 ;
        RECT 123.555 87.925 123.825 88.695 ;
        RECT 122.695 87.755 123.825 87.925 ;
        RECT 122.695 87.255 122.945 87.755 ;
        RECT 122.185 86.915 122.870 87.085 ;
        RECT 123.125 87.005 123.485 87.585 ;
        RECT 122.160 86.345 122.495 86.745 ;
        RECT 122.665 86.515 122.870 86.915 ;
        RECT 123.655 86.845 123.825 87.755 ;
        RECT 123.995 87.805 125.205 88.895 ;
        RECT 123.995 87.265 124.515 87.805 ;
        RECT 124.685 87.095 125.205 87.635 ;
        RECT 123.080 86.345 123.355 86.825 ;
        RECT 123.565 86.515 123.825 86.845 ;
        RECT 123.995 86.345 125.205 87.095 ;
        RECT 53.990 86.175 125.290 86.345 ;
        RECT 54.075 85.425 55.285 86.175 ;
        RECT 55.455 85.630 60.800 86.175 ;
        RECT 60.975 85.630 66.320 86.175 ;
        RECT 66.495 85.630 71.840 86.175 ;
        RECT 72.105 85.835 72.275 85.870 ;
        RECT 72.075 85.665 72.275 85.835 ;
        RECT 54.075 84.885 54.595 85.425 ;
        RECT 54.765 84.715 55.285 85.255 ;
        RECT 57.040 84.800 57.380 85.630 ;
        RECT 54.075 83.625 55.285 84.715 ;
        RECT 58.860 84.060 59.210 85.310 ;
        RECT 62.560 84.800 62.900 85.630 ;
        RECT 64.380 84.060 64.730 85.310 ;
        RECT 68.080 84.800 68.420 85.630 ;
        RECT 69.900 84.060 70.250 85.310 ;
        RECT 72.105 85.305 72.275 85.665 ;
        RECT 72.465 85.645 72.695 85.950 ;
        RECT 72.865 85.815 73.195 86.175 ;
        RECT 73.390 85.645 73.680 85.995 ;
        RECT 72.465 85.475 73.680 85.645 ;
        RECT 73.855 85.715 74.415 86.005 ;
        RECT 74.585 85.715 74.835 86.175 ;
        RECT 72.105 85.135 72.625 85.305 ;
        RECT 72.020 84.605 72.265 84.965 ;
        RECT 72.455 84.755 72.625 85.135 ;
        RECT 72.795 84.935 73.180 85.265 ;
        RECT 73.360 85.155 73.620 85.265 ;
        RECT 73.360 84.985 73.625 85.155 ;
        RECT 73.360 84.935 73.620 84.985 ;
        RECT 72.455 84.475 72.805 84.755 ;
        RECT 55.455 83.625 60.800 84.060 ;
        RECT 60.975 83.625 66.320 84.060 ;
        RECT 66.495 83.625 71.840 84.060 ;
        RECT 72.020 83.625 72.275 84.425 ;
        RECT 72.475 83.795 72.805 84.475 ;
        RECT 72.985 83.885 73.180 84.935 ;
        RECT 73.360 83.625 73.680 84.765 ;
        RECT 73.855 84.345 74.105 85.715 ;
        RECT 75.455 85.545 75.785 85.905 ;
        RECT 77.095 85.665 77.335 86.175 ;
        RECT 77.505 85.665 77.795 86.005 ;
        RECT 78.025 85.665 78.340 86.175 ;
        RECT 74.395 85.355 75.785 85.545 ;
        RECT 74.395 85.265 74.565 85.355 ;
        RECT 74.275 84.935 74.565 85.265 ;
        RECT 74.735 84.935 75.075 85.185 ;
        RECT 75.295 84.935 75.970 85.185 ;
        RECT 77.140 85.155 77.335 85.495 ;
        RECT 77.135 84.985 77.335 85.155 ;
        RECT 77.140 84.935 77.335 84.985 ;
        RECT 74.395 84.685 74.565 84.935 ;
        RECT 74.395 84.515 75.335 84.685 ;
        RECT 75.705 84.575 75.970 84.935 ;
        RECT 77.505 84.765 77.685 85.665 ;
        RECT 78.510 85.605 78.680 85.875 ;
        RECT 78.850 85.775 79.180 86.175 ;
        RECT 77.855 84.935 78.265 85.495 ;
        RECT 78.510 85.435 79.205 85.605 ;
        RECT 79.835 85.450 80.125 86.175 ;
        RECT 80.300 85.775 80.635 86.175 ;
        RECT 80.805 85.605 81.010 86.005 ;
        RECT 81.220 85.695 81.495 86.175 ;
        RECT 81.705 85.675 81.965 86.005 ;
        RECT 78.435 84.765 78.605 85.265 ;
        RECT 77.145 84.595 78.605 84.765 ;
        RECT 73.855 83.795 74.315 84.345 ;
        RECT 74.505 83.625 74.835 84.345 ;
        RECT 75.035 83.965 75.335 84.515 ;
        RECT 77.145 84.420 77.505 84.595 ;
        RECT 78.775 84.425 79.205 85.435 ;
        RECT 80.325 85.435 81.010 85.605 ;
        RECT 75.505 83.625 75.785 84.295 ;
        RECT 78.090 83.625 78.260 84.425 ;
        RECT 78.430 84.255 79.205 84.425 ;
        RECT 78.430 83.795 78.760 84.255 ;
        RECT 78.930 83.625 79.100 84.085 ;
        RECT 79.835 83.625 80.125 84.790 ;
        RECT 80.325 84.405 80.665 85.435 ;
        RECT 80.835 84.765 81.085 85.265 ;
        RECT 81.265 84.935 81.625 85.515 ;
        RECT 81.795 84.765 81.965 85.675 ;
        RECT 82.225 85.625 82.395 86.005 ;
        RECT 82.575 85.795 82.905 86.175 ;
        RECT 82.225 85.455 82.890 85.625 ;
        RECT 83.085 85.500 83.345 86.005 ;
        RECT 83.515 85.630 88.860 86.175 ;
        RECT 89.035 85.630 94.380 86.175 ;
        RECT 82.155 84.905 82.485 85.275 ;
        RECT 82.720 85.200 82.890 85.455 ;
        RECT 80.835 84.595 81.965 84.765 ;
        RECT 82.720 84.870 83.005 85.200 ;
        RECT 82.720 84.725 82.890 84.870 ;
        RECT 80.325 84.230 80.990 84.405 ;
        RECT 80.300 83.625 80.635 84.050 ;
        RECT 80.805 83.825 80.990 84.230 ;
        RECT 81.195 83.625 81.525 84.405 ;
        RECT 81.695 83.825 81.965 84.595 ;
        RECT 82.225 84.555 82.890 84.725 ;
        RECT 83.175 84.700 83.345 85.500 ;
        RECT 85.100 84.800 85.440 85.630 ;
        RECT 82.225 83.795 82.395 84.555 ;
        RECT 82.575 83.625 82.905 84.385 ;
        RECT 83.075 83.795 83.345 84.700 ;
        RECT 86.920 84.060 87.270 85.310 ;
        RECT 90.620 84.800 90.960 85.630 ;
        RECT 94.555 85.405 98.065 86.175 ;
        RECT 98.700 85.795 100.750 86.005 ;
        RECT 92.440 84.060 92.790 85.310 ;
        RECT 94.555 84.885 96.205 85.405 ;
        RECT 98.700 85.355 99.490 85.625 ;
        RECT 99.660 85.355 99.830 85.795 ;
        RECT 100.940 85.715 101.190 86.175 ;
        RECT 100.000 85.545 100.750 85.625 ;
        RECT 101.360 85.545 101.690 86.005 ;
        RECT 100.000 85.355 101.690 85.545 ;
        RECT 101.860 85.355 102.170 86.175 ;
        RECT 102.340 85.605 102.660 86.005 ;
        RECT 98.700 85.325 98.925 85.355 ;
        RECT 96.375 84.715 98.065 85.235 ;
        RECT 83.515 83.625 88.860 84.060 ;
        RECT 89.035 83.625 94.380 84.060 ;
        RECT 94.555 83.625 98.065 84.715 ;
        RECT 98.700 84.475 98.900 85.325 ;
        RECT 99.100 84.815 99.430 85.185 ;
        RECT 99.610 84.985 100.800 85.185 ;
        RECT 101.010 84.985 101.690 85.185 ;
        RECT 101.970 84.985 102.320 85.185 ;
        RECT 102.490 84.815 102.660 85.605 ;
        RECT 102.835 85.405 105.425 86.175 ;
        RECT 105.595 85.450 105.885 86.175 ;
        RECT 106.055 85.630 111.400 86.175 ;
        RECT 111.575 85.630 116.920 86.175 ;
        RECT 117.095 85.630 122.440 86.175 ;
        RECT 102.835 84.885 104.045 85.405 ;
        RECT 99.100 84.645 102.660 84.815 ;
        RECT 104.215 84.715 105.425 85.235 ;
        RECT 107.640 84.800 107.980 85.630 ;
        RECT 98.700 84.305 101.690 84.475 ;
        RECT 98.700 84.255 99.490 84.305 ;
        RECT 98.700 83.625 98.990 84.085 ;
        RECT 99.240 83.795 99.490 84.255 ;
        RECT 100.520 84.255 101.690 84.305 ;
        RECT 99.660 83.625 99.910 84.085 ;
        RECT 100.100 83.625 100.350 84.085 ;
        RECT 100.520 83.795 100.850 84.255 ;
        RECT 101.020 83.625 101.190 84.085 ;
        RECT 101.360 83.795 101.690 84.255 ;
        RECT 101.860 83.625 102.170 84.425 ;
        RECT 102.490 84.195 102.660 84.645 ;
        RECT 102.340 83.795 102.660 84.195 ;
        RECT 102.835 83.625 105.425 84.715 ;
        RECT 105.595 83.625 105.885 84.790 ;
        RECT 109.460 84.060 109.810 85.310 ;
        RECT 113.160 84.800 113.500 85.630 ;
        RECT 114.980 84.060 115.330 85.310 ;
        RECT 118.680 84.800 119.020 85.630 ;
        RECT 122.795 85.515 123.135 86.175 ;
        RECT 120.500 84.060 120.850 85.310 ;
        RECT 106.055 83.625 111.400 84.060 ;
        RECT 111.575 83.625 116.920 84.060 ;
        RECT 117.095 83.625 122.440 84.060 ;
        RECT 122.615 83.795 123.135 85.345 ;
        RECT 123.305 84.520 123.825 86.005 ;
        RECT 123.995 85.425 125.205 86.175 ;
        RECT 123.995 84.715 124.515 85.255 ;
        RECT 124.685 84.885 125.205 85.425 ;
        RECT 123.305 83.625 123.635 84.350 ;
        RECT 123.995 83.625 125.205 84.715 ;
        RECT 53.990 83.455 125.290 83.625 ;
        RECT 54.075 82.365 55.285 83.455 ;
        RECT 55.455 83.020 60.800 83.455 ;
        RECT 54.075 81.655 54.595 82.195 ;
        RECT 54.765 81.825 55.285 82.365 ;
        RECT 54.075 80.905 55.285 81.655 ;
        RECT 57.040 81.450 57.380 82.280 ;
        RECT 58.860 81.770 59.210 83.020 ;
        RECT 61.895 81.735 62.415 83.285 ;
        RECT 62.585 82.730 62.915 83.455 ;
        RECT 55.455 80.905 60.800 81.450 ;
        RECT 62.075 80.905 62.415 81.565 ;
        RECT 62.585 81.075 63.105 82.560 ;
        RECT 63.275 82.365 66.785 83.455 ;
        RECT 63.275 81.675 64.925 82.195 ;
        RECT 65.095 81.845 66.785 82.365 ;
        RECT 66.955 82.290 67.245 83.455 ;
        RECT 67.415 82.365 70.925 83.455 ;
        RECT 67.415 81.675 69.065 82.195 ;
        RECT 69.235 81.845 70.925 82.365 ;
        RECT 71.555 82.380 71.825 83.285 ;
        RECT 71.995 82.695 72.325 83.455 ;
        RECT 72.505 82.525 72.675 83.285 ;
        RECT 63.275 80.905 66.785 81.675 ;
        RECT 66.955 80.905 67.245 81.630 ;
        RECT 67.415 80.905 70.925 81.675 ;
        RECT 71.555 81.580 71.725 82.380 ;
        RECT 72.010 82.355 72.675 82.525 ;
        RECT 72.935 82.365 74.605 83.455 ;
        RECT 72.010 82.210 72.180 82.355 ;
        RECT 71.895 81.880 72.180 82.210 ;
        RECT 72.010 81.625 72.180 81.880 ;
        RECT 72.415 81.805 72.745 82.175 ;
        RECT 72.935 81.675 73.685 82.195 ;
        RECT 73.855 81.845 74.605 82.365 ;
        RECT 74.865 82.525 75.035 83.285 ;
        RECT 75.250 82.695 75.580 83.455 ;
        RECT 74.865 82.355 75.580 82.525 ;
        RECT 75.750 82.380 76.005 83.285 ;
        RECT 74.775 81.805 75.130 82.175 ;
        RECT 75.410 82.145 75.580 82.355 ;
        RECT 75.410 81.815 75.665 82.145 ;
        RECT 71.555 81.075 71.815 81.580 ;
        RECT 72.010 81.455 72.675 81.625 ;
        RECT 71.995 80.905 72.325 81.285 ;
        RECT 72.505 81.075 72.675 81.455 ;
        RECT 72.935 80.905 74.605 81.675 ;
        RECT 75.410 81.625 75.580 81.815 ;
        RECT 75.835 81.650 76.005 82.380 ;
        RECT 76.180 82.305 76.440 83.455 ;
        RECT 76.615 82.315 76.875 83.455 ;
        RECT 77.045 82.305 77.375 83.285 ;
        RECT 77.545 82.315 77.825 83.455 ;
        RECT 78.075 82.525 78.255 83.285 ;
        RECT 78.435 82.695 78.765 83.455 ;
        RECT 78.075 82.355 78.750 82.525 ;
        RECT 78.935 82.380 79.205 83.285 ;
        RECT 76.635 81.895 76.970 82.145 ;
        RECT 74.865 81.455 75.580 81.625 ;
        RECT 74.865 81.075 75.035 81.455 ;
        RECT 75.250 80.905 75.580 81.285 ;
        RECT 75.750 81.075 76.005 81.650 ;
        RECT 76.180 80.905 76.440 81.745 ;
        RECT 77.140 81.705 77.310 82.305 ;
        RECT 78.580 82.210 78.750 82.355 ;
        RECT 77.480 81.875 77.815 82.145 ;
        RECT 78.015 81.805 78.355 82.175 ;
        RECT 78.580 81.880 78.855 82.210 ;
        RECT 76.615 81.075 77.310 81.705 ;
        RECT 77.515 80.905 77.825 81.705 ;
        RECT 78.580 81.625 78.750 81.880 ;
        RECT 78.085 81.455 78.750 81.625 ;
        RECT 79.025 81.580 79.205 82.380 ;
        RECT 79.835 82.290 80.125 83.455 ;
        RECT 81.215 82.485 81.485 83.255 ;
        RECT 81.655 82.675 81.985 83.455 ;
        RECT 82.190 82.850 82.375 83.255 ;
        RECT 82.545 83.030 82.880 83.455 ;
        RECT 82.190 82.675 82.855 82.850 ;
        RECT 81.215 82.315 82.345 82.485 ;
        RECT 78.085 81.075 78.255 81.455 ;
        RECT 78.435 80.905 78.765 81.285 ;
        RECT 78.945 81.075 79.205 81.580 ;
        RECT 79.835 80.905 80.125 81.630 ;
        RECT 81.215 81.405 81.385 82.315 ;
        RECT 81.555 81.565 81.915 82.145 ;
        RECT 82.095 81.815 82.345 82.315 ;
        RECT 82.515 81.645 82.855 82.675 ;
        RECT 83.055 82.365 84.265 83.455 ;
        RECT 82.170 81.475 82.855 81.645 ;
        RECT 83.055 81.655 83.575 82.195 ;
        RECT 83.745 81.825 84.265 82.365 ;
        RECT 84.525 82.525 84.695 83.285 ;
        RECT 84.910 82.695 85.240 83.455 ;
        RECT 84.525 82.355 85.240 82.525 ;
        RECT 85.410 82.380 85.665 83.285 ;
        RECT 84.435 81.805 84.790 82.175 ;
        RECT 85.070 82.145 85.240 82.355 ;
        RECT 85.070 81.815 85.325 82.145 ;
        RECT 81.215 81.075 81.475 81.405 ;
        RECT 81.685 80.905 81.960 81.385 ;
        RECT 82.170 81.075 82.375 81.475 ;
        RECT 82.545 80.905 82.880 81.305 ;
        RECT 83.055 80.905 84.265 81.655 ;
        RECT 85.070 81.625 85.240 81.815 ;
        RECT 85.495 81.650 85.665 82.380 ;
        RECT 85.840 82.305 86.100 83.455 ;
        RECT 86.275 83.020 91.620 83.455 ;
        RECT 84.525 81.455 85.240 81.625 ;
        RECT 84.525 81.075 84.695 81.455 ;
        RECT 84.910 80.905 85.240 81.285 ;
        RECT 85.410 81.075 85.665 81.650 ;
        RECT 85.840 80.905 86.100 81.745 ;
        RECT 87.860 81.450 88.200 82.280 ;
        RECT 89.680 81.770 90.030 83.020 ;
        RECT 92.715 82.290 93.005 83.455 ;
        RECT 93.175 83.020 98.520 83.455 ;
        RECT 98.695 83.020 104.040 83.455 ;
        RECT 86.275 80.905 91.620 81.450 ;
        RECT 92.715 80.905 93.005 81.630 ;
        RECT 94.760 81.450 95.100 82.280 ;
        RECT 96.580 81.770 96.930 83.020 ;
        RECT 100.280 81.450 100.620 82.280 ;
        RECT 102.100 81.770 102.450 83.020 ;
        RECT 104.215 82.365 105.425 83.455 ;
        RECT 104.215 81.655 104.735 82.195 ;
        RECT 104.905 81.825 105.425 82.365 ;
        RECT 105.595 82.290 105.885 83.455 ;
        RECT 106.055 83.020 111.400 83.455 ;
        RECT 111.575 83.020 116.920 83.455 ;
        RECT 93.175 80.905 98.520 81.450 ;
        RECT 98.695 80.905 104.040 81.450 ;
        RECT 104.215 80.905 105.425 81.655 ;
        RECT 105.595 80.905 105.885 81.630 ;
        RECT 107.640 81.450 107.980 82.280 ;
        RECT 109.460 81.770 109.810 83.020 ;
        RECT 113.160 81.450 113.500 82.280 ;
        RECT 114.980 81.770 115.330 83.020 ;
        RECT 117.095 82.365 118.305 83.455 ;
        RECT 117.095 81.655 117.615 82.195 ;
        RECT 117.785 81.825 118.305 82.365 ;
        RECT 118.475 82.290 118.765 83.455 ;
        RECT 118.935 82.365 122.445 83.455 ;
        RECT 122.615 82.365 123.825 83.455 ;
        RECT 118.935 81.675 120.585 82.195 ;
        RECT 120.755 81.845 122.445 82.365 ;
        RECT 106.055 80.905 111.400 81.450 ;
        RECT 111.575 80.905 116.920 81.450 ;
        RECT 117.095 80.905 118.305 81.655 ;
        RECT 118.475 80.905 118.765 81.630 ;
        RECT 118.935 80.905 122.445 81.675 ;
        RECT 122.615 81.655 123.135 82.195 ;
        RECT 123.305 81.825 123.825 82.365 ;
        RECT 123.995 82.365 125.205 83.455 ;
        RECT 123.995 81.825 124.515 82.365 ;
        RECT 124.685 81.655 125.205 82.195 ;
        RECT 122.615 80.905 123.825 81.655 ;
        RECT 123.995 80.905 125.205 81.655 ;
        RECT 53.990 80.735 125.290 80.905 ;
      LAYER met1 ;
        RECT 57.740 155.860 58.060 155.920 ;
        RECT 77.520 155.860 77.840 155.920 ;
        RECT 57.740 155.720 77.840 155.860 ;
        RECT 57.740 155.660 58.060 155.720 ;
        RECT 77.520 155.660 77.840 155.720 ;
        RECT 60.500 154.840 60.820 154.900 ;
        RECT 116.160 154.840 116.480 154.900 ;
        RECT 60.500 154.700 116.480 154.840 ;
        RECT 60.500 154.640 60.820 154.700 ;
        RECT 116.160 154.640 116.480 154.700 ;
        RECT 62.340 154.500 62.660 154.560 ;
        RECT 68.320 154.500 68.640 154.560 ;
        RECT 117.540 154.500 117.860 154.560 ;
        RECT 62.340 154.360 117.860 154.500 ;
        RECT 62.340 154.300 62.660 154.360 ;
        RECT 68.320 154.300 68.640 154.360 ;
        RECT 117.540 154.300 117.860 154.360 ;
        RECT 60.960 154.160 61.280 154.220 ;
        RECT 90.400 154.160 90.720 154.220 ;
        RECT 60.960 154.020 90.720 154.160 ;
        RECT 60.960 153.960 61.280 154.020 ;
        RECT 90.400 153.960 90.720 154.020 ;
        RECT 55.440 153.820 55.760 153.880 ;
        RECT 67.860 153.820 68.180 153.880 ;
        RECT 55.440 153.680 68.180 153.820 ;
        RECT 55.440 153.620 55.760 153.680 ;
        RECT 67.860 153.620 68.180 153.680 ;
        RECT 72.460 153.820 72.780 153.880 ;
        RECT 95.000 153.820 95.320 153.880 ;
        RECT 72.460 153.680 95.320 153.820 ;
        RECT 72.460 153.620 72.780 153.680 ;
        RECT 95.000 153.620 95.320 153.680 ;
        RECT 52.680 153.140 53.000 153.200 ;
        RECT 58.200 153.140 58.520 153.200 ;
        RECT 52.680 153.000 58.520 153.140 ;
        RECT 52.680 152.940 53.000 153.000 ;
        RECT 58.200 152.940 58.520 153.000 ;
        RECT 71.080 153.140 71.400 153.200 ;
        RECT 77.980 153.140 78.300 153.200 ;
        RECT 71.080 153.000 78.300 153.140 ;
        RECT 71.080 152.940 71.400 153.000 ;
        RECT 77.980 152.940 78.300 153.000 ;
        RECT 95.460 153.140 95.780 153.200 ;
        RECT 118.460 153.140 118.780 153.200 ;
        RECT 95.460 153.000 118.780 153.140 ;
        RECT 95.460 152.940 95.780 153.000 ;
        RECT 118.460 152.940 118.780 153.000 ;
        RECT 65.560 152.800 65.880 152.860 ;
        RECT 97.300 152.800 97.620 152.860 ;
        RECT 65.560 152.660 97.620 152.800 ;
        RECT 65.560 152.600 65.880 152.660 ;
        RECT 97.300 152.600 97.620 152.660 ;
        RECT 66.940 152.460 67.260 152.520 ;
        RECT 107.420 152.460 107.740 152.520 ;
        RECT 66.940 152.320 107.740 152.460 ;
        RECT 66.940 152.260 67.260 152.320 ;
        RECT 107.420 152.260 107.740 152.320 ;
        RECT 60.040 152.120 60.360 152.180 ;
        RECT 77.520 152.120 77.840 152.180 ;
        RECT 60.040 151.980 77.840 152.120 ;
        RECT 60.040 151.920 60.360 151.980 ;
        RECT 77.520 151.920 77.840 151.980 ;
        RECT 53.990 151.300 125.290 151.780 ;
        RECT 57.740 150.900 58.060 151.160 ;
        RECT 60.960 150.900 61.280 151.160 ;
        RECT 65.100 151.100 65.420 151.160 ;
        RECT 98.680 151.100 99.000 151.160 ;
        RECT 103.280 151.100 103.600 151.160 ;
        RECT 61.970 150.960 65.420 151.100 ;
        RECT 55.915 150.760 56.205 150.805 ;
        RECT 61.970 150.760 62.110 150.960 ;
        RECT 65.100 150.900 65.420 150.960 ;
        RECT 68.410 150.960 103.600 151.100 ;
        RECT 55.915 150.620 57.050 150.760 ;
        RECT 55.915 150.575 56.205 150.620 ;
        RECT 56.910 150.480 57.050 150.620 ;
        RECT 60.130 150.620 62.110 150.760 ;
        RECT 56.375 150.235 56.665 150.465 ;
        RECT 56.450 150.080 56.590 150.235 ;
        RECT 56.820 150.220 57.140 150.480 ;
        RECT 60.130 150.465 60.270 150.620 ;
        RECT 62.340 150.560 62.660 150.820 ;
        RECT 60.055 150.235 60.345 150.465 ;
        RECT 61.880 150.220 62.200 150.480 ;
        RECT 63.260 150.220 63.580 150.480 ;
        RECT 65.560 150.220 65.880 150.480 ;
        RECT 66.480 150.220 66.800 150.480 ;
        RECT 68.410 150.465 68.550 150.960 ;
        RECT 98.680 150.900 99.000 150.960 ;
        RECT 103.280 150.900 103.600 150.960 ;
        RECT 103.830 150.960 110.640 151.100 ;
        RECT 72.920 150.760 73.240 150.820 ;
        RECT 81.215 150.760 81.505 150.805 ;
        RECT 69.330 150.620 81.505 150.760 ;
        RECT 69.330 150.465 69.470 150.620 ;
        RECT 72.920 150.560 73.240 150.620 ;
        RECT 81.215 150.575 81.505 150.620 ;
        RECT 89.955 150.760 90.245 150.805 ;
        RECT 92.700 150.760 93.020 150.820 ;
        RECT 89.955 150.620 93.020 150.760 ;
        RECT 89.955 150.575 90.245 150.620 ;
        RECT 92.700 150.560 93.020 150.620 ;
        RECT 101.900 150.760 102.220 150.820 ;
        RECT 103.830 150.760 103.970 150.960 ;
        RECT 101.900 150.620 103.970 150.760 ;
        RECT 107.420 150.760 107.740 150.820 ;
        RECT 109.260 150.760 109.580 150.820 ;
        RECT 107.420 150.620 109.580 150.760 ;
        RECT 110.500 150.760 110.640 150.960 ;
        RECT 117.540 150.900 117.860 151.160 ;
        RECT 110.500 150.620 120.990 150.760 ;
        RECT 101.900 150.560 102.220 150.620 ;
        RECT 107.420 150.560 107.740 150.620 ;
        RECT 109.260 150.560 109.580 150.620 ;
        RECT 68.335 150.235 68.625 150.465 ;
        RECT 69.255 150.235 69.545 150.465 ;
        RECT 70.635 150.235 70.925 150.465 ;
        RECT 72.460 150.420 72.780 150.480 ;
        RECT 73.395 150.420 73.685 150.465 ;
        RECT 72.460 150.280 73.685 150.420 ;
        RECT 66.940 150.080 67.260 150.140 ;
        RECT 56.450 149.940 67.260 150.080 ;
        RECT 66.940 149.880 67.260 149.940 ;
        RECT 67.860 150.080 68.180 150.140 ;
        RECT 67.860 149.940 69.470 150.080 ;
        RECT 67.860 149.880 68.180 149.940 ;
        RECT 59.135 149.740 59.425 149.785 ;
        RECT 67.400 149.740 67.720 149.800 ;
        RECT 59.135 149.600 67.720 149.740 ;
        RECT 59.135 149.555 59.425 149.600 ;
        RECT 67.400 149.540 67.720 149.600 ;
        RECT 68.780 149.540 69.100 149.800 ;
        RECT 69.330 149.740 69.470 149.940 ;
        RECT 69.700 149.880 70.020 150.140 ;
        RECT 70.710 149.740 70.850 150.235 ;
        RECT 72.460 150.220 72.780 150.280 ;
        RECT 73.395 150.235 73.685 150.280 ;
        RECT 73.840 150.220 74.160 150.480 ;
        RECT 74.300 150.220 74.620 150.480 ;
        RECT 75.680 150.220 76.000 150.480 ;
        RECT 76.435 150.235 76.725 150.465 ;
        RECT 71.080 150.080 71.400 150.140 ;
        RECT 74.760 150.080 75.080 150.140 ;
        RECT 71.080 149.940 75.080 150.080 ;
        RECT 71.080 149.880 71.400 149.940 ;
        RECT 69.330 149.600 70.850 149.740 ;
        RECT 71.540 149.540 71.860 149.800 ;
        RECT 72.550 149.785 72.690 149.940 ;
        RECT 74.760 149.880 75.080 149.940 ;
        RECT 72.475 149.555 72.765 149.785 ;
        RECT 76.510 149.740 76.650 150.235 ;
        RECT 77.520 150.220 77.840 150.480 ;
        RECT 78.440 150.220 78.760 150.480 ;
        RECT 90.415 150.420 90.705 150.465 ;
        RECT 90.860 150.420 91.180 150.480 ;
        RECT 90.415 150.280 91.180 150.420 ;
        RECT 90.415 150.235 90.705 150.280 ;
        RECT 90.860 150.220 91.180 150.280 ;
        RECT 91.335 150.420 91.625 150.465 ;
        RECT 96.840 150.420 97.160 150.480 ;
        RECT 91.335 150.280 97.160 150.420 ;
        RECT 91.335 150.235 91.625 150.280 ;
        RECT 96.840 150.220 97.160 150.280 ;
        RECT 105.120 150.220 105.440 150.480 ;
        RECT 105.580 150.420 105.900 150.480 ;
        RECT 106.055 150.420 106.345 150.465 ;
        RECT 105.580 150.280 106.345 150.420 ;
        RECT 105.580 150.220 105.900 150.280 ;
        RECT 106.055 150.235 106.345 150.280 ;
        RECT 106.500 150.220 106.820 150.480 ;
        RECT 107.895 150.420 108.185 150.465 ;
        RECT 111.100 150.420 111.420 150.480 ;
        RECT 107.895 150.280 111.420 150.420 ;
        RECT 107.895 150.235 108.185 150.280 ;
        RECT 111.100 150.220 111.420 150.280 ;
        RECT 117.080 150.220 117.400 150.480 ;
        RECT 120.850 150.465 120.990 150.620 ;
        RECT 120.775 150.235 121.065 150.465 ;
        RECT 123.520 150.220 123.840 150.480 ;
        RECT 77.060 149.880 77.380 150.140 ;
        RECT 93.620 149.880 93.940 150.140 ;
        RECT 94.080 149.880 94.400 150.140 ;
        RECT 94.540 149.880 94.860 150.140 ;
        RECT 95.015 149.895 95.305 150.125 ;
        RECT 95.935 150.080 96.225 150.125 ;
        RECT 95.935 149.940 116.390 150.080 ;
        RECT 95.935 149.895 96.225 149.940 ;
        RECT 73.010 149.600 76.650 149.740 ;
        RECT 79.375 149.740 79.665 149.785 ;
        RECT 85.800 149.740 86.120 149.800 ;
        RECT 95.090 149.740 95.230 149.895 ;
        RECT 79.375 149.600 86.120 149.740 ;
        RECT 64.180 149.200 64.500 149.460 ;
        RECT 66.020 149.200 66.340 149.460 ;
        RECT 66.480 149.400 66.800 149.460 ;
        RECT 73.010 149.400 73.150 149.600 ;
        RECT 79.375 149.555 79.665 149.600 ;
        RECT 85.800 149.540 86.120 149.600 ;
        RECT 86.350 149.600 95.230 149.740 ;
        RECT 98.695 149.740 98.985 149.785 ;
        RECT 111.100 149.740 111.420 149.800 ;
        RECT 98.695 149.600 111.420 149.740 ;
        RECT 66.480 149.260 73.150 149.400 ;
        RECT 66.480 149.200 66.800 149.260 ;
        RECT 75.220 149.200 75.540 149.460 ;
        RECT 76.600 149.400 76.920 149.460 ;
        RECT 86.350 149.400 86.490 149.600 ;
        RECT 98.695 149.555 98.985 149.600 ;
        RECT 111.100 149.540 111.420 149.600 ;
        RECT 76.600 149.260 86.490 149.400 ;
        RECT 76.600 149.200 76.920 149.260 ;
        RECT 91.780 149.200 92.100 149.460 ;
        RECT 104.200 149.400 104.520 149.460 ;
        RECT 107.435 149.400 107.725 149.445 ;
        RECT 104.200 149.260 107.725 149.400 ;
        RECT 116.250 149.400 116.390 149.940 ;
        RECT 116.620 149.880 116.940 150.140 ;
        RECT 118.920 149.880 119.240 150.140 ;
        RECT 121.235 150.080 121.525 150.125 ;
        RECT 123.060 150.080 123.380 150.140 ;
        RECT 121.235 149.940 123.380 150.080 ;
        RECT 121.235 149.895 121.525 149.940 ;
        RECT 123.060 149.880 123.380 149.940 ;
        RECT 118.000 149.740 118.320 149.800 ;
        RECT 122.615 149.740 122.905 149.785 ;
        RECT 118.000 149.600 122.905 149.740 ;
        RECT 118.000 149.540 118.320 149.600 ;
        RECT 122.615 149.555 122.905 149.600 ;
        RECT 120.300 149.400 120.620 149.460 ;
        RECT 116.250 149.260 120.620 149.400 ;
        RECT 104.200 149.200 104.520 149.260 ;
        RECT 107.435 149.215 107.725 149.260 ;
        RECT 120.300 149.200 120.620 149.260 ;
        RECT 121.220 149.400 121.540 149.460 ;
        RECT 122.155 149.400 122.445 149.445 ;
        RECT 121.220 149.260 122.445 149.400 ;
        RECT 121.220 149.200 121.540 149.260 ;
        RECT 122.155 149.215 122.445 149.260 ;
        RECT 53.990 148.580 125.290 149.060 ;
        RECT 53.600 148.380 53.920 148.440 ;
        RECT 59.135 148.380 59.425 148.425 ;
        RECT 53.600 148.240 59.425 148.380 ;
        RECT 53.600 148.180 53.920 148.240 ;
        RECT 59.135 148.195 59.425 148.240 ;
        RECT 62.800 148.380 63.120 148.440 ;
        RECT 64.655 148.380 64.945 148.425 ;
        RECT 62.800 148.240 64.945 148.380 ;
        RECT 62.800 148.180 63.120 148.240 ;
        RECT 64.655 148.195 64.945 148.240 ;
        RECT 65.100 148.380 65.420 148.440 ;
        RECT 67.400 148.380 67.720 148.440 ;
        RECT 71.080 148.380 71.400 148.440 ;
        RECT 65.100 148.240 67.720 148.380 ;
        RECT 65.100 148.180 65.420 148.240 ;
        RECT 67.400 148.180 67.720 148.240 ;
        RECT 68.970 148.240 71.400 148.380 ;
        RECT 57.740 148.040 58.060 148.100 ;
        RECT 61.420 148.040 61.740 148.100 ;
        RECT 65.560 148.040 65.880 148.100 ;
        RECT 68.970 148.040 69.110 148.240 ;
        RECT 71.080 148.180 71.400 148.240 ;
        RECT 103.280 148.380 103.600 148.440 ;
        RECT 106.975 148.380 107.265 148.425 ;
        RECT 103.280 148.240 107.265 148.380 ;
        RECT 103.280 148.180 103.600 148.240 ;
        RECT 106.975 148.195 107.265 148.240 ;
        RECT 108.800 148.380 109.120 148.440 ;
        RECT 108.800 148.240 119.150 148.380 ;
        RECT 108.800 148.180 109.120 148.240 ;
        RECT 77.535 148.040 77.825 148.085 ;
        RECT 78.440 148.040 78.760 148.100 ;
        RECT 85.340 148.040 85.660 148.100 ;
        RECT 57.740 147.900 61.190 148.040 ;
        RECT 57.740 147.840 58.060 147.900 ;
        RECT 58.215 147.700 58.505 147.745 ;
        RECT 61.050 147.700 61.190 147.900 ;
        RECT 61.420 147.900 69.110 148.040 ;
        RECT 69.330 147.900 76.650 148.040 ;
        RECT 61.420 147.840 61.740 147.900 ;
        RECT 65.560 147.840 65.880 147.900 ;
        RECT 66.480 147.700 66.800 147.760 ;
        RECT 58.215 147.560 60.730 147.700 ;
        RECT 61.050 147.560 66.800 147.700 ;
        RECT 58.215 147.515 58.505 147.560 ;
        RECT 57.280 147.160 57.600 147.420 ;
        RECT 60.055 147.175 60.345 147.405 ;
        RECT 60.590 147.360 60.730 147.560 ;
        RECT 66.480 147.500 66.800 147.560 ;
        RECT 60.975 147.360 61.265 147.405 ;
        RECT 60.590 147.220 61.265 147.360 ;
        RECT 60.975 147.175 61.265 147.220 ;
        RECT 61.435 147.360 61.725 147.405 ;
        RECT 62.340 147.360 62.660 147.420 ;
        RECT 61.435 147.220 62.660 147.360 ;
        RECT 61.435 147.175 61.725 147.220 ;
        RECT 53.140 147.020 53.460 147.080 ;
        RECT 60.130 147.020 60.270 147.175 ;
        RECT 53.140 146.880 60.270 147.020 ;
        RECT 61.050 147.020 61.190 147.175 ;
        RECT 62.340 147.160 62.660 147.220 ;
        RECT 62.815 147.360 63.105 147.405 ;
        RECT 64.180 147.360 64.500 147.420 ;
        RECT 62.815 147.220 64.500 147.360 ;
        RECT 62.815 147.175 63.105 147.220 ;
        RECT 64.180 147.160 64.500 147.220 ;
        RECT 66.020 147.160 66.340 147.420 ;
        RECT 69.330 147.405 69.470 147.900 ;
        RECT 70.160 147.700 70.480 147.760 ;
        RECT 74.760 147.700 75.080 147.760 ;
        RECT 76.510 147.700 76.650 147.900 ;
        RECT 77.535 147.900 85.660 148.040 ;
        RECT 77.535 147.855 77.825 147.900 ;
        RECT 78.440 147.840 78.760 147.900 ;
        RECT 85.340 147.840 85.660 147.900 ;
        RECT 90.400 148.040 90.720 148.100 ;
        RECT 94.540 148.040 94.860 148.100 ;
        RECT 113.400 148.040 113.720 148.100 ;
        RECT 116.635 148.040 116.925 148.085 ;
        RECT 90.400 147.900 113.720 148.040 ;
        RECT 90.400 147.840 90.720 147.900 ;
        RECT 94.540 147.840 94.860 147.900 ;
        RECT 113.400 147.840 113.720 147.900 ;
        RECT 114.410 147.900 116.925 148.040 ;
        RECT 95.935 147.700 96.225 147.745 ;
        RECT 96.380 147.700 96.700 147.760 ;
        RECT 106.040 147.700 106.360 147.760 ;
        RECT 70.160 147.560 73.610 147.700 ;
        RECT 70.160 147.500 70.480 147.560 ;
        RECT 73.470 147.420 73.610 147.560 ;
        RECT 74.760 147.560 76.365 147.700 ;
        RECT 76.510 147.560 90.170 147.700 ;
        RECT 74.760 147.500 75.080 147.560 ;
        RECT 69.255 147.175 69.545 147.405 ;
        RECT 63.260 147.020 63.580 147.080 ;
        RECT 61.050 146.880 63.580 147.020 ;
        RECT 53.140 146.820 53.460 146.880 ;
        RECT 63.260 146.820 63.580 146.880 ;
        RECT 63.720 147.020 64.040 147.080 ;
        RECT 64.885 147.020 65.175 147.065 ;
        RECT 69.330 147.020 69.470 147.175 ;
        RECT 69.700 147.160 70.020 147.420 ;
        RECT 70.635 147.175 70.925 147.405 ;
        RECT 71.095 147.360 71.385 147.405 ;
        RECT 72.015 147.360 72.305 147.405 ;
        RECT 71.095 147.220 72.305 147.360 ;
        RECT 71.095 147.175 71.385 147.220 ;
        RECT 72.015 147.175 72.305 147.220 ;
        RECT 63.720 146.880 69.470 147.020 ;
        RECT 70.710 147.020 70.850 147.175 ;
        RECT 73.380 147.160 73.700 147.420 ;
        RECT 73.840 147.160 74.160 147.420 ;
        RECT 75.680 147.160 76.000 147.420 ;
        RECT 76.225 147.360 76.365 147.560 ;
        RECT 79.360 147.360 79.680 147.420 ;
        RECT 76.225 147.220 79.680 147.360 ;
        RECT 79.360 147.160 79.680 147.220 ;
        RECT 83.040 147.360 83.360 147.420 ;
        RECT 83.975 147.360 84.265 147.405 ;
        RECT 83.040 147.220 84.265 147.360 ;
        RECT 83.040 147.160 83.360 147.220 ;
        RECT 83.975 147.175 84.265 147.220 ;
        RECT 84.435 147.175 84.725 147.405 ;
        RECT 72.460 147.020 72.780 147.080 ;
        RECT 70.710 146.880 72.780 147.020 ;
        RECT 63.720 146.820 64.040 146.880 ;
        RECT 64.885 146.835 65.175 146.880 ;
        RECT 72.460 146.820 72.780 146.880 ;
        RECT 74.775 147.020 75.065 147.065 ;
        RECT 75.770 147.020 75.910 147.160 ;
        RECT 77.520 147.020 77.840 147.080 ;
        RECT 74.775 146.880 77.840 147.020 ;
        RECT 74.775 146.835 75.065 146.880 ;
        RECT 77.520 146.820 77.840 146.880 ;
        RECT 83.500 147.020 83.820 147.080 ;
        RECT 84.510 147.020 84.650 147.175 ;
        RECT 84.880 147.160 85.200 147.420 ;
        RECT 85.800 147.160 86.120 147.420 ;
        RECT 86.835 147.405 86.975 147.560 ;
        RECT 90.030 147.420 90.170 147.560 ;
        RECT 95.935 147.560 96.700 147.700 ;
        RECT 95.935 147.515 96.225 147.560 ;
        RECT 96.380 147.500 96.700 147.560 ;
        RECT 96.930 147.560 106.360 147.700 ;
        RECT 86.760 147.175 87.050 147.405 ;
        RECT 88.560 147.160 88.880 147.420 ;
        RECT 89.020 147.160 89.340 147.420 ;
        RECT 89.940 147.160 90.260 147.420 ;
        RECT 90.415 147.360 90.705 147.405 ;
        RECT 96.930 147.360 97.070 147.560 ;
        RECT 106.040 147.500 106.360 147.560 ;
        RECT 112.035 147.700 112.325 147.745 ;
        RECT 114.410 147.700 114.550 147.900 ;
        RECT 116.635 147.855 116.925 147.900 ;
        RECT 112.035 147.560 114.550 147.700 ;
        RECT 112.035 147.515 112.325 147.560 ;
        RECT 115.240 147.500 115.560 147.760 ;
        RECT 119.010 147.745 119.150 148.240 ;
        RECT 122.155 148.040 122.445 148.085 ;
        RECT 119.470 147.900 122.445 148.040 ;
        RECT 115.715 147.700 116.005 147.745 ;
        RECT 115.715 147.560 118.690 147.700 ;
        RECT 115.715 147.515 116.005 147.560 ;
        RECT 90.415 147.220 97.070 147.360 ;
        RECT 90.415 147.175 90.705 147.220 ;
        RECT 97.300 147.160 97.620 147.420 ;
        RECT 103.740 147.360 104.060 147.420 ;
        RECT 109.735 147.360 110.025 147.405 ;
        RECT 103.740 147.220 110.025 147.360 ;
        RECT 103.740 147.160 104.060 147.220 ;
        RECT 109.735 147.175 110.025 147.220 ;
        RECT 111.560 147.160 111.880 147.420 ;
        RECT 113.400 147.160 113.720 147.420 ;
        RECT 118.000 147.160 118.320 147.420 ;
        RECT 118.550 147.360 118.690 147.560 ;
        RECT 118.935 147.515 119.225 147.745 ;
        RECT 119.470 147.360 119.610 147.900 ;
        RECT 122.155 147.855 122.445 147.900 ;
        RECT 121.220 147.500 121.540 147.760 ;
        RECT 118.550 147.220 119.610 147.360 ;
        RECT 120.760 147.160 121.080 147.420 ;
        RECT 123.520 147.160 123.840 147.420 ;
        RECT 83.500 146.880 84.650 147.020 ;
        RECT 83.500 146.820 83.820 146.880 ;
        RECT 86.260 146.820 86.580 147.080 ;
        RECT 87.180 147.020 87.500 147.080 ;
        RECT 93.635 147.020 93.925 147.065 ;
        RECT 96.840 147.020 97.160 147.080 ;
        RECT 99.600 147.020 99.920 147.080 ;
        RECT 87.180 146.880 92.010 147.020 ;
        RECT 87.180 146.820 87.500 146.880 ;
        RECT 54.060 146.680 54.380 146.740 ;
        RECT 56.375 146.680 56.665 146.725 ;
        RECT 54.060 146.540 56.665 146.680 ;
        RECT 54.060 146.480 54.380 146.540 ;
        RECT 56.375 146.495 56.665 146.540 ;
        RECT 57.280 146.680 57.600 146.740 ;
        RECT 61.420 146.680 61.740 146.740 ;
        RECT 57.280 146.540 61.740 146.680 ;
        RECT 57.280 146.480 57.600 146.540 ;
        RECT 61.420 146.480 61.740 146.540 ;
        RECT 62.355 146.680 62.645 146.725 ;
        RECT 66.940 146.680 67.260 146.740 ;
        RECT 62.355 146.540 67.260 146.680 ;
        RECT 62.355 146.495 62.645 146.540 ;
        RECT 66.940 146.480 67.260 146.540 ;
        RECT 68.335 146.680 68.625 146.725 ;
        RECT 68.780 146.680 69.100 146.740 ;
        RECT 68.335 146.540 69.100 146.680 ;
        RECT 68.335 146.495 68.625 146.540 ;
        RECT 68.780 146.480 69.100 146.540 ;
        RECT 71.080 146.680 71.400 146.740 ;
        RECT 72.935 146.680 73.225 146.725 ;
        RECT 80.280 146.680 80.600 146.740 ;
        RECT 71.080 146.540 80.600 146.680 ;
        RECT 71.080 146.480 71.400 146.540 ;
        RECT 72.935 146.495 73.225 146.540 ;
        RECT 80.280 146.480 80.600 146.540 ;
        RECT 84.420 146.680 84.740 146.740 ;
        RECT 87.655 146.680 87.945 146.725 ;
        RECT 84.420 146.540 87.945 146.680 ;
        RECT 84.420 146.480 84.740 146.540 ;
        RECT 87.655 146.495 87.945 146.540 ;
        RECT 91.320 146.480 91.640 146.740 ;
        RECT 91.870 146.680 92.010 146.880 ;
        RECT 93.635 146.880 99.920 147.020 ;
        RECT 93.635 146.835 93.925 146.880 ;
        RECT 96.840 146.820 97.160 146.880 ;
        RECT 99.600 146.820 99.920 146.880 ;
        RECT 100.535 146.835 100.825 147.065 ;
        RECT 106.960 147.020 107.280 147.080 ;
        RECT 112.955 147.020 113.245 147.065 ;
        RECT 121.680 147.020 122.000 147.080 ;
        RECT 106.960 146.880 113.245 147.020 ;
        RECT 100.610 146.680 100.750 146.835 ;
        RECT 106.960 146.820 107.280 146.880 ;
        RECT 112.955 146.835 113.245 146.880 ;
        RECT 113.490 146.880 122.000 147.020 ;
        RECT 91.870 146.540 100.750 146.680 ;
        RECT 107.420 146.680 107.740 146.740 ;
        RECT 113.490 146.680 113.630 146.880 ;
        RECT 121.680 146.820 122.000 146.880 ;
        RECT 107.420 146.540 113.630 146.680 ;
        RECT 107.420 146.480 107.740 146.540 ;
        RECT 117.540 146.480 117.860 146.740 ;
        RECT 122.140 146.680 122.460 146.740 ;
        RECT 122.615 146.680 122.905 146.725 ;
        RECT 122.140 146.540 122.905 146.680 ;
        RECT 122.140 146.480 122.460 146.540 ;
        RECT 122.615 146.495 122.905 146.540 ;
        RECT 53.990 145.860 125.290 146.340 ;
        RECT 54.520 145.660 54.840 145.720 ;
        RECT 55.915 145.660 56.205 145.705 ;
        RECT 54.520 145.520 56.205 145.660 ;
        RECT 54.520 145.460 54.840 145.520 ;
        RECT 55.915 145.475 56.205 145.520 ;
        RECT 57.740 145.460 58.060 145.720 ;
        RECT 61.880 145.660 62.200 145.720 ;
        RECT 58.750 145.520 62.200 145.660 ;
        RECT 56.360 144.980 56.680 145.040 ;
        RECT 56.835 144.980 57.125 145.025 ;
        RECT 56.360 144.840 57.125 144.980 ;
        RECT 56.360 144.780 56.680 144.840 ;
        RECT 56.835 144.795 57.125 144.840 ;
        RECT 57.280 144.780 57.600 145.040 ;
        RECT 58.750 145.025 58.890 145.520 ;
        RECT 61.880 145.460 62.200 145.520 ;
        RECT 63.720 145.460 64.040 145.720 ;
        RECT 93.620 145.660 93.940 145.720 ;
        RECT 105.120 145.660 105.440 145.720 ;
        RECT 64.255 145.520 93.940 145.660 ;
        RECT 59.135 145.320 59.425 145.365 ;
        RECT 64.255 145.320 64.395 145.520 ;
        RECT 93.620 145.460 93.940 145.520 ;
        RECT 94.170 145.520 105.440 145.660 ;
        RECT 59.135 145.180 64.395 145.320 ;
        RECT 59.135 145.135 59.425 145.180 ;
        RECT 64.655 145.135 64.945 145.365 ;
        RECT 66.480 145.320 66.800 145.380 ;
        RECT 70.160 145.320 70.480 145.380 ;
        RECT 66.480 145.180 70.480 145.320 ;
        RECT 58.215 144.795 58.505 145.025 ;
        RECT 58.675 144.795 58.965 145.025 ;
        RECT 58.290 144.640 58.430 144.795 ;
        RECT 59.580 144.780 59.900 145.040 ;
        RECT 60.040 144.780 60.360 145.040 ;
        RECT 61.430 144.795 61.720 145.025 ;
        RECT 61.895 144.980 62.185 145.025 ;
        RECT 62.340 144.980 62.660 145.040 ;
        RECT 63.720 144.980 64.040 145.040 ;
        RECT 61.895 144.840 62.660 144.980 ;
        RECT 61.895 144.795 62.185 144.840 ;
        RECT 61.505 144.640 61.645 144.795 ;
        RECT 62.340 144.780 62.660 144.840 ;
        RECT 62.890 144.840 64.040 144.980 ;
        RECT 62.890 144.640 63.030 144.840 ;
        RECT 63.720 144.780 64.040 144.840 ;
        RECT 64.180 144.980 64.500 145.040 ;
        RECT 64.730 144.980 64.870 145.135 ;
        RECT 66.480 145.120 66.800 145.180 ;
        RECT 70.160 145.120 70.480 145.180 ;
        RECT 70.620 145.320 70.940 145.380 ;
        RECT 81.215 145.320 81.505 145.365 ;
        RECT 70.620 145.180 81.505 145.320 ;
        RECT 70.620 145.120 70.940 145.180 ;
        RECT 81.215 145.135 81.505 145.180 ;
        RECT 83.040 145.320 83.360 145.380 ;
        RECT 89.480 145.320 89.800 145.380 ;
        RECT 83.040 145.180 89.800 145.320 ;
        RECT 83.040 145.120 83.360 145.180 ;
        RECT 89.480 145.120 89.800 145.180 ;
        RECT 64.180 144.840 64.870 144.980 ;
        RECT 64.180 144.780 64.500 144.840 ;
        RECT 66.035 144.795 66.325 145.025 ;
        RECT 66.940 144.980 67.260 145.040 ;
        RECT 69.240 144.980 69.560 145.040 ;
        RECT 66.940 144.840 69.560 144.980 ;
        RECT 58.290 144.500 63.030 144.640 ;
        RECT 63.260 144.640 63.580 144.700 ;
        RECT 65.115 144.640 65.405 144.685 ;
        RECT 63.260 144.500 65.405 144.640 ;
        RECT 66.110 144.640 66.250 144.795 ;
        RECT 66.940 144.780 67.260 144.840 ;
        RECT 69.240 144.780 69.560 144.840 ;
        RECT 69.715 144.980 70.005 145.025 ;
        RECT 72.920 144.980 73.240 145.040 ;
        RECT 69.715 144.840 73.240 144.980 ;
        RECT 69.715 144.795 70.005 144.840 ;
        RECT 72.920 144.780 73.240 144.840 ;
        RECT 79.375 144.980 79.665 145.025 ;
        RECT 87.180 144.980 87.500 145.040 ;
        RECT 79.375 144.840 87.500 144.980 ;
        RECT 79.375 144.795 79.665 144.840 ;
        RECT 87.180 144.780 87.500 144.840 ;
        RECT 87.640 144.980 87.960 145.040 ;
        RECT 94.170 144.980 94.310 145.520 ;
        RECT 105.120 145.460 105.440 145.520 ;
        RECT 106.040 145.460 106.360 145.720 ;
        RECT 107.420 145.660 107.740 145.720 ;
        RECT 121.695 145.660 121.985 145.705 ;
        RECT 106.590 145.520 107.740 145.660 ;
        RECT 94.540 145.320 94.860 145.380 ;
        RECT 103.280 145.320 103.600 145.380 ;
        RECT 106.590 145.320 106.730 145.520 ;
        RECT 107.420 145.460 107.740 145.520 ;
        RECT 117.170 145.520 121.985 145.660 ;
        RECT 117.170 145.320 117.310 145.520 ;
        RECT 121.695 145.475 121.985 145.520 ;
        RECT 122.140 145.660 122.460 145.720 ;
        RECT 122.615 145.660 122.905 145.705 ;
        RECT 122.140 145.520 122.905 145.660 ;
        RECT 122.140 145.460 122.460 145.520 ;
        RECT 122.615 145.475 122.905 145.520 ;
        RECT 94.540 145.180 103.600 145.320 ;
        RECT 94.540 145.120 94.860 145.180 ;
        RECT 103.280 145.120 103.600 145.180 ;
        RECT 104.290 145.180 106.730 145.320 ;
        RECT 107.510 145.180 117.310 145.320 ;
        RECT 121.145 145.320 121.435 145.365 ;
        RECT 121.145 145.180 123.750 145.320 ;
        RECT 87.640 144.840 94.310 144.980 ;
        RECT 96.840 144.980 97.160 145.040 ;
        RECT 99.155 144.980 99.445 145.025 ;
        RECT 96.840 144.840 99.445 144.980 ;
        RECT 87.640 144.780 87.960 144.840 ;
        RECT 96.840 144.780 97.160 144.840 ;
        RECT 99.155 144.795 99.445 144.840 ;
        RECT 99.615 144.795 99.905 145.025 ;
        RECT 100.535 144.795 100.825 145.025 ;
        RECT 67.860 144.640 68.180 144.700 ;
        RECT 72.000 144.640 72.320 144.700 ;
        RECT 66.110 144.500 72.320 144.640 ;
        RECT 63.260 144.440 63.580 144.500 ;
        RECT 65.115 144.455 65.405 144.500 ;
        RECT 65.190 144.300 65.330 144.455 ;
        RECT 67.860 144.440 68.180 144.500 ;
        RECT 72.000 144.440 72.320 144.500 ;
        RECT 73.380 144.640 73.700 144.700 ;
        RECT 78.440 144.640 78.760 144.700 ;
        RECT 73.380 144.500 78.760 144.640 ;
        RECT 73.380 144.440 73.700 144.500 ;
        RECT 78.440 144.440 78.760 144.500 ;
        RECT 89.480 144.640 89.800 144.700 ;
        RECT 96.380 144.640 96.700 144.700 ;
        RECT 89.480 144.500 96.700 144.640 ;
        RECT 89.480 144.440 89.800 144.500 ;
        RECT 96.380 144.440 96.700 144.500 ;
        RECT 97.300 144.640 97.620 144.700 ;
        RECT 99.690 144.640 99.830 144.795 ;
        RECT 97.300 144.500 99.830 144.640 ;
        RECT 97.300 144.440 97.620 144.500 ;
        RECT 100.060 144.440 100.380 144.700 ;
        RECT 100.610 144.640 100.750 144.795 ;
        RECT 100.980 144.780 101.300 145.040 ;
        RECT 102.375 144.980 102.665 145.025 ;
        RECT 103.740 144.980 104.060 145.040 ;
        RECT 104.290 145.025 104.430 145.180 ;
        RECT 102.375 144.840 104.060 144.980 ;
        RECT 102.375 144.795 102.665 144.840 ;
        RECT 103.740 144.780 104.060 144.840 ;
        RECT 104.215 144.795 104.505 145.025 ;
        RECT 107.510 144.700 107.650 145.180 ;
        RECT 121.145 145.135 121.435 145.180 ;
        RECT 109.720 144.780 110.040 145.040 ;
        RECT 110.180 144.980 110.500 145.040 ;
        RECT 110.180 144.780 110.640 144.980 ;
        RECT 119.840 144.780 120.160 145.040 ;
        RECT 120.315 144.795 120.605 145.025 ;
        RECT 121.680 144.980 122.000 145.040 ;
        RECT 122.155 144.980 122.445 145.025 ;
        RECT 121.680 144.840 122.445 144.980 ;
        RECT 101.440 144.640 101.760 144.700 ;
        RECT 100.610 144.500 101.760 144.640 ;
        RECT 101.440 144.440 101.760 144.500 ;
        RECT 102.820 144.440 103.140 144.700 ;
        RECT 105.120 144.640 105.440 144.700 ;
        RECT 106.500 144.640 106.820 144.700 ;
        RECT 105.120 144.500 106.820 144.640 ;
        RECT 105.120 144.440 105.440 144.500 ;
        RECT 106.500 144.440 106.820 144.500 ;
        RECT 106.960 144.440 107.280 144.700 ;
        RECT 107.420 144.440 107.740 144.700 ;
        RECT 109.275 144.640 109.565 144.685 ;
        RECT 110.500 144.640 110.640 144.780 ;
        RECT 116.620 144.640 116.940 144.700 ;
        RECT 120.390 144.640 120.530 144.795 ;
        RECT 121.680 144.780 122.000 144.840 ;
        RECT 122.155 144.795 122.445 144.840 ;
        RECT 109.275 144.500 116.390 144.640 ;
        RECT 109.275 144.455 109.565 144.500 ;
        RECT 66.020 144.300 66.340 144.360 ;
        RECT 65.190 144.160 66.340 144.300 ;
        RECT 66.020 144.100 66.340 144.160 ;
        RECT 69.240 144.300 69.560 144.360 ;
        RECT 74.760 144.300 75.080 144.360 ;
        RECT 69.240 144.160 75.080 144.300 ;
        RECT 69.240 144.100 69.560 144.160 ;
        RECT 74.760 144.100 75.080 144.160 ;
        RECT 75.220 144.300 75.540 144.360 ;
        RECT 97.760 144.300 98.080 144.360 ;
        RECT 110.195 144.300 110.485 144.345 ;
        RECT 75.220 144.160 96.840 144.300 ;
        RECT 75.220 144.100 75.540 144.160 ;
        RECT 61.880 143.960 62.200 144.020 ;
        RECT 62.815 143.960 63.105 144.005 ;
        RECT 61.880 143.820 63.105 143.960 ;
        RECT 61.880 143.760 62.200 143.820 ;
        RECT 62.815 143.775 63.105 143.820 ;
        RECT 63.735 143.960 64.025 144.005 ;
        RECT 64.180 143.960 64.500 144.020 ;
        RECT 63.735 143.820 64.500 143.960 ;
        RECT 63.735 143.775 64.025 143.820 ;
        RECT 64.180 143.760 64.500 143.820 ;
        RECT 65.560 143.960 65.880 144.020 ;
        RECT 66.480 143.960 66.800 144.020 ;
        RECT 65.560 143.820 66.800 143.960 ;
        RECT 65.560 143.760 65.880 143.820 ;
        RECT 66.480 143.760 66.800 143.820 ;
        RECT 66.940 143.760 67.260 144.020 ;
        RECT 72.920 143.960 73.240 144.020 ;
        RECT 77.060 143.960 77.380 144.020 ;
        RECT 86.260 143.960 86.580 144.020 ;
        RECT 72.920 143.820 86.580 143.960 ;
        RECT 72.920 143.760 73.240 143.820 ;
        RECT 77.060 143.760 77.380 143.820 ;
        RECT 86.260 143.760 86.580 143.820 ;
        RECT 92.700 143.760 93.020 144.020 ;
        RECT 96.700 143.960 96.840 144.160 ;
        RECT 97.760 144.160 110.485 144.300 ;
        RECT 116.250 144.300 116.390 144.500 ;
        RECT 116.620 144.500 120.530 144.640 ;
        RECT 116.620 144.440 116.940 144.500 ;
        RECT 123.610 144.300 123.750 145.180 ;
        RECT 116.250 144.160 123.750 144.300 ;
        RECT 97.760 144.100 98.080 144.160 ;
        RECT 110.195 144.115 110.485 144.160 ;
        RECT 102.360 143.960 102.680 144.020 ;
        RECT 109.720 143.960 110.040 144.020 ;
        RECT 96.700 143.820 110.040 143.960 ;
        RECT 102.360 143.760 102.680 143.820 ;
        RECT 109.720 143.760 110.040 143.820 ;
        RECT 112.480 143.760 112.800 144.020 ;
        RECT 53.990 143.140 125.290 143.620 ;
        RECT 60.500 142.940 60.820 143.000 ;
        RECT 61.435 142.940 61.725 142.985 ;
        RECT 73.380 142.940 73.700 143.000 ;
        RECT 60.500 142.800 61.725 142.940 ;
        RECT 60.500 142.740 60.820 142.800 ;
        RECT 61.435 142.755 61.725 142.800 ;
        RECT 66.570 142.800 73.700 142.940 ;
        RECT 53.600 142.600 53.920 142.660 ;
        RECT 58.675 142.600 58.965 142.645 ;
        RECT 53.600 142.460 58.965 142.600 ;
        RECT 53.600 142.400 53.920 142.460 ;
        RECT 58.675 142.415 58.965 142.460 ;
        RECT 62.355 142.260 62.645 142.305 ;
        RECT 65.560 142.260 65.880 142.320 ;
        RECT 66.570 142.260 66.710 142.800 ;
        RECT 73.380 142.740 73.700 142.800 ;
        RECT 73.840 142.940 74.160 143.000 ;
        RECT 75.680 142.940 76.000 143.000 ;
        RECT 73.840 142.800 76.000 142.940 ;
        RECT 73.840 142.740 74.160 142.800 ;
        RECT 75.680 142.740 76.000 142.800 ;
        RECT 76.615 142.940 76.905 142.985 ;
        RECT 112.020 142.940 112.340 143.000 ;
        RECT 76.615 142.800 112.340 142.940 ;
        RECT 76.615 142.755 76.905 142.800 ;
        RECT 112.020 142.740 112.340 142.800 ;
        RECT 67.400 142.400 67.720 142.660 ;
        RECT 69.240 142.600 69.560 142.660 ;
        RECT 82.580 142.600 82.900 142.660 ;
        RECT 69.240 142.460 82.900 142.600 ;
        RECT 69.240 142.400 69.560 142.460 ;
        RECT 82.580 142.400 82.900 142.460 ;
        RECT 85.815 142.600 86.105 142.645 ;
        RECT 87.180 142.600 87.500 142.660 ;
        RECT 85.815 142.460 87.500 142.600 ;
        RECT 85.815 142.415 86.105 142.460 ;
        RECT 87.180 142.400 87.500 142.460 ;
        RECT 94.540 142.400 94.860 142.660 ;
        RECT 95.000 142.600 95.320 142.660 ;
        RECT 114.335 142.600 114.625 142.645 ;
        RECT 95.000 142.460 114.625 142.600 ;
        RECT 95.000 142.400 95.320 142.460 ;
        RECT 114.335 142.415 114.625 142.460 ;
        RECT 115.700 142.600 116.020 142.660 ;
        RECT 123.075 142.600 123.365 142.645 ;
        RECT 115.700 142.460 123.365 142.600 ;
        RECT 115.700 142.400 116.020 142.460 ;
        RECT 123.075 142.415 123.365 142.460 ;
        RECT 57.830 142.120 62.645 142.260 ;
        RECT 57.830 141.980 57.970 142.120 ;
        RECT 62.355 142.075 62.645 142.120 ;
        RECT 63.350 142.120 65.880 142.260 ;
        RECT 56.375 141.920 56.665 141.965 ;
        RECT 57.740 141.920 58.060 141.980 ;
        RECT 56.375 141.780 58.060 141.920 ;
        RECT 56.375 141.735 56.665 141.780 ;
        RECT 57.740 141.720 58.060 141.780 ;
        RECT 59.580 141.720 59.900 141.980 ;
        RECT 60.960 141.720 61.280 141.980 ;
        RECT 61.420 141.920 61.740 141.980 ;
        RECT 63.350 141.965 63.490 142.120 ;
        RECT 65.560 142.060 65.880 142.120 ;
        RECT 66.110 142.120 66.710 142.260 ;
        RECT 67.860 142.260 68.180 142.320 ;
        RECT 81.200 142.260 81.520 142.320 ;
        RECT 94.630 142.260 94.770 142.400 ;
        RECT 67.860 142.120 81.520 142.260 ;
        RECT 66.110 141.965 66.250 142.120 ;
        RECT 67.860 142.060 68.180 142.120 ;
        RECT 81.200 142.060 81.520 142.120 ;
        RECT 93.710 142.120 94.770 142.260 ;
        RECT 96.395 142.260 96.685 142.305 ;
        RECT 108.800 142.260 109.120 142.320 ;
        RECT 96.395 142.120 109.120 142.260 ;
        RECT 61.895 141.920 62.185 141.965 ;
        RECT 61.420 141.780 62.185 141.920 ;
        RECT 61.420 141.720 61.740 141.780 ;
        RECT 61.895 141.735 62.185 141.780 ;
        RECT 63.275 141.735 63.565 141.965 ;
        RECT 64.655 141.920 64.945 141.965 ;
        RECT 63.810 141.780 64.945 141.920 ;
        RECT 62.340 141.580 62.660 141.640 ;
        RECT 63.810 141.580 63.950 141.780 ;
        RECT 64.655 141.735 64.945 141.780 ;
        RECT 66.035 141.735 66.325 141.965 ;
        RECT 66.495 141.920 66.785 141.965 ;
        RECT 66.495 141.780 68.090 141.920 ;
        RECT 66.495 141.735 66.785 141.780 ;
        RECT 62.340 141.440 63.950 141.580 ;
        RECT 64.195 141.580 64.485 141.625 ;
        RECT 67.400 141.580 67.720 141.640 ;
        RECT 64.195 141.440 67.720 141.580 ;
        RECT 67.950 141.580 68.090 141.780 ;
        RECT 68.320 141.720 68.640 141.980 ;
        RECT 68.795 141.920 69.085 141.965 ;
        RECT 69.700 141.920 70.020 141.980 ;
        RECT 68.795 141.780 70.020 141.920 ;
        RECT 68.795 141.735 69.085 141.780 ;
        RECT 69.700 141.720 70.020 141.780 ;
        RECT 70.160 141.720 70.480 141.980 ;
        RECT 90.400 141.920 90.720 141.980 ;
        RECT 70.710 141.780 90.720 141.920 ;
        RECT 70.710 141.580 70.850 141.780 ;
        RECT 90.400 141.720 90.720 141.780 ;
        RECT 91.320 141.920 91.640 141.980 ;
        RECT 93.175 141.920 93.465 141.965 ;
        RECT 93.710 141.920 93.850 142.120 ;
        RECT 96.395 142.075 96.685 142.120 ;
        RECT 108.800 142.060 109.120 142.120 ;
        RECT 91.320 141.780 93.850 141.920 ;
        RECT 91.320 141.720 91.640 141.780 ;
        RECT 93.175 141.735 93.465 141.780 ;
        RECT 94.080 141.720 94.400 141.980 ;
        RECT 94.540 141.720 94.860 141.980 ;
        RECT 95.475 141.735 95.765 141.965 ;
        RECT 95.920 141.920 96.240 141.980 ;
        RECT 97.315 141.920 97.605 141.965 ;
        RECT 95.920 141.780 97.605 141.920 ;
        RECT 67.950 141.440 70.850 141.580 ;
        RECT 72.015 141.580 72.305 141.625 ;
        RECT 74.300 141.580 74.620 141.640 ;
        RECT 72.015 141.440 74.620 141.580 ;
        RECT 62.340 141.380 62.660 141.440 ;
        RECT 64.195 141.395 64.485 141.440 ;
        RECT 67.400 141.380 67.720 141.440 ;
        RECT 72.015 141.395 72.305 141.440 ;
        RECT 74.300 141.380 74.620 141.440 ;
        RECT 74.760 141.580 75.080 141.640 ;
        RECT 82.580 141.580 82.900 141.640 ;
        RECT 74.760 141.440 82.900 141.580 ;
        RECT 74.760 141.380 75.080 141.440 ;
        RECT 82.580 141.380 82.900 141.440 ;
        RECT 83.040 141.380 83.360 141.640 ;
        RECT 89.480 141.580 89.800 141.640 ;
        RECT 92.255 141.580 92.545 141.625 ;
        RECT 89.480 141.440 92.545 141.580 ;
        RECT 89.480 141.380 89.800 141.440 ;
        RECT 92.255 141.395 92.545 141.440 ;
        RECT 57.295 141.240 57.585 141.285 ;
        RECT 58.200 141.240 58.520 141.300 ;
        RECT 57.295 141.100 58.520 141.240 ;
        RECT 57.295 141.055 57.585 141.100 ;
        RECT 58.200 141.040 58.520 141.100 ;
        RECT 61.420 141.240 61.740 141.300 ;
        RECT 62.800 141.240 63.120 141.300 ;
        RECT 61.420 141.100 63.120 141.240 ;
        RECT 61.420 141.040 61.740 141.100 ;
        RECT 62.800 141.040 63.120 141.100 ;
        RECT 63.260 141.240 63.580 141.300 ;
        RECT 64.655 141.240 64.945 141.285 ;
        RECT 63.260 141.100 64.945 141.240 ;
        RECT 63.260 141.040 63.580 141.100 ;
        RECT 64.655 141.055 64.945 141.100 ;
        RECT 65.575 141.240 65.865 141.285 ;
        RECT 68.320 141.240 68.640 141.300 ;
        RECT 65.575 141.100 68.640 141.240 ;
        RECT 65.575 141.055 65.865 141.100 ;
        RECT 68.320 141.040 68.640 141.100 ;
        RECT 69.255 141.240 69.545 141.285 ;
        RECT 69.700 141.240 70.020 141.300 ;
        RECT 69.255 141.100 70.020 141.240 ;
        RECT 69.255 141.055 69.545 141.100 ;
        RECT 69.700 141.040 70.020 141.100 ;
        RECT 71.095 141.240 71.385 141.285 ;
        RECT 77.520 141.240 77.840 141.300 ;
        RECT 71.095 141.100 77.840 141.240 ;
        RECT 71.095 141.055 71.385 141.100 ;
        RECT 77.520 141.040 77.840 141.100 ;
        RECT 81.660 141.240 81.980 141.300 ;
        RECT 95.550 141.240 95.690 141.735 ;
        RECT 95.920 141.720 96.240 141.780 ;
        RECT 97.315 141.735 97.605 141.780 ;
        RECT 98.235 141.920 98.525 141.965 ;
        RECT 99.140 141.920 99.460 141.980 ;
        RECT 117.095 141.920 117.385 141.965 ;
        RECT 117.540 141.920 117.860 141.980 ;
        RECT 98.235 141.780 108.570 141.920 ;
        RECT 98.235 141.735 98.525 141.780 ;
        RECT 99.140 141.720 99.460 141.780 ;
        RECT 96.380 141.580 96.700 141.640 ;
        RECT 98.695 141.580 98.985 141.625 ;
        RECT 107.895 141.580 108.185 141.625 ;
        RECT 96.380 141.440 98.985 141.580 ;
        RECT 96.380 141.380 96.700 141.440 ;
        RECT 98.695 141.395 98.985 141.440 ;
        RECT 99.230 141.440 108.185 141.580 ;
        RECT 108.430 141.580 108.570 141.780 ;
        RECT 117.095 141.780 117.860 141.920 ;
        RECT 117.095 141.735 117.385 141.780 ;
        RECT 117.170 141.580 117.310 141.735 ;
        RECT 117.540 141.720 117.860 141.780 ;
        RECT 118.460 141.920 118.780 141.980 ;
        RECT 118.935 141.920 119.225 141.965 ;
        RECT 118.460 141.780 119.225 141.920 ;
        RECT 118.460 141.720 118.780 141.780 ;
        RECT 118.935 141.735 119.225 141.780 ;
        RECT 119.380 141.920 119.700 141.980 ;
        RECT 121.235 141.920 121.525 141.965 ;
        RECT 122.155 141.920 122.445 141.965 ;
        RECT 119.380 141.780 121.525 141.920 ;
        RECT 119.380 141.720 119.700 141.780 ;
        RECT 121.235 141.735 121.525 141.780 ;
        RECT 121.770 141.780 122.445 141.920 ;
        RECT 108.430 141.440 117.310 141.580 ;
        RECT 81.660 141.100 95.690 141.240 ;
        RECT 97.300 141.240 97.620 141.300 ;
        RECT 97.775 141.240 98.065 141.285 ;
        RECT 97.300 141.100 98.065 141.240 ;
        RECT 81.660 141.040 81.980 141.100 ;
        RECT 97.300 141.040 97.620 141.100 ;
        RECT 97.775 141.055 98.065 141.100 ;
        RECT 98.220 141.240 98.540 141.300 ;
        RECT 99.230 141.240 99.370 141.440 ;
        RECT 107.895 141.395 108.185 141.440 ;
        RECT 120.300 141.380 120.620 141.640 ;
        RECT 98.220 141.100 99.370 141.240 ;
        RECT 99.600 141.240 99.920 141.300 ;
        RECT 105.135 141.240 105.425 141.285 ;
        RECT 99.600 141.100 105.425 141.240 ;
        RECT 98.220 141.040 98.540 141.100 ;
        RECT 99.600 141.040 99.920 141.100 ;
        RECT 105.135 141.055 105.425 141.100 ;
        RECT 118.015 141.240 118.305 141.285 ;
        RECT 121.770 141.240 121.910 141.780 ;
        RECT 122.155 141.735 122.445 141.780 ;
        RECT 118.015 141.100 121.910 141.240 ;
        RECT 118.015 141.055 118.305 141.100 ;
        RECT 53.990 140.420 125.290 140.900 ;
        RECT 58.215 140.220 58.505 140.265 ;
        RECT 58.660 140.220 58.980 140.280 ;
        RECT 58.215 140.080 58.980 140.220 ;
        RECT 58.215 140.035 58.505 140.080 ;
        RECT 58.660 140.020 58.980 140.080 ;
        RECT 59.120 140.220 59.440 140.280 ;
        RECT 59.595 140.220 59.885 140.265 ;
        RECT 59.120 140.080 59.885 140.220 ;
        RECT 59.120 140.020 59.440 140.080 ;
        RECT 59.595 140.035 59.885 140.080 ;
        RECT 66.495 140.220 66.785 140.265 ;
        RECT 67.860 140.220 68.180 140.280 ;
        RECT 66.495 140.080 68.180 140.220 ;
        RECT 66.495 140.035 66.785 140.080 ;
        RECT 67.860 140.020 68.180 140.080 ;
        RECT 71.540 140.220 71.860 140.280 ;
        RECT 71.540 140.080 73.610 140.220 ;
        RECT 71.540 140.020 71.860 140.080 ;
        RECT 56.820 139.340 57.140 139.600 ;
        RECT 58.750 139.585 58.890 140.020 ;
        RECT 60.500 139.880 60.820 139.940 ;
        RECT 61.895 139.880 62.185 139.925 ;
        RECT 60.500 139.740 62.185 139.880 ;
        RECT 60.500 139.680 60.820 139.740 ;
        RECT 61.895 139.695 62.185 139.740 ;
        RECT 63.260 139.880 63.580 139.940 ;
        RECT 63.260 139.740 64.410 139.880 ;
        RECT 63.260 139.680 63.580 139.740 ;
        RECT 58.675 139.355 58.965 139.585 ;
        RECT 60.960 139.340 61.280 139.600 ;
        RECT 61.420 139.340 61.740 139.600 ;
        RECT 62.340 139.585 62.660 139.600 ;
        RECT 62.340 139.540 62.875 139.585 ;
        RECT 63.735 139.540 64.025 139.585 ;
        RECT 62.340 139.400 64.025 139.540 ;
        RECT 64.270 139.540 64.410 139.740 ;
        RECT 67.400 139.680 67.720 139.940 ;
        RECT 73.470 139.925 73.610 140.080 ;
        RECT 75.220 140.020 75.540 140.280 ;
        RECT 76.600 140.020 76.920 140.280 ;
        RECT 77.060 140.220 77.380 140.280 ;
        RECT 83.975 140.220 84.265 140.265 ;
        RECT 84.880 140.220 85.200 140.280 ;
        RECT 91.320 140.220 91.640 140.280 ;
        RECT 77.060 140.080 83.730 140.220 ;
        RECT 77.060 140.020 77.380 140.080 ;
        RECT 67.990 139.740 73.150 139.880 ;
        RECT 64.655 139.540 64.945 139.585 ;
        RECT 64.270 139.400 64.945 139.540 ;
        RECT 62.340 139.355 62.875 139.400 ;
        RECT 63.735 139.355 64.025 139.400 ;
        RECT 64.655 139.355 64.945 139.400 ;
        RECT 66.035 139.540 66.325 139.585 ;
        RECT 67.990 139.540 68.130 139.740 ;
        RECT 68.870 139.585 69.010 139.740 ;
        RECT 73.010 139.600 73.150 139.740 ;
        RECT 73.395 139.695 73.685 139.925 ;
        RECT 74.300 139.880 74.620 139.940 ;
        RECT 83.590 139.880 83.730 140.080 ;
        RECT 83.975 140.080 85.200 140.220 ;
        RECT 83.975 140.035 84.265 140.080 ;
        RECT 84.880 140.020 85.200 140.080 ;
        RECT 85.430 140.080 91.640 140.220 ;
        RECT 85.430 139.880 85.570 140.080 ;
        RECT 91.320 140.020 91.640 140.080 ;
        RECT 92.700 140.220 93.020 140.280 ;
        RECT 104.215 140.220 104.505 140.265 ;
        RECT 105.120 140.220 105.440 140.280 ;
        RECT 92.700 140.080 103.050 140.220 ;
        RECT 92.700 140.020 93.020 140.080 ;
        RECT 88.115 139.880 88.405 139.925 ;
        RECT 89.020 139.880 89.340 139.940 ;
        RECT 74.300 139.740 83.270 139.880 ;
        RECT 83.590 139.740 85.570 139.880 ;
        RECT 74.300 139.680 74.620 139.740 ;
        RECT 66.035 139.400 68.130 139.540 ;
        RECT 66.035 139.355 66.325 139.400 ;
        RECT 68.335 139.355 68.625 139.585 ;
        RECT 68.795 139.355 69.085 139.585 ;
        RECT 69.240 139.540 69.560 139.600 ;
        RECT 69.715 139.540 70.005 139.585 ;
        RECT 69.240 139.400 70.005 139.540 ;
        RECT 62.340 139.340 62.660 139.355 ;
        RECT 60.040 139.000 60.360 139.260 ;
        RECT 63.260 139.000 63.580 139.260 ;
        RECT 64.180 139.200 64.500 139.260 ;
        RECT 65.575 139.200 65.865 139.245 ;
        RECT 64.180 139.060 65.865 139.200 ;
        RECT 64.180 139.000 64.500 139.060 ;
        RECT 65.575 139.015 65.865 139.060 ;
        RECT 67.400 139.200 67.720 139.260 ;
        RECT 68.410 139.200 68.550 139.355 ;
        RECT 69.240 139.340 69.560 139.400 ;
        RECT 69.715 139.355 70.005 139.400 ;
        RECT 70.160 139.340 70.480 139.600 ;
        RECT 70.635 139.540 70.925 139.585 ;
        RECT 70.635 139.400 72.760 139.540 ;
        RECT 70.635 139.355 70.925 139.400 ;
        RECT 67.400 139.060 68.550 139.200 ;
        RECT 65.650 138.860 65.790 139.015 ;
        RECT 67.400 139.000 67.720 139.060 ;
        RECT 70.710 138.860 70.850 139.355 ;
        RECT 72.620 139.200 72.760 139.400 ;
        RECT 72.920 139.340 73.240 139.600 ;
        RECT 73.855 139.355 74.145 139.585 ;
        RECT 73.930 139.200 74.070 139.355 ;
        RECT 74.760 139.340 75.080 139.600 ;
        RECT 75.310 139.585 75.450 139.740 ;
        RECT 75.235 139.355 75.525 139.585 ;
        RECT 76.155 139.540 76.445 139.585 ;
        RECT 77.060 139.540 77.380 139.600 ;
        RECT 76.155 139.400 77.380 139.540 ;
        RECT 76.155 139.355 76.445 139.400 ;
        RECT 77.060 139.340 77.380 139.400 ;
        RECT 77.520 139.340 77.840 139.600 ;
        RECT 77.995 139.540 78.285 139.585 ;
        RECT 79.820 139.540 80.140 139.600 ;
        RECT 77.995 139.400 80.140 139.540 ;
        RECT 77.995 139.355 78.285 139.400 ;
        RECT 79.820 139.340 80.140 139.400 ;
        RECT 80.280 139.540 80.600 139.600 ;
        RECT 80.755 139.540 81.045 139.585 ;
        RECT 80.280 139.400 81.045 139.540 ;
        RECT 80.280 139.340 80.600 139.400 ;
        RECT 80.755 139.355 81.045 139.400 ;
        RECT 81.200 139.340 81.520 139.600 ;
        RECT 83.130 139.585 83.270 139.740 ;
        RECT 83.055 139.355 83.345 139.585 ;
        RECT 84.895 139.540 85.185 139.585 ;
        RECT 85.430 139.540 85.570 139.740 ;
        RECT 86.350 139.740 87.395 139.880 ;
        RECT 84.895 139.400 85.570 139.540 ;
        RECT 84.895 139.355 85.185 139.400 ;
        RECT 85.800 139.340 86.120 139.600 ;
        RECT 86.350 139.585 86.490 139.740 ;
        RECT 86.275 139.355 86.565 139.585 ;
        RECT 86.740 139.305 87.030 139.535 ;
        RECT 76.600 139.200 76.920 139.260 ;
        RECT 72.620 139.060 76.920 139.200 ;
        RECT 76.600 139.000 76.920 139.060 ;
        RECT 78.440 139.000 78.760 139.260 ;
        RECT 78.900 139.000 79.220 139.260 ;
        RECT 65.650 138.720 70.850 138.860 ;
        RECT 71.555 138.860 71.845 138.905 ;
        RECT 75.680 138.860 76.000 138.920 ;
        RECT 86.815 138.860 86.955 139.305 ;
        RECT 71.555 138.720 73.150 138.860 ;
        RECT 71.555 138.675 71.845 138.720 ;
        RECT 55.900 138.320 56.220 138.580 ;
        RECT 67.860 138.520 68.180 138.580 ;
        RECT 72.015 138.520 72.305 138.565 ;
        RECT 67.860 138.380 72.305 138.520 ;
        RECT 73.010 138.520 73.150 138.720 ;
        RECT 75.680 138.720 86.955 138.860 ;
        RECT 75.680 138.660 76.000 138.720 ;
        RECT 74.300 138.520 74.620 138.580 ;
        RECT 73.010 138.380 74.620 138.520 ;
        RECT 67.860 138.320 68.180 138.380 ;
        RECT 72.015 138.335 72.305 138.380 ;
        RECT 74.300 138.320 74.620 138.380 ;
        RECT 78.440 138.520 78.760 138.580 ;
        RECT 83.055 138.520 83.345 138.565 ;
        RECT 87.255 138.520 87.395 139.740 ;
        RECT 88.115 139.740 89.340 139.880 ;
        RECT 88.115 139.695 88.405 139.740 ;
        RECT 89.020 139.680 89.340 139.740 ;
        RECT 94.080 139.880 94.400 139.940 ;
        RECT 102.375 139.880 102.665 139.925 ;
        RECT 94.080 139.740 102.665 139.880 ;
        RECT 102.910 139.880 103.050 140.080 ;
        RECT 104.215 140.080 105.440 140.220 ;
        RECT 104.215 140.035 104.505 140.080 ;
        RECT 105.120 140.020 105.440 140.080 ;
        RECT 106.040 140.220 106.360 140.280 ;
        RECT 112.495 140.220 112.785 140.265 ;
        RECT 106.040 140.080 112.785 140.220 ;
        RECT 106.040 140.020 106.360 140.080 ;
        RECT 112.495 140.035 112.785 140.080 ;
        RECT 116.620 140.220 116.940 140.280 ;
        RECT 120.300 140.220 120.620 140.280 ;
        RECT 116.620 140.080 120.620 140.220 ;
        RECT 116.620 140.020 116.940 140.080 ;
        RECT 120.300 140.020 120.620 140.080 ;
        RECT 122.615 140.220 122.905 140.265 ;
        RECT 125.360 140.220 125.680 140.280 ;
        RECT 122.615 140.080 125.680 140.220 ;
        RECT 122.615 140.035 122.905 140.080 ;
        RECT 125.360 140.020 125.680 140.080 ;
        RECT 107.880 139.880 108.200 139.940 ;
        RECT 102.910 139.740 106.270 139.880 ;
        RECT 94.080 139.680 94.400 139.740 ;
        RECT 102.375 139.695 102.665 139.740 ;
        RECT 88.575 139.540 88.865 139.585 ;
        RECT 91.780 139.540 92.100 139.600 ;
        RECT 88.575 139.400 92.100 139.540 ;
        RECT 88.575 139.355 88.865 139.400 ;
        RECT 91.780 139.340 92.100 139.400 ;
        RECT 97.760 139.340 98.080 139.600 ;
        RECT 98.680 139.340 99.000 139.600 ;
        RECT 99.600 139.340 99.920 139.600 ;
        RECT 100.995 139.540 101.285 139.585 ;
        RECT 103.295 139.540 103.585 139.585 ;
        RECT 100.995 139.400 103.585 139.540 ;
        RECT 100.995 139.355 101.285 139.400 ;
        RECT 103.295 139.355 103.585 139.400 ;
        RECT 104.675 139.540 104.965 139.585 ;
        RECT 105.580 139.540 105.900 139.600 ;
        RECT 106.130 139.585 106.270 139.740 ;
        RECT 107.880 139.740 117.770 139.880 ;
        RECT 107.880 139.680 108.200 139.740 ;
        RECT 104.675 139.400 105.900 139.540 ;
        RECT 104.675 139.355 104.965 139.400 ;
        RECT 96.380 139.200 96.700 139.260 ;
        RECT 98.220 139.200 98.540 139.260 ;
        RECT 96.380 139.060 98.540 139.200 ;
        RECT 96.380 139.000 96.700 139.060 ;
        RECT 98.220 139.000 98.540 139.060 ;
        RECT 99.155 139.015 99.445 139.245 ;
        RECT 100.075 139.015 100.365 139.245 ;
        RECT 92.700 138.860 93.020 138.920 ;
        RECT 98.680 138.860 99.000 138.920 ;
        RECT 99.230 138.860 99.370 139.015 ;
        RECT 92.700 138.720 95.230 138.860 ;
        RECT 92.700 138.660 93.020 138.720 ;
        RECT 78.440 138.380 87.395 138.520 ;
        RECT 90.400 138.520 90.720 138.580 ;
        RECT 94.540 138.520 94.860 138.580 ;
        RECT 90.400 138.380 94.860 138.520 ;
        RECT 95.090 138.520 95.230 138.720 ;
        RECT 98.680 138.720 99.370 138.860 ;
        RECT 99.600 138.860 99.920 138.920 ;
        RECT 100.150 138.860 100.290 139.015 ;
        RECT 99.600 138.720 100.290 138.860 ;
        RECT 98.680 138.660 99.000 138.720 ;
        RECT 99.600 138.660 99.920 138.720 ;
        RECT 104.750 138.520 104.890 139.355 ;
        RECT 105.580 139.340 105.900 139.400 ;
        RECT 106.055 139.355 106.345 139.585 ;
        RECT 106.500 139.540 106.820 139.600 ;
        RECT 115.255 139.540 115.545 139.585 ;
        RECT 106.500 139.400 115.545 139.540 ;
        RECT 106.500 139.340 106.820 139.400 ;
        RECT 115.255 139.355 115.545 139.400 ;
        RECT 116.620 139.340 116.940 139.600 ;
        RECT 117.080 139.340 117.400 139.600 ;
        RECT 117.630 139.585 117.770 139.740 ;
        RECT 118.090 139.740 121.910 139.880 ;
        RECT 118.090 139.585 118.230 139.740 ;
        RECT 121.770 139.600 121.910 139.740 ;
        RECT 117.555 139.355 117.845 139.585 ;
        RECT 118.015 139.355 118.305 139.585 ;
        RECT 120.300 139.340 120.620 139.600 ;
        RECT 121.680 139.340 122.000 139.600 ;
        RECT 123.535 139.540 123.825 139.585 ;
        RECT 123.980 139.540 124.300 139.600 ;
        RECT 123.535 139.400 124.300 139.540 ;
        RECT 123.535 139.355 123.825 139.400 ;
        RECT 123.980 139.340 124.300 139.400 ;
        RECT 114.780 139.200 115.100 139.260 ;
        RECT 119.395 139.200 119.685 139.245 ;
        RECT 121.235 139.200 121.525 139.245 ;
        RECT 114.780 139.060 119.685 139.200 ;
        RECT 114.780 139.000 115.100 139.060 ;
        RECT 119.395 139.015 119.685 139.060 ;
        RECT 119.930 139.060 121.525 139.200 ;
        RECT 117.080 138.860 117.400 138.920 ;
        RECT 119.930 138.860 120.070 139.060 ;
        RECT 121.235 139.015 121.525 139.060 ;
        RECT 117.080 138.720 120.070 138.860 ;
        RECT 117.080 138.660 117.400 138.720 ;
        RECT 120.795 138.675 121.085 138.905 ;
        RECT 95.090 138.380 104.890 138.520 ;
        RECT 116.160 138.520 116.480 138.580 ;
        RECT 120.850 138.520 120.990 138.675 ;
        RECT 116.160 138.380 120.990 138.520 ;
        RECT 78.440 138.320 78.760 138.380 ;
        RECT 83.055 138.335 83.345 138.380 ;
        RECT 90.400 138.320 90.720 138.380 ;
        RECT 94.540 138.320 94.860 138.380 ;
        RECT 116.160 138.320 116.480 138.380 ;
        RECT 53.990 137.700 125.290 138.180 ;
        RECT 60.515 137.500 60.805 137.545 ;
        RECT 60.960 137.500 61.280 137.560 ;
        RECT 60.515 137.360 61.280 137.500 ;
        RECT 60.515 137.315 60.805 137.360 ;
        RECT 60.960 137.300 61.280 137.360 ;
        RECT 65.100 137.500 65.420 137.560 ;
        RECT 65.575 137.500 65.865 137.545 ;
        RECT 65.100 137.360 65.865 137.500 ;
        RECT 65.100 137.300 65.420 137.360 ;
        RECT 65.575 137.315 65.865 137.360 ;
        RECT 66.480 137.500 66.800 137.560 ;
        RECT 67.875 137.500 68.165 137.545 ;
        RECT 66.480 137.360 68.165 137.500 ;
        RECT 66.480 137.300 66.800 137.360 ;
        RECT 67.875 137.315 68.165 137.360 ;
        RECT 69.715 137.500 70.005 137.545 ;
        RECT 80.280 137.500 80.600 137.560 ;
        RECT 69.715 137.360 80.600 137.500 ;
        RECT 69.715 137.315 70.005 137.360 ;
        RECT 80.280 137.300 80.600 137.360 ;
        RECT 85.800 137.500 86.120 137.560 ;
        RECT 88.115 137.500 88.405 137.545 ;
        RECT 85.800 137.360 88.405 137.500 ;
        RECT 85.800 137.300 86.120 137.360 ;
        RECT 88.115 137.315 88.405 137.360 ;
        RECT 90.400 137.500 90.720 137.560 ;
        RECT 95.920 137.500 96.240 137.560 ;
        RECT 116.620 137.500 116.940 137.560 ;
        RECT 90.400 137.360 96.240 137.500 ;
        RECT 90.400 137.300 90.720 137.360 ;
        RECT 95.920 137.300 96.240 137.360 ;
        RECT 101.990 137.360 116.940 137.500 ;
        RECT 61.420 137.160 61.740 137.220 ;
        RECT 67.400 137.160 67.720 137.220 ;
        RECT 69.240 137.160 69.560 137.220 ;
        RECT 72.000 137.160 72.320 137.220 ;
        RECT 61.420 137.020 63.030 137.160 ;
        RECT 61.420 136.960 61.740 137.020 ;
        RECT 58.200 136.620 58.520 136.880 ;
        RECT 62.340 136.820 62.660 136.880 ;
        RECT 62.200 136.620 62.660 136.820 ;
        RECT 57.295 136.345 57.585 136.575 ;
        RECT 57.740 136.480 58.060 136.540 ;
        RECT 59.595 136.480 59.885 136.525 ;
        RECT 57.370 136.200 57.510 136.345 ;
        RECT 57.740 136.340 59.885 136.480 ;
        RECT 57.740 136.280 58.060 136.340 ;
        RECT 59.595 136.295 59.885 136.340 ;
        RECT 60.960 136.280 61.280 136.540 ;
        RECT 61.765 136.480 62.055 136.525 ;
        RECT 62.200 136.480 62.340 136.620 ;
        RECT 62.890 136.525 63.030 137.020 ;
        RECT 67.400 137.020 69.560 137.160 ;
        RECT 67.400 136.960 67.720 137.020 ;
        RECT 69.240 136.960 69.560 137.020 ;
        RECT 70.250 137.020 72.320 137.160 ;
        RECT 70.250 136.865 70.390 137.020 ;
        RECT 72.000 136.960 72.320 137.020 ;
        RECT 74.760 136.960 75.080 137.220 ;
        RECT 77.995 137.160 78.285 137.205 ;
        RECT 83.040 137.160 83.360 137.220 ;
        RECT 77.995 137.020 83.360 137.160 ;
        RECT 77.995 136.975 78.285 137.020 ;
        RECT 83.040 136.960 83.360 137.020 ;
        RECT 86.260 137.160 86.580 137.220 ;
        RECT 86.260 137.020 90.630 137.160 ;
        RECT 86.260 136.960 86.580 137.020 ;
        RECT 63.350 136.680 69.930 136.820 ;
        RECT 63.350 136.540 63.490 136.680 ;
        RECT 61.765 136.340 62.340 136.480 ;
        RECT 61.765 136.295 62.055 136.340 ;
        RECT 62.815 136.295 63.105 136.525 ;
        RECT 57.280 135.940 57.600 136.200 ;
        RECT 58.660 135.940 58.980 136.200 ;
        RECT 62.350 135.955 62.640 136.185 ;
        RECT 62.890 136.140 63.030 136.295 ;
        RECT 63.260 136.280 63.580 136.540 ;
        RECT 64.180 136.280 64.500 136.540 ;
        RECT 66.480 136.280 66.800 136.540 ;
        RECT 67.415 136.295 67.705 136.525 ;
        RECT 68.335 136.295 68.625 136.525 ;
        RECT 68.795 136.480 69.085 136.525 ;
        RECT 69.240 136.480 69.560 136.540 ;
        RECT 68.795 136.340 69.560 136.480 ;
        RECT 69.790 136.480 69.930 136.680 ;
        RECT 70.175 136.635 70.465 136.865 ;
        RECT 74.850 136.820 74.990 136.960 ;
        RECT 72.090 136.680 74.990 136.820 ;
        RECT 77.520 136.820 77.840 136.880 ;
        RECT 80.280 136.820 80.600 136.880 ;
        RECT 77.520 136.680 80.600 136.820 ;
        RECT 70.635 136.480 70.925 136.525 ;
        RECT 69.790 136.340 70.925 136.480 ;
        RECT 68.795 136.295 69.085 136.340 ;
        RECT 64.270 136.140 64.410 136.280 ;
        RECT 62.890 136.000 64.410 136.140 ;
        RECT 65.100 136.140 65.420 136.200 ;
        RECT 67.490 136.140 67.630 136.295 ;
        RECT 65.100 136.000 67.630 136.140 ;
        RECT 68.410 136.140 68.550 136.295 ;
        RECT 69.240 136.280 69.560 136.340 ;
        RECT 70.635 136.295 70.925 136.340 ;
        RECT 71.080 136.480 71.400 136.540 ;
        RECT 72.090 136.525 72.230 136.680 ;
        RECT 77.520 136.620 77.840 136.680 ;
        RECT 80.280 136.620 80.600 136.680 ;
        RECT 85.340 136.820 85.660 136.880 ;
        RECT 90.490 136.865 90.630 137.020 ;
        RECT 89.495 136.820 89.785 136.865 ;
        RECT 85.340 136.680 89.785 136.820 ;
        RECT 85.340 136.620 85.660 136.680 ;
        RECT 89.495 136.635 89.785 136.680 ;
        RECT 90.415 136.635 90.705 136.865 ;
        RECT 98.680 136.820 99.000 136.880 ;
        RECT 90.950 136.680 99.000 136.820 ;
        RECT 71.555 136.480 71.845 136.525 ;
        RECT 71.080 136.340 71.845 136.480 ;
        RECT 71.080 136.280 71.400 136.340 ;
        RECT 71.555 136.295 71.845 136.340 ;
        RECT 72.015 136.295 72.305 136.525 ;
        RECT 72.460 136.280 72.780 136.540 ;
        RECT 73.395 136.480 73.685 136.525 ;
        RECT 74.760 136.480 75.080 136.540 ;
        RECT 73.395 136.340 75.080 136.480 ;
        RECT 73.395 136.295 73.685 136.340 ;
        RECT 74.760 136.280 75.080 136.340 ;
        RECT 75.235 136.480 75.525 136.525 ;
        RECT 75.680 136.480 76.000 136.540 ;
        RECT 75.235 136.340 76.000 136.480 ;
        RECT 75.235 136.295 75.525 136.340 ;
        RECT 75.680 136.280 76.000 136.340 ;
        RECT 77.075 136.480 77.365 136.525 ;
        RECT 79.360 136.480 79.680 136.540 ;
        RECT 77.075 136.340 79.680 136.480 ;
        RECT 77.075 136.295 77.365 136.340 ;
        RECT 79.360 136.280 79.680 136.340 ;
        RECT 81.200 136.480 81.520 136.540 ;
        RECT 83.500 136.480 83.820 136.540 ;
        RECT 89.035 136.480 89.325 136.525 ;
        RECT 81.200 136.340 83.820 136.480 ;
        RECT 81.200 136.280 81.520 136.340 ;
        RECT 83.500 136.280 83.820 136.340 ;
        RECT 84.050 136.340 89.325 136.480 ;
        RECT 76.155 136.140 76.445 136.185 ;
        RECT 68.410 136.000 76.445 136.140 ;
        RECT 56.375 135.800 56.665 135.845 ;
        RECT 62.430 135.800 62.570 135.955 ;
        RECT 65.100 135.940 65.420 136.000 ;
        RECT 76.155 135.955 76.445 136.000 ;
        RECT 76.600 136.140 76.920 136.200 ;
        RECT 84.050 136.140 84.190 136.340 ;
        RECT 89.035 136.295 89.325 136.340 ;
        RECT 89.955 136.480 90.245 136.525 ;
        RECT 90.950 136.480 91.090 136.680 ;
        RECT 98.680 136.620 99.000 136.680 ;
        RECT 89.955 136.340 91.090 136.480 ;
        RECT 91.320 136.480 91.640 136.540 ;
        RECT 97.760 136.480 98.080 136.540 ;
        RECT 101.990 136.525 102.130 137.360 ;
        RECT 116.620 137.300 116.940 137.360 ;
        RECT 122.155 137.500 122.445 137.545 ;
        RECT 123.060 137.500 123.380 137.560 ;
        RECT 122.155 137.360 123.380 137.500 ;
        RECT 122.155 137.315 122.445 137.360 ;
        RECT 123.060 137.300 123.380 137.360 ;
        RECT 111.575 137.160 111.865 137.205 ;
        RECT 120.760 137.160 121.080 137.220 ;
        RECT 111.575 137.020 121.080 137.160 ;
        RECT 111.575 136.975 111.865 137.020 ;
        RECT 120.760 136.960 121.080 137.020 ;
        RECT 106.500 136.820 106.820 136.880 ;
        RECT 107.880 136.820 108.200 136.880 ;
        RECT 114.780 136.820 115.100 136.880 ;
        RECT 103.830 136.680 106.820 136.820 ;
        RECT 91.320 136.340 98.080 136.480 ;
        RECT 89.955 136.295 90.245 136.340 ;
        RECT 76.600 136.000 84.190 136.140 ;
        RECT 62.800 135.800 63.120 135.860 ;
        RECT 56.375 135.660 63.120 135.800 ;
        RECT 56.375 135.615 56.665 135.660 ;
        RECT 62.800 135.600 63.120 135.660 ;
        RECT 63.260 135.800 63.580 135.860 ;
        RECT 64.195 135.800 64.485 135.845 ;
        RECT 63.260 135.660 64.485 135.800 ;
        RECT 63.260 135.600 63.580 135.660 ;
        RECT 64.195 135.615 64.485 135.660 ;
        RECT 66.480 135.800 66.800 135.860 ;
        RECT 69.240 135.800 69.560 135.860 ;
        RECT 66.480 135.660 69.560 135.800 ;
        RECT 66.480 135.600 66.800 135.660 ;
        RECT 69.240 135.600 69.560 135.660 ;
        RECT 69.700 135.800 70.020 135.860 ;
        RECT 73.840 135.800 74.160 135.860 ;
        RECT 69.700 135.660 74.160 135.800 ;
        RECT 69.700 135.600 70.020 135.660 ;
        RECT 73.840 135.600 74.160 135.660 ;
        RECT 74.315 135.800 74.605 135.845 ;
        RECT 75.680 135.800 76.000 135.860 ;
        RECT 74.315 135.660 76.000 135.800 ;
        RECT 76.230 135.800 76.370 135.955 ;
        RECT 76.600 135.940 76.920 136.000 ;
        RECT 87.195 135.955 87.485 136.185 ;
        RECT 87.640 136.140 87.960 136.200 ;
        RECT 90.030 136.140 90.170 136.295 ;
        RECT 91.320 136.280 91.640 136.340 ;
        RECT 97.760 136.280 98.080 136.340 ;
        RECT 101.915 136.295 102.205 136.525 ;
        RECT 102.375 136.480 102.665 136.525 ;
        RECT 103.830 136.480 103.970 136.680 ;
        RECT 106.500 136.620 106.820 136.680 ;
        RECT 107.050 136.680 108.200 136.820 ;
        RECT 107.050 136.525 107.190 136.680 ;
        RECT 107.880 136.620 108.200 136.680 ;
        RECT 108.430 136.680 115.100 136.820 ;
        RECT 102.375 136.340 103.970 136.480 ;
        RECT 102.375 136.295 102.665 136.340 ;
        RECT 106.975 136.295 107.265 136.525 ;
        RECT 107.420 136.280 107.740 136.540 ;
        RECT 108.430 136.525 108.570 136.680 ;
        RECT 114.780 136.620 115.100 136.680 ;
        RECT 108.355 136.295 108.645 136.525 ;
        RECT 108.800 136.280 109.120 136.540 ;
        RECT 118.460 136.280 118.780 136.540 ;
        RECT 118.920 136.480 119.240 136.540 ;
        RECT 120.775 136.480 121.065 136.525 ;
        RECT 118.920 136.340 121.065 136.480 ;
        RECT 118.920 136.280 119.240 136.340 ;
        RECT 120.775 136.295 121.065 136.340 ;
        RECT 121.220 136.280 121.540 136.540 ;
        RECT 122.600 136.280 122.920 136.540 ;
        RECT 87.640 136.000 90.170 136.140 ;
        RECT 77.060 135.800 77.380 135.860 ;
        RECT 79.820 135.800 80.140 135.860 ;
        RECT 76.230 135.660 80.140 135.800 ;
        RECT 74.315 135.615 74.605 135.660 ;
        RECT 75.680 135.600 76.000 135.660 ;
        RECT 77.060 135.600 77.380 135.660 ;
        RECT 79.820 135.600 80.140 135.660 ;
        RECT 80.280 135.800 80.600 135.860 ;
        RECT 80.755 135.800 81.045 135.845 ;
        RECT 82.120 135.800 82.440 135.860 ;
        RECT 80.280 135.660 82.440 135.800 ;
        RECT 80.280 135.600 80.600 135.660 ;
        RECT 80.755 135.615 81.045 135.660 ;
        RECT 82.120 135.600 82.440 135.660 ;
        RECT 82.580 135.800 82.900 135.860 ;
        RECT 85.800 135.800 86.120 135.860 ;
        RECT 82.580 135.660 86.120 135.800 ;
        RECT 87.270 135.800 87.410 135.955 ;
        RECT 87.640 135.940 87.960 136.000 ;
        RECT 93.175 135.955 93.465 136.185 ;
        RECT 102.450 136.000 103.970 136.140 ;
        RECT 93.250 135.800 93.390 135.955 ;
        RECT 102.450 135.860 102.590 136.000 ;
        RECT 100.060 135.800 100.380 135.860 ;
        RECT 87.270 135.660 100.380 135.800 ;
        RECT 82.580 135.600 82.900 135.660 ;
        RECT 85.800 135.600 86.120 135.660 ;
        RECT 100.060 135.600 100.380 135.660 ;
        RECT 102.360 135.600 102.680 135.860 ;
        RECT 103.280 135.600 103.600 135.860 ;
        RECT 103.830 135.845 103.970 136.000 ;
        RECT 104.200 135.940 104.520 136.200 ;
        RECT 105.135 136.140 105.425 136.185 ;
        RECT 105.135 136.000 110.640 136.140 ;
        RECT 105.135 135.955 105.425 136.000 ;
        RECT 103.755 135.615 104.045 135.845 ;
        RECT 104.660 135.800 104.980 135.860 ;
        RECT 106.055 135.800 106.345 135.845 ;
        RECT 104.660 135.660 106.345 135.800 ;
        RECT 110.500 135.800 110.640 136.000 ;
        RECT 118.000 135.940 118.320 136.200 ;
        RECT 118.550 136.140 118.690 136.280 ;
        RECT 118.550 136.000 119.150 136.140 ;
        RECT 118.460 135.800 118.780 135.860 ;
        RECT 119.010 135.845 119.150 136.000 ;
        RECT 110.500 135.660 118.780 135.800 ;
        RECT 104.660 135.600 104.980 135.660 ;
        RECT 106.055 135.615 106.345 135.660 ;
        RECT 118.460 135.600 118.780 135.660 ;
        RECT 118.935 135.615 119.225 135.845 ;
        RECT 123.060 135.600 123.380 135.860 ;
        RECT 53.990 134.980 125.290 135.460 ;
        RECT 56.820 134.780 57.140 134.840 ;
        RECT 58.675 134.780 58.965 134.825 ;
        RECT 56.820 134.640 58.965 134.780 ;
        RECT 56.820 134.580 57.140 134.640 ;
        RECT 58.675 134.595 58.965 134.640 ;
        RECT 59.120 134.780 59.440 134.840 ;
        RECT 60.515 134.780 60.805 134.825 ;
        RECT 61.420 134.780 61.740 134.840 ;
        RECT 59.120 134.640 61.740 134.780 ;
        RECT 59.120 134.580 59.440 134.640 ;
        RECT 60.515 134.595 60.805 134.640 ;
        RECT 61.420 134.580 61.740 134.640 ;
        RECT 63.720 134.780 64.040 134.840 ;
        RECT 64.655 134.780 64.945 134.825 ;
        RECT 72.920 134.780 73.240 134.840 ;
        RECT 63.720 134.640 64.945 134.780 ;
        RECT 63.720 134.580 64.040 134.640 ;
        RECT 64.655 134.595 64.945 134.640 ;
        RECT 65.650 134.640 69.470 134.780 ;
        RECT 53.140 134.440 53.460 134.500 ;
        RECT 65.650 134.440 65.790 134.640 ;
        RECT 53.140 134.300 57.510 134.440 ;
        RECT 53.140 134.240 53.460 134.300 ;
        RECT 56.820 133.900 57.140 134.160 ;
        RECT 57.370 134.145 57.510 134.300 ;
        RECT 63.810 134.300 65.790 134.440 ;
        RECT 57.295 133.915 57.585 134.145 ;
        RECT 59.595 134.100 59.885 134.145 ;
        RECT 60.500 134.100 60.820 134.160 ;
        RECT 59.595 133.960 60.820 134.100 ;
        RECT 59.595 133.915 59.885 133.960 ;
        RECT 55.900 133.760 56.220 133.820 ;
        RECT 59.670 133.760 59.810 133.915 ;
        RECT 60.500 133.900 60.820 133.960 ;
        RECT 60.975 133.915 61.265 134.145 ;
        RECT 62.815 134.100 63.105 134.145 ;
        RECT 63.260 134.100 63.580 134.160 ;
        RECT 63.810 134.145 63.950 134.300 ;
        RECT 66.480 134.240 66.800 134.500 ;
        RECT 62.815 133.960 63.580 134.100 ;
        RECT 62.815 133.915 63.105 133.960 ;
        RECT 55.900 133.620 59.810 133.760 ;
        RECT 55.900 133.560 56.220 133.620 ;
        RECT 61.050 133.420 61.190 133.915 ;
        RECT 63.260 133.900 63.580 133.960 ;
        RECT 63.735 133.915 64.025 134.145 ;
        RECT 64.195 133.915 64.485 134.145 ;
        RECT 64.640 134.100 64.960 134.160 ;
        RECT 65.575 134.100 65.865 134.145 ;
        RECT 64.640 133.960 65.865 134.100 ;
        RECT 61.420 133.760 61.740 133.820 ;
        RECT 63.810 133.760 63.950 133.915 ;
        RECT 61.420 133.620 63.950 133.760 ;
        RECT 64.270 133.760 64.410 133.915 ;
        RECT 64.640 133.900 64.960 133.960 ;
        RECT 65.575 133.915 65.865 133.960 ;
        RECT 67.400 133.900 67.720 134.160 ;
        RECT 67.860 134.100 68.180 134.160 ;
        RECT 69.330 134.145 69.470 134.640 ;
        RECT 69.790 134.640 73.240 134.780 ;
        RECT 69.790 134.500 69.930 134.640 ;
        RECT 72.920 134.580 73.240 134.640 ;
        RECT 76.155 134.595 76.445 134.825 ;
        RECT 78.915 134.780 79.205 134.825 ;
        RECT 81.200 134.780 81.520 134.840 ;
        RECT 86.260 134.780 86.580 134.840 ;
        RECT 78.915 134.640 81.520 134.780 ;
        RECT 78.915 134.595 79.205 134.640 ;
        RECT 69.700 134.240 70.020 134.500 ;
        RECT 70.175 134.440 70.465 134.485 ;
        RECT 75.680 134.440 76.000 134.500 ;
        RECT 70.175 134.300 76.000 134.440 ;
        RECT 76.230 134.440 76.370 134.595 ;
        RECT 81.200 134.580 81.520 134.640 ;
        RECT 81.750 134.640 86.580 134.780 ;
        RECT 81.750 134.485 81.890 134.640 ;
        RECT 86.260 134.580 86.580 134.640 ;
        RECT 89.035 134.780 89.325 134.825 ;
        RECT 89.940 134.780 90.260 134.840 ;
        RECT 89.035 134.640 90.260 134.780 ;
        RECT 89.035 134.595 89.325 134.640 ;
        RECT 89.940 134.580 90.260 134.640 ;
        RECT 98.695 134.595 98.985 134.825 ;
        RECT 103.740 134.780 104.060 134.840 ;
        RECT 106.975 134.780 107.265 134.825 ;
        RECT 122.600 134.780 122.920 134.840 ;
        RECT 103.740 134.640 107.265 134.780 ;
        RECT 76.230 134.300 81.430 134.440 ;
        RECT 70.175 134.255 70.465 134.300 ;
        RECT 75.680 134.240 76.000 134.300 ;
        RECT 81.290 134.160 81.430 134.300 ;
        RECT 81.675 134.255 81.965 134.485 ;
        RECT 82.135 134.440 82.425 134.485 ;
        RECT 82.580 134.440 82.900 134.500 ;
        RECT 82.135 134.300 82.900 134.440 ;
        RECT 82.135 134.255 82.425 134.300 ;
        RECT 82.580 134.240 82.900 134.300 ;
        RECT 83.500 134.440 83.820 134.500 ;
        RECT 87.640 134.440 87.960 134.500 ;
        RECT 83.500 134.300 87.960 134.440 ;
        RECT 83.500 134.240 83.820 134.300 ;
        RECT 87.640 134.240 87.960 134.300 ;
        RECT 95.920 134.440 96.240 134.500 ;
        RECT 98.770 134.440 98.910 134.595 ;
        RECT 103.740 134.580 104.060 134.640 ;
        RECT 106.975 134.595 107.265 134.640 ;
        RECT 110.500 134.640 122.920 134.780 ;
        RECT 110.500 134.440 110.640 134.640 ;
        RECT 122.600 134.580 122.920 134.640 ;
        RECT 123.060 134.440 123.380 134.500 ;
        RECT 95.920 134.300 110.640 134.440 ;
        RECT 112.110 134.300 123.380 134.440 ;
        RECT 95.920 134.240 96.240 134.300 ;
        RECT 68.795 134.100 69.085 134.145 ;
        RECT 67.860 133.960 69.085 134.100 ;
        RECT 67.860 133.900 68.180 133.960 ;
        RECT 68.795 133.915 69.085 133.960 ;
        RECT 69.255 134.100 69.545 134.145 ;
        RECT 71.540 134.100 71.860 134.160 ;
        RECT 69.255 133.960 71.860 134.100 ;
        RECT 69.255 133.915 69.545 133.960 ;
        RECT 71.540 133.900 71.860 133.960 ;
        RECT 72.000 134.100 72.320 134.160 ;
        RECT 72.475 134.100 72.765 134.145 ;
        RECT 72.000 133.960 72.765 134.100 ;
        RECT 72.000 133.900 72.320 133.960 ;
        RECT 72.475 133.915 72.765 133.960 ;
        RECT 67.950 133.760 68.090 133.900 ;
        RECT 64.270 133.620 68.090 133.760 ;
        RECT 72.550 133.760 72.690 133.915 ;
        RECT 73.380 133.900 73.700 134.160 ;
        RECT 76.615 134.100 76.905 134.145 ;
        RECT 78.900 134.100 79.220 134.160 ;
        RECT 76.615 133.960 79.220 134.100 ;
        RECT 76.615 133.915 76.905 133.960 ;
        RECT 78.900 133.900 79.220 133.960 ;
        RECT 81.200 133.900 81.520 134.160 ;
        RECT 83.040 133.900 83.360 134.160 ;
        RECT 84.435 134.120 84.725 134.145 ;
        RECT 84.050 133.980 84.725 134.120 ;
        RECT 73.840 133.760 74.160 133.820 ;
        RECT 72.550 133.620 74.160 133.760 ;
        RECT 61.420 133.560 61.740 133.620 ;
        RECT 73.840 133.560 74.160 133.620 ;
        RECT 75.220 133.760 75.540 133.820 ;
        RECT 77.995 133.760 78.285 133.805 ;
        RECT 80.280 133.760 80.600 133.820 ;
        RECT 75.220 133.620 75.910 133.760 ;
        RECT 75.220 133.560 75.540 133.620 ;
        RECT 64.640 133.420 64.960 133.480 ;
        RECT 61.050 133.280 64.960 133.420 ;
        RECT 64.640 133.220 64.960 133.280 ;
        RECT 67.860 133.420 68.180 133.480 ;
        RECT 68.335 133.420 68.625 133.465 ;
        RECT 67.860 133.280 68.625 133.420 ;
        RECT 67.860 133.220 68.180 133.280 ;
        RECT 68.335 133.235 68.625 133.280 ;
        RECT 70.175 133.420 70.465 133.465 ;
        RECT 72.000 133.420 72.320 133.480 ;
        RECT 70.175 133.280 72.320 133.420 ;
        RECT 70.175 133.235 70.465 133.280 ;
        RECT 72.000 133.220 72.320 133.280 ;
        RECT 72.920 133.420 73.240 133.480 ;
        RECT 75.770 133.465 75.910 133.620 ;
        RECT 77.995 133.620 80.600 133.760 ;
        RECT 84.050 133.760 84.190 133.980 ;
        RECT 84.435 133.915 84.725 133.980 ;
        RECT 84.895 134.100 85.185 134.145 ;
        RECT 85.800 134.100 86.120 134.160 ;
        RECT 84.895 133.960 86.120 134.100 ;
        RECT 84.895 133.915 85.185 133.960 ;
        RECT 85.800 133.900 86.120 133.960 ;
        RECT 86.260 133.900 86.580 134.160 ;
        RECT 95.460 133.900 95.780 134.160 ;
        RECT 105.135 134.100 105.425 134.145 ;
        RECT 106.960 134.100 107.280 134.160 ;
        RECT 112.110 134.145 112.250 134.300 ;
        RECT 123.060 134.240 123.380 134.300 ;
        RECT 105.135 133.960 107.280 134.100 ;
        RECT 105.135 133.915 105.425 133.960 ;
        RECT 106.960 133.900 107.280 133.960 ;
        RECT 107.510 133.960 108.570 134.100 ;
        RECT 94.080 133.760 94.400 133.820 ;
        RECT 84.050 133.620 94.400 133.760 ;
        RECT 77.995 133.575 78.285 133.620 ;
        RECT 80.280 133.560 80.600 133.620 ;
        RECT 94.080 133.560 94.400 133.620 ;
        RECT 103.740 133.760 104.060 133.820 ;
        RECT 106.040 133.760 106.360 133.820 ;
        RECT 103.740 133.620 106.360 133.760 ;
        RECT 103.740 133.560 104.060 133.620 ;
        RECT 106.040 133.560 106.360 133.620 ;
        RECT 72.920 133.280 75.450 133.420 ;
        RECT 72.920 133.220 73.240 133.280 ;
        RECT 52.680 133.080 53.000 133.140 ;
        RECT 55.915 133.080 56.205 133.125 ;
        RECT 52.680 132.940 56.205 133.080 ;
        RECT 52.680 132.880 53.000 132.940 ;
        RECT 55.915 132.895 56.205 132.940 ;
        RECT 57.280 133.080 57.600 133.140 ;
        RECT 58.215 133.080 58.505 133.125 ;
        RECT 58.660 133.080 58.980 133.140 ;
        RECT 57.280 132.940 58.980 133.080 ;
        RECT 57.280 132.880 57.600 132.940 ;
        RECT 58.215 132.895 58.505 132.940 ;
        RECT 58.660 132.880 58.980 132.940 ;
        RECT 61.895 133.080 62.185 133.125 ;
        RECT 62.340 133.080 62.660 133.140 ;
        RECT 61.895 132.940 62.660 133.080 ;
        RECT 61.895 132.895 62.185 132.940 ;
        RECT 62.340 132.880 62.660 132.940 ;
        RECT 64.180 133.080 64.500 133.140 ;
        RECT 71.555 133.080 71.845 133.125 ;
        RECT 74.300 133.080 74.620 133.140 ;
        RECT 64.180 132.940 74.620 133.080 ;
        RECT 75.310 133.080 75.450 133.280 ;
        RECT 75.695 133.235 75.985 133.465 ;
        RECT 77.075 133.420 77.365 133.465 ;
        RECT 77.520 133.420 77.840 133.480 ;
        RECT 83.500 133.420 83.820 133.480 ;
        RECT 77.075 133.280 77.840 133.420 ;
        RECT 77.075 133.235 77.365 133.280 ;
        RECT 77.520 133.220 77.840 133.280 ;
        RECT 79.450 133.280 83.820 133.420 ;
        RECT 79.450 133.080 79.590 133.280 ;
        RECT 83.500 133.220 83.820 133.280 ;
        RECT 85.815 133.420 86.105 133.465 ;
        RECT 107.510 133.420 107.650 133.960 ;
        RECT 107.895 133.575 108.185 133.805 ;
        RECT 85.815 133.280 107.650 133.420 ;
        RECT 85.815 133.235 86.105 133.280 ;
        RECT 75.310 132.940 79.590 133.080 ;
        RECT 79.820 133.080 80.140 133.140 ;
        RECT 80.295 133.080 80.585 133.125 ;
        RECT 79.820 132.940 80.585 133.080 ;
        RECT 64.180 132.880 64.500 132.940 ;
        RECT 71.555 132.895 71.845 132.940 ;
        RECT 74.300 132.880 74.620 132.940 ;
        RECT 79.820 132.880 80.140 132.940 ;
        RECT 80.295 132.895 80.585 132.940 ;
        RECT 86.260 133.080 86.580 133.140 ;
        RECT 92.700 133.080 93.020 133.140 ;
        RECT 86.260 132.940 93.020 133.080 ;
        RECT 86.260 132.880 86.580 132.940 ;
        RECT 92.700 132.880 93.020 132.940 ;
        RECT 93.620 133.080 93.940 133.140 ;
        RECT 96.840 133.080 97.160 133.140 ;
        RECT 93.620 132.940 97.160 133.080 ;
        RECT 93.620 132.880 93.940 132.940 ;
        RECT 96.840 132.880 97.160 132.940 ;
        RECT 97.760 133.080 98.080 133.140 ;
        RECT 107.970 133.080 108.110 133.575 ;
        RECT 108.430 133.420 108.570 133.960 ;
        RECT 112.035 133.915 112.325 134.145 ;
        RECT 112.480 133.900 112.800 134.160 ;
        RECT 113.400 133.900 113.720 134.160 ;
        RECT 123.520 133.900 123.840 134.160 ;
        RECT 110.640 133.760 110.960 133.820 ;
        RECT 111.115 133.760 111.405 133.805 ;
        RECT 110.640 133.620 111.405 133.760 ;
        RECT 110.640 133.560 110.960 133.620 ;
        RECT 111.115 133.575 111.405 133.620 ;
        RECT 111.575 133.760 111.865 133.805 ;
        RECT 111.575 133.620 111.975 133.760 ;
        RECT 111.575 133.575 111.865 133.620 ;
        RECT 111.650 133.420 111.790 133.575 ;
        RECT 115.700 133.420 116.020 133.480 ;
        RECT 108.430 133.280 116.020 133.420 ;
        RECT 115.700 133.220 116.020 133.280 ;
        RECT 117.095 133.420 117.385 133.465 ;
        RECT 117.540 133.420 117.860 133.480 ;
        RECT 117.095 133.280 117.860 133.420 ;
        RECT 117.095 133.235 117.385 133.280 ;
        RECT 117.540 133.220 117.860 133.280 ;
        RECT 118.000 133.420 118.320 133.480 ;
        RECT 120.300 133.420 120.620 133.480 ;
        RECT 118.000 133.280 120.620 133.420 ;
        RECT 118.000 133.220 118.320 133.280 ;
        RECT 120.300 133.220 120.620 133.280 ;
        RECT 97.760 132.940 108.110 133.080 ;
        RECT 108.815 133.080 109.105 133.125 ;
        RECT 109.260 133.080 109.580 133.140 ;
        RECT 108.815 132.940 109.580 133.080 ;
        RECT 97.760 132.880 98.080 132.940 ;
        RECT 108.815 132.895 109.105 132.940 ;
        RECT 109.260 132.880 109.580 132.940 ;
        RECT 110.180 132.880 110.500 133.140 ;
        RECT 53.990 132.260 125.290 132.740 ;
        RECT 59.135 132.060 59.425 132.105 ;
        RECT 59.580 132.060 59.900 132.120 ;
        RECT 59.135 131.920 59.900 132.060 ;
        RECT 59.135 131.875 59.425 131.920 ;
        RECT 59.580 131.860 59.900 131.920 ;
        RECT 65.100 132.060 65.420 132.120 ;
        RECT 77.520 132.060 77.840 132.120 ;
        RECT 65.100 131.920 77.840 132.060 ;
        RECT 65.100 131.860 65.420 131.920 ;
        RECT 77.520 131.860 77.840 131.920 ;
        RECT 78.440 131.860 78.760 132.120 ;
        RECT 79.360 132.060 79.680 132.120 ;
        RECT 86.260 132.060 86.580 132.120 ;
        RECT 79.360 131.920 86.580 132.060 ;
        RECT 79.360 131.860 79.680 131.920 ;
        RECT 86.260 131.860 86.580 131.920 ;
        RECT 88.560 131.860 88.880 132.120 ;
        RECT 89.940 132.060 90.260 132.120 ;
        RECT 91.320 132.060 91.640 132.120 ;
        RECT 89.940 131.920 91.640 132.060 ;
        RECT 89.940 131.860 90.260 131.920 ;
        RECT 91.320 131.860 91.640 131.920 ;
        RECT 92.255 132.060 92.545 132.105 ;
        RECT 92.700 132.060 93.020 132.120 ;
        RECT 92.255 131.920 93.020 132.060 ;
        RECT 92.255 131.875 92.545 131.920 ;
        RECT 92.700 131.860 93.020 131.920 ;
        RECT 93.620 132.060 93.940 132.120 ;
        RECT 96.395 132.060 96.685 132.105 ;
        RECT 107.420 132.060 107.740 132.120 ;
        RECT 93.620 131.920 96.685 132.060 ;
        RECT 93.620 131.860 93.940 131.920 ;
        RECT 96.395 131.875 96.685 131.920 ;
        RECT 97.850 131.920 107.740 132.060 ;
        RECT 55.440 131.720 55.760 131.780 ;
        RECT 61.435 131.720 61.725 131.765 ;
        RECT 55.440 131.580 61.725 131.720 ;
        RECT 55.440 131.520 55.760 131.580 ;
        RECT 61.435 131.535 61.725 131.580 ;
        RECT 61.880 131.720 62.200 131.780 ;
        RECT 64.655 131.720 64.945 131.765 ;
        RECT 73.380 131.720 73.700 131.780 ;
        RECT 73.855 131.720 74.145 131.765 ;
        RECT 61.880 131.580 73.150 131.720 ;
        RECT 61.880 131.520 62.200 131.580 ;
        RECT 64.655 131.535 64.945 131.580 ;
        RECT 60.960 131.380 61.280 131.440 ;
        RECT 57.370 131.240 61.280 131.380 ;
        RECT 56.820 130.840 57.140 131.100 ;
        RECT 57.370 131.085 57.510 131.240 ;
        RECT 60.960 131.180 61.280 131.240 ;
        RECT 67.400 131.380 67.720 131.440 ;
        RECT 69.240 131.380 69.560 131.440 ;
        RECT 67.400 131.240 69.560 131.380 ;
        RECT 67.400 131.180 67.720 131.240 ;
        RECT 69.240 131.180 69.560 131.240 ;
        RECT 70.620 131.380 70.940 131.440 ;
        RECT 71.555 131.380 71.845 131.425 ;
        RECT 72.000 131.380 72.320 131.440 ;
        RECT 70.620 131.240 72.320 131.380 ;
        RECT 73.010 131.380 73.150 131.580 ;
        RECT 73.380 131.580 74.145 131.720 ;
        RECT 73.380 131.520 73.700 131.580 ;
        RECT 73.855 131.535 74.145 131.580 ;
        RECT 74.760 131.520 75.080 131.780 ;
        RECT 75.220 131.720 75.540 131.780 ;
        RECT 75.695 131.720 75.985 131.765 ;
        RECT 75.220 131.580 75.985 131.720 ;
        RECT 75.220 131.520 75.540 131.580 ;
        RECT 75.695 131.535 75.985 131.580 ;
        RECT 80.740 131.720 81.060 131.780 ;
        RECT 83.040 131.720 83.360 131.780 ;
        RECT 86.720 131.720 87.040 131.780 ;
        RECT 80.740 131.580 83.360 131.720 ;
        RECT 80.740 131.520 81.060 131.580 ;
        RECT 83.040 131.520 83.360 131.580 ;
        RECT 84.050 131.580 87.040 131.720 ;
        RECT 73.010 131.240 74.070 131.380 ;
        RECT 70.620 131.180 70.940 131.240 ;
        RECT 71.555 131.195 71.845 131.240 ;
        RECT 72.000 131.180 72.320 131.240 ;
        RECT 57.295 130.855 57.585 131.085 ;
        RECT 58.200 131.040 58.520 131.100 ;
        RECT 58.675 131.040 58.965 131.085 ;
        RECT 59.120 131.040 59.440 131.100 ;
        RECT 58.200 130.900 59.440 131.040 ;
        RECT 58.200 130.840 58.520 130.900 ;
        RECT 58.675 130.855 58.965 130.900 ;
        RECT 59.120 130.840 59.440 130.900 ;
        RECT 60.055 131.040 60.345 131.085 ;
        RECT 64.640 131.040 64.960 131.100 ;
        RECT 60.055 130.900 64.960 131.040 ;
        RECT 60.055 130.855 60.345 130.900 ;
        RECT 64.640 130.840 64.960 130.900 ;
        RECT 65.575 130.855 65.865 131.085 ;
        RECT 56.910 130.700 57.050 130.840 ;
        RECT 61.895 130.700 62.185 130.745 ;
        RECT 56.910 130.560 57.970 130.700 ;
        RECT 56.375 130.360 56.665 130.405 ;
        RECT 56.820 130.360 57.140 130.420 ;
        RECT 57.830 130.405 57.970 130.560 ;
        RECT 61.050 130.560 62.185 130.700 ;
        RECT 56.375 130.220 57.140 130.360 ;
        RECT 56.375 130.175 56.665 130.220 ;
        RECT 56.820 130.160 57.140 130.220 ;
        RECT 57.755 130.175 58.045 130.405 ;
        RECT 60.500 130.360 60.820 130.420 ;
        RECT 61.050 130.360 61.190 130.560 ;
        RECT 61.895 130.515 62.185 130.560 ;
        RECT 62.340 130.700 62.660 130.760 ;
        RECT 62.815 130.700 63.105 130.745 ;
        RECT 62.340 130.560 63.105 130.700 ;
        RECT 65.650 130.700 65.790 130.855 ;
        RECT 72.920 130.840 73.240 131.100 ;
        RECT 66.020 130.700 66.340 130.760 ;
        RECT 65.650 130.560 66.340 130.700 ;
        RECT 73.930 130.700 74.070 131.240 ;
        RECT 74.315 131.040 74.605 131.085 ;
        RECT 74.850 131.040 74.990 131.520 ;
        RECT 74.315 130.900 74.990 131.040 ;
        RECT 74.315 130.855 74.605 130.900 ;
        RECT 75.680 130.840 76.000 131.100 ;
        RECT 79.360 131.040 79.680 131.100 ;
        RECT 84.050 131.040 84.190 131.580 ;
        RECT 86.720 131.520 87.040 131.580 ;
        RECT 87.180 131.520 87.500 131.780 ;
        RECT 87.270 131.380 87.410 131.520 ;
        RECT 88.650 131.425 88.790 131.860 ;
        RECT 85.430 131.240 87.410 131.380 ;
        RECT 79.360 130.900 84.190 131.040 ;
        RECT 79.360 130.840 79.680 130.900 ;
        RECT 84.880 130.840 85.200 131.100 ;
        RECT 85.430 131.085 85.570 131.240 ;
        RECT 88.575 131.195 88.865 131.425 ;
        RECT 85.355 130.855 85.645 131.085 ;
        RECT 86.275 130.855 86.565 131.085 ;
        RECT 82.580 130.700 82.900 130.760 ;
        RECT 73.930 130.560 82.900 130.700 ;
        RECT 62.340 130.500 62.660 130.560 ;
        RECT 62.815 130.515 63.105 130.560 ;
        RECT 66.020 130.500 66.340 130.560 ;
        RECT 82.580 130.500 82.900 130.560 ;
        RECT 86.350 130.420 86.490 130.855 ;
        RECT 86.720 130.840 87.040 131.100 ;
        RECT 87.280 131.040 87.570 131.085 ;
        RECT 87.280 130.900 87.870 131.040 ;
        RECT 87.280 130.855 87.570 130.900 ;
        RECT 87.730 130.700 87.870 130.900 ;
        RECT 89.020 130.840 89.340 131.100 ;
        RECT 90.030 131.085 90.170 131.860 ;
        RECT 96.840 131.720 97.160 131.780 ;
        RECT 90.950 131.580 97.160 131.720 ;
        RECT 90.950 131.085 91.090 131.580 ;
        RECT 96.840 131.520 97.160 131.580 ;
        RECT 97.850 131.380 97.990 131.920 ;
        RECT 107.420 131.860 107.740 131.920 ;
        RECT 119.380 132.060 119.700 132.120 ;
        RECT 120.300 132.060 120.620 132.120 ;
        RECT 119.380 131.920 120.620 132.060 ;
        RECT 119.380 131.860 119.700 131.920 ;
        RECT 120.300 131.860 120.620 131.920 ;
        RECT 121.220 132.060 121.540 132.120 ;
        RECT 122.615 132.060 122.905 132.105 ;
        RECT 121.220 131.920 122.905 132.060 ;
        RECT 121.220 131.860 121.540 131.920 ;
        RECT 122.615 131.875 122.905 131.920 ;
        RECT 114.780 131.720 115.100 131.780 ;
        RECT 114.780 131.580 123.750 131.720 ;
        RECT 114.780 131.520 115.100 131.580 ;
        RECT 92.790 131.240 97.990 131.380 ;
        RECT 98.235 131.420 98.525 131.425 ;
        RECT 98.235 131.380 99.370 131.420 ;
        RECT 104.200 131.380 104.520 131.440 ;
        RECT 113.400 131.380 113.720 131.440 ;
        RECT 117.080 131.380 117.400 131.440 ;
        RECT 98.235 131.280 117.400 131.380 ;
        RECT 89.825 130.900 90.170 131.085 ;
        RECT 89.825 130.855 90.115 130.900 ;
        RECT 90.875 130.855 91.165 131.085 ;
        RECT 91.335 131.040 91.625 131.085 ;
        RECT 92.240 131.040 92.560 131.100 ;
        RECT 91.335 130.900 92.560 131.040 ;
        RECT 91.335 130.855 91.625 130.900 ;
        RECT 92.240 130.840 92.560 130.900 ;
        RECT 88.560 130.700 88.880 130.760 ;
        RECT 87.730 130.560 88.880 130.700 ;
        RECT 88.560 130.500 88.880 130.560 ;
        RECT 90.400 130.500 90.720 130.760 ;
        RECT 60.500 130.220 61.190 130.360 ;
        RECT 63.735 130.360 64.025 130.405 ;
        RECT 64.180 130.360 64.500 130.420 ;
        RECT 63.735 130.220 64.500 130.360 ;
        RECT 60.500 130.160 60.820 130.220 ;
        RECT 63.735 130.175 64.025 130.220 ;
        RECT 64.180 130.160 64.500 130.220 ;
        RECT 65.100 130.360 65.420 130.420 ;
        RECT 68.335 130.360 68.625 130.405 ;
        RECT 65.100 130.220 68.625 130.360 ;
        RECT 65.100 130.160 65.420 130.220 ;
        RECT 68.335 130.175 68.625 130.220 ;
        RECT 70.160 130.160 70.480 130.420 ;
        RECT 70.635 130.360 70.925 130.405 ;
        RECT 71.080 130.360 71.400 130.420 ;
        RECT 70.635 130.220 71.400 130.360 ;
        RECT 70.635 130.175 70.925 130.220 ;
        RECT 71.080 130.160 71.400 130.220 ;
        RECT 71.540 130.360 71.860 130.420 ;
        RECT 74.775 130.360 75.065 130.405 ;
        RECT 71.540 130.220 75.065 130.360 ;
        RECT 71.540 130.160 71.860 130.220 ;
        RECT 74.775 130.175 75.065 130.220 ;
        RECT 86.260 130.160 86.580 130.420 ;
        RECT 87.180 130.360 87.500 130.420 ;
        RECT 92.790 130.360 92.930 131.240 ;
        RECT 98.235 131.195 98.525 131.280 ;
        RECT 99.230 131.240 117.400 131.280 ;
        RECT 104.200 131.180 104.520 131.240 ;
        RECT 113.400 131.180 113.720 131.240 ;
        RECT 117.080 131.180 117.400 131.240 ;
        RECT 118.920 131.380 119.240 131.440 ;
        RECT 122.155 131.380 122.445 131.425 ;
        RECT 118.920 131.240 122.445 131.380 ;
        RECT 118.920 131.180 119.240 131.240 ;
        RECT 122.155 131.195 122.445 131.240 ;
        RECT 95.000 130.840 95.320 131.100 ;
        RECT 96.855 131.040 97.145 131.085 ;
        RECT 97.300 131.040 97.620 131.100 ;
        RECT 96.855 130.900 97.620 131.040 ;
        RECT 96.855 130.855 97.145 130.900 ;
        RECT 87.180 130.220 92.930 130.360 ;
        RECT 96.930 130.360 97.070 130.855 ;
        RECT 97.300 130.840 97.620 130.900 ;
        RECT 97.760 130.840 98.080 131.100 ;
        RECT 98.875 130.910 99.165 131.055 ;
        RECT 98.875 130.825 99.370 130.910 ;
        RECT 99.600 130.840 99.920 131.100 ;
        RECT 100.060 130.840 100.380 131.100 ;
        RECT 107.420 131.040 107.740 131.100 ;
        RECT 108.815 131.040 109.105 131.085 ;
        RECT 118.460 131.040 118.780 131.100 ;
        RECT 120.315 131.040 120.605 131.085 ;
        RECT 107.420 130.900 114.090 131.040 ;
        RECT 107.420 130.840 107.740 130.900 ;
        RECT 108.815 130.855 109.105 130.900 ;
        RECT 98.950 130.770 99.370 130.825 ;
        RECT 99.230 130.700 99.370 130.770 ;
        RECT 113.400 130.700 113.720 130.760 ;
        RECT 99.230 130.560 113.720 130.700 ;
        RECT 113.400 130.500 113.720 130.560 ;
        RECT 105.580 130.360 105.900 130.420 ;
        RECT 96.930 130.220 105.900 130.360 ;
        RECT 87.180 130.160 87.500 130.220 ;
        RECT 105.580 130.160 105.900 130.220 ;
        RECT 106.960 130.360 107.280 130.420 ;
        RECT 110.655 130.360 110.945 130.405 ;
        RECT 106.960 130.220 110.945 130.360 ;
        RECT 113.950 130.360 114.090 130.900 ;
        RECT 118.460 130.900 120.605 131.040 ;
        RECT 118.460 130.840 118.780 130.900 ;
        RECT 120.315 130.855 120.605 130.900 ;
        RECT 123.060 130.840 123.380 131.100 ;
        RECT 123.610 131.085 123.750 131.580 ;
        RECT 123.535 130.855 123.825 131.085 ;
        RECT 118.000 130.500 118.320 130.760 ;
        RECT 118.935 130.700 119.225 130.745 ;
        RECT 118.935 130.560 120.070 130.700 ;
        RECT 118.935 130.515 119.225 130.560 ;
        RECT 119.395 130.360 119.685 130.405 ;
        RECT 113.950 130.220 119.685 130.360 ;
        RECT 119.930 130.360 120.070 130.560 ;
        RECT 121.220 130.500 121.540 130.760 ;
        RECT 122.600 130.360 122.920 130.420 ;
        RECT 119.930 130.220 122.920 130.360 ;
        RECT 106.960 130.160 107.280 130.220 ;
        RECT 110.655 130.175 110.945 130.220 ;
        RECT 119.395 130.175 119.685 130.220 ;
        RECT 122.600 130.160 122.920 130.220 ;
        RECT 53.990 129.540 125.290 130.020 ;
        RECT 52.680 129.340 53.000 129.400 ;
        RECT 55.915 129.340 56.205 129.385 ;
        RECT 60.040 129.340 60.360 129.400 ;
        RECT 52.680 129.200 56.205 129.340 ;
        RECT 52.680 129.140 53.000 129.200 ;
        RECT 55.915 129.155 56.205 129.200 ;
        RECT 57.370 129.200 60.360 129.340 ;
        RECT 56.820 128.460 57.140 128.720 ;
        RECT 57.370 128.705 57.510 129.200 ;
        RECT 60.040 129.140 60.360 129.200 ;
        RECT 61.880 129.340 62.200 129.400 ;
        RECT 63.735 129.340 64.025 129.385 ;
        RECT 73.840 129.340 74.160 129.400 ;
        RECT 79.360 129.340 79.680 129.400 ;
        RECT 61.880 129.200 64.025 129.340 ;
        RECT 61.880 129.140 62.200 129.200 ;
        RECT 63.735 129.155 64.025 129.200 ;
        RECT 66.570 129.200 73.610 129.340 ;
        RECT 57.755 129.000 58.045 129.045 ;
        RECT 59.580 129.000 59.900 129.060 ;
        RECT 61.435 129.000 61.725 129.045 ;
        RECT 66.570 129.000 66.710 129.200 ;
        RECT 57.755 128.860 59.350 129.000 ;
        RECT 57.755 128.815 58.045 128.860 ;
        RECT 59.210 128.705 59.350 128.860 ;
        RECT 59.580 128.860 61.190 129.000 ;
        RECT 59.580 128.800 59.900 128.860 ;
        RECT 57.295 128.475 57.585 128.705 ;
        RECT 58.215 128.660 58.505 128.705 ;
        RECT 58.215 128.520 58.890 128.660 ;
        RECT 58.215 128.475 58.505 128.520 ;
        RECT 58.750 127.980 58.890 128.520 ;
        RECT 59.135 128.475 59.425 128.705 ;
        RECT 60.040 128.460 60.360 128.720 ;
        RECT 60.500 128.460 60.820 128.720 ;
        RECT 61.050 128.660 61.190 128.860 ;
        RECT 61.435 128.860 66.710 129.000 ;
        RECT 71.095 129.000 71.385 129.045 ;
        RECT 73.470 129.000 73.610 129.200 ;
        RECT 73.840 129.200 79.680 129.340 ;
        RECT 73.840 129.140 74.160 129.200 ;
        RECT 79.360 129.140 79.680 129.200 ;
        RECT 79.820 129.340 80.140 129.400 ;
        RECT 80.755 129.340 81.045 129.385 ;
        RECT 79.820 129.200 81.045 129.340 ;
        RECT 79.820 129.140 80.140 129.200 ;
        RECT 80.755 129.155 81.045 129.200 ;
        RECT 82.120 129.140 82.440 129.400 ;
        RECT 84.880 129.140 85.200 129.400 ;
        RECT 87.180 129.140 87.500 129.400 ;
        RECT 100.980 129.340 101.300 129.400 ;
        RECT 90.950 129.200 101.300 129.340 ;
        RECT 87.270 129.000 87.410 129.140 ;
        RECT 71.095 128.860 72.690 129.000 ;
        RECT 73.470 128.860 84.690 129.000 ;
        RECT 61.435 128.815 61.725 128.860 ;
        RECT 71.095 128.815 71.385 128.860 ;
        RECT 63.440 128.660 63.730 128.705 ;
        RECT 61.050 128.520 63.730 128.660 ;
        RECT 63.440 128.475 63.730 128.520 ;
        RECT 64.180 128.660 64.500 128.720 ;
        RECT 65.575 128.660 65.865 128.705 ;
        RECT 64.180 128.520 65.865 128.660 ;
        RECT 64.180 128.460 64.500 128.520 ;
        RECT 65.575 128.475 65.865 128.520 ;
        RECT 66.020 128.460 66.340 128.720 ;
        RECT 66.480 128.460 66.800 128.720 ;
        RECT 67.415 128.475 67.705 128.705 ;
        RECT 67.875 128.660 68.165 128.705 ;
        RECT 69.240 128.660 69.560 128.720 ;
        RECT 67.875 128.520 69.560 128.660 ;
        RECT 67.875 128.475 68.165 128.520 ;
        RECT 59.595 128.320 59.885 128.365 ;
        RECT 60.960 128.320 61.280 128.380 ;
        RECT 59.595 128.180 61.280 128.320 ;
        RECT 59.595 128.135 59.885 128.180 ;
        RECT 60.960 128.120 61.280 128.180 ;
        RECT 62.340 128.320 62.660 128.380 ;
        RECT 67.490 128.320 67.630 128.475 ;
        RECT 62.340 128.180 67.630 128.320 ;
        RECT 62.340 128.120 62.660 128.180 ;
        RECT 61.420 127.980 61.740 128.040 ;
        RECT 58.750 127.840 61.740 127.980 ;
        RECT 61.420 127.780 61.740 127.840 ;
        RECT 66.495 127.980 66.785 128.025 ;
        RECT 67.950 127.980 68.090 128.475 ;
        RECT 69.240 128.460 69.560 128.520 ;
        RECT 70.620 128.660 70.940 128.720 ;
        RECT 72.550 128.660 72.690 128.860 ;
        RECT 73.380 128.660 73.700 128.720 ;
        RECT 75.235 128.660 75.525 128.705 ;
        RECT 70.620 128.650 71.770 128.660 ;
        RECT 70.620 128.520 72.230 128.650 ;
        RECT 72.550 128.520 75.525 128.660 ;
        RECT 70.620 128.460 70.940 128.520 ;
        RECT 71.630 128.510 72.230 128.520 ;
        RECT 68.320 128.320 68.640 128.380 ;
        RECT 72.090 128.365 72.230 128.510 ;
        RECT 73.380 128.460 73.700 128.520 ;
        RECT 75.235 128.475 75.525 128.520 ;
        RECT 75.695 128.660 75.985 128.705 ;
        RECT 77.980 128.660 78.300 128.720 ;
        RECT 81.200 128.660 81.520 128.720 ;
        RECT 75.695 128.520 77.750 128.660 ;
        RECT 75.695 128.475 75.985 128.520 ;
        RECT 68.320 128.180 69.930 128.320 ;
        RECT 68.320 128.120 68.640 128.180 ;
        RECT 66.495 127.840 68.090 127.980 ;
        RECT 69.790 127.980 69.930 128.180 ;
        RECT 71.555 128.135 71.845 128.365 ;
        RECT 72.015 128.135 72.305 128.365 ;
        RECT 75.770 128.320 75.910 128.475 ;
        RECT 72.550 128.180 75.910 128.320 ;
        RECT 71.630 127.980 71.770 128.135 ;
        RECT 72.550 127.980 72.690 128.180 ;
        RECT 76.155 128.135 76.445 128.365 ;
        RECT 69.790 127.840 71.310 127.980 ;
        RECT 71.630 127.840 72.690 127.980 ;
        RECT 75.220 127.980 75.540 128.040 ;
        RECT 76.230 127.980 76.370 128.135 ;
        RECT 75.220 127.840 76.370 127.980 ;
        RECT 77.610 127.980 77.750 128.520 ;
        RECT 77.980 128.520 81.520 128.660 ;
        RECT 77.980 128.460 78.300 128.520 ;
        RECT 81.200 128.460 81.520 128.520 ;
        RECT 79.360 128.320 79.680 128.380 ;
        RECT 81.675 128.320 81.965 128.365 ;
        RECT 79.360 128.180 81.965 128.320 ;
        RECT 79.360 128.120 79.680 128.180 ;
        RECT 81.675 128.135 81.965 128.180 ;
        RECT 82.580 128.320 82.900 128.380 ;
        RECT 83.055 128.320 83.345 128.365 ;
        RECT 82.580 128.180 83.345 128.320 ;
        RECT 84.550 128.320 84.690 128.860 ;
        RECT 86.350 128.860 87.410 129.000 ;
        RECT 88.560 129.000 88.880 129.060 ;
        RECT 90.950 129.045 91.090 129.200 ;
        RECT 100.980 129.140 101.300 129.200 ;
        RECT 107.420 129.140 107.740 129.400 ;
        RECT 112.940 129.340 113.260 129.400 ;
        RECT 121.220 129.340 121.540 129.400 ;
        RECT 112.940 129.200 121.540 129.340 ;
        RECT 112.940 129.140 113.260 129.200 ;
        RECT 121.220 129.140 121.540 129.200 ;
        RECT 88.560 128.860 89.710 129.000 ;
        RECT 84.895 128.660 85.185 128.705 ;
        RECT 85.340 128.660 85.660 128.720 ;
        RECT 84.895 128.520 85.660 128.660 ;
        RECT 84.895 128.475 85.185 128.520 ;
        RECT 85.340 128.460 85.660 128.520 ;
        RECT 85.800 128.460 86.120 128.720 ;
        RECT 86.350 128.705 86.490 128.860 ;
        RECT 88.560 128.800 88.880 128.860 ;
        RECT 86.275 128.475 86.565 128.705 ;
        RECT 87.015 128.475 87.305 128.705 ;
        RECT 89.035 128.475 89.325 128.705 ;
        RECT 87.090 128.320 87.230 128.475 ;
        RECT 84.550 128.180 87.230 128.320 ;
        RECT 82.580 128.120 82.900 128.180 ;
        RECT 83.055 128.135 83.345 128.180 ;
        RECT 87.655 128.135 87.945 128.365 ;
        RECT 79.820 127.980 80.140 128.040 ;
        RECT 77.610 127.840 80.140 127.980 ;
        RECT 66.495 127.795 66.785 127.840 ;
        RECT 62.815 127.640 63.105 127.685 ;
        RECT 63.720 127.640 64.040 127.700 ;
        RECT 62.815 127.500 64.040 127.640 ;
        RECT 62.815 127.455 63.105 127.500 ;
        RECT 63.720 127.440 64.040 127.500 ;
        RECT 67.860 127.640 68.180 127.700 ;
        RECT 68.335 127.640 68.625 127.685 ;
        RECT 67.860 127.500 68.625 127.640 ;
        RECT 67.860 127.440 68.180 127.500 ;
        RECT 68.335 127.455 68.625 127.500 ;
        RECT 69.255 127.640 69.545 127.685 ;
        RECT 69.700 127.640 70.020 127.700 ;
        RECT 69.255 127.500 70.020 127.640 ;
        RECT 71.170 127.640 71.310 127.840 ;
        RECT 75.220 127.780 75.540 127.840 ;
        RECT 79.820 127.780 80.140 127.840 ;
        RECT 84.475 127.980 84.765 128.025 ;
        RECT 85.800 127.980 86.120 128.040 ;
        RECT 87.730 127.980 87.870 128.135 ;
        RECT 88.100 128.120 88.420 128.380 ;
        RECT 88.560 128.320 88.880 128.380 ;
        RECT 89.110 128.320 89.250 128.475 ;
        RECT 88.560 128.180 89.250 128.320 ;
        RECT 89.570 128.320 89.710 128.860 ;
        RECT 90.875 128.815 91.165 129.045 ;
        RECT 91.320 129.000 91.640 129.060 ;
        RECT 95.000 129.000 95.320 129.060 ;
        RECT 91.320 128.860 95.320 129.000 ;
        RECT 91.320 128.800 91.640 128.860 ;
        RECT 95.000 128.800 95.320 128.860 ;
        RECT 95.475 129.000 95.765 129.045 ;
        RECT 95.920 129.000 96.240 129.060 ;
        RECT 95.475 128.860 96.240 129.000 ;
        RECT 95.475 128.815 95.765 128.860 ;
        RECT 95.920 128.800 96.240 128.860 ;
        RECT 105.135 129.000 105.425 129.045 ;
        RECT 111.100 129.000 111.420 129.060 ;
        RECT 105.135 128.860 111.420 129.000 ;
        RECT 105.135 128.815 105.425 128.860 ;
        RECT 111.100 128.800 111.420 128.860 ;
        RECT 122.140 129.000 122.460 129.060 ;
        RECT 123.075 129.000 123.365 129.045 ;
        RECT 122.140 128.860 123.365 129.000 ;
        RECT 122.140 128.800 122.460 128.860 ;
        RECT 123.075 128.815 123.365 128.860 ;
        RECT 89.955 128.660 90.245 128.705 ;
        RECT 90.415 128.660 90.705 128.705 ;
        RECT 89.955 128.520 90.705 128.660 ;
        RECT 89.955 128.475 90.245 128.520 ;
        RECT 90.415 128.475 90.705 128.520 ;
        RECT 92.255 128.660 92.545 128.705 ;
        RECT 93.160 128.660 93.480 128.720 ;
        RECT 107.125 128.660 107.415 128.705 ;
        RECT 92.255 128.520 93.480 128.660 ;
        RECT 92.255 128.475 92.545 128.520 ;
        RECT 93.160 128.460 93.480 128.520 ;
        RECT 101.530 128.520 107.415 128.660 ;
        RECT 101.530 128.380 101.670 128.520 ;
        RECT 107.125 128.475 107.415 128.520 ;
        RECT 109.735 128.660 110.025 128.705 ;
        RECT 110.180 128.660 110.500 128.720 ;
        RECT 109.735 128.520 110.500 128.660 ;
        RECT 109.735 128.475 110.025 128.520 ;
        RECT 110.180 128.460 110.500 128.520 ;
        RECT 111.575 128.475 111.865 128.705 ;
        RECT 112.020 128.660 112.340 128.720 ;
        RECT 113.860 128.660 114.180 128.720 ;
        RECT 112.020 128.520 114.180 128.660 ;
        RECT 91.335 128.320 91.625 128.365 ;
        RECT 92.700 128.320 93.020 128.380 ;
        RECT 89.570 128.180 93.020 128.320 ;
        RECT 88.560 128.120 88.880 128.180 ;
        RECT 91.335 128.135 91.625 128.180 ;
        RECT 92.700 128.120 93.020 128.180 ;
        RECT 94.080 128.320 94.400 128.380 ;
        RECT 95.920 128.320 96.240 128.380 ;
        RECT 94.080 128.180 96.240 128.320 ;
        RECT 94.080 128.120 94.400 128.180 ;
        RECT 95.920 128.120 96.240 128.180 ;
        RECT 101.440 128.120 101.760 128.380 ;
        RECT 109.260 128.320 109.580 128.380 ;
        RECT 111.650 128.320 111.790 128.475 ;
        RECT 112.020 128.460 112.340 128.520 ;
        RECT 113.860 128.460 114.180 128.520 ;
        RECT 121.220 128.660 121.540 128.720 ;
        RECT 121.695 128.660 121.985 128.705 ;
        RECT 121.220 128.520 121.985 128.660 ;
        RECT 121.220 128.460 121.540 128.520 ;
        RECT 121.695 128.475 121.985 128.520 ;
        RECT 122.155 128.320 122.445 128.365 ;
        RECT 109.260 128.180 122.445 128.320 ;
        RECT 109.260 128.120 109.580 128.180 ;
        RECT 122.155 128.135 122.445 128.180 ;
        RECT 84.475 127.840 87.870 127.980 ;
        RECT 89.480 127.980 89.800 128.040 ;
        RECT 106.515 127.980 106.805 128.025 ;
        RECT 89.480 127.840 106.805 127.980 ;
        RECT 84.475 127.795 84.765 127.840 ;
        RECT 85.800 127.780 86.120 127.840 ;
        RECT 89.480 127.780 89.800 127.840 ;
        RECT 106.515 127.795 106.805 127.840 ;
        RECT 73.395 127.640 73.685 127.685 ;
        RECT 71.170 127.500 73.685 127.640 ;
        RECT 69.255 127.455 69.545 127.500 ;
        RECT 69.700 127.440 70.020 127.500 ;
        RECT 73.395 127.455 73.685 127.500 ;
        RECT 77.520 127.640 77.840 127.700 ;
        RECT 78.915 127.640 79.205 127.685 ;
        RECT 77.520 127.500 79.205 127.640 ;
        RECT 77.520 127.440 77.840 127.500 ;
        RECT 78.915 127.455 79.205 127.500 ;
        RECT 81.200 127.640 81.520 127.700 ;
        RECT 83.515 127.640 83.805 127.685 ;
        RECT 81.200 127.500 83.805 127.640 ;
        RECT 81.200 127.440 81.520 127.500 ;
        RECT 83.515 127.455 83.805 127.500 ;
        RECT 89.020 127.640 89.340 127.700 ;
        RECT 97.300 127.640 97.620 127.700 ;
        RECT 89.020 127.500 97.620 127.640 ;
        RECT 89.020 127.440 89.340 127.500 ;
        RECT 97.300 127.440 97.620 127.500 ;
        RECT 98.680 127.440 99.000 127.700 ;
        RECT 100.520 127.640 100.840 127.700 ;
        RECT 109.275 127.640 109.565 127.685 ;
        RECT 100.520 127.500 109.565 127.640 ;
        RECT 100.520 127.440 100.840 127.500 ;
        RECT 109.275 127.455 109.565 127.500 ;
        RECT 110.640 127.440 110.960 127.700 ;
        RECT 115.255 127.640 115.545 127.685 ;
        RECT 120.300 127.640 120.620 127.700 ;
        RECT 115.255 127.500 120.620 127.640 ;
        RECT 115.255 127.455 115.545 127.500 ;
        RECT 120.300 127.440 120.620 127.500 ;
        RECT 53.990 126.820 125.290 127.300 ;
        RECT 56.375 126.620 56.665 126.665 ;
        RECT 57.740 126.620 58.060 126.680 ;
        RECT 65.100 126.620 65.420 126.680 ;
        RECT 56.375 126.480 58.060 126.620 ;
        RECT 56.375 126.435 56.665 126.480 ;
        RECT 57.740 126.420 58.060 126.480 ;
        RECT 59.670 126.480 65.420 126.620 ;
        RECT 59.670 126.325 59.810 126.480 ;
        RECT 65.100 126.420 65.420 126.480 ;
        RECT 67.415 126.620 67.705 126.665 ;
        RECT 67.860 126.620 68.180 126.680 ;
        RECT 67.415 126.480 68.180 126.620 ;
        RECT 67.415 126.435 67.705 126.480 ;
        RECT 67.860 126.420 68.180 126.480 ;
        RECT 68.795 126.620 69.085 126.665 ;
        RECT 69.240 126.620 69.560 126.680 ;
        RECT 68.795 126.480 69.560 126.620 ;
        RECT 68.795 126.435 69.085 126.480 ;
        RECT 69.240 126.420 69.560 126.480 ;
        RECT 71.080 126.620 71.400 126.680 ;
        RECT 73.380 126.620 73.700 126.680 ;
        RECT 71.080 126.480 73.700 126.620 ;
        RECT 71.080 126.420 71.400 126.480 ;
        RECT 73.380 126.420 73.700 126.480 ;
        RECT 73.840 126.420 74.160 126.680 ;
        RECT 74.775 126.620 75.065 126.665 ;
        RECT 76.140 126.620 76.460 126.680 ;
        RECT 74.775 126.480 76.460 126.620 ;
        RECT 74.775 126.435 75.065 126.480 ;
        RECT 76.140 126.420 76.460 126.480 ;
        RECT 79.360 126.420 79.680 126.680 ;
        RECT 85.355 126.620 85.645 126.665 ;
        RECT 86.260 126.620 86.580 126.680 ;
        RECT 81.750 126.480 85.110 126.620 ;
        RECT 59.595 126.095 59.885 126.325 ;
        RECT 60.040 126.080 60.360 126.340 ;
        RECT 62.355 126.280 62.645 126.325 ;
        RECT 63.260 126.280 63.580 126.340 ;
        RECT 62.355 126.140 63.580 126.280 ;
        RECT 62.355 126.095 62.645 126.140 ;
        RECT 63.260 126.080 63.580 126.140 ;
        RECT 63.720 126.280 64.040 126.340 ;
        RECT 66.940 126.280 67.260 126.340 ;
        RECT 63.720 126.140 66.710 126.280 ;
        RECT 63.720 126.080 64.040 126.140 ;
        RECT 57.755 125.940 58.045 125.985 ;
        RECT 57.755 125.800 59.350 125.940 ;
        RECT 57.755 125.755 58.045 125.800 ;
        RECT 55.440 125.400 55.760 125.660 ;
        RECT 57.295 125.415 57.585 125.645 ;
        RECT 58.215 125.600 58.505 125.645 ;
        RECT 58.660 125.600 58.980 125.660 ;
        RECT 59.210 125.645 59.350 125.800 ;
        RECT 61.420 125.740 61.740 126.000 ;
        RECT 64.180 125.940 64.500 126.000 ;
        RECT 65.575 125.940 65.865 125.985 ;
        RECT 64.180 125.800 65.865 125.940 ;
        RECT 66.570 125.940 66.710 126.140 ;
        RECT 66.940 126.140 75.910 126.280 ;
        RECT 66.940 126.080 67.260 126.140 ;
        RECT 72.015 125.940 72.305 125.985 ;
        RECT 75.220 125.940 75.540 126.000 ;
        RECT 66.570 125.800 71.770 125.940 ;
        RECT 64.180 125.740 64.500 125.800 ;
        RECT 65.575 125.755 65.865 125.800 ;
        RECT 58.215 125.460 58.980 125.600 ;
        RECT 58.215 125.415 58.505 125.460 ;
        RECT 57.370 125.260 57.510 125.415 ;
        RECT 58.660 125.400 58.980 125.460 ;
        RECT 59.135 125.415 59.425 125.645 ;
        RECT 60.500 125.400 60.820 125.660 ;
        RECT 61.510 125.600 61.650 125.740 ;
        RECT 62.980 125.600 63.270 125.645 ;
        RECT 61.510 125.460 63.270 125.600 ;
        RECT 62.980 125.415 63.270 125.460 ;
        RECT 65.115 125.600 65.405 125.645 ;
        RECT 67.860 125.600 68.180 125.660 ;
        RECT 65.115 125.460 68.180 125.600 ;
        RECT 65.115 125.415 65.405 125.460 ;
        RECT 67.860 125.400 68.180 125.460 ;
        RECT 68.335 125.600 68.625 125.645 ;
        RECT 70.160 125.600 70.480 125.660 ;
        RECT 68.335 125.460 70.480 125.600 ;
        RECT 71.630 125.600 71.770 125.800 ;
        RECT 72.015 125.800 75.540 125.940 ;
        RECT 72.015 125.755 72.305 125.800 ;
        RECT 75.220 125.740 75.540 125.800 ;
        RECT 75.770 125.725 75.910 126.140 ;
        RECT 80.280 126.080 80.600 126.340 ;
        RECT 72.935 125.600 73.225 125.645 ;
        RECT 73.840 125.600 74.160 125.660 ;
        RECT 71.630 125.460 72.760 125.600 ;
        RECT 68.335 125.415 68.625 125.460 ;
        RECT 70.160 125.400 70.480 125.460 ;
        RECT 60.040 125.260 60.360 125.320 ;
        RECT 57.370 125.120 60.360 125.260 ;
        RECT 60.040 125.060 60.360 125.120 ;
        RECT 61.435 125.260 61.725 125.305 ;
        RECT 70.635 125.260 70.925 125.305 ;
        RECT 71.540 125.260 71.860 125.320 ;
        RECT 61.435 125.120 66.250 125.260 ;
        RECT 61.435 125.075 61.725 125.120 ;
        RECT 61.880 124.920 62.200 124.980 ;
        RECT 63.275 124.920 63.565 124.965 ;
        RECT 61.880 124.780 63.565 124.920 ;
        RECT 61.880 124.720 62.200 124.780 ;
        RECT 63.275 124.735 63.565 124.780 ;
        RECT 64.180 124.920 64.500 124.980 ;
        RECT 65.560 124.920 65.880 124.980 ;
        RECT 64.180 124.780 65.880 124.920 ;
        RECT 66.110 124.920 66.250 125.120 ;
        RECT 70.635 125.120 71.860 125.260 ;
        RECT 72.620 125.260 72.760 125.460 ;
        RECT 72.935 125.460 74.160 125.600 ;
        RECT 75.695 125.495 75.985 125.725 ;
        RECT 72.935 125.415 73.225 125.460 ;
        RECT 73.840 125.400 74.160 125.460 ;
        RECT 77.060 125.400 77.380 125.660 ;
        RECT 77.520 125.400 77.840 125.660 ;
        RECT 78.455 125.600 78.745 125.645 ;
        RECT 78.900 125.600 79.220 125.660 ;
        RECT 78.455 125.460 79.220 125.600 ;
        RECT 78.455 125.415 78.745 125.460 ;
        RECT 78.900 125.400 79.220 125.460 ;
        RECT 81.215 125.600 81.505 125.645 ;
        RECT 81.750 125.600 81.890 126.480 ;
        RECT 82.120 126.280 82.440 126.340 ;
        RECT 84.970 126.280 85.110 126.480 ;
        RECT 85.355 126.480 86.580 126.620 ;
        RECT 85.355 126.435 85.645 126.480 ;
        RECT 86.260 126.420 86.580 126.480 ;
        RECT 89.955 126.620 90.245 126.665 ;
        RECT 90.860 126.620 91.180 126.680 ;
        RECT 89.955 126.480 91.180 126.620 ;
        RECT 89.955 126.435 90.245 126.480 ;
        RECT 90.860 126.420 91.180 126.480 ;
        RECT 91.795 126.620 92.085 126.665 ;
        RECT 92.700 126.620 93.020 126.680 ;
        RECT 101.440 126.620 101.760 126.680 ;
        RECT 91.795 126.480 101.760 126.620 ;
        RECT 91.795 126.435 92.085 126.480 ;
        RECT 92.700 126.420 93.020 126.480 ;
        RECT 101.440 126.420 101.760 126.480 ;
        RECT 103.280 126.620 103.600 126.680 ;
        RECT 108.800 126.620 109.120 126.680 ;
        RECT 103.280 126.480 105.810 126.620 ;
        RECT 103.280 126.420 103.600 126.480 ;
        RECT 85.800 126.280 86.120 126.340 ;
        RECT 88.560 126.280 88.880 126.340 ;
        RECT 95.460 126.280 95.780 126.340 ;
        RECT 105.670 126.280 105.810 126.480 ;
        RECT 108.800 126.480 116.390 126.620 ;
        RECT 108.800 126.420 109.120 126.480 ;
        RECT 111.100 126.280 111.420 126.340 ;
        RECT 115.700 126.280 116.020 126.340 ;
        RECT 82.120 126.140 84.190 126.280 ;
        RECT 84.970 126.140 86.120 126.280 ;
        RECT 82.120 126.080 82.440 126.140 ;
        RECT 83.500 125.645 83.820 125.670 ;
        RECT 84.050 125.645 84.190 126.140 ;
        RECT 85.800 126.080 86.120 126.140 ;
        RECT 87.255 126.140 88.880 126.280 ;
        RECT 87.255 125.940 87.395 126.140 ;
        RECT 88.560 126.080 88.880 126.140 ;
        RECT 90.030 126.140 95.230 126.280 ;
        RECT 85.430 125.800 87.395 125.940 ;
        RECT 81.215 125.460 81.890 125.600 ;
        RECT 81.215 125.415 81.505 125.460 ;
        RECT 82.135 125.415 82.425 125.645 ;
        RECT 82.595 125.415 82.885 125.645 ;
        RECT 83.235 125.415 83.820 125.645 ;
        RECT 83.975 125.415 84.265 125.645 ;
        RECT 82.210 125.260 82.350 125.415 ;
        RECT 72.620 125.120 82.350 125.260 ;
        RECT 82.670 125.260 82.810 125.415 ;
        RECT 83.500 125.410 83.820 125.415 ;
        RECT 85.430 125.260 85.570 125.800 ;
        RECT 86.260 125.400 86.580 125.660 ;
        RECT 86.735 125.415 87.025 125.645 ;
        RECT 87.255 125.600 87.395 125.800 ;
        RECT 87.640 125.740 87.960 126.000 ;
        RECT 88.115 125.600 88.405 125.645 ;
        RECT 87.255 125.460 88.405 125.600 ;
        RECT 88.115 125.415 88.405 125.460 ;
        RECT 82.670 125.120 85.570 125.260 ;
        RECT 85.800 125.260 86.120 125.320 ;
        RECT 86.810 125.260 86.950 125.415 ;
        RECT 88.560 125.400 88.880 125.660 ;
        RECT 89.020 125.400 89.340 125.660 ;
        RECT 90.030 125.645 90.170 126.140 ;
        RECT 90.400 125.940 90.720 126.000 ;
        RECT 95.090 125.940 95.230 126.140 ;
        RECT 95.460 126.140 105.350 126.280 ;
        RECT 105.670 126.140 116.020 126.280 ;
        RECT 95.460 126.080 95.780 126.140 ;
        RECT 101.900 125.940 102.220 126.000 ;
        RECT 90.400 125.800 91.090 125.940 ;
        RECT 95.090 125.800 102.220 125.940 ;
        RECT 90.400 125.740 90.720 125.800 ;
        RECT 90.950 125.645 91.090 125.800 ;
        RECT 101.900 125.740 102.220 125.800 ;
        RECT 89.955 125.415 90.245 125.645 ;
        RECT 90.875 125.415 91.165 125.645 ;
        RECT 92.255 125.600 92.545 125.645 ;
        RECT 96.840 125.600 97.160 125.660 ;
        RECT 92.255 125.460 97.160 125.600 ;
        RECT 92.255 125.415 92.545 125.460 ;
        RECT 96.840 125.400 97.160 125.460 ;
        RECT 103.740 125.600 104.060 125.660 ;
        RECT 105.210 125.645 105.350 126.140 ;
        RECT 111.100 126.080 111.420 126.140 ;
        RECT 115.700 126.080 116.020 126.140 ;
        RECT 113.400 125.940 113.720 126.000 ;
        RECT 116.250 125.940 116.390 126.480 ;
        RECT 121.220 126.420 121.540 126.680 ;
        RECT 113.400 125.800 115.470 125.940 ;
        RECT 116.250 125.800 122.370 125.940 ;
        RECT 113.400 125.740 113.720 125.800 ;
        RECT 104.215 125.600 104.505 125.645 ;
        RECT 103.740 125.460 104.505 125.600 ;
        RECT 103.740 125.400 104.060 125.460 ;
        RECT 104.215 125.415 104.505 125.460 ;
        RECT 105.135 125.415 105.425 125.645 ;
        RECT 110.640 125.600 110.960 125.660 ;
        RECT 115.330 125.645 115.470 125.800 ;
        RECT 110.500 125.400 110.960 125.600 ;
        RECT 114.335 125.415 114.625 125.645 ;
        RECT 115.255 125.415 115.545 125.645 ;
        RECT 101.915 125.260 102.205 125.305 ;
        RECT 110.500 125.260 110.640 125.400 ;
        RECT 85.800 125.120 101.670 125.260 ;
        RECT 70.635 125.075 70.925 125.120 ;
        RECT 71.540 125.060 71.860 125.120 ;
        RECT 68.320 124.920 68.640 124.980 ;
        RECT 66.110 124.780 68.640 124.920 ;
        RECT 64.180 124.720 64.500 124.780 ;
        RECT 65.560 124.720 65.880 124.780 ;
        RECT 68.320 124.720 68.640 124.780 ;
        RECT 71.095 124.920 71.385 124.965 ;
        RECT 72.460 124.920 72.780 124.980 ;
        RECT 71.095 124.780 72.780 124.920 ;
        RECT 71.095 124.735 71.385 124.780 ;
        RECT 72.460 124.720 72.780 124.780 ;
        RECT 72.920 124.920 73.240 124.980 ;
        RECT 75.680 124.920 76.000 124.980 ;
        RECT 72.920 124.780 76.000 124.920 ;
        RECT 72.920 124.720 73.240 124.780 ;
        RECT 75.680 124.720 76.000 124.780 ;
        RECT 79.820 124.920 80.140 124.980 ;
        RECT 82.670 124.920 82.810 125.120 ;
        RECT 85.800 125.060 86.120 125.120 ;
        RECT 79.820 124.780 82.810 124.920 ;
        RECT 89.480 124.920 89.800 124.980 ;
        RECT 91.780 124.920 92.100 124.980 ;
        RECT 89.480 124.780 92.100 124.920 ;
        RECT 79.820 124.720 80.140 124.780 ;
        RECT 89.480 124.720 89.800 124.780 ;
        RECT 91.780 124.720 92.100 124.780 ;
        RECT 95.000 124.920 95.320 124.980 ;
        RECT 100.060 124.920 100.380 124.980 ;
        RECT 95.000 124.780 100.380 124.920 ;
        RECT 101.530 124.920 101.670 125.120 ;
        RECT 101.915 125.120 110.640 125.260 ;
        RECT 114.410 125.260 114.550 125.415 ;
        RECT 115.700 125.400 116.020 125.660 ;
        RECT 116.160 125.400 116.480 125.660 ;
        RECT 118.920 125.600 119.240 125.660 ;
        RECT 122.230 125.645 122.370 125.800 ;
        RECT 119.395 125.600 119.685 125.645 ;
        RECT 118.920 125.460 119.685 125.600 ;
        RECT 118.920 125.400 119.240 125.460 ;
        RECT 119.395 125.415 119.685 125.460 ;
        RECT 121.695 125.415 121.985 125.645 ;
        RECT 122.155 125.415 122.445 125.645 ;
        RECT 117.555 125.260 117.845 125.305 ;
        RECT 121.220 125.260 121.540 125.320 ;
        RECT 114.410 125.120 116.390 125.260 ;
        RECT 101.915 125.075 102.205 125.120 ;
        RECT 116.250 124.980 116.390 125.120 ;
        RECT 117.555 125.120 121.540 125.260 ;
        RECT 121.770 125.260 121.910 125.415 ;
        RECT 123.060 125.400 123.380 125.660 ;
        RECT 124.440 125.260 124.760 125.320 ;
        RECT 125.360 125.260 125.680 125.320 ;
        RECT 121.770 125.120 125.680 125.260 ;
        RECT 117.555 125.075 117.845 125.120 ;
        RECT 121.220 125.060 121.540 125.120 ;
        RECT 124.440 125.060 124.760 125.120 ;
        RECT 125.360 125.060 125.680 125.120 ;
        RECT 106.500 124.920 106.820 124.980 ;
        RECT 101.530 124.780 106.820 124.920 ;
        RECT 95.000 124.720 95.320 124.780 ;
        RECT 100.060 124.720 100.380 124.780 ;
        RECT 106.500 124.720 106.820 124.780 ;
        RECT 112.020 124.920 112.340 124.980 ;
        RECT 112.495 124.920 112.785 124.965 ;
        RECT 112.020 124.780 112.785 124.920 ;
        RECT 112.020 124.720 112.340 124.780 ;
        RECT 112.495 124.735 112.785 124.780 ;
        RECT 116.160 124.720 116.480 124.980 ;
        RECT 117.080 124.920 117.400 124.980 ;
        RECT 119.840 124.920 120.160 124.980 ;
        RECT 122.615 124.920 122.905 124.965 ;
        RECT 117.080 124.780 122.905 124.920 ;
        RECT 117.080 124.720 117.400 124.780 ;
        RECT 119.840 124.720 120.160 124.780 ;
        RECT 122.615 124.735 122.905 124.780 ;
        RECT 53.990 124.100 125.290 124.580 ;
        RECT 54.520 123.900 54.840 123.960 ;
        RECT 57.755 123.900 58.045 123.945 ;
        RECT 54.520 123.760 58.045 123.900 ;
        RECT 54.520 123.700 54.840 123.760 ;
        RECT 57.755 123.715 58.045 123.760 ;
        RECT 60.500 123.900 60.820 123.960 ;
        RECT 61.435 123.900 61.725 123.945 ;
        RECT 60.500 123.760 61.725 123.900 ;
        RECT 60.500 123.700 60.820 123.760 ;
        RECT 61.435 123.715 61.725 123.760 ;
        RECT 62.355 123.900 62.645 123.945 ;
        RECT 63.720 123.900 64.040 123.960 ;
        RECT 62.355 123.760 64.040 123.900 ;
        RECT 62.355 123.715 62.645 123.760 ;
        RECT 63.720 123.700 64.040 123.760 ;
        RECT 64.655 123.715 64.945 123.945 ;
        RECT 56.820 123.560 57.140 123.620 ;
        RECT 59.595 123.560 59.885 123.605 ;
        RECT 56.820 123.420 59.885 123.560 ;
        RECT 64.730 123.560 64.870 123.715 ;
        RECT 66.020 123.700 66.340 123.960 ;
        RECT 66.480 123.900 66.800 123.960 ;
        RECT 66.955 123.900 67.245 123.945 ;
        RECT 66.480 123.760 67.245 123.900 ;
        RECT 66.480 123.700 66.800 123.760 ;
        RECT 66.955 123.715 67.245 123.760 ;
        RECT 71.080 123.700 71.400 123.960 ;
        RECT 72.000 123.900 72.320 123.960 ;
        RECT 72.920 123.900 73.240 123.960 ;
        RECT 72.000 123.760 73.240 123.900 ;
        RECT 72.000 123.700 72.320 123.760 ;
        RECT 72.920 123.700 73.240 123.760 ;
        RECT 77.060 123.900 77.380 123.960 ;
        RECT 80.295 123.900 80.585 123.945 ;
        RECT 77.060 123.760 80.585 123.900 ;
        RECT 77.060 123.700 77.380 123.760 ;
        RECT 80.295 123.715 80.585 123.760 ;
        RECT 83.040 123.700 83.360 123.960 ;
        RECT 83.960 123.900 84.280 123.960 ;
        RECT 84.435 123.900 84.725 123.945 ;
        RECT 83.960 123.760 84.725 123.900 ;
        RECT 83.960 123.700 84.280 123.760 ;
        RECT 84.435 123.715 84.725 123.760 ;
        RECT 86.735 123.900 87.025 123.945 ;
        RECT 89.940 123.900 90.260 123.960 ;
        RECT 86.735 123.760 90.260 123.900 ;
        RECT 86.735 123.715 87.025 123.760 ;
        RECT 89.940 123.700 90.260 123.760 ;
        RECT 95.920 123.900 96.240 123.960 ;
        RECT 96.840 123.900 97.160 123.960 ;
        RECT 95.920 123.760 97.160 123.900 ;
        RECT 95.920 123.700 96.240 123.760 ;
        RECT 96.840 123.700 97.160 123.760 ;
        RECT 97.300 123.700 97.620 123.960 ;
        RECT 98.220 123.900 98.540 123.960 ;
        RECT 99.600 123.900 99.920 123.960 ;
        RECT 101.455 123.900 101.745 123.945 ;
        RECT 98.220 123.760 98.910 123.900 ;
        RECT 98.220 123.700 98.540 123.760 ;
        RECT 67.400 123.560 67.720 123.620 ;
        RECT 64.730 123.420 67.720 123.560 ;
        RECT 56.820 123.360 57.140 123.420 ;
        RECT 59.595 123.375 59.885 123.420 ;
        RECT 67.400 123.360 67.720 123.420 ;
        RECT 69.700 123.560 70.020 123.620 ;
        RECT 81.200 123.560 81.520 123.620 ;
        RECT 90.875 123.560 91.165 123.605 ;
        RECT 92.700 123.560 93.020 123.620 ;
        RECT 97.390 123.560 97.530 123.700 ;
        RECT 98.770 123.605 98.910 123.760 ;
        RECT 99.600 123.760 101.745 123.900 ;
        RECT 99.600 123.700 99.920 123.760 ;
        RECT 101.455 123.715 101.745 123.760 ;
        RECT 104.200 123.900 104.520 123.960 ;
        RECT 104.675 123.900 104.965 123.945 ;
        RECT 104.200 123.760 104.965 123.900 ;
        RECT 104.200 123.700 104.520 123.760 ;
        RECT 104.675 123.715 104.965 123.760 ;
        RECT 109.720 123.900 110.040 123.960 ;
        RECT 114.335 123.900 114.625 123.945 ;
        RECT 123.060 123.900 123.380 123.960 ;
        RECT 109.720 123.760 123.380 123.900 ;
        RECT 109.720 123.700 110.040 123.760 ;
        RECT 114.335 123.715 114.625 123.760 ;
        RECT 123.060 123.700 123.380 123.760 ;
        RECT 69.700 123.420 81.520 123.560 ;
        RECT 69.700 123.360 70.020 123.420 ;
        RECT 81.200 123.360 81.520 123.420 ;
        RECT 82.210 123.420 90.170 123.560 ;
        RECT 54.060 123.220 54.380 123.280 ;
        RECT 57.295 123.220 57.585 123.265 ;
        RECT 54.060 123.080 57.585 123.220 ;
        RECT 54.060 123.020 54.380 123.080 ;
        RECT 57.295 123.035 57.585 123.080 ;
        RECT 58.660 123.020 58.980 123.280 ;
        RECT 60.960 123.020 61.280 123.280 ;
        RECT 61.880 123.020 62.200 123.280 ;
        RECT 62.800 123.220 63.120 123.280 ;
        RECT 63.275 123.220 63.565 123.265 ;
        RECT 62.800 123.080 63.565 123.220 ;
        RECT 62.800 123.020 63.120 123.080 ;
        RECT 63.275 123.035 63.565 123.080 ;
        RECT 63.720 123.020 64.040 123.280 ;
        RECT 65.100 123.020 65.420 123.280 ;
        RECT 66.495 123.035 66.785 123.265 ;
        RECT 57.740 122.880 58.060 122.940 ;
        RECT 66.570 122.880 66.710 123.035 ;
        RECT 68.780 123.020 69.100 123.280 ;
        RECT 70.175 123.035 70.465 123.265 ;
        RECT 71.095 123.220 71.385 123.265 ;
        RECT 76.600 123.220 76.920 123.280 ;
        RECT 71.095 123.080 76.920 123.220 ;
        RECT 71.095 123.035 71.385 123.080 ;
        RECT 57.740 122.740 66.710 122.880 ;
        RECT 70.250 122.880 70.390 123.035 ;
        RECT 76.600 123.020 76.920 123.080 ;
        RECT 79.820 123.220 80.140 123.280 ;
        RECT 82.210 123.220 82.350 123.420 ;
        RECT 90.030 123.280 90.170 123.420 ;
        RECT 90.875 123.420 94.310 123.560 ;
        RECT 90.875 123.375 91.165 123.420 ;
        RECT 92.700 123.360 93.020 123.420 ;
        RECT 79.820 123.080 82.350 123.220 ;
        RECT 79.820 123.020 80.140 123.080 ;
        RECT 82.580 123.020 82.900 123.280 ;
        RECT 83.975 123.220 84.265 123.265 ;
        RECT 84.420 123.220 84.740 123.280 ;
        RECT 83.975 123.080 84.740 123.220 ;
        RECT 83.975 123.035 84.265 123.080 ;
        RECT 84.420 123.020 84.740 123.080 ;
        RECT 85.340 123.020 85.660 123.280 ;
        RECT 85.815 123.035 86.105 123.265 ;
        RECT 88.115 123.220 88.405 123.265 ;
        RECT 89.020 123.220 89.340 123.280 ;
        RECT 88.115 123.080 89.340 123.220 ;
        RECT 88.115 123.035 88.405 123.080 ;
        RECT 72.000 122.880 72.320 122.940 ;
        RECT 80.755 122.880 81.045 122.925 ;
        RECT 70.250 122.740 81.045 122.880 ;
        RECT 57.740 122.680 58.060 122.740 ;
        RECT 72.000 122.680 72.320 122.740 ;
        RECT 80.755 122.695 81.045 122.740 ;
        RECT 81.215 122.695 81.505 122.925 ;
        RECT 85.890 122.880 86.030 123.035 ;
        RECT 89.020 123.020 89.340 123.080 ;
        RECT 89.480 123.020 89.800 123.280 ;
        RECT 89.940 123.020 90.260 123.280 ;
        RECT 90.400 123.220 90.720 123.280 ;
        RECT 91.335 123.220 91.625 123.265 ;
        RECT 90.400 123.080 91.625 123.220 ;
        RECT 90.400 123.020 90.720 123.080 ;
        RECT 91.335 123.035 91.625 123.080 ;
        RECT 91.780 123.020 92.100 123.280 ;
        RECT 94.170 123.265 94.310 123.420 ;
        RECT 94.630 123.420 97.530 123.560 ;
        RECT 94.095 123.035 94.385 123.265 ;
        RECT 88.560 122.880 88.880 122.940 ;
        RECT 93.175 122.880 93.465 122.925 ;
        RECT 85.890 122.740 88.330 122.880 ;
        RECT 54.980 122.540 55.300 122.600 ;
        RECT 67.875 122.540 68.165 122.585 ;
        RECT 54.980 122.400 68.165 122.540 ;
        RECT 54.980 122.340 55.300 122.400 ;
        RECT 67.875 122.355 68.165 122.400 ;
        RECT 68.320 122.540 68.640 122.600 ;
        RECT 79.820 122.540 80.140 122.600 ;
        RECT 81.290 122.540 81.430 122.695 ;
        RECT 68.320 122.400 80.140 122.540 ;
        RECT 68.320 122.340 68.640 122.400 ;
        RECT 79.820 122.340 80.140 122.400 ;
        RECT 80.370 122.400 81.430 122.540 ;
        RECT 81.660 122.540 81.980 122.600 ;
        RECT 87.195 122.540 87.485 122.585 ;
        RECT 81.660 122.400 87.485 122.540 ;
        RECT 88.190 122.540 88.330 122.740 ;
        RECT 88.560 122.740 93.465 122.880 ;
        RECT 88.560 122.680 88.880 122.740 ;
        RECT 93.175 122.695 93.465 122.740 ;
        RECT 94.630 122.540 94.770 123.420 ;
        RECT 98.695 123.375 98.985 123.605 ;
        RECT 110.640 123.560 110.960 123.620 ;
        RECT 120.300 123.560 120.620 123.620 ;
        RECT 123.535 123.560 123.825 123.605 ;
        RECT 110.640 123.420 112.710 123.560 ;
        RECT 110.640 123.360 110.960 123.420 ;
        RECT 95.935 123.035 96.225 123.265 ;
        RECT 96.855 123.220 97.145 123.265 ;
        RECT 97.300 123.220 97.620 123.280 ;
        RECT 96.855 123.080 97.620 123.220 ;
        RECT 96.855 123.035 97.145 123.080 ;
        RECT 95.015 122.695 95.305 122.925 ;
        RECT 88.190 122.400 94.770 122.540 ;
        RECT 95.090 122.540 95.230 122.695 ;
        RECT 95.460 122.680 95.780 122.940 ;
        RECT 96.010 122.880 96.150 123.035 ;
        RECT 97.300 123.020 97.620 123.080 ;
        RECT 98.235 123.035 98.525 123.265 ;
        RECT 99.155 123.220 99.445 123.265 ;
        RECT 99.600 123.220 99.920 123.280 ;
        RECT 99.155 123.080 99.920 123.220 ;
        RECT 99.155 123.035 99.445 123.080 ;
        RECT 97.760 122.880 98.080 122.940 ;
        RECT 96.010 122.740 98.080 122.880 ;
        RECT 98.310 122.880 98.450 123.035 ;
        RECT 99.600 123.020 99.920 123.080 ;
        RECT 100.075 123.220 100.365 123.265 ;
        RECT 100.520 123.220 100.840 123.280 ;
        RECT 100.075 123.080 100.840 123.220 ;
        RECT 100.075 123.035 100.365 123.080 ;
        RECT 100.520 123.020 100.840 123.080 ;
        RECT 101.440 123.220 101.760 123.280 ;
        RECT 102.835 123.220 103.125 123.265 ;
        RECT 101.440 123.080 103.125 123.220 ;
        RECT 101.440 123.020 101.760 123.080 ;
        RECT 102.835 123.035 103.125 123.080 ;
        RECT 112.020 123.020 112.340 123.280 ;
        RECT 112.570 123.265 112.710 123.420 ;
        RECT 120.300 123.420 123.825 123.560 ;
        RECT 120.300 123.360 120.620 123.420 ;
        RECT 123.535 123.375 123.825 123.420 ;
        RECT 112.495 123.035 112.785 123.265 ;
        RECT 112.940 123.020 113.260 123.280 ;
        RECT 98.310 122.740 101.210 122.880 ;
        RECT 97.760 122.680 98.080 122.740 ;
        RECT 97.850 122.540 97.990 122.680 ;
        RECT 101.070 122.600 101.210 122.740 ;
        RECT 102.375 122.695 102.665 122.925 ;
        RECT 112.110 122.880 112.250 123.020 ;
        RECT 122.140 122.880 122.460 122.940 ;
        RECT 112.110 122.740 122.460 122.880 ;
        RECT 100.520 122.540 100.840 122.600 ;
        RECT 95.090 122.400 96.290 122.540 ;
        RECT 97.850 122.400 100.840 122.540 ;
        RECT 80.370 122.260 80.510 122.400 ;
        RECT 81.660 122.340 81.980 122.400 ;
        RECT 87.195 122.355 87.485 122.400 ;
        RECT 56.360 122.000 56.680 122.260 ;
        RECT 60.055 122.200 60.345 122.245 ;
        RECT 60.960 122.200 61.280 122.260 ;
        RECT 62.340 122.200 62.660 122.260 ;
        RECT 60.055 122.060 62.660 122.200 ;
        RECT 60.055 122.015 60.345 122.060 ;
        RECT 60.960 122.000 61.280 122.060 ;
        RECT 62.340 122.000 62.660 122.060 ;
        RECT 65.100 122.200 65.420 122.260 ;
        RECT 80.280 122.200 80.600 122.260 ;
        RECT 65.100 122.060 80.600 122.200 ;
        RECT 65.100 122.000 65.420 122.060 ;
        RECT 80.280 122.000 80.600 122.060 ;
        RECT 80.740 122.200 81.060 122.260 ;
        RECT 82.135 122.200 82.425 122.245 ;
        RECT 80.740 122.060 82.425 122.200 ;
        RECT 80.740 122.000 81.060 122.060 ;
        RECT 82.135 122.015 82.425 122.060 ;
        RECT 86.260 122.200 86.580 122.260 ;
        RECT 88.560 122.200 88.880 122.260 ;
        RECT 86.260 122.060 88.880 122.200 ;
        RECT 86.260 122.000 86.580 122.060 ;
        RECT 88.560 122.000 88.880 122.060 ;
        RECT 91.780 122.200 92.100 122.260 ;
        RECT 92.715 122.200 93.005 122.245 ;
        RECT 91.780 122.060 93.005 122.200 ;
        RECT 96.150 122.200 96.290 122.400 ;
        RECT 100.520 122.340 100.840 122.400 ;
        RECT 100.980 122.340 101.300 122.600 ;
        RECT 102.450 122.540 102.590 122.695 ;
        RECT 122.140 122.680 122.460 122.740 ;
        RECT 105.120 122.540 105.440 122.600 ;
        RECT 117.080 122.540 117.400 122.600 ;
        RECT 102.450 122.400 105.440 122.540 ;
        RECT 105.120 122.340 105.440 122.400 ;
        RECT 110.500 122.400 117.400 122.540 ;
        RECT 96.840 122.200 97.160 122.260 ;
        RECT 96.150 122.060 97.160 122.200 ;
        RECT 91.780 122.000 92.100 122.060 ;
        RECT 92.715 122.015 93.005 122.060 ;
        RECT 96.840 122.000 97.160 122.060 ;
        RECT 97.315 122.200 97.605 122.245 ;
        RECT 97.760 122.200 98.080 122.260 ;
        RECT 97.315 122.060 98.080 122.200 ;
        RECT 97.315 122.015 97.605 122.060 ;
        RECT 97.760 122.000 98.080 122.060 ;
        RECT 102.820 122.200 103.140 122.260 ;
        RECT 110.500 122.200 110.640 122.400 ;
        RECT 117.080 122.340 117.400 122.400 ;
        RECT 102.820 122.060 110.640 122.200 ;
        RECT 102.820 122.000 103.140 122.060 ;
        RECT 116.160 122.000 116.480 122.260 ;
        RECT 53.990 121.380 125.290 121.860 ;
        RECT 59.120 120.980 59.440 121.240 ;
        RECT 62.800 121.180 63.120 121.240 ;
        RECT 65.100 121.180 65.420 121.240 ;
        RECT 62.800 121.040 65.420 121.180 ;
        RECT 62.800 120.980 63.120 121.040 ;
        RECT 65.100 120.980 65.420 121.040 ;
        RECT 66.495 121.180 66.785 121.225 ;
        RECT 68.780 121.180 69.100 121.240 ;
        RECT 77.075 121.180 77.365 121.225 ;
        RECT 66.495 121.040 69.100 121.180 ;
        RECT 66.495 120.995 66.785 121.040 ;
        RECT 68.780 120.980 69.100 121.040 ;
        RECT 70.710 121.040 77.365 121.180 ;
        RECT 60.055 120.840 60.345 120.885 ;
        RECT 62.340 120.840 62.660 120.900 ;
        RECT 63.260 120.840 63.580 120.900 ;
        RECT 60.055 120.700 61.230 120.840 ;
        RECT 60.055 120.655 60.345 120.700 ;
        RECT 57.295 120.160 57.585 120.205 ;
        RECT 58.200 120.160 58.520 120.220 ;
        RECT 57.295 120.020 58.520 120.160 ;
        RECT 61.090 120.160 61.230 120.700 ;
        RECT 62.200 120.700 63.580 120.840 ;
        RECT 62.200 120.640 62.660 120.700 ;
        RECT 63.260 120.640 63.580 120.700 ;
        RECT 64.180 120.640 64.500 120.900 ;
        RECT 61.435 120.500 61.725 120.545 ;
        RECT 62.200 120.500 62.340 120.640 ;
        RECT 61.435 120.360 62.340 120.500 ;
        RECT 62.800 120.500 63.120 120.560 ;
        RECT 66.480 120.500 66.800 120.560 ;
        RECT 70.710 120.545 70.850 121.040 ;
        RECT 77.075 120.995 77.365 121.040 ;
        RECT 80.740 120.980 81.060 121.240 ;
        RECT 85.800 120.980 86.120 121.240 ;
        RECT 90.400 121.180 90.720 121.240 ;
        RECT 91.795 121.180 92.085 121.225 ;
        RECT 87.275 121.040 92.085 121.180 ;
        RECT 72.460 120.640 72.780 120.900 ;
        RECT 73.395 120.840 73.685 120.885 ;
        RECT 79.820 120.840 80.140 120.900 ;
        RECT 87.275 120.840 87.415 121.040 ;
        RECT 90.400 120.980 90.720 121.040 ;
        RECT 91.795 120.995 92.085 121.040 ;
        RECT 94.080 121.180 94.400 121.240 ;
        RECT 100.060 121.180 100.380 121.240 ;
        RECT 100.995 121.180 101.285 121.225 ;
        RECT 94.080 121.040 98.910 121.180 ;
        RECT 73.395 120.700 80.140 120.840 ;
        RECT 73.395 120.655 73.685 120.700 ;
        RECT 79.820 120.640 80.140 120.700 ;
        RECT 80.370 120.700 87.415 120.840 ;
        RECT 80.370 120.545 80.510 120.700 ;
        RECT 87.655 120.655 87.945 120.885 ;
        RECT 90.875 120.840 91.165 120.885 ;
        RECT 90.030 120.700 91.165 120.840 ;
        RECT 62.800 120.360 66.800 120.500 ;
        RECT 61.435 120.315 61.725 120.360 ;
        RECT 62.800 120.300 63.120 120.360 ;
        RECT 66.480 120.300 66.800 120.360 ;
        RECT 68.335 120.315 68.625 120.545 ;
        RECT 70.635 120.315 70.925 120.545 ;
        RECT 72.935 120.500 73.225 120.545 ;
        RECT 80.295 120.500 80.585 120.545 ;
        RECT 72.935 120.360 80.585 120.500 ;
        RECT 72.935 120.315 73.225 120.360 ;
        RECT 80.295 120.315 80.585 120.360 ;
        RECT 81.200 120.500 81.520 120.560 ;
        RECT 83.515 120.500 83.805 120.545 ;
        RECT 83.960 120.500 84.280 120.560 ;
        RECT 81.200 120.360 84.280 120.500 ;
        RECT 61.880 120.160 62.200 120.220 ;
        RECT 61.090 120.020 62.200 120.160 ;
        RECT 57.295 119.975 57.585 120.020 ;
        RECT 58.200 119.960 58.520 120.020 ;
        RECT 61.880 119.960 62.200 120.020 ;
        RECT 65.115 120.160 65.405 120.205 ;
        RECT 68.410 120.160 68.550 120.315 ;
        RECT 81.200 120.300 81.520 120.360 ;
        RECT 83.515 120.315 83.805 120.360 ;
        RECT 83.960 120.300 84.280 120.360 ;
        RECT 84.895 120.500 85.185 120.545 ;
        RECT 87.180 120.500 87.500 120.560 ;
        RECT 87.730 120.500 87.870 120.655 ;
        RECT 89.495 120.500 89.785 120.545 ;
        RECT 84.895 120.360 86.950 120.500 ;
        RECT 84.895 120.315 85.185 120.360 ;
        RECT 65.115 120.020 68.550 120.160 ;
        RECT 65.115 119.975 65.405 120.020 ;
        RECT 69.240 119.960 69.560 120.220 ;
        RECT 69.700 119.960 70.020 120.220 ;
        RECT 70.160 119.960 70.480 120.220 ;
        RECT 71.555 119.975 71.845 120.205 ;
        RECT 72.015 120.160 72.305 120.205 ;
        RECT 73.380 120.160 73.700 120.220 ;
        RECT 72.015 120.020 73.700 120.160 ;
        RECT 72.015 119.975 72.305 120.020 ;
        RECT 56.375 119.820 56.665 119.865 ;
        RECT 60.500 119.820 60.820 119.880 ;
        RECT 56.375 119.680 60.820 119.820 ;
        RECT 56.375 119.635 56.665 119.680 ;
        RECT 57.830 119.540 57.970 119.680 ;
        RECT 60.500 119.620 60.820 119.680 ;
        RECT 66.495 119.820 66.785 119.865 ;
        RECT 71.080 119.820 71.400 119.880 ;
        RECT 66.495 119.680 71.400 119.820 ;
        RECT 66.495 119.635 66.785 119.680 ;
        RECT 71.080 119.620 71.400 119.680 ;
        RECT 57.740 119.280 58.060 119.540 ;
        RECT 58.200 119.280 58.520 119.540 ;
        RECT 65.100 119.480 65.420 119.540 ;
        RECT 65.575 119.480 65.865 119.525 ;
        RECT 65.100 119.340 65.865 119.480 ;
        RECT 71.630 119.480 71.770 119.975 ;
        RECT 73.380 119.960 73.700 120.020 ;
        RECT 73.840 120.210 74.160 120.220 ;
        RECT 73.840 120.205 74.300 120.210 ;
        RECT 73.840 119.975 74.385 120.205 ;
        RECT 73.840 119.960 74.160 119.975 ;
        RECT 74.760 119.960 75.080 120.220 ;
        RECT 76.140 120.160 76.460 120.220 ;
        RECT 75.945 120.020 76.460 120.160 ;
        RECT 76.140 119.960 76.460 120.020 ;
        RECT 76.600 119.960 76.920 120.220 ;
        RECT 77.980 119.960 78.300 120.220 ;
        RECT 78.900 119.960 79.220 120.220 ;
        RECT 79.820 120.205 80.140 120.220 ;
        RECT 79.605 119.975 80.140 120.205 ;
        RECT 79.820 119.960 80.140 119.975 ;
        RECT 80.740 120.160 81.060 120.220 ;
        RECT 81.675 120.160 81.965 120.205 ;
        RECT 80.740 120.020 81.965 120.160 ;
        RECT 80.740 119.960 81.060 120.020 ;
        RECT 81.675 119.975 81.965 120.020 ;
        RECT 82.135 119.975 82.425 120.205 ;
        RECT 85.800 120.160 86.120 120.220 ;
        RECT 86.275 120.160 86.565 120.205 ;
        RECT 85.800 120.020 86.565 120.160 ;
        RECT 75.235 119.820 75.525 119.865 ;
        RECT 75.235 119.680 75.910 119.820 ;
        RECT 75.235 119.635 75.525 119.680 ;
        RECT 75.770 119.540 75.910 119.680 ;
        RECT 74.760 119.480 75.080 119.540 ;
        RECT 71.630 119.340 75.080 119.480 ;
        RECT 65.100 119.280 65.420 119.340 ;
        RECT 65.575 119.295 65.865 119.340 ;
        RECT 74.760 119.280 75.080 119.340 ;
        RECT 75.680 119.280 76.000 119.540 ;
        RECT 76.230 119.480 76.370 119.960 ;
        RECT 78.440 119.620 78.760 119.880 ;
        RECT 81.200 119.480 81.520 119.540 ;
        RECT 76.230 119.340 81.520 119.480 ;
        RECT 82.210 119.480 82.350 119.975 ;
        RECT 85.800 119.960 86.120 120.020 ;
        RECT 86.275 119.975 86.565 120.020 ;
        RECT 83.975 119.820 84.265 119.865 ;
        RECT 84.420 119.820 84.740 119.880 ;
        RECT 83.975 119.680 84.740 119.820 ;
        RECT 83.975 119.635 84.265 119.680 ;
        RECT 84.420 119.620 84.740 119.680 ;
        RECT 84.895 119.820 85.185 119.865 ;
        RECT 85.340 119.820 85.660 119.880 ;
        RECT 84.895 119.680 85.660 119.820 ;
        RECT 84.895 119.635 85.185 119.680 ;
        RECT 85.340 119.620 85.660 119.680 ;
        RECT 82.580 119.480 82.900 119.540 ;
        RECT 86.810 119.525 86.950 120.360 ;
        RECT 87.180 120.360 89.785 120.500 ;
        RECT 87.180 120.300 87.500 120.360 ;
        RECT 89.495 120.315 89.785 120.360 ;
        RECT 87.640 120.160 87.960 120.220 ;
        RECT 88.560 120.160 88.880 120.220 ;
        RECT 90.030 120.160 90.170 120.700 ;
        RECT 90.875 120.655 91.165 120.700 ;
        RECT 91.870 120.500 92.010 120.995 ;
        RECT 94.080 120.980 94.400 121.040 ;
        RECT 95.460 120.840 95.780 120.900 ;
        RECT 95.090 120.700 95.780 120.840 ;
        RECT 95.090 120.500 95.230 120.700 ;
        RECT 95.460 120.640 95.780 120.700 ;
        RECT 95.935 120.655 96.225 120.885 ;
        RECT 96.380 120.840 96.700 120.900 ;
        RECT 97.315 120.840 97.605 120.885 ;
        RECT 96.380 120.700 97.605 120.840 ;
        RECT 98.770 120.840 98.910 121.040 ;
        RECT 100.060 121.040 101.285 121.180 ;
        RECT 100.060 120.980 100.380 121.040 ;
        RECT 100.995 120.995 101.285 121.040 ;
        RECT 101.900 120.980 102.220 121.240 ;
        RECT 107.420 121.180 107.740 121.240 ;
        RECT 119.395 121.180 119.685 121.225 ;
        RECT 107.420 121.040 119.685 121.180 ;
        RECT 107.420 120.980 107.740 121.040 ;
        RECT 119.395 120.995 119.685 121.040 ;
        RECT 108.800 120.840 109.120 120.900 ;
        RECT 98.770 120.700 100.290 120.840 ;
        RECT 96.010 120.500 96.150 120.655 ;
        RECT 96.380 120.640 96.700 120.700 ;
        RECT 97.315 120.655 97.605 120.700 ;
        RECT 99.600 120.500 99.920 120.560 ;
        RECT 91.870 120.360 95.230 120.500 ;
        RECT 92.700 120.160 93.020 120.220 ;
        RECT 95.090 120.205 95.230 120.360 ;
        RECT 95.550 120.360 96.150 120.500 ;
        RECT 96.470 120.360 99.920 120.500 ;
        RECT 95.550 120.220 95.690 120.360 ;
        RECT 93.175 120.160 93.465 120.205 ;
        RECT 87.640 120.020 88.880 120.160 ;
        RECT 87.640 119.960 87.960 120.020 ;
        RECT 88.560 119.960 88.880 120.020 ;
        RECT 89.110 120.020 90.170 120.160 ;
        RECT 90.490 120.020 93.465 120.160 ;
        RECT 89.110 119.880 89.250 120.020 ;
        RECT 89.020 119.620 89.340 119.880 ;
        RECT 82.210 119.340 82.900 119.480 ;
        RECT 81.200 119.280 81.520 119.340 ;
        RECT 82.580 119.280 82.900 119.340 ;
        RECT 86.735 119.480 87.025 119.525 ;
        RECT 90.490 119.480 90.630 120.020 ;
        RECT 92.700 119.960 93.020 120.020 ;
        RECT 93.175 119.975 93.465 120.020 ;
        RECT 95.015 119.975 95.305 120.205 ;
        RECT 95.460 119.960 95.780 120.220 ;
        RECT 90.860 119.820 91.180 119.880 ;
        RECT 94.095 119.820 94.385 119.865 ;
        RECT 90.860 119.680 94.385 119.820 ;
        RECT 90.860 119.620 91.180 119.680 ;
        RECT 94.095 119.635 94.385 119.680 ;
        RECT 86.735 119.340 90.630 119.480 ;
        RECT 94.170 119.480 94.310 119.635 ;
        RECT 94.540 119.620 94.860 119.880 ;
        RECT 96.470 119.480 96.610 120.360 ;
        RECT 99.600 120.300 99.920 120.360 ;
        RECT 97.300 119.960 97.620 120.220 ;
        RECT 97.760 120.160 98.080 120.220 ;
        RECT 99.140 120.205 99.460 120.220 ;
        RECT 100.150 120.205 100.290 120.700 ;
        RECT 104.290 120.700 109.120 120.840 ;
        RECT 102.820 120.500 103.140 120.560 ;
        RECT 104.290 120.500 104.430 120.700 ;
        RECT 108.800 120.640 109.120 120.700 ;
        RECT 113.400 120.640 113.720 120.900 ;
        RECT 116.620 120.840 116.940 120.900 ;
        RECT 117.555 120.840 117.845 120.885 ;
        RECT 116.620 120.700 117.845 120.840 ;
        RECT 116.620 120.640 116.940 120.700 ;
        RECT 117.555 120.655 117.845 120.700 ;
        RECT 119.840 120.840 120.160 120.900 ;
        RECT 119.840 120.700 120.990 120.840 ;
        RECT 119.840 120.640 120.160 120.700 ;
        RECT 102.820 120.360 104.430 120.500 ;
        RECT 102.820 120.300 103.140 120.360 ;
        RECT 98.695 120.160 98.985 120.205 ;
        RECT 97.760 120.020 98.985 120.160 ;
        RECT 97.760 119.960 98.080 120.020 ;
        RECT 98.695 119.975 98.985 120.020 ;
        RECT 99.140 119.975 99.470 120.205 ;
        RECT 100.075 119.975 100.365 120.205 ;
        RECT 101.440 120.160 101.760 120.220 ;
        RECT 104.290 120.205 104.430 120.360 ;
        RECT 105.210 120.360 120.530 120.500 ;
        RECT 105.210 120.220 105.350 120.360 ;
        RECT 120.390 120.220 120.530 120.360 ;
        RECT 103.295 120.160 103.585 120.205 ;
        RECT 101.440 120.020 103.585 120.160 ;
        RECT 99.140 119.960 99.460 119.975 ;
        RECT 101.440 119.960 101.760 120.020 ;
        RECT 103.295 119.975 103.585 120.020 ;
        RECT 103.755 119.975 104.045 120.205 ;
        RECT 104.215 119.975 104.505 120.205 ;
        RECT 98.220 119.620 98.540 119.880 ;
        RECT 103.830 119.820 103.970 119.975 ;
        RECT 105.120 119.960 105.440 120.220 ;
        RECT 105.580 119.960 105.900 120.220 ;
        RECT 106.960 119.960 107.280 120.220 ;
        RECT 109.720 120.160 110.040 120.220 ;
        RECT 108.430 120.020 110.040 120.160 ;
        RECT 108.430 119.820 108.570 120.020 ;
        RECT 109.720 119.960 110.040 120.020 ;
        RECT 110.180 120.160 110.500 120.220 ;
        RECT 113.860 120.160 114.180 120.220 ;
        RECT 116.175 120.160 116.465 120.205 ;
        RECT 110.180 120.020 116.465 120.160 ;
        RECT 110.180 119.960 110.500 120.020 ;
        RECT 113.860 119.960 114.180 120.020 ;
        RECT 116.175 119.975 116.465 120.020 ;
        RECT 117.080 119.960 117.400 120.220 ;
        RECT 120.300 119.960 120.620 120.220 ;
        RECT 120.850 120.160 120.990 120.700 ;
        RECT 121.220 120.640 121.540 120.900 ;
        RECT 121.695 120.160 121.985 120.205 ;
        RECT 120.850 120.020 121.985 120.160 ;
        RECT 121.695 119.975 121.985 120.020 ;
        RECT 122.155 119.975 122.445 120.205 ;
        RECT 103.830 119.680 108.570 119.820 ;
        RECT 108.800 119.820 109.120 119.880 ;
        RECT 122.230 119.820 122.370 119.975 ;
        RECT 108.800 119.680 122.370 119.820 ;
        RECT 105.210 119.540 105.350 119.680 ;
        RECT 108.800 119.620 109.120 119.680 ;
        RECT 94.170 119.340 96.610 119.480 ;
        RECT 86.735 119.295 87.025 119.340 ;
        RECT 105.120 119.280 105.440 119.540 ;
        RECT 106.055 119.480 106.345 119.525 ;
        RECT 106.500 119.480 106.820 119.540 ;
        RECT 106.055 119.340 106.820 119.480 ;
        RECT 106.055 119.295 106.345 119.340 ;
        RECT 106.500 119.280 106.820 119.340 ;
        RECT 123.060 119.280 123.380 119.540 ;
        RECT 53.990 118.660 125.290 119.140 ;
        RECT 61.895 118.275 62.185 118.505 ;
        RECT 69.240 118.460 69.560 118.520 ;
        RECT 76.140 118.460 76.460 118.520 ;
        RECT 82.135 118.460 82.425 118.505 ;
        RECT 69.240 118.320 82.425 118.460 ;
        RECT 53.600 118.120 53.920 118.180 ;
        RECT 61.970 118.120 62.110 118.275 ;
        RECT 69.240 118.260 69.560 118.320 ;
        RECT 76.140 118.260 76.460 118.320 ;
        RECT 82.135 118.275 82.425 118.320 ;
        RECT 83.040 118.260 83.360 118.520 ;
        RECT 84.420 118.310 84.740 118.520 ;
        RECT 87.195 118.460 87.485 118.505 ;
        RECT 89.020 118.460 89.340 118.520 ;
        RECT 84.970 118.320 85.570 118.460 ;
        RECT 84.970 118.310 85.110 118.320 ;
        RECT 84.420 118.260 85.110 118.310 ;
        RECT 53.600 117.980 62.110 118.120 ;
        RECT 69.715 118.120 70.005 118.165 ;
        RECT 71.540 118.120 71.860 118.180 ;
        RECT 69.715 117.980 71.860 118.120 ;
        RECT 53.600 117.920 53.920 117.980 ;
        RECT 69.715 117.935 70.005 117.980 ;
        RECT 71.540 117.920 71.860 117.980 ;
        RECT 78.440 118.120 78.760 118.180 ;
        RECT 84.515 118.170 85.110 118.260 ;
        RECT 85.430 118.120 85.570 118.320 ;
        RECT 87.195 118.320 89.340 118.460 ;
        RECT 87.195 118.275 87.485 118.320 ;
        RECT 89.020 118.260 89.340 118.320 ;
        RECT 99.140 118.460 99.460 118.520 ;
        RECT 100.995 118.460 101.285 118.505 ;
        RECT 99.140 118.320 101.285 118.460 ;
        RECT 99.140 118.260 99.460 118.320 ;
        RECT 95.920 118.120 96.240 118.180 ;
        RECT 97.775 118.120 98.065 118.165 ;
        RECT 78.440 117.980 81.890 118.120 ;
        RECT 85.430 117.980 92.930 118.120 ;
        RECT 78.440 117.920 78.760 117.980 ;
        RECT 81.750 117.840 81.890 117.980 ;
        RECT 55.440 117.580 55.760 117.840 ;
        RECT 57.740 117.580 58.060 117.840 ;
        RECT 58.525 117.780 58.815 117.825 ;
        RECT 60.500 117.780 60.820 117.840 ;
        RECT 58.525 117.640 60.820 117.780 ;
        RECT 58.525 117.595 58.815 117.640 ;
        RECT 60.500 117.580 60.820 117.640 ;
        RECT 60.960 117.780 61.280 117.840 ;
        RECT 61.435 117.780 61.725 117.825 ;
        RECT 60.960 117.640 61.725 117.780 ;
        RECT 60.960 117.580 61.280 117.640 ;
        RECT 61.435 117.595 61.725 117.640 ;
        RECT 62.800 117.580 63.120 117.840 ;
        RECT 63.275 117.595 63.565 117.825 ;
        RECT 69.255 117.595 69.545 117.825 ;
        RECT 70.160 117.780 70.480 117.840 ;
        RECT 75.680 117.780 76.000 117.840 ;
        RECT 70.160 117.640 76.000 117.780 ;
        RECT 53.140 117.440 53.460 117.500 ;
        RECT 63.350 117.440 63.490 117.595 ;
        RECT 53.140 117.300 63.490 117.440 ;
        RECT 69.330 117.440 69.470 117.595 ;
        RECT 70.160 117.580 70.480 117.640 ;
        RECT 75.680 117.580 76.000 117.640 ;
        RECT 81.215 117.595 81.505 117.825 ;
        RECT 69.700 117.440 70.020 117.500 ;
        RECT 72.000 117.440 72.320 117.500 ;
        RECT 69.330 117.300 72.320 117.440 ;
        RECT 53.140 117.240 53.460 117.300 ;
        RECT 69.700 117.240 70.020 117.300 ;
        RECT 72.000 117.240 72.320 117.300 ;
        RECT 80.740 117.440 81.060 117.500 ;
        RECT 81.290 117.440 81.430 117.595 ;
        RECT 81.660 117.580 81.980 117.840 ;
        RECT 83.040 117.780 83.360 117.840 ;
        RECT 83.515 117.780 83.805 117.825 ;
        RECT 83.040 117.640 83.805 117.780 ;
        RECT 84.880 117.700 85.200 117.960 ;
        RECT 83.040 117.580 83.360 117.640 ;
        RECT 83.515 117.595 83.805 117.640 ;
        RECT 84.895 117.595 85.185 117.700 ;
        RECT 85.815 117.595 86.105 117.825 ;
        RECT 86.260 117.780 86.580 117.840 ;
        RECT 86.735 117.780 87.025 117.825 ;
        RECT 86.260 117.640 87.025 117.780 ;
        RECT 80.740 117.300 81.430 117.440 ;
        RECT 81.750 117.300 85.115 117.440 ;
        RECT 80.740 117.240 81.060 117.300 ;
        RECT 81.750 117.160 81.890 117.300 ;
        RECT 59.580 116.900 59.900 117.160 ;
        RECT 64.180 116.900 64.500 117.160 ;
        RECT 80.295 117.100 80.585 117.145 ;
        RECT 81.660 117.100 81.980 117.160 ;
        RECT 80.295 116.960 81.980 117.100 ;
        RECT 80.295 116.915 80.585 116.960 ;
        RECT 81.660 116.900 81.980 116.960 ;
        RECT 56.360 116.560 56.680 116.820 ;
        RECT 60.500 116.560 60.820 116.820 ;
        RECT 74.760 116.760 75.080 116.820 ;
        RECT 76.600 116.760 76.920 116.820 ;
        RECT 74.760 116.620 76.920 116.760 ;
        RECT 74.760 116.560 75.080 116.620 ;
        RECT 76.600 116.560 76.920 116.620 ;
        RECT 82.580 116.760 82.900 116.820 ;
        RECT 83.515 116.760 83.805 116.805 ;
        RECT 82.580 116.620 83.805 116.760 ;
        RECT 84.975 116.760 85.115 117.300 ;
        RECT 85.340 117.100 85.660 117.160 ;
        RECT 85.890 117.100 86.030 117.595 ;
        RECT 86.260 117.580 86.580 117.640 ;
        RECT 86.735 117.595 87.025 117.640 ;
        RECT 88.115 117.780 88.405 117.825 ;
        RECT 89.020 117.780 89.340 117.840 ;
        RECT 88.115 117.640 89.340 117.780 ;
        RECT 88.115 117.595 88.405 117.640 ;
        RECT 89.020 117.580 89.340 117.640 ;
        RECT 89.480 117.580 89.800 117.840 ;
        RECT 89.940 117.580 90.260 117.840 ;
        RECT 90.875 117.780 91.165 117.825 ;
        RECT 91.780 117.780 92.100 117.840 ;
        RECT 90.875 117.640 92.100 117.780 ;
        RECT 90.875 117.595 91.165 117.640 ;
        RECT 91.780 117.580 92.100 117.640 ;
        RECT 92.240 117.580 92.560 117.840 ;
        RECT 92.790 117.780 92.930 117.980 ;
        RECT 95.920 117.980 98.065 118.120 ;
        RECT 95.920 117.920 96.240 117.980 ;
        RECT 97.775 117.935 98.065 117.980 ;
        RECT 99.690 117.935 99.830 118.320 ;
        RECT 100.995 118.275 101.285 118.320 ;
        RECT 106.960 118.460 107.280 118.520 ;
        RECT 114.320 118.460 114.640 118.520 ;
        RECT 106.960 118.320 114.640 118.460 ;
        RECT 106.960 118.260 107.280 118.320 ;
        RECT 100.520 118.120 100.840 118.180 ;
        RECT 105.120 118.120 105.440 118.180 ;
        RECT 107.970 118.165 108.110 118.320 ;
        RECT 114.320 118.260 114.640 118.320 ;
        RECT 117.080 118.460 117.400 118.520 ;
        RECT 120.300 118.460 120.620 118.520 ;
        RECT 117.080 118.320 120.620 118.460 ;
        RECT 117.080 118.260 117.400 118.320 ;
        RECT 120.300 118.260 120.620 118.320 ;
        RECT 107.435 118.120 107.725 118.165 ;
        RECT 100.520 117.980 104.890 118.120 ;
        RECT 96.395 117.780 96.685 117.825 ;
        RECT 96.840 117.780 97.160 117.840 ;
        RECT 92.790 117.640 95.690 117.780 ;
        RECT 90.415 117.440 90.705 117.485 ;
        RECT 86.810 117.300 90.705 117.440 ;
        RECT 86.810 117.160 86.950 117.300 ;
        RECT 90.415 117.255 90.705 117.300 ;
        RECT 93.635 117.255 93.925 117.485 ;
        RECT 94.095 117.440 94.385 117.485 ;
        RECT 95.000 117.440 95.320 117.500 ;
        RECT 94.095 117.300 95.320 117.440 ;
        RECT 95.550 117.440 95.690 117.640 ;
        RECT 96.395 117.640 97.160 117.780 ;
        RECT 96.395 117.595 96.685 117.640 ;
        RECT 96.840 117.580 97.160 117.640 ;
        RECT 97.300 117.580 97.620 117.840 ;
        RECT 98.220 117.780 98.540 117.840 ;
        RECT 98.695 117.780 98.985 117.825 ;
        RECT 98.220 117.640 98.985 117.780 ;
        RECT 98.220 117.580 98.540 117.640 ;
        RECT 98.695 117.595 98.985 117.640 ;
        RECT 95.935 117.440 96.225 117.485 ;
        RECT 95.550 117.300 98.450 117.440 ;
        RECT 94.095 117.255 94.385 117.300 ;
        RECT 85.340 116.960 86.030 117.100 ;
        RECT 85.340 116.900 85.660 116.960 ;
        RECT 86.260 116.900 86.580 117.160 ;
        RECT 86.720 116.900 87.040 117.160 ;
        RECT 88.575 117.100 88.865 117.145 ;
        RECT 90.860 117.100 91.180 117.160 ;
        RECT 88.575 116.960 91.180 117.100 ;
        RECT 88.575 116.915 88.865 116.960 ;
        RECT 90.860 116.900 91.180 116.960 ;
        RECT 91.335 117.100 91.625 117.145 ;
        RECT 93.710 117.100 93.850 117.255 ;
        RECT 95.000 117.240 95.320 117.300 ;
        RECT 95.935 117.255 96.225 117.300 ;
        RECT 97.775 117.100 98.065 117.145 ;
        RECT 91.335 116.960 93.390 117.100 ;
        RECT 93.710 116.960 98.065 117.100 ;
        RECT 91.335 116.915 91.625 116.960 ;
        RECT 87.180 116.760 87.500 116.820 ;
        RECT 84.975 116.620 87.500 116.760 ;
        RECT 82.580 116.560 82.900 116.620 ;
        RECT 83.515 116.575 83.805 116.620 ;
        RECT 87.180 116.560 87.500 116.620 ;
        RECT 91.780 116.760 92.100 116.820 ;
        RECT 92.715 116.760 93.005 116.805 ;
        RECT 91.780 116.620 93.005 116.760 ;
        RECT 93.250 116.760 93.390 116.960 ;
        RECT 97.775 116.915 98.065 116.960 ;
        RECT 94.080 116.760 94.400 116.820 ;
        RECT 93.250 116.620 94.400 116.760 ;
        RECT 91.780 116.560 92.100 116.620 ;
        RECT 92.715 116.575 93.005 116.620 ;
        RECT 94.080 116.560 94.400 116.620 ;
        RECT 95.000 116.760 95.320 116.820 ;
        RECT 96.855 116.760 97.145 116.805 ;
        RECT 95.000 116.620 97.145 116.760 ;
        RECT 95.000 116.560 95.320 116.620 ;
        RECT 96.855 116.575 97.145 116.620 ;
        RECT 97.300 116.760 97.620 116.820 ;
        RECT 98.310 116.760 98.450 117.300 ;
        RECT 98.770 117.100 98.910 117.595 ;
        RECT 99.140 117.580 99.460 117.840 ;
        RECT 99.640 117.705 99.930 117.935 ;
        RECT 100.520 117.920 100.840 117.980 ;
        RECT 102.375 117.780 102.665 117.825 ;
        RECT 100.610 117.640 102.665 117.780 ;
        RECT 100.610 117.500 100.750 117.640 ;
        RECT 102.375 117.595 102.665 117.640 ;
        RECT 103.280 117.780 103.600 117.840 ;
        RECT 103.755 117.780 104.045 117.825 ;
        RECT 103.280 117.640 104.045 117.780 ;
        RECT 103.280 117.580 103.600 117.640 ;
        RECT 103.755 117.595 104.045 117.640 ;
        RECT 100.520 117.240 100.840 117.500 ;
        RECT 101.440 117.440 101.760 117.500 ;
        RECT 101.915 117.440 102.205 117.485 ;
        RECT 101.440 117.300 102.205 117.440 ;
        RECT 101.440 117.240 101.760 117.300 ;
        RECT 101.915 117.255 102.205 117.300 ;
        RECT 102.820 117.440 103.140 117.500 ;
        RECT 104.215 117.440 104.505 117.485 ;
        RECT 102.820 117.300 104.505 117.440 ;
        RECT 104.750 117.440 104.890 117.980 ;
        RECT 105.120 117.980 107.725 118.120 ;
        RECT 105.120 117.920 105.440 117.980 ;
        RECT 107.435 117.935 107.725 117.980 ;
        RECT 107.895 117.935 108.185 118.165 ;
        RECT 113.875 118.120 114.165 118.165 ;
        RECT 117.540 118.120 117.860 118.180 ;
        RECT 113.875 117.980 117.860 118.120 ;
        RECT 113.875 117.935 114.165 117.980 ;
        RECT 117.540 117.920 117.860 117.980 ;
        RECT 106.960 117.580 107.280 117.840 ;
        RECT 108.815 117.595 109.105 117.825 ;
        RECT 110.195 117.780 110.485 117.825 ;
        RECT 111.100 117.780 111.420 117.840 ;
        RECT 112.940 117.780 113.260 117.840 ;
        RECT 110.195 117.640 113.260 117.780 ;
        RECT 110.195 117.595 110.485 117.640 ;
        RECT 108.890 117.440 109.030 117.595 ;
        RECT 111.100 117.580 111.420 117.640 ;
        RECT 112.940 117.580 113.260 117.640 ;
        RECT 110.640 117.440 110.960 117.500 ;
        RECT 111.575 117.440 111.865 117.485 ;
        RECT 104.750 117.300 110.410 117.440 ;
        RECT 102.820 117.240 103.140 117.300 ;
        RECT 104.215 117.255 104.505 117.300 ;
        RECT 106.055 117.100 106.345 117.145 ;
        RECT 98.770 116.960 106.345 117.100 ;
        RECT 106.055 116.915 106.345 116.960 ;
        RECT 107.420 117.100 107.740 117.160 ;
        RECT 109.260 117.100 109.580 117.160 ;
        RECT 107.420 116.960 109.580 117.100 ;
        RECT 110.270 117.100 110.410 117.300 ;
        RECT 110.640 117.300 111.865 117.440 ;
        RECT 110.640 117.240 110.960 117.300 ;
        RECT 111.575 117.255 111.865 117.300 ;
        RECT 112.020 117.440 112.340 117.500 ;
        RECT 115.240 117.440 115.560 117.500 ;
        RECT 112.020 117.300 115.560 117.440 ;
        RECT 112.020 117.240 112.340 117.300 ;
        RECT 115.240 117.240 115.560 117.300 ;
        RECT 119.840 117.100 120.160 117.160 ;
        RECT 110.270 116.960 120.160 117.100 ;
        RECT 107.420 116.900 107.740 116.960 ;
        RECT 109.260 116.900 109.580 116.960 ;
        RECT 119.840 116.900 120.160 116.960 ;
        RECT 97.300 116.620 98.450 116.760 ;
        RECT 99.600 116.760 99.920 116.820 ;
        RECT 100.520 116.760 100.840 116.820 ;
        RECT 99.600 116.620 100.840 116.760 ;
        RECT 97.300 116.560 97.620 116.620 ;
        RECT 99.600 116.560 99.920 116.620 ;
        RECT 100.520 116.560 100.840 116.620 ;
        RECT 101.440 116.760 101.760 116.820 ;
        RECT 102.820 116.760 103.140 116.820 ;
        RECT 101.440 116.620 103.140 116.760 ;
        RECT 101.440 116.560 101.760 116.620 ;
        RECT 102.820 116.560 103.140 116.620 ;
        RECT 106.960 116.760 107.280 116.820 ;
        RECT 112.020 116.760 112.340 116.820 ;
        RECT 106.960 116.620 112.340 116.760 ;
        RECT 106.960 116.560 107.280 116.620 ;
        RECT 112.020 116.560 112.340 116.620 ;
        RECT 118.920 116.760 119.240 116.820 ;
        RECT 120.300 116.760 120.620 116.820 ;
        RECT 118.920 116.620 120.620 116.760 ;
        RECT 118.920 116.560 119.240 116.620 ;
        RECT 120.300 116.560 120.620 116.620 ;
        RECT 53.990 115.940 125.290 116.420 ;
        RECT 69.715 115.740 70.005 115.785 ;
        RECT 77.520 115.740 77.840 115.800 ;
        RECT 91.320 115.740 91.640 115.800 ;
        RECT 97.775 115.740 98.065 115.785 ;
        RECT 99.140 115.740 99.460 115.800 ;
        RECT 69.715 115.600 77.840 115.740 ;
        RECT 69.715 115.555 70.005 115.600 ;
        RECT 77.520 115.540 77.840 115.600 ;
        RECT 87.090 115.600 91.640 115.740 ;
        RECT 70.160 115.400 70.480 115.460 ;
        RECT 57.830 115.260 70.480 115.400 ;
        RECT 55.900 115.060 56.220 115.120 ;
        RECT 57.830 115.060 57.970 115.260 ;
        RECT 70.160 115.200 70.480 115.260 ;
        RECT 75.220 115.400 75.540 115.460 ;
        RECT 87.090 115.400 87.230 115.600 ;
        RECT 91.320 115.540 91.640 115.600 ;
        RECT 91.870 115.600 94.770 115.740 ;
        RECT 75.220 115.260 87.230 115.400 ;
        RECT 87.655 115.400 87.945 115.445 ;
        RECT 89.020 115.400 89.340 115.460 ;
        RECT 87.655 115.260 89.340 115.400 ;
        RECT 75.220 115.200 75.540 115.260 ;
        RECT 87.655 115.215 87.945 115.260 ;
        RECT 89.020 115.200 89.340 115.260 ;
        RECT 90.415 115.215 90.705 115.445 ;
        RECT 90.860 115.400 91.180 115.460 ;
        RECT 91.870 115.400 92.010 115.600 ;
        RECT 90.860 115.260 92.010 115.400 ;
        RECT 93.635 115.400 93.925 115.445 ;
        RECT 94.080 115.400 94.400 115.460 ;
        RECT 93.635 115.260 94.400 115.400 ;
        RECT 94.630 115.400 94.770 115.600 ;
        RECT 97.775 115.600 99.460 115.740 ;
        RECT 97.775 115.555 98.065 115.600 ;
        RECT 99.140 115.540 99.460 115.600 ;
        RECT 100.520 115.740 100.840 115.800 ;
        RECT 101.455 115.740 101.745 115.785 ;
        RECT 100.520 115.600 101.745 115.740 ;
        RECT 100.520 115.540 100.840 115.600 ;
        RECT 101.455 115.555 101.745 115.600 ;
        RECT 103.755 115.740 104.045 115.785 ;
        RECT 106.040 115.740 106.360 115.800 ;
        RECT 109.260 115.740 109.580 115.800 ;
        RECT 103.755 115.600 106.360 115.740 ;
        RECT 103.755 115.555 104.045 115.600 ;
        RECT 106.040 115.540 106.360 115.600 ;
        RECT 107.050 115.600 109.580 115.740 ;
        RECT 94.630 115.260 104.430 115.400 ;
        RECT 55.900 114.920 57.970 115.060 ;
        RECT 55.900 114.860 56.220 114.920 ;
        RECT 57.280 114.520 57.600 114.780 ;
        RECT 57.830 114.765 57.970 114.920 ;
        RECT 58.660 114.860 58.980 115.120 ;
        RECT 60.500 115.060 60.820 115.120 ;
        RECT 79.360 115.060 79.680 115.120 ;
        RECT 90.490 115.060 90.630 115.215 ;
        RECT 90.860 115.200 91.180 115.260 ;
        RECT 93.635 115.215 93.925 115.260 ;
        RECT 94.080 115.200 94.400 115.260 ;
        RECT 60.500 114.920 79.680 115.060 ;
        RECT 60.500 114.860 60.820 114.920 ;
        RECT 79.360 114.860 79.680 114.920 ;
        RECT 87.730 114.920 90.630 115.060 ;
        RECT 91.320 115.060 91.640 115.120 ;
        RECT 99.140 115.060 99.460 115.120 ;
        RECT 91.320 114.920 95.230 115.060 ;
        RECT 57.755 114.535 58.045 114.765 ;
        RECT 59.135 114.720 59.425 114.765 ;
        RECT 63.720 114.720 64.040 114.780 ;
        RECT 59.135 114.580 64.040 114.720 ;
        RECT 59.135 114.535 59.425 114.580 ;
        RECT 63.720 114.520 64.040 114.580 ;
        RECT 64.640 114.520 64.960 114.780 ;
        RECT 67.400 114.520 67.720 114.780 ;
        RECT 68.795 114.535 69.085 114.765 ;
        RECT 72.000 114.720 72.320 114.780 ;
        RECT 74.315 114.720 74.605 114.765 ;
        RECT 72.000 114.580 74.605 114.720 ;
        RECT 64.730 114.380 64.870 114.520 ;
        RECT 68.870 114.380 69.010 114.535 ;
        RECT 72.000 114.520 72.320 114.580 ;
        RECT 74.315 114.535 74.605 114.580 ;
        RECT 75.235 114.720 75.525 114.765 ;
        RECT 77.980 114.720 78.300 114.780 ;
        RECT 87.730 114.765 87.870 114.920 ;
        RECT 91.320 114.860 91.640 114.920 ;
        RECT 75.235 114.580 78.300 114.720 ;
        RECT 75.235 114.535 75.525 114.580 ;
        RECT 77.980 114.520 78.300 114.580 ;
        RECT 87.655 114.535 87.945 114.765 ;
        RECT 89.020 114.520 89.340 114.780 ;
        RECT 91.780 114.520 92.100 114.780 ;
        RECT 95.090 114.765 95.230 114.920 ;
        RECT 97.390 114.920 99.460 115.060 ;
        RECT 94.555 114.720 94.845 114.765 ;
        RECT 94.170 114.580 94.845 114.720 ;
        RECT 64.730 114.240 69.010 114.380 ;
        RECT 90.400 114.180 90.720 114.440 ;
        RECT 92.240 114.180 92.560 114.440 ;
        RECT 94.170 114.380 94.310 114.580 ;
        RECT 94.555 114.535 94.845 114.580 ;
        RECT 95.015 114.535 95.305 114.765 ;
        RECT 95.475 114.535 95.765 114.765 ;
        RECT 95.920 114.720 96.240 114.780 ;
        RECT 97.390 114.765 97.530 114.920 ;
        RECT 99.140 114.860 99.460 114.920 ;
        RECT 99.600 115.060 99.920 115.120 ;
        RECT 99.600 114.920 102.130 115.060 ;
        RECT 99.600 114.860 99.920 114.920 ;
        RECT 96.395 114.720 96.685 114.765 ;
        RECT 95.920 114.580 96.685 114.720 ;
        RECT 95.550 114.380 95.690 114.535 ;
        RECT 95.920 114.520 96.240 114.580 ;
        RECT 96.395 114.535 96.685 114.580 ;
        RECT 97.315 114.535 97.605 114.765 ;
        RECT 98.220 114.720 98.540 114.780 ;
        RECT 98.695 114.720 98.985 114.765 ;
        RECT 98.220 114.580 98.985 114.720 ;
        RECT 98.220 114.520 98.540 114.580 ;
        RECT 98.695 114.535 98.985 114.580 ;
        RECT 100.060 114.520 100.380 114.780 ;
        RECT 100.520 114.520 100.840 114.780 ;
        RECT 94.170 114.240 94.770 114.380 ;
        RECT 95.550 114.240 96.150 114.380 ;
        RECT 56.375 114.040 56.665 114.085 ;
        RECT 64.640 114.040 64.960 114.100 ;
        RECT 56.375 113.900 64.960 114.040 ;
        RECT 56.375 113.855 56.665 113.900 ;
        RECT 64.640 113.840 64.960 113.900 ;
        RECT 66.480 114.040 66.800 114.100 ;
        RECT 67.875 114.040 68.165 114.085 ;
        RECT 66.480 113.900 68.165 114.040 ;
        RECT 66.480 113.840 66.800 113.900 ;
        RECT 67.875 113.855 68.165 113.900 ;
        RECT 74.760 113.840 75.080 114.100 ;
        RECT 80.280 114.040 80.600 114.100 ;
        RECT 87.640 114.040 87.960 114.100 ;
        RECT 88.575 114.040 88.865 114.085 ;
        RECT 80.280 113.900 88.865 114.040 ;
        RECT 80.280 113.840 80.600 113.900 ;
        RECT 87.640 113.840 87.960 113.900 ;
        RECT 88.575 113.855 88.865 113.900 ;
        RECT 89.480 114.040 89.800 114.100 ;
        RECT 89.940 114.040 90.260 114.100 ;
        RECT 89.480 113.900 90.260 114.040 ;
        RECT 89.480 113.840 89.800 113.900 ;
        RECT 89.940 113.840 90.260 113.900 ;
        RECT 91.320 113.840 91.640 114.100 ;
        RECT 92.330 114.040 92.470 114.180 ;
        RECT 94.080 114.040 94.400 114.100 ;
        RECT 92.330 113.900 94.400 114.040 ;
        RECT 94.630 114.040 94.770 114.240 ;
        RECT 96.010 114.100 96.150 114.240 ;
        RECT 99.140 114.180 99.460 114.440 ;
        RECT 99.615 114.380 99.905 114.425 ;
        RECT 100.150 114.380 100.290 114.520 ;
        RECT 99.615 114.240 100.290 114.380 ;
        RECT 101.990 114.380 102.130 114.920 ;
        RECT 102.375 114.780 102.665 114.845 ;
        RECT 102.360 114.520 102.680 114.780 ;
        RECT 102.820 114.520 103.140 114.780 ;
        RECT 103.740 114.520 104.060 114.780 ;
        RECT 104.290 114.765 104.430 115.260 ;
        RECT 105.580 114.860 105.900 115.120 ;
        RECT 107.050 115.060 107.190 115.600 ;
        RECT 109.260 115.540 109.580 115.600 ;
        RECT 110.180 115.540 110.500 115.800 ;
        RECT 110.640 115.740 110.960 115.800 ;
        RECT 113.400 115.740 113.720 115.800 ;
        RECT 110.640 115.600 113.720 115.740 ;
        RECT 110.640 115.540 110.960 115.600 ;
        RECT 113.400 115.540 113.720 115.600 ;
        RECT 116.635 115.740 116.925 115.785 ;
        RECT 118.000 115.740 118.320 115.800 ;
        RECT 116.635 115.600 118.320 115.740 ;
        RECT 116.635 115.555 116.925 115.600 ;
        RECT 118.000 115.540 118.320 115.600 ;
        RECT 119.395 115.740 119.685 115.785 ;
        RECT 119.840 115.740 120.160 115.800 ;
        RECT 119.395 115.600 120.160 115.740 ;
        RECT 119.395 115.555 119.685 115.600 ;
        RECT 119.840 115.540 120.160 115.600 ;
        RECT 121.680 115.740 122.000 115.800 ;
        RECT 124.900 115.740 125.220 115.800 ;
        RECT 121.680 115.600 125.220 115.740 ;
        RECT 121.680 115.540 122.000 115.600 ;
        RECT 124.900 115.540 125.220 115.600 ;
        RECT 107.880 115.200 108.200 115.460 ;
        RECT 110.730 115.400 110.870 115.540 ;
        RECT 114.780 115.400 115.100 115.460 ;
        RECT 109.810 115.260 110.870 115.400 ;
        RECT 111.190 115.260 115.100 115.400 ;
        RECT 106.590 114.920 107.190 115.060 ;
        RECT 109.275 115.060 109.565 115.105 ;
        RECT 109.810 115.060 109.950 115.260 ;
        RECT 110.640 115.105 110.960 115.120 ;
        RECT 111.190 115.105 111.330 115.260 ;
        RECT 114.780 115.200 115.100 115.260 ;
        RECT 115.240 115.400 115.560 115.460 ;
        RECT 115.240 115.260 122.370 115.400 ;
        RECT 115.240 115.200 115.560 115.260 ;
        RECT 109.275 114.920 109.950 115.060 ;
        RECT 106.590 114.765 106.730 114.920 ;
        RECT 109.275 114.875 109.565 114.920 ;
        RECT 110.615 114.875 110.960 115.105 ;
        RECT 111.115 114.875 111.405 115.105 ;
        RECT 120.300 115.060 120.620 115.120 ;
        RECT 121.680 115.060 122.000 115.120 ;
        RECT 114.870 114.920 120.620 115.060 ;
        RECT 110.640 114.860 110.960 114.875 ;
        RECT 104.215 114.535 104.505 114.765 ;
        RECT 106.515 114.535 106.805 114.765 ;
        RECT 107.420 114.520 107.740 114.780 ;
        RECT 108.355 114.535 108.645 114.765 ;
        RECT 104.675 114.380 104.965 114.425 ;
        RECT 108.430 114.380 108.570 114.535 ;
        RECT 112.020 114.520 112.340 114.780 ;
        RECT 112.480 114.520 112.800 114.780 ;
        RECT 113.415 114.535 113.705 114.765 ;
        RECT 113.860 114.720 114.180 114.780 ;
        RECT 114.870 114.765 115.010 114.920 ;
        RECT 120.300 114.860 120.620 114.920 ;
        RECT 120.850 114.920 122.000 115.060 ;
        RECT 114.795 114.720 115.085 114.765 ;
        RECT 113.860 114.580 115.085 114.720 ;
        RECT 113.490 114.380 113.630 114.535 ;
        RECT 113.860 114.520 114.180 114.580 ;
        RECT 114.795 114.535 115.085 114.580 ;
        RECT 117.095 114.535 117.385 114.765 ;
        RECT 119.855 114.720 120.145 114.765 ;
        RECT 120.850 114.720 120.990 114.920 ;
        RECT 121.680 114.860 122.000 114.920 ;
        RECT 119.855 114.580 120.990 114.720 ;
        RECT 119.855 114.535 120.145 114.580 ;
        RECT 101.990 114.240 113.630 114.380 ;
        RECT 117.170 114.380 117.310 114.535 ;
        RECT 121.220 114.520 121.540 114.780 ;
        RECT 122.230 114.765 122.370 115.260 ;
        RECT 122.155 114.535 122.445 114.765 ;
        RECT 124.440 114.380 124.760 114.440 ;
        RECT 117.170 114.240 124.760 114.380 ;
        RECT 99.615 114.195 99.905 114.240 ;
        RECT 104.675 114.195 104.965 114.240 ;
        RECT 124.440 114.180 124.760 114.240 ;
        RECT 95.460 114.040 95.780 114.100 ;
        RECT 94.630 113.900 95.780 114.040 ;
        RECT 94.080 113.840 94.400 113.900 ;
        RECT 95.460 113.840 95.780 113.900 ;
        RECT 95.920 113.840 96.240 114.100 ;
        RECT 96.840 113.840 97.160 114.100 ;
        RECT 97.760 114.040 98.080 114.100 ;
        RECT 102.820 114.040 103.140 114.100 ;
        RECT 97.760 113.900 103.140 114.040 ;
        RECT 97.760 113.840 98.080 113.900 ;
        RECT 102.820 113.840 103.140 113.900 ;
        RECT 106.040 114.040 106.360 114.100 ;
        RECT 108.815 114.040 109.105 114.085 ;
        RECT 112.955 114.040 113.245 114.085 ;
        RECT 106.040 113.900 113.245 114.040 ;
        RECT 106.040 113.840 106.360 113.900 ;
        RECT 108.815 113.855 109.105 113.900 ;
        RECT 112.955 113.855 113.245 113.900 ;
        RECT 113.875 114.040 114.165 114.085 ;
        RECT 122.600 114.040 122.920 114.100 ;
        RECT 113.875 113.900 122.920 114.040 ;
        RECT 113.875 113.855 114.165 113.900 ;
        RECT 122.600 113.840 122.920 113.900 ;
        RECT 123.060 113.840 123.380 114.100 ;
        RECT 53.990 113.220 125.290 113.700 ;
        RECT 57.755 113.020 58.045 113.065 ;
        RECT 58.660 113.020 58.980 113.080 ;
        RECT 57.755 112.880 58.980 113.020 ;
        RECT 57.755 112.835 58.045 112.880 ;
        RECT 58.660 112.820 58.980 112.880 ;
        RECT 59.580 112.820 59.900 113.080 ;
        RECT 65.115 113.020 65.405 113.065 ;
        RECT 66.480 113.020 66.800 113.080 ;
        RECT 65.115 112.880 66.800 113.020 ;
        RECT 65.115 112.835 65.405 112.880 ;
        RECT 66.480 112.820 66.800 112.880 ;
        RECT 67.400 113.020 67.720 113.080 ;
        RECT 71.555 113.020 71.845 113.065 ;
        RECT 67.400 112.880 71.845 113.020 ;
        RECT 67.400 112.820 67.720 112.880 ;
        RECT 71.555 112.835 71.845 112.880 ;
        RECT 74.760 113.020 75.080 113.080 ;
        RECT 75.235 113.020 75.525 113.065 ;
        RECT 74.760 112.880 75.525 113.020 ;
        RECT 74.760 112.820 75.080 112.880 ;
        RECT 75.235 112.835 75.525 112.880 ;
        RECT 80.280 113.020 80.600 113.080 ;
        RECT 80.755 113.020 81.045 113.065 ;
        RECT 80.280 112.880 81.045 113.020 ;
        RECT 80.280 112.820 80.600 112.880 ;
        RECT 80.755 112.835 81.045 112.880 ;
        RECT 82.120 113.020 82.440 113.080 ;
        RECT 82.595 113.020 82.885 113.065 ;
        RECT 92.700 113.020 93.020 113.080 ;
        RECT 82.120 112.880 82.885 113.020 ;
        RECT 82.120 112.820 82.440 112.880 ;
        RECT 82.595 112.835 82.885 112.880 ;
        RECT 84.050 112.880 93.020 113.020 ;
        RECT 63.720 112.680 64.040 112.740 ;
        RECT 81.675 112.680 81.965 112.725 ;
        RECT 63.720 112.540 69.110 112.680 ;
        RECT 63.720 112.480 64.040 112.540 ;
        RECT 64.640 112.140 64.960 112.400 ;
        RECT 65.100 112.340 65.420 112.400 ;
        RECT 66.035 112.340 66.325 112.385 ;
        RECT 65.100 112.200 66.325 112.340 ;
        RECT 65.100 112.140 65.420 112.200 ;
        RECT 66.035 112.155 66.325 112.200 ;
        RECT 67.400 112.140 67.720 112.400 ;
        RECT 68.225 112.140 68.545 112.400 ;
        RECT 68.970 112.385 69.110 112.540 ;
        RECT 73.930 112.540 81.965 112.680 ;
        RECT 68.795 112.200 69.110 112.385 ;
        RECT 68.795 112.155 69.085 112.200 ;
        RECT 70.160 112.140 70.480 112.400 ;
        RECT 70.635 112.340 70.925 112.385 ;
        RECT 72.920 112.340 73.240 112.400 ;
        RECT 70.635 112.200 73.240 112.340 ;
        RECT 70.635 112.155 70.925 112.200 ;
        RECT 72.920 112.140 73.240 112.200 ;
        RECT 60.040 111.800 60.360 112.060 ;
        RECT 60.500 111.800 60.820 112.060 ;
        RECT 73.930 112.000 74.070 112.540 ;
        RECT 81.675 112.495 81.965 112.540 ;
        RECT 74.775 112.340 75.065 112.385 ;
        RECT 77.060 112.340 77.380 112.400 ;
        RECT 74.775 112.200 77.380 112.340 ;
        RECT 74.775 112.155 75.065 112.200 ;
        RECT 77.060 112.140 77.380 112.200 ;
        RECT 79.360 112.340 79.680 112.400 ;
        RECT 80.295 112.340 80.585 112.385 ;
        RECT 79.360 112.200 80.585 112.340 ;
        RECT 79.360 112.140 79.680 112.200 ;
        RECT 80.295 112.155 80.585 112.200 ;
        RECT 83.040 112.340 83.360 112.400 ;
        RECT 83.515 112.340 83.805 112.385 ;
        RECT 83.040 112.200 83.805 112.340 ;
        RECT 83.040 112.140 83.360 112.200 ;
        RECT 83.515 112.155 83.805 112.200 ;
        RECT 66.110 111.860 74.070 112.000 ;
        RECT 75.220 112.000 75.540 112.060 ;
        RECT 75.695 112.000 75.985 112.045 ;
        RECT 75.220 111.860 75.985 112.000 ;
        RECT 66.110 111.705 66.250 111.860 ;
        RECT 75.220 111.800 75.540 111.860 ;
        RECT 75.695 111.815 75.985 111.860 ;
        RECT 76.140 112.000 76.460 112.060 ;
        RECT 82.580 112.000 82.900 112.060 ;
        RECT 76.140 111.860 82.900 112.000 ;
        RECT 76.140 111.800 76.460 111.860 ;
        RECT 82.580 111.800 82.900 111.860 ;
        RECT 66.035 111.475 66.325 111.705 ;
        RECT 69.255 111.660 69.545 111.705 ;
        RECT 72.935 111.660 73.225 111.705 ;
        RECT 69.255 111.520 73.225 111.660 ;
        RECT 69.255 111.475 69.545 111.520 ;
        RECT 72.935 111.475 73.225 111.520 ;
        RECT 81.675 111.660 81.965 111.705 ;
        RECT 84.050 111.660 84.190 112.880 ;
        RECT 92.700 112.820 93.020 112.880 ;
        RECT 93.620 112.820 93.940 113.080 ;
        RECT 94.080 113.020 94.400 113.080 ;
        RECT 100.075 113.020 100.365 113.065 ;
        RECT 104.200 113.020 104.520 113.080 ;
        RECT 94.080 112.880 100.365 113.020 ;
        RECT 94.080 112.820 94.400 112.880 ;
        RECT 100.075 112.835 100.365 112.880 ;
        RECT 101.070 112.880 104.520 113.020 ;
        RECT 84.435 112.680 84.725 112.725 ;
        RECT 88.560 112.680 88.880 112.740 ;
        RECT 84.435 112.540 88.880 112.680 ;
        RECT 84.435 112.495 84.725 112.540 ;
        RECT 88.560 112.480 88.880 112.540 ;
        RECT 89.035 112.680 89.325 112.725 ;
        RECT 89.940 112.680 90.260 112.740 ;
        RECT 89.035 112.540 90.260 112.680 ;
        RECT 89.035 112.495 89.325 112.540 ;
        RECT 89.940 112.480 90.260 112.540 ;
        RECT 90.400 112.680 90.720 112.740 ;
        RECT 90.875 112.680 91.165 112.725 ;
        RECT 90.400 112.540 91.165 112.680 ;
        RECT 90.400 112.480 90.720 112.540 ;
        RECT 90.875 112.495 91.165 112.540 ;
        RECT 84.880 112.140 85.200 112.400 ;
        RECT 88.115 112.155 88.405 112.385 ;
        RECT 88.190 112.000 88.330 112.155 ;
        RECT 89.480 112.140 89.800 112.400 ;
        RECT 91.780 112.140 92.100 112.400 ;
        RECT 92.255 112.155 92.545 112.385 ;
        RECT 92.330 112.000 92.470 112.155 ;
        RECT 94.540 112.140 94.860 112.400 ;
        RECT 95.920 112.140 96.240 112.400 ;
        RECT 96.395 112.340 96.685 112.385 ;
        RECT 96.840 112.340 97.160 112.400 ;
        RECT 96.395 112.200 97.160 112.340 ;
        RECT 96.395 112.155 96.685 112.200 ;
        RECT 96.840 112.140 97.160 112.200 ;
        RECT 98.695 112.340 98.985 112.385 ;
        RECT 99.600 112.340 99.920 112.400 ;
        RECT 101.070 112.385 101.210 112.880 ;
        RECT 104.200 112.820 104.520 112.880 ;
        RECT 105.135 112.835 105.425 113.065 ;
        RECT 107.435 113.020 107.725 113.065 ;
        RECT 118.460 113.020 118.780 113.080 ;
        RECT 107.435 112.880 118.780 113.020 ;
        RECT 107.435 112.835 107.725 112.880 ;
        RECT 104.660 112.680 104.980 112.740 ;
        RECT 101.530 112.540 104.980 112.680 ;
        RECT 105.210 112.680 105.350 112.835 ;
        RECT 118.460 112.820 118.780 112.880 ;
        RECT 119.380 113.020 119.700 113.080 ;
        RECT 121.235 113.020 121.525 113.065 ;
        RECT 119.380 112.880 121.525 113.020 ;
        RECT 119.380 112.820 119.700 112.880 ;
        RECT 121.235 112.835 121.525 112.880 ;
        RECT 107.880 112.680 108.200 112.740 ;
        RECT 113.860 112.680 114.180 112.740 ;
        RECT 105.210 112.540 108.200 112.680 ;
        RECT 101.530 112.385 101.670 112.540 ;
        RECT 104.660 112.480 104.980 112.540 ;
        RECT 107.880 112.480 108.200 112.540 ;
        RECT 108.890 112.540 114.180 112.680 ;
        RECT 98.695 112.200 99.920 112.340 ;
        RECT 98.695 112.155 98.985 112.200 ;
        RECT 99.600 112.140 99.920 112.200 ;
        RECT 100.995 112.155 101.285 112.385 ;
        RECT 101.455 112.155 101.745 112.385 ;
        RECT 103.740 112.140 104.060 112.400 ;
        RECT 104.215 112.340 104.505 112.385 ;
        RECT 105.580 112.340 105.900 112.400 ;
        RECT 104.215 112.200 105.900 112.340 ;
        RECT 104.215 112.155 104.505 112.200 ;
        RECT 105.580 112.140 105.900 112.200 ;
        RECT 106.500 112.140 106.820 112.400 ;
        RECT 108.890 112.385 109.030 112.540 ;
        RECT 113.860 112.480 114.180 112.540 ;
        RECT 108.815 112.155 109.105 112.385 ;
        RECT 109.260 112.140 109.580 112.400 ;
        RECT 109.720 112.340 110.040 112.400 ;
        RECT 110.195 112.340 110.485 112.385 ;
        RECT 109.720 112.200 110.485 112.340 ;
        RECT 109.720 112.140 110.040 112.200 ;
        RECT 110.195 112.155 110.485 112.200 ;
        RECT 111.575 112.340 111.865 112.385 ;
        RECT 112.480 112.340 112.800 112.400 ;
        RECT 111.575 112.200 112.800 112.340 ;
        RECT 111.575 112.155 111.865 112.200 ;
        RECT 112.480 112.140 112.800 112.200 ;
        RECT 112.955 112.360 113.245 112.385 ;
        RECT 112.955 112.220 113.630 112.360 ;
        RECT 112.955 112.155 113.245 112.220 ;
        RECT 95.015 112.000 95.305 112.045 ;
        RECT 88.190 111.860 91.090 112.000 ;
        RECT 92.330 111.860 95.305 112.000 ;
        RECT 81.675 111.520 84.190 111.660 ;
        RECT 84.510 111.520 87.870 111.660 ;
        RECT 81.675 111.475 81.965 111.520 ;
        RECT 70.160 111.320 70.480 111.380 ;
        RECT 73.380 111.320 73.700 111.380 ;
        RECT 70.160 111.180 73.700 111.320 ;
        RECT 70.160 111.120 70.480 111.180 ;
        RECT 73.380 111.120 73.700 111.180 ;
        RECT 75.680 111.320 76.000 111.380 ;
        RECT 82.120 111.320 82.440 111.380 ;
        RECT 75.680 111.180 82.440 111.320 ;
        RECT 75.680 111.120 76.000 111.180 ;
        RECT 82.120 111.120 82.440 111.180 ;
        RECT 82.580 111.320 82.900 111.380 ;
        RECT 84.510 111.320 84.650 111.520 ;
        RECT 82.580 111.180 84.650 111.320 ;
        RECT 87.730 111.320 87.870 111.520 ;
        RECT 88.100 111.460 88.420 111.720 ;
        RECT 90.950 111.705 91.090 111.860 ;
        RECT 95.015 111.815 95.305 111.860 ;
        RECT 97.300 112.000 97.620 112.060 ;
        RECT 98.235 112.000 98.525 112.045 ;
        RECT 113.490 112.000 113.630 112.220 ;
        RECT 114.320 112.340 114.640 112.400 ;
        RECT 114.795 112.340 115.085 112.385 ;
        RECT 114.320 112.200 115.085 112.340 ;
        RECT 114.320 112.140 114.640 112.200 ;
        RECT 114.795 112.155 115.085 112.200 ;
        RECT 97.300 111.860 98.525 112.000 ;
        RECT 97.300 111.800 97.620 111.860 ;
        RECT 98.235 111.815 98.525 111.860 ;
        RECT 99.690 111.860 113.630 112.000 ;
        RECT 90.875 111.475 91.165 111.705 ;
        RECT 97.760 111.660 98.080 111.720 ;
        RECT 99.690 111.705 99.830 111.860 ;
        RECT 91.410 111.520 98.080 111.660 ;
        RECT 91.410 111.320 91.550 111.520 ;
        RECT 97.760 111.460 98.080 111.520 ;
        RECT 99.615 111.475 99.905 111.705 ;
        RECT 100.520 111.660 100.840 111.720 ;
        RECT 101.900 111.660 102.220 111.720 ;
        RECT 100.520 111.520 102.220 111.660 ;
        RECT 100.520 111.460 100.840 111.520 ;
        RECT 101.900 111.460 102.220 111.520 ;
        RECT 102.820 111.460 103.140 111.720 ;
        RECT 111.560 111.660 111.880 111.720 ;
        RECT 103.370 111.520 111.880 111.660 ;
        RECT 87.730 111.180 91.550 111.320 ;
        RECT 102.375 111.320 102.665 111.365 ;
        RECT 103.370 111.320 103.510 111.520 ;
        RECT 111.560 111.460 111.880 111.520 ;
        RECT 112.020 111.660 112.340 111.720 ;
        RECT 112.495 111.660 112.785 111.705 ;
        RECT 112.020 111.520 112.785 111.660 ;
        RECT 112.020 111.460 112.340 111.520 ;
        RECT 112.495 111.475 112.785 111.520 ;
        RECT 113.860 111.460 114.180 111.720 ;
        RECT 102.375 111.180 103.510 111.320 ;
        RECT 82.580 111.120 82.900 111.180 ;
        RECT 102.375 111.135 102.665 111.180 ;
        RECT 53.990 110.500 125.290 110.980 ;
        RECT 57.280 110.100 57.600 110.360 ;
        RECT 69.240 110.300 69.560 110.360 ;
        RECT 62.200 110.160 69.560 110.300 ;
        RECT 59.580 109.420 59.900 109.680 ;
        RECT 60.055 109.620 60.345 109.665 ;
        RECT 60.500 109.620 60.820 109.680 ;
        RECT 62.200 109.620 62.340 110.160 ;
        RECT 69.240 110.100 69.560 110.160 ;
        RECT 71.095 110.300 71.385 110.345 ;
        RECT 71.540 110.300 71.860 110.360 ;
        RECT 71.095 110.160 71.860 110.300 ;
        RECT 71.095 110.115 71.385 110.160 ;
        RECT 71.540 110.100 71.860 110.160 ;
        RECT 72.475 110.300 72.765 110.345 ;
        RECT 72.920 110.300 73.240 110.360 ;
        RECT 72.475 110.160 73.240 110.300 ;
        RECT 72.475 110.115 72.765 110.160 ;
        RECT 72.920 110.100 73.240 110.160 ;
        RECT 73.840 110.300 74.160 110.360 ;
        RECT 78.900 110.300 79.220 110.360 ;
        RECT 82.580 110.300 82.900 110.360 ;
        RECT 73.840 110.160 82.900 110.300 ;
        RECT 73.840 110.100 74.160 110.160 ;
        RECT 78.900 110.100 79.220 110.160 ;
        RECT 82.580 110.100 82.900 110.160 ;
        RECT 84.880 110.300 85.200 110.360 ;
        RECT 85.355 110.300 85.645 110.345 ;
        RECT 84.880 110.160 85.645 110.300 ;
        RECT 84.880 110.100 85.200 110.160 ;
        RECT 85.355 110.115 85.645 110.160 ;
        RECT 94.080 110.100 94.400 110.360 ;
        RECT 100.980 110.300 101.300 110.360 ;
        RECT 111.115 110.300 111.405 110.345 ;
        RECT 100.980 110.160 111.405 110.300 ;
        RECT 100.980 110.100 101.300 110.160 ;
        RECT 111.115 110.115 111.405 110.160 ;
        RECT 65.575 109.960 65.865 110.005 ;
        RECT 66.940 109.960 67.260 110.020 ;
        RECT 65.575 109.820 67.260 109.960 ;
        RECT 65.575 109.775 65.865 109.820 ;
        RECT 66.940 109.760 67.260 109.820 ;
        RECT 67.400 109.960 67.720 110.020 ;
        RECT 67.400 109.820 76.370 109.960 ;
        RECT 67.400 109.760 67.720 109.820 ;
        RECT 60.055 109.480 62.340 109.620 ;
        RECT 60.055 109.435 60.345 109.480 ;
        RECT 59.120 109.280 59.440 109.340 ;
        RECT 60.130 109.280 60.270 109.435 ;
        RECT 60.500 109.420 60.820 109.480 ;
        RECT 74.760 109.420 75.080 109.680 ;
        RECT 75.680 109.420 76.000 109.680 ;
        RECT 59.120 109.140 60.270 109.280 ;
        RECT 64.195 109.280 64.485 109.325 ;
        RECT 65.100 109.280 65.420 109.340 ;
        RECT 64.195 109.140 65.420 109.280 ;
        RECT 59.120 109.080 59.440 109.140 ;
        RECT 64.195 109.095 64.485 109.140 ;
        RECT 65.100 109.080 65.420 109.140 ;
        RECT 65.560 109.080 65.880 109.340 ;
        RECT 67.400 109.280 67.720 109.340 ;
        RECT 68.335 109.280 68.625 109.325 ;
        RECT 67.400 109.140 68.625 109.280 ;
        RECT 67.400 109.080 67.720 109.140 ;
        RECT 68.335 109.095 68.625 109.140 ;
        RECT 69.240 109.080 69.560 109.340 ;
        RECT 69.715 109.280 70.005 109.325 ;
        RECT 71.540 109.280 71.860 109.340 ;
        RECT 69.715 109.140 71.860 109.280 ;
        RECT 69.715 109.095 70.005 109.140 ;
        RECT 71.540 109.080 71.860 109.140 ;
        RECT 76.230 109.290 76.370 109.820 ;
        RECT 76.600 109.760 76.920 110.020 ;
        RECT 78.440 109.960 78.760 110.020 ;
        RECT 81.675 109.960 81.965 110.005 ;
        RECT 86.720 109.960 87.040 110.020 ;
        RECT 78.440 109.820 79.590 109.960 ;
        RECT 78.440 109.760 78.760 109.820 ;
        RECT 76.690 109.620 76.830 109.760 ;
        RECT 76.690 109.480 78.210 109.620 ;
        RECT 78.070 109.335 78.210 109.480 ;
        RECT 76.575 109.290 76.865 109.335 ;
        RECT 76.230 109.105 76.865 109.290 ;
        RECT 77.995 109.105 78.285 109.335 ;
        RECT 76.230 109.090 76.830 109.105 ;
        RECT 65.650 108.940 65.790 109.080 ;
        RECT 68.780 108.940 69.100 109.000 ;
        RECT 71.095 108.940 71.385 108.985 ;
        RECT 65.650 108.800 71.385 108.940 ;
        RECT 68.780 108.740 69.100 108.800 ;
        RECT 71.095 108.755 71.385 108.800 ;
        RECT 57.280 108.600 57.600 108.660 ;
        RECT 59.135 108.600 59.425 108.645 ;
        RECT 60.040 108.600 60.360 108.660 ;
        RECT 57.280 108.460 60.360 108.600 ;
        RECT 57.280 108.400 57.600 108.460 ;
        RECT 59.135 108.415 59.425 108.460 ;
        RECT 60.040 108.400 60.360 108.460 ;
        RECT 64.655 108.600 64.945 108.645 ;
        RECT 67.415 108.600 67.705 108.645 ;
        RECT 70.175 108.600 70.465 108.645 ;
        RECT 64.655 108.460 70.465 108.600 ;
        RECT 64.655 108.415 64.945 108.460 ;
        RECT 67.415 108.415 67.705 108.460 ;
        RECT 70.175 108.415 70.465 108.460 ;
        RECT 73.840 108.600 74.160 108.660 ;
        RECT 74.315 108.600 74.605 108.645 ;
        RECT 73.840 108.460 74.605 108.600 ;
        RECT 76.690 108.600 76.830 109.090 ;
        RECT 78.900 109.080 79.220 109.340 ;
        RECT 77.075 108.940 77.365 108.985 ;
        RECT 79.450 108.940 79.590 109.820 ;
        RECT 81.675 109.820 87.040 109.960 ;
        RECT 81.675 109.775 81.965 109.820 ;
        RECT 86.720 109.760 87.040 109.820 ;
        RECT 89.020 109.960 89.340 110.020 ;
        RECT 101.915 109.960 102.205 110.005 ;
        RECT 89.020 109.820 102.205 109.960 ;
        RECT 89.020 109.760 89.340 109.820 ;
        RECT 101.915 109.775 102.205 109.820 ;
        RECT 102.820 109.760 103.140 110.020 ;
        RECT 106.975 109.960 107.265 110.005 ;
        RECT 105.210 109.820 107.265 109.960 ;
        RECT 79.820 109.620 80.140 109.680 ;
        RECT 97.760 109.620 98.080 109.680 ;
        RECT 99.140 109.620 99.460 109.680 ;
        RECT 79.820 109.480 85.110 109.620 ;
        RECT 79.820 109.420 80.140 109.480 ;
        RECT 80.280 109.080 80.600 109.340 ;
        RECT 80.830 109.325 80.970 109.480 ;
        RECT 80.755 109.095 81.045 109.325 ;
        RECT 82.120 109.080 82.440 109.340 ;
        RECT 84.970 109.325 85.110 109.480 ;
        RECT 97.760 109.480 100.290 109.620 ;
        RECT 97.760 109.420 98.080 109.480 ;
        RECT 99.140 109.420 99.460 109.480 ;
        RECT 84.895 109.095 85.185 109.325 ;
        RECT 85.815 109.280 86.105 109.325 ;
        RECT 86.260 109.280 86.580 109.340 ;
        RECT 94.540 109.280 94.860 109.340 ;
        RECT 85.815 109.140 86.580 109.280 ;
        RECT 85.815 109.095 86.105 109.140 ;
        RECT 86.260 109.080 86.580 109.140 ;
        RECT 86.810 109.140 94.860 109.280 ;
        RECT 81.675 108.940 81.965 108.985 ;
        RECT 77.075 108.800 78.670 108.940 ;
        RECT 79.450 108.800 81.965 108.940 ;
        RECT 77.075 108.755 77.365 108.800 ;
        RECT 77.995 108.600 78.285 108.645 ;
        RECT 76.690 108.460 78.285 108.600 ;
        RECT 78.530 108.600 78.670 108.800 ;
        RECT 81.675 108.755 81.965 108.800 ;
        RECT 81.200 108.600 81.520 108.660 ;
        RECT 78.530 108.460 81.520 108.600 ;
        RECT 82.210 108.600 82.350 109.080 ;
        RECT 82.595 108.940 82.885 108.985 ;
        RECT 83.040 108.940 83.360 109.000 ;
        RECT 86.810 108.940 86.950 109.140 ;
        RECT 94.540 109.080 94.860 109.140 ;
        RECT 95.920 109.080 96.240 109.340 ;
        RECT 100.150 109.325 100.290 109.480 ;
        RECT 99.615 109.095 99.905 109.325 ;
        RECT 100.075 109.095 100.365 109.325 ;
        RECT 82.595 108.800 86.950 108.940 ;
        RECT 89.480 108.940 89.800 109.000 ;
        RECT 98.695 108.940 98.985 108.985 ;
        RECT 89.480 108.800 98.985 108.940 ;
        RECT 99.690 108.940 99.830 109.095 ;
        RECT 100.980 109.080 101.300 109.340 ;
        RECT 101.440 109.080 101.760 109.340 ;
        RECT 102.910 109.325 103.050 109.760 ;
        RECT 102.810 109.095 103.100 109.325 ;
        RECT 103.280 109.080 103.600 109.340 ;
        RECT 104.660 109.280 104.980 109.340 ;
        RECT 105.210 109.325 105.350 109.820 ;
        RECT 106.975 109.775 107.265 109.820 ;
        RECT 109.260 109.960 109.580 110.020 ;
        RECT 109.735 109.960 110.025 110.005 ;
        RECT 113.400 109.960 113.720 110.020 ;
        RECT 109.260 109.820 113.720 109.960 ;
        RECT 109.260 109.760 109.580 109.820 ;
        RECT 109.735 109.775 110.025 109.820 ;
        RECT 113.400 109.760 113.720 109.820 ;
        RECT 114.320 109.760 114.640 110.020 ;
        RECT 106.500 109.620 106.820 109.680 ;
        RECT 118.935 109.620 119.225 109.665 ;
        RECT 120.760 109.620 121.080 109.680 ;
        RECT 106.500 109.480 119.225 109.620 ;
        RECT 106.500 109.420 106.820 109.480 ;
        RECT 118.935 109.435 119.225 109.480 ;
        RECT 119.930 109.480 121.080 109.620 ;
        RECT 104.465 109.140 104.980 109.280 ;
        RECT 104.660 109.080 104.980 109.140 ;
        RECT 105.135 109.095 105.425 109.325 ;
        RECT 105.580 109.130 105.900 109.390 ;
        RECT 107.880 109.280 108.200 109.340 ;
        RECT 108.815 109.280 109.105 109.325 ;
        RECT 107.880 109.140 109.105 109.280 ;
        RECT 107.880 109.080 108.200 109.140 ;
        RECT 108.815 109.095 109.105 109.140 ;
        RECT 109.275 109.280 109.565 109.325 ;
        RECT 109.720 109.280 110.040 109.340 ;
        RECT 109.275 109.140 110.040 109.280 ;
        RECT 109.275 109.095 109.565 109.140 ;
        RECT 109.720 109.080 110.040 109.140 ;
        RECT 110.195 109.280 110.485 109.325 ;
        RECT 110.640 109.280 110.960 109.340 ;
        RECT 110.195 109.140 110.960 109.280 ;
        RECT 110.195 109.095 110.485 109.140 ;
        RECT 110.640 109.080 110.960 109.140 ;
        RECT 112.480 109.280 112.800 109.340 ;
        RECT 119.930 109.325 120.070 109.480 ;
        RECT 120.760 109.420 121.080 109.480 ;
        RECT 112.480 109.140 117.310 109.280 ;
        RECT 112.480 109.080 112.800 109.140 ;
        RECT 103.755 108.940 104.045 108.985 ;
        RECT 99.690 108.800 106.730 108.940 ;
        RECT 82.595 108.755 82.885 108.800 ;
        RECT 83.040 108.740 83.360 108.800 ;
        RECT 89.480 108.740 89.800 108.800 ;
        RECT 98.695 108.755 98.985 108.800 ;
        RECT 103.755 108.755 104.045 108.800 ;
        RECT 89.020 108.600 89.340 108.660 ;
        RECT 82.210 108.460 89.340 108.600 ;
        RECT 73.840 108.400 74.160 108.460 ;
        RECT 74.315 108.415 74.605 108.460 ;
        RECT 77.995 108.415 78.285 108.460 ;
        RECT 81.200 108.400 81.520 108.460 ;
        RECT 89.020 108.400 89.340 108.460 ;
        RECT 90.860 108.600 91.180 108.660 ;
        RECT 93.175 108.600 93.465 108.645 ;
        RECT 90.860 108.460 93.465 108.600 ;
        RECT 90.860 108.400 91.180 108.460 ;
        RECT 93.175 108.415 93.465 108.460 ;
        RECT 102.820 108.600 103.140 108.660 ;
        RECT 106.055 108.600 106.345 108.645 ;
        RECT 102.820 108.460 106.345 108.600 ;
        RECT 106.590 108.600 106.730 108.800 ;
        RECT 106.960 108.740 107.280 109.000 ;
        RECT 113.415 108.940 113.705 108.985 ;
        RECT 113.860 108.940 114.180 109.000 ;
        RECT 113.415 108.800 114.180 108.940 ;
        RECT 113.415 108.755 113.705 108.800 ;
        RECT 113.860 108.740 114.180 108.800 ;
        RECT 116.160 108.940 116.480 109.000 ;
        RECT 116.635 108.940 116.925 108.985 ;
        RECT 116.160 108.800 116.925 108.940 ;
        RECT 117.170 108.940 117.310 109.140 ;
        RECT 119.855 109.095 120.145 109.325 ;
        RECT 120.300 109.080 120.620 109.340 ;
        RECT 121.695 108.940 121.985 108.985 ;
        RECT 117.170 108.800 121.985 108.940 ;
        RECT 116.160 108.740 116.480 108.800 ;
        RECT 116.635 108.755 116.925 108.800 ;
        RECT 121.695 108.755 121.985 108.800 ;
        RECT 111.560 108.600 111.880 108.660 ;
        RECT 106.590 108.460 111.880 108.600 ;
        RECT 102.820 108.400 103.140 108.460 ;
        RECT 106.055 108.415 106.345 108.460 ;
        RECT 111.560 108.400 111.880 108.460 ;
        RECT 53.990 107.780 125.290 108.260 ;
        RECT 58.200 107.580 58.520 107.640 ;
        RECT 59.595 107.580 59.885 107.625 ;
        RECT 58.200 107.440 59.885 107.580 ;
        RECT 58.200 107.380 58.520 107.440 ;
        RECT 59.595 107.395 59.885 107.440 ;
        RECT 65.100 107.380 65.420 107.640 ;
        RECT 69.240 107.580 69.560 107.640 ;
        RECT 75.680 107.580 76.000 107.640 ;
        RECT 69.240 107.440 76.000 107.580 ;
        RECT 69.240 107.380 69.560 107.440 ;
        RECT 75.680 107.380 76.000 107.440 ;
        RECT 83.500 107.380 83.820 107.640 ;
        RECT 84.420 107.380 84.740 107.640 ;
        RECT 88.560 107.580 88.880 107.640 ;
        RECT 89.035 107.580 89.325 107.625 ;
        RECT 91.320 107.580 91.640 107.640 ;
        RECT 97.775 107.580 98.065 107.625 ;
        RECT 104.200 107.580 104.520 107.640 ;
        RECT 88.560 107.440 89.325 107.580 ;
        RECT 88.560 107.380 88.880 107.440 ;
        RECT 89.035 107.395 89.325 107.440 ;
        RECT 90.030 107.440 98.065 107.580 ;
        RECT 74.760 107.240 75.080 107.300 ;
        RECT 62.430 107.100 75.080 107.240 ;
        RECT 59.580 106.900 59.900 106.960 ;
        RECT 62.430 106.945 62.570 107.100 ;
        RECT 74.760 107.040 75.080 107.100 ;
        RECT 60.055 106.900 60.345 106.945 ;
        RECT 59.580 106.760 60.345 106.900 ;
        RECT 59.580 106.700 59.900 106.760 ;
        RECT 60.055 106.715 60.345 106.760 ;
        RECT 62.355 106.715 62.645 106.945 ;
        RECT 63.720 106.700 64.040 106.960 ;
        RECT 64.180 106.700 64.500 106.960 ;
        RECT 79.820 106.900 80.140 106.960 ;
        RECT 90.030 106.945 90.170 107.440 ;
        RECT 91.320 107.380 91.640 107.440 ;
        RECT 97.775 107.395 98.065 107.440 ;
        RECT 102.450 107.440 104.520 107.580 ;
        RECT 90.400 107.240 90.720 107.300 ;
        RECT 96.840 107.240 97.160 107.300 ;
        RECT 102.450 107.285 102.590 107.440 ;
        RECT 104.200 107.380 104.520 107.440 ;
        RECT 105.135 107.580 105.425 107.625 ;
        RECT 119.840 107.580 120.160 107.640 ;
        RECT 105.135 107.440 120.160 107.580 ;
        RECT 105.135 107.395 105.425 107.440 ;
        RECT 119.840 107.380 120.160 107.440 ;
        RECT 120.775 107.580 121.065 107.625 ;
        RECT 122.140 107.580 122.460 107.640 ;
        RECT 120.775 107.440 122.460 107.580 ;
        RECT 120.775 107.395 121.065 107.440 ;
        RECT 122.140 107.380 122.460 107.440 ;
        RECT 90.400 107.100 91.550 107.240 ;
        RECT 90.400 107.040 90.720 107.100 ;
        RECT 84.140 106.900 84.430 106.945 ;
        RECT 79.820 106.760 84.430 106.900 ;
        RECT 79.820 106.700 80.140 106.760 ;
        RECT 84.140 106.715 84.430 106.760 ;
        RECT 89.955 106.715 90.245 106.945 ;
        RECT 90.860 106.700 91.180 106.960 ;
        RECT 91.410 106.945 91.550 107.100 ;
        RECT 93.710 107.100 95.230 107.240 ;
        RECT 91.335 106.715 91.625 106.945 ;
        RECT 91.780 106.900 92.100 106.960 ;
        RECT 92.255 106.900 92.545 106.945 ;
        RECT 91.780 106.760 92.545 106.900 ;
        RECT 91.780 106.700 92.100 106.760 ;
        RECT 92.255 106.715 92.545 106.760 ;
        RECT 93.160 106.700 93.480 106.960 ;
        RECT 93.710 106.945 93.850 107.100 ;
        RECT 95.090 106.960 95.230 107.100 ;
        RECT 96.840 107.100 99.370 107.240 ;
        RECT 96.840 107.040 97.160 107.100 ;
        RECT 93.635 106.715 93.925 106.945 ;
        RECT 94.080 106.700 94.400 106.960 ;
        RECT 95.000 106.900 95.320 106.960 ;
        RECT 95.935 106.900 96.225 106.945 ;
        RECT 95.000 106.760 96.225 106.900 ;
        RECT 95.000 106.700 95.320 106.760 ;
        RECT 95.935 106.715 96.225 106.760 ;
        RECT 96.380 106.900 96.700 106.960 ;
        RECT 99.230 106.945 99.370 107.100 ;
        RECT 102.375 107.055 102.665 107.285 ;
        RECT 102.820 107.240 103.140 107.300 ;
        RECT 103.295 107.240 103.585 107.285 ;
        RECT 102.820 107.100 103.585 107.240 ;
        RECT 102.820 107.040 103.140 107.100 ;
        RECT 103.295 107.055 103.585 107.100 ;
        RECT 106.040 107.240 106.360 107.300 ;
        RECT 109.260 107.240 109.580 107.300 ;
        RECT 113.860 107.240 114.180 107.300 ;
        RECT 121.695 107.240 121.985 107.285 ;
        RECT 123.520 107.240 123.840 107.300 ;
        RECT 106.040 107.100 108.570 107.240 ;
        RECT 98.235 106.900 98.525 106.945 ;
        RECT 96.380 106.760 98.525 106.900 ;
        RECT 96.380 106.700 96.700 106.760 ;
        RECT 98.235 106.715 98.525 106.760 ;
        RECT 99.155 106.715 99.445 106.945 ;
        RECT 103.735 106.825 104.025 107.055 ;
        RECT 106.040 107.040 106.360 107.100 ;
        RECT 59.120 106.360 59.440 106.620 ;
        RECT 68.780 106.560 69.100 106.620 ;
        RECT 86.735 106.560 87.025 106.605 ;
        RECT 89.480 106.560 89.800 106.620 ;
        RECT 68.780 106.420 89.800 106.560 ;
        RECT 68.780 106.360 69.100 106.420 ;
        RECT 86.735 106.375 87.025 106.420 ;
        RECT 89.480 106.360 89.800 106.420 ;
        RECT 90.415 106.560 90.705 106.605 ;
        RECT 92.700 106.560 93.020 106.620 ;
        RECT 90.415 106.420 93.020 106.560 ;
        RECT 94.170 106.560 94.310 106.700 ;
        RECT 103.830 106.620 103.970 106.825 ;
        RECT 104.215 106.715 104.505 106.945 ;
        RECT 106.975 106.900 107.265 106.945 ;
        RECT 107.880 106.900 108.200 106.960 ;
        RECT 108.430 106.945 108.570 107.100 ;
        RECT 109.260 107.100 113.630 107.240 ;
        RECT 109.260 107.040 109.580 107.100 ;
        RECT 106.975 106.760 108.200 106.900 ;
        RECT 106.975 106.715 107.265 106.760 ;
        RECT 98.695 106.560 98.985 106.605 ;
        RECT 94.170 106.420 98.985 106.560 ;
        RECT 90.415 106.375 90.705 106.420 ;
        RECT 92.700 106.360 93.020 106.420 ;
        RECT 98.695 106.375 98.985 106.420 ;
        RECT 103.740 106.360 104.060 106.620 ;
        RECT 104.290 106.560 104.430 106.715 ;
        RECT 107.880 106.700 108.200 106.760 ;
        RECT 108.355 106.715 108.645 106.945 ;
        RECT 109.735 106.900 110.025 106.945 ;
        RECT 110.180 106.900 110.500 106.960 ;
        RECT 109.735 106.760 110.500 106.900 ;
        RECT 109.735 106.715 110.025 106.760 ;
        RECT 110.180 106.700 110.500 106.760 ;
        RECT 110.655 106.900 110.945 106.945 ;
        RECT 111.100 106.900 111.420 106.960 ;
        RECT 110.655 106.760 111.420 106.900 ;
        RECT 110.655 106.715 110.945 106.760 ;
        RECT 111.100 106.700 111.420 106.760 ;
        RECT 112.020 106.700 112.340 106.960 ;
        RECT 112.480 106.900 112.800 106.960 ;
        RECT 113.490 106.945 113.630 107.100 ;
        RECT 113.860 107.100 123.840 107.240 ;
        RECT 113.860 107.040 114.180 107.100 ;
        RECT 121.695 107.055 121.985 107.100 ;
        RECT 123.520 107.040 123.840 107.100 ;
        RECT 112.955 106.900 113.245 106.945 ;
        RECT 112.480 106.760 113.245 106.900 ;
        RECT 112.480 106.700 112.800 106.760 ;
        RECT 112.955 106.715 113.245 106.760 ;
        RECT 113.415 106.715 113.705 106.945 ;
        RECT 114.320 106.700 114.640 106.960 ;
        RECT 122.155 106.900 122.445 106.945 ;
        RECT 118.090 106.760 122.445 106.900 ;
        RECT 118.090 106.620 118.230 106.760 ;
        RECT 122.155 106.715 122.445 106.760 ;
        RECT 116.160 106.560 116.480 106.620 ;
        RECT 104.290 106.420 116.480 106.560 ;
        RECT 116.160 106.360 116.480 106.420 ;
        RECT 116.620 106.360 116.940 106.620 ;
        RECT 118.000 106.360 118.320 106.620 ;
        RECT 118.920 106.560 119.240 106.620 ;
        RECT 120.300 106.560 120.620 106.620 ;
        RECT 118.920 106.420 120.620 106.560 ;
        RECT 118.920 106.360 119.240 106.420 ;
        RECT 120.300 106.360 120.620 106.420 ;
        RECT 86.275 106.220 86.565 106.265 ;
        RECT 95.475 106.220 95.765 106.265 ;
        RECT 86.275 106.080 95.765 106.220 ;
        RECT 86.275 106.035 86.565 106.080 ;
        RECT 95.475 106.035 95.765 106.080 ;
        RECT 101.440 106.220 101.760 106.280 ;
        RECT 102.375 106.220 102.665 106.265 ;
        RECT 101.440 106.080 102.665 106.220 ;
        RECT 103.830 106.220 103.970 106.360 ;
        RECT 105.580 106.220 105.900 106.280 ;
        RECT 103.830 106.080 105.900 106.220 ;
        RECT 101.440 106.020 101.760 106.080 ;
        RECT 102.375 106.035 102.665 106.080 ;
        RECT 105.580 106.020 105.900 106.080 ;
        RECT 107.880 106.020 108.200 106.280 ;
        RECT 108.800 106.220 109.120 106.280 ;
        RECT 109.275 106.220 109.565 106.265 ;
        RECT 108.800 106.080 109.565 106.220 ;
        RECT 108.800 106.020 109.120 106.080 ;
        RECT 109.275 106.035 109.565 106.080 ;
        RECT 110.640 106.220 110.960 106.280 ;
        RECT 114.320 106.220 114.640 106.280 ;
        RECT 110.640 106.080 114.640 106.220 ;
        RECT 110.640 106.020 110.960 106.080 ;
        RECT 114.320 106.020 114.640 106.080 ;
        RECT 115.240 106.020 115.560 106.280 ;
        RECT 118.475 106.220 118.765 106.265 ;
        RECT 121.220 106.220 121.540 106.280 ;
        RECT 123.075 106.220 123.365 106.265 ;
        RECT 118.475 106.080 123.365 106.220 ;
        RECT 118.475 106.035 118.765 106.080 ;
        RECT 121.220 106.020 121.540 106.080 ;
        RECT 123.075 106.035 123.365 106.080 ;
        RECT 61.895 105.880 62.185 105.925 ;
        RECT 62.815 105.880 63.105 105.925 ;
        RECT 61.895 105.740 63.105 105.880 ;
        RECT 61.895 105.695 62.185 105.740 ;
        RECT 62.815 105.695 63.105 105.740 ;
        RECT 66.020 105.880 66.340 105.940 ;
        RECT 86.720 105.880 87.040 105.940 ;
        RECT 66.020 105.740 87.040 105.880 ;
        RECT 66.020 105.680 66.340 105.740 ;
        RECT 86.720 105.680 87.040 105.740 ;
        RECT 111.100 105.880 111.420 105.940 ;
        RECT 113.400 105.880 113.720 105.940 ;
        RECT 111.100 105.740 113.720 105.880 ;
        RECT 111.100 105.680 111.420 105.740 ;
        RECT 113.400 105.680 113.720 105.740 ;
        RECT 117.540 105.880 117.860 105.940 ;
        RECT 118.920 105.880 119.240 105.940 ;
        RECT 117.540 105.740 119.240 105.880 ;
        RECT 117.540 105.680 117.860 105.740 ;
        RECT 118.920 105.680 119.240 105.740 ;
        RECT 119.840 105.680 120.160 105.940 ;
        RECT 120.300 105.880 120.620 105.940 ;
        RECT 120.775 105.880 121.065 105.925 ;
        RECT 122.600 105.880 122.920 105.940 ;
        RECT 120.300 105.740 122.920 105.880 ;
        RECT 120.300 105.680 120.620 105.740 ;
        RECT 120.775 105.695 121.065 105.740 ;
        RECT 122.600 105.680 122.920 105.740 ;
        RECT 53.990 105.060 125.290 105.540 ;
        RECT 63.720 104.860 64.040 104.920 ;
        RECT 66.035 104.860 66.325 104.905 ;
        RECT 63.720 104.720 66.325 104.860 ;
        RECT 63.720 104.660 64.040 104.720 ;
        RECT 66.035 104.675 66.325 104.720 ;
        RECT 70.175 104.860 70.465 104.905 ;
        RECT 71.540 104.860 71.860 104.920 ;
        RECT 70.175 104.720 71.860 104.860 ;
        RECT 70.175 104.675 70.465 104.720 ;
        RECT 59.120 103.980 59.440 104.240 ;
        RECT 66.110 104.180 66.250 104.675 ;
        RECT 71.540 104.660 71.860 104.720 ;
        RECT 79.360 104.660 79.680 104.920 ;
        RECT 81.200 104.860 81.520 104.920 ;
        RECT 83.500 104.860 83.820 104.920 ;
        RECT 81.200 104.720 83.820 104.860 ;
        RECT 81.200 104.660 81.520 104.720 ;
        RECT 83.500 104.660 83.820 104.720 ;
        RECT 91.780 104.860 92.100 104.920 ;
        RECT 93.175 104.860 93.465 104.905 ;
        RECT 91.780 104.720 93.465 104.860 ;
        RECT 91.780 104.660 92.100 104.720 ;
        RECT 93.175 104.675 93.465 104.720 ;
        RECT 95.475 104.860 95.765 104.905 ;
        RECT 96.380 104.860 96.700 104.920 ;
        RECT 95.475 104.720 96.700 104.860 ;
        RECT 95.475 104.675 95.765 104.720 ;
        RECT 96.380 104.660 96.700 104.720 ;
        RECT 107.435 104.860 107.725 104.905 ;
        RECT 108.340 104.860 108.660 104.920 ;
        RECT 107.435 104.720 108.660 104.860 ;
        RECT 107.435 104.675 107.725 104.720 ;
        RECT 108.340 104.660 108.660 104.720 ;
        RECT 108.800 104.860 109.120 104.920 ;
        RECT 110.640 104.860 110.960 104.920 ;
        RECT 111.115 104.860 111.405 104.905 ;
        RECT 108.800 104.720 110.410 104.860 ;
        RECT 108.800 104.660 109.120 104.720 ;
        RECT 71.095 104.335 71.385 104.565 ;
        RECT 67.875 104.180 68.165 104.225 ;
        RECT 71.170 104.180 71.310 104.335 ;
        RECT 66.110 104.040 67.630 104.180 ;
        RECT 58.200 103.840 58.520 103.900 ;
        RECT 60.055 103.840 60.345 103.885 ;
        RECT 58.200 103.700 60.345 103.840 ;
        RECT 58.200 103.640 58.520 103.700 ;
        RECT 60.055 103.655 60.345 103.700 ;
        RECT 65.575 103.655 65.865 103.885 ;
        RECT 65.650 103.500 65.790 103.655 ;
        RECT 66.480 103.640 66.800 103.900 ;
        RECT 67.490 103.885 67.630 104.040 ;
        RECT 67.875 104.040 71.310 104.180 ;
        RECT 74.315 104.180 74.605 104.225 ;
        RECT 74.760 104.180 75.080 104.240 ;
        RECT 74.315 104.040 75.080 104.180 ;
        RECT 67.875 103.995 68.165 104.040 ;
        RECT 74.315 103.995 74.605 104.040 ;
        RECT 74.760 103.980 75.080 104.040 ;
        RECT 78.440 104.180 78.760 104.240 ;
        RECT 84.880 104.180 85.200 104.240 ;
        RECT 78.440 104.040 85.200 104.180 ;
        RECT 78.440 103.980 78.760 104.040 ;
        RECT 67.415 103.655 67.705 103.885 ;
        RECT 68.795 103.655 69.085 103.885 ;
        RECT 69.255 103.840 69.545 103.885 ;
        RECT 70.620 103.840 70.940 103.900 ;
        RECT 69.255 103.700 70.940 103.840 ;
        RECT 69.255 103.655 69.545 103.700 ;
        RECT 67.860 103.500 68.180 103.560 ;
        RECT 65.650 103.360 68.180 103.500 ;
        RECT 68.870 103.500 69.010 103.655 ;
        RECT 70.620 103.640 70.940 103.700 ;
        RECT 71.540 103.840 71.860 103.900 ;
        RECT 75.235 103.840 75.525 103.885 ;
        RECT 71.540 103.700 75.525 103.840 ;
        RECT 71.540 103.640 71.860 103.700 ;
        RECT 75.235 103.655 75.525 103.700 ;
        RECT 76.140 103.640 76.460 103.900 ;
        RECT 80.830 103.885 80.970 104.040 ;
        RECT 84.880 103.980 85.200 104.040 ;
        RECT 94.540 103.980 94.860 104.240 ;
        RECT 101.900 104.180 102.220 104.240 ;
        RECT 95.550 104.040 102.220 104.180 ;
        RECT 80.295 103.655 80.585 103.885 ;
        RECT 80.755 103.655 81.045 103.885 ;
        RECT 74.300 103.500 74.620 103.560 ;
        RECT 68.870 103.360 74.620 103.500 ;
        RECT 80.370 103.500 80.510 103.655 ;
        RECT 81.660 103.640 81.980 103.900 ;
        RECT 82.135 103.840 82.425 103.885 ;
        RECT 87.640 103.840 87.960 103.900 ;
        RECT 82.135 103.700 87.960 103.840 ;
        RECT 82.135 103.655 82.425 103.700 ;
        RECT 87.640 103.640 87.960 103.700 ;
        RECT 89.940 103.840 90.260 103.900 ;
        RECT 95.550 103.840 95.690 104.040 ;
        RECT 101.900 103.980 102.220 104.040 ;
        RECT 89.940 103.700 95.690 103.840 ;
        RECT 89.940 103.640 90.260 103.700 ;
        RECT 95.920 103.640 96.240 103.900 ;
        RECT 110.270 103.885 110.410 104.720 ;
        RECT 110.640 104.720 111.405 104.860 ;
        RECT 110.640 104.660 110.960 104.720 ;
        RECT 111.115 104.675 111.405 104.720 ;
        RECT 112.020 104.860 112.340 104.920 ;
        RECT 113.400 104.860 113.720 104.920 ;
        RECT 112.020 104.720 113.720 104.860 ;
        RECT 112.020 104.660 112.340 104.720 ;
        RECT 113.400 104.660 113.720 104.720 ;
        RECT 111.560 104.520 111.880 104.580 ;
        RECT 115.255 104.520 115.545 104.565 ;
        RECT 111.560 104.380 115.545 104.520 ;
        RECT 111.560 104.320 111.880 104.380 ;
        RECT 115.255 104.335 115.545 104.380 ;
        RECT 112.480 104.180 112.800 104.240 ;
        RECT 113.875 104.180 114.165 104.225 ;
        RECT 112.480 104.040 114.165 104.180 ;
        RECT 112.480 103.980 112.800 104.040 ;
        RECT 113.875 103.995 114.165 104.040 ;
        RECT 116.160 103.980 116.480 104.240 ;
        RECT 117.170 104.040 121.450 104.180 ;
        RECT 110.195 103.655 110.485 103.885 ;
        RECT 110.640 103.840 110.960 103.900 ;
        RECT 111.115 103.840 111.405 103.885 ;
        RECT 110.640 103.700 111.405 103.840 ;
        RECT 110.640 103.640 110.960 103.700 ;
        RECT 111.115 103.655 111.405 103.700 ;
        RECT 112.020 103.640 112.340 103.900 ;
        RECT 90.860 103.500 91.180 103.560 ;
        RECT 80.370 103.360 99.830 103.500 ;
        RECT 67.860 103.300 68.180 103.360 ;
        RECT 74.300 103.300 74.620 103.360 ;
        RECT 90.860 103.300 91.180 103.360 ;
        RECT 99.690 103.220 99.830 103.360 ;
        RECT 107.880 103.300 108.200 103.560 ;
        RECT 112.570 103.500 112.710 103.980 ;
        RECT 113.415 103.840 113.705 103.885 ;
        RECT 114.780 103.840 115.100 103.900 ;
        RECT 117.170 103.885 117.310 104.040 ;
        RECT 121.310 103.900 121.450 104.040 ;
        RECT 113.415 103.700 115.100 103.840 ;
        RECT 113.415 103.655 113.705 103.700 ;
        RECT 114.780 103.640 115.100 103.700 ;
        RECT 117.095 103.655 117.385 103.885 ;
        RECT 118.015 103.840 118.305 103.885 ;
        RECT 118.460 103.840 118.780 103.900 ;
        RECT 118.015 103.700 118.780 103.840 ;
        RECT 118.015 103.655 118.305 103.700 ;
        RECT 118.460 103.640 118.780 103.700 ;
        RECT 118.935 103.840 119.225 103.885 ;
        RECT 120.760 103.840 121.080 103.900 ;
        RECT 118.935 103.700 121.080 103.840 ;
        RECT 118.935 103.655 119.225 103.700 ;
        RECT 120.760 103.640 121.080 103.700 ;
        RECT 121.220 103.640 121.540 103.900 ;
        RECT 122.155 103.840 122.445 103.885 ;
        RECT 122.600 103.840 122.920 103.900 ;
        RECT 122.155 103.700 122.920 103.840 ;
        RECT 122.155 103.655 122.445 103.700 ;
        RECT 122.600 103.640 122.920 103.700 ;
        RECT 123.075 103.655 123.365 103.885 ;
        RECT 109.810 103.360 112.710 103.500 ;
        RECT 116.620 103.500 116.940 103.560 ;
        RECT 123.150 103.500 123.290 103.655 ;
        RECT 116.620 103.360 123.290 103.500 ;
        RECT 59.580 102.960 59.900 103.220 ;
        RECT 61.895 103.160 62.185 103.205 ;
        RECT 64.180 103.160 64.500 103.220 ;
        RECT 61.895 103.020 64.500 103.160 ;
        RECT 61.895 102.975 62.185 103.020 ;
        RECT 64.180 102.960 64.500 103.020 ;
        RECT 72.000 103.160 72.320 103.220 ;
        RECT 72.935 103.160 73.225 103.205 ;
        RECT 72.000 103.020 73.225 103.160 ;
        RECT 72.000 102.960 72.320 103.020 ;
        RECT 72.935 102.975 73.225 103.020 ;
        RECT 73.395 103.160 73.685 103.205 ;
        RECT 74.760 103.160 75.080 103.220 ;
        RECT 75.235 103.160 75.525 103.205 ;
        RECT 73.395 103.020 75.525 103.160 ;
        RECT 73.395 102.975 73.685 103.020 ;
        RECT 74.760 102.960 75.080 103.020 ;
        RECT 75.235 102.975 75.525 103.020 ;
        RECT 85.800 103.160 86.120 103.220 ;
        RECT 88.100 103.160 88.420 103.220 ;
        RECT 89.480 103.160 89.800 103.220 ;
        RECT 99.140 103.160 99.460 103.220 ;
        RECT 85.800 103.020 99.460 103.160 ;
        RECT 85.800 102.960 86.120 103.020 ;
        RECT 88.100 102.960 88.420 103.020 ;
        RECT 89.480 102.960 89.800 103.020 ;
        RECT 99.140 102.960 99.460 103.020 ;
        RECT 99.600 103.160 99.920 103.220 ;
        RECT 109.810 103.205 109.950 103.360 ;
        RECT 116.620 103.300 116.940 103.360 ;
        RECT 108.895 103.160 109.185 103.205 ;
        RECT 99.600 103.020 109.185 103.160 ;
        RECT 99.600 102.960 99.920 103.020 ;
        RECT 108.895 102.975 109.185 103.020 ;
        RECT 109.735 102.975 110.025 103.205 ;
        RECT 112.940 102.960 113.260 103.220 ;
        RECT 117.080 103.160 117.400 103.220 ;
        RECT 120.775 103.160 121.065 103.205 ;
        RECT 117.080 103.020 121.065 103.160 ;
        RECT 117.080 102.960 117.400 103.020 ;
        RECT 120.775 102.975 121.065 103.020 ;
        RECT 53.990 102.340 125.290 102.820 ;
        RECT 58.660 102.140 58.980 102.200 ;
        RECT 60.500 102.140 60.820 102.200 ;
        RECT 58.660 102.000 70.390 102.140 ;
        RECT 58.660 101.940 58.980 102.000 ;
        RECT 60.500 101.940 60.820 102.000 ;
        RECT 66.480 101.800 66.800 101.860 ;
        RECT 70.250 101.800 70.390 102.000 ;
        RECT 70.620 101.940 70.940 102.200 ;
        RECT 72.935 102.140 73.225 102.185 ;
        RECT 74.760 102.140 75.080 102.200 ;
        RECT 72.935 102.000 75.080 102.140 ;
        RECT 72.935 101.955 73.225 102.000 ;
        RECT 74.760 101.940 75.080 102.000 ;
        RECT 80.295 102.140 80.585 102.185 ;
        RECT 81.660 102.140 81.980 102.200 ;
        RECT 80.295 102.000 81.980 102.140 ;
        RECT 80.295 101.955 80.585 102.000 ;
        RECT 81.660 101.940 81.980 102.000 ;
        RECT 82.120 102.140 82.440 102.200 ;
        RECT 82.120 102.000 86.490 102.140 ;
        RECT 82.120 101.940 82.440 102.000 ;
        RECT 75.680 101.800 76.000 101.860 ;
        RECT 76.615 101.800 76.905 101.845 ;
        RECT 83.500 101.800 83.820 101.860 ;
        RECT 66.480 101.660 69.010 101.800 ;
        RECT 70.250 101.660 75.450 101.800 ;
        RECT 66.480 101.600 66.800 101.660 ;
        RECT 56.835 101.275 57.125 101.505 ;
        RECT 56.910 101.120 57.050 101.275 ;
        RECT 57.740 101.260 58.060 101.520 ;
        RECT 67.030 101.505 67.170 101.660 ;
        RECT 60.055 101.460 60.345 101.505 ;
        RECT 66.955 101.460 67.245 101.505 ;
        RECT 60.055 101.320 67.245 101.460 ;
        RECT 60.055 101.275 60.345 101.320 ;
        RECT 66.955 101.275 67.245 101.320 ;
        RECT 67.400 101.260 67.720 101.520 ;
        RECT 67.860 101.460 68.180 101.520 ;
        RECT 68.870 101.505 69.010 101.660 ;
        RECT 68.335 101.460 68.625 101.505 ;
        RECT 67.860 101.320 68.625 101.460 ;
        RECT 67.860 101.260 68.180 101.320 ;
        RECT 68.335 101.275 68.625 101.320 ;
        RECT 68.795 101.275 69.085 101.505 ;
        RECT 72.000 101.460 72.320 101.520 ;
        RECT 72.475 101.460 72.765 101.505 ;
        RECT 74.300 101.460 74.620 101.520 ;
        RECT 72.000 101.320 74.620 101.460 ;
        RECT 75.310 101.460 75.450 101.660 ;
        RECT 75.680 101.660 82.810 101.800 ;
        RECT 75.680 101.600 76.000 101.660 ;
        RECT 76.615 101.615 76.905 101.660 ;
        RECT 77.535 101.460 77.825 101.505 ;
        RECT 78.440 101.460 78.760 101.520 ;
        RECT 75.310 101.320 77.290 101.460 ;
        RECT 68.410 101.120 68.550 101.275 ;
        RECT 72.000 101.260 72.320 101.320 ;
        RECT 72.475 101.275 72.765 101.320 ;
        RECT 74.300 101.260 74.620 101.320 ;
        RECT 73.855 101.120 74.145 101.165 ;
        RECT 74.760 101.120 75.080 101.180 ;
        RECT 76.140 101.120 76.460 101.180 ;
        RECT 56.910 100.980 59.350 101.120 ;
        RECT 68.410 100.980 70.390 101.120 ;
        RECT 55.900 100.580 56.220 100.840 ;
        RECT 59.210 100.825 59.350 100.980 ;
        RECT 59.135 100.595 59.425 100.825 ;
        RECT 70.250 100.780 70.390 100.980 ;
        RECT 73.855 100.980 76.460 101.120 ;
        RECT 77.150 101.120 77.290 101.320 ;
        RECT 77.535 101.320 78.760 101.460 ;
        RECT 77.535 101.275 77.825 101.320 ;
        RECT 78.440 101.260 78.760 101.320 ;
        RECT 78.900 101.460 79.220 101.520 ;
        RECT 82.670 101.505 82.810 101.660 ;
        RECT 83.500 101.660 84.650 101.800 ;
        RECT 83.500 101.600 83.820 101.660 ;
        RECT 81.215 101.460 81.505 101.505 ;
        RECT 78.900 101.320 81.505 101.460 ;
        RECT 78.900 101.260 79.220 101.320 ;
        RECT 81.215 101.275 81.505 101.320 ;
        RECT 82.595 101.275 82.885 101.505 ;
        RECT 83.040 101.260 83.360 101.520 ;
        RECT 83.960 101.460 84.280 101.520 ;
        RECT 84.510 101.505 84.650 101.660 ;
        RECT 85.800 101.600 86.120 101.860 ;
        RECT 86.350 101.845 86.490 102.000 ;
        RECT 87.640 101.940 87.960 102.200 ;
        RECT 88.650 102.000 90.630 102.140 ;
        RECT 86.275 101.800 86.565 101.845 ;
        RECT 88.650 101.800 88.790 102.000 ;
        RECT 86.275 101.660 88.790 101.800 ;
        RECT 86.275 101.615 86.565 101.660 ;
        RECT 89.020 101.600 89.340 101.860 ;
        RECT 89.480 101.600 89.800 101.860 ;
        RECT 90.490 101.800 90.630 102.000 ;
        RECT 90.860 101.940 91.180 102.200 ;
        RECT 92.240 102.140 92.560 102.200 ;
        RECT 99.140 102.140 99.460 102.200 ;
        RECT 101.915 102.140 102.205 102.185 ;
        RECT 92.240 102.000 98.910 102.140 ;
        RECT 92.240 101.940 92.560 102.000 ;
        RECT 96.380 101.800 96.700 101.860 ;
        RECT 98.770 101.800 98.910 102.000 ;
        RECT 99.140 102.000 102.205 102.140 ;
        RECT 99.140 101.940 99.460 102.000 ;
        RECT 101.915 101.955 102.205 102.000 ;
        RECT 103.740 102.140 104.060 102.200 ;
        RECT 106.055 102.140 106.345 102.185 ;
        RECT 103.740 102.000 106.345 102.140 ;
        RECT 103.740 101.940 104.060 102.000 ;
        RECT 106.055 101.955 106.345 102.000 ;
        RECT 111.100 101.940 111.420 102.200 ;
        RECT 113.400 101.940 113.720 102.200 ;
        RECT 121.220 101.940 121.540 102.200 ;
        RECT 100.520 101.800 100.840 101.860 ;
        RECT 107.880 101.800 108.200 101.860 ;
        RECT 109.260 101.800 109.580 101.860 ;
        RECT 90.490 101.660 96.700 101.800 ;
        RECT 96.380 101.600 96.700 101.660 ;
        RECT 96.930 101.660 98.450 101.800 ;
        RECT 98.770 101.660 100.290 101.800 ;
        RECT 83.590 101.320 84.280 101.460 ;
        RECT 81.660 101.120 81.980 101.180 ;
        RECT 82.135 101.120 82.425 101.165 ;
        RECT 83.590 101.120 83.730 101.320 ;
        RECT 83.960 101.260 84.280 101.320 ;
        RECT 84.435 101.275 84.725 101.505 ;
        RECT 85.125 101.275 85.415 101.505 ;
        RECT 86.735 101.460 87.025 101.505 ;
        RECT 88.115 101.460 88.405 101.505 ;
        RECT 86.735 101.320 88.405 101.460 ;
        RECT 86.735 101.275 87.025 101.320 ;
        RECT 88.115 101.275 88.405 101.320 ;
        RECT 89.955 101.460 90.245 101.505 ;
        RECT 92.240 101.460 92.560 101.520 ;
        RECT 96.930 101.505 97.070 101.660 ;
        RECT 89.955 101.320 92.560 101.460 ;
        RECT 89.955 101.275 90.245 101.320 ;
        RECT 85.200 101.120 85.340 101.275 ;
        RECT 77.150 100.980 82.425 101.120 ;
        RECT 73.855 100.935 74.145 100.980 ;
        RECT 74.760 100.920 75.080 100.980 ;
        RECT 76.140 100.920 76.460 100.980 ;
        RECT 81.660 100.920 81.980 100.980 ;
        RECT 82.135 100.935 82.425 100.980 ;
        RECT 83.130 100.980 83.730 101.120 ;
        RECT 84.215 100.980 85.340 101.120 ;
        RECT 85.800 101.120 86.120 101.180 ;
        RECT 86.810 101.120 86.950 101.275 ;
        RECT 85.800 100.980 86.950 101.120 ;
        RECT 88.190 101.120 88.330 101.275 ;
        RECT 92.240 101.260 92.560 101.320 ;
        RECT 96.855 101.275 97.145 101.505 ;
        RECT 97.775 101.275 98.065 101.505 ;
        RECT 94.080 101.120 94.400 101.180 ;
        RECT 96.930 101.120 97.070 101.275 ;
        RECT 88.190 100.980 97.070 101.120 ;
        RECT 76.600 100.780 76.920 100.840 ;
        RECT 70.250 100.640 76.920 100.780 ;
        RECT 76.600 100.580 76.920 100.640 ;
        RECT 78.455 100.780 78.745 100.825 ;
        RECT 79.360 100.780 79.680 100.840 ;
        RECT 78.455 100.640 79.680 100.780 ;
        RECT 78.455 100.595 78.745 100.640 ;
        RECT 79.360 100.580 79.680 100.640 ;
        RECT 58.200 100.240 58.520 100.500 ;
        RECT 69.715 100.440 70.005 100.485 ;
        RECT 83.130 100.440 83.270 100.980 ;
        RECT 84.215 100.840 84.355 100.980 ;
        RECT 85.800 100.920 86.120 100.980 ;
        RECT 94.080 100.920 94.400 100.980 ;
        RECT 83.960 100.640 84.355 100.840 ;
        RECT 89.020 100.780 89.340 100.840 ;
        RECT 91.320 100.780 91.640 100.840 ;
        RECT 94.540 100.780 94.860 100.840 ;
        RECT 97.850 100.780 97.990 101.275 ;
        RECT 98.310 101.180 98.450 101.660 ;
        RECT 99.140 101.260 99.460 101.520 ;
        RECT 100.150 101.505 100.290 101.660 ;
        RECT 100.520 101.660 103.050 101.800 ;
        RECT 100.520 101.600 100.840 101.660 ;
        RECT 102.910 101.505 103.050 101.660 ;
        RECT 107.880 101.660 109.580 101.800 ;
        RECT 107.880 101.600 108.200 101.660 ;
        RECT 100.075 101.275 100.365 101.505 ;
        RECT 101.455 101.460 101.745 101.505 ;
        RECT 100.610 101.320 101.745 101.460 ;
        RECT 98.220 101.120 98.540 101.180 ;
        RECT 100.610 101.120 100.750 101.320 ;
        RECT 101.455 101.275 101.745 101.320 ;
        RECT 102.835 101.275 103.125 101.505 ;
        RECT 106.500 101.460 106.820 101.520 ;
        RECT 106.975 101.460 107.265 101.505 ;
        RECT 106.500 101.320 107.265 101.460 ;
        RECT 106.500 101.260 106.820 101.320 ;
        RECT 106.975 101.275 107.265 101.320 ;
        RECT 107.435 101.460 107.725 101.505 ;
        RECT 108.340 101.460 108.660 101.520 ;
        RECT 108.890 101.505 109.030 101.660 ;
        RECT 109.260 101.600 109.580 101.660 ;
        RECT 107.435 101.320 108.660 101.460 ;
        RECT 107.435 101.275 107.725 101.320 ;
        RECT 108.340 101.260 108.660 101.320 ;
        RECT 108.815 101.275 109.105 101.505 ;
        RECT 110.425 101.460 110.715 101.675 ;
        RECT 111.560 101.600 111.880 101.860 ;
        RECT 112.480 101.845 112.800 101.860 ;
        RECT 112.480 101.615 112.865 101.845 ;
        RECT 114.795 101.800 115.085 101.845 ;
        RECT 119.380 101.800 119.700 101.860 ;
        RECT 114.795 101.660 119.700 101.800 ;
        RECT 114.795 101.615 115.085 101.660 ;
        RECT 112.480 101.600 112.800 101.615 ;
        RECT 119.380 101.600 119.700 101.660 ;
        RECT 109.350 101.445 110.715 101.460 ;
        RECT 109.350 101.320 110.640 101.445 ;
        RECT 98.220 100.980 100.750 101.120 ;
        RECT 100.980 101.120 101.300 101.180 ;
        RECT 103.755 101.120 104.045 101.165 ;
        RECT 109.350 101.120 109.490 101.320 ;
        RECT 100.980 100.980 109.490 101.120 ;
        RECT 98.220 100.920 98.540 100.980 ;
        RECT 100.980 100.920 101.300 100.980 ;
        RECT 103.755 100.935 104.045 100.980 ;
        RECT 89.020 100.640 97.990 100.780 ;
        RECT 98.695 100.780 98.985 100.825 ;
        RECT 107.880 100.780 108.200 100.840 ;
        RECT 108.355 100.780 108.645 100.825 ;
        RECT 110.640 100.780 110.960 100.840 ;
        RECT 98.695 100.640 112.710 100.780 ;
        RECT 83.960 100.580 84.280 100.640 ;
        RECT 89.020 100.580 89.340 100.640 ;
        RECT 91.320 100.580 91.640 100.640 ;
        RECT 94.540 100.580 94.860 100.640 ;
        RECT 98.695 100.595 98.985 100.640 ;
        RECT 107.880 100.580 108.200 100.640 ;
        RECT 108.355 100.595 108.645 100.640 ;
        RECT 110.640 100.580 110.960 100.640 ;
        RECT 69.715 100.300 83.270 100.440 ;
        RECT 83.500 100.440 83.820 100.500 ;
        RECT 85.340 100.440 85.660 100.500 ;
        RECT 83.500 100.300 85.660 100.440 ;
        RECT 69.715 100.255 70.005 100.300 ;
        RECT 83.500 100.240 83.820 100.300 ;
        RECT 85.340 100.240 85.660 100.300 ;
        RECT 86.720 100.440 87.040 100.500 ;
        RECT 89.940 100.440 90.260 100.500 ;
        RECT 86.720 100.300 90.260 100.440 ;
        RECT 86.720 100.240 87.040 100.300 ;
        RECT 89.940 100.240 90.260 100.300 ;
        RECT 96.380 100.440 96.700 100.500 ;
        RECT 104.660 100.440 104.980 100.500 ;
        RECT 107.420 100.440 107.740 100.500 ;
        RECT 96.380 100.300 107.740 100.440 ;
        RECT 96.380 100.240 96.700 100.300 ;
        RECT 104.660 100.240 104.980 100.300 ;
        RECT 107.420 100.240 107.740 100.300 ;
        RECT 108.800 100.440 109.120 100.500 ;
        RECT 112.570 100.485 112.710 100.640 ;
        RECT 110.195 100.440 110.485 100.485 ;
        RECT 108.800 100.300 110.485 100.440 ;
        RECT 108.800 100.240 109.120 100.300 ;
        RECT 110.195 100.255 110.485 100.300 ;
        RECT 112.495 100.255 112.785 100.485 ;
        RECT 53.990 99.620 125.290 100.100 ;
        RECT 57.280 99.220 57.600 99.480 ;
        RECT 59.580 99.420 59.900 99.480 ;
        RECT 61.895 99.420 62.185 99.465 ;
        RECT 59.580 99.280 62.185 99.420 ;
        RECT 59.580 99.220 59.900 99.280 ;
        RECT 61.895 99.235 62.185 99.280 ;
        RECT 62.340 99.220 62.660 99.480 ;
        RECT 65.100 99.420 65.420 99.480 ;
        RECT 67.860 99.420 68.180 99.480 ;
        RECT 65.100 99.280 68.180 99.420 ;
        RECT 65.100 99.220 65.420 99.280 ;
        RECT 67.860 99.220 68.180 99.280 ;
        RECT 75.680 99.220 76.000 99.480 ;
        RECT 81.660 99.420 81.980 99.480 ;
        RECT 85.355 99.420 85.645 99.465 ;
        RECT 81.660 99.280 91.090 99.420 ;
        RECT 81.660 99.220 81.980 99.280 ;
        RECT 85.355 99.235 85.645 99.280 ;
        RECT 58.200 99.080 58.520 99.140 ;
        RECT 60.055 99.080 60.345 99.125 ;
        RECT 63.260 99.080 63.580 99.140 ;
        RECT 56.450 98.940 63.580 99.080 ;
        RECT 56.450 98.445 56.590 98.940 ;
        RECT 58.200 98.880 58.520 98.940 ;
        RECT 60.055 98.895 60.345 98.940 ;
        RECT 63.260 98.880 63.580 98.940 ;
        RECT 72.460 99.080 72.780 99.140 ;
        RECT 74.300 99.080 74.620 99.140 ;
        RECT 83.960 99.080 84.280 99.140 ;
        RECT 72.460 98.940 74.070 99.080 ;
        RECT 72.460 98.880 72.780 98.940 ;
        RECT 57.755 98.555 58.045 98.785 ;
        RECT 60.500 98.740 60.820 98.800 ;
        RECT 73.930 98.785 74.070 98.940 ;
        RECT 74.300 98.940 84.280 99.080 ;
        RECT 74.300 98.880 74.620 98.940 ;
        RECT 83.960 98.880 84.280 98.940 ;
        RECT 89.480 98.880 89.800 99.140 ;
        RECT 90.415 99.080 90.705 99.125 ;
        RECT 90.030 98.940 90.705 99.080 ;
        RECT 90.950 99.080 91.090 99.280 ;
        RECT 101.440 99.220 101.760 99.480 ;
        RECT 102.820 99.420 103.140 99.480 ;
        RECT 103.295 99.420 103.585 99.465 ;
        RECT 102.820 99.280 103.585 99.420 ;
        RECT 102.820 99.220 103.140 99.280 ;
        RECT 103.295 99.235 103.585 99.280 ;
        RECT 107.880 99.220 108.200 99.480 ;
        RECT 108.815 99.420 109.105 99.465 ;
        RECT 109.720 99.420 110.040 99.480 ;
        RECT 108.815 99.280 110.040 99.420 ;
        RECT 108.815 99.235 109.105 99.280 ;
        RECT 109.720 99.220 110.040 99.280 ;
        RECT 110.195 99.420 110.485 99.465 ;
        RECT 114.780 99.420 115.100 99.480 ;
        RECT 110.195 99.280 115.100 99.420 ;
        RECT 110.195 99.235 110.485 99.280 ;
        RECT 114.780 99.220 115.100 99.280 ;
        RECT 116.160 99.220 116.480 99.480 ;
        RECT 100.075 99.080 100.365 99.125 ;
        RECT 106.500 99.080 106.820 99.140 ;
        RECT 90.950 98.940 95.690 99.080 ;
        RECT 61.435 98.740 61.725 98.785 ;
        RECT 73.855 98.740 74.145 98.785 ;
        RECT 75.680 98.740 76.000 98.800 ;
        RECT 90.030 98.740 90.170 98.940 ;
        RECT 90.415 98.895 90.705 98.940 ;
        RECT 91.320 98.740 91.640 98.800 ;
        RECT 95.015 98.740 95.305 98.785 ;
        RECT 60.500 98.600 61.725 98.740 ;
        RECT 56.375 98.215 56.665 98.445 ;
        RECT 56.835 98.215 57.125 98.445 ;
        RECT 57.830 98.400 57.970 98.555 ;
        RECT 60.500 98.540 60.820 98.600 ;
        RECT 61.435 98.555 61.725 98.600 ;
        RECT 62.430 98.600 73.610 98.740 ;
        RECT 62.430 98.400 62.570 98.600 ;
        RECT 57.830 98.260 62.570 98.400 ;
        RECT 62.815 98.400 63.105 98.445 ;
        RECT 63.260 98.400 63.580 98.460 ;
        RECT 62.815 98.260 63.580 98.400 ;
        RECT 62.815 98.215 63.105 98.260 ;
        RECT 56.910 98.060 57.050 98.215 ;
        RECT 63.260 98.200 63.580 98.260 ;
        RECT 68.795 98.400 69.085 98.445 ;
        RECT 72.460 98.400 72.780 98.460 ;
        RECT 68.795 98.260 72.780 98.400 ;
        RECT 73.470 98.400 73.610 98.600 ;
        RECT 73.855 98.600 76.000 98.740 ;
        RECT 73.855 98.555 74.145 98.600 ;
        RECT 75.680 98.540 76.000 98.600 ;
        RECT 84.970 98.600 89.250 98.740 ;
        RECT 90.030 98.600 91.640 98.740 ;
        RECT 84.970 98.460 85.110 98.600 ;
        RECT 74.775 98.400 75.065 98.445 ;
        RECT 78.900 98.400 79.220 98.460 ;
        RECT 73.470 98.260 79.220 98.400 ;
        RECT 68.795 98.215 69.085 98.260 ;
        RECT 72.460 98.200 72.780 98.260 ;
        RECT 74.775 98.215 75.065 98.260 ;
        RECT 78.900 98.200 79.220 98.260 ;
        RECT 84.435 98.400 84.725 98.445 ;
        RECT 84.880 98.400 85.200 98.460 ;
        RECT 84.435 98.260 85.200 98.400 ;
        RECT 84.435 98.215 84.725 98.260 ;
        RECT 84.880 98.200 85.200 98.260 ;
        RECT 85.815 98.400 86.105 98.445 ;
        RECT 86.720 98.400 87.040 98.460 ;
        RECT 85.815 98.260 87.040 98.400 ;
        RECT 85.815 98.215 86.105 98.260 ;
        RECT 86.720 98.200 87.040 98.260 ;
        RECT 88.100 98.200 88.420 98.460 ;
        RECT 89.110 98.400 89.250 98.600 ;
        RECT 91.320 98.540 91.640 98.600 ;
        RECT 93.250 98.600 95.305 98.740 ;
        RECT 93.250 98.400 93.390 98.600 ;
        RECT 95.015 98.555 95.305 98.600 ;
        RECT 89.110 98.260 93.390 98.400 ;
        RECT 93.635 98.400 93.925 98.445 ;
        RECT 94.080 98.400 94.400 98.460 ;
        RECT 93.635 98.260 94.400 98.400 ;
        RECT 93.635 98.215 93.925 98.260 ;
        RECT 94.080 98.200 94.400 98.260 ;
        RECT 58.215 98.060 58.505 98.105 ;
        RECT 62.340 98.060 62.660 98.120 ;
        RECT 56.910 97.920 62.660 98.060 ;
        RECT 78.990 98.060 79.130 98.200 ;
        RECT 95.090 98.060 95.230 98.555 ;
        RECT 95.550 98.400 95.690 98.940 ;
        RECT 100.075 98.940 106.820 99.080 ;
        RECT 100.075 98.895 100.365 98.940 ;
        RECT 106.500 98.880 106.820 98.940 ;
        RECT 107.050 98.940 116.850 99.080 ;
        RECT 99.600 98.740 99.920 98.800 ;
        RECT 101.455 98.740 101.745 98.785 ;
        RECT 99.600 98.600 101.745 98.740 ;
        RECT 99.600 98.540 99.920 98.600 ;
        RECT 101.455 98.555 101.745 98.600 ;
        RECT 101.900 98.740 102.220 98.800 ;
        RECT 107.050 98.740 107.190 98.940 ;
        RECT 116.710 98.785 116.850 98.940 ;
        RECT 101.900 98.600 107.190 98.740 ;
        RECT 116.635 98.740 116.925 98.785 ;
        RECT 116.635 98.600 122.830 98.740 ;
        RECT 101.900 98.540 102.220 98.600 ;
        RECT 116.635 98.555 116.925 98.600 ;
        RECT 122.690 98.460 122.830 98.600 ;
        RECT 95.935 98.400 96.225 98.445 ;
        RECT 97.760 98.400 98.080 98.460 ;
        RECT 95.550 98.260 98.080 98.400 ;
        RECT 95.935 98.215 96.225 98.260 ;
        RECT 97.760 98.200 98.080 98.260 ;
        RECT 98.220 98.400 98.540 98.460 ;
        RECT 98.695 98.400 98.985 98.445 ;
        RECT 98.220 98.260 98.985 98.400 ;
        RECT 98.220 98.200 98.540 98.260 ;
        RECT 98.695 98.215 98.985 98.260 ;
        RECT 99.140 98.200 99.460 98.460 ;
        RECT 100.980 98.200 101.300 98.460 ;
        RECT 102.375 98.215 102.665 98.445 ;
        RECT 106.040 98.400 106.360 98.460 ;
        RECT 109.260 98.400 109.580 98.460 ;
        RECT 106.040 98.260 109.580 98.400 ;
        RECT 100.075 98.060 100.365 98.105 ;
        RECT 100.520 98.060 100.840 98.120 ;
        RECT 102.450 98.060 102.590 98.215 ;
        RECT 106.040 98.200 106.360 98.260 ;
        RECT 109.260 98.200 109.580 98.260 ;
        RECT 110.195 98.400 110.485 98.445 ;
        RECT 112.480 98.400 112.800 98.460 ;
        RECT 110.195 98.260 112.800 98.400 ;
        RECT 110.195 98.215 110.485 98.260 ;
        RECT 106.975 98.060 107.265 98.105 ;
        RECT 110.270 98.060 110.410 98.215 ;
        RECT 112.480 98.200 112.800 98.260 ;
        RECT 115.255 98.400 115.545 98.445 ;
        RECT 117.080 98.400 117.400 98.460 ;
        RECT 115.255 98.260 117.400 98.400 ;
        RECT 115.255 98.215 115.545 98.260 ;
        RECT 117.080 98.200 117.400 98.260 ;
        RECT 119.395 98.215 119.685 98.445 ;
        RECT 78.990 97.920 90.170 98.060 ;
        RECT 95.090 97.920 100.840 98.060 ;
        RECT 58.215 97.875 58.505 97.920 ;
        RECT 62.340 97.860 62.660 97.920 ;
        RECT 60.515 97.720 60.805 97.765 ;
        RECT 66.940 97.720 67.260 97.780 ;
        RECT 60.515 97.580 67.260 97.720 ;
        RECT 60.515 97.535 60.805 97.580 ;
        RECT 66.940 97.520 67.260 97.580 ;
        RECT 83.500 97.520 83.820 97.780 ;
        RECT 90.030 97.720 90.170 97.920 ;
        RECT 100.075 97.875 100.365 97.920 ;
        RECT 100.520 97.860 100.840 97.920 ;
        RECT 101.070 97.920 107.265 98.060 ;
        RECT 101.070 97.780 101.210 97.920 ;
        RECT 106.975 97.875 107.265 97.920 ;
        RECT 108.430 97.920 110.410 98.060 ;
        RECT 117.555 98.060 117.845 98.105 ;
        RECT 118.000 98.060 118.320 98.120 ;
        RECT 117.555 97.920 118.320 98.060 ;
        RECT 94.095 97.720 94.385 97.765 ;
        RECT 90.030 97.580 94.385 97.720 ;
        RECT 94.095 97.535 94.385 97.580 ;
        RECT 94.540 97.520 94.860 97.780 ;
        RECT 95.000 97.520 95.320 97.780 ;
        RECT 100.980 97.520 101.300 97.780 ;
        RECT 106.500 97.720 106.820 97.780 ;
        RECT 107.975 97.720 108.265 97.765 ;
        RECT 108.430 97.720 108.570 97.920 ;
        RECT 117.555 97.875 117.845 97.920 ;
        RECT 118.000 97.860 118.320 97.920 ;
        RECT 106.500 97.580 108.570 97.720 ;
        RECT 117.080 97.720 117.400 97.780 ;
        RECT 119.470 97.720 119.610 98.215 ;
        RECT 122.140 98.200 122.460 98.460 ;
        RECT 122.600 98.400 122.920 98.460 ;
        RECT 123.075 98.400 123.365 98.445 ;
        RECT 122.600 98.260 123.365 98.400 ;
        RECT 122.600 98.200 122.920 98.260 ;
        RECT 123.075 98.215 123.365 98.260 ;
        RECT 117.080 97.580 119.610 97.720 ;
        RECT 120.315 97.720 120.605 97.765 ;
        RECT 120.760 97.720 121.080 97.780 ;
        RECT 120.315 97.580 121.080 97.720 ;
        RECT 106.500 97.520 106.820 97.580 ;
        RECT 107.975 97.535 108.265 97.580 ;
        RECT 117.080 97.520 117.400 97.580 ;
        RECT 120.315 97.535 120.605 97.580 ;
        RECT 120.760 97.520 121.080 97.580 ;
        RECT 122.615 97.720 122.905 97.765 ;
        RECT 123.520 97.720 123.840 97.780 ;
        RECT 122.615 97.580 123.840 97.720 ;
        RECT 122.615 97.535 122.905 97.580 ;
        RECT 123.520 97.520 123.840 97.580 ;
        RECT 53.990 96.900 125.290 97.380 ;
        RECT 61.420 96.700 61.740 96.760 ;
        RECT 62.355 96.700 62.645 96.745 ;
        RECT 61.420 96.560 62.645 96.700 ;
        RECT 61.420 96.500 61.740 96.560 ;
        RECT 62.355 96.515 62.645 96.560 ;
        RECT 64.195 96.700 64.485 96.745 ;
        RECT 78.440 96.700 78.760 96.760 ;
        RECT 64.195 96.560 78.760 96.700 ;
        RECT 64.195 96.515 64.485 96.560 ;
        RECT 78.440 96.500 78.760 96.560 ;
        RECT 80.280 96.500 80.600 96.760 ;
        RECT 95.920 96.700 96.240 96.760 ;
        RECT 82.210 96.560 96.240 96.700 ;
        RECT 65.100 96.160 65.420 96.420 ;
        RECT 65.560 96.360 65.880 96.420 ;
        RECT 75.235 96.360 75.525 96.405 ;
        RECT 82.210 96.360 82.350 96.560 ;
        RECT 95.920 96.500 96.240 96.560 ;
        RECT 106.960 96.700 107.280 96.760 ;
        RECT 106.960 96.560 108.110 96.700 ;
        RECT 106.960 96.500 107.280 96.560 ;
        RECT 83.500 96.360 83.820 96.420 ;
        RECT 65.560 96.220 74.530 96.360 ;
        RECT 65.560 96.160 65.880 96.220 ;
        RECT 65.650 95.880 68.090 96.020 ;
        RECT 55.440 95.480 55.760 95.740 ;
        RECT 56.835 95.680 57.125 95.725 ;
        RECT 60.975 95.680 61.265 95.725 ;
        RECT 56.835 95.540 61.265 95.680 ;
        RECT 56.835 95.495 57.125 95.540 ;
        RECT 60.975 95.495 61.265 95.540 ;
        RECT 61.050 95.340 61.190 95.495 ;
        RECT 62.800 95.480 63.120 95.740 ;
        RECT 63.260 95.725 63.580 95.740 ;
        RECT 63.260 95.680 63.690 95.725 ;
        RECT 65.650 95.680 65.790 95.880 ;
        RECT 67.950 95.740 68.090 95.880 ;
        RECT 72.000 95.820 72.320 96.080 ;
        RECT 72.920 95.820 73.240 96.080 ;
        RECT 74.390 96.065 74.530 96.220 ;
        RECT 75.235 96.220 82.350 96.360 ;
        RECT 82.670 96.220 83.820 96.360 ;
        RECT 75.235 96.175 75.525 96.220 ;
        RECT 74.315 96.020 74.605 96.065 ;
        RECT 75.680 96.020 76.000 96.080 ;
        RECT 74.315 95.880 76.000 96.020 ;
        RECT 74.315 95.835 74.605 95.880 ;
        RECT 75.680 95.820 76.000 95.880 ;
        RECT 81.215 95.835 81.505 96.065 ;
        RECT 81.675 96.020 81.965 96.065 ;
        RECT 82.120 96.020 82.440 96.080 ;
        RECT 82.670 96.065 82.810 96.220 ;
        RECT 83.500 96.160 83.820 96.220 ;
        RECT 83.960 96.360 84.280 96.420 ;
        RECT 88.560 96.360 88.880 96.420 ;
        RECT 100.535 96.360 100.825 96.405 ;
        RECT 83.960 96.220 88.330 96.360 ;
        RECT 83.960 96.160 84.280 96.220 ;
        RECT 81.675 95.880 82.440 96.020 ;
        RECT 81.675 95.835 81.965 95.880 ;
        RECT 63.260 95.540 65.790 95.680 ;
        RECT 63.260 95.495 63.690 95.540 ;
        RECT 63.260 95.480 63.580 95.495 ;
        RECT 67.400 95.480 67.720 95.740 ;
        RECT 67.860 95.480 68.180 95.740 ;
        RECT 81.290 95.680 81.430 95.835 ;
        RECT 82.120 95.820 82.440 95.880 ;
        RECT 82.595 95.835 82.885 96.065 ;
        RECT 83.040 95.820 83.360 96.080 ;
        RECT 84.435 96.020 84.725 96.065 ;
        RECT 84.880 96.020 85.200 96.080 ;
        RECT 84.435 95.880 85.200 96.020 ;
        RECT 84.435 95.835 84.725 95.880 ;
        RECT 83.515 95.680 83.805 95.725 ;
        RECT 81.290 95.540 83.805 95.680 ;
        RECT 83.515 95.495 83.805 95.540 ;
        RECT 62.340 95.340 62.660 95.400 ;
        RECT 65.100 95.340 65.420 95.400 ;
        RECT 61.050 95.200 65.420 95.340 ;
        RECT 67.490 95.340 67.630 95.480 ;
        RECT 68.795 95.340 69.085 95.385 ;
        RECT 84.510 95.340 84.650 95.835 ;
        RECT 84.880 95.820 85.200 95.880 ;
        RECT 85.340 95.820 85.660 96.080 ;
        RECT 85.800 95.820 86.120 96.080 ;
        RECT 88.190 96.065 88.330 96.220 ;
        RECT 88.560 96.220 100.825 96.360 ;
        RECT 88.560 96.160 88.880 96.220 ;
        RECT 100.535 96.175 100.825 96.220 ;
        RECT 88.115 95.835 88.405 96.065 ;
        RECT 89.035 96.020 89.325 96.065 ;
        RECT 89.940 96.020 90.260 96.080 ;
        RECT 89.035 95.880 90.260 96.020 ;
        RECT 89.035 95.835 89.325 95.880 ;
        RECT 88.190 95.680 88.330 95.835 ;
        RECT 89.940 95.820 90.260 95.880 ;
        RECT 100.995 95.835 101.285 96.065 ;
        RECT 105.580 96.020 105.900 96.080 ;
        RECT 106.055 96.020 106.345 96.065 ;
        RECT 105.580 95.880 106.345 96.020 ;
        RECT 89.480 95.680 89.800 95.740 ;
        RECT 88.190 95.540 89.800 95.680 ;
        RECT 101.070 95.680 101.210 95.835 ;
        RECT 105.580 95.820 105.900 95.880 ;
        RECT 106.055 95.835 106.345 95.880 ;
        RECT 106.515 96.020 106.805 96.065 ;
        RECT 106.960 96.020 107.280 96.080 ;
        RECT 106.515 95.880 107.280 96.020 ;
        RECT 106.515 95.835 106.805 95.880 ;
        RECT 106.590 95.680 106.730 95.835 ;
        RECT 106.960 95.820 107.280 95.880 ;
        RECT 107.435 95.835 107.725 96.065 ;
        RECT 107.970 96.020 108.110 96.560 ;
        RECT 108.340 96.500 108.660 96.760 ;
        RECT 119.855 96.700 120.145 96.745 ;
        RECT 120.300 96.700 120.620 96.760 ;
        RECT 119.855 96.560 120.620 96.700 ;
        RECT 119.855 96.515 120.145 96.560 ;
        RECT 120.300 96.500 120.620 96.560 ;
        RECT 120.775 96.515 121.065 96.745 ;
        RECT 117.080 96.360 117.400 96.420 ;
        RECT 120.850 96.360 120.990 96.515 ;
        RECT 123.060 96.500 123.380 96.760 ;
        RECT 122.600 96.360 122.920 96.420 ;
        RECT 124.900 96.360 125.220 96.420 ;
        RECT 110.270 96.220 120.990 96.360 ;
        RECT 121.770 96.220 125.220 96.360 ;
        RECT 109.735 96.020 110.025 96.065 ;
        RECT 107.970 95.880 110.025 96.020 ;
        RECT 109.735 95.835 110.025 95.880 ;
        RECT 107.510 95.680 107.650 95.835 ;
        RECT 107.880 95.680 108.200 95.740 ;
        RECT 101.070 95.540 106.730 95.680 ;
        RECT 107.050 95.540 108.200 95.680 ;
        RECT 89.480 95.480 89.800 95.540 ;
        RECT 90.860 95.340 91.180 95.400 ;
        RECT 67.490 95.200 68.090 95.340 ;
        RECT 62.340 95.140 62.660 95.200 ;
        RECT 65.100 95.140 65.420 95.200 ;
        RECT 67.950 95.000 68.090 95.200 ;
        RECT 68.795 95.200 84.650 95.340 ;
        RECT 84.970 95.200 91.180 95.340 ;
        RECT 68.795 95.155 69.085 95.200 ;
        RECT 79.820 95.000 80.140 95.060 ;
        RECT 84.970 95.000 85.110 95.200 ;
        RECT 90.860 95.140 91.180 95.200 ;
        RECT 91.320 95.340 91.640 95.400 ;
        RECT 95.920 95.340 96.240 95.400 ;
        RECT 104.200 95.340 104.520 95.400 ;
        RECT 107.050 95.340 107.190 95.540 ;
        RECT 107.880 95.480 108.200 95.540 ;
        RECT 91.320 95.200 107.190 95.340 ;
        RECT 107.420 95.340 107.740 95.400 ;
        RECT 108.815 95.340 109.105 95.385 ;
        RECT 107.420 95.200 109.105 95.340 ;
        RECT 91.320 95.140 91.640 95.200 ;
        RECT 95.920 95.140 96.240 95.200 ;
        RECT 104.200 95.140 104.520 95.200 ;
        RECT 107.420 95.140 107.740 95.200 ;
        RECT 108.815 95.155 109.105 95.200 ;
        RECT 67.950 94.860 85.110 95.000 ;
        RECT 79.820 94.800 80.140 94.860 ;
        RECT 89.020 94.800 89.340 95.060 ;
        RECT 89.480 95.000 89.800 95.060 ;
        RECT 91.410 95.000 91.550 95.140 ;
        RECT 89.480 94.860 91.550 95.000 ;
        RECT 96.840 95.000 97.160 95.060 ;
        RECT 110.270 95.000 110.410 96.220 ;
        RECT 117.080 96.160 117.400 96.220 ;
        RECT 118.460 95.820 118.780 96.080 ;
        RECT 118.935 96.020 119.225 96.065 ;
        RECT 119.840 96.020 120.160 96.080 ;
        RECT 121.770 96.065 121.910 96.220 ;
        RECT 122.600 96.160 122.920 96.220 ;
        RECT 124.900 96.160 125.220 96.220 ;
        RECT 118.935 95.880 120.160 96.020 ;
        RECT 118.935 95.835 119.225 95.880 ;
        RECT 119.840 95.820 120.160 95.880 ;
        RECT 121.695 95.835 121.985 96.065 ;
        RECT 122.155 95.835 122.445 96.065 ;
        RECT 110.655 95.495 110.945 95.725 ;
        RECT 119.380 95.680 119.700 95.740 ;
        RECT 122.230 95.680 122.370 95.835 ;
        RECT 119.380 95.540 122.370 95.680 ;
        RECT 110.730 95.340 110.870 95.495 ;
        RECT 119.380 95.480 119.700 95.540 ;
        RECT 123.520 95.340 123.840 95.400 ;
        RECT 110.730 95.200 123.840 95.340 ;
        RECT 123.520 95.140 123.840 95.200 ;
        RECT 96.840 94.860 110.410 95.000 ;
        RECT 89.480 94.800 89.800 94.860 ;
        RECT 96.840 94.800 97.160 94.860 ;
        RECT 117.540 94.800 117.860 95.060 ;
        RECT 53.990 94.180 125.290 94.660 ;
        RECT 60.515 93.980 60.805 94.025 ;
        RECT 60.960 93.980 61.280 94.040 ;
        RECT 60.515 93.840 61.280 93.980 ;
        RECT 60.515 93.795 60.805 93.840 ;
        RECT 60.960 93.780 61.280 93.840 ;
        RECT 61.420 93.980 61.740 94.040 ;
        RECT 65.115 93.980 65.405 94.025 ;
        RECT 68.320 93.980 68.640 94.040 ;
        RECT 69.255 93.980 69.545 94.025 ;
        RECT 61.420 93.840 65.405 93.980 ;
        RECT 61.420 93.780 61.740 93.840 ;
        RECT 65.115 93.795 65.405 93.840 ;
        RECT 65.650 93.840 69.545 93.980 ;
        RECT 60.055 93.640 60.345 93.685 ;
        RECT 62.340 93.640 62.660 93.700 ;
        RECT 60.055 93.500 62.660 93.640 ;
        RECT 60.055 93.455 60.345 93.500 ;
        RECT 60.130 93.300 60.270 93.455 ;
        RECT 62.340 93.440 62.660 93.500 ;
        RECT 62.800 93.640 63.120 93.700 ;
        RECT 63.275 93.640 63.565 93.685 ;
        RECT 65.650 93.640 65.790 93.840 ;
        RECT 68.320 93.780 68.640 93.840 ;
        RECT 69.255 93.795 69.545 93.840 ;
        RECT 72.920 93.980 73.240 94.040 ;
        RECT 81.215 93.980 81.505 94.025 ;
        RECT 83.040 93.980 83.360 94.040 ;
        RECT 72.920 93.840 80.510 93.980 ;
        RECT 72.920 93.780 73.240 93.840 ;
        RECT 62.800 93.500 65.790 93.640 ;
        RECT 70.175 93.640 70.465 93.685 ;
        RECT 72.000 93.640 72.320 93.700 ;
        RECT 70.175 93.500 73.150 93.640 ;
        RECT 62.800 93.440 63.120 93.500 ;
        RECT 63.275 93.455 63.565 93.500 ;
        RECT 70.175 93.455 70.465 93.500 ;
        RECT 72.000 93.440 72.320 93.500 ;
        RECT 56.910 93.160 60.270 93.300 ;
        RECT 67.490 93.160 72.690 93.300 ;
        RECT 56.910 93.005 57.050 93.160 ;
        RECT 56.835 92.775 57.125 93.005 ;
        RECT 57.755 92.775 58.045 93.005 ;
        RECT 61.420 92.960 61.740 93.020 ;
        RECT 67.490 93.005 67.630 93.160 ;
        RECT 67.415 92.960 67.705 93.005 ;
        RECT 61.420 92.820 67.705 92.960 ;
        RECT 57.280 92.620 57.600 92.680 ;
        RECT 57.830 92.620 57.970 92.775 ;
        RECT 61.420 92.760 61.740 92.820 ;
        RECT 67.415 92.775 67.705 92.820 ;
        RECT 71.540 92.760 71.860 93.020 ;
        RECT 72.000 92.960 72.320 93.020 ;
        RECT 72.550 93.005 72.690 93.160 ;
        RECT 72.475 92.960 72.765 93.005 ;
        RECT 72.000 92.820 72.765 92.960 ;
        RECT 73.010 92.960 73.150 93.500 ;
        RECT 73.395 93.300 73.685 93.345 ;
        RECT 73.395 93.160 78.670 93.300 ;
        RECT 73.395 93.115 73.685 93.160 ;
        RECT 78.530 93.020 78.670 93.160 ;
        RECT 73.855 92.960 74.145 93.005 ;
        RECT 77.535 92.960 77.825 93.005 ;
        RECT 73.010 92.820 77.825 92.960 ;
        RECT 72.000 92.760 72.320 92.820 ;
        RECT 72.475 92.775 72.765 92.820 ;
        RECT 73.855 92.775 74.145 92.820 ;
        RECT 77.535 92.775 77.825 92.820 ;
        RECT 58.215 92.620 58.505 92.665 ;
        RECT 63.260 92.620 63.580 92.680 ;
        RECT 57.280 92.480 63.580 92.620 ;
        RECT 57.280 92.420 57.600 92.480 ;
        RECT 58.215 92.435 58.505 92.480 ;
        RECT 63.260 92.420 63.580 92.480 ;
        RECT 65.100 92.420 65.420 92.680 ;
        RECT 67.860 92.620 68.180 92.680 ;
        RECT 69.255 92.620 69.545 92.665 ;
        RECT 67.860 92.480 69.545 92.620 ;
        RECT 72.550 92.620 72.690 92.775 ;
        RECT 78.440 92.760 78.760 93.020 ;
        RECT 79.820 92.760 80.140 93.020 ;
        RECT 80.370 93.005 80.510 93.840 ;
        RECT 81.215 93.840 83.360 93.980 ;
        RECT 81.215 93.795 81.505 93.840 ;
        RECT 83.040 93.780 83.360 93.840 ;
        RECT 84.420 93.980 84.740 94.040 ;
        RECT 86.275 93.980 86.565 94.025 ;
        RECT 84.420 93.840 86.565 93.980 ;
        RECT 84.420 93.780 84.740 93.840 ;
        RECT 86.275 93.795 86.565 93.840 ;
        RECT 90.875 93.980 91.165 94.025 ;
        RECT 91.320 93.980 91.640 94.040 ;
        RECT 90.875 93.840 91.640 93.980 ;
        RECT 90.875 93.795 91.165 93.840 ;
        RECT 91.320 93.780 91.640 93.840 ;
        RECT 93.160 93.780 93.480 94.040 ;
        RECT 94.540 93.980 94.860 94.040 ;
        RECT 95.475 93.980 95.765 94.025 ;
        RECT 94.540 93.840 95.765 93.980 ;
        RECT 94.540 93.780 94.860 93.840 ;
        RECT 95.475 93.795 95.765 93.840 ;
        RECT 99.155 93.980 99.445 94.025 ;
        RECT 101.900 93.980 102.220 94.040 ;
        RECT 99.155 93.840 102.220 93.980 ;
        RECT 99.155 93.795 99.445 93.840 ;
        RECT 101.900 93.780 102.220 93.840 ;
        RECT 106.040 93.780 106.360 94.040 ;
        RECT 121.680 93.780 122.000 94.040 ;
        RECT 83.515 93.640 83.805 93.685 ;
        RECT 87.180 93.640 87.500 93.700 ;
        RECT 90.400 93.640 90.720 93.700 ;
        RECT 83.515 93.500 90.720 93.640 ;
        RECT 83.515 93.455 83.805 93.500 ;
        RECT 87.180 93.440 87.500 93.500 ;
        RECT 90.400 93.440 90.720 93.500 ;
        RECT 91.780 93.640 92.100 93.700 ;
        RECT 91.780 93.500 97.530 93.640 ;
        RECT 91.780 93.440 92.100 93.500 ;
        RECT 88.100 93.300 88.420 93.360 ;
        RECT 81.750 93.160 88.420 93.300 ;
        RECT 80.295 92.775 80.585 93.005 ;
        RECT 81.200 92.960 81.520 93.020 ;
        RECT 81.750 93.005 81.890 93.160 ;
        RECT 88.100 93.100 88.420 93.160 ;
        RECT 89.570 93.160 96.610 93.300 ;
        RECT 82.580 93.005 82.900 93.020 ;
        RECT 81.675 92.960 81.965 93.005 ;
        RECT 81.200 92.820 81.965 92.960 ;
        RECT 81.200 92.760 81.520 92.820 ;
        RECT 81.675 92.775 81.965 92.820 ;
        RECT 82.445 92.775 82.900 93.005 ;
        RECT 87.195 92.960 87.485 93.005 ;
        RECT 87.195 92.820 88.790 92.960 ;
        RECT 87.195 92.775 87.485 92.820 ;
        RECT 82.580 92.760 82.900 92.775 ;
        RECT 72.550 92.480 76.370 92.620 ;
        RECT 67.860 92.420 68.180 92.480 ;
        RECT 69.255 92.435 69.545 92.480 ;
        RECT 55.915 92.280 56.205 92.325 ;
        RECT 65.560 92.280 65.880 92.340 ;
        RECT 55.915 92.140 65.880 92.280 ;
        RECT 55.915 92.095 56.205 92.140 ;
        RECT 65.560 92.080 65.880 92.140 ;
        RECT 66.035 92.280 66.325 92.325 ;
        RECT 71.080 92.280 71.400 92.340 ;
        RECT 72.920 92.280 73.240 92.340 ;
        RECT 66.035 92.140 73.240 92.280 ;
        RECT 66.035 92.095 66.325 92.140 ;
        RECT 71.080 92.080 71.400 92.140 ;
        RECT 72.920 92.080 73.240 92.140 ;
        RECT 75.235 92.280 75.525 92.325 ;
        RECT 75.680 92.280 76.000 92.340 ;
        RECT 76.230 92.325 76.370 92.480 ;
        RECT 76.600 92.420 76.920 92.680 ;
        RECT 82.670 92.620 82.810 92.760 ;
        RECT 87.640 92.620 87.960 92.680 ;
        RECT 82.670 92.480 87.960 92.620 ;
        RECT 87.640 92.420 87.960 92.480 ;
        RECT 88.100 92.420 88.420 92.680 ;
        RECT 88.650 92.620 88.790 92.820 ;
        RECT 89.020 92.760 89.340 93.020 ;
        RECT 89.570 93.005 89.710 93.160 ;
        RECT 89.495 92.775 89.785 93.005 ;
        RECT 89.955 92.970 90.245 93.005 ;
        RECT 89.955 92.960 90.630 92.970 ;
        RECT 90.860 92.960 91.180 93.020 ;
        RECT 89.955 92.830 91.180 92.960 ;
        RECT 89.955 92.775 90.245 92.830 ;
        RECT 90.490 92.820 91.180 92.830 ;
        RECT 90.860 92.760 91.180 92.820 ;
        RECT 94.080 92.760 94.400 93.020 ;
        RECT 94.555 92.960 94.845 93.005 ;
        RECT 95.000 92.960 95.320 93.020 ;
        RECT 94.555 92.820 95.320 92.960 ;
        RECT 94.555 92.775 94.845 92.820 ;
        RECT 93.160 92.620 93.480 92.680 ;
        RECT 94.630 92.620 94.770 92.775 ;
        RECT 95.000 92.760 95.320 92.820 ;
        RECT 95.920 92.760 96.240 93.020 ;
        RECT 88.650 92.480 89.940 92.620 ;
        RECT 75.235 92.140 76.000 92.280 ;
        RECT 75.235 92.095 75.525 92.140 ;
        RECT 75.680 92.080 76.000 92.140 ;
        RECT 76.155 92.095 76.445 92.325 ;
        RECT 77.980 92.080 78.300 92.340 ;
        RECT 89.800 92.280 89.940 92.480 ;
        RECT 93.160 92.480 94.770 92.620 ;
        RECT 96.470 92.620 96.610 93.160 ;
        RECT 96.840 92.760 97.160 93.020 ;
        RECT 97.390 93.005 97.530 93.500 ;
        RECT 100.075 93.455 100.365 93.685 ;
        RECT 101.440 93.640 101.760 93.700 ;
        RECT 107.895 93.640 108.185 93.685 ;
        RECT 111.560 93.640 111.880 93.700 ;
        RECT 101.440 93.500 111.880 93.640 ;
        RECT 100.150 93.300 100.290 93.455 ;
        RECT 101.440 93.440 101.760 93.500 ;
        RECT 107.895 93.455 108.185 93.500 ;
        RECT 111.560 93.440 111.880 93.500 ;
        RECT 123.520 93.440 123.840 93.700 ;
        RECT 100.150 93.160 107.190 93.300 ;
        RECT 97.315 92.775 97.605 93.005 ;
        RECT 99.140 92.760 99.460 93.020 ;
        RECT 101.070 93.005 101.210 93.160 ;
        RECT 107.050 93.020 107.190 93.160 ;
        RECT 100.995 92.775 101.285 93.005 ;
        RECT 101.965 92.960 102.255 93.005 ;
        RECT 101.965 92.820 102.590 92.960 ;
        RECT 101.965 92.775 102.255 92.820 ;
        RECT 100.520 92.620 100.840 92.680 ;
        RECT 96.470 92.480 100.840 92.620 ;
        RECT 102.450 92.620 102.590 92.820 ;
        RECT 103.740 92.760 104.060 93.020 ;
        RECT 105.120 92.760 105.440 93.020 ;
        RECT 105.580 92.960 105.900 93.020 ;
        RECT 106.515 92.960 106.805 93.005 ;
        RECT 105.580 92.820 106.805 92.960 ;
        RECT 105.580 92.760 105.900 92.820 ;
        RECT 106.515 92.775 106.805 92.820 ;
        RECT 106.960 92.760 107.280 93.020 ;
        RECT 107.880 92.760 108.200 93.020 ;
        RECT 120.760 92.760 121.080 93.020 ;
        RECT 102.820 92.620 103.140 92.680 ;
        RECT 105.670 92.620 105.810 92.760 ;
        RECT 102.450 92.480 105.810 92.620 ;
        RECT 117.540 92.620 117.860 92.680 ;
        RECT 122.615 92.620 122.905 92.665 ;
        RECT 117.540 92.480 122.905 92.620 ;
        RECT 93.160 92.420 93.480 92.480 ;
        RECT 100.520 92.420 100.840 92.480 ;
        RECT 102.820 92.420 103.140 92.480 ;
        RECT 117.540 92.420 117.860 92.480 ;
        RECT 122.615 92.435 122.905 92.480 ;
        RECT 91.780 92.280 92.100 92.340 ;
        RECT 100.995 92.280 101.285 92.325 ;
        RECT 89.800 92.140 101.285 92.280 ;
        RECT 91.780 92.080 92.100 92.140 ;
        RECT 100.995 92.095 101.285 92.140 ;
        RECT 104.200 92.080 104.520 92.340 ;
        RECT 53.990 91.460 125.290 91.940 ;
        RECT 72.000 91.060 72.320 91.320 ;
        RECT 73.855 91.260 74.145 91.305 ;
        RECT 85.800 91.260 86.120 91.320 ;
        RECT 101.440 91.260 101.760 91.320 ;
        RECT 72.550 91.120 86.120 91.260 ;
        RECT 71.080 90.720 71.400 90.980 ;
        RECT 71.540 90.920 71.860 90.980 ;
        RECT 72.550 90.920 72.690 91.120 ;
        RECT 73.855 91.075 74.145 91.120 ;
        RECT 85.800 91.060 86.120 91.120 ;
        RECT 89.570 91.120 101.760 91.260 ;
        RECT 71.540 90.780 72.690 90.920 ;
        RECT 71.540 90.720 71.860 90.780 ;
        RECT 56.835 90.395 57.125 90.625 ;
        RECT 56.910 90.240 57.050 90.395 ;
        RECT 57.280 90.380 57.600 90.640 ;
        RECT 72.550 90.625 72.690 90.780 ;
        RECT 87.640 90.720 87.960 90.980 ;
        RECT 57.755 90.580 58.045 90.625 ;
        RECT 59.595 90.580 59.885 90.625 ;
        RECT 57.755 90.440 59.885 90.580 ;
        RECT 57.755 90.395 58.045 90.440 ;
        RECT 59.595 90.395 59.885 90.440 ;
        RECT 72.475 90.395 72.765 90.625 ;
        RECT 72.935 90.395 73.225 90.625 ;
        RECT 87.195 90.395 87.485 90.625 ;
        RECT 60.960 90.240 61.280 90.300 ;
        RECT 73.010 90.240 73.150 90.395 ;
        RECT 56.910 90.100 58.890 90.240 ;
        RECT 55.900 89.700 56.220 89.960 ;
        RECT 58.750 89.945 58.890 90.100 ;
        RECT 60.960 90.100 73.150 90.240 ;
        RECT 60.960 90.040 61.280 90.100 ;
        RECT 58.675 89.715 58.965 89.945 ;
        RECT 86.260 89.700 86.580 89.960 ;
        RECT 71.095 89.560 71.385 89.605 ;
        RECT 71.540 89.560 71.860 89.620 ;
        RECT 71.095 89.420 71.860 89.560 ;
        RECT 87.270 89.560 87.410 90.395 ;
        RECT 88.100 90.380 88.420 90.640 ;
        RECT 89.570 90.625 89.710 91.120 ;
        RECT 101.440 91.060 101.760 91.120 ;
        RECT 101.990 91.120 105.350 91.260 ;
        RECT 92.700 90.920 93.020 90.980 ;
        RECT 93.635 90.920 93.925 90.965 ;
        RECT 95.920 90.920 96.240 90.980 ;
        RECT 101.990 90.920 102.130 91.120 ;
        RECT 105.210 90.980 105.350 91.120 ;
        RECT 104.200 90.920 104.520 90.980 ;
        RECT 90.030 90.780 92.470 90.920 ;
        RECT 90.030 90.640 90.170 90.780 ;
        RECT 89.035 90.395 89.325 90.625 ;
        RECT 89.495 90.395 89.785 90.625 ;
        RECT 89.110 90.240 89.250 90.395 ;
        RECT 89.940 90.380 90.260 90.640 ;
        RECT 90.860 90.380 91.180 90.640 ;
        RECT 91.780 90.380 92.100 90.640 ;
        RECT 92.330 90.625 92.470 90.780 ;
        RECT 92.700 90.780 93.925 90.920 ;
        RECT 92.700 90.720 93.020 90.780 ;
        RECT 93.635 90.735 93.925 90.780 ;
        RECT 95.090 90.780 96.240 90.920 ;
        RECT 92.255 90.395 92.545 90.625 ;
        RECT 93.160 90.380 93.480 90.640 ;
        RECT 94.080 90.580 94.400 90.640 ;
        RECT 95.090 90.625 95.230 90.780 ;
        RECT 95.920 90.720 96.240 90.780 ;
        RECT 96.470 90.780 102.130 90.920 ;
        RECT 103.370 90.780 104.520 90.920 ;
        RECT 94.555 90.580 94.845 90.625 ;
        RECT 94.080 90.440 94.845 90.580 ;
        RECT 94.080 90.380 94.400 90.440 ;
        RECT 94.555 90.395 94.845 90.440 ;
        RECT 95.015 90.395 95.305 90.625 ;
        RECT 95.460 90.580 95.780 90.640 ;
        RECT 96.470 90.625 96.610 90.780 ;
        RECT 96.395 90.580 96.685 90.625 ;
        RECT 95.460 90.440 96.685 90.580 ;
        RECT 92.715 90.240 93.005 90.285 ;
        RECT 89.110 90.100 93.005 90.240 ;
        RECT 94.630 90.240 94.770 90.395 ;
        RECT 95.460 90.380 95.780 90.440 ;
        RECT 96.395 90.395 96.685 90.440 ;
        RECT 96.855 90.395 97.145 90.625 ;
        RECT 97.760 90.580 98.080 90.640 ;
        RECT 103.370 90.580 103.510 90.780 ;
        RECT 104.200 90.720 104.520 90.780 ;
        RECT 105.120 90.720 105.440 90.980 ;
        RECT 97.760 90.440 103.510 90.580 ;
        RECT 95.920 90.240 96.240 90.300 ;
        RECT 96.930 90.240 97.070 90.395 ;
        RECT 97.760 90.380 98.080 90.440 ;
        RECT 103.740 90.380 104.060 90.640 ;
        RECT 123.520 90.380 123.840 90.640 ;
        RECT 103.830 90.240 103.970 90.380 ;
        RECT 94.630 90.100 103.970 90.240 ;
        RECT 92.715 90.055 93.005 90.100 ;
        RECT 95.920 90.040 96.240 90.100 ;
        RECT 97.315 89.900 97.605 89.945 ;
        RECT 94.170 89.760 97.605 89.900 ;
        RECT 90.860 89.560 91.180 89.620 ;
        RECT 94.170 89.560 94.310 89.760 ;
        RECT 97.315 89.715 97.605 89.760 ;
        RECT 100.520 89.900 100.840 89.960 ;
        RECT 105.135 89.900 105.425 89.945 ;
        RECT 100.520 89.760 105.425 89.900 ;
        RECT 100.520 89.700 100.840 89.760 ;
        RECT 105.135 89.715 105.425 89.760 ;
        RECT 118.000 89.900 118.320 89.960 ;
        RECT 122.615 89.900 122.905 89.945 ;
        RECT 118.000 89.760 122.905 89.900 ;
        RECT 118.000 89.700 118.320 89.760 ;
        RECT 122.615 89.715 122.905 89.760 ;
        RECT 87.270 89.420 94.310 89.560 ;
        RECT 94.540 89.560 94.860 89.620 ;
        RECT 95.935 89.560 96.225 89.605 ;
        RECT 102.820 89.560 103.140 89.620 ;
        RECT 94.540 89.420 103.140 89.560 ;
        RECT 71.095 89.375 71.385 89.420 ;
        RECT 71.540 89.360 71.860 89.420 ;
        RECT 90.860 89.360 91.180 89.420 ;
        RECT 94.540 89.360 94.860 89.420 ;
        RECT 95.935 89.375 96.225 89.420 ;
        RECT 102.820 89.360 103.140 89.420 ;
        RECT 53.990 88.740 125.290 89.220 ;
        RECT 71.540 88.340 71.860 88.600 ;
        RECT 74.775 88.540 75.065 88.585 ;
        RECT 75.220 88.540 75.540 88.600 ;
        RECT 74.775 88.400 75.540 88.540 ;
        RECT 74.775 88.355 75.065 88.400 ;
        RECT 75.220 88.340 75.540 88.400 ;
        RECT 77.060 88.540 77.380 88.600 ;
        RECT 83.055 88.540 83.345 88.585 ;
        RECT 93.160 88.540 93.480 88.600 ;
        RECT 77.060 88.400 93.480 88.540 ;
        RECT 77.060 88.340 77.380 88.400 ;
        RECT 83.055 88.355 83.345 88.400 ;
        RECT 93.160 88.340 93.480 88.400 ;
        RECT 95.935 88.540 96.225 88.585 ;
        RECT 96.840 88.540 97.160 88.600 ;
        RECT 95.935 88.400 97.160 88.540 ;
        RECT 95.935 88.355 96.225 88.400 ;
        RECT 96.840 88.340 97.160 88.400 ;
        RECT 97.315 88.540 97.605 88.585 ;
        RECT 97.760 88.540 98.080 88.600 ;
        RECT 97.315 88.400 98.080 88.540 ;
        RECT 97.315 88.355 97.605 88.400 ;
        RECT 97.760 88.340 98.080 88.400 ;
        RECT 98.695 88.540 98.985 88.585 ;
        RECT 99.140 88.540 99.460 88.600 ;
        RECT 98.695 88.400 99.460 88.540 ;
        RECT 98.695 88.355 98.985 88.400 ;
        RECT 70.175 87.860 70.465 87.905 ;
        RECT 73.855 87.860 74.145 87.905 ;
        RECT 74.760 87.860 75.080 87.920 ;
        RECT 70.175 87.720 72.690 87.860 ;
        RECT 70.175 87.675 70.465 87.720 ;
        RECT 69.700 87.320 70.020 87.580 ;
        RECT 72.550 87.565 72.690 87.720 ;
        RECT 73.855 87.720 75.080 87.860 ;
        RECT 73.855 87.675 74.145 87.720 ;
        RECT 74.760 87.660 75.080 87.720 ;
        RECT 93.620 87.860 93.940 87.920 ;
        RECT 94.095 87.860 94.385 87.905 ;
        RECT 98.770 87.860 98.910 88.355 ;
        RECT 99.140 88.340 99.460 88.400 ;
        RECT 122.600 88.340 122.920 88.600 ;
        RECT 102.820 88.000 103.140 88.260 ;
        RECT 93.620 87.720 94.385 87.860 ;
        RECT 93.620 87.660 93.940 87.720 ;
        RECT 94.095 87.675 94.385 87.720 ;
        RECT 96.470 87.720 100.750 87.860 ;
        RECT 70.635 87.335 70.925 87.565 ;
        RECT 71.095 87.335 71.385 87.565 ;
        RECT 72.475 87.335 72.765 87.565 ;
        RECT 72.935 87.520 73.225 87.565 ;
        RECT 75.680 87.520 76.000 87.580 ;
        RECT 72.935 87.380 76.000 87.520 ;
        RECT 72.935 87.335 73.225 87.380 ;
        RECT 70.710 86.840 70.850 87.335 ;
        RECT 71.170 87.180 71.310 87.335 ;
        RECT 75.680 87.320 76.000 87.380 ;
        RECT 76.140 87.320 76.460 87.580 ;
        RECT 76.600 87.320 76.920 87.580 ;
        RECT 77.075 87.335 77.365 87.565 ;
        RECT 72.000 87.180 72.320 87.240 ;
        RECT 77.150 87.180 77.290 87.335 ;
        RECT 77.980 87.320 78.300 87.580 ;
        RECT 81.200 87.320 81.520 87.580 ;
        RECT 82.580 87.520 82.900 87.580 ;
        RECT 83.515 87.520 83.805 87.565 ;
        RECT 82.580 87.380 83.805 87.520 ;
        RECT 82.580 87.320 82.900 87.380 ;
        RECT 83.515 87.335 83.805 87.380 ;
        RECT 91.320 87.520 91.640 87.580 ;
        RECT 96.470 87.565 96.610 87.720 ;
        RECT 94.555 87.520 94.845 87.565 ;
        RECT 91.320 87.380 94.845 87.520 ;
        RECT 91.320 87.320 91.640 87.380 ;
        RECT 94.555 87.335 94.845 87.380 ;
        RECT 96.395 87.335 96.685 87.565 ;
        RECT 97.300 87.520 97.620 87.580 ;
        RECT 100.610 87.565 100.750 87.720 ;
        RECT 97.775 87.520 98.065 87.565 ;
        RECT 97.300 87.380 98.065 87.520 ;
        RECT 97.300 87.320 97.620 87.380 ;
        RECT 97.775 87.335 98.065 87.380 ;
        RECT 100.075 87.335 100.365 87.565 ;
        RECT 100.535 87.520 100.825 87.565 ;
        RECT 100.980 87.520 101.300 87.580 ;
        RECT 100.535 87.380 101.300 87.520 ;
        RECT 100.535 87.335 100.825 87.380 ;
        RECT 71.170 87.040 77.290 87.180 ;
        RECT 96.840 87.180 97.160 87.240 ;
        RECT 100.150 87.180 100.290 87.335 ;
        RECT 100.980 87.320 101.300 87.380 ;
        RECT 101.900 87.320 102.220 87.580 ;
        RECT 96.840 87.040 100.290 87.180 ;
        RECT 72.000 86.980 72.320 87.040 ;
        RECT 96.840 86.980 97.160 87.040 ;
        RECT 123.060 86.980 123.380 87.240 ;
        RECT 76.140 86.840 76.460 86.900 ;
        RECT 70.710 86.700 76.460 86.840 ;
        RECT 76.140 86.640 76.460 86.700 ;
        RECT 53.990 86.020 125.290 86.500 ;
        RECT 72.000 85.620 72.320 85.880 ;
        RECT 81.200 85.820 81.520 85.880 ;
        RECT 78.070 85.680 81.520 85.820 ;
        RECT 69.700 85.480 70.020 85.540 ;
        RECT 73.855 85.480 74.145 85.525 ;
        RECT 76.600 85.480 76.920 85.540 ;
        RECT 78.070 85.525 78.210 85.680 ;
        RECT 81.200 85.620 81.520 85.680 ;
        RECT 69.700 85.340 76.920 85.480 ;
        RECT 69.700 85.280 70.020 85.340 ;
        RECT 73.855 85.295 74.145 85.340 ;
        RECT 76.600 85.280 76.920 85.340 ;
        RECT 77.995 85.295 78.285 85.525 ;
        RECT 80.295 85.480 80.585 85.525 ;
        RECT 82.580 85.480 82.900 85.540 ;
        RECT 80.295 85.340 82.900 85.480 ;
        RECT 80.295 85.295 80.585 85.340 ;
        RECT 64.640 85.140 64.960 85.200 ;
        RECT 73.395 85.140 73.685 85.185 ;
        RECT 64.640 85.000 73.685 85.140 ;
        RECT 64.640 84.940 64.960 85.000 ;
        RECT 73.395 84.955 73.685 85.000 ;
        RECT 74.775 85.140 75.065 85.185 ;
        RECT 77.075 85.140 77.365 85.185 ;
        RECT 80.370 85.140 80.510 85.295 ;
        RECT 82.580 85.280 82.900 85.340 ;
        RECT 95.920 85.480 96.240 85.540 ;
        RECT 98.695 85.480 98.985 85.525 ;
        RECT 95.920 85.340 98.985 85.480 ;
        RECT 95.920 85.280 96.240 85.340 ;
        RECT 98.695 85.295 98.985 85.340 ;
        RECT 74.775 85.000 80.510 85.140 ;
        RECT 80.740 85.140 81.060 85.200 ;
        RECT 81.215 85.140 81.505 85.185 ;
        RECT 80.740 85.000 81.505 85.140 ;
        RECT 74.775 84.955 75.065 85.000 ;
        RECT 77.075 84.955 77.365 85.000 ;
        RECT 71.540 84.800 71.860 84.860 ;
        RECT 72.015 84.800 72.305 84.845 ;
        RECT 71.540 84.660 72.305 84.800 ;
        RECT 73.470 84.800 73.610 84.955 ;
        RECT 80.740 84.940 81.060 85.000 ;
        RECT 81.215 84.955 81.505 85.000 ;
        RECT 82.135 85.140 82.425 85.185 ;
        RECT 85.340 85.140 85.660 85.200 ;
        RECT 82.135 85.000 85.660 85.140 ;
        RECT 82.135 84.955 82.425 85.000 ;
        RECT 85.340 84.940 85.660 85.000 ;
        RECT 99.615 84.955 99.905 85.185 ;
        RECT 75.695 84.800 75.985 84.845 ;
        RECT 96.840 84.800 97.160 84.860 ;
        RECT 99.690 84.800 99.830 84.955 ;
        RECT 100.980 84.940 101.300 85.200 ;
        RECT 101.900 84.940 102.220 85.200 ;
        RECT 73.470 84.660 99.830 84.800 ;
        RECT 71.540 84.600 71.860 84.660 ;
        RECT 72.015 84.615 72.305 84.660 ;
        RECT 75.695 84.615 75.985 84.660 ;
        RECT 72.090 84.460 72.230 84.615 ;
        RECT 96.840 84.600 97.160 84.660 ;
        RECT 123.520 84.600 123.840 84.860 ;
        RECT 78.915 84.460 79.205 84.505 ;
        RECT 93.620 84.460 93.940 84.520 ;
        RECT 72.090 84.320 79.205 84.460 ;
        RECT 78.915 84.275 79.205 84.320 ;
        RECT 82.670 84.320 93.940 84.460 ;
        RECT 72.935 84.120 73.225 84.165 ;
        RECT 78.440 84.120 78.760 84.180 ;
        RECT 82.670 84.120 82.810 84.320 ;
        RECT 93.620 84.260 93.940 84.320 ;
        RECT 72.935 83.980 82.810 84.120 ;
        RECT 83.055 84.120 83.345 84.165 ;
        RECT 84.420 84.120 84.740 84.180 ;
        RECT 83.055 83.980 84.740 84.120 ;
        RECT 72.935 83.935 73.225 83.980 ;
        RECT 78.440 83.920 78.760 83.980 ;
        RECT 83.055 83.935 83.345 83.980 ;
        RECT 84.420 83.920 84.740 83.980 ;
        RECT 53.990 83.300 125.290 83.780 ;
        RECT 71.555 83.100 71.845 83.145 ;
        RECT 72.460 83.100 72.780 83.160 ;
        RECT 71.555 82.960 72.780 83.100 ;
        RECT 71.555 82.915 71.845 82.960 ;
        RECT 72.460 82.900 72.780 82.960 ;
        RECT 76.140 83.100 76.460 83.160 ;
        RECT 77.075 83.100 77.365 83.145 ;
        RECT 76.140 82.960 77.365 83.100 ;
        RECT 76.140 82.900 76.460 82.960 ;
        RECT 77.075 82.915 77.365 82.960 ;
        RECT 78.915 83.100 79.205 83.145 ;
        RECT 80.740 83.100 81.060 83.160 ;
        RECT 78.915 82.960 81.060 83.100 ;
        RECT 78.915 82.915 79.205 82.960 ;
        RECT 80.740 82.900 81.060 82.960 ;
        RECT 81.200 83.100 81.520 83.160 ;
        RECT 82.135 83.100 82.425 83.145 ;
        RECT 81.200 82.960 82.425 83.100 ;
        RECT 81.200 82.900 81.520 82.960 ;
        RECT 82.135 82.915 82.425 82.960 ;
        RECT 75.695 82.760 75.985 82.805 ;
        RECT 79.820 82.760 80.140 82.820 ;
        RECT 75.695 82.620 80.140 82.760 ;
        RECT 75.695 82.575 75.985 82.620 ;
        RECT 79.820 82.560 80.140 82.620 ;
        RECT 78.440 82.420 78.760 82.480 ;
        RECT 76.690 82.280 78.760 82.420 ;
        RECT 61.420 82.080 61.740 82.140 ;
        RECT 61.895 82.080 62.185 82.125 ;
        RECT 61.420 81.940 62.185 82.080 ;
        RECT 61.420 81.880 61.740 81.940 ;
        RECT 61.895 81.895 62.185 81.940 ;
        RECT 71.080 82.080 71.400 82.140 ;
        RECT 72.475 82.080 72.765 82.125 ;
        RECT 71.080 81.940 72.765 82.080 ;
        RECT 71.080 81.880 71.400 81.940 ;
        RECT 72.475 81.895 72.765 81.940 ;
        RECT 74.760 81.880 75.080 82.140 ;
        RECT 76.690 82.125 76.830 82.280 ;
        RECT 78.440 82.220 78.760 82.280 ;
        RECT 76.615 81.895 76.905 82.125 ;
        RECT 77.535 81.895 77.825 82.125 ;
        RECT 77.610 81.740 77.750 81.895 ;
        RECT 77.980 81.880 78.300 82.140 ;
        RECT 81.200 82.080 81.520 82.140 ;
        RECT 78.530 81.940 81.520 82.080 ;
        RECT 78.530 81.740 78.670 81.940 ;
        RECT 81.200 81.880 81.520 81.940 ;
        RECT 84.420 81.880 84.740 82.140 ;
        RECT 77.610 81.600 78.670 81.740 ;
        RECT 80.740 81.740 81.060 81.800 ;
        RECT 81.675 81.740 81.965 81.785 ;
        RECT 80.740 81.600 81.965 81.740 ;
        RECT 80.740 81.540 81.060 81.600 ;
        RECT 81.675 81.555 81.965 81.600 ;
        RECT 83.960 81.400 84.280 81.460 ;
        RECT 85.355 81.400 85.645 81.445 ;
        RECT 83.960 81.260 85.645 81.400 ;
        RECT 83.960 81.200 84.280 81.260 ;
        RECT 85.355 81.215 85.645 81.260 ;
        RECT 53.990 80.580 125.290 81.060 ;
      LAYER met2 ;
        RECT 48.560 159.010 48.840 163.010 ;
        RECT 51.780 159.010 52.060 163.010 ;
        RECT 55.000 159.010 55.280 163.010 ;
        RECT 58.220 159.010 58.500 163.010 ;
        RECT 61.440 159.010 61.720 163.010 ;
        RECT 64.660 159.010 64.940 163.010 ;
        RECT 67.880 159.010 68.160 163.010 ;
        RECT 71.100 159.010 71.380 163.010 ;
        RECT 74.320 159.010 74.600 163.010 ;
        RECT 74.850 159.290 76.370 159.430 ;
        RECT 48.630 156.145 48.770 159.010 ;
        RECT 48.560 155.775 48.840 156.145 ;
        RECT 51.850 122.825 51.990 159.010 ;
        RECT 52.710 152.910 52.970 153.230 ;
        RECT 52.770 133.590 52.910 152.910 ;
        RECT 53.620 151.695 53.900 152.065 ;
        RECT 53.690 148.470 53.830 151.695 ;
        RECT 55.070 149.910 55.210 159.010 ;
        RECT 57.770 155.630 58.030 155.950 ;
        RECT 55.470 153.590 55.730 153.910 ;
        RECT 54.610 149.770 55.210 149.910 ;
        RECT 53.630 148.150 53.890 148.470 ;
        RECT 53.170 146.790 53.430 147.110 ;
        RECT 53.230 139.710 53.370 146.790 ;
        RECT 54.090 146.450 54.350 146.770 ;
        RECT 53.630 142.370 53.890 142.690 ;
        RECT 53.690 141.865 53.830 142.370 ;
        RECT 53.620 141.495 53.900 141.865 ;
        RECT 53.230 139.570 53.830 139.710 ;
        RECT 53.160 134.695 53.440 135.065 ;
        RECT 53.230 134.530 53.370 134.695 ;
        RECT 53.170 134.210 53.430 134.530 ;
        RECT 52.770 133.450 53.370 133.590 ;
        RECT 52.710 132.850 52.970 133.170 ;
        RECT 52.770 132.345 52.910 132.850 ;
        RECT 52.700 131.975 52.980 132.345 ;
        RECT 52.700 129.255 52.980 129.625 ;
        RECT 52.710 129.110 52.970 129.255 ;
        RECT 51.780 122.455 52.060 122.825 ;
        RECT 53.230 117.530 53.370 133.450 ;
        RECT 53.690 118.210 53.830 139.570 ;
        RECT 54.150 123.310 54.290 146.450 ;
        RECT 54.610 145.750 54.750 149.770 ;
        RECT 55.000 148.295 55.280 148.665 ;
        RECT 54.550 145.430 54.810 145.750 ;
        RECT 54.540 144.895 54.820 145.265 ;
        RECT 54.610 123.990 54.750 144.895 ;
        RECT 54.550 123.670 54.810 123.990 ;
        RECT 54.090 122.990 54.350 123.310 ;
        RECT 55.070 122.630 55.210 148.295 ;
        RECT 55.530 131.810 55.670 153.590 ;
        RECT 56.840 152.375 57.120 152.745 ;
        RECT 56.910 150.510 57.050 152.375 ;
        RECT 57.830 151.190 57.970 155.630 ;
        RECT 58.290 153.230 58.430 159.010 ;
        RECT 58.680 158.495 58.960 158.865 ;
        RECT 58.230 152.910 58.490 153.230 ;
        RECT 57.770 150.870 58.030 151.190 ;
        RECT 56.850 150.190 57.110 150.510 ;
        RECT 57.770 147.810 58.030 148.130 ;
        RECT 57.310 147.305 57.570 147.450 ;
        RECT 57.300 146.935 57.580 147.305 ;
        RECT 57.310 146.450 57.570 146.770 ;
        RECT 57.370 145.070 57.510 146.450 ;
        RECT 57.830 145.750 57.970 147.810 ;
        RECT 57.770 145.430 58.030 145.750 ;
        RECT 56.390 144.750 56.650 145.070 ;
        RECT 57.310 144.750 57.570 145.070 ;
        RECT 55.930 138.465 56.190 138.610 ;
        RECT 55.920 138.095 56.200 138.465 ;
        RECT 55.930 133.530 56.190 133.850 ;
        RECT 55.470 131.490 55.730 131.810 ;
        RECT 55.470 125.370 55.730 125.690 ;
        RECT 55.530 124.865 55.670 125.370 ;
        RECT 55.460 124.495 55.740 124.865 ;
        RECT 55.010 122.310 55.270 122.630 ;
        RECT 53.630 117.890 53.890 118.210 ;
        RECT 55.460 117.695 55.740 118.065 ;
        RECT 55.470 117.550 55.730 117.695 ;
        RECT 53.170 117.210 53.430 117.530 ;
        RECT 55.990 115.150 56.130 133.530 ;
        RECT 56.450 122.290 56.590 144.750 ;
        RECT 57.770 141.690 58.030 142.010 ;
        RECT 56.850 139.310 57.110 139.630 ;
        RECT 56.910 134.870 57.050 139.310 ;
        RECT 57.830 136.570 57.970 141.690 ;
        RECT 58.230 141.010 58.490 141.330 ;
        RECT 58.290 136.910 58.430 141.010 ;
        RECT 58.750 140.310 58.890 158.495 ;
        RECT 60.530 154.610 60.790 154.930 ;
        RECT 60.070 151.890 60.330 152.210 ;
        RECT 59.140 151.015 59.420 151.385 ;
        RECT 59.210 140.310 59.350 151.015 ;
        RECT 60.130 145.070 60.270 151.890 ;
        RECT 59.610 144.750 59.870 145.070 ;
        RECT 60.070 144.750 60.330 145.070 ;
        RECT 59.670 143.225 59.810 144.750 ;
        RECT 59.600 142.855 59.880 143.225 ;
        RECT 60.590 143.030 60.730 154.610 ;
        RECT 60.990 153.930 61.250 154.250 ;
        RECT 61.050 151.190 61.190 153.930 ;
        RECT 61.510 153.425 61.650 159.010 ;
        RECT 62.370 154.270 62.630 154.590 ;
        RECT 61.440 153.055 61.720 153.425 ;
        RECT 60.990 150.870 61.250 151.190 ;
        RECT 62.430 150.850 62.570 154.270 ;
        RECT 62.370 150.530 62.630 150.850 ;
        RECT 61.910 150.190 62.170 150.510 ;
        RECT 61.970 150.025 62.110 150.190 ;
        RECT 61.900 149.655 62.180 150.025 ;
        RECT 61.450 147.810 61.710 148.130 ;
        RECT 61.510 146.770 61.650 147.810 ;
        RECT 62.430 147.450 62.570 150.530 ;
        RECT 63.290 150.190 63.550 150.510 ;
        RECT 62.830 148.150 63.090 148.470 ;
        RECT 62.370 147.130 62.630 147.450 ;
        RECT 61.450 146.450 61.710 146.770 ;
        RECT 61.900 146.255 62.180 146.625 ;
        RECT 61.440 145.575 61.720 145.945 ;
        RECT 61.970 145.750 62.110 146.255 ;
        RECT 60.530 142.710 60.790 143.030 ;
        RECT 61.510 142.010 61.650 145.575 ;
        RECT 61.910 145.430 62.170 145.750 ;
        RECT 62.370 144.750 62.630 145.070 ;
        RECT 61.910 143.730 62.170 144.050 ;
        RECT 59.610 141.690 59.870 142.010 ;
        RECT 60.990 141.865 61.250 142.010 ;
        RECT 58.690 139.990 58.950 140.310 ;
        RECT 59.150 139.990 59.410 140.310 ;
        RECT 58.230 136.590 58.490 136.910 ;
        RECT 57.770 136.250 58.030 136.570 ;
        RECT 57.310 135.910 57.570 136.230 ;
        RECT 56.850 134.550 57.110 134.870 ;
        RECT 56.850 133.870 57.110 134.190 ;
        RECT 56.910 131.130 57.050 133.870 ;
        RECT 57.370 133.170 57.510 135.910 ;
        RECT 57.310 132.850 57.570 133.170 ;
        RECT 56.850 130.810 57.110 131.130 ;
        RECT 56.850 130.130 57.110 130.450 ;
        RECT 56.910 128.750 57.050 130.130 ;
        RECT 56.850 128.430 57.110 128.750 ;
        RECT 56.850 123.330 57.110 123.650 ;
        RECT 56.390 121.970 56.650 122.290 ;
        RECT 56.910 121.350 57.050 123.330 ;
        RECT 57.370 122.880 57.510 132.850 ;
        RECT 57.830 126.710 57.970 136.250 ;
        RECT 58.290 131.550 58.430 136.590 ;
        RECT 58.690 135.910 58.950 136.230 ;
        RECT 58.750 133.170 58.890 135.910 ;
        RECT 59.150 134.550 59.410 134.870 ;
        RECT 58.690 132.850 58.950 133.170 ;
        RECT 58.290 131.410 58.890 131.550 ;
        RECT 58.230 130.810 58.490 131.130 ;
        RECT 57.770 126.390 58.030 126.710 ;
        RECT 57.770 122.880 58.030 122.970 ;
        RECT 57.370 122.740 58.030 122.880 ;
        RECT 57.770 122.650 58.030 122.740 ;
        RECT 56.450 121.210 57.050 121.350 ;
        RECT 56.450 116.850 56.590 121.210 ;
        RECT 58.290 120.250 58.430 130.810 ;
        RECT 58.750 129.625 58.890 131.410 ;
        RECT 59.210 131.130 59.350 134.550 ;
        RECT 59.670 132.150 59.810 141.690 ;
        RECT 60.980 141.495 61.260 141.865 ;
        RECT 61.450 141.690 61.710 142.010 ;
        RECT 61.450 141.010 61.710 141.330 ;
        RECT 60.530 139.650 60.790 139.970 ;
        RECT 60.070 138.970 60.330 139.290 ;
        RECT 59.610 131.830 59.870 132.150 ;
        RECT 59.150 130.810 59.410 131.130 ;
        RECT 58.680 129.255 58.960 129.625 ;
        RECT 60.130 129.430 60.270 138.970 ;
        RECT 60.590 136.480 60.730 139.650 ;
        RECT 61.510 139.630 61.650 141.010 ;
        RECT 60.990 139.310 61.250 139.630 ;
        RECT 61.450 139.310 61.710 139.630 ;
        RECT 61.050 137.590 61.190 139.310 ;
        RECT 60.990 137.270 61.250 137.590 ;
        RECT 61.510 137.250 61.650 139.310 ;
        RECT 61.450 136.930 61.710 137.250 ;
        RECT 60.990 136.480 61.250 136.570 ;
        RECT 60.590 136.340 61.250 136.480 ;
        RECT 60.990 136.250 61.250 136.340 ;
        RECT 60.520 135.375 60.800 135.745 ;
        RECT 60.590 134.190 60.730 135.375 ;
        RECT 60.530 133.870 60.790 134.190 ;
        RECT 61.050 133.760 61.190 136.250 ;
        RECT 61.440 134.695 61.720 135.065 ;
        RECT 61.450 134.550 61.710 134.695 ;
        RECT 61.450 133.760 61.710 133.850 ;
        RECT 61.050 133.620 61.710 133.760 ;
        RECT 61.050 131.470 61.190 133.620 ;
        RECT 61.450 133.530 61.710 133.620 ;
        RECT 61.970 133.590 62.110 143.730 ;
        RECT 62.430 143.225 62.570 144.750 ;
        RECT 62.360 142.855 62.640 143.225 ;
        RECT 62.370 141.350 62.630 141.670 ;
        RECT 62.430 141.185 62.570 141.350 ;
        RECT 62.890 141.330 63.030 148.150 ;
        RECT 63.350 147.110 63.490 150.190 ;
        RECT 64.210 149.170 64.470 149.490 ;
        RECT 64.270 147.985 64.410 149.170 ;
        RECT 64.200 147.615 64.480 147.985 ;
        RECT 64.210 147.130 64.470 147.450 ;
        RECT 63.290 146.790 63.550 147.110 ;
        RECT 63.750 146.790 64.010 147.110 ;
        RECT 63.350 144.730 63.490 146.790 ;
        RECT 63.810 145.750 63.950 146.790 ;
        RECT 63.750 145.430 64.010 145.750 ;
        RECT 63.740 144.895 64.020 145.265 ;
        RECT 64.270 145.070 64.410 147.130 ;
        RECT 63.750 144.750 64.010 144.895 ;
        RECT 64.210 144.750 64.470 145.070 ;
        RECT 63.290 144.410 63.550 144.730 ;
        RECT 64.270 144.470 64.410 144.750 ;
        RECT 63.810 144.330 64.410 144.470 ;
        RECT 63.280 143.535 63.560 143.905 ;
        RECT 63.350 141.330 63.490 143.535 ;
        RECT 62.360 140.815 62.640 141.185 ;
        RECT 62.830 141.010 63.090 141.330 ;
        RECT 63.290 141.010 63.550 141.330 ;
        RECT 63.810 140.505 63.950 144.330 ;
        RECT 64.210 143.730 64.470 144.050 ;
        RECT 63.740 140.135 64.020 140.505 ;
        RECT 63.290 139.880 63.550 139.970 ;
        RECT 63.290 139.740 63.950 139.880 ;
        RECT 63.290 139.650 63.550 139.740 ;
        RECT 62.370 139.310 62.630 139.630 ;
        RECT 62.430 136.910 62.570 139.310 ;
        RECT 63.290 138.970 63.550 139.290 ;
        RECT 62.820 137.415 63.100 137.785 ;
        RECT 62.370 136.590 62.630 136.910 ;
        RECT 62.890 135.890 63.030 137.415 ;
        RECT 63.350 136.570 63.490 138.970 ;
        RECT 63.810 137.785 63.950 139.740 ;
        RECT 64.270 139.290 64.410 143.730 ;
        RECT 64.210 138.970 64.470 139.290 ;
        RECT 63.740 137.415 64.020 137.785 ;
        RECT 63.290 136.480 63.550 136.570 ;
        RECT 63.290 136.340 63.950 136.480 ;
        RECT 63.290 136.250 63.550 136.340 ;
        RECT 62.830 135.570 63.090 135.890 ;
        RECT 63.290 135.570 63.550 135.890 ;
        RECT 63.350 134.190 63.490 135.570 ;
        RECT 63.810 134.870 63.950 136.340 ;
        RECT 64.210 136.250 64.470 136.570 ;
        RECT 64.730 136.425 64.870 159.010 ;
        RECT 67.420 153.735 67.700 154.105 ;
        RECT 67.950 153.910 68.090 159.010 ;
        RECT 68.350 154.270 68.610 154.590 ;
        RECT 66.040 153.055 66.320 153.425 ;
        RECT 65.590 152.570 65.850 152.890 ;
        RECT 65.130 150.870 65.390 151.190 ;
        RECT 65.190 148.470 65.330 150.870 ;
        RECT 65.650 150.510 65.790 152.570 ;
        RECT 65.590 150.190 65.850 150.510 ;
        RECT 66.110 149.490 66.250 153.055 ;
        RECT 66.970 152.230 67.230 152.550 ;
        RECT 66.500 150.335 66.780 150.705 ;
        RECT 66.510 150.190 66.770 150.335 ;
        RECT 67.030 150.170 67.170 152.230 ;
        RECT 66.970 149.850 67.230 150.170 ;
        RECT 67.490 149.830 67.630 153.735 ;
        RECT 67.890 153.590 68.150 153.910 ;
        RECT 67.890 149.850 68.150 150.170 ;
        RECT 67.430 149.510 67.690 149.830 ;
        RECT 66.050 149.170 66.310 149.490 ;
        RECT 66.510 149.170 66.770 149.490 ;
        RECT 65.130 148.150 65.390 148.470 ;
        RECT 65.590 147.810 65.850 148.130 ;
        RECT 65.120 146.935 65.400 147.305 ;
        RECT 65.190 137.590 65.330 146.935 ;
        RECT 65.650 144.050 65.790 147.810 ;
        RECT 66.570 147.790 66.710 149.170 ;
        RECT 67.430 148.150 67.690 148.470 ;
        RECT 66.510 147.470 66.770 147.790 ;
        RECT 66.050 147.130 66.310 147.450 ;
        RECT 66.110 146.625 66.250 147.130 ;
        RECT 66.040 146.255 66.320 146.625 ;
        RECT 66.970 146.450 67.230 146.770 ;
        RECT 66.510 145.265 66.770 145.410 ;
        RECT 66.500 144.895 66.780 145.265 ;
        RECT 67.030 145.070 67.170 146.450 ;
        RECT 66.970 144.750 67.230 145.070 ;
        RECT 66.050 144.070 66.310 144.390 ;
        RECT 65.590 143.730 65.850 144.050 ;
        RECT 65.590 142.030 65.850 142.350 ;
        RECT 65.130 137.270 65.390 137.590 ;
        RECT 63.750 134.550 64.010 134.870 ;
        RECT 63.290 133.870 63.550 134.190 ;
        RECT 61.970 133.450 63.030 133.590 ;
        RECT 62.370 132.850 62.630 133.170 ;
        RECT 61.910 131.720 62.170 131.810 ;
        RECT 61.510 131.580 62.170 131.720 ;
        RECT 60.990 131.150 61.250 131.470 ;
        RECT 60.980 130.615 61.260 130.985 ;
        RECT 60.530 130.130 60.790 130.450 ;
        RECT 60.070 129.110 60.330 129.430 ;
        RECT 59.610 129.000 59.870 129.090 ;
        RECT 58.750 128.860 59.870 129.000 ;
        RECT 58.750 125.690 58.890 128.860 ;
        RECT 59.610 128.770 59.870 128.860 ;
        RECT 60.130 128.750 60.270 129.110 ;
        RECT 60.590 128.750 60.730 130.130 ;
        RECT 60.070 128.430 60.330 128.750 ;
        RECT 60.530 128.430 60.790 128.750 ;
        RECT 60.130 126.370 60.270 128.430 ;
        RECT 60.070 126.050 60.330 126.370 ;
        RECT 58.690 125.600 58.950 125.690 ;
        RECT 58.690 125.460 59.350 125.600 ;
        RECT 58.690 125.370 58.950 125.460 ;
        RECT 58.680 123.135 58.960 123.505 ;
        RECT 58.690 122.990 58.950 123.135 ;
        RECT 59.210 121.270 59.350 125.460 ;
        RECT 60.130 125.350 60.270 126.050 ;
        RECT 60.590 125.690 60.730 128.430 ;
        RECT 61.050 128.410 61.190 130.615 ;
        RECT 60.990 128.090 61.250 128.410 ;
        RECT 61.510 128.070 61.650 131.580 ;
        RECT 61.910 131.490 62.170 131.580 ;
        RECT 62.430 130.790 62.570 132.850 ;
        RECT 62.370 130.700 62.630 130.790 ;
        RECT 61.970 130.560 62.630 130.700 ;
        RECT 61.970 129.430 62.110 130.560 ;
        RECT 62.370 130.470 62.630 130.560 ;
        RECT 61.910 129.110 62.170 129.430 ;
        RECT 62.360 129.255 62.640 129.625 ;
        RECT 61.450 127.750 61.710 128.070 ;
        RECT 61.510 126.030 61.650 127.750 ;
        RECT 61.450 125.710 61.710 126.030 ;
        RECT 60.530 125.370 60.790 125.690 ;
        RECT 60.070 125.030 60.330 125.350 ;
        RECT 60.590 123.990 60.730 125.370 ;
        RECT 61.970 125.010 62.110 129.110 ;
        RECT 62.430 128.410 62.570 129.255 ;
        RECT 62.370 128.090 62.630 128.410 ;
        RECT 61.910 124.690 62.170 125.010 ;
        RECT 60.530 123.670 60.790 123.990 ;
        RECT 61.900 123.815 62.180 124.185 ;
        RECT 59.150 120.950 59.410 121.270 ;
        RECT 58.230 119.930 58.490 120.250 ;
        RECT 57.770 119.250 58.030 119.570 ;
        RECT 58.230 119.250 58.490 119.570 ;
        RECT 57.830 117.870 57.970 119.250 ;
        RECT 57.770 117.550 58.030 117.870 ;
        RECT 56.390 116.530 56.650 116.850 ;
        RECT 55.930 114.830 56.190 115.150 ;
        RECT 56.450 111.945 56.590 116.530 ;
        RECT 57.310 114.490 57.570 114.810 ;
        RECT 56.380 111.575 56.660 111.945 ;
        RECT 57.370 110.390 57.510 114.490 ;
        RECT 57.310 110.070 57.570 110.390 ;
        RECT 57.310 108.370 57.570 108.690 ;
        RECT 55.920 100.695 56.200 101.065 ;
        RECT 55.930 100.550 56.190 100.695 ;
        RECT 57.370 99.510 57.510 108.370 ;
        RECT 58.290 107.670 58.430 119.250 ;
        RECT 58.690 114.830 58.950 115.150 ;
        RECT 58.750 113.110 58.890 114.830 ;
        RECT 58.690 112.790 58.950 113.110 ;
        RECT 59.210 112.510 59.350 120.950 ;
        RECT 60.590 119.910 60.730 123.670 ;
        RECT 61.970 123.310 62.110 123.815 ;
        RECT 60.990 122.990 61.250 123.310 ;
        RECT 61.910 122.990 62.170 123.310 ;
        RECT 61.050 122.290 61.190 122.990 ;
        RECT 60.990 121.970 61.250 122.290 ;
        RECT 61.970 120.250 62.110 122.990 ;
        RECT 62.430 122.710 62.570 128.090 ;
        RECT 62.890 123.310 63.030 133.450 ;
        RECT 64.270 133.170 64.410 136.250 ;
        RECT 64.660 136.055 64.940 136.425 ;
        RECT 65.130 135.910 65.390 136.230 ;
        RECT 64.670 133.870 64.930 134.190 ;
        RECT 64.730 133.510 64.870 133.870 ;
        RECT 64.670 133.190 64.930 133.510 ;
        RECT 64.210 132.850 64.470 133.170 ;
        RECT 64.730 131.665 64.870 133.190 ;
        RECT 65.190 132.150 65.330 135.910 ;
        RECT 65.130 131.830 65.390 132.150 ;
        RECT 64.660 131.295 64.940 131.665 ;
        RECT 64.670 131.040 64.930 131.130 ;
        RECT 65.190 131.040 65.330 131.830 ;
        RECT 65.650 131.380 65.790 142.030 ;
        RECT 66.110 132.345 66.250 144.070 ;
        RECT 66.510 143.730 66.770 144.050 ;
        RECT 66.970 143.730 67.230 144.050 ;
        RECT 66.570 137.590 66.710 143.730 ;
        RECT 66.510 137.270 66.770 137.590 ;
        RECT 66.500 136.735 66.780 137.105 ;
        RECT 66.570 136.570 66.710 136.735 ;
        RECT 66.510 136.250 66.770 136.570 ;
        RECT 66.510 135.570 66.770 135.890 ;
        RECT 66.570 134.530 66.710 135.570 ;
        RECT 66.510 134.210 66.770 134.530 ;
        RECT 66.040 131.975 66.320 132.345 ;
        RECT 65.650 131.240 66.710 131.380 ;
        RECT 64.670 130.900 65.330 131.040 ;
        RECT 64.670 130.810 64.930 130.900 ;
        RECT 64.210 130.130 64.470 130.450 ;
        RECT 64.270 128.750 64.410 130.130 ;
        RECT 64.210 128.430 64.470 128.750 ;
        RECT 63.750 127.410 64.010 127.730 ;
        RECT 63.810 126.370 63.950 127.410 ;
        RECT 63.290 126.225 63.550 126.370 ;
        RECT 63.280 125.855 63.560 126.225 ;
        RECT 63.750 126.050 64.010 126.370 ;
        RECT 64.270 126.030 64.410 128.430 ;
        RECT 64.210 125.710 64.470 126.030 ;
        RECT 63.740 125.175 64.020 125.545 ;
        RECT 63.810 123.990 63.950 125.175 ;
        RECT 64.210 124.690 64.470 125.010 ;
        RECT 63.750 123.670 64.010 123.990 ;
        RECT 62.830 122.990 63.090 123.310 ;
        RECT 63.750 122.990 64.010 123.310 ;
        RECT 63.810 122.825 63.950 122.990 ;
        RECT 62.430 122.570 63.030 122.710 ;
        RECT 62.370 121.970 62.630 122.290 ;
        RECT 62.430 120.930 62.570 121.970 ;
        RECT 62.890 121.270 63.030 122.570 ;
        RECT 63.740 122.455 64.020 122.825 ;
        RECT 63.740 121.775 64.020 122.145 ;
        RECT 62.830 120.950 63.090 121.270 ;
        RECT 62.370 120.610 62.630 120.930 ;
        RECT 63.290 120.610 63.550 120.930 ;
        RECT 62.830 120.270 63.090 120.590 ;
        RECT 61.910 119.930 62.170 120.250 ;
        RECT 60.530 119.590 60.790 119.910 ;
        RECT 61.970 118.310 62.110 119.930 ;
        RECT 61.510 118.170 62.110 118.310 ;
        RECT 60.530 117.550 60.790 117.870 ;
        RECT 60.990 117.550 61.250 117.870 ;
        RECT 59.610 116.870 59.870 117.190 ;
        RECT 59.670 113.110 59.810 116.870 ;
        RECT 60.590 116.850 60.730 117.550 ;
        RECT 60.530 116.530 60.790 116.850 ;
        RECT 60.590 115.150 60.730 116.530 ;
        RECT 60.530 114.830 60.790 115.150 ;
        RECT 59.610 112.790 59.870 113.110 ;
        RECT 58.750 112.370 59.350 112.510 ;
        RECT 58.230 107.350 58.490 107.670 ;
        RECT 58.290 103.930 58.430 107.350 ;
        RECT 58.230 103.610 58.490 103.930 ;
        RECT 58.750 102.230 58.890 112.370 ;
        RECT 59.670 109.710 59.810 112.790 ;
        RECT 60.070 111.770 60.330 112.090 ;
        RECT 60.530 111.770 60.790 112.090 ;
        RECT 59.610 109.390 59.870 109.710 ;
        RECT 59.150 109.050 59.410 109.370 ;
        RECT 59.210 106.650 59.350 109.050 ;
        RECT 60.130 108.690 60.270 111.770 ;
        RECT 60.590 109.710 60.730 111.770 ;
        RECT 60.530 109.390 60.790 109.710 ;
        RECT 60.070 108.370 60.330 108.690 ;
        RECT 59.610 106.670 59.870 106.990 ;
        RECT 59.150 106.330 59.410 106.650 ;
        RECT 59.210 104.270 59.350 106.330 ;
        RECT 59.150 103.950 59.410 104.270 ;
        RECT 59.670 103.250 59.810 106.670 ;
        RECT 59.610 102.930 59.870 103.250 ;
        RECT 58.690 101.910 58.950 102.230 ;
        RECT 57.770 101.230 58.030 101.550 ;
        RECT 57.310 99.190 57.570 99.510 ;
        RECT 57.830 97.665 57.970 101.230 ;
        RECT 58.230 100.210 58.490 100.530 ;
        RECT 58.290 99.170 58.430 100.210 ;
        RECT 59.670 99.510 59.810 102.930 ;
        RECT 60.530 101.910 60.790 102.230 ;
        RECT 59.610 99.190 59.870 99.510 ;
        RECT 58.230 98.850 58.490 99.170 ;
        RECT 60.590 98.830 60.730 101.910 ;
        RECT 60.530 98.510 60.790 98.830 ;
        RECT 57.760 97.295 58.040 97.665 ;
        RECT 55.470 95.450 55.730 95.770 ;
        RECT 55.530 94.945 55.670 95.450 ;
        RECT 55.460 94.575 55.740 94.945 ;
        RECT 61.050 94.070 61.190 117.550 ;
        RECT 61.510 96.790 61.650 118.170 ;
        RECT 62.890 117.870 63.030 120.270 ;
        RECT 62.830 117.550 63.090 117.870 ;
        RECT 63.350 107.185 63.490 120.610 ;
        RECT 63.810 115.230 63.950 121.775 ;
        RECT 64.270 120.930 64.410 124.690 ;
        RECT 64.210 120.610 64.470 120.930 ;
        RECT 64.200 119.735 64.480 120.105 ;
        RECT 64.270 117.190 64.410 119.735 ;
        RECT 64.210 116.870 64.470 117.190 ;
        RECT 63.810 115.090 64.410 115.230 ;
        RECT 63.750 114.490 64.010 114.810 ;
        RECT 63.810 112.770 63.950 114.490 ;
        RECT 63.750 112.450 64.010 112.770 ;
        RECT 63.280 106.815 63.560 107.185 ;
        RECT 63.810 106.990 63.950 112.450 ;
        RECT 64.270 107.750 64.410 115.090 ;
        RECT 64.730 114.810 64.870 130.810 ;
        RECT 66.050 130.470 66.310 130.790 ;
        RECT 65.130 130.130 65.390 130.450 ;
        RECT 65.190 126.710 65.330 130.130 ;
        RECT 66.110 129.340 66.250 130.470 ;
        RECT 65.650 129.200 66.250 129.340 ;
        RECT 65.130 126.390 65.390 126.710 ;
        RECT 65.650 125.010 65.790 129.200 ;
        RECT 66.570 128.750 66.710 131.240 ;
        RECT 66.050 128.430 66.310 128.750 ;
        RECT 66.510 128.430 66.770 128.750 ;
        RECT 66.110 126.225 66.250 128.430 ;
        RECT 66.040 125.855 66.320 126.225 ;
        RECT 65.120 124.495 65.400 124.865 ;
        RECT 65.590 124.690 65.850 125.010 ;
        RECT 65.190 123.310 65.330 124.495 ;
        RECT 65.130 122.990 65.390 123.310 ;
        RECT 65.130 121.970 65.390 122.290 ;
        RECT 65.190 121.270 65.330 121.970 ;
        RECT 65.130 120.950 65.390 121.270 ;
        RECT 65.190 119.570 65.330 120.950 ;
        RECT 65.130 119.250 65.390 119.570 ;
        RECT 64.670 114.720 64.930 114.810 ;
        RECT 64.670 114.580 65.330 114.720 ;
        RECT 64.670 114.490 64.930 114.580 ;
        RECT 64.670 113.810 64.930 114.130 ;
        RECT 64.730 112.430 64.870 113.810 ;
        RECT 65.190 112.430 65.330 114.580 ;
        RECT 65.650 113.190 65.790 124.690 ;
        RECT 66.040 123.815 66.320 124.185 ;
        RECT 66.570 123.990 66.710 128.430 ;
        RECT 67.030 126.370 67.170 143.730 ;
        RECT 67.490 142.690 67.630 148.150 ;
        RECT 67.950 144.730 68.090 149.850 ;
        RECT 67.890 144.410 68.150 144.730 ;
        RECT 67.880 142.855 68.160 143.225 ;
        RECT 67.430 142.370 67.690 142.690 ;
        RECT 67.950 142.350 68.090 142.855 ;
        RECT 67.890 142.030 68.150 142.350 ;
        RECT 67.430 141.350 67.690 141.670 ;
        RECT 67.490 139.970 67.630 141.350 ;
        RECT 67.950 140.310 68.090 142.030 ;
        RECT 68.410 142.010 68.550 154.270 ;
        RECT 71.170 153.230 71.310 159.010 ;
        RECT 74.390 158.750 74.530 159.010 ;
        RECT 74.850 158.750 74.990 159.290 ;
        RECT 74.390 158.610 74.990 158.750 ;
        RECT 72.490 153.590 72.750 153.910 ;
        RECT 71.110 152.910 71.370 153.230 ;
        RECT 71.100 151.015 71.380 151.385 ;
        RECT 71.170 150.170 71.310 151.015 ;
        RECT 72.550 150.510 72.690 153.590 ;
        RECT 75.700 152.375 75.980 152.745 ;
        RECT 72.840 151.355 74.380 151.725 ;
        RECT 74.780 151.100 75.060 151.385 ;
        RECT 73.470 151.015 75.060 151.100 ;
        RECT 73.470 150.960 74.990 151.015 ;
        RECT 72.950 150.530 73.210 150.850 ;
        RECT 72.490 150.190 72.750 150.510 ;
        RECT 69.730 150.025 69.990 150.170 ;
        RECT 68.810 149.510 69.070 149.830 ;
        RECT 69.720 149.655 70.000 150.025 ;
        RECT 71.110 149.850 71.370 150.170 ;
        RECT 71.570 149.510 71.830 149.830 ;
        RECT 68.870 148.380 69.010 149.510 ;
        RECT 69.540 148.635 71.080 149.005 ;
        RECT 68.870 148.240 70.850 148.380 ;
        RECT 70.190 147.470 70.450 147.790 ;
        RECT 69.730 147.130 69.990 147.450 ;
        RECT 68.810 146.450 69.070 146.770 ;
        RECT 68.870 142.545 69.010 146.450 ;
        RECT 69.270 144.750 69.530 145.070 ;
        RECT 69.330 144.390 69.470 144.750 ;
        RECT 69.790 144.585 69.930 147.130 ;
        RECT 70.250 145.410 70.390 147.470 ;
        RECT 70.710 145.410 70.850 148.240 ;
        RECT 71.110 148.150 71.370 148.470 ;
        RECT 71.170 146.770 71.310 148.150 ;
        RECT 71.110 146.450 71.370 146.770 ;
        RECT 70.190 145.090 70.450 145.410 ;
        RECT 70.650 145.090 70.910 145.410 ;
        RECT 69.270 144.070 69.530 144.390 ;
        RECT 69.720 144.215 70.000 144.585 ;
        RECT 69.540 143.195 71.080 143.565 ;
        RECT 68.800 142.175 69.080 142.545 ;
        RECT 69.270 142.370 69.530 142.690 ;
        RECT 68.350 141.690 68.610 142.010 ;
        RECT 68.350 141.240 68.610 141.330 ;
        RECT 69.330 141.240 69.470 142.370 ;
        RECT 69.720 142.175 70.000 142.545 ;
        RECT 69.790 142.010 69.930 142.175 ;
        RECT 69.730 141.690 69.990 142.010 ;
        RECT 70.190 141.690 70.450 142.010 ;
        RECT 71.630 141.865 71.770 149.510 ;
        RECT 73.010 148.550 73.150 150.530 ;
        RECT 73.470 150.025 73.610 150.960 ;
        RECT 75.770 150.510 75.910 152.375 ;
        RECT 73.870 150.190 74.130 150.510 ;
        RECT 74.330 150.190 74.590 150.510 ;
        RECT 75.710 150.190 75.970 150.510 ;
        RECT 73.400 149.655 73.680 150.025 ;
        RECT 73.930 149.345 74.070 150.190 ;
        RECT 74.390 150.025 74.530 150.190 ;
        RECT 74.320 149.655 74.600 150.025 ;
        RECT 74.790 149.850 75.050 150.170 ;
        RECT 73.860 148.975 74.140 149.345 ;
        RECT 73.010 148.410 74.070 148.550 ;
        RECT 72.090 147.560 73.150 147.700 ;
        RECT 73.400 147.615 73.680 147.985 ;
        RECT 72.090 145.945 72.230 147.560 ;
        RECT 72.490 146.790 72.750 147.110 ;
        RECT 72.020 145.575 72.300 145.945 ;
        RECT 72.030 144.410 72.290 144.730 ;
        RECT 72.090 143.225 72.230 144.410 ;
        RECT 72.550 143.905 72.690 146.790 ;
        RECT 73.010 146.680 73.150 147.560 ;
        RECT 73.470 147.450 73.610 147.615 ;
        RECT 73.930 147.450 74.070 148.410 ;
        RECT 74.850 147.790 74.990 149.850 ;
        RECT 75.250 149.170 75.510 149.490 ;
        RECT 74.790 147.470 75.050 147.790 ;
        RECT 73.410 147.130 73.670 147.450 ;
        RECT 73.870 147.130 74.130 147.450 ;
        RECT 73.010 146.540 74.990 146.680 ;
        RECT 75.310 146.625 75.450 149.170 ;
        RECT 75.770 147.450 75.910 150.190 ;
        RECT 75.710 147.130 75.970 147.450 ;
        RECT 72.840 145.915 74.380 146.285 ;
        RECT 74.850 145.945 74.990 146.540 ;
        RECT 75.240 146.255 75.520 146.625 ;
        RECT 74.780 145.575 75.060 145.945 ;
        RECT 72.950 144.750 73.210 145.070 ;
        RECT 73.010 144.050 73.150 144.750 ;
        RECT 73.410 144.410 73.670 144.730 ;
        RECT 72.480 143.535 72.760 143.905 ;
        RECT 72.950 143.730 73.210 144.050 ;
        RECT 72.020 142.855 72.300 143.225 ;
        RECT 73.470 143.030 73.610 144.410 ;
        RECT 74.790 144.070 75.050 144.390 ;
        RECT 75.250 144.070 75.510 144.390 ;
        RECT 73.410 142.710 73.670 143.030 ;
        RECT 73.870 142.710 74.130 143.030 ;
        RECT 74.320 142.855 74.600 143.225 ;
        RECT 73.930 142.260 74.070 142.710 ;
        RECT 72.090 142.120 74.070 142.260 ;
        RECT 68.350 141.100 69.470 141.240 ;
        RECT 68.350 141.010 68.610 141.100 ;
        RECT 69.730 141.010 69.990 141.330 ;
        RECT 69.790 140.390 69.930 141.010 ;
        RECT 70.250 140.505 70.390 141.690 ;
        RECT 71.560 141.495 71.840 141.865 ;
        RECT 72.090 141.185 72.230 142.120 ;
        RECT 74.390 141.670 74.530 142.855 ;
        RECT 74.850 141.670 74.990 144.070 ;
        RECT 74.330 141.350 74.590 141.670 ;
        RECT 74.790 141.350 75.050 141.670 ;
        RECT 72.020 140.815 72.300 141.185 ;
        RECT 67.890 139.990 68.150 140.310 ;
        RECT 69.330 140.250 69.930 140.390 ;
        RECT 69.330 140.220 69.470 140.250 ;
        RECT 68.870 140.080 69.470 140.220 ;
        RECT 70.180 140.135 70.460 140.505 ;
        RECT 72.840 140.475 74.380 140.845 ;
        RECT 67.430 139.825 67.690 139.970 ;
        RECT 67.420 139.455 67.700 139.825 ;
        RECT 67.430 138.970 67.690 139.290 ;
        RECT 67.490 137.250 67.630 138.970 ;
        RECT 68.870 138.860 69.010 140.080 ;
        RECT 71.570 139.990 71.830 140.310 ;
        RECT 74.780 140.135 75.060 140.505 ;
        RECT 75.310 140.310 75.450 144.070 ;
        RECT 75.710 142.710 75.970 143.030 ;
        RECT 75.770 141.185 75.910 142.710 ;
        RECT 75.700 140.815 75.980 141.185 ;
        RECT 69.260 139.455 69.540 139.825 ;
        RECT 69.270 139.310 69.530 139.455 ;
        RECT 70.190 139.310 70.450 139.630 ;
        RECT 68.315 138.720 69.010 138.860 ;
        RECT 67.890 138.290 68.150 138.610 ;
        RECT 67.430 136.930 67.690 137.250 ;
        RECT 67.420 136.055 67.700 136.425 ;
        RECT 67.490 134.190 67.630 136.055 ;
        RECT 67.950 134.190 68.090 138.290 ;
        RECT 68.315 137.670 68.455 138.720 ;
        RECT 70.250 138.520 70.390 139.310 ;
        RECT 71.630 138.520 71.770 139.990 ;
        RECT 74.330 139.880 74.590 139.970 ;
        RECT 73.930 139.740 74.590 139.880 ;
        RECT 72.950 139.310 73.210 139.630 ;
        RECT 70.250 138.380 71.770 138.520 ;
        RECT 69.540 137.755 71.080 138.125 ;
        RECT 68.315 137.530 68.550 137.670 ;
        RECT 67.430 133.870 67.690 134.190 ;
        RECT 67.890 133.870 68.150 134.190 ;
        RECT 67.420 133.335 67.700 133.705 ;
        RECT 67.890 133.420 68.150 133.510 ;
        RECT 68.410 133.420 68.550 137.530 ;
        RECT 69.270 137.160 69.530 137.250 ;
        RECT 69.270 137.020 70.390 137.160 ;
        RECT 69.270 136.930 69.530 137.020 ;
        RECT 69.270 136.250 69.530 136.570 ;
        RECT 69.330 135.890 69.470 136.250 ;
        RECT 69.270 135.570 69.530 135.890 ;
        RECT 69.730 135.570 69.990 135.890 ;
        RECT 69.330 134.385 69.470 135.570 ;
        RECT 69.790 135.065 69.930 135.570 ;
        RECT 69.720 134.695 70.000 135.065 ;
        RECT 69.730 134.440 69.990 134.530 ;
        RECT 70.250 134.440 70.390 137.020 ;
        RECT 71.110 136.480 71.370 136.570 ;
        RECT 71.630 136.480 71.770 138.380 ;
        RECT 72.020 137.415 72.300 137.785 ;
        RECT 72.090 137.250 72.230 137.415 ;
        RECT 72.030 136.930 72.290 137.250 ;
        RECT 72.490 136.480 72.750 136.570 ;
        RECT 71.110 136.340 71.770 136.480 ;
        RECT 72.090 136.340 72.750 136.480 ;
        RECT 71.110 136.250 71.370 136.340 ;
        RECT 69.260 134.015 69.540 134.385 ;
        RECT 69.730 134.300 70.390 134.440 ;
        RECT 69.730 134.210 69.990 134.300 ;
        RECT 71.170 133.705 71.310 136.250 ;
        RECT 72.090 134.190 72.230 136.340 ;
        RECT 72.490 136.250 72.750 136.340 ;
        RECT 73.010 135.800 73.150 139.310 ;
        RECT 73.930 135.890 74.070 139.740 ;
        RECT 74.330 139.650 74.590 139.740 ;
        RECT 74.850 139.630 74.990 140.135 ;
        RECT 75.250 139.990 75.510 140.310 ;
        RECT 74.790 139.310 75.050 139.630 ;
        RECT 74.330 138.290 74.590 138.610 ;
        RECT 72.550 135.660 73.150 135.800 ;
        RECT 71.570 133.870 71.830 134.190 ;
        RECT 72.030 133.870 72.290 134.190 ;
        RECT 67.490 131.470 67.630 133.335 ;
        RECT 67.890 133.280 68.550 133.420 ;
        RECT 71.100 133.335 71.380 133.705 ;
        RECT 67.890 133.190 68.150 133.280 ;
        RECT 67.430 131.150 67.690 131.470 ;
        RECT 67.950 129.625 68.090 133.190 ;
        RECT 68.800 132.655 69.080 133.025 ;
        RECT 68.340 131.975 68.620 132.345 ;
        RECT 67.880 129.255 68.160 129.625 ;
        RECT 68.410 129.000 68.550 131.975 ;
        RECT 67.490 128.860 68.550 129.000 ;
        RECT 66.970 126.050 67.230 126.370 ;
        RECT 66.050 123.670 66.310 123.815 ;
        RECT 66.510 123.670 66.770 123.990 ;
        RECT 66.570 120.590 66.710 123.670 ;
        RECT 67.490 123.650 67.630 128.860 ;
        RECT 67.880 127.895 68.160 128.265 ;
        RECT 68.350 128.090 68.610 128.410 ;
        RECT 67.950 127.730 68.090 127.895 ;
        RECT 67.890 127.410 68.150 127.730 ;
        RECT 67.880 126.535 68.160 126.905 ;
        RECT 67.890 126.390 68.150 126.535 ;
        RECT 67.890 125.600 68.150 125.690 ;
        RECT 68.410 125.600 68.550 128.090 ;
        RECT 67.890 125.460 68.550 125.600 ;
        RECT 67.890 125.370 68.150 125.460 ;
        RECT 68.350 124.690 68.610 125.010 ;
        RECT 68.410 124.185 68.550 124.690 ;
        RECT 68.340 123.815 68.620 124.185 ;
        RECT 67.430 123.330 67.690 123.650 ;
        RECT 68.870 123.310 69.010 132.655 ;
        RECT 69.540 132.315 71.080 132.685 ;
        RECT 69.270 131.150 69.530 131.470 ;
        RECT 70.650 131.150 70.910 131.470 ;
        RECT 69.330 128.750 69.470 131.150 ;
        RECT 69.720 130.615 70.000 130.985 ;
        RECT 69.270 128.430 69.530 128.750 ;
        RECT 69.790 127.730 69.930 130.615 ;
        RECT 70.190 130.305 70.450 130.450 ;
        RECT 70.180 129.935 70.460 130.305 ;
        RECT 70.710 128.750 70.850 131.150 ;
        RECT 71.630 130.450 71.770 133.870 ;
        RECT 72.030 133.190 72.290 133.510 ;
        RECT 72.090 131.470 72.230 133.190 ;
        RECT 72.030 131.150 72.290 131.470 ;
        RECT 71.110 130.130 71.370 130.450 ;
        RECT 71.570 130.130 71.830 130.450 ;
        RECT 71.170 129.625 71.310 130.130 ;
        RECT 71.100 129.255 71.380 129.625 ;
        RECT 70.650 128.430 70.910 128.750 ;
        RECT 69.730 127.410 69.990 127.730 ;
        RECT 71.630 127.640 71.770 130.130 ;
        RECT 72.020 129.255 72.300 129.625 ;
        RECT 72.550 129.340 72.690 135.660 ;
        RECT 73.870 135.570 74.130 135.890 ;
        RECT 74.390 135.800 74.530 138.290 ;
        RECT 74.850 137.250 74.990 139.310 ;
        RECT 75.310 137.785 75.450 139.990 ;
        RECT 75.710 138.630 75.970 138.950 ;
        RECT 75.240 137.415 75.520 137.785 ;
        RECT 74.790 136.930 75.050 137.250 ;
        RECT 75.770 136.570 75.910 138.630 ;
        RECT 74.790 136.310 75.050 136.570 ;
        RECT 75.710 136.425 75.970 136.570 ;
        RECT 74.790 136.250 75.450 136.310 ;
        RECT 74.850 136.170 75.450 136.250 ;
        RECT 74.390 135.660 74.990 135.800 ;
        RECT 72.840 135.035 74.380 135.405 ;
        RECT 72.950 134.550 73.210 134.870 ;
        RECT 73.010 133.510 73.150 134.550 ;
        RECT 73.410 133.870 73.670 134.190 ;
        RECT 72.950 133.190 73.210 133.510 ;
        RECT 73.470 133.025 73.610 133.870 ;
        RECT 73.870 133.530 74.130 133.850 ;
        RECT 73.400 132.655 73.680 133.025 ;
        RECT 73.400 131.975 73.680 132.345 ;
        RECT 73.470 131.810 73.610 131.975 ;
        RECT 72.940 131.295 73.220 131.665 ;
        RECT 73.410 131.490 73.670 131.810 ;
        RECT 73.010 131.130 73.150 131.295 ;
        RECT 72.950 130.810 73.210 131.130 ;
        RECT 73.930 130.985 74.070 133.530 ;
        RECT 74.330 132.850 74.590 133.170 ;
        RECT 74.390 131.040 74.530 132.850 ;
        RECT 74.850 131.810 74.990 135.660 ;
        RECT 75.310 133.850 75.450 136.170 ;
        RECT 75.700 136.055 75.980 136.425 ;
        RECT 75.710 135.570 75.970 135.890 ;
        RECT 75.770 134.530 75.910 135.570 ;
        RECT 75.710 134.210 75.970 134.530 ;
        RECT 75.250 133.705 75.510 133.850 ;
        RECT 75.240 133.335 75.520 133.705 ;
        RECT 74.790 131.490 75.050 131.810 ;
        RECT 75.250 131.490 75.510 131.810 ;
        RECT 73.860 130.615 74.140 130.985 ;
        RECT 74.390 130.900 74.990 131.040 ;
        RECT 72.840 129.595 74.380 129.965 ;
        RECT 72.090 128.150 72.230 129.255 ;
        RECT 72.550 129.200 73.150 129.340 ;
        RECT 72.090 128.010 72.690 128.150 ;
        RECT 71.630 127.500 72.230 127.640 ;
        RECT 69.540 126.875 71.080 127.245 ;
        RECT 69.270 126.390 69.530 126.710 ;
        RECT 71.110 126.390 71.370 126.710 ;
        RECT 69.330 126.225 69.470 126.390 ;
        RECT 69.260 125.855 69.540 126.225 ;
        RECT 70.180 125.855 70.460 126.225 ;
        RECT 70.250 125.690 70.390 125.855 ;
        RECT 69.720 125.175 70.000 125.545 ;
        RECT 70.190 125.370 70.450 125.690 ;
        RECT 69.790 123.650 69.930 125.175 ;
        RECT 71.170 123.990 71.310 126.390 ;
        RECT 71.570 125.030 71.830 125.350 ;
        RECT 71.630 124.865 71.770 125.030 ;
        RECT 71.560 124.495 71.840 124.865 ;
        RECT 71.110 123.670 71.370 123.990 ;
        RECT 69.730 123.330 69.990 123.650 ;
        RECT 68.810 122.990 69.070 123.310 ;
        RECT 67.880 122.540 68.160 122.825 ;
        RECT 68.350 122.540 68.610 122.630 ;
        RECT 67.880 122.455 68.610 122.540 ;
        RECT 68.800 122.455 69.080 122.825 ;
        RECT 67.950 122.400 68.610 122.455 ;
        RECT 66.510 120.270 66.770 120.590 ;
        RECT 67.430 114.490 67.690 114.810 ;
        RECT 66.510 113.810 66.770 114.130 ;
        RECT 65.650 113.050 66.250 113.190 ;
        RECT 66.570 113.110 66.710 113.810 ;
        RECT 67.490 113.110 67.630 114.490 ;
        RECT 64.670 112.110 64.930 112.430 ;
        RECT 65.130 112.340 65.390 112.430 ;
        RECT 65.130 112.200 65.790 112.340 ;
        RECT 65.130 112.110 65.390 112.200 ;
        RECT 65.650 109.370 65.790 112.200 ;
        RECT 65.130 109.050 65.390 109.370 ;
        RECT 65.590 109.050 65.850 109.370 ;
        RECT 64.270 107.610 64.870 107.750 ;
        RECT 65.190 107.670 65.330 109.050 ;
        RECT 63.750 106.670 64.010 106.990 ;
        RECT 64.210 106.670 64.470 106.990 ;
        RECT 63.810 104.950 63.950 106.670 ;
        RECT 63.750 104.630 64.010 104.950 ;
        RECT 64.270 103.250 64.410 106.670 ;
        RECT 64.210 102.930 64.470 103.250 ;
        RECT 62.370 99.190 62.630 99.510 ;
        RECT 62.430 98.150 62.570 99.190 ;
        RECT 63.290 98.850 63.550 99.170 ;
        RECT 63.350 98.490 63.490 98.850 ;
        RECT 63.290 98.170 63.550 98.490 ;
        RECT 62.370 97.830 62.630 98.150 ;
        RECT 61.450 96.470 61.710 96.790 ;
        RECT 61.510 94.070 61.650 96.470 ;
        RECT 62.430 95.430 62.570 97.830 ;
        RECT 63.350 95.770 63.490 98.170 ;
        RECT 62.830 95.450 63.090 95.770 ;
        RECT 63.290 95.450 63.550 95.770 ;
        RECT 62.370 95.110 62.630 95.430 ;
        RECT 60.990 93.750 61.250 94.070 ;
        RECT 61.450 93.750 61.710 94.070 ;
        RECT 57.310 92.390 57.570 92.710 ;
        RECT 57.370 90.670 57.510 92.390 ;
        RECT 57.310 90.350 57.570 90.670 ;
        RECT 61.050 90.330 61.190 93.750 ;
        RECT 61.510 93.050 61.650 93.750 ;
        RECT 62.430 93.730 62.570 95.110 ;
        RECT 62.890 93.730 63.030 95.450 ;
        RECT 62.370 93.410 62.630 93.730 ;
        RECT 62.830 93.410 63.090 93.730 ;
        RECT 61.450 92.730 61.710 93.050 ;
        RECT 63.350 92.710 63.490 95.450 ;
        RECT 63.290 92.390 63.550 92.710 ;
        RECT 55.920 89.815 56.200 90.185 ;
        RECT 60.990 90.010 61.250 90.330 ;
        RECT 55.930 89.670 56.190 89.815 ;
        RECT 64.730 85.230 64.870 107.610 ;
        RECT 65.130 107.350 65.390 107.670 ;
        RECT 66.110 105.970 66.250 113.050 ;
        RECT 66.510 112.790 66.770 113.110 ;
        RECT 67.430 112.790 67.690 113.110 ;
        RECT 67.430 112.110 67.690 112.430 ;
        RECT 67.490 110.050 67.630 112.110 ;
        RECT 66.970 109.905 67.230 110.050 ;
        RECT 66.960 109.535 67.240 109.905 ;
        RECT 67.430 109.730 67.690 110.050 ;
        RECT 67.490 109.370 67.630 109.730 ;
        RECT 67.430 109.050 67.690 109.370 ;
        RECT 66.050 105.650 66.310 105.970 ;
        RECT 67.950 104.180 68.090 122.400 ;
        RECT 68.350 122.310 68.610 122.400 ;
        RECT 68.870 121.270 69.010 122.455 ;
        RECT 69.540 121.435 71.080 121.805 ;
        RECT 68.810 120.950 69.070 121.270 ;
        RECT 69.270 119.930 69.530 120.250 ;
        RECT 69.730 119.930 69.990 120.250 ;
        RECT 70.190 119.930 70.450 120.250 ;
        RECT 69.330 118.550 69.470 119.930 ;
        RECT 69.270 118.230 69.530 118.550 ;
        RECT 69.790 117.530 69.930 119.930 ;
        RECT 70.250 117.870 70.390 119.930 ;
        RECT 71.110 119.590 71.370 119.910 ;
        RECT 70.190 117.550 70.450 117.870 ;
        RECT 69.730 117.210 69.990 117.530 ;
        RECT 71.170 117.440 71.310 119.590 ;
        RECT 71.630 118.210 71.770 124.495 ;
        RECT 72.090 123.990 72.230 127.500 ;
        RECT 72.550 125.010 72.690 128.010 ;
        RECT 73.010 125.010 73.150 129.200 ;
        RECT 73.870 129.110 74.130 129.430 ;
        RECT 73.410 128.430 73.670 128.750 ;
        RECT 73.470 126.710 73.610 128.430 ;
        RECT 73.930 126.710 74.070 129.110 ;
        RECT 73.410 126.390 73.670 126.710 ;
        RECT 73.870 126.390 74.130 126.710 ;
        RECT 73.860 125.855 74.140 126.225 ;
        RECT 73.930 125.690 74.070 125.855 ;
        RECT 73.870 125.370 74.130 125.690 ;
        RECT 72.490 124.690 72.750 125.010 ;
        RECT 72.950 124.690 73.210 125.010 ;
        RECT 72.030 123.670 72.290 123.990 ;
        RECT 72.030 122.650 72.290 122.970 ;
        RECT 71.570 117.890 71.830 118.210 ;
        RECT 72.090 117.530 72.230 122.650 ;
        RECT 72.550 120.930 72.690 124.690 ;
        RECT 72.840 124.155 74.380 124.525 ;
        RECT 72.950 123.670 73.210 123.990 ;
        RECT 74.850 123.900 74.990 130.900 ;
        RECT 75.310 128.070 75.450 131.490 ;
        RECT 75.770 131.130 75.910 134.210 ;
        RECT 75.710 130.810 75.970 131.130 ;
        RECT 75.700 128.575 75.980 128.945 ;
        RECT 75.250 127.750 75.510 128.070 ;
        RECT 75.310 126.030 75.450 127.750 ;
        RECT 75.250 125.710 75.510 126.030 ;
        RECT 75.770 125.430 75.910 128.575 ;
        RECT 76.230 126.710 76.370 159.290 ;
        RECT 77.540 159.010 77.820 163.010 ;
        RECT 80.760 159.010 81.040 163.010 ;
        RECT 83.980 159.010 84.260 163.010 ;
        RECT 87.200 159.010 87.480 163.010 ;
        RECT 90.420 159.010 90.700 163.010 ;
        RECT 93.640 159.010 93.920 163.010 ;
        RECT 96.860 159.010 97.140 163.010 ;
        RECT 100.080 159.010 100.360 163.010 ;
        RECT 103.300 159.010 103.580 163.010 ;
        RECT 106.520 159.010 106.800 163.010 ;
        RECT 107.050 159.290 108.570 159.430 ;
        RECT 77.610 155.950 77.750 159.010 ;
        RECT 77.550 155.630 77.810 155.950 ;
        RECT 78.010 152.910 78.270 153.230 ;
        RECT 77.550 151.890 77.810 152.210 ;
        RECT 77.610 150.510 77.750 151.890 ;
        RECT 77.550 150.190 77.810 150.510 ;
        RECT 77.090 149.850 77.350 150.170 ;
        RECT 76.630 149.170 76.890 149.490 ;
        RECT 76.690 140.310 76.830 149.170 ;
        RECT 77.150 144.050 77.290 149.850 ;
        RECT 77.550 146.790 77.810 147.110 ;
        RECT 77.090 143.730 77.350 144.050 ;
        RECT 77.610 143.110 77.750 146.790 ;
        RECT 77.150 142.970 77.750 143.110 ;
        RECT 77.150 140.310 77.290 142.970 ;
        RECT 77.550 141.010 77.810 141.330 ;
        RECT 76.630 139.990 76.890 140.310 ;
        RECT 77.090 139.990 77.350 140.310 ;
        RECT 77.610 139.630 77.750 141.010 ;
        RECT 77.090 139.310 77.350 139.630 ;
        RECT 77.550 139.310 77.810 139.630 ;
        RECT 76.630 138.970 76.890 139.290 ;
        RECT 76.690 137.785 76.830 138.970 ;
        RECT 76.620 137.415 76.900 137.785 ;
        RECT 76.630 135.910 76.890 136.230 ;
        RECT 76.170 126.390 76.430 126.710 ;
        RECT 73.930 123.760 74.990 123.900 ;
        RECT 75.310 125.290 75.910 125.430 ;
        RECT 72.490 120.610 72.750 120.930 ;
        RECT 73.010 120.160 73.150 123.670 ;
        RECT 73.400 121.095 73.680 121.465 ;
        RECT 73.470 120.250 73.610 121.095 ;
        RECT 73.930 120.250 74.070 123.760 ;
        RECT 74.780 121.095 75.060 121.465 ;
        RECT 74.850 120.250 74.990 121.095 ;
        RECT 72.550 120.020 73.150 120.160 ;
        RECT 71.170 117.300 71.770 117.440 ;
        RECT 69.540 115.995 71.080 116.365 ;
        RECT 70.190 115.170 70.450 115.490 ;
        RECT 68.340 112.430 68.620 112.625 ;
        RECT 70.250 112.430 70.390 115.170 ;
        RECT 68.255 112.255 68.620 112.430 ;
        RECT 68.255 112.200 68.550 112.255 ;
        RECT 68.255 112.110 68.515 112.200 ;
        RECT 70.190 112.110 70.450 112.430 ;
        RECT 70.250 111.410 70.390 112.110 ;
        RECT 70.190 111.090 70.450 111.410 ;
        RECT 69.540 110.555 71.080 110.925 ;
        RECT 71.630 110.390 71.770 117.300 ;
        RECT 72.030 117.210 72.290 117.530 ;
        RECT 72.090 114.810 72.230 117.210 ;
        RECT 72.030 114.490 72.290 114.810 ;
        RECT 69.270 110.070 69.530 110.390 ;
        RECT 71.570 110.070 71.830 110.390 ;
        RECT 69.330 109.370 69.470 110.070 ;
        RECT 69.270 109.050 69.530 109.370 ;
        RECT 71.570 109.050 71.830 109.370 ;
        RECT 68.810 108.710 69.070 109.030 ;
        RECT 68.340 106.815 68.620 107.185 ;
        RECT 67.030 104.040 68.090 104.180 ;
        RECT 66.510 103.610 66.770 103.930 ;
        RECT 66.570 101.890 66.710 103.610 ;
        RECT 66.510 101.570 66.770 101.890 ;
        RECT 65.130 99.190 65.390 99.510 ;
        RECT 65.190 96.450 65.330 99.190 ;
        RECT 67.030 97.810 67.170 104.040 ;
        RECT 67.890 103.270 68.150 103.590 ;
        RECT 67.950 101.550 68.090 103.270 ;
        RECT 67.430 101.230 67.690 101.550 ;
        RECT 67.890 101.230 68.150 101.550 ;
        RECT 66.970 97.490 67.230 97.810 ;
        RECT 65.130 96.130 65.390 96.450 ;
        RECT 65.590 96.130 65.850 96.450 ;
        RECT 65.130 95.110 65.390 95.430 ;
        RECT 65.190 92.710 65.330 95.110 ;
        RECT 65.130 92.390 65.390 92.710 ;
        RECT 65.650 92.370 65.790 96.130 ;
        RECT 67.490 95.770 67.630 101.230 ;
        RECT 67.950 99.510 68.090 101.230 ;
        RECT 67.890 99.190 68.150 99.510 ;
        RECT 67.430 95.450 67.690 95.770 ;
        RECT 67.890 95.450 68.150 95.770 ;
        RECT 67.950 92.710 68.090 95.450 ;
        RECT 68.410 94.070 68.550 106.815 ;
        RECT 68.870 106.650 69.010 108.710 ;
        RECT 69.330 107.670 69.470 109.050 ;
        RECT 69.270 107.350 69.530 107.670 ;
        RECT 68.810 106.330 69.070 106.650 ;
        RECT 69.540 105.115 71.080 105.485 ;
        RECT 71.630 104.950 71.770 109.050 ;
        RECT 71.570 104.630 71.830 104.950 ;
        RECT 70.650 103.610 70.910 103.930 ;
        RECT 71.570 103.840 71.830 103.930 ;
        RECT 72.090 103.840 72.230 114.490 ;
        RECT 71.570 103.700 72.230 103.840 ;
        RECT 71.570 103.610 71.830 103.700 ;
        RECT 70.710 102.230 70.850 103.610 ;
        RECT 70.650 101.910 70.910 102.230 ;
        RECT 69.540 99.675 71.080 100.045 ;
        RECT 69.540 94.235 71.080 94.605 ;
        RECT 68.350 93.750 68.610 94.070 ;
        RECT 71.630 93.980 71.770 103.610 ;
        RECT 72.030 102.930 72.290 103.250 ;
        RECT 72.090 101.550 72.230 102.930 ;
        RECT 72.030 101.230 72.290 101.550 ;
        RECT 72.550 99.170 72.690 120.020 ;
        RECT 73.410 119.930 73.670 120.250 ;
        RECT 73.870 119.930 74.130 120.250 ;
        RECT 74.790 119.930 75.050 120.250 ;
        RECT 74.790 119.250 75.050 119.570 ;
        RECT 72.840 118.715 74.380 119.085 ;
        RECT 74.850 118.745 74.990 119.250 ;
        RECT 74.780 118.375 75.060 118.745 ;
        RECT 74.850 116.850 74.990 118.375 ;
        RECT 74.790 116.530 75.050 116.850 ;
        RECT 75.310 115.490 75.450 125.290 ;
        RECT 75.710 124.690 75.970 125.010 ;
        RECT 75.770 119.570 75.910 124.690 ;
        RECT 76.690 123.310 76.830 135.910 ;
        RECT 77.150 135.890 77.290 139.310 ;
        RECT 77.540 138.775 77.820 139.145 ;
        RECT 77.610 136.910 77.750 138.775 ;
        RECT 77.550 136.590 77.810 136.910 ;
        RECT 77.090 135.570 77.350 135.890 ;
        RECT 78.070 134.100 78.210 152.910 ;
        RECT 78.470 150.190 78.730 150.510 ;
        RECT 78.530 148.130 78.670 150.190 ;
        RECT 79.840 149.655 80.120 150.025 ;
        RECT 78.920 148.975 79.200 149.345 ;
        RECT 78.470 147.810 78.730 148.130 ;
        RECT 78.470 144.585 78.730 144.730 ;
        RECT 78.460 144.215 78.740 144.585 ;
        RECT 78.460 143.110 78.740 143.225 ;
        RECT 78.990 143.110 79.130 148.975 ;
        RECT 79.390 147.130 79.650 147.450 ;
        RECT 78.460 142.970 79.130 143.110 ;
        RECT 78.460 142.855 78.740 142.970 ;
        RECT 78.530 139.290 78.670 142.855 ;
        RECT 78.470 138.970 78.730 139.290 ;
        RECT 78.930 139.145 79.190 139.290 ;
        RECT 78.920 138.775 79.200 139.145 ;
        RECT 78.470 138.290 78.730 138.610 ;
        RECT 79.450 138.520 79.590 147.130 ;
        RECT 79.910 139.630 80.050 149.655 ;
        RECT 80.310 146.450 80.570 146.770 ;
        RECT 80.370 139.630 80.510 146.450 ;
        RECT 79.850 139.310 80.110 139.630 ;
        RECT 80.310 139.310 80.570 139.630 ;
        RECT 78.990 138.380 79.590 138.520 ;
        RECT 77.150 133.960 78.210 134.100 ;
        RECT 77.150 126.905 77.290 133.960 ;
        RECT 77.550 133.420 77.810 133.510 ;
        RECT 77.550 133.280 78.210 133.420 ;
        RECT 77.550 133.190 77.810 133.280 ;
        RECT 77.550 131.830 77.810 132.150 ;
        RECT 77.610 127.730 77.750 131.830 ;
        RECT 78.070 129.340 78.210 133.280 ;
        RECT 78.530 132.150 78.670 138.290 ;
        RECT 78.990 135.745 79.130 138.380 ;
        RECT 79.390 136.250 79.650 136.570 ;
        RECT 79.910 136.425 80.050 139.310 ;
        RECT 80.300 138.775 80.580 139.145 ;
        RECT 80.370 137.590 80.510 138.775 ;
        RECT 80.310 137.270 80.570 137.590 ;
        RECT 80.310 136.590 80.570 136.910 ;
        RECT 78.920 135.375 79.200 135.745 ;
        RECT 78.930 133.870 79.190 134.190 ;
        RECT 78.470 131.830 78.730 132.150 ;
        RECT 78.990 129.625 79.130 133.870 ;
        RECT 79.450 132.150 79.590 136.250 ;
        RECT 79.840 136.055 80.120 136.425 ;
        RECT 80.370 135.890 80.510 136.590 ;
        RECT 79.850 135.570 80.110 135.890 ;
        RECT 80.310 135.570 80.570 135.890 ;
        RECT 79.910 133.170 80.050 135.570 ;
        RECT 80.310 133.530 80.570 133.850 ;
        RECT 79.850 132.850 80.110 133.170 ;
        RECT 79.390 131.830 79.650 132.150 ;
        RECT 79.390 130.810 79.650 131.130 ;
        RECT 78.070 129.200 78.670 129.340 ;
        RECT 78.920 129.255 79.200 129.625 ;
        RECT 79.450 129.430 79.590 130.810 ;
        RECT 79.840 129.935 80.120 130.305 ;
        RECT 79.910 129.430 80.050 129.935 ;
        RECT 78.010 128.430 78.270 128.750 ;
        RECT 78.070 128.265 78.210 128.430 ;
        RECT 78.000 127.895 78.280 128.265 ;
        RECT 77.550 127.410 77.810 127.730 ;
        RECT 77.080 126.535 77.360 126.905 ;
        RECT 77.090 125.370 77.350 125.690 ;
        RECT 77.550 125.370 77.810 125.690 ;
        RECT 77.150 123.990 77.290 125.370 ;
        RECT 77.090 123.670 77.350 123.990 ;
        RECT 76.630 122.990 76.890 123.310 ;
        RECT 76.690 120.670 76.830 122.990 ;
        RECT 77.080 121.095 77.360 121.465 ;
        RECT 76.230 120.530 76.830 120.670 ;
        RECT 76.230 120.250 76.370 120.530 ;
        RECT 76.170 119.930 76.430 120.250 ;
        RECT 76.630 119.930 76.890 120.250 ;
        RECT 75.710 119.480 75.970 119.570 ;
        RECT 75.710 119.340 76.370 119.480 ;
        RECT 75.710 119.250 75.970 119.340 ;
        RECT 76.230 118.550 76.370 119.340 ;
        RECT 76.170 118.230 76.430 118.550 ;
        RECT 75.710 117.550 75.970 117.870 ;
        RECT 75.250 115.170 75.510 115.490 ;
        RECT 74.790 113.810 75.050 114.130 ;
        RECT 72.840 113.275 74.380 113.645 ;
        RECT 74.850 113.110 74.990 113.810 ;
        RECT 74.790 112.790 75.050 113.110 ;
        RECT 72.950 112.110 73.210 112.430 ;
        RECT 73.010 110.390 73.150 112.110 ;
        RECT 73.410 111.090 73.670 111.410 ;
        RECT 72.950 110.070 73.210 110.390 ;
        RECT 73.470 109.225 73.610 111.090 ;
        RECT 73.870 110.070 74.130 110.390 ;
        RECT 73.400 108.855 73.680 109.225 ;
        RECT 73.930 108.690 74.070 110.070 ;
        RECT 74.850 109.710 74.990 112.790 ;
        RECT 75.240 112.255 75.520 112.625 ;
        RECT 75.310 112.090 75.450 112.255 ;
        RECT 75.250 111.770 75.510 112.090 ;
        RECT 74.790 109.390 75.050 109.710 ;
        RECT 74.780 108.855 75.060 109.225 ;
        RECT 73.870 108.370 74.130 108.690 ;
        RECT 72.840 107.835 74.380 108.205 ;
        RECT 74.850 107.330 74.990 108.855 ;
        RECT 74.790 107.010 75.050 107.330 ;
        RECT 74.850 104.860 74.990 107.010 ;
        RECT 74.390 104.720 74.990 104.860 ;
        RECT 74.390 103.590 74.530 104.720 ;
        RECT 74.790 104.180 75.050 104.270 ;
        RECT 75.310 104.180 75.450 111.770 ;
        RECT 75.770 111.410 75.910 117.550 ;
        RECT 76.230 112.090 76.370 118.230 ;
        RECT 76.690 118.065 76.830 119.930 ;
        RECT 76.620 117.695 76.900 118.065 ;
        RECT 76.630 116.530 76.890 116.850 ;
        RECT 76.170 111.770 76.430 112.090 ;
        RECT 75.710 111.090 75.970 111.410 ;
        RECT 75.710 109.390 75.970 109.710 ;
        RECT 75.770 107.670 75.910 109.390 ;
        RECT 75.710 107.350 75.970 107.670 ;
        RECT 74.790 104.040 75.450 104.180 ;
        RECT 74.790 103.950 75.050 104.040 ;
        RECT 74.330 103.270 74.590 103.590 ;
        RECT 74.790 102.930 75.050 103.250 ;
        RECT 72.840 102.395 74.380 102.765 ;
        RECT 74.850 102.230 74.990 102.930 ;
        RECT 74.790 101.910 75.050 102.230 ;
        RECT 74.330 101.230 74.590 101.550 ;
        RECT 74.390 99.170 74.530 101.230 ;
        RECT 74.790 100.890 75.050 101.210 ;
        RECT 72.490 98.850 72.750 99.170 ;
        RECT 74.330 98.850 74.590 99.170 ;
        RECT 72.490 98.170 72.750 98.490 ;
        RECT 72.030 95.790 72.290 96.110 ;
        RECT 70.710 93.840 71.770 93.980 ;
        RECT 67.890 92.390 68.150 92.710 ;
        RECT 65.590 92.050 65.850 92.370 ;
        RECT 70.710 90.240 70.850 93.840 ;
        RECT 72.090 93.730 72.230 95.790 ;
        RECT 72.030 93.410 72.290 93.730 ;
        RECT 71.570 92.730 71.830 93.050 ;
        RECT 72.030 92.730 72.290 93.050 ;
        RECT 71.110 92.050 71.370 92.370 ;
        RECT 71.170 91.010 71.310 92.050 ;
        RECT 71.630 91.010 71.770 92.730 ;
        RECT 72.090 91.350 72.230 92.730 ;
        RECT 72.030 91.030 72.290 91.350 ;
        RECT 71.110 90.690 71.370 91.010 ;
        RECT 71.570 90.690 71.830 91.010 ;
        RECT 70.710 90.100 72.230 90.240 ;
        RECT 71.570 89.330 71.830 89.650 ;
        RECT 69.540 88.795 71.080 89.165 ;
        RECT 71.630 88.630 71.770 89.330 ;
        RECT 71.570 88.310 71.830 88.630 ;
        RECT 72.090 88.030 72.230 90.100 ;
        RECT 71.630 87.890 72.230 88.030 ;
        RECT 69.730 87.290 69.990 87.610 ;
        RECT 69.790 85.570 69.930 87.290 ;
        RECT 69.730 85.250 69.990 85.570 ;
        RECT 64.670 84.910 64.930 85.230 ;
        RECT 71.630 84.890 71.770 87.890 ;
        RECT 72.030 86.950 72.290 87.270 ;
        RECT 72.090 85.910 72.230 86.950 ;
        RECT 72.030 85.590 72.290 85.910 ;
        RECT 71.570 84.570 71.830 84.890 ;
        RECT 69.540 83.355 71.080 83.725 ;
        RECT 72.550 83.190 72.690 98.170 ;
        RECT 72.840 96.955 74.380 97.325 ;
        RECT 72.950 95.790 73.210 96.110 ;
        RECT 73.010 94.070 73.150 95.790 ;
        RECT 72.950 93.750 73.210 94.070 ;
        RECT 73.010 92.370 73.150 93.750 ;
        RECT 72.950 92.050 73.210 92.370 ;
        RECT 72.840 91.515 74.380 91.885 ;
        RECT 74.850 87.950 74.990 100.890 ;
        RECT 75.310 88.630 75.450 104.040 ;
        RECT 75.770 102.310 75.910 107.350 ;
        RECT 76.230 103.930 76.370 111.770 ;
        RECT 76.690 110.050 76.830 116.530 ;
        RECT 77.150 114.040 77.290 121.095 ;
        RECT 77.610 115.830 77.750 125.370 ;
        RECT 78.530 122.825 78.670 129.200 ;
        RECT 78.990 125.690 79.130 129.255 ;
        RECT 79.390 129.110 79.650 129.430 ;
        RECT 79.850 129.110 80.110 129.430 ;
        RECT 79.390 128.090 79.650 128.410 ;
        RECT 79.450 126.710 79.590 128.090 ;
        RECT 79.850 127.750 80.110 128.070 ;
        RECT 79.390 126.390 79.650 126.710 ;
        RECT 78.930 125.370 79.190 125.690 ;
        RECT 79.910 125.600 80.050 127.750 ;
        RECT 80.370 126.370 80.510 133.530 ;
        RECT 80.830 131.810 80.970 159.010 ;
        RECT 82.140 148.295 82.420 148.665 ;
        RECT 81.230 142.030 81.490 142.350 ;
        RECT 81.290 139.630 81.430 142.030 ;
        RECT 81.690 141.010 81.950 141.330 ;
        RECT 81.230 139.310 81.490 139.630 ;
        RECT 81.230 136.250 81.490 136.570 ;
        RECT 81.290 134.870 81.430 136.250 ;
        RECT 81.230 134.550 81.490 134.870 ;
        RECT 81.230 133.870 81.490 134.190 ;
        RECT 80.770 131.490 81.030 131.810 ;
        RECT 81.290 129.340 81.430 133.870 ;
        RECT 80.830 129.200 81.430 129.340 ;
        RECT 80.310 126.050 80.570 126.370 ;
        RECT 79.380 125.175 79.660 125.545 ;
        RECT 79.910 125.460 80.510 125.600 ;
        RECT 78.460 122.455 78.740 122.825 ;
        RECT 78.000 120.415 78.280 120.785 ;
        RECT 78.070 120.250 78.210 120.415 ;
        RECT 78.010 119.930 78.270 120.250 ;
        RECT 78.930 120.105 79.190 120.250 ;
        RECT 77.550 115.510 77.810 115.830 ;
        RECT 78.070 114.810 78.210 119.930 ;
        RECT 78.470 119.590 78.730 119.910 ;
        RECT 78.920 119.735 79.200 120.105 ;
        RECT 78.530 118.210 78.670 119.590 ;
        RECT 78.470 117.890 78.730 118.210 ;
        RECT 78.010 114.490 78.270 114.810 ;
        RECT 77.150 113.900 78.210 114.040 ;
        RECT 77.090 112.110 77.350 112.430 ;
        RECT 76.630 109.730 76.890 110.050 ;
        RECT 76.170 103.610 76.430 103.930 ;
        RECT 75.770 102.170 76.370 102.310 ;
        RECT 75.710 101.570 75.970 101.890 ;
        RECT 75.770 99.510 75.910 101.570 ;
        RECT 76.230 101.210 76.370 102.170 ;
        RECT 76.170 100.890 76.430 101.210 ;
        RECT 76.690 100.870 76.830 109.730 ;
        RECT 76.630 100.550 76.890 100.870 ;
        RECT 75.710 99.190 75.970 99.510 ;
        RECT 75.710 98.510 75.970 98.830 ;
        RECT 75.770 96.110 75.910 98.510 ;
        RECT 75.710 95.790 75.970 96.110 ;
        RECT 76.620 92.535 76.900 92.905 ;
        RECT 76.630 92.390 76.890 92.535 ;
        RECT 75.710 92.050 75.970 92.370 ;
        RECT 75.250 88.310 75.510 88.630 ;
        RECT 74.790 87.630 75.050 87.950 ;
        RECT 75.770 87.610 75.910 92.050 ;
        RECT 77.150 88.630 77.290 112.110 ;
        RECT 78.070 109.280 78.210 113.900 ;
        RECT 78.990 110.390 79.130 119.735 ;
        RECT 79.450 115.150 79.590 125.175 ;
        RECT 79.850 124.865 80.110 125.010 ;
        RECT 79.840 124.495 80.120 124.865 ;
        RECT 79.850 122.990 80.110 123.310 ;
        RECT 79.910 122.630 80.050 122.990 ;
        RECT 80.370 122.825 80.510 125.460 ;
        RECT 80.830 124.185 80.970 129.200 ;
        RECT 81.230 128.660 81.490 128.750 ;
        RECT 81.750 128.660 81.890 141.010 ;
        RECT 82.210 136.425 82.350 148.295 ;
        RECT 83.070 147.130 83.330 147.450 ;
        RECT 83.130 145.410 83.270 147.130 ;
        RECT 83.530 146.790 83.790 147.110 ;
        RECT 83.070 145.090 83.330 145.410 ;
        RECT 82.600 143.535 82.880 143.905 ;
        RECT 82.670 142.690 82.810 143.535 ;
        RECT 82.610 142.370 82.870 142.690 ;
        RECT 82.610 141.350 82.870 141.670 ;
        RECT 83.070 141.350 83.330 141.670 ;
        RECT 82.140 136.055 82.420 136.425 ;
        RECT 82.670 135.890 82.810 141.350 ;
        RECT 83.130 139.825 83.270 141.350 ;
        RECT 83.060 139.455 83.340 139.825 ;
        RECT 83.070 136.930 83.330 137.250 ;
        RECT 82.150 135.570 82.410 135.890 ;
        RECT 82.610 135.570 82.870 135.890 ;
        RECT 82.210 129.430 82.350 135.570 ;
        RECT 82.670 134.530 82.810 135.570 ;
        RECT 83.130 135.065 83.270 136.930 ;
        RECT 83.590 136.570 83.730 146.790 ;
        RECT 83.530 136.250 83.790 136.570 ;
        RECT 83.060 134.695 83.340 135.065 ;
        RECT 82.610 134.210 82.870 134.530 ;
        RECT 83.530 134.210 83.790 134.530 ;
        RECT 83.070 133.870 83.330 134.190 ;
        RECT 83.130 132.110 83.270 133.870 ;
        RECT 83.590 133.510 83.730 134.210 ;
        RECT 83.530 133.190 83.790 133.510 ;
        RECT 82.670 131.970 83.270 132.110 ;
        RECT 83.520 131.975 83.800 132.345 ;
        RECT 82.670 130.790 82.810 131.970 ;
        RECT 83.070 131.490 83.330 131.810 ;
        RECT 82.610 130.470 82.870 130.790 ;
        RECT 82.150 129.110 82.410 129.430 ;
        RECT 81.230 128.520 81.890 128.660 ;
        RECT 81.230 128.430 81.490 128.520 ;
        RECT 81.230 127.410 81.490 127.730 ;
        RECT 80.760 123.815 81.040 124.185 ;
        RECT 81.290 123.650 81.430 127.410 ;
        RECT 81.680 126.535 81.960 126.905 ;
        RECT 81.230 123.330 81.490 123.650 ;
        RECT 79.850 122.310 80.110 122.630 ;
        RECT 80.300 122.455 80.580 122.825 ;
        RECT 81.750 122.630 81.890 126.535 ;
        RECT 82.210 126.370 82.350 129.110 ;
        RECT 82.670 128.945 82.810 130.470 ;
        RECT 82.600 128.575 82.880 128.945 ;
        RECT 82.610 128.090 82.870 128.410 ;
        RECT 82.150 126.050 82.410 126.370 ;
        RECT 82.670 123.900 82.810 128.090 ;
        RECT 83.130 123.990 83.270 131.490 ;
        RECT 83.590 126.225 83.730 131.975 ;
        RECT 83.520 125.855 83.800 126.225 ;
        RECT 83.530 125.380 83.790 125.700 ;
        RECT 82.210 123.760 82.810 123.900 ;
        RECT 81.690 122.310 81.950 122.630 ;
        RECT 80.310 121.970 80.570 122.290 ;
        RECT 80.770 121.970 81.030 122.290 ;
        RECT 79.850 120.610 80.110 120.930 ;
        RECT 79.910 120.250 80.050 120.610 ;
        RECT 79.850 119.930 80.110 120.250 ;
        RECT 79.390 114.830 79.650 115.150 ;
        RECT 80.370 114.130 80.510 121.970 ;
        RECT 80.830 121.270 80.970 121.970 ;
        RECT 80.770 120.950 81.030 121.270 ;
        RECT 81.230 120.270 81.490 120.590 ;
        RECT 80.770 119.930 81.030 120.250 ;
        RECT 80.830 117.530 80.970 119.930 ;
        RECT 81.290 119.570 81.430 120.270 ;
        RECT 81.230 119.250 81.490 119.570 ;
        RECT 82.210 118.630 82.350 123.760 ;
        RECT 83.070 123.670 83.330 123.990 ;
        RECT 82.610 122.990 82.870 123.310 ;
        RECT 82.670 119.990 82.810 122.990 ;
        RECT 82.670 119.850 83.270 119.990 ;
        RECT 82.610 119.250 82.870 119.570 ;
        RECT 81.750 118.490 82.350 118.630 ;
        RECT 81.750 118.310 81.890 118.490 ;
        RECT 81.750 118.170 82.350 118.310 ;
        RECT 81.690 117.780 81.950 117.870 ;
        RECT 81.290 117.640 81.950 117.780 ;
        RECT 80.770 117.210 81.030 117.530 ;
        RECT 80.310 113.810 80.570 114.130 ;
        RECT 80.370 113.110 80.510 113.810 ;
        RECT 80.310 112.790 80.570 113.110 ;
        RECT 79.390 112.110 79.650 112.430 ;
        RECT 78.930 110.070 79.190 110.390 ;
        RECT 78.470 109.905 78.730 110.050 ;
        RECT 78.460 109.535 78.740 109.905 ;
        RECT 78.930 109.280 79.190 109.370 ;
        RECT 78.070 109.140 79.190 109.280 ;
        RECT 78.930 109.050 79.190 109.140 ;
        RECT 78.470 103.950 78.730 104.270 ;
        RECT 78.530 103.160 78.670 103.950 ;
        RECT 78.990 103.670 79.130 109.050 ;
        RECT 79.450 104.950 79.590 112.110 ;
        RECT 80.370 109.790 80.510 112.790 ;
        RECT 79.910 109.710 80.510 109.790 ;
        RECT 79.850 109.650 80.510 109.710 ;
        RECT 79.850 109.390 80.110 109.650 ;
        RECT 79.910 106.990 80.050 109.390 ;
        RECT 80.310 109.050 80.570 109.370 ;
        RECT 79.850 106.670 80.110 106.990 ;
        RECT 79.390 104.630 79.650 104.950 ;
        RECT 78.990 103.530 80.050 103.670 ;
        RECT 78.530 103.020 79.130 103.160 ;
        RECT 78.990 101.550 79.130 103.020 ;
        RECT 78.470 101.230 78.730 101.550 ;
        RECT 78.930 101.230 79.190 101.550 ;
        RECT 78.530 96.790 78.670 101.230 ;
        RECT 78.990 98.490 79.130 101.230 ;
        RECT 79.380 100.695 79.660 101.065 ;
        RECT 79.390 100.550 79.650 100.695 ;
        RECT 78.930 98.170 79.190 98.490 ;
        RECT 78.470 96.470 78.730 96.790 ;
        RECT 78.530 93.050 78.670 96.470 ;
        RECT 79.910 95.090 80.050 103.530 ;
        RECT 80.370 96.790 80.510 109.050 ;
        RECT 80.310 96.470 80.570 96.790 ;
        RECT 79.850 94.770 80.110 95.090 ;
        RECT 79.910 93.050 80.050 94.770 ;
        RECT 78.470 92.730 78.730 93.050 ;
        RECT 79.850 92.730 80.110 93.050 ;
        RECT 78.010 92.050 78.270 92.370 ;
        RECT 77.090 88.310 77.350 88.630 ;
        RECT 78.070 87.610 78.210 92.050 ;
        RECT 75.710 87.290 75.970 87.610 ;
        RECT 76.170 87.290 76.430 87.610 ;
        RECT 76.630 87.290 76.890 87.610 ;
        RECT 78.010 87.290 78.270 87.610 ;
        RECT 76.230 86.930 76.370 87.290 ;
        RECT 76.170 86.610 76.430 86.930 ;
        RECT 72.840 86.075 74.380 86.445 ;
        RECT 76.230 83.190 76.370 86.610 ;
        RECT 76.690 85.570 76.830 87.290 ;
        RECT 76.630 85.250 76.890 85.570 ;
        RECT 78.470 83.890 78.730 84.210 ;
        RECT 72.490 82.870 72.750 83.190 ;
        RECT 76.170 82.870 76.430 83.190 ;
        RECT 78.530 82.510 78.670 83.890 ;
        RECT 79.910 82.850 80.050 92.730 ;
        RECT 80.830 85.230 80.970 117.210 ;
        RECT 81.290 108.690 81.430 117.640 ;
        RECT 81.690 117.550 81.950 117.640 ;
        RECT 81.690 116.870 81.950 117.190 ;
        RECT 81.230 108.370 81.490 108.690 ;
        RECT 81.290 104.950 81.430 108.370 ;
        RECT 81.230 104.630 81.490 104.950 ;
        RECT 81.750 104.350 81.890 116.870 ;
        RECT 82.210 113.110 82.350 118.170 ;
        RECT 82.670 116.850 82.810 119.250 ;
        RECT 83.130 118.550 83.270 119.850 ;
        RECT 83.070 118.230 83.330 118.550 ;
        RECT 83.060 117.695 83.340 118.065 ;
        RECT 83.070 117.550 83.330 117.695 ;
        RECT 82.610 116.530 82.870 116.850 ;
        RECT 83.130 115.910 83.270 117.550 ;
        RECT 82.670 115.770 83.270 115.910 ;
        RECT 82.150 112.790 82.410 113.110 ;
        RECT 82.670 112.625 82.810 115.770 ;
        RECT 83.060 112.935 83.340 113.305 ;
        RECT 82.600 112.255 82.880 112.625 ;
        RECT 83.130 112.430 83.270 112.935 ;
        RECT 83.070 112.110 83.330 112.430 ;
        RECT 82.610 111.770 82.870 112.090 ;
        RECT 82.670 111.410 82.810 111.770 ;
        RECT 82.150 111.090 82.410 111.410 ;
        RECT 82.610 111.090 82.870 111.410 ;
        RECT 83.130 111.265 83.270 112.110 ;
        RECT 82.210 109.370 82.350 111.090 ;
        RECT 83.060 110.895 83.340 111.265 ;
        RECT 82.610 110.070 82.870 110.390 ;
        RECT 82.150 109.050 82.410 109.370 ;
        RECT 81.290 104.210 81.890 104.350 ;
        RECT 81.290 93.050 81.430 104.210 ;
        RECT 81.690 103.610 81.950 103.930 ;
        RECT 81.750 102.230 81.890 103.610 ;
        RECT 81.690 101.910 81.950 102.230 ;
        RECT 82.150 101.910 82.410 102.230 ;
        RECT 81.690 100.890 81.950 101.210 ;
        RECT 81.750 99.510 81.890 100.890 ;
        RECT 81.690 99.190 81.950 99.510 ;
        RECT 82.210 96.110 82.350 101.910 ;
        RECT 82.150 95.790 82.410 96.110 ;
        RECT 82.670 93.050 82.810 110.070 ;
        RECT 83.060 108.855 83.340 109.225 ;
        RECT 83.070 108.710 83.330 108.855 ;
        RECT 83.590 107.670 83.730 125.380 ;
        RECT 84.050 123.990 84.190 159.010 ;
        RECT 87.270 154.105 87.410 159.010 ;
        RECT 90.490 154.250 90.630 159.010 ;
        RECT 87.200 153.735 87.480 154.105 ;
        RECT 90.430 153.930 90.690 154.250 ;
        RECT 92.260 152.375 92.540 152.745 ;
        RECT 90.890 150.190 91.150 150.510 ;
        RECT 85.830 149.510 86.090 149.830 ;
        RECT 85.370 147.810 85.630 148.130 ;
        RECT 84.910 147.130 85.170 147.450 ;
        RECT 84.450 146.450 84.710 146.770 ;
        RECT 83.990 123.670 84.250 123.990 ;
        RECT 84.510 123.310 84.650 146.450 ;
        RECT 84.970 140.310 85.110 147.130 ;
        RECT 84.910 139.990 85.170 140.310 ;
        RECT 84.900 138.095 85.180 138.465 ;
        RECT 84.970 131.130 85.110 138.095 ;
        RECT 85.430 136.910 85.570 147.810 ;
        RECT 85.890 147.450 86.030 149.510 ;
        RECT 90.430 147.810 90.690 148.130 ;
        RECT 85.830 147.130 86.090 147.450 ;
        RECT 88.590 147.130 88.850 147.450 ;
        RECT 89.050 147.130 89.310 147.450 ;
        RECT 89.970 147.130 90.230 147.450 ;
        RECT 86.290 147.020 86.550 147.110 ;
        RECT 86.290 146.880 86.950 147.020 ;
        RECT 86.290 146.790 86.550 146.880 ;
        RECT 86.290 143.730 86.550 144.050 ;
        RECT 85.830 139.310 86.090 139.630 ;
        RECT 85.890 137.590 86.030 139.310 ;
        RECT 85.830 137.270 86.090 137.590 ;
        RECT 86.350 137.250 86.490 143.730 ;
        RECT 86.290 136.930 86.550 137.250 ;
        RECT 85.370 136.590 85.630 136.910 ;
        RECT 86.280 136.055 86.560 136.425 ;
        RECT 85.830 135.570 86.090 135.890 ;
        RECT 85.360 134.015 85.640 134.385 ;
        RECT 85.890 134.190 86.030 135.570 ;
        RECT 86.350 134.870 86.490 136.055 ;
        RECT 86.290 134.550 86.550 134.870 ;
        RECT 86.350 134.190 86.490 134.550 ;
        RECT 84.910 130.810 85.170 131.130 ;
        RECT 84.900 129.255 85.180 129.625 ;
        RECT 84.910 129.110 85.170 129.255 ;
        RECT 85.430 128.945 85.570 134.015 ;
        RECT 85.830 133.870 86.090 134.190 ;
        RECT 86.290 133.870 86.550 134.190 ;
        RECT 86.290 132.850 86.550 133.170 ;
        RECT 86.350 132.150 86.490 132.850 ;
        RECT 86.290 131.830 86.550 132.150 ;
        RECT 86.350 130.870 86.490 131.830 ;
        RECT 86.810 131.810 86.950 146.880 ;
        RECT 87.210 146.790 87.470 147.110 ;
        RECT 87.270 145.070 87.410 146.790 ;
        RECT 87.210 144.750 87.470 145.070 ;
        RECT 87.670 144.750 87.930 145.070 ;
        RECT 87.270 142.690 87.410 144.750 ;
        RECT 87.210 142.370 87.470 142.690 ;
        RECT 87.730 140.505 87.870 144.750 ;
        RECT 88.120 142.175 88.400 142.545 ;
        RECT 87.660 140.135 87.940 140.505 ;
        RECT 87.670 135.910 87.930 136.230 ;
        RECT 87.730 134.530 87.870 135.910 ;
        RECT 87.670 134.210 87.930 134.530 ;
        RECT 86.750 131.490 87.010 131.810 ;
        RECT 87.210 131.490 87.470 131.810 ;
        RECT 88.190 131.550 88.330 142.175 ;
        RECT 88.650 132.150 88.790 147.130 ;
        RECT 89.110 139.970 89.250 147.130 ;
        RECT 89.510 145.090 89.770 145.410 ;
        RECT 89.570 144.730 89.710 145.090 ;
        RECT 89.510 144.410 89.770 144.730 ;
        RECT 89.510 141.350 89.770 141.670 ;
        RECT 89.050 139.650 89.310 139.970 ;
        RECT 89.040 137.415 89.320 137.785 ;
        RECT 89.110 132.175 89.250 137.415 ;
        RECT 88.590 131.830 88.850 132.150 ;
        RECT 89.040 131.805 89.320 132.175 ;
        RECT 85.890 130.730 86.490 130.870 ;
        RECT 86.750 130.810 87.010 131.130 ;
        RECT 85.360 128.575 85.640 128.945 ;
        RECT 85.890 128.750 86.030 130.730 ;
        RECT 86.290 130.130 86.550 130.450 ;
        RECT 85.370 128.430 85.630 128.575 ;
        RECT 85.830 128.430 86.090 128.750 ;
        RECT 85.430 125.545 85.570 128.430 ;
        RECT 85.830 127.750 86.090 128.070 ;
        RECT 85.890 126.370 86.030 127.750 ;
        RECT 86.350 126.710 86.490 130.130 ;
        RECT 86.290 126.390 86.550 126.710 ;
        RECT 85.830 126.050 86.090 126.370 ;
        RECT 85.360 125.175 85.640 125.545 ;
        RECT 85.890 125.350 86.030 126.050 ;
        RECT 86.290 125.370 86.550 125.690 ;
        RECT 85.830 125.030 86.090 125.350 ;
        RECT 85.360 124.495 85.640 124.865 ;
        RECT 86.350 124.750 86.490 125.370 ;
        RECT 85.890 124.610 86.490 124.750 ;
        RECT 85.430 123.310 85.570 124.495 ;
        RECT 84.450 122.990 84.710 123.310 ;
        RECT 85.370 122.990 85.630 123.310 ;
        RECT 85.360 122.455 85.640 122.825 ;
        RECT 83.990 120.270 84.250 120.590 ;
        RECT 84.440 120.415 84.720 120.785 ;
        RECT 83.530 107.350 83.790 107.670 ;
        RECT 83.530 104.630 83.790 104.950 ;
        RECT 83.590 101.890 83.730 104.630 ;
        RECT 83.530 101.570 83.790 101.890 ;
        RECT 84.050 101.745 84.190 120.270 ;
        RECT 84.510 119.910 84.650 120.415 ;
        RECT 85.430 119.910 85.570 122.455 ;
        RECT 85.890 122.145 86.030 124.610 ;
        RECT 85.820 121.775 86.100 122.145 ;
        RECT 86.290 121.970 86.550 122.290 ;
        RECT 85.820 121.095 86.100 121.465 ;
        RECT 85.830 120.950 86.090 121.095 ;
        RECT 85.830 119.930 86.090 120.250 ;
        RECT 84.450 119.590 84.710 119.910 ;
        RECT 85.370 119.590 85.630 119.910 ;
        RECT 84.900 119.055 85.180 119.425 ;
        RECT 84.440 118.375 84.720 118.745 ;
        RECT 84.450 118.230 84.710 118.375 ;
        RECT 84.970 117.990 85.110 119.055 ;
        RECT 84.910 117.670 85.170 117.990 ;
        RECT 85.370 116.870 85.630 117.190 ;
        RECT 85.430 115.345 85.570 116.870 ;
        RECT 85.360 114.975 85.640 115.345 ;
        RECT 84.440 113.615 84.720 113.985 ;
        RECT 84.510 108.430 84.650 113.615 ;
        RECT 84.910 112.110 85.170 112.430 ;
        RECT 84.970 110.390 85.110 112.110 ;
        RECT 84.910 110.070 85.170 110.390 ;
        RECT 84.510 108.290 85.110 108.430 ;
        RECT 84.450 107.350 84.710 107.670 ;
        RECT 83.070 101.230 83.330 101.550 ;
        RECT 83.130 99.705 83.270 101.230 ;
        RECT 83.590 100.530 83.730 101.570 ;
        RECT 83.980 101.375 84.260 101.745 ;
        RECT 83.990 101.230 84.250 101.375 ;
        RECT 83.980 100.695 84.260 101.065 ;
        RECT 83.990 100.550 84.250 100.695 ;
        RECT 83.530 100.210 83.790 100.530 ;
        RECT 83.060 99.335 83.340 99.705 ;
        RECT 83.990 98.850 84.250 99.170 ;
        RECT 83.530 97.490 83.790 97.810 ;
        RECT 83.590 96.450 83.730 97.490 ;
        RECT 84.050 96.450 84.190 98.850 ;
        RECT 83.530 96.130 83.790 96.450 ;
        RECT 83.990 96.130 84.250 96.450 ;
        RECT 83.070 95.790 83.330 96.110 ;
        RECT 83.130 94.070 83.270 95.790 ;
        RECT 84.510 94.070 84.650 107.350 ;
        RECT 84.970 104.270 85.110 108.290 ;
        RECT 84.910 103.950 85.170 104.270 ;
        RECT 85.890 103.250 86.030 119.930 ;
        RECT 86.350 117.870 86.490 121.970 ;
        RECT 86.810 118.745 86.950 130.810 ;
        RECT 87.270 130.450 87.410 131.490 ;
        RECT 87.730 131.410 88.330 131.550 ;
        RECT 87.210 130.130 87.470 130.450 ;
        RECT 87.270 129.430 87.410 130.130 ;
        RECT 87.730 129.625 87.870 131.410 ;
        RECT 89.050 130.810 89.310 131.130 ;
        RECT 88.590 130.470 88.850 130.790 ;
        RECT 88.650 130.305 88.790 130.470 ;
        RECT 88.580 129.935 88.860 130.305 ;
        RECT 87.210 129.110 87.470 129.430 ;
        RECT 87.660 129.255 87.940 129.625 ;
        RECT 88.650 129.090 88.790 129.935 ;
        RECT 88.590 128.770 88.850 129.090 ;
        RECT 88.130 128.090 88.390 128.410 ;
        RECT 88.590 128.090 88.850 128.410 ;
        RECT 89.110 128.265 89.250 130.810 ;
        RECT 87.670 125.710 87.930 126.030 ;
        RECT 87.210 120.270 87.470 120.590 ;
        RECT 86.740 118.375 87.020 118.745 ;
        RECT 86.290 117.550 86.550 117.870 ;
        RECT 86.280 117.015 86.560 117.385 ;
        RECT 86.290 116.870 86.550 117.015 ;
        RECT 86.750 116.870 87.010 117.190 ;
        RECT 86.810 116.705 86.950 116.870 ;
        RECT 87.270 116.850 87.410 120.270 ;
        RECT 87.730 120.250 87.870 125.710 ;
        RECT 87.670 119.930 87.930 120.250 ;
        RECT 86.740 116.335 87.020 116.705 ;
        RECT 87.210 116.530 87.470 116.850 ;
        RECT 88.190 115.400 88.330 128.090 ;
        RECT 88.650 126.370 88.790 128.090 ;
        RECT 89.040 127.895 89.320 128.265 ;
        RECT 89.570 128.070 89.710 141.350 ;
        RECT 90.030 134.870 90.170 147.130 ;
        RECT 90.490 142.010 90.630 147.810 ;
        RECT 90.430 141.690 90.690 142.010 ;
        RECT 90.490 138.610 90.630 141.690 ;
        RECT 90.430 138.290 90.690 138.610 ;
        RECT 90.430 137.270 90.690 137.590 ;
        RECT 89.970 134.550 90.230 134.870 ;
        RECT 89.960 132.655 90.240 133.025 ;
        RECT 90.030 132.150 90.170 132.655 ;
        RECT 89.970 131.830 90.230 132.150 ;
        RECT 89.960 131.295 90.240 131.665 ;
        RECT 89.510 127.750 89.770 128.070 ;
        RECT 89.050 127.410 89.310 127.730 ;
        RECT 88.590 126.050 88.850 126.370 ;
        RECT 89.110 125.690 89.250 127.410 ;
        RECT 88.590 125.370 88.850 125.690 ;
        RECT 89.050 125.370 89.310 125.690 ;
        RECT 88.650 122.970 88.790 125.370 ;
        RECT 89.040 124.495 89.320 124.865 ;
        RECT 89.510 124.690 89.770 125.010 ;
        RECT 89.110 123.310 89.250 124.495 ;
        RECT 89.570 123.310 89.710 124.690 ;
        RECT 90.030 123.990 90.170 131.295 ;
        RECT 90.490 130.790 90.630 137.270 ;
        RECT 90.430 130.470 90.690 130.790 ;
        RECT 90.490 126.030 90.630 130.470 ;
        RECT 90.950 126.710 91.090 150.190 ;
        RECT 91.810 149.170 92.070 149.490 ;
        RECT 91.350 146.625 91.610 146.770 ;
        RECT 91.340 146.255 91.620 146.625 ;
        RECT 91.350 141.690 91.610 142.010 ;
        RECT 91.410 140.310 91.550 141.690 ;
        RECT 91.350 139.990 91.610 140.310 ;
        RECT 91.870 139.630 92.010 149.170 ;
        RECT 91.810 139.310 92.070 139.630 ;
        RECT 91.350 136.250 91.610 136.570 ;
        RECT 91.410 135.065 91.550 136.250 ;
        RECT 91.340 134.695 91.620 135.065 ;
        RECT 91.350 131.830 91.610 132.150 ;
        RECT 92.330 132.110 92.470 152.375 ;
        RECT 93.710 152.065 93.850 159.010 ;
        RECT 95.030 153.590 95.290 153.910 ;
        RECT 93.640 151.695 93.920 152.065 ;
        RECT 92.730 150.530 92.990 150.850 ;
        RECT 92.790 144.050 92.930 150.530 ;
        RECT 93.650 149.850 93.910 150.170 ;
        RECT 94.110 149.850 94.370 150.170 ;
        RECT 94.570 149.850 94.830 150.170 ;
        RECT 93.180 145.575 93.460 145.945 ;
        RECT 93.710 145.750 93.850 149.850 ;
        RECT 94.170 149.345 94.310 149.850 ;
        RECT 94.100 148.975 94.380 149.345 ;
        RECT 94.630 148.130 94.770 149.850 ;
        RECT 94.570 147.810 94.830 148.130 ;
        RECT 92.730 143.730 92.990 144.050 ;
        RECT 92.790 140.310 92.930 143.730 ;
        RECT 92.730 139.990 92.990 140.310 ;
        RECT 92.730 138.630 92.990 138.950 ;
        RECT 92.790 133.170 92.930 138.630 ;
        RECT 92.730 132.850 92.990 133.170 ;
        RECT 92.790 132.150 92.930 132.850 ;
        RECT 91.870 131.970 92.470 132.110 ;
        RECT 91.410 129.090 91.550 131.830 ;
        RECT 91.350 128.770 91.610 129.090 ;
        RECT 91.340 127.895 91.620 128.265 ;
        RECT 90.890 126.390 91.150 126.710 ;
        RECT 90.430 125.710 90.690 126.030 ;
        RECT 90.880 125.175 91.160 125.545 ;
        RECT 89.970 123.670 90.230 123.990 ;
        RECT 89.050 122.990 89.310 123.310 ;
        RECT 89.510 122.990 89.770 123.310 ;
        RECT 89.970 122.990 90.230 123.310 ;
        RECT 90.430 122.990 90.690 123.310 ;
        RECT 88.590 122.650 88.850 122.970 ;
        RECT 88.590 122.145 88.850 122.290 ;
        RECT 88.580 121.775 88.860 122.145 ;
        RECT 88.590 119.930 88.850 120.250 ;
        RECT 88.650 115.910 88.790 119.930 ;
        RECT 89.040 119.735 89.320 120.105 ;
        RECT 89.050 119.590 89.310 119.735 ;
        RECT 90.030 118.745 90.170 122.990 ;
        RECT 90.490 121.270 90.630 122.990 ;
        RECT 90.950 122.825 91.090 125.175 ;
        RECT 90.880 122.455 91.160 122.825 ;
        RECT 90.430 120.950 90.690 121.270 ;
        RECT 90.950 119.910 91.090 122.455 ;
        RECT 90.890 119.590 91.150 119.910 ;
        RECT 89.040 118.375 89.320 118.745 ;
        RECT 89.960 118.375 90.240 118.745 ;
        RECT 89.050 118.230 89.310 118.375 ;
        RECT 89.050 117.550 89.310 117.870 ;
        RECT 89.510 117.550 89.770 117.870 ;
        RECT 89.960 117.695 90.240 118.065 ;
        RECT 89.970 117.550 90.230 117.695 ;
        RECT 89.110 117.385 89.250 117.550 ;
        RECT 89.040 117.015 89.320 117.385 ;
        RECT 88.650 115.770 89.250 115.910 ;
        RECT 89.110 115.490 89.250 115.770 ;
        RECT 88.190 115.260 88.790 115.400 ;
        RECT 87.200 113.615 87.480 113.985 ;
        RECT 87.670 113.810 87.930 114.130 ;
        RECT 88.650 114.040 88.790 115.260 ;
        RECT 89.050 115.170 89.310 115.490 ;
        RECT 89.050 114.490 89.310 114.810 ;
        RECT 89.570 114.665 89.710 117.550 ;
        RECT 91.410 117.270 91.550 127.895 ;
        RECT 91.870 125.010 92.010 131.970 ;
        RECT 92.730 131.830 92.990 132.150 ;
        RECT 93.250 131.550 93.390 145.575 ;
        RECT 93.650 145.430 93.910 145.750 ;
        RECT 93.710 140.505 93.850 145.430 ;
        RECT 94.570 145.090 94.830 145.410 ;
        RECT 94.630 142.690 94.770 145.090 ;
        RECT 95.090 144.585 95.230 153.590 ;
        RECT 96.930 153.310 97.070 159.010 ;
        RECT 100.150 156.145 100.290 159.010 ;
        RECT 100.080 155.775 100.360 156.145 ;
        RECT 103.370 155.465 103.510 159.010 ;
        RECT 106.590 158.750 106.730 159.010 ;
        RECT 107.050 158.750 107.190 159.290 ;
        RECT 106.590 158.610 107.190 158.750 ;
        RECT 103.300 155.095 103.580 155.465 ;
        RECT 104.680 155.095 104.960 155.465 ;
        RECT 95.490 152.910 95.750 153.230 ;
        RECT 96.470 153.170 97.070 153.310 ;
        RECT 95.020 144.215 95.300 144.585 ;
        RECT 94.570 142.370 94.830 142.690 ;
        RECT 95.030 142.370 95.290 142.690 ;
        RECT 94.110 141.690 94.370 142.010 ;
        RECT 94.570 141.690 94.830 142.010 ;
        RECT 93.640 140.135 93.920 140.505 ;
        RECT 94.170 139.970 94.310 141.690 ;
        RECT 94.110 139.650 94.370 139.970 ;
        RECT 94.630 139.145 94.770 141.690 ;
        RECT 94.560 138.775 94.840 139.145 ;
        RECT 94.570 138.290 94.830 138.610 ;
        RECT 94.110 133.530 94.370 133.850 ;
        RECT 93.650 132.850 93.910 133.170 ;
        RECT 93.710 132.150 93.850 132.850 ;
        RECT 93.650 131.830 93.910 132.150 ;
        RECT 93.250 131.410 93.850 131.550 ;
        RECT 92.270 130.810 92.530 131.130 ;
        RECT 92.330 127.585 92.470 130.810 ;
        RECT 93.190 128.430 93.450 128.750 ;
        RECT 92.730 128.090 92.990 128.410 ;
        RECT 92.260 127.215 92.540 127.585 ;
        RECT 92.790 126.710 92.930 128.090 ;
        RECT 92.730 126.390 92.990 126.710 ;
        RECT 92.260 125.175 92.540 125.545 ;
        RECT 91.810 124.690 92.070 125.010 ;
        RECT 91.810 122.990 92.070 123.310 ;
        RECT 91.870 122.825 92.010 122.990 ;
        RECT 91.800 122.455 92.080 122.825 ;
        RECT 91.810 121.970 92.070 122.290 ;
        RECT 91.870 121.465 92.010 121.970 ;
        RECT 91.800 121.095 92.080 121.465 ;
        RECT 91.800 120.415 92.080 120.785 ;
        RECT 91.870 117.870 92.010 120.415 ;
        RECT 92.330 117.870 92.470 125.175 ;
        RECT 92.730 123.330 92.990 123.650 ;
        RECT 92.790 120.250 92.930 123.330 ;
        RECT 92.730 119.930 92.990 120.250 ;
        RECT 93.250 118.630 93.390 128.430 ;
        RECT 92.790 118.490 93.390 118.630 ;
        RECT 91.810 117.550 92.070 117.870 ;
        RECT 92.270 117.550 92.530 117.870 ;
        RECT 90.950 117.190 91.550 117.270 ;
        RECT 90.890 117.130 91.550 117.190 ;
        RECT 91.870 117.270 92.010 117.550 ;
        RECT 91.870 117.130 92.470 117.270 ;
        RECT 90.890 116.870 91.150 117.130 ;
        RECT 91.810 116.530 92.070 116.850 ;
        RECT 91.350 115.510 91.610 115.830 ;
        RECT 90.890 115.170 91.150 115.490 ;
        RECT 88.190 113.900 88.790 114.040 ;
        RECT 86.740 112.935 87.020 113.305 ;
        RECT 86.810 110.050 86.950 112.935 ;
        RECT 86.750 109.730 87.010 110.050 ;
        RECT 86.290 109.050 86.550 109.370 ;
        RECT 85.830 102.930 86.090 103.250 ;
        RECT 85.830 101.745 86.090 101.890 ;
        RECT 85.820 101.375 86.100 101.745 ;
        RECT 85.830 100.890 86.090 101.210 ;
        RECT 85.370 100.210 85.630 100.530 ;
        RECT 84.910 98.170 85.170 98.490 ;
        RECT 84.970 96.110 85.110 98.170 ;
        RECT 85.430 96.110 85.570 100.210 ;
        RECT 85.890 99.705 86.030 100.890 ;
        RECT 85.820 99.335 86.100 99.705 ;
        RECT 85.890 96.110 86.030 99.335 ;
        RECT 84.910 95.790 85.170 96.110 ;
        RECT 85.370 95.790 85.630 96.110 ;
        RECT 85.830 95.790 86.090 96.110 ;
        RECT 83.070 93.750 83.330 94.070 ;
        RECT 84.450 93.750 84.710 94.070 ;
        RECT 81.230 92.730 81.490 93.050 ;
        RECT 82.610 92.730 82.870 93.050 ;
        RECT 81.290 87.610 81.430 92.730 ;
        RECT 82.670 87.610 82.810 92.730 ;
        RECT 81.230 87.290 81.490 87.610 ;
        RECT 82.610 87.290 82.870 87.610 ;
        RECT 81.290 85.910 81.430 87.290 ;
        RECT 81.230 85.590 81.490 85.910 ;
        RECT 80.770 84.910 81.030 85.230 ;
        RECT 80.830 83.190 80.970 84.910 ;
        RECT 81.290 83.190 81.430 85.590 ;
        RECT 82.670 85.570 82.810 87.290 ;
        RECT 82.610 85.250 82.870 85.570 ;
        RECT 85.430 85.230 85.570 95.790 ;
        RECT 85.890 91.350 86.030 95.790 ;
        RECT 85.830 91.030 86.090 91.350 ;
        RECT 86.350 89.990 86.490 109.050 ;
        RECT 86.750 105.650 87.010 105.970 ;
        RECT 86.810 100.530 86.950 105.650 ;
        RECT 86.750 100.210 87.010 100.530 ;
        RECT 86.810 98.490 86.950 100.210 ;
        RECT 86.750 98.170 87.010 98.490 ;
        RECT 87.270 93.730 87.410 113.615 ;
        RECT 87.730 113.305 87.870 113.810 ;
        RECT 87.660 112.935 87.940 113.305 ;
        RECT 87.660 112.255 87.940 112.625 ;
        RECT 87.730 107.070 87.870 112.255 ;
        RECT 88.190 111.750 88.330 113.900 ;
        RECT 88.590 112.450 88.850 112.770 ;
        RECT 88.130 111.430 88.390 111.750 ;
        RECT 88.650 107.670 88.790 112.450 ;
        RECT 89.110 110.050 89.250 114.490 ;
        RECT 89.500 114.295 89.780 114.665 ;
        RECT 90.430 114.150 90.690 114.470 ;
        RECT 89.510 113.810 89.770 114.130 ;
        RECT 89.970 113.810 90.230 114.130 ;
        RECT 89.570 113.305 89.710 113.810 ;
        RECT 89.500 112.935 89.780 113.305 ;
        RECT 90.030 112.770 90.170 113.810 ;
        RECT 90.490 112.770 90.630 114.150 ;
        RECT 89.970 112.450 90.230 112.770 ;
        RECT 90.430 112.450 90.690 112.770 ;
        RECT 89.510 112.110 89.770 112.430 ;
        RECT 89.050 109.730 89.310 110.050 ;
        RECT 89.570 109.030 89.710 112.110 ;
        RECT 89.510 108.710 89.770 109.030 ;
        RECT 89.050 108.370 89.310 108.690 ;
        RECT 88.590 107.350 88.850 107.670 ;
        RECT 87.730 106.930 88.790 107.070 ;
        RECT 87.670 103.610 87.930 103.930 ;
        RECT 87.730 102.230 87.870 103.610 ;
        RECT 88.130 102.930 88.390 103.250 ;
        RECT 87.670 101.910 87.930 102.230 ;
        RECT 88.190 98.490 88.330 102.930 ;
        RECT 88.130 98.170 88.390 98.490 ;
        RECT 88.650 96.450 88.790 106.930 ;
        RECT 89.110 101.890 89.250 108.370 ;
        RECT 90.490 107.330 90.630 112.450 ;
        RECT 90.950 111.265 91.090 115.170 ;
        RECT 91.410 115.150 91.550 115.510 ;
        RECT 91.350 114.830 91.610 115.150 ;
        RECT 91.870 114.810 92.010 116.530 ;
        RECT 91.810 114.490 92.070 114.810 ;
        RECT 92.330 114.470 92.470 117.130 ;
        RECT 92.270 114.150 92.530 114.470 ;
        RECT 91.350 113.810 91.610 114.130 ;
        RECT 90.880 110.895 91.160 111.265 ;
        RECT 90.890 108.370 91.150 108.690 ;
        RECT 90.430 107.070 90.690 107.330 ;
        RECT 89.570 107.010 90.690 107.070 ;
        RECT 89.570 106.930 90.630 107.010 ;
        RECT 90.950 106.990 91.090 108.370 ;
        RECT 91.410 107.670 91.550 113.810 ;
        RECT 92.260 113.615 92.540 113.985 ;
        RECT 91.810 112.110 92.070 112.430 ;
        RECT 91.350 107.350 91.610 107.670 ;
        RECT 91.870 106.990 92.010 112.110 ;
        RECT 89.570 106.650 89.710 106.930 ;
        RECT 90.890 106.670 91.150 106.990 ;
        RECT 91.810 106.670 92.070 106.990 ;
        RECT 89.510 106.330 89.770 106.650 ;
        RECT 91.870 104.950 92.010 106.670 ;
        RECT 91.810 104.630 92.070 104.950 ;
        RECT 89.970 103.610 90.230 103.930 ;
        RECT 89.510 102.930 89.770 103.250 ;
        RECT 89.570 101.890 89.710 102.930 ;
        RECT 89.050 101.570 89.310 101.890 ;
        RECT 89.510 101.570 89.770 101.890 ;
        RECT 89.110 100.870 89.250 101.570 ;
        RECT 89.050 100.550 89.310 100.870 ;
        RECT 90.030 100.530 90.170 103.610 ;
        RECT 90.890 103.270 91.150 103.590 ;
        RECT 90.950 102.230 91.090 103.270 ;
        RECT 92.330 102.230 92.470 113.615 ;
        RECT 92.790 113.110 92.930 118.490 ;
        RECT 93.180 114.295 93.460 114.665 ;
        RECT 92.730 112.790 92.990 113.110 ;
        RECT 93.250 107.750 93.390 114.295 ;
        RECT 93.710 113.110 93.850 131.410 ;
        RECT 94.170 128.410 94.310 133.530 ;
        RECT 94.110 128.090 94.370 128.410 ;
        RECT 94.100 123.815 94.380 124.185 ;
        RECT 94.170 121.270 94.310 123.815 ;
        RECT 94.110 120.950 94.370 121.270 ;
        RECT 94.630 120.670 94.770 138.290 ;
        RECT 95.090 131.130 95.230 142.370 ;
        RECT 95.550 141.865 95.690 152.910 ;
        RECT 96.470 147.790 96.610 153.170 ;
        RECT 97.330 152.570 97.590 152.890 ;
        RECT 96.870 150.190 97.130 150.510 ;
        RECT 96.410 147.470 96.670 147.790 ;
        RECT 96.930 147.110 97.070 150.190 ;
        RECT 97.390 147.450 97.530 152.570 ;
        RECT 98.710 150.870 98.970 151.190 ;
        RECT 103.310 150.870 103.570 151.190 ;
        RECT 97.330 147.130 97.590 147.450 ;
        RECT 96.870 146.790 97.130 147.110 ;
        RECT 97.390 145.660 97.530 147.130 ;
        RECT 96.010 145.520 97.530 145.660 ;
        RECT 96.010 142.010 96.150 145.520 ;
        RECT 96.870 144.750 97.130 145.070 ;
        RECT 96.410 144.410 96.670 144.730 ;
        RECT 95.480 141.495 95.760 141.865 ;
        RECT 95.950 141.690 96.210 142.010 ;
        RECT 96.010 137.590 96.150 141.690 ;
        RECT 96.470 141.670 96.610 144.410 ;
        RECT 96.410 141.350 96.670 141.670 ;
        RECT 96.410 138.970 96.670 139.290 ;
        RECT 96.470 138.465 96.610 138.970 ;
        RECT 96.400 138.095 96.680 138.465 ;
        RECT 95.950 137.270 96.210 137.590 ;
        RECT 95.950 134.210 96.210 134.530 ;
        RECT 95.490 133.870 95.750 134.190 ;
        RECT 95.030 130.810 95.290 131.130 ;
        RECT 95.030 128.770 95.290 129.090 ;
        RECT 95.090 125.010 95.230 128.770 ;
        RECT 95.550 126.370 95.690 133.870 ;
        RECT 96.010 129.090 96.150 134.210 ;
        RECT 96.930 133.170 97.070 144.750 ;
        RECT 97.330 144.410 97.590 144.730 ;
        RECT 97.390 141.330 97.530 144.410 ;
        RECT 97.790 144.070 98.050 144.390 ;
        RECT 97.330 141.010 97.590 141.330 ;
        RECT 96.870 132.850 97.130 133.170 ;
        RECT 96.860 131.975 97.140 132.345 ;
        RECT 96.930 131.810 97.070 131.975 ;
        RECT 96.870 131.490 97.130 131.810 ;
        RECT 95.950 128.770 96.210 129.090 ;
        RECT 95.950 128.090 96.210 128.410 ;
        RECT 95.490 126.050 95.750 126.370 ;
        RECT 95.030 124.690 95.290 125.010 ;
        RECT 96.010 123.990 96.150 128.090 ;
        RECT 96.930 125.690 97.070 131.490 ;
        RECT 97.390 131.130 97.530 141.010 ;
        RECT 97.850 139.630 97.990 144.070 ;
        RECT 98.250 141.010 98.510 141.330 ;
        RECT 97.790 139.310 98.050 139.630 ;
        RECT 98.310 139.290 98.450 141.010 ;
        RECT 98.770 139.630 98.910 150.870 ;
        RECT 101.930 150.530 102.190 150.850 ;
        RECT 99.630 146.790 99.890 147.110 ;
        RECT 99.170 141.690 99.430 142.010 ;
        RECT 98.710 139.310 98.970 139.630 ;
        RECT 98.250 138.970 98.510 139.290 ;
        RECT 98.710 138.630 98.970 138.950 ;
        RECT 98.770 136.910 98.910 138.630 ;
        RECT 98.710 136.590 98.970 136.910 ;
        RECT 97.790 136.250 98.050 136.570 ;
        RECT 97.850 133.170 97.990 136.250 ;
        RECT 97.790 132.850 98.050 133.170 ;
        RECT 99.230 133.025 99.370 141.690 ;
        RECT 99.690 141.330 99.830 146.790 ;
        RECT 101.010 144.750 101.270 145.070 ;
        RECT 100.090 144.410 100.350 144.730 ;
        RECT 99.630 141.010 99.890 141.330 ;
        RECT 99.690 139.630 99.830 141.010 ;
        RECT 99.630 139.310 99.890 139.630 ;
        RECT 99.630 138.630 99.890 138.950 ;
        RECT 99.160 132.655 99.440 133.025 ;
        RECT 97.780 131.975 98.060 132.345 ;
        RECT 97.850 131.130 97.990 131.975 ;
        RECT 99.690 131.550 99.830 138.630 ;
        RECT 100.150 138.350 100.290 144.410 ;
        RECT 100.150 138.210 100.750 138.350 ;
        RECT 100.090 135.570 100.350 135.890 ;
        RECT 99.230 131.410 99.830 131.550 ;
        RECT 97.330 130.810 97.590 131.130 ;
        RECT 97.790 130.810 98.050 131.130 ;
        RECT 97.390 127.730 97.530 130.810 ;
        RECT 97.330 127.410 97.590 127.730 ;
        RECT 97.320 126.535 97.600 126.905 ;
        RECT 96.870 125.370 97.130 125.690 ;
        RECT 97.390 123.990 97.530 126.535 ;
        RECT 95.950 123.670 96.210 123.990 ;
        RECT 96.870 123.670 97.130 123.990 ;
        RECT 97.330 123.670 97.590 123.990 ;
        RECT 95.490 122.650 95.750 122.970 ;
        RECT 95.550 120.930 95.690 122.650 ;
        RECT 96.930 122.290 97.070 123.670 ;
        RECT 97.320 123.135 97.600 123.505 ;
        RECT 97.330 122.990 97.590 123.135 ;
        RECT 97.850 122.970 97.990 130.810 ;
        RECT 99.230 128.945 99.370 131.410 ;
        RECT 100.150 131.130 100.290 135.570 ;
        RECT 99.630 130.810 99.890 131.130 ;
        RECT 100.090 130.810 100.350 131.130 ;
        RECT 99.160 128.575 99.440 128.945 ;
        RECT 98.240 127.215 98.520 127.585 ;
        RECT 98.710 127.410 98.970 127.730 ;
        RECT 98.310 123.990 98.450 127.215 ;
        RECT 98.250 123.670 98.510 123.990 ;
        RECT 97.790 122.650 98.050 122.970 ;
        RECT 96.870 121.970 97.130 122.290 ;
        RECT 97.790 121.970 98.050 122.290 ;
        RECT 94.170 120.530 94.770 120.670 ;
        RECT 95.490 120.610 95.750 120.930 ;
        RECT 96.410 120.610 96.670 120.930 ;
        RECT 96.930 120.785 97.070 121.970 ;
        RECT 97.320 121.095 97.600 121.465 ;
        RECT 94.170 116.850 94.310 120.530 ;
        RECT 94.560 119.735 94.840 120.105 ;
        RECT 95.490 119.930 95.750 120.250 ;
        RECT 94.570 119.590 94.830 119.735 ;
        RECT 94.630 118.745 94.770 119.590 ;
        RECT 94.560 118.375 94.840 118.745 ;
        RECT 95.550 118.120 95.690 119.930 ;
        RECT 96.470 118.745 96.610 120.610 ;
        RECT 96.860 120.415 97.140 120.785 ;
        RECT 97.390 120.250 97.530 121.095 ;
        RECT 97.850 120.250 97.990 121.970 ;
        RECT 97.330 120.160 97.590 120.250 ;
        RECT 96.930 120.020 97.590 120.160 ;
        RECT 96.400 118.375 96.680 118.745 ;
        RECT 95.950 118.120 96.210 118.210 ;
        RECT 94.560 117.695 94.840 118.065 ;
        RECT 95.550 117.980 96.210 118.120 ;
        RECT 95.950 117.890 96.210 117.980 ;
        RECT 94.110 116.530 94.370 116.850 ;
        RECT 94.110 115.170 94.370 115.490 ;
        RECT 94.170 114.665 94.310 115.170 ;
        RECT 94.100 114.295 94.380 114.665 ;
        RECT 94.110 113.810 94.370 114.130 ;
        RECT 94.170 113.110 94.310 113.810 ;
        RECT 93.650 112.790 93.910 113.110 ;
        RECT 94.110 112.790 94.370 113.110 ;
        RECT 94.630 112.430 94.770 117.695 ;
        RECT 95.030 117.210 95.290 117.530 ;
        RECT 95.090 116.850 95.230 117.210 ;
        RECT 95.480 117.015 95.760 117.385 ;
        RECT 95.030 116.530 95.290 116.850 ;
        RECT 94.570 112.110 94.830 112.430 ;
        RECT 95.090 111.830 95.230 116.530 ;
        RECT 95.550 114.130 95.690 117.015 ;
        RECT 96.010 114.810 96.150 117.890 ;
        RECT 96.400 117.695 96.680 118.065 ;
        RECT 96.930 117.870 97.070 120.020 ;
        RECT 97.330 119.930 97.590 120.020 ;
        RECT 97.790 119.930 98.050 120.250 ;
        RECT 95.950 114.490 96.210 114.810 ;
        RECT 95.490 113.810 95.750 114.130 ;
        RECT 95.950 113.985 96.210 114.130 ;
        RECT 95.940 113.615 96.220 113.985 ;
        RECT 95.950 112.340 96.210 112.430 ;
        RECT 96.470 112.340 96.610 117.695 ;
        RECT 96.870 117.550 97.130 117.870 ;
        RECT 97.330 117.780 97.590 117.870 ;
        RECT 97.850 117.780 97.990 119.930 ;
        RECT 98.250 119.590 98.510 119.910 ;
        RECT 98.310 117.870 98.450 119.590 ;
        RECT 97.330 117.640 97.990 117.780 ;
        RECT 97.330 117.550 97.590 117.640 ;
        RECT 98.250 117.550 98.510 117.870 ;
        RECT 97.330 116.530 97.590 116.850 ;
        RECT 96.870 113.810 97.130 114.130 ;
        RECT 96.930 112.430 97.070 113.810 ;
        RECT 95.950 112.200 96.610 112.340 ;
        RECT 95.950 112.110 96.210 112.200 ;
        RECT 96.870 112.110 97.130 112.430 ;
        RECT 95.090 111.690 96.610 111.830 ;
        RECT 94.110 110.070 94.370 110.390 ;
        RECT 93.250 107.610 93.850 107.750 ;
        RECT 93.190 106.670 93.450 106.990 ;
        RECT 92.730 106.330 92.990 106.650 ;
        RECT 90.890 101.910 91.150 102.230 ;
        RECT 92.270 101.910 92.530 102.230 ;
        RECT 92.330 101.550 92.470 101.910 ;
        RECT 92.270 101.230 92.530 101.550 ;
        RECT 91.350 100.550 91.610 100.870 ;
        RECT 89.970 100.210 90.230 100.530 ;
        RECT 89.510 99.080 89.770 99.170 ;
        RECT 89.510 98.940 91.090 99.080 ;
        RECT 89.510 98.850 89.770 98.940 ;
        RECT 88.590 96.130 88.850 96.450 ;
        RECT 89.970 95.790 90.230 96.110 ;
        RECT 89.510 95.450 89.770 95.770 ;
        RECT 89.570 95.090 89.710 95.450 ;
        RECT 89.050 94.770 89.310 95.090 ;
        RECT 89.510 94.770 89.770 95.090 ;
        RECT 87.210 93.410 87.470 93.730 ;
        RECT 88.130 93.070 88.390 93.390 ;
        RECT 88.190 92.710 88.330 93.070 ;
        RECT 89.110 93.050 89.250 94.770 ;
        RECT 89.050 92.730 89.310 93.050 ;
        RECT 87.670 92.390 87.930 92.710 ;
        RECT 88.130 92.390 88.390 92.710 ;
        RECT 87.730 91.010 87.870 92.390 ;
        RECT 87.670 90.690 87.930 91.010 ;
        RECT 88.190 90.670 88.330 92.390 ;
        RECT 90.030 90.670 90.170 95.790 ;
        RECT 90.950 95.430 91.090 98.940 ;
        RECT 91.410 98.830 91.550 100.550 ;
        RECT 91.350 98.510 91.610 98.830 ;
        RECT 90.890 95.110 91.150 95.430 ;
        RECT 91.350 95.110 91.610 95.430 ;
        RECT 90.430 93.410 90.690 93.730 ;
        RECT 90.950 93.470 91.090 95.110 ;
        RECT 91.410 94.070 91.550 95.110 ;
        RECT 91.350 93.750 91.610 94.070 ;
        RECT 91.810 93.470 92.070 93.730 ;
        RECT 90.950 93.410 92.070 93.470 ;
        RECT 90.490 92.960 90.630 93.410 ;
        RECT 90.950 93.330 92.010 93.410 ;
        RECT 90.890 92.960 91.150 93.050 ;
        RECT 90.490 92.820 91.150 92.960 ;
        RECT 90.890 92.730 91.150 92.820 ;
        RECT 88.130 90.350 88.390 90.670 ;
        RECT 89.970 90.350 90.230 90.670 ;
        RECT 90.890 90.350 91.150 90.670 ;
        RECT 86.290 89.670 86.550 89.990 ;
        RECT 90.950 89.650 91.090 90.350 ;
        RECT 90.890 89.330 91.150 89.650 ;
        RECT 91.410 87.610 91.550 93.330 ;
        RECT 91.810 92.050 92.070 92.370 ;
        RECT 91.870 90.670 92.010 92.050 ;
        RECT 92.790 91.010 92.930 106.330 ;
        RECT 93.250 94.070 93.390 106.670 ;
        RECT 93.190 93.750 93.450 94.070 ;
        RECT 93.190 92.390 93.450 92.710 ;
        RECT 92.730 90.690 92.990 91.010 ;
        RECT 93.250 90.670 93.390 92.390 ;
        RECT 91.810 90.350 92.070 90.670 ;
        RECT 93.190 90.350 93.450 90.670 ;
        RECT 93.250 88.630 93.390 90.350 ;
        RECT 93.190 88.310 93.450 88.630 ;
        RECT 93.710 87.950 93.850 107.610 ;
        RECT 94.170 106.990 94.310 110.070 ;
        RECT 94.570 109.050 94.830 109.370 ;
        RECT 95.950 109.050 96.210 109.370 ;
        RECT 94.110 106.670 94.370 106.990 ;
        RECT 94.630 104.270 94.770 109.050 ;
        RECT 95.030 106.670 95.290 106.990 ;
        RECT 94.570 103.950 94.830 104.270 ;
        RECT 94.110 100.890 94.370 101.210 ;
        RECT 94.170 98.490 94.310 100.890 ;
        RECT 94.570 100.550 94.830 100.870 ;
        RECT 94.110 98.170 94.370 98.490 ;
        RECT 94.630 97.810 94.770 100.550 ;
        RECT 95.090 97.810 95.230 106.670 ;
        RECT 96.010 103.930 96.150 109.050 ;
        RECT 96.470 106.990 96.610 111.690 ;
        RECT 96.930 107.330 97.070 112.110 ;
        RECT 97.390 112.090 97.530 116.530 ;
        RECT 97.780 115.655 98.060 116.025 ;
        RECT 97.850 114.130 97.990 115.655 ;
        RECT 98.250 114.490 98.510 114.810 ;
        RECT 97.790 113.810 98.050 114.130 ;
        RECT 98.310 112.625 98.450 114.490 ;
        RECT 98.240 112.255 98.520 112.625 ;
        RECT 97.330 111.770 97.590 112.090 ;
        RECT 96.870 107.010 97.130 107.330 ;
        RECT 96.410 106.670 96.670 106.990 ;
        RECT 96.470 104.950 96.610 106.670 ;
        RECT 96.410 104.630 96.670 104.950 ;
        RECT 95.950 103.610 96.210 103.930 ;
        RECT 94.570 97.490 94.830 97.810 ;
        RECT 95.030 97.490 95.290 97.810 ;
        RECT 96.010 96.790 96.150 103.610 ;
        RECT 96.410 101.570 96.670 101.890 ;
        RECT 96.470 100.530 96.610 101.570 ;
        RECT 96.410 100.210 96.670 100.530 ;
        RECT 95.950 96.470 96.210 96.790 ;
        RECT 95.950 95.110 96.210 95.430 ;
        RECT 94.570 93.750 94.830 94.070 ;
        RECT 94.110 92.730 94.370 93.050 ;
        RECT 94.170 90.670 94.310 92.730 ;
        RECT 94.110 90.350 94.370 90.670 ;
        RECT 94.630 89.650 94.770 93.750 ;
        RECT 96.010 93.050 96.150 95.110 ;
        RECT 96.870 94.770 97.130 95.090 ;
        RECT 96.930 93.050 97.070 94.770 ;
        RECT 95.030 92.960 95.290 93.050 ;
        RECT 95.030 92.820 95.690 92.960 ;
        RECT 95.030 92.730 95.290 92.820 ;
        RECT 95.550 90.670 95.690 92.820 ;
        RECT 95.950 92.730 96.210 93.050 ;
        RECT 96.870 92.730 97.130 93.050 ;
        RECT 96.010 91.010 96.150 92.730 ;
        RECT 95.950 90.690 96.210 91.010 ;
        RECT 95.490 90.350 95.750 90.670 ;
        RECT 95.950 90.010 96.210 90.330 ;
        RECT 94.570 89.330 94.830 89.650 ;
        RECT 93.650 87.630 93.910 87.950 ;
        RECT 91.350 87.290 91.610 87.610 ;
        RECT 85.370 84.910 85.630 85.230 ;
        RECT 93.710 84.550 93.850 87.630 ;
        RECT 96.010 85.570 96.150 90.010 ;
        RECT 96.930 88.630 97.070 92.730 ;
        RECT 96.870 88.310 97.130 88.630 ;
        RECT 96.930 87.270 97.070 88.310 ;
        RECT 97.390 87.610 97.530 111.770 ;
        RECT 97.790 111.660 98.050 111.750 ;
        RECT 98.310 111.660 98.450 112.255 ;
        RECT 97.790 111.520 98.450 111.660 ;
        RECT 97.790 111.430 98.050 111.520 ;
        RECT 98.770 110.585 98.910 127.410 ;
        RECT 99.690 123.990 99.830 130.810 ;
        RECT 100.610 127.730 100.750 138.210 ;
        RECT 101.070 129.430 101.210 144.750 ;
        RECT 101.470 144.410 101.730 144.730 ;
        RECT 101.530 132.345 101.670 144.410 ;
        RECT 101.990 143.225 102.130 150.530 ;
        RECT 103.370 148.470 103.510 150.870 ;
        RECT 104.230 149.170 104.490 149.490 ;
        RECT 103.310 148.150 103.570 148.470 ;
        RECT 103.770 147.305 104.030 147.450 ;
        RECT 103.760 146.935 104.040 147.305 ;
        RECT 103.310 145.090 103.570 145.410 ;
        RECT 102.850 144.410 103.110 144.730 ;
        RECT 102.390 143.730 102.650 144.050 ;
        RECT 101.920 142.855 102.200 143.225 ;
        RECT 102.450 135.890 102.590 143.730 ;
        RECT 102.910 139.145 103.050 144.410 ;
        RECT 102.840 138.775 103.120 139.145 ;
        RECT 103.370 138.350 103.510 145.090 ;
        RECT 103.770 144.750 104.030 145.070 ;
        RECT 102.910 138.210 103.510 138.350 ;
        RECT 102.390 135.570 102.650 135.890 ;
        RECT 101.460 131.975 101.740 132.345 ;
        RECT 101.010 129.110 101.270 129.430 ;
        RECT 101.470 128.090 101.730 128.410 ;
        RECT 100.550 127.410 100.810 127.730 ;
        RECT 101.530 126.710 101.670 128.090 ;
        RECT 101.470 126.390 101.730 126.710 ;
        RECT 100.090 124.690 100.350 125.010 ;
        RECT 99.630 123.670 99.890 123.990 ;
        RECT 99.630 123.220 99.890 123.310 ;
        RECT 100.150 123.220 100.290 124.690 ;
        RECT 99.630 123.080 100.290 123.220 ;
        RECT 100.540 123.135 100.820 123.505 ;
        RECT 101.530 123.310 101.670 126.390 ;
        RECT 101.930 125.710 102.190 126.030 ;
        RECT 99.630 122.990 99.890 123.080 ;
        RECT 100.150 121.270 100.290 123.080 ;
        RECT 100.550 122.990 100.810 123.135 ;
        RECT 101.470 122.990 101.730 123.310 ;
        RECT 100.550 122.310 100.810 122.630 ;
        RECT 101.010 122.310 101.270 122.630 ;
        RECT 100.090 120.950 100.350 121.270 ;
        RECT 99.630 120.270 99.890 120.590 ;
        RECT 99.170 119.930 99.430 120.250 ;
        RECT 99.230 118.550 99.370 119.930 ;
        RECT 99.170 118.230 99.430 118.550 ;
        RECT 99.170 117.550 99.430 117.870 ;
        RECT 99.230 115.830 99.370 117.550 ;
        RECT 99.690 116.850 99.830 120.270 ;
        RECT 99.630 116.530 99.890 116.850 ;
        RECT 99.170 115.510 99.430 115.830 ;
        RECT 99.230 115.150 99.370 115.510 ;
        RECT 99.170 114.830 99.430 115.150 ;
        RECT 99.630 114.830 99.890 115.150 ;
        RECT 99.160 114.295 99.440 114.665 ;
        RECT 99.170 114.150 99.430 114.295 ;
        RECT 98.700 110.215 98.980 110.585 ;
        RECT 99.230 109.710 99.370 114.150 ;
        RECT 99.690 112.430 99.830 114.830 ;
        RECT 100.150 114.810 100.290 120.950 ;
        RECT 100.610 118.210 100.750 122.310 ;
        RECT 100.550 117.890 100.810 118.210 ;
        RECT 100.550 117.210 100.810 117.530 ;
        RECT 100.610 116.850 100.750 117.210 ;
        RECT 100.550 116.530 100.810 116.850 ;
        RECT 100.550 115.510 100.810 115.830 ;
        RECT 100.610 115.345 100.750 115.510 ;
        RECT 100.540 114.975 100.820 115.345 ;
        RECT 100.090 114.490 100.350 114.810 ;
        RECT 100.550 114.490 100.810 114.810 ;
        RECT 99.630 112.110 99.890 112.430 ;
        RECT 100.610 111.750 100.750 114.490 ;
        RECT 101.070 112.625 101.210 122.310 ;
        RECT 101.530 120.250 101.670 122.990 ;
        RECT 101.990 121.270 102.130 125.710 ;
        RECT 102.910 122.290 103.050 138.210 ;
        RECT 103.310 135.570 103.570 135.890 ;
        RECT 103.370 134.270 103.510 135.570 ;
        RECT 103.830 134.870 103.970 144.750 ;
        RECT 104.290 136.230 104.430 149.170 ;
        RECT 104.750 138.465 104.890 155.095 ;
        RECT 107.450 152.230 107.710 152.550 ;
        RECT 107.510 150.850 107.650 152.230 ;
        RECT 107.900 151.015 108.180 151.385 ;
        RECT 107.450 150.530 107.710 150.850 ;
        RECT 105.150 150.190 105.410 150.510 ;
        RECT 105.610 150.190 105.870 150.510 ;
        RECT 106.530 150.190 106.790 150.510 ;
        RECT 105.210 146.625 105.350 150.190 ;
        RECT 105.140 146.255 105.420 146.625 ;
        RECT 105.150 145.430 105.410 145.750 ;
        RECT 105.210 144.730 105.350 145.430 ;
        RECT 105.150 144.410 105.410 144.730 ;
        RECT 105.210 140.310 105.350 144.410 ;
        RECT 105.150 139.990 105.410 140.310 ;
        RECT 105.670 139.630 105.810 150.190 ;
        RECT 106.070 147.470 106.330 147.790 ;
        RECT 106.130 145.750 106.270 147.470 ;
        RECT 106.070 145.430 106.330 145.750 ;
        RECT 106.590 144.730 106.730 150.190 ;
        RECT 107.970 147.305 108.110 151.015 ;
        RECT 106.990 146.790 107.250 147.110 ;
        RECT 107.900 146.935 108.180 147.305 ;
        RECT 107.050 144.730 107.190 146.790 ;
        RECT 107.450 146.450 107.710 146.770 ;
        RECT 107.510 145.750 107.650 146.450 ;
        RECT 107.450 145.430 107.710 145.750 ;
        RECT 107.900 144.895 108.180 145.265 ;
        RECT 106.530 144.410 106.790 144.730 ;
        RECT 106.990 144.410 107.250 144.730 ;
        RECT 107.450 144.410 107.710 144.730 ;
        RECT 107.510 141.185 107.650 144.410 ;
        RECT 107.440 140.815 107.720 141.185 ;
        RECT 106.070 139.990 106.330 140.310 ;
        RECT 105.610 139.310 105.870 139.630 ;
        RECT 104.680 138.095 104.960 138.465 ;
        RECT 105.140 136.735 105.420 137.105 ;
        RECT 104.230 135.910 104.490 136.230 ;
        RECT 104.690 135.570 104.950 135.890 ;
        RECT 103.770 134.550 104.030 134.870 ;
        RECT 103.370 134.130 103.970 134.270 ;
        RECT 103.830 133.850 103.970 134.130 ;
        RECT 103.770 133.530 104.030 133.850 ;
        RECT 103.310 126.390 103.570 126.710 ;
        RECT 103.370 124.920 103.510 126.390 ;
        RECT 103.830 125.690 103.970 133.530 ;
        RECT 104.230 131.150 104.490 131.470 ;
        RECT 103.770 125.370 104.030 125.690 ;
        RECT 103.370 124.780 103.970 124.920 ;
        RECT 102.850 121.970 103.110 122.290 ;
        RECT 101.930 120.950 102.190 121.270 ;
        RECT 102.850 120.270 103.110 120.590 ;
        RECT 101.470 119.930 101.730 120.250 ;
        RECT 101.920 119.735 102.200 120.105 ;
        RECT 101.990 119.310 102.130 119.735 ;
        RECT 101.530 119.170 102.130 119.310 ;
        RECT 101.530 117.530 101.670 119.170 ;
        RECT 102.910 117.530 103.050 120.270 ;
        RECT 103.830 118.630 103.970 124.780 ;
        RECT 104.290 123.990 104.430 131.150 ;
        RECT 104.230 123.670 104.490 123.990 ;
        RECT 103.370 118.490 103.970 118.630 ;
        RECT 103.370 117.870 103.510 118.490 ;
        RECT 104.220 118.375 104.500 118.745 ;
        RECT 103.310 117.550 103.570 117.870 ;
        RECT 103.760 117.695 104.040 118.065 ;
        RECT 101.470 117.210 101.730 117.530 ;
        RECT 102.850 117.210 103.110 117.530 ;
        RECT 102.910 116.850 103.050 117.210 ;
        RECT 101.470 116.530 101.730 116.850 ;
        RECT 102.850 116.530 103.110 116.850 ;
        RECT 101.000 112.255 101.280 112.625 ;
        RECT 100.550 111.430 100.810 111.750 ;
        RECT 101.530 111.265 101.670 116.530 ;
        RECT 102.390 114.665 102.650 114.810 ;
        RECT 102.380 114.295 102.660 114.665 ;
        RECT 102.850 114.490 103.110 114.810 ;
        RECT 102.910 114.130 103.050 114.490 ;
        RECT 102.850 113.810 103.110 114.130 ;
        RECT 102.840 112.935 103.120 113.305 ;
        RECT 102.910 111.750 103.050 112.935 ;
        RECT 103.370 111.830 103.510 117.550 ;
        RECT 103.830 114.810 103.970 117.695 ;
        RECT 103.770 114.490 104.030 114.810 ;
        RECT 103.760 113.615 104.040 113.985 ;
        RECT 103.830 112.430 103.970 113.615 ;
        RECT 104.290 113.110 104.430 118.375 ;
        RECT 104.230 112.790 104.490 113.110 ;
        RECT 104.750 112.770 104.890 135.570 ;
        RECT 105.210 123.505 105.350 136.735 ;
        RECT 106.130 133.850 106.270 139.990 ;
        RECT 107.970 139.970 108.110 144.895 ;
        RECT 107.910 139.650 108.170 139.970 ;
        RECT 106.530 139.310 106.790 139.630 ;
        RECT 106.590 136.910 106.730 139.310 ;
        RECT 106.530 136.590 106.790 136.910 ;
        RECT 107.910 136.590 108.170 136.910 ;
        RECT 107.450 136.250 107.710 136.570 ;
        RECT 106.990 133.870 107.250 134.190 ;
        RECT 106.070 133.530 106.330 133.850 ;
        RECT 106.060 131.975 106.340 132.345 ;
        RECT 105.610 130.130 105.870 130.450 ;
        RECT 105.140 123.135 105.420 123.505 ;
        RECT 105.150 122.310 105.410 122.630 ;
        RECT 105.210 120.250 105.350 122.310 ;
        RECT 105.670 120.250 105.810 130.130 ;
        RECT 105.150 119.930 105.410 120.250 ;
        RECT 105.610 119.930 105.870 120.250 ;
        RECT 105.150 119.250 105.410 119.570 ;
        RECT 105.210 118.210 105.350 119.250 ;
        RECT 105.150 117.890 105.410 118.210 ;
        RECT 104.690 112.450 104.950 112.770 ;
        RECT 103.770 112.110 104.030 112.430 ;
        RECT 105.210 112.000 105.350 117.890 ;
        RECT 105.600 117.695 105.880 118.065 ;
        RECT 105.670 115.150 105.810 117.695 ;
        RECT 106.130 115.830 106.270 131.975 ;
        RECT 107.050 130.450 107.190 133.870 ;
        RECT 107.510 132.150 107.650 136.250 ;
        RECT 107.450 131.830 107.710 132.150 ;
        RECT 107.510 131.130 107.650 131.830 ;
        RECT 107.450 130.810 107.710 131.130 ;
        RECT 106.990 130.130 107.250 130.450 ;
        RECT 106.530 124.690 106.790 125.010 ;
        RECT 106.590 119.570 106.730 124.690 ;
        RECT 107.050 120.250 107.190 130.130 ;
        RECT 107.450 129.110 107.710 129.430 ;
        RECT 107.510 121.270 107.650 129.110 ;
        RECT 107.450 120.950 107.710 121.270 ;
        RECT 107.440 120.415 107.720 120.785 ;
        RECT 106.990 119.930 107.250 120.250 ;
        RECT 106.530 119.250 106.790 119.570 ;
        RECT 106.070 115.510 106.330 115.830 ;
        RECT 105.610 114.830 105.870 115.150 ;
        RECT 106.590 114.550 106.730 119.250 ;
        RECT 106.990 118.460 107.250 118.550 ;
        RECT 107.510 118.460 107.650 120.415 ;
        RECT 106.990 118.320 107.650 118.460 ;
        RECT 106.990 118.230 107.250 118.320 ;
        RECT 106.990 117.550 107.250 117.870 ;
        RECT 107.050 116.850 107.190 117.550 ;
        RECT 107.450 116.870 107.710 117.190 ;
        RECT 106.990 116.530 107.250 116.850 ;
        RECT 105.670 114.410 106.730 114.550 ;
        RECT 105.670 112.430 105.810 114.410 ;
        RECT 106.070 113.985 106.330 114.130 ;
        RECT 106.060 113.615 106.340 113.985 ;
        RECT 105.610 112.110 105.870 112.430 ;
        RECT 104.290 111.860 105.350 112.000 ;
        RECT 101.930 111.430 102.190 111.750 ;
        RECT 102.850 111.430 103.110 111.750 ;
        RECT 103.370 111.690 103.970 111.830 ;
        RECT 101.460 110.895 101.740 111.265 ;
        RECT 101.010 110.070 101.270 110.390 ;
        RECT 97.790 109.390 98.050 109.710 ;
        RECT 99.170 109.390 99.430 109.710 ;
        RECT 97.850 98.490 97.990 109.390 ;
        RECT 101.070 109.370 101.210 110.070 ;
        RECT 101.010 109.050 101.270 109.370 ;
        RECT 101.470 109.050 101.730 109.370 ;
        RECT 101.990 109.280 102.130 111.430 ;
        RECT 102.850 109.905 103.110 110.050 ;
        RECT 102.840 109.535 103.120 109.905 ;
        RECT 103.310 109.280 103.570 109.370 ;
        RECT 101.990 109.140 103.570 109.280 ;
        RECT 101.530 106.310 101.670 109.050 ;
        RECT 101.470 105.990 101.730 106.310 ;
        RECT 101.990 104.270 102.130 109.140 ;
        RECT 103.310 109.050 103.570 109.140 ;
        RECT 102.850 108.370 103.110 108.690 ;
        RECT 102.910 107.330 103.050 108.370 ;
        RECT 102.850 107.010 103.110 107.330 ;
        RECT 103.830 107.070 103.970 111.690 ;
        RECT 104.290 107.670 104.430 111.860 ;
        RECT 105.140 110.895 105.420 111.265 ;
        RECT 104.690 109.050 104.950 109.370 ;
        RECT 104.230 107.350 104.490 107.670 ;
        RECT 101.930 103.950 102.190 104.270 ;
        RECT 99.170 102.930 99.430 103.250 ;
        RECT 99.630 102.930 99.890 103.250 ;
        RECT 99.230 102.230 99.370 102.930 ;
        RECT 99.170 101.910 99.430 102.230 ;
        RECT 99.230 101.550 99.370 101.910 ;
        RECT 99.170 101.230 99.430 101.550 ;
        RECT 98.250 100.890 98.510 101.210 ;
        RECT 98.310 98.490 98.450 100.890 ;
        RECT 99.230 98.490 99.370 101.230 ;
        RECT 99.690 98.830 99.830 102.930 ;
        RECT 100.550 101.570 100.810 101.890 ;
        RECT 99.630 98.510 99.890 98.830 ;
        RECT 97.790 98.170 98.050 98.490 ;
        RECT 98.250 98.170 98.510 98.490 ;
        RECT 99.170 98.170 99.430 98.490 ;
        RECT 99.230 93.050 99.370 98.170 ;
        RECT 100.610 98.150 100.750 101.570 ;
        RECT 101.010 100.890 101.270 101.210 ;
        RECT 101.070 98.490 101.210 100.890 ;
        RECT 102.910 99.510 103.050 107.010 ;
        RECT 103.830 106.930 104.430 107.070 ;
        RECT 103.770 106.330 104.030 106.650 ;
        RECT 103.830 102.230 103.970 106.330 ;
        RECT 103.770 101.910 104.030 102.230 ;
        RECT 101.470 99.190 101.730 99.510 ;
        RECT 102.850 99.190 103.110 99.510 ;
        RECT 101.010 98.170 101.270 98.490 ;
        RECT 100.550 97.830 100.810 98.150 ;
        RECT 101.010 97.490 101.270 97.810 ;
        RECT 99.170 92.730 99.430 93.050 ;
        RECT 97.790 90.350 98.050 90.670 ;
        RECT 97.850 88.630 97.990 90.350 ;
        RECT 99.230 88.630 99.370 92.730 ;
        RECT 100.550 92.620 100.810 92.710 ;
        RECT 101.070 92.620 101.210 97.490 ;
        RECT 101.530 93.730 101.670 99.190 ;
        RECT 101.930 98.510 102.190 98.830 ;
        RECT 101.990 94.070 102.130 98.510 ;
        RECT 104.290 95.430 104.430 106.930 ;
        RECT 104.750 100.530 104.890 109.050 ;
        RECT 104.690 100.210 104.950 100.530 ;
        RECT 104.230 95.110 104.490 95.430 ;
        RECT 101.930 93.750 102.190 94.070 ;
        RECT 101.470 93.410 101.730 93.730 ;
        RECT 100.550 92.480 101.210 92.620 ;
        RECT 100.550 92.390 100.810 92.480 ;
        RECT 100.610 89.990 100.750 92.390 ;
        RECT 101.530 91.350 101.670 93.410 ;
        RECT 101.470 91.030 101.730 91.350 ;
        RECT 100.550 89.670 100.810 89.990 ;
        RECT 97.790 88.310 98.050 88.630 ;
        RECT 99.170 88.310 99.430 88.630 ;
        RECT 101.990 87.610 102.130 93.750 ;
        RECT 105.210 93.050 105.350 110.895 ;
        RECT 105.610 109.100 105.870 109.420 ;
        RECT 105.670 106.310 105.810 109.100 ;
        RECT 106.130 107.330 106.270 113.615 ;
        RECT 106.530 112.110 106.790 112.430 ;
        RECT 106.590 109.710 106.730 112.110 ;
        RECT 106.530 109.390 106.790 109.710 ;
        RECT 107.050 109.030 107.190 116.530 ;
        RECT 107.510 114.810 107.650 116.870 ;
        RECT 107.970 115.490 108.110 136.590 ;
        RECT 107.910 115.170 108.170 115.490 ;
        RECT 107.450 114.490 107.710 114.810 ;
        RECT 107.910 112.625 108.170 112.770 ;
        RECT 107.900 112.255 108.180 112.625 ;
        RECT 107.910 109.280 108.170 109.370 ;
        RECT 107.510 109.140 108.170 109.280 ;
        RECT 106.990 108.710 107.250 109.030 ;
        RECT 106.070 107.010 106.330 107.330 ;
        RECT 106.980 106.815 107.260 107.185 ;
        RECT 105.610 105.990 105.870 106.310 ;
        RECT 106.530 101.230 106.790 101.550 ;
        RECT 106.590 99.170 106.730 101.230 ;
        RECT 106.530 98.850 106.790 99.170 ;
        RECT 106.070 98.170 106.330 98.490 ;
        RECT 105.610 95.790 105.870 96.110 ;
        RECT 105.670 93.050 105.810 95.790 ;
        RECT 106.130 94.070 106.270 98.170 ;
        RECT 106.590 97.810 106.730 98.850 ;
        RECT 106.530 97.490 106.790 97.810 ;
        RECT 107.050 96.790 107.190 106.815 ;
        RECT 107.510 100.530 107.650 109.140 ;
        RECT 107.910 109.050 108.170 109.140 ;
        RECT 107.910 106.900 108.170 106.990 ;
        RECT 108.430 106.900 108.570 159.290 ;
        RECT 109.740 159.010 110.020 163.010 ;
        RECT 112.960 159.010 113.240 163.010 ;
        RECT 114.410 159.290 115.930 159.430 ;
        RECT 109.810 153.425 109.950 159.010 ;
        RECT 113.030 158.185 113.170 159.010 ;
        RECT 112.960 157.815 113.240 158.185 ;
        RECT 109.740 153.055 110.020 153.425 ;
        RECT 109.290 150.530 109.550 150.850 ;
        RECT 108.830 148.150 109.090 148.470 ;
        RECT 108.890 143.905 109.030 148.150 ;
        RECT 108.820 143.535 109.100 143.905 ;
        RECT 108.830 142.030 109.090 142.350 ;
        RECT 108.890 136.570 109.030 142.030 ;
        RECT 108.830 136.250 109.090 136.570 ;
        RECT 109.350 133.170 109.490 150.530 ;
        RECT 111.130 150.190 111.390 150.510 ;
        RECT 111.190 149.830 111.330 150.190 ;
        RECT 111.130 149.510 111.390 149.830 ;
        RECT 109.750 144.750 110.010 145.070 ;
        RECT 110.200 144.895 110.480 145.265 ;
        RECT 110.210 144.750 110.470 144.895 ;
        RECT 109.810 144.050 109.950 144.750 ;
        RECT 109.750 143.730 110.010 144.050 ;
        RECT 110.670 133.530 110.930 133.850 ;
        RECT 109.290 132.850 109.550 133.170 ;
        RECT 110.210 132.850 110.470 133.170 ;
        RECT 109.350 128.410 109.490 132.850 ;
        RECT 110.270 128.750 110.410 132.850 ;
        RECT 110.210 128.430 110.470 128.750 ;
        RECT 109.290 128.090 109.550 128.410 ;
        RECT 110.730 128.150 110.870 133.530 ;
        RECT 111.190 129.090 111.330 149.510 ;
        RECT 113.430 147.810 113.690 148.130 ;
        RECT 113.490 147.450 113.630 147.810 ;
        RECT 111.590 147.130 111.850 147.450 ;
        RECT 113.430 147.130 113.690 147.450 ;
        RECT 111.650 143.225 111.790 147.130 ;
        RECT 112.510 143.730 112.770 144.050 ;
        RECT 111.580 142.855 111.860 143.225 ;
        RECT 112.050 142.710 112.310 143.030 ;
        RECT 111.580 134.695 111.860 135.065 ;
        RECT 111.130 128.770 111.390 129.090 ;
        RECT 108.830 126.390 109.090 126.710 ;
        RECT 108.890 120.930 109.030 126.390 ;
        RECT 108.830 120.610 109.090 120.930 ;
        RECT 108.830 119.590 109.090 119.910 ;
        RECT 107.910 106.760 108.570 106.900 ;
        RECT 107.910 106.670 108.170 106.760 ;
        RECT 107.900 106.135 108.180 106.505 ;
        RECT 107.910 105.990 108.170 106.135 ;
        RECT 108.430 104.950 108.570 106.760 ;
        RECT 108.890 106.310 109.030 119.590 ;
        RECT 109.350 117.190 109.490 128.090 ;
        RECT 110.730 128.010 111.330 128.150 ;
        RECT 110.670 127.410 110.930 127.730 ;
        RECT 110.730 125.690 110.870 127.410 ;
        RECT 111.190 126.370 111.330 128.010 ;
        RECT 111.130 126.050 111.390 126.370 ;
        RECT 110.670 125.370 110.930 125.690 ;
        RECT 109.750 123.670 110.010 123.990 ;
        RECT 109.810 120.250 109.950 123.670 ;
        RECT 110.670 123.330 110.930 123.650 ;
        RECT 109.750 119.930 110.010 120.250 ;
        RECT 110.210 119.930 110.470 120.250 ;
        RECT 109.290 116.870 109.550 117.190 ;
        RECT 110.270 116.590 110.410 119.930 ;
        RECT 110.730 117.530 110.870 123.330 ;
        RECT 111.130 117.550 111.390 117.870 ;
        RECT 110.670 117.210 110.930 117.530 ;
        RECT 109.350 116.450 110.410 116.590 ;
        RECT 109.350 115.830 109.490 116.450 ;
        RECT 110.730 115.830 110.870 117.210 ;
        RECT 109.290 115.510 109.550 115.830 ;
        RECT 110.210 115.510 110.470 115.830 ;
        RECT 110.670 115.510 110.930 115.830 ;
        RECT 109.290 112.110 109.550 112.430 ;
        RECT 109.750 112.110 110.010 112.430 ;
        RECT 109.350 110.050 109.490 112.110 ;
        RECT 109.290 109.730 109.550 110.050 ;
        RECT 109.810 109.370 109.950 112.110 ;
        RECT 109.750 109.050 110.010 109.370 ;
        RECT 109.290 107.240 109.550 107.330 ;
        RECT 109.810 107.240 109.950 109.050 ;
        RECT 109.290 107.100 109.950 107.240 ;
        RECT 109.290 107.010 109.550 107.100 ;
        RECT 108.830 105.990 109.090 106.310 ;
        RECT 108.370 104.630 108.630 104.950 ;
        RECT 108.830 104.630 109.090 104.950 ;
        RECT 107.910 103.270 108.170 103.590 ;
        RECT 107.970 101.890 108.110 103.270 ;
        RECT 107.910 101.570 108.170 101.890 ;
        RECT 108.370 101.230 108.630 101.550 ;
        RECT 107.910 100.550 108.170 100.870 ;
        RECT 107.450 100.210 107.710 100.530 ;
        RECT 106.990 96.470 107.250 96.790 ;
        RECT 106.990 95.790 107.250 96.110 ;
        RECT 106.070 93.750 106.330 94.070 ;
        RECT 107.050 93.050 107.190 95.790 ;
        RECT 107.510 95.430 107.650 100.210 ;
        RECT 107.970 99.510 108.110 100.550 ;
        RECT 108.430 100.440 108.570 101.230 ;
        RECT 108.890 100.530 109.030 104.630 ;
        RECT 109.290 101.570 109.550 101.890 ;
        RECT 108.830 100.440 109.090 100.530 ;
        RECT 108.430 100.300 109.090 100.440 ;
        RECT 107.910 99.190 108.170 99.510 ;
        RECT 108.430 96.790 108.570 100.300 ;
        RECT 108.830 100.210 109.090 100.300 ;
        RECT 109.350 98.490 109.490 101.570 ;
        RECT 109.810 99.510 109.950 107.100 ;
        RECT 110.270 106.990 110.410 115.510 ;
        RECT 110.670 114.830 110.930 115.150 ;
        RECT 110.730 109.370 110.870 114.830 ;
        RECT 110.670 109.050 110.930 109.370 ;
        RECT 110.210 106.670 110.470 106.990 ;
        RECT 110.730 106.310 110.870 109.050 ;
        RECT 111.190 107.185 111.330 117.550 ;
        RECT 111.650 111.750 111.790 134.695 ;
        RECT 112.110 128.750 112.250 142.710 ;
        RECT 112.570 134.190 112.710 143.730 ;
        RECT 112.510 133.870 112.770 134.190 ;
        RECT 113.430 133.870 113.690 134.190 ;
        RECT 112.500 132.655 112.780 133.025 ;
        RECT 112.050 128.430 112.310 128.750 ;
        RECT 112.570 125.545 112.710 132.655 ;
        RECT 113.490 131.470 113.630 133.870 ;
        RECT 113.430 131.150 113.690 131.470 ;
        RECT 113.430 130.470 113.690 130.790 ;
        RECT 112.970 129.110 113.230 129.430 ;
        RECT 113.030 126.905 113.170 129.110 ;
        RECT 112.960 126.535 113.240 126.905 ;
        RECT 113.490 126.030 113.630 130.470 ;
        RECT 113.890 128.430 114.150 128.750 ;
        RECT 113.430 125.710 113.690 126.030 ;
        RECT 112.500 125.175 112.780 125.545 ;
        RECT 112.050 124.690 112.310 125.010 ;
        RECT 112.110 123.310 112.250 124.690 ;
        RECT 112.050 122.990 112.310 123.310 ;
        RECT 112.970 122.990 113.230 123.310 ;
        RECT 113.030 117.870 113.170 122.990 ;
        RECT 113.490 120.930 113.630 125.710 ;
        RECT 113.430 120.610 113.690 120.930 ;
        RECT 113.950 120.250 114.090 128.430 ;
        RECT 113.890 119.930 114.150 120.250 ;
        RECT 114.410 119.310 114.550 159.290 ;
        RECT 115.790 158.750 115.930 159.290 ;
        RECT 116.180 159.010 116.460 163.010 ;
        RECT 119.400 159.010 119.680 163.010 ;
        RECT 122.620 159.010 122.900 163.010 ;
        RECT 125.840 159.010 126.120 163.010 ;
        RECT 129.060 159.010 129.340 163.010 ;
        RECT 116.250 158.750 116.390 159.010 ;
        RECT 115.790 158.610 116.390 158.750 ;
        RECT 115.720 155.775 116.000 156.145 ;
        RECT 115.260 148.975 115.540 149.345 ;
        RECT 115.330 147.790 115.470 148.975 ;
        RECT 115.270 147.470 115.530 147.790 ;
        RECT 115.790 142.690 115.930 155.775 ;
        RECT 116.190 154.610 116.450 154.930 ;
        RECT 116.250 143.960 116.390 154.610 ;
        RECT 117.570 154.270 117.830 154.590 ;
        RECT 117.630 151.190 117.770 154.270 ;
        RECT 119.470 154.105 119.610 159.010 ;
        RECT 119.400 153.735 119.680 154.105 ;
        RECT 118.490 152.910 118.750 153.230 ;
        RECT 117.570 150.870 117.830 151.190 ;
        RECT 117.110 150.190 117.370 150.510 ;
        RECT 118.020 150.335 118.300 150.705 ;
        RECT 116.650 149.850 116.910 150.170 ;
        RECT 116.710 144.730 116.850 149.850 ;
        RECT 117.170 147.305 117.310 150.190 ;
        RECT 118.090 149.830 118.230 150.335 ;
        RECT 118.030 149.510 118.290 149.830 ;
        RECT 118.090 147.450 118.230 149.510 ;
        RECT 117.100 146.935 117.380 147.305 ;
        RECT 118.030 147.130 118.290 147.450 ;
        RECT 117.570 146.450 117.830 146.770 ;
        RECT 116.650 144.410 116.910 144.730 ;
        RECT 116.250 143.820 117.310 143.960 ;
        RECT 115.730 142.370 115.990 142.690 ;
        RECT 117.170 141.070 117.310 143.820 ;
        RECT 117.630 142.010 117.770 146.450 ;
        RECT 118.550 142.010 118.690 152.910 ;
        RECT 118.950 150.025 119.210 150.170 ;
        RECT 118.940 149.655 119.220 150.025 ;
        RECT 122.160 149.655 122.440 150.025 ;
        RECT 120.330 149.170 120.590 149.490 ;
        RECT 121.250 149.170 121.510 149.490 ;
        RECT 119.870 144.750 120.130 145.070 ;
        RECT 120.390 144.980 120.530 149.170 ;
        RECT 121.310 147.790 121.450 149.170 ;
        RECT 121.250 147.470 121.510 147.790 ;
        RECT 120.790 147.130 121.050 147.450 ;
        RECT 120.850 146.625 120.990 147.130 ;
        RECT 121.710 146.790 121.970 147.110 ;
        RECT 120.780 146.255 121.060 146.625 ;
        RECT 121.770 145.830 121.910 146.790 ;
        RECT 122.230 146.770 122.370 149.655 ;
        RECT 122.170 146.450 122.430 146.770 ;
        RECT 121.770 145.750 122.370 145.830 ;
        RECT 121.770 145.690 122.430 145.750 ;
        RECT 122.170 145.430 122.430 145.690 ;
        RECT 121.710 144.980 121.970 145.070 ;
        RECT 120.390 144.840 121.970 144.980 ;
        RECT 121.710 144.750 121.970 144.840 ;
        RECT 117.570 141.690 117.830 142.010 ;
        RECT 118.490 141.690 118.750 142.010 ;
        RECT 119.410 141.690 119.670 142.010 ;
        RECT 116.250 140.930 117.310 141.070 ;
        RECT 114.810 138.970 115.070 139.290 ;
        RECT 114.870 136.910 115.010 138.970 ;
        RECT 116.250 138.610 116.390 140.930 ;
        RECT 116.640 140.135 116.920 140.505 ;
        RECT 116.650 139.990 116.910 140.135 ;
        RECT 116.710 139.630 116.850 139.990 ;
        RECT 117.170 139.630 117.310 140.930 ;
        RECT 116.650 139.310 116.910 139.630 ;
        RECT 117.110 139.310 117.370 139.630 ;
        RECT 117.560 139.455 117.840 139.825 ;
        RECT 117.110 138.630 117.370 138.950 ;
        RECT 116.190 138.290 116.450 138.610 ;
        RECT 116.650 137.270 116.910 137.590 ;
        RECT 114.810 136.590 115.070 136.910 ;
        RECT 115.730 133.190 115.990 133.510 ;
        RECT 115.790 132.110 115.930 133.190 ;
        RECT 115.330 131.970 115.930 132.110 ;
        RECT 114.810 131.490 115.070 131.810 ;
        RECT 113.950 119.170 114.550 119.310 ;
        RECT 112.970 117.550 113.230 117.870 ;
        RECT 112.050 117.210 112.310 117.530 ;
        RECT 113.950 117.385 114.090 119.170 ;
        RECT 114.350 118.230 114.610 118.550 ;
        RECT 112.110 116.850 112.250 117.210 ;
        RECT 113.880 117.015 114.160 117.385 ;
        RECT 112.050 116.530 112.310 116.850 ;
        RECT 113.430 115.510 113.690 115.830 ;
        RECT 112.050 114.490 112.310 114.810 ;
        RECT 112.510 114.490 112.770 114.810 ;
        RECT 112.110 111.750 112.250 114.490 ;
        RECT 112.570 113.190 112.710 114.490 ;
        RECT 112.570 113.050 113.170 113.190 ;
        RECT 112.510 112.110 112.770 112.430 ;
        RECT 111.590 111.430 111.850 111.750 ;
        RECT 112.050 111.430 112.310 111.750 ;
        RECT 112.570 111.410 112.710 112.110 ;
        RECT 113.030 111.945 113.170 113.050 ;
        RECT 112.960 111.575 113.240 111.945 ;
        RECT 113.490 111.410 113.630 115.510 ;
        RECT 114.410 115.345 114.550 118.230 ;
        RECT 114.870 116.705 115.010 131.490 ;
        RECT 115.330 125.430 115.470 131.970 ;
        RECT 115.730 126.110 115.990 126.370 ;
        RECT 115.730 126.050 116.390 126.110 ;
        RECT 115.790 125.970 116.390 126.050 ;
        RECT 116.250 125.690 116.390 125.970 ;
        RECT 115.730 125.430 115.990 125.690 ;
        RECT 115.330 125.370 115.990 125.430 ;
        RECT 116.190 125.370 116.450 125.690 ;
        RECT 115.330 125.290 115.930 125.370 ;
        RECT 115.330 117.530 115.470 125.290 ;
        RECT 116.190 124.690 116.450 125.010 ;
        RECT 116.250 122.290 116.390 124.690 ;
        RECT 116.190 121.970 116.450 122.290 ;
        RECT 115.270 117.210 115.530 117.530 ;
        RECT 114.800 116.335 115.080 116.705 ;
        RECT 114.340 114.975 114.620 115.345 ;
        RECT 114.810 115.170 115.070 115.490 ;
        RECT 115.270 115.170 115.530 115.490 ;
        RECT 113.890 114.490 114.150 114.810 ;
        RECT 113.950 112.770 114.090 114.490 ;
        RECT 113.890 112.450 114.150 112.770 ;
        RECT 114.350 112.110 114.610 112.430 ;
        RECT 113.890 111.430 114.150 111.750 ;
        RECT 112.570 111.270 113.630 111.410 ;
        RECT 112.500 110.215 112.780 110.585 ;
        RECT 113.490 110.470 113.630 111.270 ;
        RECT 113.950 111.265 114.090 111.430 ;
        RECT 113.880 110.895 114.160 111.265 ;
        RECT 113.490 110.330 114.090 110.470 ;
        RECT 112.570 109.370 112.710 110.215 ;
        RECT 113.430 109.730 113.690 110.050 ;
        RECT 112.510 109.050 112.770 109.370 ;
        RECT 111.590 108.370 111.850 108.690 ;
        RECT 111.120 106.815 111.400 107.185 ;
        RECT 111.130 106.670 111.390 106.815 ;
        RECT 110.670 105.990 110.930 106.310 ;
        RECT 110.730 104.950 110.870 105.990 ;
        RECT 111.130 105.650 111.390 105.970 ;
        RECT 110.670 104.630 110.930 104.950 ;
        RECT 110.670 103.610 110.930 103.930 ;
        RECT 110.730 100.870 110.870 103.610 ;
        RECT 111.190 102.230 111.330 105.650 ;
        RECT 111.650 104.610 111.790 108.370 ;
        RECT 112.050 106.670 112.310 106.990 ;
        RECT 112.510 106.670 112.770 106.990 ;
        RECT 112.110 104.950 112.250 106.670 ;
        RECT 112.050 104.630 112.310 104.950 ;
        RECT 111.590 104.290 111.850 104.610 ;
        RECT 112.040 104.095 112.320 104.465 ;
        RECT 112.570 104.270 112.710 106.670 ;
        RECT 113.490 105.970 113.630 109.730 ;
        RECT 113.950 109.030 114.090 110.330 ;
        RECT 114.410 110.050 114.550 112.110 ;
        RECT 114.350 109.730 114.610 110.050 ;
        RECT 113.890 108.710 114.150 109.030 ;
        RECT 113.950 107.330 114.090 108.710 ;
        RECT 113.890 107.010 114.150 107.330 ;
        RECT 114.350 106.670 114.610 106.990 ;
        RECT 114.410 106.310 114.550 106.670 ;
        RECT 114.350 105.990 114.610 106.310 ;
        RECT 113.430 105.650 113.690 105.970 ;
        RECT 113.430 104.630 113.690 104.950 ;
        RECT 112.110 103.930 112.250 104.095 ;
        RECT 112.510 103.950 112.770 104.270 ;
        RECT 112.050 103.610 112.310 103.930 ;
        RECT 112.960 103.415 113.240 103.785 ;
        RECT 113.030 103.250 113.170 103.415 ;
        RECT 112.970 102.930 113.230 103.250 ;
        RECT 113.490 102.230 113.630 104.630 ;
        RECT 114.870 103.930 115.010 115.170 ;
        RECT 115.330 112.625 115.470 115.170 ;
        RECT 115.260 112.255 115.540 112.625 ;
        RECT 115.260 109.535 115.540 109.905 ;
        RECT 115.330 106.310 115.470 109.535 ;
        RECT 116.250 109.030 116.390 121.970 ;
        RECT 116.710 120.930 116.850 137.270 ;
        RECT 117.170 132.345 117.310 138.630 ;
        RECT 117.630 133.510 117.770 139.455 ;
        RECT 118.490 136.425 118.750 136.570 ;
        RECT 118.030 135.910 118.290 136.230 ;
        RECT 118.480 136.055 118.760 136.425 ;
        RECT 118.950 136.250 119.210 136.570 ;
        RECT 118.090 133.510 118.230 135.910 ;
        RECT 118.490 135.570 118.750 135.890 ;
        RECT 119.010 135.745 119.150 136.250 ;
        RECT 117.570 133.190 117.830 133.510 ;
        RECT 118.030 133.190 118.290 133.510 ;
        RECT 117.100 131.975 117.380 132.345 ;
        RECT 117.110 131.150 117.370 131.470 ;
        RECT 117.170 125.010 117.310 131.150 ;
        RECT 117.110 124.690 117.370 125.010 ;
        RECT 117.110 122.310 117.370 122.630 ;
        RECT 116.650 120.610 116.910 120.930 ;
        RECT 117.170 120.250 117.310 122.310 ;
        RECT 117.110 119.930 117.370 120.250 ;
        RECT 117.110 118.230 117.370 118.550 ;
        RECT 117.170 117.440 117.310 118.230 ;
        RECT 117.630 118.210 117.770 133.190 ;
        RECT 118.550 131.130 118.690 135.570 ;
        RECT 118.940 135.375 119.220 135.745 ;
        RECT 119.470 133.705 119.610 141.690 ;
        RECT 119.400 133.335 119.680 133.705 ;
        RECT 119.410 131.830 119.670 132.150 ;
        RECT 118.950 131.150 119.210 131.470 ;
        RECT 118.490 130.810 118.750 131.130 ;
        RECT 118.030 130.470 118.290 130.790 ;
        RECT 117.570 117.890 117.830 118.210 ;
        RECT 117.170 117.300 117.770 117.440 ;
        RECT 116.190 108.710 116.450 109.030 ;
        RECT 116.190 106.330 116.450 106.650 ;
        RECT 116.650 106.330 116.910 106.650 ;
        RECT 115.270 105.990 115.530 106.310 ;
        RECT 116.250 104.270 116.390 106.330 ;
        RECT 116.190 103.950 116.450 104.270 ;
        RECT 114.810 103.610 115.070 103.930 ;
        RECT 111.130 101.910 111.390 102.230 ;
        RECT 113.430 101.910 113.690 102.230 ;
        RECT 111.590 101.570 111.850 101.890 ;
        RECT 112.510 101.570 112.770 101.890 ;
        RECT 110.670 100.550 110.930 100.870 ;
        RECT 109.750 99.190 110.010 99.510 ;
        RECT 109.290 98.170 109.550 98.490 ;
        RECT 108.370 96.470 108.630 96.790 ;
        RECT 107.910 95.450 108.170 95.770 ;
        RECT 107.450 95.110 107.710 95.430 ;
        RECT 107.970 93.050 108.110 95.450 ;
        RECT 111.650 93.730 111.790 101.570 ;
        RECT 112.570 98.490 112.710 101.570 ;
        RECT 114.870 99.510 115.010 103.610 ;
        RECT 116.710 103.590 116.850 106.330 ;
        RECT 117.630 105.970 117.770 117.300 ;
        RECT 118.090 115.830 118.230 130.470 ;
        RECT 119.010 130.305 119.150 131.150 ;
        RECT 118.940 129.935 119.220 130.305 ;
        RECT 118.480 127.895 118.760 128.265 ;
        RECT 118.030 115.510 118.290 115.830 ;
        RECT 118.020 114.975 118.300 115.345 ;
        RECT 118.090 107.240 118.230 114.975 ;
        RECT 118.550 113.110 118.690 127.895 ;
        RECT 118.950 125.370 119.210 125.690 ;
        RECT 119.010 116.850 119.150 125.370 ;
        RECT 118.950 116.530 119.210 116.850 ;
        RECT 118.940 115.655 119.220 116.025 ;
        RECT 118.490 112.790 118.750 113.110 ;
        RECT 118.090 107.100 118.690 107.240 ;
        RECT 118.030 106.330 118.290 106.650 ;
        RECT 117.570 105.650 117.830 105.970 ;
        RECT 116.650 103.270 116.910 103.590 ;
        RECT 116.180 100.695 116.460 101.065 ;
        RECT 116.250 99.510 116.390 100.695 ;
        RECT 114.810 99.190 115.070 99.510 ;
        RECT 116.190 99.190 116.450 99.510 ;
        RECT 112.510 98.170 112.770 98.490 ;
        RECT 116.710 97.550 116.850 103.270 ;
        RECT 117.110 102.930 117.370 103.250 ;
        RECT 117.170 98.490 117.310 102.930 ;
        RECT 117.110 98.170 117.370 98.490 ;
        RECT 118.090 98.150 118.230 106.330 ;
        RECT 118.550 103.930 118.690 107.100 ;
        RECT 119.010 106.650 119.150 115.655 ;
        RECT 119.470 113.110 119.610 131.830 ;
        RECT 119.930 131.550 120.070 144.750 ;
        RECT 122.690 144.470 122.830 159.010 ;
        RECT 123.540 151.695 123.820 152.065 ;
        RECT 123.610 150.510 123.750 151.695 ;
        RECT 123.550 150.190 123.810 150.510 ;
        RECT 123.090 149.850 123.350 150.170 ;
        RECT 122.230 144.330 122.830 144.470 ;
        RECT 120.330 141.350 120.590 141.670 ;
        RECT 120.390 141.185 120.530 141.350 ;
        RECT 120.320 140.815 120.600 141.185 ;
        RECT 120.330 139.990 120.590 140.310 ;
        RECT 120.390 139.630 120.530 139.990 ;
        RECT 120.330 139.310 120.590 139.630 ;
        RECT 121.710 139.310 121.970 139.630 ;
        RECT 120.790 136.930 121.050 137.250 ;
        RECT 120.330 133.190 120.590 133.510 ;
        RECT 120.390 132.150 120.530 133.190 ;
        RECT 120.330 131.830 120.590 132.150 ;
        RECT 119.930 131.410 120.530 131.550 ;
        RECT 120.390 127.730 120.530 131.410 ;
        RECT 120.330 127.410 120.590 127.730 ;
        RECT 119.870 124.690 120.130 125.010 ;
        RECT 119.930 120.930 120.070 124.690 ;
        RECT 120.390 123.650 120.530 127.410 ;
        RECT 120.330 123.330 120.590 123.650 ;
        RECT 119.870 120.610 120.130 120.930 ;
        RECT 120.330 119.930 120.590 120.250 ;
        RECT 120.390 118.550 120.530 119.930 ;
        RECT 120.330 118.230 120.590 118.550 ;
        RECT 119.870 116.870 120.130 117.190 ;
        RECT 119.930 115.830 120.070 116.870 ;
        RECT 120.330 116.530 120.590 116.850 ;
        RECT 119.870 115.510 120.130 115.830 ;
        RECT 119.410 112.790 119.670 113.110 ;
        RECT 118.950 106.330 119.210 106.650 ;
        RECT 118.950 105.650 119.210 105.970 ;
        RECT 118.490 103.610 118.750 103.930 ;
        RECT 119.010 100.950 119.150 105.650 ;
        RECT 119.470 101.890 119.610 112.790 ;
        RECT 119.930 109.280 120.070 115.510 ;
        RECT 120.390 115.150 120.530 116.530 ;
        RECT 120.330 114.830 120.590 115.150 ;
        RECT 120.850 109.710 120.990 136.930 ;
        RECT 121.250 136.250 121.510 136.570 ;
        RECT 121.310 132.150 121.450 136.250 ;
        RECT 121.250 131.830 121.510 132.150 ;
        RECT 121.250 130.470 121.510 130.790 ;
        RECT 121.310 129.430 121.450 130.470 ;
        RECT 121.250 129.110 121.510 129.430 ;
        RECT 121.250 128.430 121.510 128.750 ;
        RECT 121.310 126.710 121.450 128.430 ;
        RECT 121.250 126.390 121.510 126.710 ;
        RECT 121.250 125.030 121.510 125.350 ;
        RECT 121.310 120.930 121.450 125.030 ;
        RECT 121.770 123.390 121.910 139.310 ;
        RECT 122.230 129.090 122.370 144.330 ;
        RECT 123.150 137.590 123.290 149.850 ;
        RECT 123.540 147.615 123.820 147.985 ;
        RECT 123.610 147.450 123.750 147.615 ;
        RECT 123.550 147.130 123.810 147.450 ;
        RECT 125.390 139.990 125.650 140.310 ;
        RECT 124.010 139.310 124.270 139.630 ;
        RECT 123.090 137.270 123.350 137.590 ;
        RECT 122.630 136.250 122.890 136.570 ;
        RECT 122.690 134.870 122.830 136.250 ;
        RECT 123.090 135.570 123.350 135.890 ;
        RECT 122.630 134.550 122.890 134.870 ;
        RECT 123.150 134.530 123.290 135.570 ;
        RECT 123.090 134.210 123.350 134.530 ;
        RECT 123.550 133.870 123.810 134.190 ;
        RECT 123.090 130.810 123.350 131.130 ;
        RECT 122.630 130.130 122.890 130.450 ;
        RECT 122.170 128.770 122.430 129.090 ;
        RECT 121.770 123.250 122.370 123.390 ;
        RECT 122.230 122.970 122.370 123.250 ;
        RECT 122.170 122.650 122.430 122.970 ;
        RECT 121.250 120.610 121.510 120.930 ;
        RECT 121.710 115.510 121.970 115.830 ;
        RECT 121.770 115.150 121.910 115.510 ;
        RECT 121.710 114.830 121.970 115.150 ;
        RECT 121.250 114.490 121.510 114.810 ;
        RECT 121.310 113.305 121.450 114.490 ;
        RECT 121.240 112.935 121.520 113.305 ;
        RECT 120.790 109.390 121.050 109.710 ;
        RECT 120.330 109.280 120.590 109.370 ;
        RECT 119.930 109.140 120.590 109.280 ;
        RECT 120.330 109.050 120.590 109.140 ;
        RECT 119.860 107.495 120.140 107.865 ;
        RECT 119.870 107.350 120.130 107.495 ;
        RECT 120.330 106.330 120.590 106.650 ;
        RECT 120.390 105.970 120.530 106.330 ;
        RECT 119.870 105.650 120.130 105.970 ;
        RECT 120.330 105.650 120.590 105.970 ;
        RECT 119.410 101.570 119.670 101.890 ;
        RECT 119.010 100.810 119.610 100.950 ;
        RECT 118.030 97.830 118.290 98.150 ;
        RECT 117.110 97.550 117.370 97.810 ;
        RECT 116.710 97.490 117.370 97.550 ;
        RECT 116.710 97.410 117.310 97.490 ;
        RECT 117.170 96.450 117.310 97.410 ;
        RECT 117.110 96.130 117.370 96.450 ;
        RECT 117.570 94.770 117.830 95.090 ;
        RECT 111.590 93.410 111.850 93.730 ;
        RECT 103.770 92.730 104.030 93.050 ;
        RECT 105.150 92.730 105.410 93.050 ;
        RECT 105.610 92.730 105.870 93.050 ;
        RECT 106.990 92.730 107.250 93.050 ;
        RECT 107.910 92.730 108.170 93.050 ;
        RECT 117.630 92.905 117.770 94.770 ;
        RECT 102.850 92.390 103.110 92.710 ;
        RECT 102.910 89.650 103.050 92.390 ;
        RECT 103.830 90.670 103.970 92.730 ;
        RECT 104.230 92.050 104.490 92.370 ;
        RECT 104.290 91.010 104.430 92.050 ;
        RECT 105.210 91.010 105.350 92.730 ;
        RECT 117.560 92.535 117.840 92.905 ;
        RECT 117.570 92.390 117.830 92.535 ;
        RECT 104.230 90.690 104.490 91.010 ;
        RECT 105.150 90.690 105.410 91.010 ;
        RECT 103.770 90.350 104.030 90.670 ;
        RECT 118.090 89.990 118.230 97.830 ;
        RECT 118.490 95.790 118.750 96.110 ;
        RECT 118.550 94.265 118.690 95.790 ;
        RECT 119.470 95.770 119.610 100.810 ;
        RECT 119.930 96.110 120.070 105.650 ;
        RECT 120.320 104.095 120.600 104.465 ;
        RECT 120.390 96.790 120.530 104.095 ;
        RECT 120.850 103.930 120.990 109.390 ;
        RECT 121.310 106.310 121.450 112.935 ;
        RECT 122.230 107.670 122.370 122.650 ;
        RECT 122.690 114.130 122.830 130.130 ;
        RECT 123.150 126.225 123.290 130.810 ;
        RECT 123.080 125.855 123.360 126.225 ;
        RECT 123.090 125.370 123.350 125.690 ;
        RECT 123.150 123.990 123.290 125.370 ;
        RECT 123.090 123.670 123.350 123.990 ;
        RECT 123.610 121.465 123.750 133.870 ;
        RECT 124.070 124.865 124.210 139.310 ;
        RECT 124.920 133.335 125.200 133.705 ;
        RECT 124.470 125.030 124.730 125.350 ;
        RECT 124.000 124.495 124.280 124.865 ;
        RECT 123.540 121.095 123.820 121.465 ;
        RECT 123.090 119.250 123.350 119.570 ;
        RECT 123.150 118.065 123.290 119.250 ;
        RECT 123.080 117.695 123.360 118.065 ;
        RECT 123.080 114.295 123.360 114.665 ;
        RECT 124.530 114.470 124.670 125.030 ;
        RECT 124.990 115.830 125.130 133.335 ;
        RECT 125.450 125.350 125.590 139.990 ;
        RECT 125.390 125.030 125.650 125.350 ;
        RECT 125.910 120.105 126.050 159.010 ;
        RECT 129.130 153.425 129.270 159.010 ;
        RECT 129.060 153.055 129.340 153.425 ;
        RECT 125.840 119.735 126.120 120.105 ;
        RECT 124.930 115.510 125.190 115.830 ;
        RECT 123.150 114.130 123.290 114.295 ;
        RECT 124.470 114.150 124.730 114.470 ;
        RECT 122.630 113.810 122.890 114.130 ;
        RECT 123.090 113.810 123.350 114.130 ;
        RECT 122.170 107.350 122.430 107.670 ;
        RECT 121.250 105.990 121.510 106.310 ;
        RECT 120.790 103.610 121.050 103.930 ;
        RECT 121.250 103.610 121.510 103.930 ;
        RECT 121.310 102.230 121.450 103.610 ;
        RECT 121.250 101.910 121.510 102.230 ;
        RECT 122.230 98.490 122.370 107.350 ;
        RECT 123.550 107.010 123.810 107.330 ;
        RECT 122.630 105.880 122.890 105.970 ;
        RECT 122.630 105.740 123.290 105.880 ;
        RECT 122.630 105.650 122.890 105.740 ;
        RECT 122.630 103.610 122.890 103.930 ;
        RECT 122.690 98.490 122.830 103.610 ;
        RECT 122.170 98.170 122.430 98.490 ;
        RECT 122.630 98.170 122.890 98.490 ;
        RECT 120.790 97.490 121.050 97.810 ;
        RECT 120.330 96.470 120.590 96.790 ;
        RECT 119.870 95.790 120.130 96.110 ;
        RECT 119.410 95.450 119.670 95.770 ;
        RECT 118.480 93.895 118.760 94.265 ;
        RECT 120.850 93.050 120.990 97.490 ;
        RECT 121.700 97.295 121.980 97.665 ;
        RECT 121.770 94.070 121.910 97.295 ;
        RECT 123.150 96.790 123.290 105.740 ;
        RECT 123.610 97.810 123.750 107.010 ;
        RECT 123.550 97.490 123.810 97.810 ;
        RECT 123.090 96.470 123.350 96.790 ;
        RECT 122.630 96.130 122.890 96.450 ;
        RECT 121.710 93.750 121.970 94.070 ;
        RECT 120.790 92.730 121.050 93.050 ;
        RECT 118.030 89.670 118.290 89.990 ;
        RECT 102.850 89.330 103.110 89.650 ;
        RECT 102.910 88.290 103.050 89.330 ;
        RECT 122.690 88.630 122.830 96.130 ;
        RECT 123.610 95.430 123.750 97.490 ;
        RECT 124.990 96.450 125.130 115.510 ;
        RECT 124.930 96.130 125.190 96.450 ;
        RECT 123.550 95.110 123.810 95.430 ;
        RECT 123.610 93.730 123.750 95.110 ;
        RECT 123.550 93.410 123.810 93.730 ;
        RECT 123.540 90.495 123.820 90.865 ;
        RECT 123.550 90.350 123.810 90.495 ;
        RECT 122.630 88.310 122.890 88.630 ;
        RECT 102.850 87.970 103.110 88.290 ;
        RECT 97.330 87.290 97.590 87.610 ;
        RECT 101.010 87.290 101.270 87.610 ;
        RECT 101.930 87.290 102.190 87.610 ;
        RECT 96.870 86.950 97.130 87.270 ;
        RECT 95.950 85.250 96.210 85.570 ;
        RECT 96.930 84.890 97.070 86.950 ;
        RECT 101.070 85.230 101.210 87.290 ;
        RECT 101.990 85.230 102.130 87.290 ;
        RECT 123.080 87.095 123.360 87.465 ;
        RECT 123.090 86.950 123.350 87.095 ;
        RECT 101.010 84.910 101.270 85.230 ;
        RECT 101.930 84.910 102.190 85.230 ;
        RECT 96.870 84.570 97.130 84.890 ;
        RECT 123.550 84.570 123.810 84.890 ;
        RECT 93.650 84.230 93.910 84.550 ;
        RECT 84.450 83.890 84.710 84.210 ;
        RECT 123.610 84.065 123.750 84.570 ;
        RECT 80.770 82.870 81.030 83.190 ;
        RECT 81.230 82.870 81.490 83.190 ;
        RECT 79.850 82.530 80.110 82.850 ;
        RECT 78.470 82.190 78.730 82.510 ;
        RECT 81.290 82.170 81.430 82.870 ;
        RECT 84.510 82.170 84.650 83.890 ;
        RECT 123.540 83.695 123.820 84.065 ;
        RECT 61.450 81.850 61.710 82.170 ;
        RECT 71.110 81.850 71.370 82.170 ;
        RECT 74.790 81.850 75.050 82.170 ;
        RECT 78.010 82.080 78.270 82.170 ;
        RECT 77.610 81.940 78.270 82.080 ;
        RECT 61.510 73.940 61.650 81.850 ;
        RECT 71.170 73.940 71.310 81.850 ;
        RECT 72.840 80.635 74.380 81.005 ;
        RECT 74.850 76.470 74.990 81.850 ;
        RECT 74.390 76.330 74.990 76.470 ;
        RECT 74.390 73.940 74.530 76.330 ;
        RECT 77.610 73.940 77.750 81.940 ;
        RECT 78.010 81.850 78.270 81.940 ;
        RECT 81.230 81.850 81.490 82.170 ;
        RECT 84.450 81.850 84.710 82.170 ;
        RECT 80.770 81.510 81.030 81.830 ;
        RECT 80.830 73.940 80.970 81.510 ;
        RECT 83.990 81.170 84.250 81.490 ;
        RECT 84.050 73.940 84.190 81.170 ;
        RECT 61.440 69.940 61.720 73.940 ;
        RECT 71.100 69.940 71.380 73.940 ;
        RECT 74.320 69.940 74.600 73.940 ;
        RECT 77.540 69.940 77.820 73.940 ;
        RECT 80.760 69.940 81.040 73.940 ;
        RECT 83.980 69.940 84.260 73.940 ;
      LAYER met3 ;
        RECT 67.140 162.230 67.520 162.240 ;
        RECT 126.820 162.230 130.820 162.380 ;
        RECT 67.140 161.930 130.820 162.230 ;
        RECT 67.140 161.920 67.520 161.930 ;
        RECT 126.820 161.780 130.820 161.930 ;
        RECT 58.655 158.830 58.985 158.845 ;
        RECT 126.820 158.830 130.820 158.980 ;
        RECT 58.655 158.530 130.820 158.830 ;
        RECT 58.655 158.515 58.985 158.530 ;
        RECT 126.820 158.380 130.820 158.530 ;
        RECT 54.260 158.150 54.640 158.160 ;
        RECT 112.935 158.150 113.265 158.165 ;
        RECT 54.260 157.850 113.265 158.150 ;
        RECT 54.260 157.840 54.640 157.850 ;
        RECT 112.935 157.835 113.265 157.850 ;
        RECT 48.535 156.110 48.865 156.125 ;
        RECT 62.540 156.110 62.920 156.120 ;
        RECT 48.535 155.810 62.920 156.110 ;
        RECT 48.535 155.795 48.865 155.810 ;
        RECT 62.540 155.800 62.920 155.810 ;
        RECT 100.055 156.110 100.385 156.125 ;
        RECT 115.695 156.110 116.025 156.125 ;
        RECT 100.055 155.810 116.025 156.110 ;
        RECT 100.055 155.795 100.385 155.810 ;
        RECT 115.695 155.795 116.025 155.810 ;
        RECT 78.180 155.430 78.560 155.440 ;
        RECT 103.275 155.430 103.605 155.445 ;
        RECT 78.180 155.130 103.605 155.430 ;
        RECT 78.180 155.120 78.560 155.130 ;
        RECT 103.275 155.115 103.605 155.130 ;
        RECT 104.655 155.430 104.985 155.445 ;
        RECT 126.820 155.430 130.820 155.580 ;
        RECT 104.655 155.130 130.820 155.430 ;
        RECT 104.655 155.115 104.985 155.130 ;
        RECT 126.820 154.980 130.820 155.130 ;
        RECT 67.395 154.070 67.725 154.085 ;
        RECT 87.175 154.070 87.505 154.085 ;
        RECT 67.395 153.770 87.505 154.070 ;
        RECT 67.395 153.755 67.725 153.770 ;
        RECT 87.175 153.755 87.505 153.770 ;
        RECT 94.740 154.070 95.120 154.080 ;
        RECT 119.375 154.070 119.705 154.085 ;
        RECT 94.740 153.770 119.705 154.070 ;
        RECT 94.740 153.760 95.120 153.770 ;
        RECT 119.375 153.755 119.705 153.770 ;
        RECT 58.860 153.390 59.240 153.400 ;
        RECT 61.415 153.390 61.745 153.405 ;
        RECT 58.860 153.090 61.745 153.390 ;
        RECT 58.860 153.080 59.240 153.090 ;
        RECT 61.415 153.075 61.745 153.090 ;
        RECT 66.015 153.390 66.345 153.405 ;
        RECT 80.940 153.390 81.320 153.400 ;
        RECT 66.015 153.090 81.320 153.390 ;
        RECT 66.015 153.075 66.345 153.090 ;
        RECT 80.940 153.080 81.320 153.090 ;
        RECT 91.980 153.390 92.360 153.400 ;
        RECT 109.715 153.390 110.045 153.405 ;
        RECT 129.035 153.390 129.365 153.405 ;
        RECT 91.980 153.090 110.045 153.390 ;
        RECT 91.980 153.080 92.360 153.090 ;
        RECT 109.715 153.075 110.045 153.090 ;
        RECT 110.420 153.090 129.365 153.390 ;
        RECT 56.815 152.710 57.145 152.725 ;
        RECT 75.675 152.710 76.005 152.725 ;
        RECT 56.815 152.410 76.005 152.710 ;
        RECT 56.815 152.395 57.145 152.410 ;
        RECT 75.675 152.395 76.005 152.410 ;
        RECT 92.235 152.710 92.565 152.725 ;
        RECT 110.420 152.710 110.720 153.090 ;
        RECT 129.035 153.075 129.365 153.090 ;
        RECT 92.235 152.410 110.720 152.710 ;
        RECT 92.235 152.395 92.565 152.410 ;
        RECT 48.470 152.030 52.470 152.180 ;
        RECT 53.595 152.030 53.925 152.045 ;
        RECT 48.470 151.730 53.925 152.030 ;
        RECT 48.470 151.580 52.470 151.730 ;
        RECT 53.595 151.715 53.925 151.730 ;
        RECT 93.615 152.030 93.945 152.045 ;
        RECT 123.515 152.030 123.845 152.045 ;
        RECT 126.820 152.030 130.820 152.180 ;
        RECT 93.615 151.730 123.845 152.030 ;
        RECT 93.615 151.715 93.945 151.730 ;
        RECT 123.515 151.715 123.845 151.730 ;
        RECT 124.220 151.730 130.820 152.030 ;
        RECT 72.820 151.375 74.400 151.705 ;
        RECT 59.115 151.350 59.445 151.365 ;
        RECT 71.075 151.350 71.405 151.365 ;
        RECT 59.115 151.050 71.405 151.350 ;
        RECT 59.115 151.035 59.445 151.050 ;
        RECT 71.075 151.035 71.405 151.050 ;
        RECT 74.755 151.350 75.085 151.365 ;
        RECT 107.875 151.350 108.205 151.365 ;
        RECT 74.755 151.050 108.205 151.350 ;
        RECT 74.755 151.035 75.085 151.050 ;
        RECT 107.875 151.035 108.205 151.050 ;
        RECT 114.980 151.350 115.360 151.360 ;
        RECT 124.220 151.350 124.520 151.730 ;
        RECT 126.820 151.580 130.820 151.730 ;
        RECT 114.980 151.050 124.520 151.350 ;
        RECT 114.980 151.040 115.360 151.050 ;
        RECT 66.475 150.670 66.805 150.685 ;
        RECT 117.995 150.670 118.325 150.685 ;
        RECT 66.475 150.370 118.325 150.670 ;
        RECT 66.475 150.355 66.805 150.370 ;
        RECT 117.995 150.355 118.325 150.370 ;
        RECT 60.700 149.990 61.080 150.000 ;
        RECT 61.875 149.990 62.205 150.005 ;
        RECT 69.695 149.990 70.025 150.005 ;
        RECT 73.375 149.990 73.705 150.005 ;
        RECT 60.700 149.690 62.205 149.990 ;
        RECT 60.700 149.680 61.080 149.690 ;
        RECT 61.875 149.675 62.205 149.690 ;
        RECT 63.500 149.690 73.705 149.990 ;
        RECT 48.470 148.630 52.470 148.780 ;
        RECT 54.975 148.630 55.305 148.645 ;
        RECT 48.470 148.330 55.305 148.630 ;
        RECT 48.470 148.180 52.470 148.330 ;
        RECT 54.975 148.315 55.305 148.330 ;
        RECT 57.275 147.270 57.605 147.285 ;
        RECT 63.500 147.280 63.800 149.690 ;
        RECT 69.695 149.675 70.025 149.690 ;
        RECT 73.375 149.675 73.705 149.690 ;
        RECT 74.295 149.990 74.625 150.005 ;
        RECT 79.815 149.990 80.145 150.005 ;
        RECT 118.915 149.990 119.245 150.005 ;
        RECT 74.295 149.690 119.245 149.990 ;
        RECT 74.295 149.675 74.625 149.690 ;
        RECT 79.815 149.675 80.145 149.690 ;
        RECT 118.915 149.675 119.245 149.690 ;
        RECT 121.420 149.990 121.800 150.000 ;
        RECT 122.135 149.990 122.465 150.005 ;
        RECT 121.420 149.690 122.465 149.990 ;
        RECT 121.420 149.680 121.800 149.690 ;
        RECT 122.135 149.675 122.465 149.690 ;
        RECT 73.835 149.310 74.165 149.325 ;
        RECT 78.895 149.310 79.225 149.325 ;
        RECT 73.835 149.010 79.225 149.310 ;
        RECT 73.835 148.995 74.165 149.010 ;
        RECT 78.895 148.995 79.225 149.010 ;
        RECT 92.900 149.310 93.280 149.320 ;
        RECT 94.075 149.310 94.405 149.325 ;
        RECT 115.235 149.310 115.565 149.325 ;
        RECT 92.900 149.010 115.565 149.310 ;
        RECT 92.900 149.000 93.280 149.010 ;
        RECT 94.075 148.995 94.405 149.010 ;
        RECT 115.235 148.995 115.565 149.010 ;
        RECT 69.520 148.655 71.100 148.985 ;
        RECT 82.115 148.630 82.445 148.645 ;
        RECT 113.140 148.630 113.520 148.640 ;
        RECT 126.820 148.630 130.820 148.780 ;
        RECT 71.780 148.330 96.920 148.630 ;
        RECT 64.175 147.950 64.505 147.965 ;
        RECT 71.780 147.950 72.080 148.330 ;
        RECT 82.115 148.315 82.445 148.330 ;
        RECT 64.175 147.650 72.080 147.950 ;
        RECT 73.375 147.950 73.705 147.965 ;
        RECT 82.780 147.950 83.160 147.960 ;
        RECT 73.375 147.650 83.160 147.950 ;
        RECT 96.620 147.950 96.920 148.330 ;
        RECT 113.140 148.330 130.820 148.630 ;
        RECT 113.140 148.320 113.520 148.330 ;
        RECT 126.820 148.180 130.820 148.330 ;
        RECT 123.515 147.950 123.845 147.965 ;
        RECT 96.620 147.650 123.845 147.950 ;
        RECT 64.175 147.635 64.505 147.650 ;
        RECT 73.375 147.635 73.705 147.650 ;
        RECT 82.780 147.640 83.160 147.650 ;
        RECT 123.515 147.635 123.845 147.650 ;
        RECT 63.460 147.270 63.840 147.280 ;
        RECT 57.275 146.970 63.840 147.270 ;
        RECT 57.275 146.955 57.605 146.970 ;
        RECT 63.460 146.960 63.840 146.970 ;
        RECT 65.095 147.270 65.425 147.285 ;
        RECT 103.735 147.270 104.065 147.285 ;
        RECT 65.095 146.970 104.065 147.270 ;
        RECT 65.095 146.955 65.425 146.970 ;
        RECT 103.735 146.955 104.065 146.970 ;
        RECT 107.875 147.270 108.205 147.285 ;
        RECT 117.075 147.270 117.405 147.285 ;
        RECT 107.875 146.970 117.405 147.270 ;
        RECT 107.875 146.955 108.205 146.970 ;
        RECT 117.075 146.955 117.405 146.970 ;
        RECT 61.875 146.590 62.205 146.605 ;
        RECT 65.110 146.590 65.410 146.955 ;
        RECT 61.875 146.290 65.410 146.590 ;
        RECT 66.015 146.590 66.345 146.605 ;
        RECT 75.215 146.600 75.545 146.605 ;
        RECT 71.740 146.590 72.120 146.600 ;
        RECT 66.015 146.290 72.120 146.590 ;
        RECT 61.875 146.275 62.205 146.290 ;
        RECT 66.015 146.275 66.345 146.290 ;
        RECT 71.740 146.280 72.120 146.290 ;
        RECT 75.215 146.590 75.800 146.600 ;
        RECT 90.140 146.590 90.520 146.600 ;
        RECT 91.315 146.590 91.645 146.605 ;
        RECT 75.215 146.290 76.000 146.590 ;
        RECT 90.140 146.290 91.645 146.590 ;
        RECT 75.215 146.280 75.800 146.290 ;
        RECT 90.140 146.280 90.520 146.290 ;
        RECT 75.215 146.275 75.545 146.280 ;
        RECT 91.315 146.275 91.645 146.290 ;
        RECT 105.115 146.590 105.445 146.605 ;
        RECT 105.780 146.590 106.160 146.600 ;
        RECT 105.115 146.290 106.160 146.590 ;
        RECT 105.115 146.275 105.445 146.290 ;
        RECT 105.780 146.280 106.160 146.290 ;
        RECT 107.620 146.590 108.000 146.600 ;
        RECT 120.755 146.590 121.085 146.605 ;
        RECT 107.620 146.290 121.085 146.590 ;
        RECT 107.620 146.280 108.000 146.290 ;
        RECT 120.755 146.275 121.085 146.290 ;
        RECT 72.820 145.935 74.400 146.265 ;
        RECT 61.415 145.910 61.745 145.925 ;
        RECT 71.995 145.910 72.325 145.925 ;
        RECT 61.415 145.610 72.325 145.910 ;
        RECT 61.415 145.595 61.745 145.610 ;
        RECT 71.995 145.595 72.325 145.610 ;
        RECT 74.755 145.910 75.085 145.925 ;
        RECT 93.155 145.910 93.485 145.925 ;
        RECT 74.755 145.610 109.800 145.910 ;
        RECT 74.755 145.595 75.085 145.610 ;
        RECT 93.155 145.595 93.485 145.610 ;
        RECT 48.470 145.230 52.470 145.380 ;
        RECT 54.515 145.230 54.845 145.245 ;
        RECT 48.470 144.930 54.845 145.230 ;
        RECT 48.470 144.780 52.470 144.930 ;
        RECT 54.515 144.915 54.845 144.930 ;
        RECT 63.715 145.230 64.045 145.245 ;
        RECT 66.475 145.230 66.805 145.245 ;
        RECT 104.860 145.230 105.240 145.240 ;
        RECT 107.875 145.230 108.205 145.245 ;
        RECT 63.715 144.930 66.805 145.230 ;
        RECT 63.715 144.915 64.045 144.930 ;
        RECT 66.475 144.915 66.805 144.930 ;
        RECT 68.100 144.930 108.205 145.230 ;
        RECT 109.500 145.230 109.800 145.610 ;
        RECT 110.175 145.230 110.505 145.245 ;
        RECT 109.500 144.930 110.505 145.230 ;
        RECT 63.255 143.870 63.585 143.885 ;
        RECT 68.100 143.870 68.400 144.930 ;
        RECT 104.860 144.920 105.240 144.930 ;
        RECT 107.875 144.915 108.205 144.930 ;
        RECT 110.175 144.915 110.505 144.930 ;
        RECT 114.060 145.230 114.440 145.240 ;
        RECT 126.820 145.230 130.820 145.380 ;
        RECT 114.060 144.930 130.820 145.230 ;
        RECT 114.060 144.920 114.440 144.930 ;
        RECT 126.820 144.780 130.820 144.930 ;
        RECT 69.695 144.550 70.025 144.565 ;
        RECT 77.260 144.550 77.640 144.560 ;
        RECT 69.695 144.250 77.640 144.550 ;
        RECT 69.695 144.235 70.025 144.250 ;
        RECT 77.260 144.240 77.640 144.250 ;
        RECT 78.435 144.550 78.765 144.565 ;
        RECT 92.900 144.550 93.280 144.560 ;
        RECT 78.435 144.250 93.280 144.550 ;
        RECT 78.435 144.235 78.765 144.250 ;
        RECT 92.900 144.240 93.280 144.250 ;
        RECT 94.995 144.550 95.325 144.565 ;
        RECT 95.660 144.550 96.040 144.560 ;
        RECT 94.995 144.250 96.040 144.550 ;
        RECT 94.995 144.235 95.325 144.250 ;
        RECT 95.660 144.240 96.040 144.250 ;
        RECT 63.255 143.570 68.400 143.870 ;
        RECT 72.455 143.870 72.785 143.885 ;
        RECT 80.020 143.870 80.400 143.880 ;
        RECT 72.455 143.570 80.400 143.870 ;
        RECT 63.255 143.555 63.585 143.570 ;
        RECT 72.455 143.555 72.785 143.570 ;
        RECT 80.020 143.560 80.400 143.570 ;
        RECT 82.575 143.870 82.905 143.885 ;
        RECT 88.300 143.870 88.680 143.880 ;
        RECT 108.795 143.870 109.125 143.885 ;
        RECT 82.575 143.570 109.125 143.870 ;
        RECT 82.575 143.555 82.905 143.570 ;
        RECT 88.300 143.560 88.680 143.570 ;
        RECT 108.795 143.555 109.125 143.570 ;
        RECT 69.520 143.215 71.100 143.545 ;
        RECT 59.575 143.190 59.905 143.205 ;
        RECT 60.700 143.190 61.080 143.200 ;
        RECT 59.575 142.890 61.080 143.190 ;
        RECT 59.575 142.875 59.905 142.890 ;
        RECT 60.700 142.880 61.080 142.890 ;
        RECT 62.335 143.190 62.665 143.205 ;
        RECT 67.855 143.190 68.185 143.205 ;
        RECT 62.335 142.890 68.185 143.190 ;
        RECT 62.335 142.875 62.665 142.890 ;
        RECT 67.855 142.875 68.185 142.890 ;
        RECT 71.995 143.190 72.325 143.205 ;
        RECT 74.295 143.190 74.625 143.205 ;
        RECT 76.340 143.190 76.720 143.200 ;
        RECT 71.995 142.890 76.720 143.190 ;
        RECT 71.995 142.875 72.325 142.890 ;
        RECT 74.295 142.875 74.625 142.890 ;
        RECT 76.340 142.880 76.720 142.890 ;
        RECT 78.435 143.190 78.765 143.205 ;
        RECT 101.180 143.190 101.560 143.200 ;
        RECT 101.895 143.190 102.225 143.205 ;
        RECT 78.435 142.890 102.225 143.190 ;
        RECT 78.435 142.875 78.765 142.890 ;
        RECT 101.180 142.880 101.560 142.890 ;
        RECT 101.895 142.875 102.225 142.890 ;
        RECT 109.460 143.190 109.840 143.200 ;
        RECT 111.555 143.190 111.885 143.205 ;
        RECT 109.460 142.890 111.885 143.190 ;
        RECT 109.460 142.880 109.840 142.890 ;
        RECT 111.555 142.875 111.885 142.890 ;
        RECT 64.380 142.510 64.760 142.520 ;
        RECT 68.775 142.510 69.105 142.525 ;
        RECT 64.380 142.210 69.105 142.510 ;
        RECT 64.380 142.200 64.760 142.210 ;
        RECT 68.775 142.195 69.105 142.210 ;
        RECT 69.695 142.510 70.025 142.525 ;
        RECT 88.095 142.510 88.425 142.525 ;
        RECT 69.695 142.210 88.425 142.510 ;
        RECT 69.695 142.195 70.025 142.210 ;
        RECT 88.095 142.195 88.425 142.210 ;
        RECT 48.470 141.830 52.470 141.980 ;
        RECT 53.595 141.830 53.925 141.845 ;
        RECT 48.470 141.530 53.925 141.830 ;
        RECT 48.470 141.380 52.470 141.530 ;
        RECT 53.595 141.515 53.925 141.530 ;
        RECT 60.955 141.830 61.285 141.845 ;
        RECT 71.535 141.830 71.865 141.845 ;
        RECT 81.860 141.830 82.240 141.840 ;
        RECT 60.955 141.530 67.710 141.830 ;
        RECT 60.955 141.515 61.285 141.530 ;
        RECT 62.335 141.150 62.665 141.165 ;
        RECT 66.220 141.150 66.600 141.160 ;
        RECT 62.335 140.850 66.600 141.150 ;
        RECT 67.410 141.150 67.710 141.530 ;
        RECT 71.535 141.530 82.240 141.830 ;
        RECT 71.535 141.515 71.865 141.530 ;
        RECT 81.860 141.520 82.240 141.530 ;
        RECT 91.060 141.830 91.440 141.840 ;
        RECT 95.455 141.830 95.785 141.845 ;
        RECT 91.060 141.530 95.785 141.830 ;
        RECT 91.060 141.520 91.440 141.530 ;
        RECT 95.455 141.515 95.785 141.530 ;
        RECT 111.300 141.830 111.680 141.840 ;
        RECT 126.820 141.830 130.820 141.980 ;
        RECT 111.300 141.530 130.820 141.830 ;
        RECT 111.300 141.520 111.680 141.530 ;
        RECT 126.820 141.380 130.820 141.530 ;
        RECT 71.995 141.150 72.325 141.165 ;
        RECT 67.410 140.850 72.325 141.150 ;
        RECT 62.335 140.835 62.665 140.850 ;
        RECT 66.220 140.840 66.600 140.850 ;
        RECT 71.995 140.835 72.325 140.850 ;
        RECT 75.675 141.150 76.005 141.165 ;
        RECT 96.580 141.150 96.960 141.160 ;
        RECT 107.415 141.150 107.745 141.165 ;
        RECT 75.675 140.850 107.745 141.150 ;
        RECT 75.675 140.835 76.005 140.850 ;
        RECT 96.580 140.840 96.960 140.850 ;
        RECT 107.415 140.835 107.745 140.850 ;
        RECT 118.660 141.150 119.040 141.160 ;
        RECT 120.295 141.150 120.625 141.165 ;
        RECT 118.660 140.850 120.625 141.150 ;
        RECT 118.660 140.840 119.040 140.850 ;
        RECT 120.295 140.835 120.625 140.850 ;
        RECT 72.820 140.495 74.400 140.825 ;
        RECT 60.700 140.470 61.080 140.480 ;
        RECT 63.715 140.470 64.045 140.485 ;
        RECT 60.700 140.170 64.045 140.470 ;
        RECT 60.700 140.160 61.080 140.170 ;
        RECT 63.715 140.155 64.045 140.170 ;
        RECT 68.060 140.470 68.440 140.480 ;
        RECT 70.155 140.470 70.485 140.485 ;
        RECT 68.060 140.170 70.485 140.470 ;
        RECT 68.060 140.160 68.440 140.170 ;
        RECT 70.155 140.155 70.485 140.170 ;
        RECT 74.755 140.470 75.085 140.485 ;
        RECT 87.635 140.470 87.965 140.485 ;
        RECT 74.755 140.170 87.965 140.470 ;
        RECT 74.755 140.155 75.085 140.170 ;
        RECT 87.635 140.155 87.965 140.170 ;
        RECT 93.615 140.470 93.945 140.485 ;
        RECT 116.615 140.470 116.945 140.485 ;
        RECT 93.615 140.170 116.945 140.470 ;
        RECT 93.615 140.155 93.945 140.170 ;
        RECT 116.615 140.155 116.945 140.170 ;
        RECT 67.395 139.790 67.725 139.805 ;
        RECT 69.235 139.790 69.565 139.805 ;
        RECT 74.770 139.790 75.070 140.155 ;
        RECT 67.395 139.490 75.070 139.790 ;
        RECT 83.035 139.790 83.365 139.805 ;
        RECT 117.535 139.790 117.865 139.805 ;
        RECT 83.035 139.490 117.865 139.790 ;
        RECT 67.395 139.475 67.725 139.490 ;
        RECT 69.235 139.475 69.565 139.490 ;
        RECT 83.035 139.475 83.365 139.490 ;
        RECT 117.535 139.475 117.865 139.490 ;
        RECT 76.340 139.110 76.720 139.120 ;
        RECT 77.515 139.110 77.845 139.125 ;
        RECT 68.100 138.810 72.080 139.110 ;
        RECT 48.470 138.430 52.470 138.580 ;
        RECT 55.895 138.430 56.225 138.445 ;
        RECT 48.470 138.130 56.225 138.430 ;
        RECT 48.470 137.980 52.470 138.130 ;
        RECT 55.895 138.115 56.225 138.130 ;
        RECT 62.795 137.750 63.125 137.765 ;
        RECT 63.715 137.750 64.045 137.765 ;
        RECT 68.100 137.750 68.400 138.810 ;
        RECT 71.780 138.430 72.080 138.810 ;
        RECT 76.340 138.810 77.845 139.110 ;
        RECT 76.340 138.800 76.720 138.810 ;
        RECT 77.515 138.795 77.845 138.810 ;
        RECT 78.895 139.120 79.225 139.125 ;
        RECT 78.895 139.110 79.480 139.120 ;
        RECT 80.275 139.110 80.605 139.125 ;
        RECT 94.535 139.110 94.865 139.125 ;
        RECT 78.895 138.810 79.680 139.110 ;
        RECT 80.275 138.810 94.865 139.110 ;
        RECT 78.895 138.800 79.480 138.810 ;
        RECT 78.895 138.795 79.225 138.800 ;
        RECT 80.275 138.795 80.605 138.810 ;
        RECT 94.535 138.795 94.865 138.810 ;
        RECT 102.815 139.120 103.145 139.125 ;
        RECT 102.815 139.110 103.400 139.120 ;
        RECT 102.815 138.810 103.600 139.110 ;
        RECT 102.815 138.800 103.400 138.810 ;
        RECT 102.815 138.795 103.145 138.800 ;
        RECT 84.875 138.430 85.205 138.445 ;
        RECT 96.375 138.430 96.705 138.445 ;
        RECT 71.780 138.130 79.440 138.430 ;
        RECT 69.520 137.775 71.100 138.105 ;
        RECT 62.795 137.450 68.400 137.750 ;
        RECT 71.995 137.750 72.325 137.765 ;
        RECT 75.215 137.750 75.545 137.765 ;
        RECT 76.595 137.760 76.925 137.765 ;
        RECT 76.340 137.750 76.925 137.760 ;
        RECT 71.995 137.450 75.545 137.750 ;
        RECT 76.140 137.450 76.925 137.750 ;
        RECT 62.795 137.435 63.125 137.450 ;
        RECT 63.715 137.435 64.045 137.450 ;
        RECT 71.995 137.435 72.325 137.450 ;
        RECT 75.215 137.435 75.545 137.450 ;
        RECT 76.340 137.440 76.925 137.450 ;
        RECT 76.595 137.435 76.925 137.440 ;
        RECT 66.475 137.070 66.805 137.085 ;
        RECT 78.180 137.070 78.560 137.080 ;
        RECT 66.475 136.770 78.560 137.070 ;
        RECT 79.140 137.070 79.440 138.130 ;
        RECT 84.875 138.130 96.705 138.430 ;
        RECT 84.875 138.115 85.205 138.130 ;
        RECT 96.375 138.115 96.705 138.130 ;
        RECT 102.100 138.430 102.480 138.440 ;
        RECT 104.655 138.430 104.985 138.445 ;
        RECT 126.820 138.430 130.820 138.580 ;
        RECT 102.100 138.130 104.985 138.430 ;
        RECT 102.100 138.120 102.480 138.130 ;
        RECT 104.655 138.115 104.985 138.130 ;
        RECT 110.420 138.130 130.820 138.430 ;
        RECT 89.015 137.750 89.345 137.765 ;
        RECT 110.420 137.750 110.720 138.130 ;
        RECT 126.820 137.980 130.820 138.130 ;
        RECT 89.015 137.450 110.720 137.750 ;
        RECT 89.015 137.435 89.345 137.450 ;
        RECT 105.115 137.070 105.445 137.085 ;
        RECT 79.140 136.770 105.445 137.070 ;
        RECT 66.475 136.755 66.805 136.770 ;
        RECT 78.180 136.760 78.560 136.770 ;
        RECT 105.115 136.755 105.445 136.770 ;
        RECT 61.620 136.390 62.000 136.400 ;
        RECT 64.635 136.390 64.965 136.405 ;
        RECT 67.395 136.400 67.725 136.405 ;
        RECT 67.140 136.390 67.725 136.400 ;
        RECT 75.675 136.390 76.005 136.405 ;
        RECT 61.620 136.090 64.965 136.390 ;
        RECT 66.940 136.090 67.725 136.390 ;
        RECT 61.620 136.080 62.000 136.090 ;
        RECT 64.635 136.075 64.965 136.090 ;
        RECT 67.140 136.080 67.725 136.090 ;
        RECT 67.395 136.075 67.725 136.080 ;
        RECT 72.010 136.090 76.005 136.390 ;
        RECT 60.495 135.710 60.825 135.725 ;
        RECT 72.010 135.710 72.310 136.090 ;
        RECT 75.675 136.075 76.005 136.090 ;
        RECT 78.180 136.390 78.560 136.400 ;
        RECT 79.815 136.390 80.145 136.405 ;
        RECT 78.180 136.090 80.145 136.390 ;
        RECT 78.180 136.080 78.560 136.090 ;
        RECT 79.815 136.075 80.145 136.090 ;
        RECT 82.115 136.390 82.445 136.405 ;
        RECT 86.255 136.390 86.585 136.405 ;
        RECT 82.115 136.090 86.585 136.390 ;
        RECT 82.115 136.075 82.445 136.090 ;
        RECT 86.255 136.075 86.585 136.090 ;
        RECT 95.660 136.390 96.040 136.400 ;
        RECT 118.455 136.390 118.785 136.405 ;
        RECT 95.660 136.090 118.785 136.390 ;
        RECT 95.660 136.080 96.040 136.090 ;
        RECT 118.455 136.075 118.785 136.090 ;
        RECT 60.495 135.410 72.310 135.710 ;
        RECT 78.895 135.710 79.225 135.725 ;
        RECT 83.700 135.710 84.080 135.720 ;
        RECT 118.915 135.710 119.245 135.725 ;
        RECT 78.895 135.410 119.245 135.710 ;
        RECT 60.495 135.395 60.825 135.410 ;
        RECT 78.895 135.395 79.225 135.410 ;
        RECT 83.700 135.400 84.080 135.410 ;
        RECT 118.915 135.395 119.245 135.410 ;
        RECT 48.470 135.030 52.470 135.180 ;
        RECT 72.820 135.055 74.400 135.385 ;
        RECT 53.135 135.030 53.465 135.045 ;
        RECT 48.470 134.730 53.465 135.030 ;
        RECT 48.470 134.580 52.470 134.730 ;
        RECT 53.135 134.715 53.465 134.730 ;
        RECT 61.415 135.030 61.745 135.045 ;
        RECT 69.695 135.030 70.025 135.045 ;
        RECT 61.415 134.730 70.025 135.030 ;
        RECT 61.415 134.715 61.745 134.730 ;
        RECT 69.695 134.715 70.025 134.730 ;
        RECT 83.035 135.030 83.365 135.045 ;
        RECT 91.315 135.030 91.645 135.045 ;
        RECT 83.035 134.730 91.645 135.030 ;
        RECT 83.035 134.715 83.365 134.730 ;
        RECT 91.315 134.715 91.645 134.730 ;
        RECT 111.555 135.030 111.885 135.045 ;
        RECT 126.820 135.030 130.820 135.180 ;
        RECT 111.555 134.730 130.820 135.030 ;
        RECT 111.555 134.715 111.885 134.730 ;
        RECT 126.820 134.580 130.820 134.730 ;
        RECT 69.235 134.350 69.565 134.365 ;
        RECT 85.335 134.350 85.665 134.365 ;
        RECT 69.235 134.050 85.665 134.350 ;
        RECT 69.235 134.035 69.565 134.050 ;
        RECT 85.335 134.035 85.665 134.050 ;
        RECT 67.395 133.670 67.725 133.685 ;
        RECT 71.075 133.670 71.405 133.685 ;
        RECT 67.395 133.370 71.405 133.670 ;
        RECT 67.395 133.355 67.725 133.370 ;
        RECT 71.075 133.355 71.405 133.370 ;
        RECT 75.215 133.670 75.545 133.685 ;
        RECT 119.375 133.670 119.705 133.685 ;
        RECT 124.895 133.670 125.225 133.685 ;
        RECT 75.215 133.370 125.225 133.670 ;
        RECT 75.215 133.355 75.545 133.370 ;
        RECT 119.375 133.355 119.705 133.370 ;
        RECT 124.895 133.355 125.225 133.370 ;
        RECT 64.380 132.990 64.760 133.000 ;
        RECT 68.775 132.990 69.105 133.005 ;
        RECT 73.375 132.990 73.705 133.005 ;
        RECT 64.380 132.690 69.105 132.990 ;
        RECT 64.380 132.680 64.760 132.690 ;
        RECT 68.775 132.675 69.105 132.690 ;
        RECT 71.550 132.690 73.705 132.990 ;
        RECT 69.520 132.335 71.100 132.665 ;
        RECT 52.675 132.310 53.005 132.325 ;
        RECT 52.460 131.995 53.005 132.310 ;
        RECT 66.015 132.310 66.345 132.325 ;
        RECT 68.315 132.310 68.645 132.325 ;
        RECT 66.015 132.010 68.645 132.310 ;
        RECT 66.015 131.995 66.345 132.010 ;
        RECT 68.315 131.995 68.645 132.010 ;
        RECT 52.460 131.780 52.760 131.995 ;
        RECT 48.470 131.330 52.760 131.780 ;
        RECT 64.635 131.640 64.965 131.645 ;
        RECT 64.380 131.630 64.965 131.640 ;
        RECT 64.180 131.330 64.965 131.630 ;
        RECT 48.470 131.180 52.470 131.330 ;
        RECT 64.380 131.320 64.965 131.330 ;
        RECT 65.300 131.630 65.680 131.640 ;
        RECT 71.550 131.630 71.850 132.690 ;
        RECT 73.375 132.675 73.705 132.690 ;
        RECT 76.340 132.990 76.720 133.000 ;
        RECT 89.935 132.990 90.265 133.005 ;
        RECT 99.135 132.990 99.465 133.005 ;
        RECT 76.340 132.690 90.265 132.990 ;
        RECT 76.340 132.680 76.720 132.690 ;
        RECT 89.935 132.675 90.265 132.690 ;
        RECT 96.850 132.690 99.465 132.990 ;
        RECT 96.850 132.325 97.150 132.690 ;
        RECT 99.135 132.675 99.465 132.690 ;
        RECT 112.475 132.990 112.805 133.005 ;
        RECT 114.980 132.990 115.360 133.000 ;
        RECT 112.475 132.690 115.360 132.990 ;
        RECT 112.475 132.675 112.805 132.690 ;
        RECT 114.980 132.680 115.360 132.690 ;
        RECT 73.375 132.310 73.705 132.325 ;
        RECT 83.495 132.310 83.825 132.325 ;
        RECT 73.375 132.010 83.825 132.310 ;
        RECT 89.015 132.140 89.345 132.155 ;
        RECT 73.375 131.995 73.705 132.010 ;
        RECT 83.495 131.995 83.825 132.010 ;
        RECT 88.340 131.840 89.345 132.140 ;
        RECT 96.835 131.995 97.165 132.325 ;
        RECT 97.755 132.310 98.085 132.325 ;
        RECT 101.435 132.310 101.765 132.325 ;
        RECT 97.755 132.010 101.765 132.310 ;
        RECT 97.755 131.995 98.085 132.010 ;
        RECT 101.435 131.995 101.765 132.010 ;
        RECT 106.035 132.310 106.365 132.325 ;
        RECT 117.075 132.310 117.405 132.325 ;
        RECT 106.035 132.010 117.405 132.310 ;
        RECT 106.035 131.995 106.365 132.010 ;
        RECT 117.075 131.995 117.405 132.010 ;
        RECT 65.300 131.330 71.850 131.630 ;
        RECT 72.915 131.630 73.245 131.645 ;
        RECT 88.340 131.630 88.640 131.840 ;
        RECT 89.015 131.825 89.345 131.840 ;
        RECT 72.915 131.330 88.640 131.630 ;
        RECT 89.935 131.630 90.265 131.645 ;
        RECT 126.820 131.630 130.820 131.780 ;
        RECT 89.935 131.330 130.820 131.630 ;
        RECT 65.300 131.320 65.680 131.330 ;
        RECT 64.635 131.315 64.965 131.320 ;
        RECT 72.915 131.315 73.245 131.330 ;
        RECT 89.935 131.315 90.265 131.330 ;
        RECT 126.820 131.180 130.820 131.330 ;
        RECT 60.955 130.950 61.285 130.965 ;
        RECT 69.695 130.950 70.025 130.965 ;
        RECT 60.955 130.650 70.025 130.950 ;
        RECT 60.955 130.635 61.285 130.650 ;
        RECT 69.695 130.635 70.025 130.650 ;
        RECT 73.835 130.950 74.165 130.965 ;
        RECT 91.060 130.950 91.440 130.960 ;
        RECT 111.300 130.950 111.680 130.960 ;
        RECT 73.835 130.650 91.440 130.950 ;
        RECT 73.835 130.635 74.165 130.650 ;
        RECT 91.060 130.640 91.440 130.650 ;
        RECT 99.380 130.650 111.680 130.950 ;
        RECT 67.140 130.270 67.520 130.280 ;
        RECT 70.155 130.270 70.485 130.285 ;
        RECT 79.815 130.280 80.145 130.285 ;
        RECT 79.815 130.270 80.400 130.280 ;
        RECT 88.555 130.270 88.885 130.285 ;
        RECT 67.140 129.970 70.485 130.270 ;
        RECT 79.590 129.970 80.400 130.270 ;
        RECT 67.140 129.960 67.520 129.970 ;
        RECT 70.155 129.955 70.485 129.970 ;
        RECT 79.815 129.960 80.400 129.970 ;
        RECT 81.210 129.970 88.885 130.270 ;
        RECT 79.815 129.955 80.145 129.960 ;
        RECT 72.820 129.615 74.400 129.945 ;
        RECT 52.675 129.600 53.005 129.605 ;
        RECT 52.420 129.590 53.005 129.600 ;
        RECT 52.220 129.290 53.005 129.590 ;
        RECT 52.420 129.280 53.005 129.290 ;
        RECT 52.675 129.275 53.005 129.280 ;
        RECT 58.655 129.590 58.985 129.605 ;
        RECT 62.335 129.590 62.665 129.605 ;
        RECT 58.655 129.290 62.665 129.590 ;
        RECT 58.655 129.275 58.985 129.290 ;
        RECT 62.335 129.275 62.665 129.290 ;
        RECT 67.855 129.275 68.185 129.605 ;
        RECT 71.075 129.590 71.405 129.605 ;
        RECT 71.995 129.590 72.325 129.605 ;
        RECT 71.075 129.290 72.325 129.590 ;
        RECT 71.075 129.275 71.405 129.290 ;
        RECT 71.995 129.275 72.325 129.290 ;
        RECT 78.895 129.590 79.225 129.605 ;
        RECT 81.210 129.590 81.510 129.970 ;
        RECT 88.555 129.955 88.885 129.970 ;
        RECT 93.820 130.270 94.200 130.280 ;
        RECT 99.380 130.270 99.680 130.650 ;
        RECT 111.300 130.640 111.680 130.650 ;
        RECT 118.915 130.270 119.245 130.285 ;
        RECT 93.820 129.970 99.680 130.270 ;
        RECT 110.420 129.970 119.245 130.270 ;
        RECT 93.820 129.960 94.200 129.970 ;
        RECT 78.895 129.290 81.510 129.590 ;
        RECT 82.780 129.590 83.160 129.600 ;
        RECT 84.875 129.590 85.205 129.605 ;
        RECT 82.780 129.290 85.205 129.590 ;
        RECT 78.895 129.275 79.225 129.290 ;
        RECT 82.780 129.280 83.160 129.290 ;
        RECT 84.875 129.275 85.205 129.290 ;
        RECT 87.635 129.590 87.965 129.605 ;
        RECT 89.220 129.590 89.600 129.600 ;
        RECT 110.420 129.590 110.720 129.970 ;
        RECT 118.915 129.955 119.245 129.970 ;
        RECT 87.635 129.290 110.720 129.590 ;
        RECT 87.635 129.275 87.965 129.290 ;
        RECT 89.220 129.280 89.600 129.290 ;
        RECT 67.870 128.910 68.170 129.275 ;
        RECT 75.675 128.910 76.005 128.925 ;
        RECT 67.870 128.610 76.005 128.910 ;
        RECT 75.675 128.595 76.005 128.610 ;
        RECT 82.575 128.910 82.905 128.925 ;
        RECT 85.335 128.910 85.665 128.925 ;
        RECT 99.135 128.910 99.465 128.925 ;
        RECT 82.575 128.610 84.960 128.910 ;
        RECT 82.575 128.595 82.905 128.610 ;
        RECT 48.470 128.240 52.470 128.380 ;
        RECT 48.470 127.920 52.800 128.240 ;
        RECT 67.855 128.230 68.185 128.245 ;
        RECT 77.975 128.230 78.305 128.245 ;
        RECT 67.855 127.930 78.305 128.230 ;
        RECT 48.470 127.780 52.470 127.920 ;
        RECT 67.855 127.915 68.185 127.930 ;
        RECT 77.975 127.915 78.305 127.930 ;
        RECT 84.660 127.560 84.960 128.610 ;
        RECT 85.335 128.610 99.465 128.910 ;
        RECT 85.335 128.595 85.665 128.610 ;
        RECT 99.135 128.595 99.465 128.610 ;
        RECT 87.380 128.230 87.760 128.240 ;
        RECT 89.015 128.230 89.345 128.245 ;
        RECT 87.380 127.930 89.345 128.230 ;
        RECT 87.380 127.920 87.760 127.930 ;
        RECT 89.015 127.915 89.345 127.930 ;
        RECT 91.315 128.230 91.645 128.245 ;
        RECT 92.900 128.230 93.280 128.240 ;
        RECT 91.315 127.930 93.280 128.230 ;
        RECT 91.315 127.915 91.645 127.930 ;
        RECT 92.900 127.920 93.280 127.930 ;
        RECT 118.455 128.230 118.785 128.245 ;
        RECT 126.820 128.230 130.820 128.380 ;
        RECT 118.455 127.930 130.820 128.230 ;
        RECT 118.455 127.915 118.785 127.930 ;
        RECT 126.820 127.780 130.820 127.930 ;
        RECT 84.620 127.550 85.000 127.560 ;
        RECT 92.235 127.550 92.565 127.565 ;
        RECT 98.215 127.550 98.545 127.565 ;
        RECT 84.620 127.250 98.545 127.550 ;
        RECT 84.620 127.240 85.000 127.250 ;
        RECT 92.235 127.235 92.565 127.250 ;
        RECT 98.215 127.235 98.545 127.250 ;
        RECT 69.520 126.895 71.100 127.225 ;
        RECT 61.620 126.870 62.000 126.880 ;
        RECT 67.855 126.870 68.185 126.885 ;
        RECT 77.055 126.870 77.385 126.885 ;
        RECT 61.620 126.570 68.185 126.870 ;
        RECT 61.620 126.560 62.000 126.570 ;
        RECT 67.855 126.555 68.185 126.570 ;
        RECT 73.850 126.570 77.385 126.870 ;
        RECT 73.850 126.205 74.150 126.570 ;
        RECT 77.055 126.555 77.385 126.570 ;
        RECT 78.180 126.870 78.560 126.880 ;
        RECT 81.655 126.870 81.985 126.885 ;
        RECT 78.180 126.570 81.985 126.870 ;
        RECT 78.180 126.560 78.560 126.570 ;
        RECT 81.655 126.555 81.985 126.570 ;
        RECT 97.295 126.870 97.625 126.885 ;
        RECT 112.935 126.870 113.265 126.885 ;
        RECT 97.295 126.570 113.265 126.870 ;
        RECT 97.295 126.555 97.625 126.570 ;
        RECT 112.935 126.555 113.265 126.570 ;
        RECT 63.255 126.190 63.585 126.205 ;
        RECT 66.015 126.190 66.345 126.205 ;
        RECT 69.235 126.190 69.565 126.205 ;
        RECT 63.255 125.890 65.640 126.190 ;
        RECT 63.255 125.875 63.585 125.890 ;
        RECT 62.540 125.510 62.920 125.520 ;
        RECT 63.715 125.510 64.045 125.525 ;
        RECT 62.540 125.210 64.045 125.510 ;
        RECT 65.340 125.510 65.640 125.890 ;
        RECT 66.015 125.890 69.565 126.190 ;
        RECT 66.015 125.875 66.345 125.890 ;
        RECT 69.235 125.875 69.565 125.890 ;
        RECT 70.155 126.190 70.485 126.205 ;
        RECT 71.740 126.190 72.120 126.200 ;
        RECT 70.155 125.890 72.120 126.190 ;
        RECT 70.155 125.875 70.485 125.890 ;
        RECT 71.740 125.880 72.120 125.890 ;
        RECT 73.835 125.875 74.165 126.205 ;
        RECT 83.495 126.190 83.825 126.205 ;
        RECT 123.055 126.190 123.385 126.205 ;
        RECT 83.495 125.890 123.385 126.190 ;
        RECT 83.495 125.875 83.825 125.890 ;
        RECT 123.055 125.875 123.385 125.890 ;
        RECT 69.695 125.510 70.025 125.525 ;
        RECT 65.340 125.210 70.025 125.510 ;
        RECT 62.540 125.200 62.920 125.210 ;
        RECT 63.715 125.195 64.045 125.210 ;
        RECT 69.695 125.195 70.025 125.210 ;
        RECT 79.355 125.510 79.685 125.525 ;
        RECT 85.335 125.510 85.665 125.525 ;
        RECT 90.855 125.510 91.185 125.525 ;
        RECT 92.235 125.520 92.565 125.525 ;
        RECT 91.980 125.510 92.565 125.520 ;
        RECT 112.475 125.510 112.805 125.525 ;
        RECT 79.355 125.210 91.185 125.510 ;
        RECT 91.780 125.210 92.565 125.510 ;
        RECT 79.355 125.195 79.685 125.210 ;
        RECT 85.335 125.195 85.665 125.210 ;
        RECT 90.855 125.195 91.185 125.210 ;
        RECT 91.980 125.200 92.565 125.210 ;
        RECT 92.235 125.195 92.565 125.200 ;
        RECT 99.380 125.210 112.805 125.510 ;
        RECT 48.470 124.830 52.470 124.980 ;
        RECT 55.435 124.830 55.765 124.845 ;
        RECT 48.470 124.530 55.765 124.830 ;
        RECT 48.470 124.380 52.470 124.530 ;
        RECT 55.435 124.515 55.765 124.530 ;
        RECT 58.860 124.830 59.240 124.840 ;
        RECT 65.095 124.830 65.425 124.845 ;
        RECT 58.860 124.530 65.425 124.830 ;
        RECT 58.860 124.520 59.240 124.530 ;
        RECT 65.095 124.515 65.425 124.530 ;
        RECT 67.140 124.830 67.520 124.840 ;
        RECT 71.535 124.830 71.865 124.845 ;
        RECT 67.140 124.530 71.865 124.830 ;
        RECT 67.140 124.520 67.520 124.530 ;
        RECT 71.535 124.515 71.865 124.530 ;
        RECT 79.815 124.830 80.145 124.845 ;
        RECT 80.940 124.830 81.320 124.840 ;
        RECT 79.815 124.530 81.320 124.830 ;
        RECT 79.815 124.515 80.145 124.530 ;
        RECT 80.940 124.520 81.320 124.530 ;
        RECT 81.860 124.830 82.240 124.840 ;
        RECT 85.335 124.830 85.665 124.845 ;
        RECT 81.860 124.530 85.665 124.830 ;
        RECT 81.860 124.520 82.240 124.530 ;
        RECT 85.335 124.515 85.665 124.530 ;
        RECT 89.015 124.830 89.345 124.845 ;
        RECT 99.380 124.830 99.680 125.210 ;
        RECT 112.475 125.195 112.805 125.210 ;
        RECT 89.015 124.530 99.680 124.830 ;
        RECT 123.975 124.830 124.305 124.845 ;
        RECT 126.820 124.830 130.820 124.980 ;
        RECT 123.975 124.530 130.820 124.830 ;
        RECT 89.015 124.515 89.345 124.530 ;
        RECT 123.975 124.515 124.305 124.530 ;
        RECT 72.820 124.175 74.400 124.505 ;
        RECT 126.820 124.380 130.820 124.530 ;
        RECT 60.700 124.150 61.080 124.160 ;
        RECT 61.875 124.150 62.205 124.165 ;
        RECT 60.700 123.850 62.205 124.150 ;
        RECT 60.700 123.840 61.080 123.850 ;
        RECT 61.875 123.835 62.205 123.850 ;
        RECT 63.460 124.150 63.840 124.160 ;
        RECT 66.015 124.150 66.345 124.165 ;
        RECT 63.460 123.850 66.345 124.150 ;
        RECT 63.460 123.840 63.840 123.850 ;
        RECT 66.015 123.835 66.345 123.850 ;
        RECT 68.315 124.150 68.645 124.165 ;
        RECT 71.740 124.150 72.120 124.160 ;
        RECT 68.315 123.850 72.120 124.150 ;
        RECT 68.315 123.835 68.645 123.850 ;
        RECT 71.740 123.840 72.120 123.850 ;
        RECT 80.735 124.150 81.065 124.165 ;
        RECT 94.075 124.150 94.405 124.165 ;
        RECT 80.735 123.850 94.405 124.150 ;
        RECT 80.735 123.835 81.065 123.850 ;
        RECT 94.075 123.835 94.405 123.850 ;
        RECT 103.020 124.150 103.400 124.160 ;
        RECT 111.300 124.150 111.680 124.160 ;
        RECT 103.020 123.850 111.680 124.150 ;
        RECT 103.020 123.840 103.400 123.850 ;
        RECT 111.300 123.840 111.680 123.850 ;
        RECT 58.655 123.470 58.985 123.485 ;
        RECT 90.140 123.470 90.520 123.480 ;
        RECT 58.655 123.170 90.520 123.470 ;
        RECT 58.655 123.155 58.985 123.170 ;
        RECT 90.140 123.160 90.520 123.170 ;
        RECT 97.295 123.470 97.625 123.485 ;
        RECT 99.340 123.470 99.720 123.480 ;
        RECT 100.515 123.470 100.845 123.485 ;
        RECT 97.295 123.170 100.845 123.470 ;
        RECT 97.295 123.155 97.625 123.170 ;
        RECT 99.340 123.160 99.720 123.170 ;
        RECT 100.515 123.155 100.845 123.170 ;
        RECT 105.115 123.470 105.445 123.485 ;
        RECT 107.620 123.470 108.000 123.480 ;
        RECT 105.115 123.170 108.000 123.470 ;
        RECT 105.115 123.155 105.445 123.170 ;
        RECT 107.620 123.160 108.000 123.170 ;
        RECT 51.755 122.790 52.085 122.805 ;
        RECT 63.715 122.790 64.045 122.805 ;
        RECT 51.755 122.490 64.045 122.790 ;
        RECT 51.755 122.475 52.085 122.490 ;
        RECT 63.715 122.475 64.045 122.490 ;
        RECT 64.380 122.790 64.760 122.800 ;
        RECT 67.855 122.790 68.185 122.805 ;
        RECT 64.380 122.490 68.185 122.790 ;
        RECT 64.380 122.480 64.760 122.490 ;
        RECT 67.855 122.475 68.185 122.490 ;
        RECT 68.775 122.790 69.105 122.805 ;
        RECT 78.435 122.790 78.765 122.805 ;
        RECT 68.775 122.490 78.765 122.790 ;
        RECT 68.775 122.475 69.105 122.490 ;
        RECT 78.435 122.475 78.765 122.490 ;
        RECT 80.275 122.790 80.605 122.805 ;
        RECT 85.335 122.790 85.665 122.805 ;
        RECT 80.275 122.490 85.665 122.790 ;
        RECT 80.275 122.475 80.605 122.490 ;
        RECT 85.335 122.475 85.665 122.490 ;
        RECT 90.855 122.790 91.185 122.805 ;
        RECT 91.775 122.790 92.105 122.805 ;
        RECT 90.855 122.490 92.105 122.790 ;
        RECT 90.855 122.475 91.185 122.490 ;
        RECT 91.775 122.475 92.105 122.490 ;
        RECT 63.715 122.110 64.045 122.125 ;
        RECT 65.300 122.110 65.680 122.120 ;
        RECT 63.715 121.810 65.680 122.110 ;
        RECT 63.715 121.795 64.045 121.810 ;
        RECT 65.300 121.800 65.680 121.810 ;
        RECT 71.740 122.110 72.120 122.120 ;
        RECT 85.795 122.110 86.125 122.125 ;
        RECT 88.555 122.120 88.885 122.125 ;
        RECT 71.740 121.810 86.125 122.110 ;
        RECT 71.740 121.800 72.120 121.810 ;
        RECT 85.795 121.795 86.125 121.810 ;
        RECT 88.300 122.110 88.885 122.120 ;
        RECT 88.300 121.810 89.110 122.110 ;
        RECT 88.300 121.800 88.885 121.810 ;
        RECT 88.555 121.795 88.885 121.800 ;
        RECT 69.520 121.455 71.100 121.785 ;
        RECT 73.375 121.430 73.705 121.445 ;
        RECT 74.755 121.430 75.085 121.445 ;
        RECT 77.055 121.430 77.385 121.445 ;
        RECT 85.795 121.430 86.125 121.445 ;
        RECT 73.375 121.130 86.125 121.430 ;
        RECT 73.375 121.115 73.705 121.130 ;
        RECT 74.755 121.115 75.085 121.130 ;
        RECT 77.055 121.115 77.385 121.130 ;
        RECT 85.795 121.115 86.125 121.130 ;
        RECT 91.775 121.430 92.105 121.445 ;
        RECT 97.295 121.430 97.625 121.445 ;
        RECT 91.775 121.130 97.625 121.430 ;
        RECT 91.775 121.115 92.105 121.130 ;
        RECT 97.295 121.115 97.625 121.130 ;
        RECT 123.515 121.430 123.845 121.445 ;
        RECT 126.820 121.430 130.820 121.580 ;
        RECT 123.515 121.130 130.820 121.430 ;
        RECT 123.515 121.115 123.845 121.130 ;
        RECT 126.820 120.980 130.820 121.130 ;
        RECT 76.340 120.750 76.720 120.760 ;
        RECT 77.975 120.750 78.305 120.765 ;
        RECT 84.415 120.750 84.745 120.765 ;
        RECT 76.340 120.450 84.745 120.750 ;
        RECT 76.340 120.440 76.720 120.450 ;
        RECT 77.975 120.435 78.305 120.450 ;
        RECT 84.415 120.435 84.745 120.450 ;
        RECT 91.775 120.750 92.105 120.765 ;
        RECT 95.660 120.750 96.040 120.760 ;
        RECT 91.775 120.450 96.040 120.750 ;
        RECT 91.775 120.435 92.105 120.450 ;
        RECT 95.660 120.440 96.040 120.450 ;
        RECT 96.835 120.750 97.165 120.765 ;
        RECT 107.415 120.750 107.745 120.765 ;
        RECT 96.835 120.450 107.745 120.750 ;
        RECT 96.835 120.435 97.165 120.450 ;
        RECT 107.415 120.435 107.745 120.450 ;
        RECT 64.175 120.070 64.505 120.085 ;
        RECT 77.260 120.070 77.640 120.080 ;
        RECT 64.175 119.770 77.640 120.070 ;
        RECT 64.175 119.755 64.505 119.770 ;
        RECT 77.260 119.760 77.640 119.770 ;
        RECT 78.895 120.070 79.225 120.085 ;
        RECT 89.015 120.070 89.345 120.085 ;
        RECT 78.895 119.770 89.345 120.070 ;
        RECT 78.895 119.755 79.225 119.770 ;
        RECT 89.015 119.755 89.345 119.770 ;
        RECT 94.535 120.070 94.865 120.085 ;
        RECT 101.895 120.070 102.225 120.085 ;
        RECT 94.535 119.770 102.225 120.070 ;
        RECT 94.535 119.755 94.865 119.770 ;
        RECT 101.895 119.755 102.225 119.770 ;
        RECT 103.020 120.070 103.400 120.080 ;
        RECT 125.815 120.070 126.145 120.085 ;
        RECT 103.020 119.770 126.145 120.070 ;
        RECT 103.020 119.760 103.400 119.770 ;
        RECT 125.815 119.755 126.145 119.770 ;
        RECT 84.875 119.390 85.205 119.405 ;
        RECT 91.060 119.390 91.440 119.400 ;
        RECT 92.900 119.390 93.280 119.400 ;
        RECT 106.700 119.390 107.080 119.400 ;
        RECT 84.875 119.090 107.080 119.390 ;
        RECT 84.875 119.075 85.205 119.090 ;
        RECT 91.060 119.080 91.440 119.090 ;
        RECT 92.900 119.080 93.280 119.090 ;
        RECT 106.700 119.080 107.080 119.090 ;
        RECT 72.820 118.735 74.400 119.065 ;
        RECT 74.755 118.710 75.085 118.725 ;
        RECT 84.415 118.710 84.745 118.725 ;
        RECT 86.715 118.720 87.045 118.725 ;
        RECT 86.460 118.710 87.045 118.720 ;
        RECT 89.015 118.720 89.345 118.725 ;
        RECT 89.015 118.710 89.600 118.720 ;
        RECT 74.755 118.410 84.745 118.710 ;
        RECT 86.260 118.410 87.045 118.710 ;
        RECT 88.790 118.410 89.600 118.710 ;
        RECT 74.755 118.395 75.085 118.410 ;
        RECT 84.415 118.395 84.745 118.410 ;
        RECT 86.460 118.400 87.045 118.410 ;
        RECT 86.715 118.395 87.045 118.400 ;
        RECT 89.015 118.400 89.600 118.410 ;
        RECT 89.935 118.710 90.265 118.725 ;
        RECT 91.980 118.710 92.360 118.720 ;
        RECT 94.535 118.710 94.865 118.725 ;
        RECT 89.935 118.410 94.865 118.710 ;
        RECT 89.015 118.395 89.345 118.400 ;
        RECT 89.935 118.395 90.265 118.410 ;
        RECT 91.980 118.400 92.360 118.410 ;
        RECT 94.535 118.395 94.865 118.410 ;
        RECT 96.375 118.395 96.705 118.725 ;
        RECT 104.195 118.710 104.525 118.725 ;
        RECT 114.060 118.710 114.440 118.720 ;
        RECT 104.195 118.410 114.440 118.710 ;
        RECT 104.195 118.395 104.525 118.410 ;
        RECT 114.060 118.400 114.440 118.410 ;
        RECT 48.470 118.030 52.470 118.180 ;
        RECT 96.390 118.045 96.690 118.395 ;
        RECT 55.435 118.030 55.765 118.045 ;
        RECT 48.470 117.730 55.765 118.030 ;
        RECT 48.470 117.580 52.470 117.730 ;
        RECT 55.435 117.715 55.765 117.730 ;
        RECT 76.595 118.030 76.925 118.045 ;
        RECT 83.035 118.030 83.365 118.045 ;
        RECT 76.595 117.730 83.365 118.030 ;
        RECT 76.595 117.715 76.925 117.730 ;
        RECT 83.035 117.715 83.365 117.730 ;
        RECT 83.700 118.030 84.080 118.040 ;
        RECT 89.935 118.030 90.265 118.045 ;
        RECT 83.700 117.730 90.265 118.030 ;
        RECT 83.700 117.720 84.080 117.730 ;
        RECT 89.935 117.715 90.265 117.730 ;
        RECT 94.535 118.040 94.865 118.045 ;
        RECT 94.535 118.030 95.120 118.040 ;
        RECT 94.535 117.730 95.320 118.030 ;
        RECT 94.535 117.720 95.120 117.730 ;
        RECT 94.535 117.715 94.865 117.720 ;
        RECT 96.375 117.715 96.705 118.045 ;
        RECT 103.735 118.030 104.065 118.045 ;
        RECT 105.575 118.040 105.905 118.045 ;
        RECT 104.860 118.030 105.240 118.040 ;
        RECT 103.735 117.730 105.240 118.030 ;
        RECT 103.735 117.715 104.065 117.730 ;
        RECT 104.860 117.720 105.240 117.730 ;
        RECT 105.575 118.030 106.160 118.040 ;
        RECT 123.055 118.030 123.385 118.045 ;
        RECT 126.820 118.030 130.820 118.180 ;
        RECT 105.575 117.730 106.360 118.030 ;
        RECT 123.055 117.730 130.820 118.030 ;
        RECT 105.575 117.720 106.160 117.730 ;
        RECT 105.575 117.715 105.905 117.720 ;
        RECT 123.055 117.715 123.385 117.730 ;
        RECT 126.820 117.580 130.820 117.730 ;
        RECT 68.060 117.350 68.440 117.360 ;
        RECT 79.100 117.350 79.480 117.360 ;
        RECT 86.255 117.350 86.585 117.365 ;
        RECT 68.060 117.050 78.750 117.350 ;
        RECT 68.060 117.040 68.440 117.050 ;
        RECT 78.450 116.670 78.750 117.050 ;
        RECT 79.100 117.050 86.585 117.350 ;
        RECT 79.100 117.040 79.480 117.050 ;
        RECT 86.255 117.035 86.585 117.050 ;
        RECT 89.015 117.350 89.345 117.365 ;
        RECT 93.820 117.350 94.200 117.360 ;
        RECT 89.015 117.050 94.200 117.350 ;
        RECT 89.015 117.035 89.345 117.050 ;
        RECT 93.820 117.040 94.200 117.050 ;
        RECT 95.455 117.350 95.785 117.365 ;
        RECT 113.855 117.350 114.185 117.365 ;
        RECT 95.455 117.050 114.185 117.350 ;
        RECT 95.455 117.035 95.785 117.050 ;
        RECT 113.855 117.035 114.185 117.050 ;
        RECT 86.715 116.670 87.045 116.685 ;
        RECT 114.775 116.670 115.105 116.685 ;
        RECT 78.450 116.370 87.045 116.670 ;
        RECT 86.715 116.355 87.045 116.370 ;
        RECT 101.220 116.370 115.105 116.670 ;
        RECT 69.520 116.015 71.100 116.345 ;
        RECT 75.420 115.990 75.800 116.000 ;
        RECT 97.755 115.990 98.085 116.005 ;
        RECT 75.420 115.690 98.085 115.990 ;
        RECT 75.420 115.680 75.800 115.690 ;
        RECT 97.755 115.675 98.085 115.690 ;
        RECT 66.220 115.310 66.600 115.320 ;
        RECT 85.335 115.310 85.665 115.325 ;
        RECT 100.515 115.310 100.845 115.325 ;
        RECT 66.220 115.010 100.845 115.310 ;
        RECT 66.220 115.000 66.600 115.010 ;
        RECT 85.335 114.995 85.665 115.010 ;
        RECT 100.515 114.995 100.845 115.010 ;
        RECT 54.260 114.630 54.640 114.640 ;
        RECT 89.475 114.630 89.805 114.645 ;
        RECT 93.155 114.640 93.485 114.645 ;
        RECT 54.260 114.330 89.805 114.630 ;
        RECT 54.260 114.320 54.640 114.330 ;
        RECT 89.475 114.315 89.805 114.330 ;
        RECT 92.900 114.630 93.485 114.640 ;
        RECT 94.075 114.630 94.405 114.645 ;
        RECT 99.135 114.640 99.465 114.645 ;
        RECT 96.580 114.630 96.960 114.640 ;
        RECT 92.900 114.330 93.710 114.630 ;
        RECT 94.075 114.330 96.960 114.630 ;
        RECT 92.900 114.320 93.485 114.330 ;
        RECT 93.155 114.315 93.485 114.320 ;
        RECT 94.075 114.315 94.405 114.330 ;
        RECT 96.580 114.320 96.960 114.330 ;
        RECT 99.135 114.630 99.720 114.640 ;
        RECT 99.135 114.330 99.920 114.630 ;
        RECT 99.135 114.320 99.720 114.330 ;
        RECT 99.135 114.315 99.465 114.320 ;
        RECT 84.415 113.960 84.745 113.965 ;
        RECT 87.175 113.960 87.505 113.965 ;
        RECT 92.235 113.960 92.565 113.965 ;
        RECT 84.415 113.950 85.000 113.960 ;
        RECT 87.175 113.950 87.760 113.960 ;
        RECT 91.980 113.950 92.565 113.960 ;
        RECT 84.190 113.650 85.000 113.950 ;
        RECT 86.950 113.650 87.760 113.950 ;
        RECT 91.780 113.650 92.565 113.950 ;
        RECT 84.415 113.640 85.000 113.650 ;
        RECT 87.175 113.640 87.760 113.650 ;
        RECT 91.980 113.640 92.565 113.650 ;
        RECT 84.415 113.635 84.745 113.640 ;
        RECT 87.175 113.635 87.505 113.640 ;
        RECT 92.235 113.635 92.565 113.640 ;
        RECT 95.915 113.950 96.245 113.965 ;
        RECT 101.220 113.950 101.520 116.370 ;
        RECT 114.775 116.355 115.105 116.370 ;
        RECT 118.915 115.990 119.245 116.005 ;
        RECT 110.420 115.690 119.245 115.990 ;
        RECT 102.355 114.630 102.685 114.645 ;
        RECT 103.020 114.630 103.400 114.640 ;
        RECT 110.420 114.630 110.720 115.690 ;
        RECT 118.915 115.675 119.245 115.690 ;
        RECT 114.315 115.310 114.645 115.325 ;
        RECT 117.995 115.310 118.325 115.325 ;
        RECT 118.660 115.310 119.040 115.320 ;
        RECT 114.315 115.010 119.040 115.310 ;
        RECT 114.315 114.995 114.645 115.010 ;
        RECT 117.995 114.995 118.325 115.010 ;
        RECT 118.660 115.000 119.040 115.010 ;
        RECT 102.355 114.330 103.400 114.630 ;
        RECT 102.355 114.315 102.685 114.330 ;
        RECT 103.020 114.320 103.400 114.330 ;
        RECT 104.900 114.330 110.720 114.630 ;
        RECT 123.055 114.630 123.385 114.645 ;
        RECT 126.820 114.630 130.820 114.780 ;
        RECT 123.055 114.330 130.820 114.630 ;
        RECT 95.915 113.650 101.520 113.950 ;
        RECT 102.100 113.950 102.480 113.960 ;
        RECT 103.735 113.950 104.065 113.965 ;
        RECT 102.100 113.650 104.065 113.950 ;
        RECT 95.915 113.635 96.245 113.650 ;
        RECT 102.100 113.640 102.480 113.650 ;
        RECT 103.735 113.635 104.065 113.650 ;
        RECT 72.820 113.295 74.400 113.625 ;
        RECT 80.940 113.270 81.320 113.280 ;
        RECT 83.035 113.270 83.365 113.285 ;
        RECT 86.715 113.280 87.045 113.285 ;
        RECT 80.940 112.970 83.365 113.270 ;
        RECT 80.940 112.960 81.320 112.970 ;
        RECT 83.035 112.955 83.365 112.970 ;
        RECT 86.460 113.270 87.045 113.280 ;
        RECT 87.635 113.270 87.965 113.285 ;
        RECT 89.475 113.270 89.805 113.285 ;
        RECT 86.460 112.970 87.270 113.270 ;
        RECT 87.635 112.970 89.805 113.270 ;
        RECT 86.460 112.960 87.045 112.970 ;
        RECT 86.715 112.955 87.045 112.960 ;
        RECT 87.635 112.955 87.965 112.970 ;
        RECT 89.475 112.955 89.805 112.970 ;
        RECT 101.180 113.270 101.560 113.280 ;
        RECT 102.815 113.270 103.145 113.285 ;
        RECT 101.180 112.970 103.145 113.270 ;
        RECT 101.180 112.960 101.560 112.970 ;
        RECT 102.815 112.955 103.145 112.970 ;
        RECT 68.315 112.590 68.645 112.605 ;
        RECT 75.215 112.590 75.545 112.605 ;
        RECT 68.315 112.290 75.545 112.590 ;
        RECT 68.315 112.275 68.645 112.290 ;
        RECT 75.215 112.275 75.545 112.290 ;
        RECT 82.575 112.590 82.905 112.605 ;
        RECT 87.635 112.590 87.965 112.605 ;
        RECT 82.575 112.290 87.965 112.590 ;
        RECT 82.575 112.275 82.905 112.290 ;
        RECT 87.635 112.275 87.965 112.290 ;
        RECT 98.215 112.590 98.545 112.605 ;
        RECT 100.975 112.590 101.305 112.605 ;
        RECT 104.900 112.590 105.200 114.330 ;
        RECT 123.055 114.315 123.385 114.330 ;
        RECT 126.820 114.180 130.820 114.330 ;
        RECT 106.035 113.950 106.365 113.965 ;
        RECT 107.620 113.950 108.000 113.960 ;
        RECT 106.035 113.650 108.000 113.950 ;
        RECT 106.035 113.635 106.365 113.650 ;
        RECT 107.620 113.640 108.000 113.650 ;
        RECT 106.700 113.270 107.080 113.280 ;
        RECT 121.215 113.270 121.545 113.285 ;
        RECT 106.700 112.970 121.545 113.270 ;
        RECT 106.700 112.960 107.080 112.970 ;
        RECT 121.215 112.955 121.545 112.970 ;
        RECT 98.215 112.290 105.200 112.590 ;
        RECT 107.875 112.590 108.205 112.605 ;
        RECT 115.235 112.590 115.565 112.605 ;
        RECT 107.875 112.290 115.565 112.590 ;
        RECT 98.215 112.275 98.545 112.290 ;
        RECT 100.975 112.275 101.305 112.290 ;
        RECT 107.875 112.275 108.205 112.290 ;
        RECT 115.235 112.275 115.565 112.290 ;
        RECT 56.355 111.910 56.685 111.925 ;
        RECT 112.935 111.910 113.265 111.925 ;
        RECT 56.355 111.610 113.265 111.910 ;
        RECT 56.355 111.595 56.685 111.610 ;
        RECT 112.935 111.595 113.265 111.610 ;
        RECT 83.035 111.230 83.365 111.245 ;
        RECT 90.855 111.230 91.185 111.245 ;
        RECT 83.035 110.930 91.185 111.230 ;
        RECT 83.035 110.915 83.365 110.930 ;
        RECT 90.855 110.915 91.185 110.930 ;
        RECT 101.435 111.230 101.765 111.245 ;
        RECT 105.115 111.230 105.445 111.245 ;
        RECT 101.435 110.930 105.445 111.230 ;
        RECT 101.435 110.915 101.765 110.930 ;
        RECT 105.115 110.915 105.445 110.930 ;
        RECT 113.855 111.230 114.185 111.245 ;
        RECT 126.820 111.230 130.820 111.380 ;
        RECT 113.855 110.930 130.820 111.230 ;
        RECT 113.855 110.915 114.185 110.930 ;
        RECT 69.520 110.575 71.100 110.905 ;
        RECT 126.820 110.780 130.820 110.930 ;
        RECT 98.675 110.550 99.005 110.565 ;
        RECT 112.475 110.550 112.805 110.565 ;
        RECT 98.675 110.250 112.805 110.550 ;
        RECT 98.675 110.235 99.005 110.250 ;
        RECT 112.475 110.235 112.805 110.250 ;
        RECT 66.935 109.870 67.265 109.885 ;
        RECT 78.435 109.870 78.765 109.885 ;
        RECT 66.935 109.570 78.765 109.870 ;
        RECT 66.935 109.555 67.265 109.570 ;
        RECT 78.435 109.555 78.765 109.570 ;
        RECT 102.815 109.870 103.145 109.885 ;
        RECT 115.235 109.870 115.565 109.885 ;
        RECT 102.815 109.570 115.565 109.870 ;
        RECT 102.815 109.555 103.145 109.570 ;
        RECT 115.235 109.555 115.565 109.570 ;
        RECT 73.375 109.190 73.705 109.205 ;
        RECT 74.755 109.190 75.085 109.205 ;
        RECT 83.035 109.190 83.365 109.205 ;
        RECT 73.375 108.890 83.365 109.190 ;
        RECT 73.375 108.875 73.705 108.890 ;
        RECT 74.755 108.875 75.085 108.890 ;
        RECT 83.035 108.875 83.365 108.890 ;
        RECT 72.820 107.855 74.400 108.185 ;
        RECT 119.835 107.830 120.165 107.845 ;
        RECT 126.820 107.830 130.820 107.980 ;
        RECT 119.835 107.530 130.820 107.830 ;
        RECT 119.835 107.515 120.165 107.530 ;
        RECT 126.820 107.380 130.820 107.530 ;
        RECT 63.255 107.150 63.585 107.165 ;
        RECT 68.315 107.150 68.645 107.165 ;
        RECT 106.955 107.150 107.285 107.165 ;
        RECT 111.095 107.150 111.425 107.165 ;
        RECT 63.255 106.850 111.425 107.150 ;
        RECT 63.255 106.835 63.585 106.850 ;
        RECT 68.315 106.835 68.645 106.850 ;
        RECT 106.955 106.835 107.285 106.850 ;
        RECT 111.095 106.835 111.425 106.850 ;
        RECT 107.875 106.470 108.205 106.485 ;
        RECT 109.460 106.470 109.840 106.480 ;
        RECT 107.875 106.170 109.840 106.470 ;
        RECT 107.875 106.155 108.205 106.170 ;
        RECT 109.460 106.160 109.840 106.170 ;
        RECT 69.520 105.135 71.100 105.465 ;
        RECT 111.300 104.430 111.680 104.440 ;
        RECT 112.015 104.430 112.345 104.445 ;
        RECT 111.300 104.130 112.345 104.430 ;
        RECT 111.300 104.120 111.680 104.130 ;
        RECT 112.015 104.115 112.345 104.130 ;
        RECT 120.295 104.430 120.625 104.445 ;
        RECT 126.820 104.430 130.820 104.580 ;
        RECT 120.295 104.130 130.820 104.430 ;
        RECT 120.295 104.115 120.625 104.130 ;
        RECT 126.820 103.980 130.820 104.130 ;
        RECT 112.935 103.760 113.265 103.765 ;
        RECT 112.935 103.750 113.520 103.760 ;
        RECT 112.710 103.450 113.520 103.750 ;
        RECT 112.935 103.440 113.520 103.450 ;
        RECT 112.935 103.435 113.265 103.440 ;
        RECT 72.820 102.415 74.400 102.745 ;
        RECT 83.955 101.710 84.285 101.725 ;
        RECT 85.795 101.710 86.125 101.725 ;
        RECT 83.955 101.410 86.125 101.710 ;
        RECT 83.955 101.395 84.285 101.410 ;
        RECT 85.795 101.395 86.125 101.410 ;
        RECT 48.470 101.030 52.470 101.180 ;
        RECT 55.895 101.030 56.225 101.045 ;
        RECT 48.470 100.730 56.225 101.030 ;
        RECT 48.470 100.580 52.470 100.730 ;
        RECT 55.895 100.715 56.225 100.730 ;
        RECT 79.355 101.030 79.685 101.045 ;
        RECT 83.955 101.030 84.285 101.045 ;
        RECT 79.355 100.730 84.285 101.030 ;
        RECT 79.355 100.715 79.685 100.730 ;
        RECT 83.955 100.715 84.285 100.730 ;
        RECT 116.155 101.030 116.485 101.045 ;
        RECT 126.820 101.030 130.820 101.180 ;
        RECT 116.155 100.730 130.820 101.030 ;
        RECT 116.155 100.715 116.485 100.730 ;
        RECT 126.820 100.580 130.820 100.730 ;
        RECT 69.520 99.695 71.100 100.025 ;
        RECT 83.035 99.670 83.365 99.685 ;
        RECT 85.795 99.670 86.125 99.685 ;
        RECT 83.035 99.370 86.125 99.670 ;
        RECT 83.035 99.355 83.365 99.370 ;
        RECT 85.795 99.355 86.125 99.370 ;
        RECT 48.470 97.630 52.470 97.780 ;
        RECT 57.735 97.630 58.065 97.645 ;
        RECT 48.470 97.330 58.065 97.630 ;
        RECT 48.470 97.180 52.470 97.330 ;
        RECT 57.735 97.315 58.065 97.330 ;
        RECT 121.675 97.630 122.005 97.645 ;
        RECT 126.820 97.630 130.820 97.780 ;
        RECT 121.675 97.330 130.820 97.630 ;
        RECT 121.675 97.315 122.005 97.330 ;
        RECT 72.820 96.975 74.400 97.305 ;
        RECT 126.820 97.180 130.820 97.330 ;
        RECT 55.435 94.910 55.765 94.925 ;
        RECT 52.460 94.610 55.765 94.910 ;
        RECT 52.460 94.380 52.760 94.610 ;
        RECT 55.435 94.595 55.765 94.610 ;
        RECT 48.470 93.930 52.760 94.380 ;
        RECT 69.520 94.255 71.100 94.585 ;
        RECT 118.455 94.230 118.785 94.245 ;
        RECT 126.820 94.230 130.820 94.380 ;
        RECT 118.455 93.930 130.820 94.230 ;
        RECT 48.470 93.780 52.470 93.930 ;
        RECT 118.455 93.915 118.785 93.930 ;
        RECT 126.820 93.780 130.820 93.930 ;
        RECT 76.595 92.870 76.925 92.885 ;
        RECT 117.535 92.870 117.865 92.885 ;
        RECT 76.595 92.570 117.865 92.870 ;
        RECT 76.595 92.555 76.925 92.570 ;
        RECT 117.535 92.555 117.865 92.570 ;
        RECT 72.820 91.535 74.400 91.865 ;
        RECT 48.470 90.830 52.470 90.980 ;
        RECT 123.515 90.830 123.845 90.845 ;
        RECT 126.820 90.830 130.820 90.980 ;
        RECT 48.470 90.380 52.760 90.830 ;
        RECT 123.515 90.530 130.820 90.830 ;
        RECT 123.515 90.515 123.845 90.530 ;
        RECT 126.820 90.380 130.820 90.530 ;
        RECT 52.460 90.150 52.760 90.380 ;
        RECT 55.895 90.150 56.225 90.165 ;
        RECT 52.460 89.850 56.225 90.150 ;
        RECT 55.895 89.835 56.225 89.850 ;
        RECT 69.520 88.815 71.100 89.145 ;
        RECT 123.055 87.430 123.385 87.445 ;
        RECT 126.820 87.430 130.820 87.580 ;
        RECT 123.055 87.130 130.820 87.430 ;
        RECT 123.055 87.115 123.385 87.130 ;
        RECT 126.820 86.980 130.820 87.130 ;
        RECT 72.820 86.095 74.400 86.425 ;
        RECT 123.515 84.030 123.845 84.045 ;
        RECT 126.820 84.030 130.820 84.180 ;
        RECT 123.515 83.730 130.820 84.030 ;
        RECT 123.515 83.715 123.845 83.730 ;
        RECT 69.520 83.375 71.100 83.705 ;
        RECT 126.820 83.580 130.820 83.730 ;
        RECT 72.820 80.655 74.400 80.985 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 67.165 161.915 67.495 162.245 ;
        RECT 54.285 157.835 54.615 158.165 ;
        RECT 52.445 129.275 52.775 129.605 ;
        RECT 52.460 128.245 52.760 129.275 ;
        RECT 52.445 127.915 52.775 128.245 ;
        RECT 54.300 114.645 54.600 157.835 ;
        RECT 62.565 155.795 62.895 156.125 ;
        RECT 58.885 153.075 59.215 153.405 ;
        RECT 58.900 124.845 59.200 153.075 ;
        RECT 60.300 149.250 61.480 150.430 ;
        RECT 60.300 142.450 61.480 143.630 ;
        RECT 60.725 140.155 61.055 140.485 ;
        RECT 58.885 124.515 59.215 124.845 ;
        RECT 60.740 124.165 61.040 140.155 ;
        RECT 61.645 136.075 61.975 136.405 ;
        RECT 61.660 126.885 61.960 136.075 ;
        RECT 61.645 126.555 61.975 126.885 ;
        RECT 62.580 125.525 62.880 155.795 ;
        RECT 63.485 146.955 63.815 147.285 ;
        RECT 62.565 125.195 62.895 125.525 ;
        RECT 63.500 124.165 63.800 146.955 ;
        RECT 64.405 142.195 64.735 142.525 ;
        RECT 64.420 133.005 64.720 142.195 ;
        RECT 66.245 140.835 66.575 141.165 ;
        RECT 66.260 133.430 66.560 140.835 ;
        RECT 67.180 136.405 67.480 161.915 ;
        RECT 78.205 155.115 78.535 155.445 ;
        RECT 68.085 140.155 68.415 140.485 ;
        RECT 67.165 136.075 67.495 136.405 ;
        RECT 64.405 132.675 64.735 133.005 ;
        RECT 65.820 132.250 67.000 133.430 ;
        RECT 64.405 131.315 64.735 131.645 ;
        RECT 65.325 131.315 65.655 131.645 ;
        RECT 60.725 123.835 61.055 124.165 ;
        RECT 63.485 123.835 63.815 124.165 ;
        RECT 64.420 122.805 64.720 131.315 ;
        RECT 64.405 122.475 64.735 122.805 ;
        RECT 65.340 122.125 65.640 131.315 ;
        RECT 65.325 121.795 65.655 122.125 ;
        RECT 66.260 115.325 66.560 132.250 ;
        RECT 67.165 129.955 67.495 130.285 ;
        RECT 67.180 124.845 67.480 129.955 ;
        RECT 67.165 124.515 67.495 124.845 ;
        RECT 68.100 117.365 68.400 140.155 ;
        RECT 68.085 117.035 68.415 117.365 ;
        RECT 66.245 114.995 66.575 115.325 ;
        RECT 54.285 114.315 54.615 114.645 ;
        RECT 69.510 80.580 71.110 151.780 ;
        RECT 71.765 146.275 72.095 146.605 ;
        RECT 71.780 126.205 72.080 146.275 ;
        RECT 71.765 125.875 72.095 126.205 ;
        RECT 71.765 123.835 72.095 124.165 ;
        RECT 71.780 122.125 72.080 123.835 ;
        RECT 71.765 121.795 72.095 122.125 ;
        RECT 72.810 80.580 74.410 151.780 ;
        RECT 75.445 146.275 75.775 146.605 ;
        RECT 75.460 116.005 75.760 146.275 ;
        RECT 77.285 144.235 77.615 144.565 ;
        RECT 76.365 142.875 76.695 143.205 ;
        RECT 76.380 139.125 76.680 142.875 ;
        RECT 76.365 138.795 76.695 139.125 ;
        RECT 76.365 137.435 76.695 137.765 ;
        RECT 76.380 133.005 76.680 137.435 ;
        RECT 76.365 132.675 76.695 133.005 ;
        RECT 76.380 120.765 76.680 132.675 ;
        RECT 76.365 120.435 76.695 120.765 ;
        RECT 77.300 120.085 77.600 144.235 ;
        RECT 78.220 137.085 78.520 155.115 ;
        RECT 94.765 153.755 95.095 154.085 ;
        RECT 80.965 153.075 81.295 153.405 ;
        RECT 92.005 153.075 92.335 153.405 ;
        RECT 80.045 143.555 80.375 143.885 ;
        RECT 79.125 138.795 79.455 139.125 ;
        RECT 78.205 136.755 78.535 137.085 ;
        RECT 78.205 136.075 78.535 136.405 ;
        RECT 78.220 126.885 78.520 136.075 ;
        RECT 78.205 126.555 78.535 126.885 ;
        RECT 77.285 119.755 77.615 120.085 ;
        RECT 79.140 117.365 79.440 138.795 ;
        RECT 80.060 130.285 80.360 143.555 ;
        RECT 80.045 129.955 80.375 130.285 ;
        RECT 80.980 124.845 81.280 153.075 ;
        RECT 82.805 147.635 83.135 147.965 ;
        RECT 81.885 141.515 82.215 141.845 ;
        RECT 81.900 124.845 82.200 141.515 ;
        RECT 82.820 129.605 83.120 147.635 ;
        RECT 90.165 146.275 90.495 146.605 ;
        RECT 88.325 143.555 88.655 143.885 ;
        RECT 83.725 135.395 84.055 135.725 ;
        RECT 82.805 129.275 83.135 129.605 ;
        RECT 80.965 124.515 81.295 124.845 ;
        RECT 81.885 124.515 82.215 124.845 ;
        RECT 79.125 117.035 79.455 117.365 ;
        RECT 75.445 115.675 75.775 116.005 ;
        RECT 80.980 113.285 81.280 124.515 ;
        RECT 83.740 118.045 84.040 135.395 ;
        RECT 87.405 127.915 87.735 128.245 ;
        RECT 84.645 127.235 84.975 127.565 ;
        RECT 83.725 117.715 84.055 118.045 ;
        RECT 84.660 113.965 84.960 127.235 ;
        RECT 86.485 118.395 86.815 118.725 ;
        RECT 84.645 113.635 84.975 113.965 ;
        RECT 86.500 113.285 86.800 118.395 ;
        RECT 87.420 113.965 87.720 127.915 ;
        RECT 88.340 122.125 88.640 143.555 ;
        RECT 89.245 129.275 89.575 129.605 ;
        RECT 88.325 121.795 88.655 122.125 ;
        RECT 89.260 118.725 89.560 129.275 ;
        RECT 90.180 123.485 90.480 146.275 ;
        RECT 91.085 141.515 91.415 141.845 ;
        RECT 91.100 130.965 91.400 141.515 ;
        RECT 91.085 130.635 91.415 130.965 ;
        RECT 90.165 123.155 90.495 123.485 ;
        RECT 91.100 119.405 91.400 130.635 ;
        RECT 92.020 125.525 92.320 153.075 ;
        RECT 92.925 148.995 93.255 149.325 ;
        RECT 92.940 144.565 93.240 148.995 ;
        RECT 92.925 144.235 93.255 144.565 ;
        RECT 92.940 128.245 93.240 144.235 ;
        RECT 93.845 129.955 94.175 130.285 ;
        RECT 92.925 127.915 93.255 128.245 ;
        RECT 92.005 125.195 92.335 125.525 ;
        RECT 91.085 119.075 91.415 119.405 ;
        RECT 92.925 119.075 93.255 119.405 ;
        RECT 89.245 118.395 89.575 118.725 ;
        RECT 92.005 118.395 92.335 118.725 ;
        RECT 92.020 113.965 92.320 118.395 ;
        RECT 92.940 114.645 93.240 119.075 ;
        RECT 93.860 117.365 94.160 129.955 ;
        RECT 94.780 118.045 95.080 153.755 ;
        RECT 115.005 151.035 115.335 151.365 ;
        RECT 113.165 148.315 113.495 148.645 ;
        RECT 105.805 146.275 106.135 146.605 ;
        RECT 107.645 146.275 107.975 146.605 ;
        RECT 104.885 144.915 105.215 145.245 ;
        RECT 95.685 144.235 96.015 144.565 ;
        RECT 95.700 136.405 96.000 144.235 ;
        RECT 101.205 142.875 101.535 143.205 ;
        RECT 96.605 140.835 96.935 141.165 ;
        RECT 95.685 136.075 96.015 136.405 ;
        RECT 95.700 120.765 96.000 136.075 ;
        RECT 95.685 120.435 96.015 120.765 ;
        RECT 94.765 117.715 95.095 118.045 ;
        RECT 93.845 117.035 94.175 117.365 ;
        RECT 96.620 114.645 96.920 140.835 ;
        RECT 99.365 123.155 99.695 123.485 ;
        RECT 99.380 114.645 99.680 123.155 ;
        RECT 92.925 114.315 93.255 114.645 ;
        RECT 96.605 114.315 96.935 114.645 ;
        RECT 99.365 114.315 99.695 114.645 ;
        RECT 87.405 113.635 87.735 113.965 ;
        RECT 92.005 113.635 92.335 113.965 ;
        RECT 101.220 113.285 101.520 142.875 ;
        RECT 103.045 138.795 103.375 139.125 ;
        RECT 102.125 138.115 102.455 138.445 ;
        RECT 102.140 113.965 102.440 138.115 ;
        RECT 103.060 124.165 103.360 138.795 ;
        RECT 103.045 123.835 103.375 124.165 ;
        RECT 103.045 119.755 103.375 120.085 ;
        RECT 103.060 114.645 103.360 119.755 ;
        RECT 104.900 118.045 105.200 144.915 ;
        RECT 105.820 118.045 106.120 146.275 ;
        RECT 107.660 133.430 107.960 146.275 ;
        RECT 109.060 142.450 110.240 143.630 ;
        RECT 107.220 132.250 108.400 133.430 ;
        RECT 107.645 123.155 107.975 123.485 ;
        RECT 106.725 119.075 107.055 119.405 ;
        RECT 104.885 117.715 105.215 118.045 ;
        RECT 105.805 117.715 106.135 118.045 ;
        RECT 103.045 114.315 103.375 114.645 ;
        RECT 102.125 113.635 102.455 113.965 ;
        RECT 106.740 113.285 107.040 119.075 ;
        RECT 107.660 113.965 107.960 123.155 ;
        RECT 107.645 113.635 107.975 113.965 ;
        RECT 80.965 112.955 81.295 113.285 ;
        RECT 86.485 112.955 86.815 113.285 ;
        RECT 101.205 112.955 101.535 113.285 ;
        RECT 106.725 112.955 107.055 113.285 ;
        RECT 109.500 106.485 109.800 142.450 ;
        RECT 111.325 141.515 111.655 141.845 ;
        RECT 111.340 130.965 111.640 141.515 ;
        RECT 111.325 130.635 111.655 130.965 ;
        RECT 111.325 123.835 111.655 124.165 ;
        RECT 109.485 106.155 109.815 106.485 ;
        RECT 111.340 104.445 111.640 123.835 ;
        RECT 111.325 104.115 111.655 104.445 ;
        RECT 113.180 103.765 113.480 148.315 ;
        RECT 114.085 144.915 114.415 145.245 ;
        RECT 114.100 118.725 114.400 144.915 ;
        RECT 115.020 133.005 115.320 151.035 ;
        RECT 121.020 149.250 122.200 150.430 ;
        RECT 118.685 140.835 119.015 141.165 ;
        RECT 115.005 132.675 115.335 133.005 ;
        RECT 114.085 118.395 114.415 118.725 ;
        RECT 118.700 115.325 119.000 140.835 ;
        RECT 118.685 114.995 119.015 115.325 ;
        RECT 113.165 103.435 113.495 103.765 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
      LAYER met5 ;
        RECT 60.090 149.040 122.410 150.640 ;
        RECT 60.090 142.240 110.450 143.840 ;
        RECT 65.610 132.040 108.610 133.640 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

