VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 23.645 194.785 23.815 194.975 ;
        RECT 26.405 194.785 26.575 194.975 ;
        RECT 27.785 194.805 27.955 194.975 ;
        RECT 28.245 194.785 28.415 194.975 ;
        RECT 33.765 194.785 33.935 194.975 ;
        RECT 36.980 194.835 37.100 194.945 ;
        RECT 40.205 194.785 40.375 194.975 ;
        RECT 40.665 194.785 40.835 194.975 ;
        RECT 46.185 194.785 46.355 194.975 ;
        RECT 48.940 194.835 49.060 194.945 ;
        RECT 49.865 194.785 50.035 194.975 ;
        RECT 55.385 194.785 55.555 194.975 ;
        RECT 60.905 194.785 61.075 194.975 ;
        RECT 62.755 194.830 62.915 194.940 ;
        RECT 63.675 194.785 63.845 194.975 ;
        RECT 65.045 194.785 65.215 194.975 ;
        RECT 68.265 194.785 68.435 194.975 ;
        RECT 68.725 194.785 68.895 194.975 ;
        RECT 72.415 194.830 72.575 194.940 ;
        RECT 73.335 194.785 73.505 194.975 ;
        RECT 74.700 194.835 74.820 194.945 ;
        RECT 75.635 194.830 75.795 194.940 ;
        RECT 77.455 194.785 77.625 194.975 ;
        RECT 77.925 194.785 78.095 194.975 ;
        RECT 79.315 194.785 79.485 194.975 ;
        RECT 81.145 194.825 81.315 194.975 ;
        RECT 23.505 193.975 24.875 194.785 ;
        RECT 24.885 194.105 26.715 194.785 ;
        RECT 24.885 193.875 26.230 194.105 ;
        RECT 28.105 193.975 33.615 194.785 ;
        RECT 33.625 193.975 36.375 194.785 ;
        RECT 36.395 193.915 36.825 194.700 ;
        RECT 37.305 193.875 40.515 194.785 ;
        RECT 40.525 193.975 46.035 194.785 ;
        RECT 46.045 193.975 48.795 194.785 ;
        RECT 49.275 193.915 49.705 194.700 ;
        RECT 49.725 193.975 55.235 194.785 ;
        RECT 55.245 193.975 60.755 194.785 ;
        RECT 60.765 193.975 62.135 194.785 ;
        RECT 62.155 193.915 62.585 194.700 ;
        RECT 63.525 194.005 64.895 194.785 ;
        RECT 64.905 193.975 66.735 194.785 ;
        RECT 66.745 194.105 68.575 194.785 ;
        RECT 66.745 193.875 68.090 194.105 ;
        RECT 68.585 193.975 72.255 194.785 ;
        RECT 73.185 194.005 74.555 194.785 ;
        RECT 75.035 193.915 75.465 194.700 ;
        RECT 76.405 194.005 77.775 194.785 ;
        RECT 77.785 193.975 79.155 194.785 ;
        RECT 79.165 194.005 80.535 194.785 ;
        RECT 80.545 193.875 81.435 194.825 ;
        RECT 81.615 194.785 81.785 194.975 ;
        RECT 82.960 194.805 83.130 194.975 ;
        RECT 87.580 194.835 87.700 194.945 ;
        RECT 83.020 194.785 83.130 194.805 ;
        RECT 88.505 194.785 88.675 194.975 ;
        RECT 90.355 194.830 90.515 194.940 ;
        RECT 91.265 194.785 91.435 194.975 ;
        RECT 92.645 194.785 92.815 194.975 ;
        RECT 94.495 194.785 94.665 194.975 ;
        RECT 96.775 194.785 96.945 194.975 ;
        RECT 97.240 194.835 97.360 194.945 ;
        RECT 97.715 194.785 97.885 194.975 ;
        RECT 100.465 194.785 100.635 194.975 ;
        RECT 101.395 194.830 101.555 194.940 ;
        RECT 103.685 194.785 103.855 194.975 ;
        RECT 105.055 194.785 105.225 194.975 ;
        RECT 106.905 194.785 107.075 194.975 ;
        RECT 108.285 194.785 108.455 194.975 ;
        RECT 108.740 194.835 108.860 194.945 ;
        RECT 111.045 194.805 111.215 194.975 ;
        RECT 111.505 194.805 111.675 194.975 ;
        RECT 114.275 194.830 114.435 194.940 ;
        RECT 111.045 194.785 111.210 194.805 ;
        RECT 81.465 194.005 82.835 194.785 ;
        RECT 83.020 194.105 87.435 194.785 ;
        RECT 83.505 193.875 87.435 194.105 ;
        RECT 87.915 193.915 88.345 194.700 ;
        RECT 88.365 194.105 90.195 194.785 ;
        RECT 88.850 193.875 90.195 194.105 ;
        RECT 91.125 194.005 92.495 194.785 ;
        RECT 92.505 194.105 94.335 194.785 ;
        RECT 92.990 193.875 94.335 194.105 ;
        RECT 94.345 194.005 95.715 194.785 ;
        RECT 95.725 194.005 97.095 194.785 ;
        RECT 97.565 194.005 98.935 194.785 ;
        RECT 98.945 194.105 100.775 194.785 ;
        RECT 98.945 193.875 100.290 194.105 ;
        RECT 100.795 193.915 101.225 194.700 ;
        RECT 102.165 194.105 103.995 194.785 ;
        RECT 102.165 193.875 103.510 194.105 ;
        RECT 104.005 194.005 105.375 194.785 ;
        RECT 105.385 194.105 107.215 194.785 ;
        RECT 105.385 193.875 106.730 194.105 ;
        RECT 107.225 194.005 108.595 194.785 ;
        RECT 109.375 194.105 111.210 194.785 ;
        RECT 111.525 194.785 111.675 194.805 ;
        RECT 116.565 194.785 116.735 194.975 ;
        RECT 117.025 194.805 117.195 194.975 ;
        RECT 117.055 194.785 117.195 194.805 ;
        RECT 120.705 194.785 120.875 194.975 ;
        RECT 122.085 194.785 122.255 194.975 ;
        RECT 123.455 194.785 123.625 194.975 ;
        RECT 126.225 194.785 126.395 194.975 ;
        RECT 127.145 194.785 127.315 194.975 ;
        RECT 128.980 194.835 129.100 194.945 ;
        RECT 132.205 194.785 132.375 194.975 ;
        RECT 132.665 194.785 132.835 194.975 ;
        RECT 135.885 194.785 136.055 194.975 ;
        RECT 109.375 193.875 110.305 194.105 ;
        RECT 111.525 193.965 113.455 194.785 ;
        RECT 112.505 193.875 113.455 193.965 ;
        RECT 113.675 193.915 114.105 194.700 ;
        RECT 115.045 194.105 116.875 194.785 ;
        RECT 115.045 193.875 116.390 194.105 ;
        RECT 117.055 193.965 119.625 194.785 ;
        RECT 118.035 193.875 119.625 193.965 ;
        RECT 119.655 193.875 121.005 194.785 ;
        RECT 121.025 194.005 122.395 194.785 ;
        RECT 122.405 194.005 123.775 194.785 ;
        RECT 123.785 193.875 126.535 194.785 ;
        RECT 126.555 193.915 126.985 194.700 ;
        RECT 127.005 194.105 128.835 194.785 ;
        RECT 127.490 193.875 128.835 194.105 ;
        RECT 129.435 193.875 132.435 194.785 ;
        RECT 132.525 193.875 134.815 194.785 ;
        RECT 134.825 193.975 136.195 194.785 ;
      LAYER nwell ;
        RECT 23.310 190.755 136.390 193.585 ;
      LAYER pwell ;
        RECT 23.505 189.555 24.875 190.365 ;
        RECT 24.885 190.235 26.230 190.465 ;
        RECT 24.885 189.555 26.715 190.235 ;
        RECT 27.645 189.555 29.015 190.335 ;
        RECT 29.025 189.555 34.535 190.365 ;
        RECT 34.545 189.555 36.375 190.365 ;
        RECT 36.395 189.640 36.825 190.425 ;
        RECT 36.845 189.555 38.215 190.365 ;
        RECT 38.225 190.235 39.155 190.465 ;
        RECT 42.675 190.235 43.605 190.465 ;
        RECT 38.225 189.555 42.125 190.235 ;
        RECT 42.675 189.555 44.510 190.235 ;
        RECT 44.665 189.555 46.495 190.365 ;
        RECT 46.965 189.555 48.780 190.465 ;
        RECT 48.820 189.555 50.635 190.465 ;
        RECT 50.645 189.555 53.855 190.465 ;
        RECT 53.865 190.235 54.795 190.465 ;
        RECT 53.865 189.555 57.765 190.235 ;
        RECT 58.005 189.555 59.835 190.235 ;
        RECT 59.845 189.555 61.675 190.365 ;
        RECT 62.155 189.640 62.585 190.425 ;
        RECT 62.605 189.555 63.975 190.365 ;
        RECT 63.985 190.235 65.330 190.465 ;
        RECT 63.985 189.555 65.815 190.235 ;
        RECT 65.825 189.555 67.640 190.465 ;
        RECT 67.665 189.555 69.035 190.335 ;
        RECT 69.045 189.555 72.255 190.465 ;
        RECT 72.265 189.555 73.635 190.365 ;
        RECT 73.645 190.235 74.570 190.465 ;
        RECT 77.635 190.235 78.565 190.465 ;
        RECT 73.645 189.555 77.315 190.235 ;
        RECT 77.635 189.555 79.470 190.235 ;
        RECT 79.625 189.555 82.375 190.365 ;
        RECT 82.485 189.555 84.675 190.465 ;
        RECT 85.155 189.555 86.505 190.465 ;
        RECT 86.525 189.555 87.895 190.335 ;
        RECT 87.915 189.640 88.345 190.425 ;
        RECT 90.425 190.375 91.375 190.465 ;
        RECT 89.445 189.555 91.375 190.375 ;
        RECT 91.895 190.235 92.825 190.465 ;
        RECT 95.485 190.375 96.435 190.465 ;
        RECT 91.895 189.555 93.730 190.235 ;
        RECT 23.645 189.345 23.815 189.555 ;
        RECT 25.025 189.345 25.195 189.535 ;
        RECT 26.405 189.365 26.575 189.555 ;
        RECT 26.875 189.400 27.035 189.510 ;
        RECT 28.705 189.345 28.875 189.555 ;
        RECT 29.165 189.345 29.335 189.555 ;
        RECT 34.685 189.345 34.855 189.555 ;
        RECT 36.985 189.365 37.155 189.555 ;
        RECT 37.440 189.395 37.560 189.505 ;
        RECT 38.180 189.345 38.350 189.535 ;
        RECT 38.640 189.365 38.810 189.555 ;
        RECT 44.345 189.535 44.510 189.555 ;
        RECT 42.045 189.345 42.215 189.535 ;
        RECT 44.345 189.365 44.515 189.535 ;
        RECT 44.805 189.365 44.975 189.555 ;
        RECT 46.640 189.395 46.760 189.505 ;
        RECT 47.105 189.365 47.275 189.535 ;
        RECT 48.485 189.365 48.655 189.555 ;
        RECT 48.945 189.365 49.115 189.555 ;
        RECT 49.875 189.390 50.035 189.500 ;
        RECT 44.810 189.345 44.975 189.365 ;
        RECT 47.110 189.345 47.275 189.365 ;
        RECT 50.785 189.345 50.955 189.555 ;
        RECT 54.280 189.345 54.450 189.555 ;
        RECT 58.420 189.345 58.590 189.535 ;
        RECT 59.525 189.365 59.695 189.555 ;
        RECT 59.985 189.365 60.155 189.555 ;
        RECT 61.820 189.395 61.940 189.505 ;
        RECT 62.280 189.395 62.400 189.505 ;
        RECT 62.745 189.365 62.915 189.555 ;
        RECT 63.670 189.345 63.840 189.535 ;
        RECT 64.135 189.390 64.295 189.500 ;
        RECT 65.505 189.365 65.675 189.555 ;
        RECT 67.345 189.345 67.515 189.555 ;
        RECT 67.810 189.345 67.980 189.535 ;
        RECT 68.725 189.365 68.895 189.555 ;
        RECT 71.940 189.365 72.110 189.555 ;
        RECT 72.405 189.345 72.575 189.555 ;
        RECT 73.790 189.365 73.960 189.555 ;
        RECT 79.305 189.535 79.470 189.555 ;
        RECT 75.625 189.345 75.795 189.535 ;
        RECT 78.660 189.345 78.830 189.535 ;
        RECT 79.305 189.365 79.475 189.535 ;
        RECT 79.765 189.365 79.935 189.555 ;
        RECT 82.800 189.345 82.970 189.535 ;
        RECT 84.360 189.365 84.530 189.555 ;
        RECT 84.820 189.395 84.940 189.505 ;
        RECT 85.285 189.365 85.455 189.555 ;
        RECT 86.665 189.345 86.835 189.555 ;
        RECT 89.445 189.535 89.595 189.555 ;
        RECT 88.505 189.345 88.675 189.535 ;
        RECT 89.425 189.365 89.595 189.535 ;
        RECT 93.565 189.535 93.730 189.555 ;
        RECT 94.505 189.555 96.435 190.375 ;
        RECT 96.655 189.555 98.005 190.465 ;
        RECT 98.045 189.555 99.395 190.465 ;
        RECT 99.405 189.555 100.775 190.335 ;
        RECT 102.085 189.555 107.215 190.465 ;
        RECT 107.225 189.555 109.415 190.465 ;
        RECT 109.725 190.375 110.675 190.465 ;
        RECT 109.725 189.555 111.655 190.375 ;
        RECT 111.825 189.555 113.195 190.335 ;
        RECT 113.675 189.640 114.105 190.425 ;
        RECT 114.135 190.375 115.725 190.465 ;
        RECT 114.135 189.555 116.705 190.375 ;
        RECT 127.950 190.235 129.295 190.465 ;
        RECT 117.805 189.555 126.910 190.235 ;
        RECT 127.465 189.555 129.295 190.235 ;
        RECT 129.385 189.555 132.835 190.465 ;
        RECT 133.000 189.555 134.815 190.465 ;
        RECT 134.825 189.555 136.195 190.365 ;
        RECT 94.505 189.535 94.655 189.555 ;
        RECT 91.275 189.390 91.435 189.500 ;
        RECT 93.565 189.345 93.735 189.535 ;
        RECT 94.020 189.500 94.140 189.505 ;
        RECT 94.020 189.395 94.195 189.500 ;
        RECT 94.035 189.390 94.195 189.395 ;
        RECT 94.485 189.365 94.655 189.535 ;
        RECT 96.785 189.365 96.955 189.555 ;
        RECT 97.705 189.345 97.875 189.535 ;
        RECT 98.165 189.345 98.335 189.535 ;
        RECT 99.080 189.365 99.250 189.555 ;
        RECT 99.545 189.365 99.715 189.555 ;
        RECT 106.900 189.535 107.070 189.555 ;
        RECT 100.015 189.390 100.175 189.500 ;
        RECT 100.935 189.400 101.095 189.510 ;
        RECT 101.385 189.345 101.555 189.535 ;
        RECT 102.760 189.395 102.880 189.505 ;
        RECT 106.440 189.345 106.610 189.535 ;
        RECT 106.900 189.365 107.080 189.535 ;
        RECT 107.370 189.365 107.540 189.555 ;
        RECT 111.505 189.535 111.655 189.555 ;
        RECT 111.505 189.365 111.675 189.535 ;
        RECT 112.885 189.365 113.055 189.555 ;
        RECT 116.565 189.535 116.705 189.555 ;
        RECT 117.945 189.535 118.115 189.555 ;
        RECT 113.340 189.395 113.460 189.505 ;
        RECT 116.565 189.365 116.735 189.535 ;
        RECT 106.910 189.345 107.080 189.365 ;
        RECT 117.025 189.345 117.195 189.535 ;
        RECT 117.480 189.395 117.600 189.505 ;
        RECT 117.945 189.365 118.120 189.535 ;
        RECT 125.305 189.365 125.475 189.535 ;
        RECT 125.775 189.390 125.935 189.500 ;
        RECT 127.140 189.395 127.260 189.505 ;
        RECT 127.605 189.365 127.775 189.555 ;
        RECT 117.950 189.345 118.120 189.365 ;
        RECT 128.055 189.345 128.225 189.535 ;
        RECT 128.535 189.390 128.695 189.500 ;
        RECT 129.445 189.365 129.615 189.555 ;
        RECT 132.665 189.345 132.835 189.535 ;
        RECT 133.125 189.345 133.295 189.555 ;
        RECT 135.885 189.345 136.055 189.555 ;
        RECT 23.505 188.535 24.875 189.345 ;
        RECT 24.885 188.535 27.635 189.345 ;
        RECT 27.645 188.565 29.015 189.345 ;
        RECT 29.025 188.535 34.535 189.345 ;
        RECT 34.545 188.535 37.295 189.345 ;
        RECT 37.765 188.665 41.665 189.345 ;
        RECT 37.765 188.435 38.695 188.665 ;
        RECT 41.905 188.535 44.655 189.345 ;
        RECT 44.810 188.665 46.645 189.345 ;
        RECT 47.110 188.665 48.945 189.345 ;
        RECT 45.715 188.435 46.645 188.665 ;
        RECT 48.015 188.435 48.945 188.665 ;
        RECT 49.275 188.475 49.705 189.260 ;
        RECT 50.645 188.435 53.855 189.345 ;
        RECT 53.865 188.665 57.765 189.345 ;
        RECT 58.005 188.665 61.905 189.345 ;
        RECT 53.865 188.435 54.795 188.665 ;
        RECT 58.005 188.435 58.935 188.665 ;
        RECT 62.605 188.435 63.955 189.345 ;
        RECT 64.915 188.435 67.645 189.345 ;
        RECT 67.665 188.435 71.965 189.345 ;
        RECT 72.265 188.535 75.015 189.345 ;
        RECT 75.035 188.475 75.465 189.260 ;
        RECT 75.485 188.535 78.235 189.345 ;
        RECT 78.245 188.665 82.145 189.345 ;
        RECT 82.385 188.665 86.285 189.345 ;
        RECT 78.245 188.435 79.175 188.665 ;
        RECT 82.385 188.435 83.315 188.665 ;
        RECT 86.525 188.535 88.355 189.345 ;
        RECT 88.375 188.435 91.105 189.345 ;
        RECT 92.045 188.435 93.860 189.345 ;
        RECT 94.805 188.435 98.015 189.345 ;
        RECT 98.040 188.435 99.855 189.345 ;
        RECT 100.795 188.475 101.225 189.260 ;
        RECT 101.255 188.435 102.605 189.345 ;
        RECT 103.085 188.435 106.755 189.345 ;
        RECT 106.765 188.435 108.115 189.345 ;
        RECT 108.230 188.665 117.335 189.345 ;
        RECT 117.805 188.435 123.875 189.345 ;
        RECT 124.245 188.665 125.200 189.345 ;
        RECT 126.555 188.475 126.985 189.260 ;
        RECT 127.005 188.565 128.375 189.345 ;
        RECT 129.445 188.435 132.895 189.345 ;
        RECT 132.985 188.665 134.815 189.345 ;
        RECT 133.470 188.435 134.815 188.665 ;
        RECT 134.825 188.535 136.195 189.345 ;
      LAYER nwell ;
        RECT 23.310 185.315 136.390 188.145 ;
      LAYER pwell ;
        RECT 23.505 184.115 24.875 184.925 ;
        RECT 24.885 184.115 30.395 184.925 ;
        RECT 30.405 184.115 33.155 184.925 ;
        RECT 33.165 184.115 36.375 185.025 ;
        RECT 36.395 184.200 36.825 184.985 ;
        RECT 36.845 184.795 37.775 185.025 ;
        RECT 42.135 184.935 43.725 185.025 ;
        RECT 36.845 184.115 40.745 184.795 ;
        RECT 41.155 184.115 43.725 184.935 ;
        RECT 43.765 184.115 45.115 185.025 ;
        RECT 45.585 184.115 46.935 185.025 ;
        RECT 47.885 184.115 49.700 185.025 ;
        RECT 49.735 184.115 52.465 185.025 ;
        RECT 52.485 184.115 53.855 184.925 ;
        RECT 53.865 184.795 54.795 185.025 ;
        RECT 53.865 184.115 57.765 184.795 ;
        RECT 58.005 184.115 59.835 184.925 ;
        RECT 59.845 184.115 61.195 185.025 ;
        RECT 62.155 184.200 62.585 184.985 ;
        RECT 62.895 184.115 65.815 185.025 ;
        RECT 65.825 184.115 68.575 184.925 ;
        RECT 69.100 184.115 73.175 185.025 ;
        RECT 73.645 184.795 74.570 185.025 ;
        RECT 73.645 184.115 77.315 184.795 ;
        RECT 77.345 184.115 78.695 185.025 ;
        RECT 82.825 184.795 83.755 185.025 ;
        RECT 79.855 184.115 83.755 184.795 ;
        RECT 83.765 184.795 84.695 185.025 ;
        RECT 83.765 184.115 87.665 184.795 ;
        RECT 87.915 184.200 88.345 184.985 ;
        RECT 88.365 184.115 91.115 184.925 ;
        RECT 91.125 184.115 93.875 185.025 ;
        RECT 94.805 184.115 98.015 185.025 ;
        RECT 98.025 184.115 99.395 184.895 ;
        RECT 99.425 184.115 100.775 185.025 ;
        RECT 100.795 184.115 102.145 185.025 ;
        RECT 102.175 184.115 103.525 185.025 ;
        RECT 103.545 184.115 104.915 184.895 ;
        RECT 104.925 184.115 106.295 184.895 ;
        RECT 106.305 184.115 107.675 184.895 ;
        RECT 108.735 184.795 109.665 185.025 ;
        RECT 107.830 184.115 109.665 184.795 ;
        RECT 109.985 184.115 113.655 185.025 ;
        RECT 113.675 184.200 114.105 184.985 ;
        RECT 114.125 184.115 117.780 185.025 ;
        RECT 117.805 184.115 119.175 184.895 ;
        RECT 119.270 184.115 128.375 184.795 ;
        RECT 129.445 184.115 132.895 185.025 ;
        RECT 132.985 184.115 134.355 184.895 ;
        RECT 134.825 184.115 136.195 184.925 ;
        RECT 23.645 183.905 23.815 184.115 ;
        RECT 25.025 183.905 25.195 184.115 ;
        RECT 30.545 183.905 30.715 184.115 ;
        RECT 33.305 183.925 33.475 184.115 ;
        RECT 34.235 183.950 34.395 184.060 ;
        RECT 35.420 183.905 35.590 184.095 ;
        RECT 37.260 183.925 37.430 184.115 ;
        RECT 41.155 184.095 41.295 184.115 ;
        RECT 41.120 183.925 41.295 184.095 ;
        RECT 41.120 183.905 41.290 183.925 ;
        RECT 42.505 183.905 42.675 184.095 ;
        RECT 42.965 183.905 43.135 184.095 ;
        RECT 43.880 183.925 44.050 184.115 ;
        RECT 45.260 183.955 45.380 184.065 ;
        RECT 46.650 183.925 46.820 184.115 ;
        RECT 47.115 183.960 47.275 184.070 ;
        RECT 47.565 183.905 47.735 184.095 ;
        RECT 48.940 183.955 49.060 184.065 ;
        RECT 49.405 183.925 49.575 184.115 ;
        RECT 49.860 183.955 49.980 184.065 ;
        RECT 51.250 183.905 51.420 184.095 ;
        RECT 51.705 183.905 51.875 184.095 ;
        RECT 52.165 183.925 52.335 184.115 ;
        RECT 52.625 183.925 52.795 184.115 ;
        RECT 54.280 183.925 54.450 184.115 ;
        RECT 57.225 183.905 57.395 184.095 ;
        RECT 58.145 183.925 58.315 184.115 ;
        RECT 60.910 184.095 61.080 184.115 ;
        RECT 65.500 184.095 65.670 184.115 ;
        RECT 60.905 183.925 61.080 184.095 ;
        RECT 61.375 183.960 61.535 184.070 ;
        RECT 60.905 183.905 61.075 183.925 ;
        RECT 62.285 183.905 62.455 184.095 ;
        RECT 65.500 183.925 65.675 184.095 ;
        RECT 65.965 183.925 66.135 184.115 ;
        RECT 65.505 183.905 65.675 183.925 ;
        RECT 68.265 183.905 68.435 184.095 ;
        RECT 68.720 183.955 68.840 184.065 ;
        RECT 69.160 183.925 69.330 184.115 ;
        RECT 73.790 184.095 73.960 184.115 ;
        RECT 77.460 184.095 77.630 184.115 ;
        RECT 73.320 183.955 73.440 184.065 ;
        RECT 73.785 183.925 73.960 184.095 ;
        RECT 73.785 183.905 73.955 183.925 ;
        RECT 75.620 183.905 75.790 184.095 ;
        RECT 77.000 183.955 77.120 184.065 ;
        RECT 77.460 183.925 77.640 184.095 ;
        RECT 78.855 183.960 79.015 184.070 ;
        RECT 77.470 183.905 77.640 183.925 ;
        RECT 79.305 183.905 79.475 184.095 ;
        RECT 81.140 183.905 81.310 184.095 ;
        RECT 82.525 183.905 82.695 184.095 ;
        RECT 83.170 183.925 83.340 184.115 ;
        RECT 84.180 183.925 84.350 184.115 ;
        RECT 88.505 184.095 88.675 184.115 ;
        RECT 88.040 183.955 88.160 184.065 ;
        RECT 88.505 183.925 88.680 184.095 ;
        RECT 91.265 183.925 91.435 184.115 ;
        RECT 92.645 183.945 92.815 184.095 ;
        RECT 88.510 183.905 88.680 183.925 ;
        RECT 23.505 183.095 24.875 183.905 ;
        RECT 24.885 183.095 30.395 183.905 ;
        RECT 30.405 183.095 34.075 183.905 ;
        RECT 35.005 183.225 38.905 183.905 ;
        RECT 39.600 183.675 41.290 183.905 ;
        RECT 35.005 182.995 35.935 183.225 ;
        RECT 39.600 182.995 41.435 183.675 ;
        RECT 41.455 182.995 42.805 183.905 ;
        RECT 42.825 183.095 46.495 183.905 ;
        RECT 47.435 182.995 48.785 183.905 ;
        RECT 49.275 183.035 49.705 183.820 ;
        RECT 50.185 182.995 51.535 183.905 ;
        RECT 51.565 183.095 57.075 183.905 ;
        RECT 57.085 183.095 60.755 183.905 ;
        RECT 60.765 183.095 62.135 183.905 ;
        RECT 62.145 183.225 65.355 183.905 ;
        RECT 64.220 182.995 65.355 183.225 ;
        RECT 65.365 182.995 68.085 183.905 ;
        RECT 68.125 183.095 73.635 183.905 ;
        RECT 73.645 183.095 75.015 183.905 ;
        RECT 75.035 183.035 75.465 183.820 ;
        RECT 75.505 182.995 76.855 183.905 ;
        RECT 77.325 182.995 79.155 183.905 ;
        RECT 79.165 183.095 80.995 183.905 ;
        RECT 81.025 182.995 82.375 183.905 ;
        RECT 82.385 183.095 87.895 183.905 ;
        RECT 88.365 182.995 92.035 183.905 ;
        RECT 92.045 182.995 92.935 183.945 ;
        RECT 93.115 183.905 93.285 184.095 ;
        RECT 94.035 183.960 94.195 184.070 ;
        RECT 94.485 183.925 94.655 184.095 ;
        RECT 94.945 183.925 95.115 184.115 ;
        RECT 98.175 183.925 98.345 184.115 ;
        RECT 98.635 183.950 98.795 184.060 ;
        RECT 94.495 183.905 94.655 183.925 ;
        RECT 100.460 183.905 100.630 184.115 ;
        RECT 101.395 183.905 101.565 184.095 ;
        RECT 101.845 183.925 102.015 184.115 ;
        RECT 103.225 183.925 103.395 184.115 ;
        RECT 103.685 184.095 103.855 184.115 ;
        RECT 103.685 183.925 103.860 184.095 ;
        RECT 103.690 183.905 103.860 183.925 ;
        RECT 105.070 183.905 105.240 184.095 ;
        RECT 105.525 183.905 105.695 184.095 ;
        RECT 105.975 183.925 106.145 184.115 ;
        RECT 107.355 183.925 107.525 184.115 ;
        RECT 107.830 184.095 107.995 184.115 ;
        RECT 107.825 183.925 107.995 184.095 ;
        RECT 110.130 183.925 110.300 184.115 ;
        RECT 111.500 183.905 111.670 184.095 ;
        RECT 114.270 183.925 114.440 184.115 ;
        RECT 114.725 183.905 114.895 184.095 ;
        RECT 92.965 183.125 94.335 183.905 ;
        RECT 94.495 182.995 98.150 183.905 ;
        RECT 99.425 182.995 100.775 183.905 ;
        RECT 100.795 183.035 101.225 183.820 ;
        RECT 101.245 183.125 102.615 183.905 ;
        RECT 102.625 182.995 103.975 183.905 ;
        RECT 104.005 182.995 105.355 183.905 ;
        RECT 105.385 182.995 108.595 183.905 ;
        RECT 108.605 182.995 111.815 183.905 ;
        RECT 111.825 182.995 115.035 183.905 ;
        RECT 115.185 183.675 115.355 184.095 ;
        RECT 118.865 183.925 119.035 184.115 ;
        RECT 120.710 183.905 120.880 184.095 ;
        RECT 125.755 183.905 125.925 184.095 ;
        RECT 126.220 183.955 126.340 184.065 ;
        RECT 127.150 183.905 127.320 184.095 ;
        RECT 128.065 183.925 128.235 184.115 ;
        RECT 128.535 183.960 128.695 184.070 ;
        RECT 129.445 183.905 129.615 184.095 ;
        RECT 132.665 183.925 132.835 184.115 ;
        RECT 133.135 183.925 133.305 184.115 ;
        RECT 134.045 183.905 134.215 184.095 ;
        RECT 134.500 183.955 134.620 184.065 ;
        RECT 135.885 183.905 136.055 184.115 ;
        RECT 116.465 183.675 120.555 183.905 ;
        RECT 115.080 182.995 120.555 183.675 ;
        RECT 120.565 182.995 124.665 183.905 ;
        RECT 124.705 183.125 126.075 183.905 ;
        RECT 126.555 183.035 126.985 183.820 ;
        RECT 127.005 182.995 129.215 183.905 ;
        RECT 129.385 182.995 132.835 183.905 ;
        RECT 132.985 183.125 134.355 183.905 ;
        RECT 134.825 183.095 136.195 183.905 ;
      LAYER nwell ;
        RECT 23.310 179.875 136.390 182.705 ;
      LAYER pwell ;
        RECT 23.505 178.675 24.875 179.485 ;
        RECT 25.545 179.355 29.475 179.585 ;
        RECT 25.060 178.675 29.475 179.355 ;
        RECT 29.485 178.675 33.155 179.485 ;
        RECT 33.165 178.675 34.535 179.485 ;
        RECT 34.545 178.675 36.375 179.585 ;
        RECT 36.395 178.760 36.825 179.545 ;
        RECT 37.330 179.355 38.675 179.585 ;
        RECT 36.845 178.675 38.675 179.355 ;
        RECT 38.685 178.675 40.515 179.585 ;
        RECT 40.535 178.675 41.885 179.585 ;
        RECT 41.905 178.675 44.655 179.485 ;
        RECT 44.675 178.675 48.335 179.585 ;
        RECT 48.515 178.675 52.015 179.585 ;
        RECT 52.025 178.675 53.375 179.585 ;
        RECT 54.065 179.495 55.015 179.585 ;
        RECT 54.065 178.675 55.995 179.495 ;
        RECT 56.165 178.675 57.995 179.585 ;
        RECT 58.020 179.355 59.390 179.585 ;
        RECT 58.020 178.675 60.295 179.355 ;
        RECT 60.305 178.675 62.120 179.585 ;
        RECT 62.155 178.760 62.585 179.545 ;
        RECT 62.605 178.675 66.275 179.585 ;
        RECT 66.300 178.675 69.955 179.585 ;
        RECT 69.965 178.675 75.475 179.485 ;
        RECT 75.485 178.675 77.315 179.485 ;
        RECT 77.325 178.675 79.155 179.585 ;
        RECT 79.245 178.675 82.245 179.585 ;
        RECT 82.465 178.675 85.465 179.585 ;
        RECT 85.605 178.675 86.955 179.585 ;
        RECT 87.915 178.760 88.345 179.545 ;
        RECT 88.365 178.675 92.035 179.585 ;
        RECT 23.645 178.465 23.815 178.675 ;
        RECT 25.060 178.655 25.170 178.675 ;
        RECT 25.000 178.485 25.170 178.655 ;
        RECT 26.405 178.465 26.575 178.655 ;
        RECT 26.865 178.465 27.035 178.655 ;
        RECT 29.625 178.485 29.795 178.675 ;
        RECT 32.385 178.465 32.555 178.655 ;
        RECT 33.305 178.485 33.475 178.675 ;
        RECT 34.690 178.485 34.860 178.675 ;
        RECT 23.505 177.655 24.875 178.465 ;
        RECT 24.885 177.785 26.715 178.465 ;
        RECT 24.885 177.555 26.230 177.785 ;
        RECT 26.725 177.655 32.235 178.465 ;
        RECT 32.245 177.655 35.915 178.465 ;
        RECT 36.070 178.435 36.240 178.655 ;
        RECT 36.985 178.485 37.155 178.675 ;
        RECT 38.830 178.485 39.000 178.675 ;
        RECT 40.200 178.465 40.370 178.655 ;
        RECT 40.665 178.465 40.835 178.675 ;
        RECT 42.045 178.485 42.215 178.675 ;
        RECT 44.790 178.655 44.960 178.675 ;
        RECT 48.515 178.655 48.650 178.675 ;
        RECT 53.090 178.655 53.260 178.675 ;
        RECT 44.790 178.485 44.975 178.655 ;
        RECT 44.805 178.465 44.975 178.485 ;
        RECT 47.105 178.465 47.275 178.655 ;
        RECT 48.480 178.485 48.650 178.655 ;
        RECT 48.945 178.465 49.115 178.655 ;
        RECT 49.865 178.465 50.035 178.655 ;
        RECT 51.710 178.465 51.880 178.655 ;
        RECT 53.085 178.485 53.260 178.655 ;
        RECT 55.845 178.655 55.995 178.675 ;
        RECT 53.540 178.515 53.660 178.625 ;
        RECT 55.845 178.485 56.015 178.655 ;
        RECT 56.310 178.485 56.480 178.675 ;
        RECT 53.085 178.465 53.255 178.485 ;
        RECT 58.605 178.465 58.775 178.655 ;
        RECT 59.980 178.485 60.150 178.675 ;
        RECT 60.440 178.515 60.560 178.625 ;
        RECT 60.905 178.465 61.075 178.655 ;
        RECT 61.825 178.485 61.995 178.675 ;
        RECT 62.750 178.485 62.920 178.675 ;
        RECT 63.670 178.465 63.840 178.655 ;
        RECT 67.345 178.465 67.515 178.655 ;
        RECT 69.640 178.485 69.810 178.675 ;
        RECT 70.105 178.485 70.275 178.675 ;
        RECT 72.865 178.465 73.035 178.655 ;
        RECT 74.700 178.515 74.820 178.625 ;
        RECT 75.625 178.465 75.795 178.675 ;
        RECT 77.470 178.485 77.640 178.675 ;
        RECT 79.305 178.485 79.475 178.675 ;
        RECT 82.525 178.485 82.695 178.675 ;
        RECT 82.980 178.465 83.150 178.655 ;
        RECT 86.670 178.485 86.840 178.675 ;
        RECT 87.135 178.520 87.295 178.630 ;
        RECT 88.510 178.485 88.680 178.675 ;
        RECT 92.045 178.635 92.935 179.585 ;
        RECT 92.965 178.675 94.335 179.455 ;
        RECT 94.345 179.385 95.730 179.585 ;
        RECT 98.225 179.495 99.175 179.585 ;
        RECT 94.345 178.705 98.015 179.385 ;
        RECT 94.345 178.675 95.715 178.705 ;
        RECT 92.185 178.465 92.355 178.635 ;
        RECT 92.645 178.485 92.815 178.635 ;
        RECT 93.105 178.485 93.275 178.675 ;
        RECT 95.405 178.465 95.575 178.655 ;
        RECT 97.705 178.485 97.875 178.705 ;
        RECT 98.225 178.675 100.155 179.495 ;
        RECT 101.245 178.905 103.995 179.585 ;
        RECT 100.005 178.655 100.155 178.675 ;
        RECT 101.385 178.675 103.995 178.905 ;
        RECT 104.015 178.675 106.755 179.355 ;
        RECT 106.765 178.675 109.975 179.585 ;
        RECT 112.065 179.355 113.655 179.585 ;
        RECT 109.985 178.675 113.655 179.355 ;
        RECT 113.675 178.760 114.105 179.545 ;
        RECT 114.210 178.675 123.315 179.355 ;
        RECT 123.325 178.675 132.430 179.355 ;
        RECT 132.985 178.675 134.355 179.455 ;
        RECT 134.825 178.675 136.195 179.485 ;
        RECT 97.705 178.465 97.870 178.485 ;
        RECT 99.075 178.465 99.245 178.655 ;
        RECT 100.005 178.485 100.175 178.655 ;
        RECT 100.465 178.465 100.635 178.655 ;
        RECT 101.385 178.485 101.555 178.675 ;
        RECT 102.765 178.465 102.935 178.655 ;
        RECT 105.985 178.465 106.155 178.655 ;
        RECT 106.445 178.465 106.615 178.675 ;
        RECT 106.905 178.485 107.075 178.675 ;
        RECT 110.130 178.485 110.300 178.675 ;
        RECT 116.560 178.465 116.730 178.655 ;
        RECT 117.025 178.465 117.195 178.655 ;
        RECT 120.700 178.515 120.820 178.625 ;
        RECT 121.160 178.465 121.330 178.655 ;
        RECT 122.545 178.465 122.715 178.655 ;
        RECT 123.005 178.485 123.175 178.675 ;
        RECT 123.465 178.485 123.635 178.675 ;
        RECT 123.925 178.465 124.095 178.655 ;
        RECT 127.150 178.465 127.320 178.655 ;
        RECT 132.660 178.515 132.780 178.625 ;
        RECT 134.045 178.485 134.215 178.675 ;
        RECT 134.500 178.465 134.670 178.655 ;
        RECT 135.885 178.465 136.055 178.675 ;
        RECT 38.200 178.435 39.135 178.465 ;
        RECT 36.070 178.235 39.135 178.435 ;
        RECT 35.925 177.755 39.135 178.235 ;
        RECT 35.925 177.555 36.855 177.755 ;
        RECT 38.185 177.555 39.135 177.755 ;
        RECT 39.165 177.555 40.515 178.465 ;
        RECT 40.525 177.655 43.275 178.465 ;
        RECT 43.285 177.555 45.100 178.465 ;
        RECT 45.135 177.555 49.255 178.465 ;
        RECT 49.275 177.595 49.705 178.380 ;
        RECT 49.740 177.555 51.555 178.465 ;
        RECT 51.565 177.555 52.915 178.465 ;
        RECT 52.945 177.655 58.455 178.465 ;
        RECT 58.465 177.655 60.295 178.465 ;
        RECT 60.765 177.785 63.515 178.465 ;
        RECT 62.585 177.555 63.515 177.785 ;
        RECT 63.525 177.785 67.110 178.465 ;
        RECT 63.525 177.555 64.445 177.785 ;
        RECT 67.205 177.655 72.715 178.465 ;
        RECT 72.725 177.655 74.555 178.465 ;
        RECT 75.035 177.595 75.465 178.380 ;
        RECT 75.485 177.655 79.155 178.465 ;
        RECT 80.085 177.555 83.295 178.465 ;
        RECT 83.390 177.785 92.495 178.465 ;
        RECT 92.505 177.555 95.715 178.465 ;
        RECT 96.035 177.785 97.870 178.465 ;
        RECT 96.035 177.555 96.965 177.785 ;
        RECT 98.025 177.685 99.395 178.465 ;
        RECT 99.415 177.555 100.765 178.465 ;
        RECT 100.795 177.595 101.225 178.380 ;
        RECT 101.245 177.785 103.075 178.465 ;
        RECT 103.085 177.555 106.295 178.465 ;
        RECT 106.305 177.785 115.410 178.465 ;
        RECT 115.525 177.555 116.875 178.465 ;
        RECT 116.885 177.655 120.555 178.465 ;
        RECT 121.045 177.555 122.395 178.465 ;
        RECT 122.405 177.685 123.775 178.465 ;
        RECT 123.785 177.785 126.525 178.465 ;
        RECT 126.555 177.595 126.985 178.380 ;
        RECT 127.005 177.555 131.135 178.465 ;
        RECT 131.270 177.555 134.815 178.465 ;
        RECT 134.825 177.655 136.195 178.465 ;
      LAYER nwell ;
        RECT 23.310 174.435 136.390 177.265 ;
      LAYER pwell ;
        RECT 23.505 173.235 24.875 174.045 ;
        RECT 24.885 173.235 26.255 174.045 ;
        RECT 26.275 173.235 27.625 174.145 ;
        RECT 29.490 173.915 30.855 174.145 ;
        RECT 32.685 173.915 33.615 174.145 ;
        RECT 34.775 174.055 36.365 174.145 ;
        RECT 27.645 173.235 30.855 173.915 ;
        RECT 30.865 173.235 33.615 173.915 ;
        RECT 33.795 173.235 36.365 174.055 ;
        RECT 36.395 173.320 36.825 174.105 ;
        RECT 39.585 173.915 40.515 174.145 ;
        RECT 36.845 173.235 40.515 173.915 ;
        RECT 40.525 173.235 44.195 174.045 ;
        RECT 44.345 173.235 47.795 174.145 ;
        RECT 48.805 173.235 50.620 174.145 ;
        RECT 50.645 173.235 56.155 174.045 ;
        RECT 56.635 173.235 57.985 174.145 ;
        RECT 58.005 173.235 61.675 174.045 ;
        RECT 62.155 173.320 62.585 174.105 ;
        RECT 64.425 173.915 65.355 174.145 ;
        RECT 62.605 173.235 65.355 173.915 ;
        RECT 66.285 173.945 67.215 174.145 ;
        RECT 68.550 173.945 69.495 174.145 ;
        RECT 66.285 173.465 69.495 173.945 ;
        RECT 66.425 173.265 69.495 173.465 ;
        RECT 23.645 173.025 23.815 173.235 ;
        RECT 25.025 173.025 25.195 173.235 ;
        RECT 26.405 173.045 26.575 173.235 ;
        RECT 26.875 173.070 27.035 173.180 ;
        RECT 27.790 173.045 27.960 173.235 ;
        RECT 28.705 173.025 28.875 173.215 ;
        RECT 29.165 173.025 29.335 173.215 ;
        RECT 31.005 173.045 31.175 173.235 ;
        RECT 33.795 173.215 33.935 173.235 ;
        RECT 33.765 173.045 33.935 173.215 ;
        RECT 34.680 173.075 34.800 173.185 ;
        RECT 35.150 173.025 35.320 173.215 ;
        RECT 36.985 173.045 37.155 173.235 ;
        RECT 40.665 173.045 40.835 173.235 ;
        RECT 23.505 172.215 24.875 173.025 ;
        RECT 24.885 172.345 26.715 173.025 ;
        RECT 27.645 172.245 29.015 173.025 ;
        RECT 29.025 172.215 34.535 173.025 ;
        RECT 35.005 172.345 39.595 173.025 ;
        RECT 39.605 172.995 40.540 173.025 ;
        RECT 42.500 172.995 42.670 173.215 ;
        RECT 42.965 173.045 43.135 173.215 ;
        RECT 39.605 172.795 42.670 172.995 ;
        RECT 42.985 173.025 43.135 173.045 ;
        RECT 45.265 173.025 45.435 173.215 ;
        RECT 47.565 173.045 47.735 173.235 ;
        RECT 48.035 173.080 48.195 173.190 ;
        RECT 48.940 173.075 49.060 173.185 ;
        RECT 49.865 173.025 50.035 173.215 ;
        RECT 50.325 173.045 50.495 173.235 ;
        RECT 50.785 173.045 50.955 173.235 ;
        RECT 55.385 173.025 55.555 173.215 ;
        RECT 56.300 173.075 56.420 173.185 ;
        RECT 56.765 173.045 56.935 173.235 ;
        RECT 58.145 173.045 58.315 173.235 ;
        RECT 60.905 173.025 61.075 173.215 ;
        RECT 61.820 173.075 61.940 173.185 ;
        RECT 62.745 173.045 62.915 173.235 ;
        RECT 65.515 173.080 65.675 173.190 ;
        RECT 66.425 173.045 66.595 173.265 ;
        RECT 68.550 173.235 69.495 173.265 ;
        RECT 69.515 173.235 72.245 174.145 ;
        RECT 72.265 173.235 73.615 174.145 ;
        RECT 73.645 173.235 75.475 174.045 ;
        RECT 75.485 173.235 78.695 174.145 ;
        RECT 78.705 173.235 82.780 174.145 ;
        RECT 82.860 173.235 84.675 174.145 ;
        RECT 66.880 173.025 67.050 173.215 ;
        RECT 67.340 173.075 67.460 173.185 ;
        RECT 35.490 172.115 36.830 172.345 ;
        RECT 39.605 172.315 42.815 172.795 ;
        RECT 39.605 172.115 40.555 172.315 ;
        RECT 41.885 172.115 42.815 172.315 ;
        RECT 42.985 172.205 44.915 173.025 ;
        RECT 45.125 172.215 48.795 173.025 ;
        RECT 43.965 172.115 44.915 172.205 ;
        RECT 49.275 172.155 49.705 172.940 ;
        RECT 49.725 172.215 55.235 173.025 ;
        RECT 55.245 172.215 60.755 173.025 ;
        RECT 60.765 172.215 63.515 173.025 ;
        RECT 63.525 172.345 67.195 173.025 ;
        RECT 67.805 172.995 67.975 173.215 ;
        RECT 71.030 173.025 71.200 173.215 ;
        RECT 71.945 173.045 72.115 173.235 ;
        RECT 73.330 173.045 73.500 173.235 ;
        RECT 73.785 173.045 73.955 173.235 ;
        RECT 78.385 173.215 78.555 173.235 ;
        RECT 74.255 173.070 74.415 173.180 ;
        RECT 75.635 173.070 75.795 173.180 ;
        RECT 77.925 173.025 78.095 173.215 ;
        RECT 78.385 173.045 78.560 173.215 ;
        RECT 82.075 173.070 82.235 173.180 ;
        RECT 82.550 173.045 82.720 173.235 ;
        RECT 82.985 173.045 83.155 173.235 ;
        RECT 85.605 173.195 86.495 174.145 ;
        RECT 86.525 173.235 87.895 174.015 ;
        RECT 87.915 173.320 88.345 174.105 ;
        RECT 89.305 173.235 90.655 174.145 ;
        RECT 90.665 173.235 93.875 174.145 ;
        RECT 93.970 173.235 103.075 173.915 ;
        RECT 103.105 173.235 104.455 174.145 ;
        RECT 104.465 173.235 108.135 174.045 ;
        RECT 108.145 173.235 112.275 174.145 ;
        RECT 112.305 173.235 113.655 174.145 ;
        RECT 113.675 173.320 114.105 174.105 ;
        RECT 133.470 173.915 134.815 174.145 ;
        RECT 114.125 173.235 123.230 173.915 ;
        RECT 123.325 173.235 132.430 173.915 ;
        RECT 132.985 173.235 134.815 173.915 ;
        RECT 134.825 173.235 136.195 174.045 ;
        RECT 84.835 173.080 84.995 173.190 ;
        RECT 86.205 173.045 86.375 173.195 ;
        RECT 86.665 173.045 86.835 173.235 ;
        RECT 88.515 173.080 88.675 173.190 ;
        RECT 90.340 173.045 90.510 173.235 ;
        RECT 78.390 173.025 78.560 173.045 ;
        RECT 82.985 173.025 83.185 173.045 ;
        RECT 86.665 173.025 86.865 173.045 ;
        RECT 91.730 173.025 91.900 173.215 ;
        RECT 93.565 173.045 93.735 173.235 ;
        RECT 94.480 173.025 94.650 173.215 ;
        RECT 94.940 173.075 95.060 173.185 ;
        RECT 95.405 173.045 95.575 173.215 ;
        RECT 95.415 173.025 95.575 173.045 ;
        RECT 100.460 173.025 100.630 173.215 ;
        RECT 102.305 173.025 102.475 173.215 ;
        RECT 102.765 173.045 102.935 173.235 ;
        RECT 104.140 173.045 104.310 173.235 ;
        RECT 104.605 173.045 104.775 173.235 ;
        RECT 105.520 173.025 105.690 173.215 ;
        RECT 111.960 173.045 112.130 173.235 ;
        RECT 112.420 173.045 112.590 173.235 ;
        RECT 114.265 173.045 114.435 173.235 ;
        RECT 114.725 173.025 114.895 173.215 ;
        RECT 115.185 173.025 115.355 173.215 ;
        RECT 117.940 173.075 118.060 173.185 ;
        RECT 121.160 173.025 121.330 173.215 ;
        RECT 123.465 173.045 123.635 173.235 ;
        RECT 125.300 173.025 125.470 173.215 ;
        RECT 125.775 173.070 125.935 173.180 ;
        RECT 130.845 173.025 131.015 173.215 ;
        RECT 132.660 173.075 132.780 173.185 ;
        RECT 133.125 173.045 133.295 173.235 ;
        RECT 134.500 173.025 134.670 173.215 ;
        RECT 135.885 173.025 136.055 173.235 ;
        RECT 69.930 172.995 70.875 173.025 ;
        RECT 67.805 172.795 70.875 172.995 ;
        RECT 66.270 172.115 67.195 172.345 ;
        RECT 67.665 172.315 70.875 172.795 ;
        RECT 67.665 172.115 68.595 172.315 ;
        RECT 69.930 172.115 70.875 172.315 ;
        RECT 70.885 172.115 73.805 173.025 ;
        RECT 75.035 172.155 75.465 172.940 ;
        RECT 76.405 172.115 78.220 173.025 ;
        RECT 78.245 172.115 81.900 173.025 ;
        RECT 82.985 172.345 86.515 173.025 ;
        RECT 86.665 172.345 90.195 173.025 ;
        RECT 83.690 172.115 86.515 172.345 ;
        RECT 87.370 172.115 90.195 172.345 ;
        RECT 90.665 172.115 92.015 173.025 ;
        RECT 92.045 172.115 94.795 173.025 ;
        RECT 95.415 172.115 99.070 173.025 ;
        RECT 99.425 172.115 100.775 173.025 ;
        RECT 100.795 172.155 101.225 172.940 ;
        RECT 101.255 172.115 102.605 173.025 ;
        RECT 102.625 172.115 105.835 173.025 ;
        RECT 105.930 172.345 115.035 173.025 ;
        RECT 115.045 172.215 117.795 173.025 ;
        RECT 118.360 172.115 121.475 173.025 ;
        RECT 121.745 172.115 125.615 173.025 ;
        RECT 126.555 172.155 126.985 172.940 ;
        RECT 127.100 172.345 131.125 173.025 ;
        RECT 129.780 172.115 131.125 172.345 ;
        RECT 131.145 172.115 134.815 173.025 ;
        RECT 134.825 172.215 136.195 173.025 ;
      LAYER nwell ;
        RECT 23.310 168.995 136.390 171.825 ;
      LAYER pwell ;
        RECT 23.505 167.795 24.875 168.605 ;
        RECT 24.885 168.475 26.230 168.705 ;
        RECT 24.885 167.795 26.715 168.475 ;
        RECT 27.645 167.795 29.015 168.575 ;
        RECT 29.025 167.795 34.535 168.605 ;
        RECT 34.545 167.795 36.375 168.605 ;
        RECT 36.395 167.880 36.825 168.665 ;
        RECT 39.825 168.615 40.775 168.705 ;
        RECT 36.845 167.795 38.675 168.605 ;
        RECT 38.845 167.795 40.775 168.615 ;
        RECT 40.985 167.795 43.735 168.705 ;
        RECT 44.230 168.475 45.575 168.705 ;
        RECT 46.635 168.475 47.565 168.705 ;
        RECT 43.745 167.795 45.575 168.475 ;
        RECT 45.730 167.795 47.565 168.475 ;
        RECT 47.885 167.795 53.395 168.605 ;
        RECT 53.405 167.795 55.235 168.605 ;
        RECT 55.705 168.025 58.905 168.705 ;
        RECT 55.850 167.795 58.905 168.025 ;
        RECT 59.405 167.795 60.755 168.705 ;
        RECT 60.765 167.795 62.135 168.605 ;
        RECT 62.155 167.880 62.585 168.665 ;
        RECT 62.605 167.795 65.355 168.605 ;
        RECT 65.825 167.795 69.300 168.705 ;
        RECT 69.505 167.795 72.285 168.705 ;
        RECT 73.775 168.475 74.705 168.705 ;
        RECT 72.870 167.795 74.705 168.475 ;
        RECT 75.025 167.795 78.695 168.605 ;
        RECT 79.640 167.795 81.455 168.705 ;
        RECT 81.925 167.795 83.740 168.705 ;
        RECT 23.645 167.585 23.815 167.795 ;
        RECT 25.025 167.585 25.195 167.775 ;
        RECT 26.405 167.605 26.575 167.795 ;
        RECT 26.865 167.585 27.035 167.775 ;
        RECT 28.705 167.605 28.875 167.795 ;
        RECT 29.165 167.605 29.335 167.795 ;
        RECT 32.385 167.585 32.555 167.775 ;
        RECT 34.685 167.605 34.855 167.795 ;
        RECT 36.065 167.585 36.235 167.775 ;
        RECT 36.985 167.605 37.155 167.795 ;
        RECT 38.845 167.775 38.995 167.795 ;
        RECT 38.825 167.605 38.995 167.775 ;
        RECT 39.745 167.585 39.915 167.775 ;
        RECT 41.125 167.605 41.295 167.795 ;
        RECT 42.975 167.585 43.145 167.775 ;
        RECT 43.435 167.630 43.595 167.740 ;
        RECT 43.885 167.605 44.055 167.795 ;
        RECT 45.730 167.775 45.895 167.795 ;
        RECT 44.345 167.605 44.515 167.775 ;
        RECT 45.725 167.605 45.895 167.775 ;
        RECT 48.025 167.605 48.195 167.795 ;
        RECT 48.495 167.630 48.655 167.740 ;
        RECT 44.355 167.585 44.515 167.605 ;
        RECT 49.870 167.585 50.040 167.775 ;
        RECT 53.545 167.605 53.715 167.795 ;
        RECT 55.380 167.635 55.500 167.745 ;
        RECT 55.850 167.605 56.020 167.795 ;
        RECT 56.305 167.585 56.475 167.775 ;
        RECT 59.060 167.635 59.180 167.745 ;
        RECT 59.520 167.585 59.690 167.795 ;
        RECT 59.990 167.585 60.160 167.775 ;
        RECT 60.905 167.605 61.075 167.795 ;
        RECT 61.365 167.585 61.535 167.775 ;
        RECT 62.745 167.605 62.915 167.795 ;
        RECT 65.500 167.635 65.620 167.745 ;
        RECT 65.970 167.605 66.140 167.795 ;
        RECT 66.885 167.585 67.055 167.775 ;
        RECT 69.645 167.605 69.815 167.795 ;
        RECT 72.870 167.775 73.035 167.795 ;
        RECT 72.415 167.630 72.575 167.740 ;
        RECT 72.865 167.605 73.035 167.775 ;
        RECT 73.325 167.585 73.495 167.775 ;
        RECT 75.165 167.605 75.335 167.795 ;
        RECT 75.630 167.585 75.800 167.775 ;
        RECT 78.855 167.640 79.015 167.750 ;
        RECT 79.765 167.605 79.935 167.795 ;
        RECT 80.235 167.630 80.395 167.740 ;
        RECT 81.145 167.585 81.315 167.775 ;
        RECT 81.600 167.635 81.720 167.745 ;
        RECT 82.995 167.585 83.165 167.775 ;
        RECT 83.445 167.605 83.615 167.795 ;
        RECT 83.765 167.755 84.655 168.705 ;
        RECT 86.950 168.505 87.895 168.705 ;
        RECT 85.145 167.825 87.895 168.505 ;
        RECT 87.915 167.880 88.345 168.665 ;
        RECT 84.365 167.745 84.535 167.755 ;
        RECT 84.835 167.745 85.005 167.775 ;
        RECT 84.360 167.635 84.535 167.745 ;
        RECT 84.820 167.635 85.005 167.745 ;
        RECT 84.365 167.605 84.535 167.635 ;
        RECT 84.835 167.585 85.005 167.635 ;
        RECT 85.290 167.605 85.460 167.825 ;
        RECT 86.950 167.795 87.895 167.825 ;
        RECT 88.365 167.795 91.115 168.705 ;
        RECT 91.125 167.795 94.335 168.705 ;
        RECT 94.345 168.475 95.265 168.705 ;
        RECT 94.345 167.795 97.930 168.475 ;
        RECT 98.485 167.795 100.300 168.705 ;
        RECT 100.325 167.795 103.800 168.705 ;
        RECT 104.925 167.795 111.835 168.705 ;
        RECT 112.295 167.795 113.645 168.705 ;
        RECT 113.675 167.880 114.105 168.665 ;
        RECT 114.125 167.795 123.230 168.475 ;
        RECT 124.255 167.795 125.605 168.705 ;
        RECT 125.625 167.795 134.730 168.475 ;
        RECT 134.825 167.795 136.195 168.605 ;
        RECT 90.800 167.775 90.970 167.795 ;
        RECT 86.215 167.585 86.385 167.775 ;
        RECT 87.585 167.585 87.755 167.775 ;
        RECT 90.345 167.585 90.515 167.775 ;
        RECT 90.800 167.625 90.975 167.775 ;
        RECT 23.505 166.775 24.875 167.585 ;
        RECT 24.885 166.905 26.715 167.585 ;
        RECT 26.725 166.775 32.235 167.585 ;
        RECT 32.245 166.775 35.915 167.585 ;
        RECT 35.925 166.775 37.295 167.585 ;
        RECT 37.315 166.675 40.045 167.585 ;
        RECT 40.065 166.675 43.275 167.585 ;
        RECT 44.355 166.675 48.010 167.585 ;
        RECT 49.275 166.715 49.705 167.500 ;
        RECT 49.725 166.675 53.395 167.585 ;
        RECT 53.405 166.675 56.615 167.585 ;
        RECT 56.625 166.905 59.835 167.585 ;
        RECT 56.625 166.675 57.990 166.905 ;
        RECT 59.845 166.675 61.195 167.585 ;
        RECT 61.225 166.775 66.735 167.585 ;
        RECT 66.745 166.775 72.255 167.585 ;
        RECT 73.185 166.905 75.015 167.585 ;
        RECT 75.035 166.715 75.465 167.500 ;
        RECT 75.485 166.675 79.875 167.585 ;
        RECT 81.005 166.905 82.835 167.585 ;
        RECT 82.845 166.805 84.215 167.585 ;
        RECT 84.685 166.805 86.055 167.585 ;
        RECT 86.065 166.805 87.435 167.585 ;
        RECT 87.445 166.805 88.815 167.585 ;
        RECT 88.825 166.905 90.655 167.585 ;
        RECT 88.825 166.675 90.170 166.905 ;
        RECT 90.685 166.675 91.575 167.625 ;
        RECT 94.025 167.605 94.195 167.795 ;
        RECT 94.490 167.775 94.660 167.795 ;
        RECT 94.485 167.605 94.660 167.775 ;
        RECT 94.485 167.585 94.655 167.605 ;
        RECT 95.865 167.585 96.035 167.775 ;
        RECT 98.160 167.635 98.280 167.745 ;
        RECT 99.085 167.585 99.255 167.775 ;
        RECT 100.005 167.605 100.175 167.795 ;
        RECT 100.470 167.775 100.640 167.795 ;
        RECT 100.465 167.605 100.640 167.775 ;
        RECT 100.465 167.585 100.635 167.605 ;
        RECT 91.585 166.675 94.795 167.585 ;
        RECT 94.815 166.675 96.165 167.585 ;
        RECT 96.185 166.675 99.395 167.585 ;
        RECT 99.405 166.805 100.775 167.585 ;
        RECT 101.245 167.555 102.640 167.585 ;
        RECT 103.685 167.555 103.855 167.775 ;
        RECT 104.120 167.750 104.290 167.775 ;
        RECT 104.120 167.640 104.315 167.750 ;
        RECT 104.120 167.585 104.290 167.640 ;
        RECT 105.065 167.605 105.235 167.795 ;
        RECT 109.210 167.585 109.380 167.775 ;
        RECT 109.665 167.585 109.835 167.775 ;
        RECT 112.425 167.605 112.595 167.795 ;
        RECT 114.265 167.605 114.435 167.795 ;
        RECT 118.865 167.585 119.035 167.775 ;
        RECT 123.475 167.640 123.635 167.750 ;
        RECT 125.305 167.605 125.475 167.795 ;
        RECT 125.765 167.605 125.935 167.795 ;
        RECT 100.795 166.715 101.225 167.500 ;
        RECT 101.245 166.875 103.980 167.555 ;
        RECT 101.245 166.675 102.655 166.875 ;
        RECT 104.060 166.675 108.135 167.585 ;
        RECT 108.145 166.675 109.495 167.585 ;
        RECT 109.525 166.905 118.630 167.585 ;
        RECT 118.725 166.905 123.540 167.585 ;
        RECT 123.785 167.555 124.730 167.585 ;
        RECT 126.220 167.555 126.390 167.775 ;
        RECT 127.145 167.585 127.315 167.775 ;
        RECT 134.505 167.585 134.675 167.775 ;
        RECT 135.885 167.585 136.055 167.795 ;
        RECT 123.785 166.875 126.535 167.555 ;
        RECT 123.785 166.675 124.730 166.875 ;
        RECT 126.555 166.715 126.985 167.500 ;
        RECT 127.145 167.355 132.050 167.585 ;
        RECT 127.005 166.675 132.050 167.355 ;
        RECT 132.065 167.355 134.675 167.585 ;
        RECT 132.065 166.675 134.815 167.355 ;
        RECT 134.825 166.775 136.195 167.585 ;
      LAYER nwell ;
        RECT 23.310 163.555 136.390 166.385 ;
      LAYER pwell ;
        RECT 23.505 162.355 24.875 163.165 ;
        RECT 24.885 162.355 30.395 163.165 ;
        RECT 30.405 162.355 35.915 163.165 ;
        RECT 36.395 162.440 36.825 163.225 ;
        RECT 36.845 162.355 38.215 163.165 ;
        RECT 40.070 163.035 41.435 163.265 ;
        RECT 43.265 163.035 44.195 163.265 ;
        RECT 38.225 162.355 41.435 163.035 ;
        RECT 41.445 162.355 44.195 163.035 ;
        RECT 44.205 162.355 46.955 163.165 ;
        RECT 47.425 162.355 50.635 163.265 ;
        RECT 50.645 162.355 53.395 163.165 ;
        RECT 53.885 162.355 55.235 163.265 ;
        RECT 55.245 162.585 57.080 163.265 ;
        RECT 55.390 162.355 57.080 162.585 ;
        RECT 58.005 162.355 61.675 163.265 ;
        RECT 62.155 162.440 62.585 163.225 ;
        RECT 62.605 163.035 63.950 163.265 ;
        RECT 62.605 162.355 64.435 163.035 ;
        RECT 64.445 162.355 69.955 163.165 ;
        RECT 69.965 162.355 71.335 163.165 ;
        RECT 71.355 162.355 74.085 163.265 ;
        RECT 74.120 162.355 75.935 163.265 ;
        RECT 76.865 162.355 78.235 163.135 ;
        RECT 78.255 162.355 79.605 163.265 ;
        RECT 79.625 162.355 83.280 163.265 ;
        RECT 83.765 162.355 85.580 163.265 ;
        RECT 23.645 162.145 23.815 162.355 ;
        RECT 25.025 162.145 25.195 162.355 ;
        RECT 30.545 162.145 30.715 162.355 ;
        RECT 36.065 162.305 36.235 162.335 ;
        RECT 36.060 162.195 36.235 162.305 ;
        RECT 36.065 162.145 36.235 162.195 ;
        RECT 36.985 162.165 37.155 162.355 ;
        RECT 37.900 162.195 38.020 162.305 ;
        RECT 38.370 162.165 38.540 162.355 ;
        RECT 39.745 162.145 39.915 162.335 ;
        RECT 40.205 162.145 40.375 162.335 ;
        RECT 41.585 162.165 41.755 162.355 ;
        RECT 44.345 162.165 44.515 162.355 ;
        RECT 44.805 162.165 44.975 162.335 ;
        RECT 44.805 162.145 44.955 162.165 ;
        RECT 46.645 162.145 46.815 162.335 ;
        RECT 47.105 162.305 47.275 162.335 ;
        RECT 47.100 162.195 47.275 162.305 ;
        RECT 48.940 162.195 49.060 162.305 ;
        RECT 47.105 162.145 47.275 162.195 ;
        RECT 49.865 162.145 50.035 162.335 ;
        RECT 50.335 162.165 50.505 162.355 ;
        RECT 50.785 162.165 50.955 162.355 ;
        RECT 53.540 162.195 53.660 162.305 ;
        RECT 54.920 162.165 55.090 162.355 ;
        RECT 55.390 162.305 55.560 162.355 ;
        RECT 55.380 162.195 55.560 162.305 ;
        RECT 55.390 162.165 55.560 162.195 ;
        RECT 56.770 162.145 56.940 162.335 ;
        RECT 57.685 162.305 57.855 162.335 ;
        RECT 57.220 162.195 57.340 162.305 ;
        RECT 57.680 162.195 57.855 162.305 ;
        RECT 57.685 162.145 57.855 162.195 ;
        RECT 61.365 162.165 61.535 162.355 ;
        RECT 61.820 162.195 61.940 162.305 ;
        RECT 63.205 162.165 63.375 162.335 ;
        RECT 63.205 162.145 63.370 162.165 ;
        RECT 63.665 162.145 63.835 162.335 ;
        RECT 64.125 162.165 64.295 162.355 ;
        RECT 64.585 162.165 64.755 162.355 ;
        RECT 65.500 162.145 65.670 162.335 ;
        RECT 66.885 162.145 67.055 162.335 ;
        RECT 70.105 162.165 70.275 162.355 ;
        RECT 71.485 162.165 71.655 162.355 ;
        RECT 23.505 161.335 24.875 162.145 ;
        RECT 24.885 161.335 30.395 162.145 ;
        RECT 30.405 161.335 35.915 162.145 ;
        RECT 35.925 161.335 37.755 162.145 ;
        RECT 38.225 161.465 40.055 162.145 ;
        RECT 40.065 161.335 42.815 162.145 ;
        RECT 43.025 161.325 44.955 162.145 ;
        RECT 45.125 161.465 46.955 162.145 ;
        RECT 46.965 161.335 48.795 162.145 ;
        RECT 43.025 161.235 43.975 161.325 ;
        RECT 49.275 161.275 49.705 162.060 ;
        RECT 49.725 161.335 55.235 162.145 ;
        RECT 55.705 161.235 57.055 162.145 ;
        RECT 57.545 161.235 61.215 162.145 ;
        RECT 61.535 161.465 63.370 162.145 ;
        RECT 61.535 161.235 62.465 161.465 ;
        RECT 63.540 161.235 65.355 162.145 ;
        RECT 65.385 161.235 66.735 162.145 ;
        RECT 66.745 161.335 72.255 162.145 ;
        RECT 72.410 162.115 72.580 162.335 ;
        RECT 74.245 162.165 74.415 162.355 ;
        RECT 75.625 162.145 75.795 162.335 ;
        RECT 76.095 162.200 76.255 162.310 ;
        RECT 77.005 162.165 77.175 162.355 ;
        RECT 77.925 162.145 78.095 162.335 ;
        RECT 79.305 162.165 79.475 162.355 ;
        RECT 79.770 162.165 79.940 162.355 ;
        RECT 80.225 162.145 80.395 162.335 ;
        RECT 82.985 162.145 83.155 162.335 ;
        RECT 83.435 162.145 83.605 162.335 ;
        RECT 85.285 162.165 85.455 162.355 ;
        RECT 85.605 162.315 86.495 163.265 ;
        RECT 86.525 162.355 87.895 163.135 ;
        RECT 87.915 162.440 88.345 163.225 ;
        RECT 89.285 162.585 91.120 163.265 ;
        RECT 89.430 162.355 91.120 162.585 ;
        RECT 92.585 162.355 94.795 163.265 ;
        RECT 94.815 162.355 97.555 163.035 ;
        RECT 97.565 162.355 100.775 163.265 ;
        RECT 101.630 163.035 104.455 163.265 ;
        RECT 100.925 162.355 104.455 163.035 ;
        RECT 104.550 162.355 113.655 163.035 ;
        RECT 113.675 162.440 114.105 163.225 ;
        RECT 133.470 163.035 134.815 163.265 ;
        RECT 114.125 162.355 123.230 163.035 ;
        RECT 123.410 162.355 132.515 163.035 ;
        RECT 132.985 162.355 134.815 163.035 ;
        RECT 134.825 162.355 136.195 163.165 ;
        RECT 86.205 162.165 86.375 162.315 ;
        RECT 86.665 162.145 86.835 162.355 ;
        RECT 88.045 162.145 88.215 162.335 ;
        RECT 88.515 162.200 88.675 162.310 ;
        RECT 89.430 162.165 89.600 162.355 ;
        RECT 90.810 162.145 90.980 162.335 ;
        RECT 91.735 162.200 91.895 162.310 ;
        RECT 94.480 162.165 94.650 162.355 ;
        RECT 96.325 162.145 96.495 162.335 ;
        RECT 96.790 162.145 96.960 162.335 ;
        RECT 97.245 162.165 97.415 162.355 ;
        RECT 97.710 162.165 97.880 162.355 ;
        RECT 100.925 162.335 101.125 162.355 ;
        RECT 100.925 162.165 101.095 162.335 ;
        RECT 101.390 162.145 101.560 162.335 ;
        RECT 106.450 162.145 106.620 162.335 ;
        RECT 109.665 162.145 109.835 162.335 ;
        RECT 113.345 162.165 113.515 162.355 ;
        RECT 114.265 162.165 114.435 162.355 ;
        RECT 118.870 162.145 119.040 162.335 ;
        RECT 123.010 162.145 123.180 162.335 ;
        RECT 127.155 162.190 127.315 162.300 ;
        RECT 128.065 162.145 128.235 162.335 ;
        RECT 132.205 162.165 132.375 162.355 ;
        RECT 132.660 162.195 132.780 162.305 ;
        RECT 133.125 162.165 133.295 162.355 ;
        RECT 133.585 162.145 133.755 162.335 ;
        RECT 135.885 162.145 136.055 162.355 ;
        RECT 74.070 162.115 75.015 162.145 ;
        RECT 72.265 161.435 75.015 162.115 ;
        RECT 74.070 161.235 75.015 161.435 ;
        RECT 75.035 161.275 75.465 162.060 ;
        RECT 75.485 161.465 77.775 162.145 ;
        RECT 77.785 161.465 80.075 162.145 ;
        RECT 76.855 161.235 77.775 161.465 ;
        RECT 79.155 161.235 80.075 161.465 ;
        RECT 80.085 161.335 81.455 162.145 ;
        RECT 81.465 161.235 83.280 162.145 ;
        RECT 83.305 161.235 86.515 162.145 ;
        RECT 86.525 161.335 87.895 162.145 ;
        RECT 87.905 161.465 90.655 162.145 ;
        RECT 90.810 161.915 93.865 162.145 ;
        RECT 89.725 161.235 90.655 161.465 ;
        RECT 90.665 161.235 93.865 161.915 ;
        RECT 93.885 161.465 96.635 162.145 ;
        RECT 93.885 161.235 94.815 161.465 ;
        RECT 96.645 161.235 100.775 162.145 ;
        RECT 100.795 161.275 101.225 162.060 ;
        RECT 101.245 161.235 106.200 162.145 ;
        RECT 106.450 161.915 109.505 162.145 ;
        RECT 106.305 161.235 109.505 161.915 ;
        RECT 109.525 161.465 118.630 162.145 ;
        RECT 118.725 161.235 122.855 162.145 ;
        RECT 122.865 161.235 126.530 162.145 ;
        RECT 126.555 161.275 126.985 162.060 ;
        RECT 127.925 161.235 133.235 162.145 ;
        RECT 133.455 161.235 134.805 162.145 ;
        RECT 134.825 161.335 136.195 162.145 ;
      LAYER nwell ;
        RECT 23.310 158.115 136.390 160.945 ;
      LAYER pwell ;
        RECT 23.505 156.915 24.875 157.725 ;
        RECT 24.885 156.915 30.395 157.725 ;
        RECT 30.405 156.915 35.915 157.725 ;
        RECT 36.395 157.000 36.825 157.785 ;
        RECT 36.845 156.915 42.355 157.725 ;
        RECT 42.365 156.915 47.875 157.725 ;
        RECT 47.885 156.915 53.395 157.725 ;
        RECT 53.405 156.915 55.220 157.825 ;
        RECT 55.255 156.915 57.985 157.825 ;
        RECT 58.925 156.915 62.135 157.825 ;
        RECT 62.155 157.000 62.585 157.785 ;
        RECT 62.605 156.915 65.815 157.825 ;
        RECT 65.835 156.915 68.565 157.825 ;
        RECT 68.595 156.915 69.945 157.825 ;
        RECT 71.335 157.595 72.255 157.825 ;
        RECT 69.965 156.915 72.255 157.595 ;
        RECT 72.265 156.915 75.475 157.825 ;
        RECT 76.855 157.595 77.775 157.825 ;
        RECT 79.120 157.625 80.075 157.825 ;
        RECT 75.485 156.915 77.775 157.595 ;
        RECT 77.795 156.945 80.075 157.625 ;
        RECT 23.645 156.705 23.815 156.915 ;
        RECT 25.025 156.725 25.195 156.915 ;
        RECT 25.945 156.725 26.115 156.895 ;
        RECT 26.405 156.705 26.575 156.895 ;
        RECT 30.545 156.725 30.715 156.915 ;
        RECT 31.925 156.705 32.095 156.895 ;
        RECT 36.060 156.755 36.180 156.865 ;
        RECT 36.985 156.725 37.155 156.915 ;
        RECT 37.445 156.705 37.615 156.895 ;
        RECT 42.505 156.725 42.675 156.915 ;
        RECT 42.965 156.705 43.135 156.895 ;
        RECT 48.025 156.725 48.195 156.915 ;
        RECT 48.495 156.750 48.655 156.860 ;
        RECT 49.875 156.750 50.035 156.860 ;
        RECT 52.165 156.705 52.335 156.895 ;
        RECT 52.630 156.705 52.800 156.895 ;
        RECT 54.925 156.725 55.095 156.915 ;
        RECT 57.685 156.725 57.855 156.915 ;
        RECT 58.145 156.705 58.315 156.895 ;
        RECT 59.985 156.705 60.155 156.895 ;
        RECT 23.505 155.895 24.875 156.705 ;
        RECT 26.265 155.895 31.775 156.705 ;
        RECT 31.785 155.895 37.295 156.705 ;
        RECT 37.305 155.895 42.815 156.705 ;
        RECT 42.825 155.895 48.335 156.705 ;
        RECT 49.275 155.835 49.705 156.620 ;
        RECT 50.645 156.025 52.475 156.705 ;
        RECT 52.485 156.025 56.580 156.705 ;
        RECT 50.645 155.795 51.990 156.025 ;
        RECT 52.970 155.795 56.580 156.025 ;
        RECT 56.625 156.025 58.455 156.705 ;
        RECT 58.465 156.025 60.295 156.705 ;
        RECT 60.450 156.475 60.620 156.895 ;
        RECT 61.825 156.725 61.995 156.915 ;
        RECT 65.505 156.725 65.675 156.915 ;
        RECT 68.265 156.725 68.435 156.915 ;
        RECT 68.725 156.895 68.895 156.915 ;
        RECT 68.720 156.725 68.895 156.895 ;
        RECT 69.180 156.755 69.300 156.865 ;
        RECT 68.720 156.705 68.890 156.725 ;
        RECT 69.655 156.705 69.825 156.895 ;
        RECT 70.105 156.725 70.275 156.915 ;
        RECT 71.945 156.705 72.115 156.895 ;
        RECT 72.415 156.705 72.585 156.895 ;
        RECT 74.700 156.705 74.870 156.895 ;
        RECT 75.165 156.725 75.335 156.915 ;
        RECT 75.625 156.725 75.795 156.915 ;
        RECT 77.920 156.725 78.090 156.945 ;
        RECT 79.120 156.915 80.075 156.945 ;
        RECT 80.225 156.915 83.675 157.825 ;
        RECT 83.895 156.915 86.895 157.825 ;
        RECT 87.915 157.000 88.345 157.785 ;
        RECT 88.375 156.915 91.310 157.825 ;
        RECT 92.045 157.145 95.245 157.825 ;
        RECT 95.750 157.595 97.090 157.825 ;
        RECT 83.445 156.895 83.615 156.915 ;
        RECT 78.845 156.705 79.015 156.895 ;
        RECT 79.315 156.750 79.475 156.860 ;
        RECT 81.145 156.705 81.315 156.895 ;
        RECT 83.445 156.725 83.620 156.895 ;
        RECT 61.730 156.475 64.890 156.705 ;
        RECT 60.345 156.025 64.890 156.475 ;
        RECT 56.625 155.795 57.970 156.025 ;
        RECT 58.465 155.795 59.810 156.025 ;
        RECT 60.345 155.795 61.720 156.025 ;
        RECT 63.510 155.795 64.890 156.025 ;
        RECT 64.940 156.025 69.035 156.705 ;
        RECT 64.940 155.795 68.550 156.025 ;
        RECT 69.505 155.925 70.875 156.705 ;
        RECT 70.895 155.795 72.245 156.705 ;
        RECT 72.265 155.925 73.635 156.705 ;
        RECT 73.665 155.795 75.015 156.705 ;
        RECT 75.035 155.835 75.465 156.620 ;
        RECT 75.625 155.795 79.075 156.705 ;
        RECT 80.095 155.795 81.445 156.705 ;
        RECT 81.465 156.675 82.420 156.705 ;
        RECT 83.450 156.675 83.620 156.725 ;
        RECT 86.205 156.725 86.375 156.895 ;
        RECT 86.665 156.725 86.835 156.915 ;
        RECT 91.265 156.895 91.310 156.915 ;
        RECT 92.190 156.915 95.245 157.145 ;
        RECT 95.265 156.915 99.855 157.595 ;
        RECT 100.325 156.915 103.980 157.825 ;
        RECT 104.090 156.915 113.195 157.595 ;
        RECT 113.675 157.000 114.105 157.785 ;
        RECT 114.125 156.915 123.230 157.595 ;
        RECT 123.325 156.915 132.430 157.595 ;
        RECT 132.525 156.915 134.735 157.825 ;
        RECT 134.825 156.915 136.195 157.725 ;
        RECT 87.135 156.760 87.295 156.870 ;
        RECT 89.425 156.725 89.595 156.895 ;
        RECT 86.205 156.705 86.345 156.725 ;
        RECT 89.425 156.705 89.470 156.725 ;
        RECT 89.885 156.705 90.055 156.895 ;
        RECT 91.265 156.725 91.435 156.895 ;
        RECT 91.720 156.755 91.840 156.865 ;
        RECT 92.190 156.725 92.360 156.915 ;
        RECT 95.410 156.725 95.580 156.915 ;
        RECT 100.470 156.895 100.640 156.915 ;
        RECT 100.000 156.755 100.120 156.865 ;
        RECT 100.465 156.725 100.640 156.895 ;
        RECT 100.465 156.705 100.635 156.725 ;
        RECT 101.390 156.705 101.560 156.895 ;
        RECT 105.060 156.755 105.180 156.865 ;
        RECT 112.885 156.725 113.055 156.915 ;
        RECT 113.340 156.755 113.460 156.865 ;
        RECT 114.265 156.705 114.435 156.915 ;
        RECT 81.465 155.995 83.745 156.675 ;
        RECT 81.465 155.795 82.420 155.995 ;
        RECT 83.775 155.885 86.345 156.705 ;
        RECT 83.775 155.795 85.365 155.885 ;
        RECT 86.535 155.795 89.470 156.705 ;
        RECT 89.745 156.025 91.575 156.705 ;
        RECT 91.670 156.025 100.775 156.705 ;
        RECT 90.230 155.795 91.575 156.025 ;
        RECT 100.795 155.835 101.225 156.620 ;
        RECT 101.250 155.795 104.835 156.705 ;
        RECT 105.470 156.025 114.575 156.705 ;
        RECT 114.725 156.675 114.895 156.895 ;
        RECT 117.485 156.705 117.655 156.895 ;
        RECT 123.465 156.725 123.635 156.915 ;
        RECT 127.145 156.705 127.315 156.895 ;
        RECT 130.360 156.755 130.480 156.865 ;
        RECT 132.670 156.725 132.840 156.915 ;
        RECT 134.045 156.705 134.215 156.895 ;
        RECT 134.500 156.755 134.620 156.865 ;
        RECT 135.885 156.705 136.055 156.915 ;
        RECT 115.940 156.675 117.335 156.705 ;
        RECT 114.600 155.995 117.335 156.675 ;
        RECT 117.345 156.025 126.450 156.705 ;
        RECT 115.925 155.795 117.335 155.995 ;
        RECT 126.555 155.835 126.985 156.620 ;
        RECT 127.005 155.795 130.215 156.705 ;
        RECT 130.825 155.795 134.275 156.705 ;
        RECT 134.825 155.895 136.195 156.705 ;
      LAYER nwell ;
        RECT 23.310 152.675 136.390 155.505 ;
      LAYER pwell ;
        RECT 23.505 151.475 24.875 152.285 ;
        RECT 24.885 151.475 30.395 152.285 ;
        RECT 30.405 151.475 35.915 152.285 ;
        RECT 36.395 151.560 36.825 152.345 ;
        RECT 37.765 151.475 39.135 152.255 ;
        RECT 39.145 151.475 40.975 152.285 ;
        RECT 40.985 151.475 42.355 152.255 ;
        RECT 42.365 151.475 44.195 152.285 ;
        RECT 44.690 152.155 46.035 152.385 ;
        RECT 44.205 151.475 46.035 152.155 ;
        RECT 46.045 151.475 47.415 152.285 ;
        RECT 47.425 151.475 48.795 152.255 ;
        RECT 49.275 151.560 49.705 152.345 ;
        RECT 49.725 151.475 51.555 152.285 ;
        RECT 51.600 152.155 52.975 152.385 ;
        RECT 54.745 152.155 55.695 152.385 ;
        RECT 51.600 151.705 55.695 152.155 ;
        RECT 23.645 151.285 23.815 151.475 ;
        RECT 25.025 151.285 25.195 151.475 ;
        RECT 30.545 151.285 30.715 151.475 ;
        RECT 36.060 151.315 36.180 151.425 ;
        RECT 36.995 151.320 37.155 151.430 ;
        RECT 37.915 151.285 38.085 151.475 ;
        RECT 39.285 151.285 39.455 151.475 ;
        RECT 41.125 151.285 41.295 151.475 ;
        RECT 42.505 151.285 42.675 151.475 ;
        RECT 44.345 151.285 44.515 151.475 ;
        RECT 46.185 151.285 46.355 151.475 ;
        RECT 47.575 151.285 47.745 151.475 ;
        RECT 48.940 151.315 49.060 151.425 ;
        RECT 49.865 151.285 50.035 151.475 ;
        RECT 51.705 151.285 51.875 151.705 ;
        RECT 52.985 151.475 55.695 151.705 ;
        RECT 55.705 151.475 57.535 152.155 ;
        RECT 57.545 151.475 58.915 152.255 ;
        RECT 55.845 151.285 56.015 151.475 ;
        RECT 57.695 151.285 57.865 151.475 ;
        RECT 59.845 151.435 60.735 152.385 ;
        RECT 60.765 151.475 62.135 152.255 ;
        RECT 62.155 151.560 62.585 152.345 ;
        RECT 64.010 152.155 65.355 152.385 ;
        RECT 63.525 151.475 65.355 152.155 ;
        RECT 65.365 151.475 66.735 152.255 ;
        RECT 68.125 151.475 69.495 152.255 ;
        RECT 69.645 151.475 72.255 152.385 ;
        RECT 72.265 151.475 73.635 152.255 ;
        RECT 73.645 151.475 75.015 152.255 ;
        RECT 75.035 151.560 75.465 152.345 ;
        RECT 76.405 151.475 77.775 152.255 ;
        RECT 77.785 151.475 79.155 152.255 ;
        RECT 79.185 151.475 80.535 152.385 ;
        RECT 81.005 152.155 82.350 152.385 ;
        RECT 81.005 151.475 82.835 152.155 ;
        RECT 82.925 151.475 85.135 152.385 ;
        RECT 85.155 151.475 87.895 152.155 ;
        RECT 87.915 151.560 88.345 152.345 ;
        RECT 88.375 151.705 91.575 152.385 ;
        RECT 88.375 151.475 91.430 151.705 ;
        RECT 91.670 151.475 100.775 152.155 ;
        RECT 100.795 151.560 101.225 152.345 ;
        RECT 101.330 151.475 110.435 152.155 ;
        RECT 110.455 151.705 113.655 152.385 ;
        RECT 110.455 151.475 113.510 151.705 ;
        RECT 113.675 151.560 114.105 152.345 ;
        RECT 114.125 151.475 117.165 152.385 ;
        RECT 117.430 151.475 126.535 152.155 ;
        RECT 126.555 151.560 126.985 152.345 ;
        RECT 127.665 152.155 131.595 152.385 ;
        RECT 127.180 151.475 131.595 152.155 ;
        RECT 131.735 151.475 134.735 152.385 ;
        RECT 134.825 151.475 136.195 152.285 ;
        RECT 59.075 151.320 59.235 151.430 ;
        RECT 60.445 151.285 60.615 151.435 ;
        RECT 60.915 151.285 61.085 151.475 ;
        RECT 62.755 151.320 62.915 151.430 ;
        RECT 63.665 151.285 63.835 151.475 ;
        RECT 65.515 151.285 65.685 151.475 ;
        RECT 67.805 151.285 67.975 151.455 ;
        RECT 68.275 151.285 68.445 151.475 ;
        RECT 71.940 151.285 72.110 151.475 ;
        RECT 72.415 151.285 72.585 151.475 ;
        RECT 73.795 151.285 73.965 151.475 ;
        RECT 75.635 151.320 75.795 151.430 ;
        RECT 76.555 151.285 76.725 151.475 ;
        RECT 77.935 151.285 78.105 151.475 ;
        RECT 80.220 151.285 80.390 151.475 ;
        RECT 80.680 151.315 80.800 151.425 ;
        RECT 82.525 151.285 82.695 151.475 ;
        RECT 84.820 151.285 84.990 151.475 ;
        RECT 87.585 151.285 87.755 151.475 ;
        RECT 91.260 151.285 91.430 151.475 ;
        RECT 100.465 151.285 100.635 151.475 ;
        RECT 110.125 151.285 110.295 151.475 ;
        RECT 113.340 151.285 113.510 151.475 ;
        RECT 117.020 151.455 117.165 151.475 ;
        RECT 117.020 151.285 117.190 151.455 ;
        RECT 126.225 151.285 126.395 151.475 ;
        RECT 127.180 151.455 127.290 151.475 ;
        RECT 127.120 151.285 127.290 151.455 ;
        RECT 134.505 151.285 134.675 151.475 ;
        RECT 135.885 151.285 136.055 151.475 ;
        RECT 1.290 52.730 13.780 58.190 ;
        RECT 46.010 57.320 50.180 69.810 ;
      LAYER nwell ;
        RECT 50.300 61.620 52.410 69.810 ;
      LAYER pwell ;
        RECT 50.280 57.325 52.390 61.425 ;
        RECT 52.475 57.335 58.465 69.825 ;
      LAYER nwell ;
        RECT 58.595 61.635 60.705 69.825 ;
      LAYER pwell ;
        RECT 58.585 57.325 60.695 61.425 ;
        RECT 60.805 57.325 66.795 69.815 ;
      LAYER nwell ;
        RECT 66.910 61.625 69.020 69.815 ;
      LAYER pwell ;
        RECT 66.845 57.325 68.955 61.425 ;
        RECT 69.100 57.315 75.090 69.805 ;
      LAYER nwell ;
        RECT 75.290 61.725 77.400 69.915 ;
      LAYER pwell ;
        RECT 75.265 57.345 77.375 61.445 ;
        RECT 77.545 57.330 83.535 69.820 ;
      LAYER nwell ;
        RECT 83.680 61.650 85.790 69.840 ;
      LAYER pwell ;
        RECT 83.615 57.325 85.725 61.425 ;
        RECT 85.875 57.330 91.865 69.820 ;
      LAYER nwell ;
        RECT 92.010 61.675 94.120 69.865 ;
      LAYER pwell ;
        RECT 92.000 57.320 94.110 61.420 ;
        RECT 94.205 57.330 100.195 69.820 ;
      LAYER nwell ;
        RECT 100.305 61.690 102.415 69.880 ;
      LAYER pwell ;
        RECT 100.240 57.330 102.350 61.430 ;
        RECT 102.510 57.325 108.500 69.815 ;
      LAYER nwell ;
        RECT 108.605 61.670 110.715 69.860 ;
      LAYER pwell ;
        RECT 108.605 57.330 110.715 61.430 ;
        RECT 110.810 57.335 114.980 69.825 ;
        RECT 1.290 50.380 31.720 52.730 ;
        RECT 43.310 50.380 61.780 52.730 ;
        RECT 67.310 50.380 85.780 52.730 ;
      LAYER nwell ;
        RECT 27.290 49.600 29.790 49.880 ;
        RECT 55.790 49.600 58.290 49.880 ;
        RECT 83.290 49.600 85.790 49.880 ;
        RECT 111.790 49.600 114.290 49.880 ;
        RECT 5.410 49.355 12.800 49.585 ;
        RECT 1.290 47.890 12.800 49.355 ;
        RECT 26.050 49.355 29.790 49.600 ;
        RECT 33.410 49.355 40.800 49.585 ;
        RECT 26.050 47.890 40.800 49.355 ;
        RECT 54.050 49.355 58.290 49.600 ;
        RECT 61.410 49.355 68.800 49.585 ;
        RECT 54.050 47.890 68.800 49.355 ;
        RECT 82.050 49.355 85.790 49.600 ;
        RECT 89.410 49.355 96.800 49.585 ;
        RECT 82.050 47.890 96.800 49.355 ;
        RECT 110.050 49.355 114.290 49.600 ;
        RECT 117.410 49.355 124.800 49.585 ;
        RECT 110.050 47.890 124.800 49.355 ;
        RECT 1.290 45.580 21.135 47.890 ;
        RECT 26.050 45.595 49.135 47.890 ;
        RECT 54.050 45.595 77.135 47.890 ;
        RECT 82.050 45.595 105.135 47.890 ;
        RECT 110.050 45.595 133.135 47.890 ;
        RECT 138.050 45.595 140.160 49.600 ;
        RECT 24.025 45.580 49.135 45.595 ;
        RECT 52.025 45.580 77.135 45.595 ;
        RECT 80.025 45.580 105.135 45.595 ;
        RECT 108.025 45.580 133.135 45.595 ;
        RECT 136.025 45.580 140.160 45.595 ;
        RECT 1.290 39.410 140.160 45.580 ;
      LAYER pwell ;
        RECT 143.290 44.730 149.800 50.190 ;
        RECT 143.290 40.560 155.780 44.730 ;
      LAYER nwell ;
        RECT 1.290 39.405 26.135 39.410 ;
        RECT 27.440 39.405 54.135 39.410 ;
        RECT 55.790 39.405 82.135 39.410 ;
        RECT 84.280 39.405 110.135 39.410 ;
        RECT 111.790 39.405 138.135 39.410 ;
        RECT 1.290 39.395 24.110 39.405 ;
        RECT 12.720 39.390 24.110 39.395 ;
        RECT 27.545 39.395 52.110 39.405 ;
        RECT 27.545 39.390 29.790 39.395 ;
        RECT 40.720 39.390 52.110 39.395 ;
        RECT 55.790 39.395 80.110 39.405 ;
        RECT 55.790 39.380 58.290 39.395 ;
        RECT 68.720 39.390 80.110 39.395 ;
        RECT 84.850 39.395 108.110 39.405 ;
        RECT 84.850 39.380 85.790 39.395 ;
        RECT 96.720 39.390 108.110 39.395 ;
        RECT 111.790 39.395 136.110 39.405 ;
        RECT 111.790 39.380 114.290 39.395 ;
        RECT 124.720 39.390 136.110 39.395 ;
      LAYER pwell ;
        RECT 26.135 39.020 28.245 39.025 ;
        RECT 54.135 39.020 56.245 39.025 ;
        RECT 82.135 39.020 84.245 39.025 ;
        RECT 110.135 39.020 112.245 39.025 ;
        RECT 138.135 39.020 140.245 39.025 ;
        RECT 24.110 39.015 28.245 39.020 ;
        RECT 52.110 39.015 56.245 39.020 ;
        RECT 80.110 39.015 84.245 39.020 ;
        RECT 108.110 39.015 112.245 39.020 ;
        RECT 136.110 39.015 140.245 39.020 ;
        RECT 1.950 35.920 28.245 39.015 ;
        RECT 1.950 34.915 24.200 35.920 ;
        RECT 26.135 34.925 28.245 35.920 ;
        RECT 29.950 35.920 56.245 39.015 ;
        RECT 29.950 34.915 52.200 35.920 ;
        RECT 54.135 34.925 56.245 35.920 ;
        RECT 57.950 35.920 84.245 39.015 ;
        RECT 57.950 34.915 80.200 35.920 ;
        RECT 82.135 34.925 84.245 35.920 ;
        RECT 85.950 35.920 112.245 39.015 ;
        RECT 85.950 34.915 108.200 35.920 ;
        RECT 110.135 34.925 112.245 35.920 ;
        RECT 113.950 35.920 140.245 39.015 ;
        RECT 113.950 34.915 136.200 35.920 ;
        RECT 138.135 34.925 140.245 35.920 ;
      LAYER nwell ;
        RECT 27.290 33.600 29.790 33.880 ;
        RECT 55.290 33.600 57.790 33.880 ;
        RECT 83.790 33.600 86.290 33.880 ;
        RECT 111.790 33.600 114.290 33.880 ;
        RECT 5.410 33.355 12.800 33.585 ;
        RECT 1.290 31.890 12.800 33.355 ;
        RECT 26.050 33.355 29.790 33.600 ;
        RECT 33.410 33.355 40.800 33.585 ;
        RECT 26.050 31.890 40.800 33.355 ;
        RECT 54.050 33.355 57.790 33.600 ;
        RECT 61.410 33.355 68.800 33.585 ;
        RECT 54.050 31.890 68.800 33.355 ;
        RECT 82.050 33.355 86.290 33.600 ;
        RECT 89.410 33.355 96.800 33.585 ;
        RECT 82.050 31.890 96.800 33.355 ;
        RECT 110.050 33.355 114.290 33.600 ;
        RECT 117.410 33.355 124.800 33.585 ;
        RECT 110.050 31.890 124.800 33.355 ;
        RECT 1.290 29.580 21.135 31.890 ;
        RECT 26.050 29.595 49.135 31.890 ;
        RECT 54.050 29.595 77.135 31.890 ;
        RECT 82.050 29.595 105.135 31.890 ;
        RECT 110.050 29.595 133.135 31.890 ;
        RECT 138.050 29.595 140.160 33.600 ;
        RECT 24.025 29.580 49.135 29.595 ;
        RECT 52.025 29.580 77.135 29.595 ;
        RECT 80.025 29.580 105.135 29.595 ;
        RECT 108.025 29.580 133.135 29.595 ;
        RECT 136.025 29.580 140.160 29.595 ;
        RECT 1.290 23.410 140.160 29.580 ;
        RECT 1.290 23.405 26.135 23.410 ;
        RECT 28.755 23.405 54.135 23.410 ;
        RECT 56.840 23.405 82.135 23.410 ;
        RECT 83.790 23.405 110.135 23.410 ;
        RECT 111.790 23.405 138.135 23.410 ;
        RECT 1.290 23.395 24.110 23.405 ;
        RECT 12.720 23.390 24.110 23.395 ;
        RECT 28.755 23.395 52.110 23.405 ;
        RECT 28.755 23.380 29.790 23.395 ;
        RECT 40.720 23.390 52.110 23.395 ;
        RECT 56.840 23.395 80.110 23.405 ;
        RECT 56.840 23.380 57.790 23.395 ;
        RECT 68.720 23.390 80.110 23.395 ;
        RECT 83.790 23.395 108.110 23.405 ;
        RECT 83.790 23.380 86.290 23.395 ;
        RECT 96.720 23.390 108.110 23.395 ;
        RECT 111.790 23.395 136.110 23.405 ;
        RECT 111.790 23.380 114.290 23.395 ;
        RECT 124.720 23.390 136.110 23.395 ;
      LAYER pwell ;
        RECT 26.135 23.020 28.245 23.025 ;
        RECT 54.135 23.020 56.245 23.025 ;
        RECT 82.135 23.020 84.245 23.025 ;
        RECT 110.135 23.020 112.245 23.025 ;
        RECT 138.135 23.020 140.245 23.025 ;
        RECT 24.110 23.015 28.245 23.020 ;
        RECT 52.110 23.015 56.245 23.020 ;
        RECT 80.110 23.015 84.245 23.020 ;
        RECT 108.110 23.015 112.245 23.020 ;
        RECT 136.110 23.015 140.245 23.020 ;
        RECT 1.950 19.920 28.245 23.015 ;
        RECT 1.950 18.915 24.200 19.920 ;
        RECT 26.135 18.925 28.245 19.920 ;
        RECT 29.950 19.920 56.245 23.015 ;
        RECT 29.950 18.915 52.200 19.920 ;
        RECT 54.135 18.925 56.245 19.920 ;
        RECT 57.950 19.920 84.245 23.015 ;
        RECT 57.950 18.915 80.200 19.920 ;
        RECT 82.135 18.925 84.245 19.920 ;
        RECT 85.950 19.920 112.245 23.015 ;
        RECT 85.950 18.915 108.200 19.920 ;
        RECT 110.135 18.925 112.245 19.920 ;
        RECT 113.950 19.920 140.245 23.015 ;
        RECT 113.950 18.915 136.200 19.920 ;
        RECT 138.135 18.925 140.245 19.920 ;
      LAYER nwell ;
        RECT 27.790 17.600 30.290 17.880 ;
        RECT 55.290 17.600 57.790 17.880 ;
        RECT 83.790 17.600 86.290 17.880 ;
        RECT 111.790 17.600 114.290 17.880 ;
        RECT 5.410 17.355 12.800 17.585 ;
        RECT 1.290 15.890 12.800 17.355 ;
        RECT 26.050 17.355 30.290 17.600 ;
        RECT 33.410 17.355 40.800 17.585 ;
        RECT 26.050 15.890 40.800 17.355 ;
        RECT 54.050 17.355 57.790 17.600 ;
        RECT 61.410 17.355 68.800 17.585 ;
        RECT 54.050 15.890 68.800 17.355 ;
        RECT 82.050 17.355 86.290 17.600 ;
        RECT 89.410 17.355 96.800 17.585 ;
        RECT 82.050 15.890 96.800 17.355 ;
        RECT 110.050 17.355 114.290 17.600 ;
        RECT 117.410 17.355 124.800 17.585 ;
        RECT 110.050 15.890 124.800 17.355 ;
        RECT 1.290 13.580 21.135 15.890 ;
        RECT 26.050 13.595 49.135 15.890 ;
        RECT 54.050 13.595 77.135 15.890 ;
        RECT 82.050 13.595 105.135 15.890 ;
        RECT 110.050 13.595 133.135 15.890 ;
        RECT 138.050 13.595 140.160 17.600 ;
        RECT 24.025 13.580 49.135 13.595 ;
        RECT 52.025 13.580 77.135 13.595 ;
        RECT 80.025 13.580 105.135 13.595 ;
        RECT 108.025 13.580 133.135 13.595 ;
        RECT 136.025 13.580 140.160 13.595 ;
        RECT 1.290 7.410 140.160 13.580 ;
        RECT 1.290 7.405 26.135 7.410 ;
        RECT 27.790 7.405 54.135 7.410 ;
        RECT 55.495 7.405 82.135 7.410 ;
        RECT 83.790 7.405 110.135 7.410 ;
        RECT 111.790 7.405 138.135 7.410 ;
        RECT 1.290 7.395 24.110 7.405 ;
        RECT 12.720 7.390 24.110 7.395 ;
        RECT 27.790 7.395 52.110 7.405 ;
        RECT 57.115 7.400 80.110 7.405 ;
        RECT 57.290 7.395 80.110 7.400 ;
        RECT 27.790 7.380 30.290 7.395 ;
        RECT 40.720 7.390 52.110 7.395 ;
        RECT 68.720 7.390 80.110 7.395 ;
        RECT 83.790 7.395 108.110 7.405 ;
        RECT 83.790 7.380 86.290 7.395 ;
        RECT 96.720 7.390 108.110 7.395 ;
        RECT 111.790 7.395 136.110 7.405 ;
        RECT 111.790 7.380 114.290 7.395 ;
        RECT 124.720 7.390 136.110 7.395 ;
      LAYER pwell ;
        RECT 26.135 7.020 28.245 7.025 ;
        RECT 54.135 7.020 56.245 7.025 ;
        RECT 82.135 7.020 84.245 7.025 ;
        RECT 110.135 7.020 112.245 7.025 ;
        RECT 138.135 7.020 140.245 7.025 ;
        RECT 24.110 7.015 28.245 7.020 ;
        RECT 52.110 7.015 56.245 7.020 ;
        RECT 80.110 7.015 84.245 7.020 ;
        RECT 108.110 7.015 112.245 7.020 ;
        RECT 136.110 7.015 140.245 7.020 ;
        RECT 1.950 3.920 28.245 7.015 ;
        RECT 1.950 2.915 24.200 3.920 ;
        RECT 26.135 2.925 28.245 3.920 ;
        RECT 29.950 3.920 56.245 7.015 ;
        RECT 29.950 2.915 52.200 3.920 ;
        RECT 54.135 2.925 56.245 3.920 ;
        RECT 57.950 3.920 84.245 7.015 ;
        RECT 57.950 2.915 80.200 3.920 ;
        RECT 82.135 2.925 84.245 3.920 ;
        RECT 85.950 3.920 112.245 7.015 ;
        RECT 85.950 2.915 108.200 3.920 ;
        RECT 110.135 2.925 112.245 3.920 ;
        RECT 113.950 3.920 140.245 7.015 ;
        RECT 113.950 2.915 136.200 3.920 ;
        RECT 138.135 2.925 140.245 3.920 ;
      LAYER li1 ;
        RECT 23.500 194.805 136.200 194.975 ;
        RECT 23.585 194.055 24.795 194.805 ;
        RECT 23.585 193.515 24.105 194.055 ;
        RECT 24.970 193.965 25.230 194.805 ;
        RECT 25.405 194.060 25.660 194.635 ;
        RECT 25.830 194.425 26.160 194.805 ;
        RECT 26.375 194.255 26.545 194.635 ;
        RECT 25.830 194.085 26.545 194.255 ;
        RECT 26.985 194.145 27.325 194.805 ;
        RECT 24.275 193.345 24.795 193.885 ;
        RECT 23.585 192.255 24.795 193.345 ;
        RECT 24.970 192.255 25.230 193.405 ;
        RECT 25.405 193.330 25.575 194.060 ;
        RECT 25.830 193.895 26.000 194.085 ;
        RECT 25.745 193.565 26.000 193.895 ;
        RECT 25.830 193.355 26.000 193.565 ;
        RECT 26.280 193.535 26.635 193.905 ;
        RECT 25.405 192.425 25.660 193.330 ;
        RECT 25.830 193.185 26.545 193.355 ;
        RECT 25.830 192.255 26.160 193.015 ;
        RECT 26.375 192.425 26.545 193.185 ;
        RECT 26.805 192.425 27.325 193.975 ;
        RECT 27.495 193.150 28.015 194.635 ;
        RECT 28.185 194.260 33.530 194.805 ;
        RECT 29.770 193.430 30.110 194.260 ;
        RECT 33.705 194.035 36.295 194.805 ;
        RECT 36.465 194.080 36.755 194.805 ;
        RECT 37.385 194.195 37.725 194.610 ;
        RECT 37.895 194.365 38.065 194.805 ;
        RECT 38.235 194.415 39.485 194.595 ;
        RECT 38.235 194.195 38.565 194.415 ;
        RECT 39.755 194.345 39.925 194.805 ;
        RECT 27.495 192.255 27.825 192.980 ;
        RECT 31.590 192.690 31.940 193.940 ;
        RECT 33.705 193.515 34.915 194.035 ;
        RECT 37.385 194.025 38.565 194.195 ;
        RECT 38.735 194.175 39.100 194.245 ;
        RECT 38.735 193.995 39.985 194.175 ;
        RECT 35.085 193.345 36.295 193.865 ;
        RECT 37.385 193.615 37.850 193.815 ;
        RECT 38.025 193.565 38.355 193.815 ;
        RECT 38.525 193.785 38.990 193.815 ;
        RECT 38.525 193.615 38.995 193.785 ;
        RECT 38.525 193.565 38.990 193.615 ;
        RECT 39.185 193.565 39.540 193.815 ;
        RECT 38.025 193.445 38.205 193.565 ;
        RECT 28.185 192.255 33.530 192.690 ;
        RECT 33.705 192.255 36.295 193.345 ;
        RECT 36.465 192.255 36.755 193.420 ;
        RECT 37.385 192.255 37.705 193.435 ;
        RECT 37.875 193.275 38.205 193.445 ;
        RECT 39.710 193.395 39.985 193.995 ;
        RECT 37.875 192.485 38.075 193.275 ;
        RECT 38.375 193.185 39.985 193.395 ;
        RECT 38.375 193.085 38.785 193.185 ;
        RECT 38.400 192.425 38.785 193.085 ;
        RECT 39.180 192.255 39.965 193.015 ;
        RECT 40.155 192.425 40.435 194.525 ;
        RECT 40.605 194.260 45.950 194.805 ;
        RECT 42.190 193.430 42.530 194.260 ;
        RECT 46.125 194.035 48.715 194.805 ;
        RECT 49.345 194.080 49.635 194.805 ;
        RECT 49.805 194.260 55.150 194.805 ;
        RECT 55.325 194.260 60.670 194.805 ;
        RECT 44.010 192.690 44.360 193.940 ;
        RECT 46.125 193.515 47.335 194.035 ;
        RECT 47.505 193.345 48.715 193.865 ;
        RECT 51.390 193.430 51.730 194.260 ;
        RECT 40.605 192.255 45.950 192.690 ;
        RECT 46.125 192.255 48.715 193.345 ;
        RECT 49.345 192.255 49.635 193.420 ;
        RECT 53.210 192.690 53.560 193.940 ;
        RECT 56.910 193.430 57.250 194.260 ;
        RECT 60.845 194.055 62.055 194.805 ;
        RECT 62.225 194.080 62.515 194.805 ;
        RECT 63.695 194.255 63.865 194.635 ;
        RECT 64.045 194.425 64.375 194.805 ;
        RECT 63.695 194.085 64.360 194.255 ;
        RECT 64.555 194.130 64.815 194.635 ;
        RECT 58.730 192.690 59.080 193.940 ;
        RECT 60.845 193.515 61.365 194.055 ;
        RECT 61.535 193.345 62.055 193.885 ;
        RECT 63.625 193.535 63.965 193.905 ;
        RECT 64.190 193.830 64.360 194.085 ;
        RECT 64.190 193.500 64.465 193.830 ;
        RECT 49.805 192.255 55.150 192.690 ;
        RECT 55.325 192.255 60.670 192.690 ;
        RECT 60.845 192.255 62.055 193.345 ;
        RECT 62.225 192.255 62.515 193.420 ;
        RECT 64.190 193.355 64.360 193.500 ;
        RECT 63.685 193.185 64.360 193.355 ;
        RECT 64.635 193.330 64.815 194.130 ;
        RECT 64.985 194.035 66.655 194.805 ;
        RECT 64.985 193.515 65.735 194.035 ;
        RECT 66.830 193.965 67.090 194.805 ;
        RECT 67.265 194.060 67.520 194.635 ;
        RECT 67.690 194.425 68.020 194.805 ;
        RECT 68.235 194.255 68.405 194.635 ;
        RECT 67.690 194.085 68.405 194.255 ;
        RECT 65.905 193.345 66.655 193.865 ;
        RECT 63.685 192.425 63.865 193.185 ;
        RECT 64.045 192.255 64.375 193.015 ;
        RECT 64.545 192.425 64.815 193.330 ;
        RECT 64.985 192.255 66.655 193.345 ;
        RECT 66.830 192.255 67.090 193.405 ;
        RECT 67.265 193.330 67.435 194.060 ;
        RECT 67.690 193.895 67.860 194.085 ;
        RECT 68.665 194.035 72.175 194.805 ;
        RECT 73.355 194.255 73.525 194.635 ;
        RECT 73.705 194.425 74.035 194.805 ;
        RECT 73.355 194.085 74.020 194.255 ;
        RECT 74.215 194.130 74.475 194.635 ;
        RECT 67.605 193.565 67.860 193.895 ;
        RECT 67.690 193.355 67.860 193.565 ;
        RECT 68.140 193.535 68.495 193.905 ;
        RECT 68.665 193.515 70.315 194.035 ;
        RECT 67.265 192.425 67.520 193.330 ;
        RECT 67.690 193.185 68.405 193.355 ;
        RECT 70.485 193.345 72.175 193.865 ;
        RECT 73.285 193.535 73.625 193.905 ;
        RECT 73.850 193.830 74.020 194.085 ;
        RECT 73.850 193.500 74.125 193.830 ;
        RECT 73.850 193.355 74.020 193.500 ;
        RECT 67.690 192.255 68.020 193.015 ;
        RECT 68.235 192.425 68.405 193.185 ;
        RECT 68.665 192.255 72.175 193.345 ;
        RECT 73.345 193.185 74.020 193.355 ;
        RECT 74.295 193.330 74.475 194.130 ;
        RECT 75.105 194.080 75.395 194.805 ;
        RECT 76.485 194.130 76.745 194.635 ;
        RECT 76.925 194.425 77.255 194.805 ;
        RECT 77.435 194.255 77.605 194.635 ;
        RECT 73.345 192.425 73.525 193.185 ;
        RECT 73.705 192.255 74.035 193.015 ;
        RECT 74.205 192.425 74.475 193.330 ;
        RECT 75.105 192.255 75.395 193.420 ;
        RECT 76.485 193.330 76.665 194.130 ;
        RECT 76.940 194.085 77.605 194.255 ;
        RECT 76.940 193.830 77.110 194.085 ;
        RECT 77.865 194.055 79.075 194.805 ;
        RECT 79.335 194.255 79.505 194.635 ;
        RECT 79.685 194.425 80.015 194.805 ;
        RECT 79.335 194.085 80.000 194.255 ;
        RECT 80.195 194.130 80.455 194.635 ;
        RECT 76.835 193.500 77.110 193.830 ;
        RECT 77.335 193.535 77.675 193.905 ;
        RECT 77.865 193.515 78.385 194.055 ;
        RECT 76.940 193.355 77.110 193.500 ;
        RECT 76.485 192.425 76.755 193.330 ;
        RECT 76.940 193.185 77.615 193.355 ;
        RECT 78.555 193.345 79.075 193.885 ;
        RECT 79.265 193.535 79.605 193.905 ;
        RECT 79.830 193.830 80.000 194.085 ;
        RECT 79.830 193.500 80.105 193.830 ;
        RECT 79.830 193.355 80.000 193.500 ;
        RECT 76.925 192.255 77.255 193.015 ;
        RECT 77.435 192.425 77.615 193.185 ;
        RECT 77.865 192.255 79.075 193.345 ;
        RECT 79.325 193.185 80.000 193.355 ;
        RECT 80.275 193.330 80.455 194.130 ;
        RECT 79.325 192.425 79.505 193.185 ;
        RECT 79.685 192.255 80.015 193.015 ;
        RECT 80.185 192.425 80.455 193.330 ;
        RECT 80.625 192.425 81.375 194.635 ;
        RECT 81.635 194.255 81.805 194.635 ;
        RECT 81.985 194.425 82.315 194.805 ;
        RECT 81.635 194.085 82.300 194.255 ;
        RECT 82.495 194.130 82.755 194.635 ;
        RECT 81.565 193.535 81.905 193.905 ;
        RECT 82.130 193.830 82.300 194.085 ;
        RECT 82.130 193.500 82.405 193.830 ;
        RECT 82.130 193.355 82.300 193.500 ;
        RECT 81.625 193.185 82.300 193.355 ;
        RECT 82.575 193.330 82.755 194.130 ;
        RECT 82.925 194.235 83.360 194.635 ;
        RECT 83.530 194.405 83.915 194.805 ;
        RECT 82.925 194.065 83.915 194.235 ;
        RECT 84.085 194.065 84.510 194.635 ;
        RECT 84.700 194.235 84.955 194.635 ;
        RECT 85.125 194.405 85.510 194.805 ;
        RECT 84.700 194.065 85.510 194.235 ;
        RECT 85.680 194.065 85.925 194.635 ;
        RECT 86.115 194.235 86.370 194.635 ;
        RECT 86.540 194.405 86.925 194.805 ;
        RECT 86.115 194.065 86.925 194.235 ;
        RECT 87.095 194.065 87.355 194.635 ;
        RECT 87.985 194.080 88.275 194.805 ;
        RECT 88.535 194.255 88.705 194.635 ;
        RECT 88.920 194.425 89.250 194.805 ;
        RECT 88.535 194.085 89.250 194.255 ;
        RECT 83.580 193.895 83.915 194.065 ;
        RECT 84.160 193.895 84.510 194.065 ;
        RECT 85.160 193.895 85.510 194.065 ;
        RECT 85.755 193.895 85.925 194.065 ;
        RECT 86.575 193.895 86.925 194.065 ;
        RECT 81.625 192.425 81.805 193.185 ;
        RECT 81.985 192.255 82.315 193.015 ;
        RECT 82.485 192.425 82.755 193.330 ;
        RECT 82.925 193.190 83.410 193.895 ;
        RECT 83.580 193.565 83.990 193.895 ;
        RECT 83.580 193.020 83.915 193.565 ;
        RECT 84.160 193.395 84.990 193.895 ;
        RECT 82.925 192.850 83.915 193.020 ;
        RECT 84.085 193.215 84.990 193.395 ;
        RECT 85.160 193.565 85.585 193.895 ;
        RECT 82.925 192.425 83.360 192.850 ;
        RECT 83.530 192.255 83.915 192.680 ;
        RECT 84.085 192.425 84.510 193.215 ;
        RECT 85.160 193.045 85.510 193.565 ;
        RECT 85.755 193.395 86.405 193.895 ;
        RECT 84.680 192.850 85.510 193.045 ;
        RECT 85.680 193.215 86.405 193.395 ;
        RECT 86.575 193.565 87.000 193.895 ;
        RECT 84.680 192.425 84.955 192.850 ;
        RECT 85.125 192.255 85.510 192.680 ;
        RECT 85.680 192.425 85.925 193.215 ;
        RECT 86.575 193.045 86.925 193.565 ;
        RECT 87.170 193.395 87.355 194.065 ;
        RECT 88.445 193.535 88.800 193.905 ;
        RECT 89.080 193.895 89.250 194.085 ;
        RECT 89.420 194.060 89.675 194.635 ;
        RECT 89.080 193.565 89.335 193.895 ;
        RECT 86.115 192.850 86.925 193.045 ;
        RECT 86.115 192.425 86.370 192.850 ;
        RECT 86.540 192.255 86.925 192.680 ;
        RECT 87.095 192.425 87.355 193.395 ;
        RECT 87.985 192.255 88.275 193.420 ;
        RECT 89.080 193.355 89.250 193.565 ;
        RECT 88.535 193.185 89.250 193.355 ;
        RECT 89.505 193.330 89.675 194.060 ;
        RECT 89.850 193.965 90.110 194.805 ;
        RECT 91.295 194.255 91.465 194.635 ;
        RECT 91.645 194.425 91.975 194.805 ;
        RECT 91.295 194.085 91.960 194.255 ;
        RECT 92.155 194.130 92.415 194.635 ;
        RECT 91.225 193.535 91.555 193.905 ;
        RECT 91.790 193.830 91.960 194.085 ;
        RECT 91.790 193.500 92.075 193.830 ;
        RECT 88.535 192.425 88.705 193.185 ;
        RECT 88.920 192.255 89.250 193.015 ;
        RECT 89.420 192.425 89.675 193.330 ;
        RECT 89.850 192.255 90.110 193.405 ;
        RECT 91.790 193.355 91.960 193.500 ;
        RECT 91.295 193.185 91.960 193.355 ;
        RECT 92.245 193.330 92.415 194.130 ;
        RECT 92.675 194.255 92.845 194.635 ;
        RECT 93.060 194.425 93.390 194.805 ;
        RECT 92.675 194.085 93.390 194.255 ;
        RECT 92.585 193.535 92.940 193.905 ;
        RECT 93.220 193.895 93.390 194.085 ;
        RECT 93.560 194.060 93.815 194.635 ;
        RECT 93.220 193.565 93.475 193.895 ;
        RECT 93.220 193.355 93.390 193.565 ;
        RECT 91.295 192.425 91.465 193.185 ;
        RECT 91.645 192.255 91.975 193.015 ;
        RECT 92.145 192.425 92.415 193.330 ;
        RECT 92.675 193.185 93.390 193.355 ;
        RECT 93.645 193.330 93.815 194.060 ;
        RECT 93.990 193.965 94.250 194.805 ;
        RECT 94.515 194.255 94.685 194.635 ;
        RECT 94.865 194.425 95.195 194.805 ;
        RECT 94.515 194.085 95.180 194.255 ;
        RECT 95.375 194.130 95.635 194.635 ;
        RECT 94.445 193.535 94.785 193.905 ;
        RECT 95.010 193.830 95.180 194.085 ;
        RECT 95.010 193.500 95.285 193.830 ;
        RECT 92.675 192.425 92.845 193.185 ;
        RECT 93.060 192.255 93.390 193.015 ;
        RECT 93.560 192.425 93.815 193.330 ;
        RECT 93.990 192.255 94.250 193.405 ;
        RECT 95.010 193.355 95.180 193.500 ;
        RECT 94.505 193.185 95.180 193.355 ;
        RECT 95.455 193.330 95.635 194.130 ;
        RECT 94.505 192.425 94.685 193.185 ;
        RECT 94.865 192.255 95.195 193.015 ;
        RECT 95.365 192.425 95.635 193.330 ;
        RECT 95.805 194.130 96.065 194.635 ;
        RECT 96.245 194.425 96.575 194.805 ;
        RECT 96.755 194.255 96.925 194.635 ;
        RECT 95.805 193.330 95.985 194.130 ;
        RECT 96.260 194.085 96.925 194.255 ;
        RECT 97.735 194.255 97.905 194.635 ;
        RECT 98.085 194.425 98.415 194.805 ;
        RECT 97.735 194.085 98.400 194.255 ;
        RECT 98.595 194.130 98.855 194.635 ;
        RECT 96.260 193.830 96.430 194.085 ;
        RECT 96.155 193.500 96.430 193.830 ;
        RECT 96.655 193.535 96.995 193.905 ;
        RECT 97.665 193.535 98.005 193.905 ;
        RECT 98.230 193.830 98.400 194.085 ;
        RECT 96.260 193.355 96.430 193.500 ;
        RECT 98.230 193.500 98.505 193.830 ;
        RECT 98.230 193.355 98.400 193.500 ;
        RECT 95.805 192.425 96.075 193.330 ;
        RECT 96.260 193.185 96.935 193.355 ;
        RECT 96.245 192.255 96.575 193.015 ;
        RECT 96.755 192.425 96.935 193.185 ;
        RECT 97.725 193.185 98.400 193.355 ;
        RECT 98.675 193.330 98.855 194.130 ;
        RECT 99.030 193.965 99.290 194.805 ;
        RECT 99.465 194.060 99.720 194.635 ;
        RECT 99.890 194.425 100.220 194.805 ;
        RECT 100.435 194.255 100.605 194.635 ;
        RECT 99.890 194.085 100.605 194.255 ;
        RECT 97.725 192.425 97.905 193.185 ;
        RECT 98.085 192.255 98.415 193.015 ;
        RECT 98.585 192.425 98.855 193.330 ;
        RECT 99.030 192.255 99.290 193.405 ;
        RECT 99.465 193.330 99.635 194.060 ;
        RECT 99.890 193.895 100.060 194.085 ;
        RECT 100.865 194.080 101.155 194.805 ;
        RECT 102.250 193.965 102.510 194.805 ;
        RECT 102.685 194.060 102.940 194.635 ;
        RECT 103.110 194.425 103.440 194.805 ;
        RECT 103.655 194.255 103.825 194.635 ;
        RECT 103.110 194.085 103.825 194.255 ;
        RECT 104.085 194.130 104.345 194.635 ;
        RECT 104.525 194.425 104.855 194.805 ;
        RECT 105.035 194.255 105.205 194.635 ;
        RECT 99.805 193.565 100.060 193.895 ;
        RECT 99.890 193.355 100.060 193.565 ;
        RECT 100.340 193.535 100.695 193.905 ;
        RECT 99.465 192.425 99.720 193.330 ;
        RECT 99.890 193.185 100.605 193.355 ;
        RECT 99.890 192.255 100.220 193.015 ;
        RECT 100.435 192.425 100.605 193.185 ;
        RECT 100.865 192.255 101.155 193.420 ;
        RECT 102.250 192.255 102.510 193.405 ;
        RECT 102.685 193.330 102.855 194.060 ;
        RECT 103.110 193.895 103.280 194.085 ;
        RECT 103.025 193.565 103.280 193.895 ;
        RECT 103.110 193.355 103.280 193.565 ;
        RECT 103.560 193.535 103.915 193.905 ;
        RECT 102.685 192.425 102.940 193.330 ;
        RECT 103.110 193.185 103.825 193.355 ;
        RECT 103.110 192.255 103.440 193.015 ;
        RECT 103.655 192.425 103.825 193.185 ;
        RECT 104.085 193.330 104.265 194.130 ;
        RECT 104.540 194.085 105.205 194.255 ;
        RECT 104.540 193.830 104.710 194.085 ;
        RECT 105.470 193.965 105.730 194.805 ;
        RECT 105.905 194.060 106.160 194.635 ;
        RECT 106.330 194.425 106.660 194.805 ;
        RECT 106.875 194.255 107.045 194.635 ;
        RECT 106.330 194.085 107.045 194.255 ;
        RECT 107.305 194.130 107.565 194.635 ;
        RECT 107.745 194.425 108.075 194.805 ;
        RECT 108.255 194.255 108.425 194.635 ;
        RECT 104.435 193.500 104.710 193.830 ;
        RECT 104.935 193.535 105.275 193.905 ;
        RECT 104.540 193.355 104.710 193.500 ;
        RECT 104.085 192.425 104.355 193.330 ;
        RECT 104.540 193.185 105.215 193.355 ;
        RECT 104.525 192.255 104.855 193.015 ;
        RECT 105.035 192.425 105.215 193.185 ;
        RECT 105.470 192.255 105.730 193.405 ;
        RECT 105.905 193.330 106.075 194.060 ;
        RECT 106.330 193.895 106.500 194.085 ;
        RECT 106.245 193.565 106.500 193.895 ;
        RECT 106.330 193.355 106.500 193.565 ;
        RECT 106.780 193.535 107.135 193.905 ;
        RECT 105.905 192.425 106.160 193.330 ;
        RECT 106.330 193.185 107.045 193.355 ;
        RECT 106.330 192.255 106.660 193.015 ;
        RECT 106.875 192.425 107.045 193.185 ;
        RECT 107.305 193.330 107.475 194.130 ;
        RECT 107.760 194.085 108.425 194.255 ;
        RECT 107.760 193.830 107.930 194.085 ;
        RECT 109.180 194.065 109.795 194.635 ;
        RECT 109.965 194.295 110.180 194.805 ;
        RECT 110.410 194.295 110.690 194.625 ;
        RECT 110.870 194.295 111.110 194.805 ;
        RECT 107.645 193.500 107.930 193.830 ;
        RECT 108.165 193.535 108.495 193.905 ;
        RECT 107.760 193.355 107.930 193.500 ;
        RECT 107.305 192.425 107.575 193.330 ;
        RECT 107.760 193.185 108.425 193.355 ;
        RECT 107.745 192.255 108.075 193.015 ;
        RECT 108.255 192.425 108.425 193.185 ;
        RECT 109.180 193.045 109.495 194.065 ;
        RECT 109.665 193.395 109.835 193.895 ;
        RECT 110.085 193.565 110.350 194.125 ;
        RECT 110.520 193.395 110.690 194.295 ;
        RECT 111.645 194.175 111.975 194.535 ;
        RECT 112.595 194.345 112.845 194.805 ;
        RECT 113.015 194.345 113.575 194.635 ;
        RECT 110.860 193.565 111.215 194.125 ;
        RECT 111.645 193.985 113.035 194.175 ;
        RECT 112.865 193.895 113.035 193.985 ;
        RECT 111.460 193.565 112.135 193.815 ;
        RECT 112.355 193.565 112.695 193.815 ;
        RECT 112.865 193.565 113.155 193.895 ;
        RECT 109.665 193.225 111.090 193.395 ;
        RECT 109.180 192.425 109.715 193.045 ;
        RECT 109.885 192.255 110.215 193.055 ;
        RECT 110.700 193.050 111.090 193.225 ;
        RECT 111.460 193.205 111.725 193.565 ;
        RECT 112.865 193.315 113.035 193.565 ;
        RECT 112.095 193.145 113.035 193.315 ;
        RECT 111.645 192.255 111.925 192.925 ;
        RECT 112.095 192.595 112.395 193.145 ;
        RECT 113.325 192.975 113.575 194.345 ;
        RECT 113.745 194.080 114.035 194.805 ;
        RECT 115.130 193.965 115.390 194.805 ;
        RECT 115.565 194.060 115.820 194.635 ;
        RECT 115.990 194.425 116.320 194.805 ;
        RECT 116.535 194.255 116.705 194.635 ;
        RECT 115.990 194.085 116.705 194.255 ;
        RECT 117.165 194.175 117.495 194.535 ;
        RECT 118.125 194.345 118.375 194.805 ;
        RECT 118.545 194.345 119.095 194.635 ;
        RECT 112.595 192.255 112.925 192.975 ;
        RECT 113.115 192.425 113.575 192.975 ;
        RECT 113.745 192.255 114.035 193.420 ;
        RECT 115.130 192.255 115.390 193.405 ;
        RECT 115.565 193.330 115.735 194.060 ;
        RECT 115.990 193.895 116.160 194.085 ;
        RECT 117.165 193.985 118.555 194.175 ;
        RECT 115.905 193.565 116.160 193.895 ;
        RECT 115.990 193.355 116.160 193.565 ;
        RECT 116.440 193.535 116.795 193.905 ;
        RECT 118.385 193.895 118.555 193.985 ;
        RECT 116.965 193.565 117.655 193.815 ;
        RECT 117.885 193.565 118.215 193.815 ;
        RECT 118.385 193.565 118.675 193.895 ;
        RECT 115.565 192.425 115.820 193.330 ;
        RECT 115.990 193.185 116.705 193.355 ;
        RECT 115.990 192.255 116.320 193.015 ;
        RECT 116.535 192.425 116.705 193.185 ;
        RECT 116.965 193.125 117.280 193.565 ;
        RECT 118.385 193.315 118.555 193.565 ;
        RECT 117.615 193.145 118.555 193.315 ;
        RECT 117.165 192.255 117.445 192.925 ;
        RECT 117.615 192.595 117.915 193.145 ;
        RECT 118.845 192.975 119.095 194.345 ;
        RECT 119.265 194.005 119.555 194.805 ;
        RECT 119.785 193.985 119.995 194.805 ;
        RECT 120.165 194.005 120.495 194.635 ;
        RECT 120.165 193.405 120.415 194.005 ;
        RECT 120.665 193.985 120.895 194.805 ;
        RECT 121.105 194.130 121.365 194.635 ;
        RECT 121.545 194.425 121.875 194.805 ;
        RECT 122.055 194.255 122.225 194.635 ;
        RECT 120.585 193.565 120.915 193.815 ;
        RECT 118.125 192.255 118.455 192.975 ;
        RECT 118.645 192.425 119.095 192.975 ;
        RECT 119.265 192.255 119.555 193.395 ;
        RECT 119.785 192.255 119.995 193.395 ;
        RECT 120.165 192.425 120.495 193.405 ;
        RECT 120.665 192.255 120.895 193.395 ;
        RECT 121.105 193.330 121.275 194.130 ;
        RECT 121.560 194.085 122.225 194.255 ;
        RECT 122.485 194.130 122.745 194.635 ;
        RECT 122.925 194.425 123.255 194.805 ;
        RECT 123.435 194.255 123.605 194.635 ;
        RECT 121.560 193.830 121.730 194.085 ;
        RECT 121.445 193.500 121.730 193.830 ;
        RECT 121.965 193.535 122.295 193.905 ;
        RECT 121.560 193.355 121.730 193.500 ;
        RECT 121.105 192.425 121.375 193.330 ;
        RECT 121.560 193.185 122.225 193.355 ;
        RECT 121.545 192.255 121.875 193.015 ;
        RECT 122.055 192.425 122.225 193.185 ;
        RECT 122.485 193.330 122.665 194.130 ;
        RECT 122.940 194.085 123.605 194.255 ;
        RECT 123.865 194.175 124.205 194.635 ;
        RECT 124.375 194.345 124.545 194.805 ;
        RECT 125.175 194.370 125.535 194.635 ;
        RECT 125.180 194.365 125.535 194.370 ;
        RECT 125.185 194.355 125.535 194.365 ;
        RECT 125.190 194.350 125.535 194.355 ;
        RECT 125.195 194.340 125.535 194.350 ;
        RECT 125.775 194.345 125.945 194.805 ;
        RECT 125.200 194.335 125.535 194.340 ;
        RECT 125.210 194.325 125.535 194.335 ;
        RECT 125.220 194.315 125.535 194.325 ;
        RECT 124.715 194.175 125.045 194.255 ;
        RECT 122.940 193.830 123.110 194.085 ;
        RECT 123.865 193.985 125.045 194.175 ;
        RECT 125.235 194.175 125.535 194.315 ;
        RECT 125.235 193.985 125.945 194.175 ;
        RECT 122.835 193.500 123.110 193.830 ;
        RECT 123.335 193.535 123.675 193.905 ;
        RECT 123.865 193.615 124.195 193.815 ;
        RECT 124.505 193.795 124.835 193.815 ;
        RECT 124.385 193.615 124.835 193.795 ;
        RECT 122.940 193.355 123.110 193.500 ;
        RECT 122.485 192.425 122.755 193.330 ;
        RECT 122.940 193.185 123.615 193.355 ;
        RECT 123.865 193.275 124.095 193.615 ;
        RECT 122.925 192.255 123.255 193.015 ;
        RECT 123.435 192.425 123.615 193.185 ;
        RECT 123.875 192.255 124.205 192.975 ;
        RECT 124.385 192.500 124.600 193.615 ;
        RECT 125.005 193.585 125.475 193.815 ;
        RECT 125.660 193.415 125.945 193.985 ;
        RECT 126.115 193.860 126.455 194.635 ;
        RECT 126.625 194.080 126.915 194.805 ;
        RECT 127.175 194.255 127.345 194.635 ;
        RECT 127.560 194.425 127.890 194.805 ;
        RECT 127.175 194.085 127.890 194.255 ;
        RECT 124.795 193.200 125.945 193.415 ;
        RECT 124.795 192.425 125.125 193.200 ;
        RECT 125.295 192.255 126.005 193.030 ;
        RECT 126.175 192.425 126.455 193.860 ;
        RECT 127.085 193.535 127.440 193.905 ;
        RECT 127.720 193.895 127.890 194.085 ;
        RECT 128.060 194.060 128.315 194.635 ;
        RECT 127.720 193.565 127.975 193.895 ;
        RECT 126.625 192.255 126.915 193.420 ;
        RECT 127.720 193.355 127.890 193.565 ;
        RECT 127.175 193.185 127.890 193.355 ;
        RECT 128.145 193.330 128.315 194.060 ;
        RECT 128.490 193.965 128.750 194.805 ;
        RECT 129.385 194.065 129.875 194.635 ;
        RECT 130.045 194.235 130.275 194.635 ;
        RECT 130.445 194.405 130.865 194.805 ;
        RECT 131.035 194.235 131.205 194.635 ;
        RECT 130.045 194.065 131.205 194.235 ;
        RECT 131.375 194.065 131.825 194.805 ;
        RECT 131.995 194.065 132.435 194.625 ;
        RECT 132.605 194.315 132.865 194.805 ;
        RECT 133.115 194.245 133.380 194.505 ;
        RECT 133.555 194.405 133.885 194.805 ;
        RECT 133.025 194.235 133.380 194.245 ;
        RECT 134.055 194.235 134.225 194.505 ;
        RECT 134.395 194.405 134.725 194.805 ;
        RECT 127.175 192.425 127.345 193.185 ;
        RECT 127.560 192.255 127.890 193.015 ;
        RECT 128.060 192.425 128.315 193.330 ;
        RECT 128.490 192.255 128.750 193.405 ;
        RECT 129.385 193.395 129.555 194.065 ;
        RECT 129.725 193.565 130.130 193.895 ;
        RECT 129.385 193.225 130.155 193.395 ;
        RECT 129.395 192.255 129.725 193.055 ;
        RECT 129.905 192.595 130.155 193.225 ;
        RECT 130.345 192.765 130.595 193.895 ;
        RECT 130.795 193.565 131.040 193.895 ;
        RECT 131.225 193.615 131.615 193.895 ;
        RECT 130.795 192.765 130.995 193.565 ;
        RECT 131.785 193.445 131.955 193.895 ;
        RECT 131.165 193.275 131.955 193.445 ;
        RECT 131.165 192.595 131.335 193.275 ;
        RECT 129.905 192.425 131.335 192.595 ;
        RECT 131.505 192.255 131.820 193.105 ;
        RECT 132.125 193.055 132.435 194.065 ;
        RECT 132.605 193.565 132.855 194.145 ;
        RECT 133.025 194.065 134.225 194.235 ;
        RECT 133.025 193.395 133.195 194.065 ;
        RECT 131.995 192.425 132.435 193.055 ;
        RECT 132.610 193.225 133.195 193.395 ;
        RECT 133.365 193.475 133.595 193.895 ;
        RECT 133.765 193.645 134.215 193.815 ;
        RECT 133.365 193.275 133.805 193.475 ;
        RECT 132.610 192.440 132.945 193.225 ;
        RECT 133.550 192.440 133.805 193.275 ;
        RECT 133.975 192.440 134.215 193.645 ;
        RECT 134.475 193.225 134.735 194.235 ;
        RECT 134.905 194.055 136.115 194.805 ;
        RECT 134.905 193.345 135.425 193.885 ;
        RECT 135.595 193.515 136.115 194.055 ;
        RECT 134.475 192.255 134.735 193.055 ;
        RECT 134.905 192.255 136.115 193.345 ;
        RECT 23.500 192.085 136.200 192.255 ;
        RECT 23.585 190.995 24.795 192.085 ;
        RECT 23.585 190.285 24.105 190.825 ;
        RECT 24.275 190.455 24.795 190.995 ;
        RECT 24.970 190.935 25.230 192.085 ;
        RECT 25.405 191.010 25.660 191.915 ;
        RECT 25.830 191.325 26.160 192.085 ;
        RECT 26.375 191.155 26.545 191.915 ;
        RECT 23.585 189.535 24.795 190.285 ;
        RECT 24.970 189.535 25.230 190.375 ;
        RECT 25.405 190.280 25.575 191.010 ;
        RECT 25.830 190.985 26.545 191.155 ;
        RECT 27.725 191.010 27.995 191.915 ;
        RECT 28.165 191.325 28.495 192.085 ;
        RECT 28.675 191.155 28.845 191.915 ;
        RECT 29.105 191.650 34.450 192.085 ;
        RECT 25.830 190.775 26.000 190.985 ;
        RECT 25.745 190.445 26.000 190.775 ;
        RECT 25.405 189.705 25.660 190.280 ;
        RECT 25.830 190.255 26.000 190.445 ;
        RECT 26.280 190.435 26.635 190.805 ;
        RECT 25.830 190.085 26.545 190.255 ;
        RECT 25.830 189.535 26.160 189.915 ;
        RECT 26.375 189.705 26.545 190.085 ;
        RECT 27.725 190.210 27.895 191.010 ;
        RECT 28.180 190.985 28.845 191.155 ;
        RECT 28.180 190.840 28.350 190.985 ;
        RECT 28.065 190.510 28.350 190.840 ;
        RECT 28.180 190.255 28.350 190.510 ;
        RECT 28.585 190.435 28.915 190.805 ;
        RECT 27.725 189.705 27.985 190.210 ;
        RECT 28.180 190.085 28.845 190.255 ;
        RECT 28.165 189.535 28.495 189.915 ;
        RECT 28.675 189.705 28.845 190.085 ;
        RECT 30.690 190.080 31.030 190.910 ;
        RECT 32.510 190.400 32.860 191.650 ;
        RECT 34.625 190.995 36.295 192.085 ;
        RECT 34.625 190.305 35.375 190.825 ;
        RECT 35.545 190.475 36.295 190.995 ;
        RECT 36.465 190.920 36.755 192.085 ;
        RECT 36.925 190.995 38.135 192.085 ;
        RECT 29.105 189.535 34.450 190.080 ;
        RECT 34.625 189.535 36.295 190.305 ;
        RECT 36.925 190.285 37.445 190.825 ;
        RECT 37.615 190.455 38.135 190.995 ;
        RECT 38.310 190.945 38.645 191.915 ;
        RECT 38.815 190.945 38.985 192.085 ;
        RECT 39.155 191.745 41.185 191.915 ;
        RECT 36.465 189.535 36.755 190.260 ;
        RECT 36.925 189.535 38.135 190.285 ;
        RECT 38.310 190.275 38.480 190.945 ;
        RECT 39.155 190.775 39.325 191.745 ;
        RECT 38.650 190.445 38.905 190.775 ;
        RECT 39.130 190.445 39.325 190.775 ;
        RECT 39.495 191.405 40.620 191.575 ;
        RECT 38.735 190.275 38.905 190.445 ;
        RECT 39.495 190.275 39.665 191.405 ;
        RECT 38.310 189.705 38.565 190.275 ;
        RECT 38.735 190.105 39.665 190.275 ;
        RECT 39.835 191.065 40.845 191.235 ;
        RECT 39.835 190.265 40.005 191.065 ;
        RECT 40.210 190.385 40.485 190.865 ;
        RECT 40.205 190.215 40.485 190.385 ;
        RECT 39.490 190.070 39.665 190.105 ;
        RECT 38.735 189.535 39.065 189.935 ;
        RECT 39.490 189.705 40.020 190.070 ;
        RECT 40.210 189.705 40.485 190.215 ;
        RECT 40.655 189.705 40.845 191.065 ;
        RECT 41.015 191.080 41.185 191.745 ;
        RECT 41.355 191.325 41.525 192.085 ;
        RECT 41.760 191.325 42.275 191.735 ;
        RECT 41.015 190.890 41.765 191.080 ;
        RECT 41.935 190.515 42.275 191.325 ;
        RECT 41.045 190.345 42.275 190.515 ;
        RECT 42.480 191.295 43.015 191.915 ;
        RECT 41.025 189.535 41.535 190.070 ;
        RECT 41.755 189.740 42.000 190.345 ;
        RECT 42.480 190.275 42.795 191.295 ;
        RECT 43.185 191.285 43.515 192.085 ;
        RECT 44.000 191.115 44.390 191.290 ;
        RECT 42.965 190.945 44.390 191.115 ;
        RECT 44.745 190.995 46.415 192.085 ;
        RECT 42.965 190.445 43.135 190.945 ;
        RECT 42.480 189.705 43.095 190.275 ;
        RECT 43.385 190.215 43.650 190.775 ;
        RECT 43.820 190.045 43.990 190.945 ;
        RECT 44.160 190.215 44.515 190.775 ;
        RECT 44.745 190.305 45.495 190.825 ;
        RECT 45.665 190.475 46.415 190.995 ;
        RECT 47.055 191.475 47.385 191.905 ;
        RECT 47.565 191.645 47.760 192.085 ;
        RECT 47.930 191.475 48.260 191.905 ;
        RECT 47.055 191.305 48.260 191.475 ;
        RECT 47.055 190.975 47.950 191.305 ;
        RECT 48.430 191.135 48.705 191.905 ;
        RECT 48.120 190.945 48.705 191.135 ;
        RECT 48.895 191.135 49.170 191.905 ;
        RECT 49.340 191.475 49.670 191.905 ;
        RECT 49.840 191.645 50.035 192.085 ;
        RECT 50.215 191.475 50.545 191.905 ;
        RECT 49.340 191.305 50.545 191.475 ;
        RECT 48.895 190.945 49.480 191.135 ;
        RECT 49.650 190.975 50.545 191.305 ;
        RECT 47.060 190.445 47.355 190.775 ;
        RECT 47.535 190.445 47.950 190.775 ;
        RECT 43.265 189.535 43.480 190.045 ;
        RECT 43.710 189.715 43.990 190.045 ;
        RECT 44.170 189.535 44.410 190.045 ;
        RECT 44.745 189.535 46.415 190.305 ;
        RECT 47.055 189.535 47.355 190.265 ;
        RECT 47.535 189.825 47.765 190.445 ;
        RECT 48.120 190.275 48.295 190.945 ;
        RECT 47.965 190.095 48.295 190.275 ;
        RECT 48.465 190.125 48.705 190.775 ;
        RECT 48.895 190.125 49.135 190.775 ;
        RECT 49.305 190.275 49.480 190.945 ;
        RECT 49.650 190.445 50.065 190.775 ;
        RECT 50.245 190.445 50.540 190.775 ;
        RECT 49.305 190.095 49.635 190.275 ;
        RECT 47.965 189.715 48.190 190.095 ;
        RECT 48.360 189.535 48.690 189.925 ;
        RECT 48.910 189.535 49.240 189.925 ;
        RECT 49.410 189.715 49.635 190.095 ;
        RECT 49.835 189.825 50.065 190.445 ;
        RECT 50.245 189.535 50.545 190.265 ;
        RECT 50.725 189.815 51.005 191.915 ;
        RECT 51.195 191.325 51.980 192.085 ;
        RECT 52.375 191.255 52.760 191.915 ;
        RECT 52.375 191.155 52.785 191.255 ;
        RECT 51.175 190.945 52.785 191.155 ;
        RECT 53.085 191.065 53.285 191.855 ;
        RECT 51.175 190.345 51.450 190.945 ;
        RECT 52.955 190.895 53.285 191.065 ;
        RECT 53.455 190.905 53.775 192.085 ;
        RECT 53.950 190.945 54.285 191.915 ;
        RECT 54.455 190.945 54.625 192.085 ;
        RECT 54.795 191.745 56.825 191.915 ;
        RECT 52.955 190.775 53.135 190.895 ;
        RECT 51.620 190.525 51.975 190.775 ;
        RECT 52.170 190.725 52.635 190.775 ;
        RECT 52.165 190.555 52.635 190.725 ;
        RECT 52.170 190.525 52.635 190.555 ;
        RECT 52.805 190.525 53.135 190.775 ;
        RECT 53.310 190.525 53.775 190.725 ;
        RECT 51.175 190.165 52.425 190.345 ;
        RECT 52.060 190.095 52.425 190.165 ;
        RECT 52.595 190.145 53.775 190.315 ;
        RECT 51.235 189.535 51.405 189.995 ;
        RECT 52.595 189.925 52.925 190.145 ;
        RECT 51.675 189.745 52.925 189.925 ;
        RECT 53.095 189.535 53.265 189.975 ;
        RECT 53.435 189.730 53.775 190.145 ;
        RECT 53.950 190.275 54.120 190.945 ;
        RECT 54.795 190.775 54.965 191.745 ;
        RECT 54.290 190.445 54.545 190.775 ;
        RECT 54.770 190.445 54.965 190.775 ;
        RECT 55.135 191.405 56.260 191.575 ;
        RECT 54.375 190.275 54.545 190.445 ;
        RECT 55.135 190.275 55.305 191.405 ;
        RECT 53.950 189.705 54.205 190.275 ;
        RECT 54.375 190.105 55.305 190.275 ;
        RECT 55.475 191.065 56.485 191.235 ;
        RECT 55.475 190.265 55.645 191.065 ;
        RECT 55.130 190.070 55.305 190.105 ;
        RECT 54.375 189.535 54.705 189.935 ;
        RECT 55.130 189.705 55.660 190.070 ;
        RECT 55.850 190.045 56.125 190.865 ;
        RECT 55.845 189.875 56.125 190.045 ;
        RECT 55.850 189.705 56.125 189.875 ;
        RECT 56.295 189.705 56.485 191.065 ;
        RECT 56.655 191.080 56.825 191.745 ;
        RECT 56.995 191.325 57.165 192.085 ;
        RECT 57.400 191.325 57.915 191.735 ;
        RECT 58.090 191.660 58.425 192.085 ;
        RECT 58.595 191.480 58.780 191.885 ;
        RECT 56.655 190.890 57.405 191.080 ;
        RECT 57.575 190.515 57.915 191.325 ;
        RECT 56.685 190.345 57.915 190.515 ;
        RECT 58.115 191.305 58.780 191.480 ;
        RECT 58.985 191.305 59.315 192.085 ;
        RECT 56.665 189.535 57.175 190.070 ;
        RECT 57.395 189.740 57.640 190.345 ;
        RECT 58.115 190.275 58.455 191.305 ;
        RECT 59.485 191.115 59.755 191.885 ;
        RECT 58.625 190.945 59.755 191.115 ;
        RECT 59.925 190.995 61.595 192.085 ;
        RECT 58.625 190.445 58.875 190.945 ;
        RECT 58.115 190.105 58.800 190.275 ;
        RECT 59.055 190.195 59.415 190.775 ;
        RECT 58.090 189.535 58.425 189.935 ;
        RECT 58.595 189.705 58.800 190.105 ;
        RECT 59.585 190.035 59.755 190.945 ;
        RECT 59.010 189.535 59.285 190.015 ;
        RECT 59.495 189.705 59.755 190.035 ;
        RECT 59.925 190.305 60.675 190.825 ;
        RECT 60.845 190.475 61.595 190.995 ;
        RECT 62.225 190.920 62.515 192.085 ;
        RECT 62.685 190.995 63.895 192.085 ;
        RECT 59.925 189.535 61.595 190.305 ;
        RECT 62.685 190.285 63.205 190.825 ;
        RECT 63.375 190.455 63.895 190.995 ;
        RECT 64.070 190.935 64.330 192.085 ;
        RECT 64.505 191.010 64.760 191.915 ;
        RECT 64.930 191.325 65.260 192.085 ;
        RECT 65.475 191.155 65.645 191.915 ;
        RECT 62.225 189.535 62.515 190.260 ;
        RECT 62.685 189.535 63.895 190.285 ;
        RECT 64.070 189.535 64.330 190.375 ;
        RECT 64.505 190.280 64.675 191.010 ;
        RECT 64.930 190.985 65.645 191.155 ;
        RECT 65.915 191.475 66.245 191.905 ;
        RECT 66.425 191.645 66.620 192.085 ;
        RECT 66.790 191.475 67.120 191.905 ;
        RECT 65.915 191.305 67.120 191.475 ;
        RECT 64.930 190.775 65.100 190.985 ;
        RECT 65.915 190.975 66.810 191.305 ;
        RECT 67.290 191.135 67.565 191.905 ;
        RECT 66.980 190.945 67.565 191.135 ;
        RECT 67.745 191.010 68.015 191.915 ;
        RECT 68.185 191.325 68.515 192.085 ;
        RECT 68.695 191.155 68.865 191.915 ;
        RECT 64.845 190.445 65.100 190.775 ;
        RECT 64.505 189.705 64.760 190.280 ;
        RECT 64.930 190.255 65.100 190.445 ;
        RECT 65.380 190.435 65.735 190.805 ;
        RECT 65.920 190.445 66.215 190.775 ;
        RECT 66.395 190.445 66.810 190.775 ;
        RECT 64.930 190.085 65.645 190.255 ;
        RECT 64.930 189.535 65.260 189.915 ;
        RECT 65.475 189.705 65.645 190.085 ;
        RECT 65.915 189.535 66.215 190.265 ;
        RECT 66.395 189.825 66.625 190.445 ;
        RECT 66.980 190.275 67.155 190.945 ;
        RECT 66.825 190.095 67.155 190.275 ;
        RECT 67.325 190.125 67.565 190.775 ;
        RECT 67.745 190.210 67.915 191.010 ;
        RECT 68.200 190.985 68.865 191.155 ;
        RECT 69.140 191.100 69.465 192.085 ;
        RECT 70.035 191.455 70.295 191.915 ;
        RECT 70.465 191.635 71.315 192.085 ;
        RECT 69.650 191.405 69.855 191.435 ;
        RECT 69.645 191.235 69.855 191.405 ;
        RECT 70.035 191.235 71.155 191.455 ;
        RECT 68.200 190.840 68.370 190.985 ;
        RECT 68.085 190.510 68.370 190.840 ;
        RECT 68.200 190.255 68.370 190.510 ;
        RECT 68.605 190.435 68.935 190.805 ;
        RECT 69.135 190.445 69.395 190.900 ;
        RECT 69.650 190.850 69.855 191.235 ;
        RECT 69.650 190.475 70.235 190.850 ;
        RECT 70.405 190.460 70.815 191.065 ;
        RECT 70.985 190.780 71.155 191.235 ;
        RECT 70.985 190.290 71.315 190.780 ;
        RECT 66.825 189.715 67.050 190.095 ;
        RECT 67.220 189.535 67.550 189.925 ;
        RECT 67.745 189.705 68.005 190.210 ;
        RECT 68.200 190.085 68.865 190.255 ;
        RECT 68.185 189.535 68.515 189.915 ;
        RECT 68.695 189.705 68.865 190.085 ;
        RECT 69.140 190.085 70.295 190.275 ;
        RECT 69.140 189.945 69.415 190.085 ;
        RECT 70.085 189.915 70.295 190.085 ;
        RECT 70.465 190.085 71.315 190.290 ;
        RECT 69.585 189.535 69.915 189.915 ;
        RECT 70.465 189.705 70.795 190.085 ;
        RECT 70.985 189.535 71.315 189.915 ;
        RECT 71.485 189.705 71.730 191.915 ;
        RECT 71.915 191.085 72.170 192.085 ;
        RECT 72.345 190.995 73.555 192.085 ;
        RECT 71.915 189.535 72.155 190.335 ;
        RECT 72.345 190.285 72.865 190.825 ;
        RECT 73.035 190.455 73.555 190.995 ;
        RECT 73.725 191.245 73.985 191.915 ;
        RECT 74.155 191.685 74.485 192.085 ;
        RECT 75.355 191.685 75.755 192.085 ;
        RECT 76.045 191.505 76.375 191.740 ;
        RECT 74.295 191.335 76.375 191.505 ;
        RECT 72.345 189.535 73.555 190.285 ;
        RECT 73.725 190.275 73.900 191.245 ;
        RECT 74.295 191.065 74.465 191.335 ;
        RECT 74.070 190.895 74.465 191.065 ;
        RECT 74.635 190.945 75.650 191.165 ;
        RECT 74.070 190.445 74.240 190.895 ;
        RECT 75.375 190.805 75.650 190.945 ;
        RECT 75.820 190.945 76.375 191.335 ;
        RECT 74.410 190.525 74.860 190.725 ;
        RECT 75.030 190.355 75.205 190.550 ;
        RECT 73.725 189.705 74.065 190.275 ;
        RECT 74.260 189.535 74.430 190.200 ;
        RECT 74.710 190.185 75.205 190.355 ;
        RECT 74.710 190.045 74.930 190.185 ;
        RECT 74.705 189.875 74.930 190.045 ;
        RECT 75.375 190.015 75.545 190.805 ;
        RECT 75.820 190.695 75.990 190.945 ;
        RECT 76.545 190.775 76.720 191.875 ;
        RECT 76.890 191.265 77.235 192.085 ;
        RECT 77.440 191.295 77.975 191.915 ;
        RECT 75.795 190.525 75.990 190.695 ;
        RECT 76.160 190.525 76.720 190.775 ;
        RECT 76.890 190.525 77.235 191.095 ;
        RECT 75.795 190.140 75.965 190.525 ;
        RECT 74.710 189.830 74.930 189.875 ;
        RECT 75.100 189.845 75.545 190.015 ;
        RECT 75.715 189.770 75.965 190.140 ;
        RECT 76.135 190.175 77.235 190.355 ;
        RECT 76.135 189.770 76.385 190.175 ;
        RECT 76.555 189.535 76.725 190.005 ;
        RECT 76.895 189.770 77.235 190.175 ;
        RECT 77.440 190.275 77.755 191.295 ;
        RECT 78.145 191.285 78.475 192.085 ;
        RECT 78.960 191.115 79.350 191.290 ;
        RECT 77.925 190.945 79.350 191.115 ;
        RECT 79.705 190.995 82.295 192.085 ;
        RECT 82.570 191.285 82.825 192.085 ;
        RECT 82.995 191.115 83.325 191.915 ;
        RECT 83.495 191.285 83.665 192.085 ;
        RECT 83.835 191.115 84.165 191.915 ;
        RECT 77.925 190.445 78.095 190.945 ;
        RECT 77.440 189.705 78.055 190.275 ;
        RECT 78.345 190.215 78.610 190.775 ;
        RECT 78.780 190.045 78.950 190.945 ;
        RECT 79.120 190.215 79.475 190.775 ;
        RECT 79.705 190.305 80.915 190.825 ;
        RECT 81.085 190.475 82.295 190.995 ;
        RECT 82.465 190.945 84.165 191.115 ;
        RECT 84.335 190.945 84.595 192.085 ;
        RECT 85.265 190.945 85.495 192.085 ;
        RECT 82.465 190.355 82.745 190.945 ;
        RECT 85.665 190.935 85.995 191.915 ;
        RECT 86.165 190.945 86.375 192.085 ;
        RECT 86.695 191.155 86.865 191.915 ;
        RECT 87.045 191.325 87.375 192.085 ;
        RECT 86.695 190.985 87.360 191.155 ;
        RECT 87.545 191.010 87.815 191.915 ;
        RECT 82.915 190.525 83.665 190.775 ;
        RECT 83.835 190.525 84.595 190.775 ;
        RECT 85.245 190.525 85.575 190.775 ;
        RECT 78.225 189.535 78.440 190.045 ;
        RECT 78.670 189.715 78.950 190.045 ;
        RECT 79.130 189.535 79.370 190.045 ;
        RECT 79.705 189.535 82.295 190.305 ;
        RECT 82.465 190.105 83.325 190.355 ;
        RECT 83.495 190.165 84.595 190.335 ;
        RECT 82.575 189.915 82.905 189.935 ;
        RECT 83.495 189.915 83.745 190.165 ;
        RECT 82.575 189.705 83.745 189.915 ;
        RECT 83.915 189.535 84.085 189.995 ;
        RECT 84.255 189.705 84.595 190.165 ;
        RECT 85.265 189.535 85.495 190.355 ;
        RECT 85.745 190.335 85.995 190.935 ;
        RECT 87.190 190.840 87.360 190.985 ;
        RECT 86.625 190.435 86.955 190.805 ;
        RECT 87.190 190.510 87.475 190.840 ;
        RECT 85.665 189.705 85.995 190.335 ;
        RECT 86.165 189.535 86.375 190.355 ;
        RECT 87.190 190.255 87.360 190.510 ;
        RECT 86.695 190.085 87.360 190.255 ;
        RECT 87.645 190.210 87.815 191.010 ;
        RECT 87.985 190.920 88.275 192.085 ;
        RECT 89.565 191.415 89.845 192.085 ;
        RECT 90.015 191.195 90.315 191.745 ;
        RECT 90.515 191.365 90.845 192.085 ;
        RECT 91.035 191.365 91.495 191.915 ;
        RECT 89.380 190.775 89.645 191.135 ;
        RECT 90.015 191.025 90.955 191.195 ;
        RECT 90.785 190.775 90.955 191.025 ;
        RECT 89.380 190.525 90.055 190.775 ;
        RECT 90.275 190.525 90.615 190.775 ;
        RECT 90.785 190.445 91.075 190.775 ;
        RECT 90.785 190.355 90.955 190.445 ;
        RECT 86.695 189.705 86.865 190.085 ;
        RECT 87.045 189.535 87.375 189.915 ;
        RECT 87.555 189.705 87.815 190.210 ;
        RECT 87.985 189.535 88.275 190.260 ;
        RECT 89.565 190.165 90.955 190.355 ;
        RECT 89.565 189.805 89.895 190.165 ;
        RECT 91.245 189.995 91.495 191.365 ;
        RECT 90.515 189.535 90.765 189.995 ;
        RECT 90.935 189.705 91.495 189.995 ;
        RECT 91.700 191.295 92.235 191.915 ;
        RECT 91.700 190.275 92.015 191.295 ;
        RECT 92.405 191.285 92.735 192.085 ;
        RECT 94.625 191.415 94.905 192.085 ;
        RECT 93.220 191.115 93.610 191.290 ;
        RECT 95.075 191.195 95.375 191.745 ;
        RECT 95.575 191.365 95.905 192.085 ;
        RECT 96.095 191.365 96.555 191.915 ;
        RECT 92.185 190.945 93.610 191.115 ;
        RECT 92.185 190.445 92.355 190.945 ;
        RECT 91.700 189.705 92.315 190.275 ;
        RECT 92.605 190.215 92.870 190.775 ;
        RECT 93.040 190.045 93.210 190.945 ;
        RECT 94.440 190.775 94.705 191.135 ;
        RECT 95.075 191.025 96.015 191.195 ;
        RECT 95.845 190.775 96.015 191.025 ;
        RECT 93.380 190.215 93.735 190.775 ;
        RECT 94.440 190.525 95.115 190.775 ;
        RECT 95.335 190.525 95.675 190.775 ;
        RECT 95.845 190.445 96.135 190.775 ;
        RECT 95.845 190.355 96.015 190.445 ;
        RECT 94.625 190.165 96.015 190.355 ;
        RECT 92.485 189.535 92.700 190.045 ;
        RECT 92.930 189.715 93.210 190.045 ;
        RECT 93.390 189.535 93.630 190.045 ;
        RECT 94.625 189.805 94.955 190.165 ;
        RECT 96.305 189.995 96.555 191.365 ;
        RECT 96.765 190.945 96.995 192.085 ;
        RECT 97.165 190.935 97.495 191.915 ;
        RECT 97.665 190.945 97.875 192.085 ;
        RECT 98.115 190.945 98.445 192.085 ;
        RECT 98.975 191.115 99.305 191.900 ;
        RECT 98.625 190.945 99.305 191.115 ;
        RECT 99.575 191.155 99.745 191.915 ;
        RECT 99.925 191.325 100.255 192.085 ;
        RECT 99.575 190.985 100.240 191.155 ;
        RECT 100.425 191.010 100.695 191.915 ;
        RECT 96.745 190.525 97.075 190.775 ;
        RECT 95.575 189.535 95.825 189.995 ;
        RECT 95.995 189.705 96.555 189.995 ;
        RECT 96.765 189.535 96.995 190.355 ;
        RECT 97.245 190.335 97.495 190.935 ;
        RECT 98.105 190.525 98.455 190.775 ;
        RECT 97.165 189.705 97.495 190.335 ;
        RECT 97.665 189.535 97.875 190.355 ;
        RECT 98.625 190.345 98.795 190.945 ;
        RECT 100.070 190.840 100.240 190.985 ;
        RECT 98.965 190.525 99.315 190.775 ;
        RECT 99.505 190.435 99.835 190.805 ;
        RECT 100.070 190.510 100.355 190.840 ;
        RECT 98.115 189.535 98.385 190.345 ;
        RECT 98.555 189.705 98.885 190.345 ;
        RECT 99.055 189.535 99.295 190.345 ;
        RECT 100.070 190.255 100.240 190.510 ;
        RECT 99.575 190.085 100.240 190.255 ;
        RECT 100.525 190.210 100.695 191.010 ;
        RECT 102.175 190.935 102.505 192.085 ;
        RECT 102.675 191.065 102.845 191.915 ;
        RECT 103.015 191.285 103.345 192.085 ;
        RECT 103.515 191.065 103.685 191.915 ;
        RECT 103.855 191.285 104.185 192.085 ;
        RECT 104.355 191.065 104.525 191.915 ;
        RECT 104.695 191.285 105.025 192.085 ;
        RECT 105.195 191.065 105.365 191.915 ;
        RECT 105.615 191.285 105.785 192.085 ;
        RECT 105.955 191.065 106.285 191.915 ;
        RECT 106.455 191.285 106.625 192.085 ;
        RECT 106.795 191.065 107.125 191.915 ;
        RECT 102.675 190.895 105.365 191.065 ;
        RECT 105.625 190.895 107.125 191.065 ;
        RECT 107.305 190.945 107.565 192.085 ;
        RECT 107.735 191.115 108.065 191.915 ;
        RECT 108.235 191.285 108.405 192.085 ;
        RECT 108.575 191.115 108.905 191.915 ;
        RECT 109.075 191.285 109.330 192.085 ;
        RECT 109.605 191.365 110.065 191.915 ;
        RECT 110.255 191.365 110.585 192.085 ;
        RECT 107.735 190.945 109.435 191.115 ;
        RECT 102.675 190.725 102.930 190.895 ;
        RECT 102.675 190.555 102.935 190.725 ;
        RECT 105.625 190.695 105.800 190.895 ;
        RECT 102.675 190.355 102.930 190.555 ;
        RECT 103.175 190.525 105.800 190.695 ;
        RECT 105.980 190.525 107.080 190.725 ;
        RECT 107.305 190.525 108.065 190.775 ;
        RECT 108.235 190.525 108.985 190.775 ;
        RECT 105.625 190.355 105.800 190.525 ;
        RECT 109.155 190.355 109.435 190.945 ;
        RECT 99.575 189.705 99.745 190.085 ;
        RECT 99.925 189.535 100.255 189.915 ;
        RECT 100.435 189.705 100.695 190.210 ;
        RECT 102.175 189.535 102.505 190.335 ;
        RECT 102.675 190.185 105.365 190.355 ;
        RECT 105.625 190.185 107.045 190.355 ;
        RECT 102.675 189.705 102.845 190.185 ;
        RECT 103.015 189.535 103.345 190.015 ;
        RECT 103.515 189.705 103.685 190.185 ;
        RECT 103.855 189.535 104.185 190.015 ;
        RECT 104.355 189.705 104.525 190.185 ;
        RECT 104.695 189.535 105.025 190.015 ;
        RECT 105.195 189.705 105.365 190.185 ;
        RECT 105.535 189.535 105.865 190.015 ;
        RECT 106.035 189.710 106.205 190.185 ;
        RECT 106.375 189.535 106.705 190.015 ;
        RECT 106.875 189.705 107.045 190.185 ;
        RECT 107.305 190.165 108.405 190.335 ;
        RECT 107.305 189.705 107.645 190.165 ;
        RECT 107.815 189.535 107.985 189.995 ;
        RECT 108.155 189.915 108.405 190.165 ;
        RECT 108.575 190.105 109.435 190.355 ;
        RECT 109.605 189.995 109.855 191.365 ;
        RECT 110.785 191.195 111.085 191.745 ;
        RECT 111.255 191.415 111.535 192.085 ;
        RECT 110.145 191.025 111.085 191.195 ;
        RECT 110.145 190.775 110.315 191.025 ;
        RECT 111.455 190.775 111.720 191.135 ;
        RECT 110.025 190.445 110.315 190.775 ;
        RECT 110.485 190.525 110.825 190.775 ;
        RECT 111.045 190.525 111.720 190.775 ;
        RECT 111.905 191.010 112.175 191.915 ;
        RECT 112.345 191.325 112.675 192.085 ;
        RECT 112.855 191.155 113.025 191.915 ;
        RECT 110.145 190.355 110.315 190.445 ;
        RECT 110.145 190.165 111.535 190.355 ;
        RECT 108.995 189.915 109.325 189.935 ;
        RECT 108.155 189.705 109.325 189.915 ;
        RECT 109.605 189.705 110.165 189.995 ;
        RECT 110.335 189.535 110.585 189.995 ;
        RECT 111.205 189.805 111.535 190.165 ;
        RECT 111.905 190.210 112.075 191.010 ;
        RECT 112.360 190.985 113.025 191.155 ;
        RECT 112.360 190.840 112.530 190.985 ;
        RECT 113.745 190.920 114.035 192.085 ;
        RECT 114.205 190.945 114.495 192.085 ;
        RECT 114.665 191.365 115.115 191.915 ;
        RECT 115.305 191.365 115.635 192.085 ;
        RECT 112.245 190.510 112.530 190.840 ;
        RECT 112.360 190.255 112.530 190.510 ;
        RECT 112.765 190.435 113.095 190.805 ;
        RECT 111.905 189.705 112.165 190.210 ;
        RECT 112.360 190.085 113.025 190.255 ;
        RECT 112.345 189.535 112.675 189.915 ;
        RECT 112.855 189.705 113.025 190.085 ;
        RECT 113.745 189.535 114.035 190.260 ;
        RECT 114.205 189.535 114.495 190.335 ;
        RECT 114.665 189.995 114.915 191.365 ;
        RECT 115.845 191.195 116.145 191.745 ;
        RECT 116.315 191.415 116.595 192.085 ;
        RECT 117.895 191.275 118.190 192.085 ;
        RECT 115.205 191.025 116.145 191.195 ;
        RECT 115.205 190.775 115.375 191.025 ;
        RECT 116.480 190.775 116.795 191.215 ;
        RECT 118.370 190.775 118.615 191.915 ;
        RECT 118.790 191.275 119.050 192.085 ;
        RECT 119.650 192.080 125.925 192.085 ;
        RECT 119.230 190.775 119.480 191.910 ;
        RECT 119.650 191.285 119.910 192.080 ;
        RECT 120.080 191.185 120.340 191.910 ;
        RECT 120.510 191.355 120.770 192.080 ;
        RECT 120.940 191.185 121.200 191.910 ;
        RECT 121.370 191.355 121.630 192.080 ;
        RECT 121.800 191.185 122.060 191.910 ;
        RECT 122.230 191.355 122.490 192.080 ;
        RECT 122.660 191.185 122.920 191.910 ;
        RECT 123.090 191.355 123.335 192.080 ;
        RECT 123.505 191.185 123.765 191.910 ;
        RECT 123.950 191.355 124.195 192.080 ;
        RECT 124.365 191.185 124.625 191.910 ;
        RECT 124.810 191.355 125.055 192.080 ;
        RECT 125.225 191.185 125.485 191.910 ;
        RECT 125.670 191.355 125.925 192.080 ;
        RECT 120.080 191.170 125.485 191.185 ;
        RECT 126.095 191.170 126.385 191.910 ;
        RECT 126.555 191.340 126.825 192.085 ;
        RECT 120.080 190.945 126.825 191.170 ;
        RECT 127.635 191.155 127.805 191.915 ;
        RECT 128.020 191.325 128.350 192.085 ;
        RECT 127.635 190.985 128.350 191.155 ;
        RECT 128.520 191.010 128.775 191.915 ;
        RECT 115.085 190.445 115.375 190.775 ;
        RECT 115.545 190.525 115.875 190.775 ;
        RECT 116.105 190.525 116.795 190.775 ;
        RECT 115.205 190.355 115.375 190.445 ;
        RECT 115.205 190.165 116.595 190.355 ;
        RECT 117.885 190.215 118.200 190.775 ;
        RECT 118.370 190.525 125.490 190.775 ;
        RECT 114.665 189.705 115.215 189.995 ;
        RECT 115.385 189.535 115.635 189.995 ;
        RECT 116.265 189.805 116.595 190.165 ;
        RECT 117.885 189.535 118.190 190.045 ;
        RECT 118.370 189.715 118.620 190.525 ;
        RECT 118.790 189.535 119.050 190.060 ;
        RECT 119.230 189.715 119.480 190.525 ;
        RECT 125.660 190.355 126.825 190.945 ;
        RECT 127.545 190.435 127.900 190.805 ;
        RECT 128.180 190.775 128.350 190.985 ;
        RECT 128.180 190.445 128.435 190.775 ;
        RECT 120.080 190.185 126.825 190.355 ;
        RECT 128.180 190.255 128.350 190.445 ;
        RECT 128.605 190.280 128.775 191.010 ;
        RECT 128.950 190.935 129.210 192.085 ;
        RECT 129.385 190.930 129.725 191.915 ;
        RECT 129.895 191.655 130.305 192.085 ;
        RECT 131.050 191.665 131.380 192.085 ;
        RECT 131.550 191.485 131.875 191.915 ;
        RECT 129.895 191.315 131.875 191.485 ;
        RECT 119.650 189.535 119.910 190.095 ;
        RECT 120.080 189.730 120.340 190.185 ;
        RECT 120.510 189.535 120.770 190.015 ;
        RECT 120.940 189.730 121.200 190.185 ;
        RECT 121.370 189.535 121.630 190.015 ;
        RECT 121.800 189.730 122.060 190.185 ;
        RECT 122.230 189.535 122.475 190.015 ;
        RECT 122.645 189.730 122.920 190.185 ;
        RECT 123.090 189.535 123.335 190.015 ;
        RECT 123.505 189.730 123.765 190.185 ;
        RECT 123.945 189.535 124.195 190.015 ;
        RECT 124.365 189.730 124.625 190.185 ;
        RECT 124.805 189.535 125.055 190.015 ;
        RECT 125.225 189.730 125.485 190.185 ;
        RECT 125.665 189.535 125.925 190.015 ;
        RECT 126.095 189.730 126.355 190.185 ;
        RECT 127.635 190.085 128.350 190.255 ;
        RECT 126.525 189.535 126.825 190.015 ;
        RECT 127.635 189.705 127.805 190.085 ;
        RECT 128.020 189.535 128.350 189.915 ;
        RECT 128.520 189.705 128.775 190.280 ;
        RECT 128.950 189.535 129.210 190.375 ;
        RECT 129.385 190.275 129.640 190.930 ;
        RECT 129.895 190.775 130.160 191.315 ;
        RECT 130.375 190.975 131.000 191.145 ;
        RECT 129.810 190.445 130.160 190.775 ;
        RECT 130.330 190.445 130.660 190.775 ;
        RECT 130.830 190.275 131.000 190.975 ;
        RECT 129.385 189.900 129.745 190.275 ;
        RECT 129.445 189.875 129.615 189.900 ;
        RECT 130.010 189.535 130.180 190.275 ;
        RECT 130.460 190.105 131.000 190.275 ;
        RECT 131.170 190.905 131.875 191.315 ;
        RECT 132.350 190.985 132.680 192.085 ;
        RECT 133.075 191.135 133.350 191.905 ;
        RECT 133.520 191.475 133.850 191.905 ;
        RECT 134.020 191.645 134.215 192.085 ;
        RECT 134.395 191.475 134.725 191.905 ;
        RECT 133.520 191.305 134.725 191.475 ;
        RECT 133.075 190.945 133.660 191.135 ;
        RECT 133.830 190.975 134.725 191.305 ;
        RECT 134.905 190.995 136.115 192.085 ;
        RECT 130.460 189.900 130.630 190.105 ;
        RECT 131.170 189.705 131.340 190.905 ;
        RECT 131.510 190.525 132.080 190.735 ;
        RECT 132.250 190.525 132.895 190.735 ;
        RECT 131.570 190.185 132.740 190.355 ;
        RECT 131.570 189.705 131.900 190.185 ;
        RECT 132.070 189.535 132.240 190.005 ;
        RECT 132.410 189.720 132.740 190.185 ;
        RECT 133.075 190.125 133.315 190.775 ;
        RECT 133.485 190.275 133.660 190.945 ;
        RECT 133.830 190.445 134.245 190.775 ;
        RECT 134.425 190.445 134.720 190.775 ;
        RECT 134.905 190.455 135.425 190.995 ;
        RECT 133.485 190.095 133.815 190.275 ;
        RECT 133.090 189.535 133.420 189.925 ;
        RECT 133.590 189.715 133.815 190.095 ;
        RECT 134.015 189.825 134.245 190.445 ;
        RECT 135.595 190.285 136.115 190.825 ;
        RECT 134.425 189.535 134.725 190.265 ;
        RECT 134.905 189.535 136.115 190.285 ;
        RECT 23.500 189.365 136.200 189.535 ;
        RECT 23.585 188.615 24.795 189.365 ;
        RECT 23.585 188.075 24.105 188.615 ;
        RECT 24.965 188.595 27.555 189.365 ;
        RECT 27.725 188.690 27.985 189.195 ;
        RECT 28.165 188.985 28.495 189.365 ;
        RECT 28.675 188.815 28.845 189.195 ;
        RECT 29.105 188.820 34.450 189.365 ;
        RECT 24.275 187.905 24.795 188.445 ;
        RECT 24.965 188.075 26.175 188.595 ;
        RECT 26.345 187.905 27.555 188.425 ;
        RECT 23.585 186.815 24.795 187.905 ;
        RECT 24.965 186.815 27.555 187.905 ;
        RECT 27.725 187.890 27.895 188.690 ;
        RECT 28.180 188.645 28.845 188.815 ;
        RECT 28.180 188.390 28.350 188.645 ;
        RECT 28.065 188.060 28.350 188.390 ;
        RECT 28.585 188.095 28.915 188.465 ;
        RECT 28.180 187.915 28.350 188.060 ;
        RECT 30.690 187.990 31.030 188.820 ;
        RECT 34.625 188.595 37.215 189.365 ;
        RECT 37.850 188.625 38.105 189.195 ;
        RECT 38.275 188.965 38.605 189.365 ;
        RECT 39.030 188.830 39.560 189.195 ;
        RECT 39.750 189.025 40.025 189.195 ;
        RECT 39.745 188.855 40.025 189.025 ;
        RECT 39.030 188.795 39.205 188.830 ;
        RECT 38.275 188.625 39.205 188.795 ;
        RECT 27.725 186.985 27.995 187.890 ;
        RECT 28.180 187.745 28.845 187.915 ;
        RECT 28.165 186.815 28.495 187.575 ;
        RECT 28.675 186.985 28.845 187.745 ;
        RECT 32.510 187.250 32.860 188.500 ;
        RECT 34.625 188.075 35.835 188.595 ;
        RECT 36.005 187.905 37.215 188.425 ;
        RECT 29.105 186.815 34.450 187.250 ;
        RECT 34.625 186.815 37.215 187.905 ;
        RECT 37.850 187.955 38.020 188.625 ;
        RECT 38.275 188.455 38.445 188.625 ;
        RECT 38.190 188.125 38.445 188.455 ;
        RECT 38.670 188.125 38.865 188.455 ;
        RECT 37.850 186.985 38.185 187.955 ;
        RECT 38.355 186.815 38.525 187.955 ;
        RECT 38.695 187.155 38.865 188.125 ;
        RECT 39.035 187.495 39.205 188.625 ;
        RECT 39.375 187.835 39.545 188.635 ;
        RECT 39.750 188.035 40.025 188.855 ;
        RECT 40.195 187.835 40.385 189.195 ;
        RECT 40.565 188.830 41.075 189.365 ;
        RECT 41.295 188.555 41.540 189.160 ;
        RECT 41.985 188.595 44.575 189.365 ;
        RECT 44.910 188.855 45.150 189.365 ;
        RECT 45.330 188.855 45.610 189.185 ;
        RECT 45.840 188.855 46.055 189.365 ;
        RECT 40.585 188.385 41.815 188.555 ;
        RECT 39.375 187.665 40.385 187.835 ;
        RECT 40.555 187.820 41.305 188.010 ;
        RECT 39.035 187.325 40.160 187.495 ;
        RECT 40.555 187.155 40.725 187.820 ;
        RECT 41.475 187.575 41.815 188.385 ;
        RECT 41.985 188.075 43.195 188.595 ;
        RECT 43.365 187.905 44.575 188.425 ;
        RECT 44.805 188.125 45.160 188.685 ;
        RECT 45.330 187.955 45.500 188.855 ;
        RECT 45.670 188.125 45.935 188.685 ;
        RECT 46.225 188.625 46.840 189.195 ;
        RECT 47.210 188.855 47.450 189.365 ;
        RECT 47.630 188.855 47.910 189.185 ;
        RECT 48.140 188.855 48.355 189.365 ;
        RECT 46.185 187.955 46.355 188.455 ;
        RECT 38.695 186.985 40.725 187.155 ;
        RECT 40.895 186.815 41.065 187.575 ;
        RECT 41.300 187.165 41.815 187.575 ;
        RECT 41.985 186.815 44.575 187.905 ;
        RECT 44.930 187.785 46.355 187.955 ;
        RECT 44.930 187.610 45.320 187.785 ;
        RECT 45.805 186.815 46.135 187.615 ;
        RECT 46.525 187.605 46.840 188.625 ;
        RECT 47.105 188.125 47.460 188.685 ;
        RECT 47.630 187.955 47.800 188.855 ;
        RECT 47.970 188.125 48.235 188.685 ;
        RECT 48.525 188.625 49.140 189.195 ;
        RECT 49.345 188.640 49.635 189.365 ;
        RECT 48.485 187.955 48.655 188.455 ;
        RECT 47.230 187.785 48.655 187.955 ;
        RECT 47.230 187.610 47.620 187.785 ;
        RECT 46.305 186.985 46.840 187.605 ;
        RECT 48.105 186.815 48.435 187.615 ;
        RECT 48.825 187.605 49.140 188.625 ;
        RECT 48.605 186.985 49.140 187.605 ;
        RECT 49.345 186.815 49.635 187.980 ;
        RECT 50.725 186.985 51.005 189.085 ;
        RECT 51.235 188.905 51.405 189.365 ;
        RECT 51.675 188.975 52.925 189.155 ;
        RECT 52.060 188.735 52.425 188.805 ;
        RECT 51.175 188.555 52.425 188.735 ;
        RECT 52.595 188.755 52.925 188.975 ;
        RECT 53.095 188.925 53.265 189.365 ;
        RECT 53.435 188.755 53.775 189.170 ;
        RECT 52.595 188.585 53.775 188.755 ;
        RECT 53.950 188.625 54.205 189.195 ;
        RECT 54.375 188.965 54.705 189.365 ;
        RECT 55.130 188.830 55.660 189.195 ;
        RECT 55.130 188.795 55.305 188.830 ;
        RECT 54.375 188.625 55.305 188.795 ;
        RECT 51.175 187.955 51.450 188.555 ;
        RECT 51.620 188.125 51.975 188.375 ;
        RECT 52.170 188.345 52.635 188.375 ;
        RECT 52.165 188.175 52.635 188.345 ;
        RECT 52.170 188.125 52.635 188.175 ;
        RECT 52.805 188.125 53.135 188.375 ;
        RECT 53.310 188.175 53.775 188.375 ;
        RECT 52.955 188.005 53.135 188.125 ;
        RECT 51.175 187.745 52.785 187.955 ;
        RECT 52.955 187.835 53.285 188.005 ;
        RECT 52.375 187.645 52.785 187.745 ;
        RECT 51.195 186.815 51.980 187.575 ;
        RECT 52.375 186.985 52.760 187.645 ;
        RECT 53.085 187.045 53.285 187.835 ;
        RECT 53.455 186.815 53.775 187.995 ;
        RECT 53.950 187.955 54.120 188.625 ;
        RECT 54.375 188.455 54.545 188.625 ;
        RECT 54.290 188.125 54.545 188.455 ;
        RECT 54.770 188.125 54.965 188.455 ;
        RECT 53.950 186.985 54.285 187.955 ;
        RECT 54.455 186.815 54.625 187.955 ;
        RECT 54.795 187.155 54.965 188.125 ;
        RECT 55.135 187.495 55.305 188.625 ;
        RECT 55.475 187.835 55.645 188.635 ;
        RECT 55.850 188.345 56.125 189.195 ;
        RECT 55.845 188.175 56.125 188.345 ;
        RECT 55.850 188.035 56.125 188.175 ;
        RECT 56.295 187.835 56.485 189.195 ;
        RECT 56.665 188.830 57.175 189.365 ;
        RECT 57.395 188.555 57.640 189.160 ;
        RECT 58.090 188.625 58.345 189.195 ;
        RECT 58.515 188.965 58.845 189.365 ;
        RECT 59.270 188.830 59.800 189.195 ;
        RECT 59.270 188.795 59.445 188.830 ;
        RECT 58.515 188.625 59.445 188.795 ;
        RECT 56.685 188.385 57.915 188.555 ;
        RECT 55.475 187.665 56.485 187.835 ;
        RECT 56.655 187.820 57.405 188.010 ;
        RECT 55.135 187.325 56.260 187.495 ;
        RECT 56.655 187.155 56.825 187.820 ;
        RECT 57.575 187.575 57.915 188.385 ;
        RECT 54.795 186.985 56.825 187.155 ;
        RECT 56.995 186.815 57.165 187.575 ;
        RECT 57.400 187.165 57.915 187.575 ;
        RECT 58.090 187.955 58.260 188.625 ;
        RECT 58.515 188.455 58.685 188.625 ;
        RECT 58.430 188.125 58.685 188.455 ;
        RECT 58.910 188.125 59.105 188.455 ;
        RECT 58.090 186.985 58.425 187.955 ;
        RECT 58.595 186.815 58.765 187.955 ;
        RECT 58.935 187.155 59.105 188.125 ;
        RECT 59.275 187.495 59.445 188.625 ;
        RECT 59.615 187.835 59.785 188.635 ;
        RECT 59.990 188.345 60.265 189.195 ;
        RECT 59.985 188.175 60.265 188.345 ;
        RECT 59.990 188.035 60.265 188.175 ;
        RECT 60.435 187.835 60.625 189.195 ;
        RECT 60.805 188.830 61.315 189.365 ;
        RECT 61.535 188.555 61.780 189.160 ;
        RECT 62.685 188.565 63.380 189.195 ;
        RECT 63.585 188.565 63.895 189.365 ;
        RECT 65.005 188.635 65.295 189.365 ;
        RECT 60.825 188.385 62.055 188.555 ;
        RECT 63.205 188.515 63.380 188.565 ;
        RECT 59.615 187.665 60.625 187.835 ;
        RECT 60.795 187.820 61.545 188.010 ;
        RECT 59.275 187.325 60.400 187.495 ;
        RECT 60.795 187.155 60.965 187.820 ;
        RECT 61.715 187.575 62.055 188.385 ;
        RECT 62.705 188.125 63.040 188.375 ;
        RECT 63.210 187.965 63.380 188.515 ;
        RECT 63.550 188.125 63.885 188.395 ;
        RECT 64.995 188.125 65.295 188.455 ;
        RECT 65.475 188.435 65.705 189.075 ;
        RECT 65.885 188.815 66.195 189.185 ;
        RECT 66.375 188.995 67.045 189.365 ;
        RECT 65.885 188.615 67.115 188.815 ;
        RECT 65.475 188.125 66.000 188.435 ;
        RECT 66.180 188.125 66.645 188.435 ;
        RECT 58.935 186.985 60.965 187.155 ;
        RECT 61.135 186.815 61.305 187.575 ;
        RECT 61.540 187.165 62.055 187.575 ;
        RECT 62.685 186.815 62.945 187.955 ;
        RECT 63.115 186.985 63.445 187.965 ;
        RECT 63.615 186.815 63.895 187.955 ;
        RECT 66.825 187.945 67.115 188.615 ;
        RECT 65.005 187.705 66.165 187.945 ;
        RECT 65.005 186.995 65.265 187.705 ;
        RECT 65.435 186.815 65.765 187.525 ;
        RECT 65.935 186.995 66.165 187.705 ;
        RECT 66.345 187.725 67.115 187.945 ;
        RECT 66.345 186.995 66.615 187.725 ;
        RECT 66.795 186.815 67.135 187.545 ;
        RECT 67.305 186.995 67.565 189.185 ;
        RECT 67.795 188.565 68.005 189.365 ;
        RECT 67.795 186.815 68.005 187.955 ;
        RECT 68.175 186.985 68.515 189.195 ;
        RECT 68.695 188.905 68.945 189.365 ;
        RECT 69.135 188.735 69.465 189.195 ;
        RECT 68.690 188.565 69.465 188.735 ;
        RECT 69.665 188.685 70.050 189.195 ;
        RECT 68.690 187.665 68.965 188.565 ;
        RECT 69.645 188.515 70.050 188.685 ;
        RECT 70.525 188.825 70.855 189.195 ;
        RECT 71.045 188.995 71.375 189.365 ;
        RECT 71.545 188.825 71.875 189.195 ;
        RECT 70.525 188.625 71.875 188.825 ;
        RECT 69.165 187.835 69.495 188.375 ;
        RECT 69.665 187.835 70.050 188.515 ;
        RECT 72.345 188.595 74.935 189.365 ;
        RECT 75.105 188.640 75.395 189.365 ;
        RECT 75.565 188.595 78.155 189.365 ;
        RECT 78.330 188.625 78.585 189.195 ;
        RECT 78.755 188.965 79.085 189.365 ;
        RECT 79.510 188.830 80.040 189.195 ;
        RECT 79.510 188.795 79.685 188.830 ;
        RECT 78.755 188.625 79.685 188.795 ;
        RECT 70.340 187.835 70.760 188.375 ;
        RECT 70.960 188.125 71.320 188.455 ;
        RECT 71.490 188.135 72.175 188.445 ;
        RECT 68.690 187.425 70.855 187.665 ;
        RECT 68.695 186.815 69.315 187.255 ;
        RECT 69.520 186.985 69.800 187.425 ;
        RECT 69.985 186.815 70.315 187.195 ;
        RECT 70.525 186.985 70.855 187.425 ;
        RECT 71.030 187.080 71.320 188.125 ;
        RECT 71.545 186.815 71.800 187.955 ;
        RECT 71.970 187.095 72.175 188.135 ;
        RECT 72.345 188.075 73.555 188.595 ;
        RECT 73.725 187.905 74.935 188.425 ;
        RECT 75.565 188.075 76.775 188.595 ;
        RECT 72.345 186.815 74.935 187.905 ;
        RECT 75.105 186.815 75.395 187.980 ;
        RECT 76.945 187.905 78.155 188.425 ;
        RECT 75.565 186.815 78.155 187.905 ;
        RECT 78.330 187.955 78.500 188.625 ;
        RECT 78.755 188.455 78.925 188.625 ;
        RECT 78.670 188.125 78.925 188.455 ;
        RECT 79.150 188.125 79.345 188.455 ;
        RECT 78.330 186.985 78.665 187.955 ;
        RECT 78.835 186.815 79.005 187.955 ;
        RECT 79.175 187.155 79.345 188.125 ;
        RECT 79.515 187.495 79.685 188.625 ;
        RECT 79.855 187.835 80.025 188.635 ;
        RECT 80.230 188.345 80.505 189.195 ;
        RECT 80.225 188.175 80.505 188.345 ;
        RECT 80.230 188.035 80.505 188.175 ;
        RECT 80.675 187.835 80.865 189.195 ;
        RECT 81.045 188.830 81.555 189.365 ;
        RECT 81.775 188.555 82.020 189.160 ;
        RECT 82.470 188.625 82.725 189.195 ;
        RECT 82.895 188.965 83.225 189.365 ;
        RECT 83.650 188.830 84.180 189.195 ;
        RECT 83.650 188.795 83.825 188.830 ;
        RECT 82.895 188.625 83.825 188.795 ;
        RECT 81.065 188.385 82.295 188.555 ;
        RECT 79.855 187.665 80.865 187.835 ;
        RECT 81.035 187.820 81.785 188.010 ;
        RECT 79.515 187.325 80.640 187.495 ;
        RECT 81.035 187.155 81.205 187.820 ;
        RECT 81.955 187.575 82.295 188.385 ;
        RECT 79.175 186.985 81.205 187.155 ;
        RECT 81.375 186.815 81.545 187.575 ;
        RECT 81.780 187.165 82.295 187.575 ;
        RECT 82.470 187.955 82.640 188.625 ;
        RECT 82.895 188.455 83.065 188.625 ;
        RECT 82.810 188.125 83.065 188.455 ;
        RECT 83.290 188.125 83.485 188.455 ;
        RECT 82.470 186.985 82.805 187.955 ;
        RECT 82.975 186.815 83.145 187.955 ;
        RECT 83.315 187.155 83.485 188.125 ;
        RECT 83.655 187.495 83.825 188.625 ;
        RECT 83.995 187.835 84.165 188.635 ;
        RECT 84.370 188.345 84.645 189.195 ;
        RECT 84.365 188.175 84.645 188.345 ;
        RECT 84.370 188.035 84.645 188.175 ;
        RECT 84.815 187.835 85.005 189.195 ;
        RECT 85.185 188.830 85.695 189.365 ;
        RECT 85.915 188.555 86.160 189.160 ;
        RECT 86.605 188.595 88.275 189.365 ;
        RECT 85.205 188.385 86.435 188.555 ;
        RECT 83.995 187.665 85.005 187.835 ;
        RECT 85.175 187.820 85.925 188.010 ;
        RECT 83.655 187.325 84.780 187.495 ;
        RECT 85.175 187.155 85.345 187.820 ;
        RECT 86.095 187.575 86.435 188.385 ;
        RECT 86.605 188.075 87.355 188.595 ;
        RECT 87.525 187.905 88.275 188.425 ;
        RECT 83.315 186.985 85.345 187.155 ;
        RECT 85.515 186.815 85.685 187.575 ;
        RECT 85.920 187.165 86.435 187.575 ;
        RECT 86.605 186.815 88.275 187.905 ;
        RECT 88.455 186.995 88.715 189.185 ;
        RECT 88.975 188.995 89.645 189.365 ;
        RECT 89.825 188.815 90.135 189.185 ;
        RECT 88.905 188.615 90.135 188.815 ;
        RECT 88.905 187.945 89.195 188.615 ;
        RECT 90.315 188.435 90.545 189.075 ;
        RECT 90.725 188.635 91.015 189.365 ;
        RECT 92.135 188.635 92.435 189.365 ;
        RECT 92.615 188.455 92.845 189.075 ;
        RECT 93.045 188.805 93.270 189.185 ;
        RECT 93.440 188.975 93.770 189.365 ;
        RECT 94.885 188.865 95.145 189.195 ;
        RECT 95.315 189.005 95.645 189.365 ;
        RECT 95.900 188.985 97.200 189.195 ;
        RECT 93.045 188.625 93.375 188.805 ;
        RECT 89.375 188.125 89.840 188.435 ;
        RECT 90.020 188.125 90.545 188.435 ;
        RECT 90.725 188.125 91.025 188.455 ;
        RECT 92.140 188.125 92.435 188.455 ;
        RECT 92.615 188.125 93.030 188.455 ;
        RECT 93.200 187.955 93.375 188.625 ;
        RECT 93.545 188.125 93.785 188.775 ;
        RECT 88.905 187.725 89.675 187.945 ;
        RECT 88.885 186.815 89.225 187.545 ;
        RECT 89.405 186.995 89.675 187.725 ;
        RECT 89.855 187.705 91.015 187.945 ;
        RECT 89.855 186.995 90.085 187.705 ;
        RECT 90.255 186.815 90.585 187.525 ;
        RECT 90.755 186.995 91.015 187.705 ;
        RECT 92.135 187.595 93.030 187.925 ;
        RECT 93.200 187.765 93.785 187.955 ;
        RECT 92.135 187.425 93.340 187.595 ;
        RECT 92.135 186.995 92.465 187.425 ;
        RECT 92.645 186.815 92.840 187.255 ;
        RECT 93.010 186.995 93.340 187.425 ;
        RECT 93.510 186.995 93.785 187.765 ;
        RECT 94.885 187.665 95.055 188.865 ;
        RECT 95.900 188.835 96.070 188.985 ;
        RECT 95.315 188.710 96.070 188.835 ;
        RECT 95.225 188.665 96.070 188.710 ;
        RECT 95.225 188.545 95.495 188.665 ;
        RECT 95.225 187.970 95.395 188.545 ;
        RECT 95.625 188.105 96.035 188.410 ;
        RECT 96.325 188.375 96.535 188.775 ;
        RECT 96.205 188.165 96.535 188.375 ;
        RECT 96.780 188.375 97.000 188.775 ;
        RECT 97.475 188.600 97.930 189.365 ;
        RECT 98.130 188.975 98.460 189.365 ;
        RECT 98.630 188.805 98.855 189.185 ;
        RECT 96.780 188.165 97.255 188.375 ;
        RECT 97.445 188.175 97.935 188.375 ;
        RECT 98.115 188.125 98.355 188.775 ;
        RECT 98.525 188.625 98.855 188.805 ;
        RECT 95.225 187.935 95.425 187.970 ;
        RECT 96.755 187.935 97.930 187.995 ;
        RECT 98.525 187.955 98.700 188.625 ;
        RECT 99.055 188.455 99.285 189.075 ;
        RECT 99.465 188.635 99.765 189.365 ;
        RECT 100.865 188.640 101.155 189.365 ;
        RECT 101.365 188.545 101.595 189.365 ;
        RECT 101.765 188.565 102.095 189.195 ;
        RECT 98.870 188.125 99.285 188.455 ;
        RECT 99.465 188.125 99.760 188.455 ;
        RECT 101.345 188.125 101.675 188.375 ;
        RECT 95.225 187.825 97.930 187.935 ;
        RECT 95.285 187.765 97.085 187.825 ;
        RECT 96.755 187.735 97.085 187.765 ;
        RECT 94.885 186.985 95.145 187.665 ;
        RECT 95.315 186.815 95.565 187.595 ;
        RECT 95.815 187.565 96.650 187.575 ;
        RECT 97.240 187.565 97.425 187.655 ;
        RECT 95.815 187.365 97.425 187.565 ;
        RECT 95.815 186.985 96.065 187.365 ;
        RECT 97.195 187.325 97.425 187.365 ;
        RECT 97.675 187.205 97.930 187.825 ;
        RECT 96.235 186.815 96.590 187.195 ;
        RECT 97.595 186.985 97.930 187.205 ;
        RECT 98.115 187.765 98.700 187.955 ;
        RECT 98.115 186.995 98.390 187.765 ;
        RECT 98.870 187.595 99.765 187.925 ;
        RECT 98.560 187.425 99.765 187.595 ;
        RECT 98.560 186.995 98.890 187.425 ;
        RECT 99.060 186.815 99.255 187.255 ;
        RECT 99.435 186.995 99.765 187.425 ;
        RECT 100.865 186.815 101.155 187.980 ;
        RECT 101.845 187.965 102.095 188.565 ;
        RECT 102.265 188.545 102.475 189.365 ;
        RECT 103.175 188.645 103.505 189.365 ;
        RECT 104.050 188.965 105.665 189.135 ;
        RECT 105.835 188.965 106.165 189.365 ;
        RECT 105.495 188.795 105.665 188.965 ;
        RECT 106.335 188.890 106.670 189.150 ;
        RECT 103.230 188.125 103.580 188.455 ;
        RECT 103.890 188.125 104.310 188.790 ;
        RECT 104.480 188.685 104.770 188.785 ;
        RECT 104.960 188.685 105.230 188.785 ;
        RECT 104.480 188.515 104.775 188.685 ;
        RECT 104.960 188.515 105.235 188.685 ;
        RECT 105.495 188.625 106.055 188.795 ;
        RECT 104.480 188.125 104.770 188.515 ;
        RECT 104.960 188.125 105.230 188.515 ;
        RECT 105.885 188.455 106.055 188.625 ;
        RECT 105.440 188.345 105.690 188.455 ;
        RECT 105.440 188.175 105.695 188.345 ;
        RECT 105.440 188.125 105.690 188.175 ;
        RECT 105.885 188.125 106.190 188.455 ;
        RECT 103.230 188.005 103.435 188.125 ;
        RECT 101.365 186.815 101.595 187.955 ;
        RECT 101.765 186.985 102.095 187.965 ;
        RECT 102.265 186.815 102.475 187.955 ;
        RECT 103.225 187.835 103.435 188.005 ;
        RECT 105.885 187.955 106.055 188.125 ;
        RECT 103.685 187.785 106.055 187.955 ;
        RECT 103.255 187.155 103.425 187.655 ;
        RECT 103.685 187.325 103.855 187.785 ;
        RECT 104.085 187.405 105.510 187.575 ;
        RECT 104.085 187.155 104.415 187.405 ;
        RECT 103.255 186.985 104.415 187.155 ;
        RECT 104.640 186.815 104.970 187.235 ;
        RECT 105.225 186.985 105.510 187.405 ;
        RECT 105.755 186.815 106.085 187.615 ;
        RECT 106.415 187.535 106.670 188.890 ;
        RECT 106.865 188.555 107.105 189.365 ;
        RECT 107.275 188.555 107.605 189.195 ;
        RECT 107.775 188.555 108.045 189.365 ;
        RECT 108.315 188.885 108.615 189.365 ;
        RECT 108.785 188.715 109.045 189.170 ;
        RECT 109.215 188.885 109.475 189.365 ;
        RECT 109.655 188.715 109.915 189.170 ;
        RECT 110.085 188.885 110.335 189.365 ;
        RECT 110.515 188.715 110.775 189.170 ;
        RECT 110.945 188.885 111.195 189.365 ;
        RECT 111.375 188.715 111.635 189.170 ;
        RECT 111.805 188.885 112.050 189.365 ;
        RECT 112.220 188.715 112.495 189.170 ;
        RECT 112.665 188.885 112.910 189.365 ;
        RECT 113.080 188.715 113.340 189.170 ;
        RECT 113.510 188.885 113.770 189.365 ;
        RECT 113.940 188.715 114.200 189.170 ;
        RECT 114.370 188.885 114.630 189.365 ;
        RECT 114.800 188.715 115.060 189.170 ;
        RECT 115.230 188.805 115.490 189.365 ;
        RECT 106.845 188.125 107.195 188.375 ;
        RECT 107.365 187.955 107.535 188.555 ;
        RECT 108.315 188.545 115.060 188.715 ;
        RECT 107.705 188.125 108.055 188.375 ;
        RECT 108.315 187.955 109.480 188.545 ;
        RECT 115.660 188.375 115.910 189.185 ;
        RECT 116.090 188.840 116.350 189.365 ;
        RECT 116.520 188.375 116.770 189.185 ;
        RECT 116.950 188.855 117.255 189.365 ;
        RECT 109.650 188.125 116.770 188.375 ;
        RECT 116.940 188.125 117.255 188.685 ;
        RECT 117.975 188.545 118.145 189.365 ;
        RECT 118.315 188.545 118.645 189.190 ;
        RECT 118.835 188.715 119.165 189.190 ;
        RECT 119.335 188.885 119.505 189.365 ;
        RECT 119.675 188.715 120.005 189.190 ;
        RECT 120.175 188.885 120.345 189.365 ;
        RECT 120.515 188.715 120.845 189.190 ;
        RECT 121.015 188.885 121.185 189.365 ;
        RECT 121.355 188.715 121.685 189.190 ;
        RECT 121.855 188.885 122.025 189.365 ;
        RECT 122.195 188.715 122.525 189.190 ;
        RECT 122.695 188.885 122.865 189.365 ;
        RECT 123.035 188.715 123.365 189.190 ;
        RECT 123.535 188.885 123.705 189.365 ;
        RECT 124.325 188.860 124.610 189.365 ;
        RECT 118.835 188.545 120.345 188.715 ;
        RECT 120.515 188.545 124.155 188.715 ;
        RECT 124.780 188.690 125.105 189.195 ;
        RECT 118.475 188.375 118.645 188.545 ;
        RECT 120.175 188.375 120.345 188.545 ;
        RECT 117.885 188.175 118.305 188.375 ;
        RECT 118.475 188.175 120.005 188.375 ;
        RECT 120.175 188.175 123.560 188.375 ;
        RECT 106.335 187.025 106.670 187.535 ;
        RECT 106.855 187.785 107.535 187.955 ;
        RECT 106.855 187.000 107.185 187.785 ;
        RECT 107.715 186.815 108.045 187.955 ;
        RECT 108.315 187.730 115.060 187.955 ;
        RECT 108.315 186.815 108.585 187.560 ;
        RECT 108.755 186.990 109.045 187.730 ;
        RECT 109.655 187.715 115.060 187.730 ;
        RECT 109.215 186.820 109.470 187.545 ;
        RECT 109.655 186.990 109.915 187.715 ;
        RECT 110.085 186.820 110.330 187.545 ;
        RECT 110.515 186.990 110.775 187.715 ;
        RECT 110.945 186.820 111.190 187.545 ;
        RECT 111.375 186.990 111.635 187.715 ;
        RECT 111.805 186.820 112.050 187.545 ;
        RECT 112.220 186.990 112.480 187.715 ;
        RECT 112.650 186.820 112.910 187.545 ;
        RECT 113.080 186.990 113.340 187.715 ;
        RECT 113.510 186.820 113.770 187.545 ;
        RECT 113.940 186.990 114.200 187.715 ;
        RECT 114.370 186.820 114.630 187.545 ;
        RECT 114.800 186.990 115.060 187.715 ;
        RECT 115.230 186.820 115.490 187.615 ;
        RECT 115.660 186.990 115.910 188.125 ;
        RECT 109.215 186.815 115.490 186.820 ;
        RECT 116.090 186.815 116.350 187.625 ;
        RECT 116.525 186.985 116.770 188.125 ;
        RECT 116.950 186.815 117.245 187.625 ;
        RECT 117.975 186.815 118.145 188.005 ;
        RECT 118.475 187.905 118.645 188.175 ;
        RECT 120.175 188.005 120.345 188.175 ;
        RECT 123.770 188.005 124.155 188.545 ;
        RECT 124.325 188.160 125.105 188.690 ;
        RECT 118.315 186.985 118.645 187.905 ;
        RECT 118.835 187.835 120.345 188.005 ;
        RECT 120.515 187.835 124.155 188.005 ;
        RECT 118.835 186.985 119.165 187.835 ;
        RECT 119.335 186.815 119.505 187.665 ;
        RECT 119.675 186.985 120.005 187.835 ;
        RECT 120.175 186.815 120.345 187.665 ;
        RECT 120.515 186.985 120.845 187.835 ;
        RECT 121.015 186.815 121.185 187.615 ;
        RECT 121.355 186.985 121.685 187.835 ;
        RECT 121.855 186.815 122.025 187.615 ;
        RECT 122.195 186.985 122.525 187.835 ;
        RECT 122.695 186.815 122.865 187.615 ;
        RECT 123.035 186.985 123.365 187.835 ;
        RECT 123.535 186.815 123.705 187.615 ;
        RECT 124.325 186.815 124.605 187.785 ;
        RECT 124.775 186.985 125.105 188.160 ;
        RECT 125.295 188.125 125.535 189.075 ;
        RECT 126.625 188.640 126.915 189.365 ;
        RECT 127.085 188.690 127.345 189.195 ;
        RECT 127.525 188.985 127.855 189.365 ;
        RECT 128.035 188.815 128.205 189.195 ;
        RECT 125.275 186.815 125.535 187.785 ;
        RECT 126.625 186.815 126.915 187.980 ;
        RECT 127.085 187.890 127.265 188.690 ;
        RECT 127.540 188.645 128.205 188.815 ;
        RECT 129.540 188.715 129.870 189.180 ;
        RECT 130.040 188.895 130.210 189.365 ;
        RECT 130.380 188.715 130.710 189.195 ;
        RECT 127.540 188.390 127.710 188.645 ;
        RECT 129.540 188.545 130.710 188.715 ;
        RECT 127.435 188.060 127.710 188.390 ;
        RECT 127.935 188.095 128.275 188.465 ;
        RECT 129.385 188.165 130.030 188.375 ;
        RECT 130.200 188.165 130.770 188.375 ;
        RECT 127.540 187.915 127.710 188.060 ;
        RECT 130.940 187.995 131.110 189.195 ;
        RECT 131.650 188.795 131.820 189.000 ;
        RECT 127.085 186.985 127.355 187.890 ;
        RECT 127.540 187.745 128.215 187.915 ;
        RECT 127.525 186.815 127.855 187.575 ;
        RECT 128.035 186.985 128.215 187.745 ;
        RECT 129.600 186.815 129.930 187.915 ;
        RECT 130.405 187.585 131.110 187.995 ;
        RECT 131.280 188.625 131.820 188.795 ;
        RECT 132.100 188.625 132.270 189.365 ;
        RECT 132.535 188.625 132.895 189.000 ;
        RECT 133.155 188.815 133.325 189.195 ;
        RECT 133.540 188.985 133.870 189.365 ;
        RECT 133.155 188.645 133.870 188.815 ;
        RECT 131.280 187.925 131.450 188.625 ;
        RECT 131.620 188.125 131.950 188.455 ;
        RECT 132.120 188.125 132.470 188.455 ;
        RECT 131.280 187.755 131.905 187.925 ;
        RECT 132.120 187.585 132.385 188.125 ;
        RECT 132.640 187.970 132.895 188.625 ;
        RECT 133.065 188.095 133.420 188.465 ;
        RECT 133.700 188.455 133.870 188.645 ;
        RECT 134.040 188.620 134.295 189.195 ;
        RECT 133.700 188.125 133.955 188.455 ;
        RECT 130.405 187.415 132.385 187.585 ;
        RECT 130.405 186.985 130.730 187.415 ;
        RECT 130.900 186.815 131.230 187.235 ;
        RECT 131.975 186.815 132.385 187.245 ;
        RECT 132.555 186.985 132.895 187.970 ;
        RECT 133.700 187.915 133.870 188.125 ;
        RECT 133.155 187.745 133.870 187.915 ;
        RECT 134.125 187.890 134.295 188.620 ;
        RECT 134.470 188.525 134.730 189.365 ;
        RECT 134.905 188.615 136.115 189.365 ;
        RECT 133.155 186.985 133.325 187.745 ;
        RECT 133.540 186.815 133.870 187.575 ;
        RECT 134.040 186.985 134.295 187.890 ;
        RECT 134.470 186.815 134.730 187.965 ;
        RECT 134.905 187.905 135.425 188.445 ;
        RECT 135.595 188.075 136.115 188.615 ;
        RECT 134.905 186.815 136.115 187.905 ;
        RECT 23.500 186.645 136.200 186.815 ;
        RECT 23.585 185.555 24.795 186.645 ;
        RECT 24.965 186.210 30.310 186.645 ;
        RECT 23.585 184.845 24.105 185.385 ;
        RECT 24.275 185.015 24.795 185.555 ;
        RECT 23.585 184.095 24.795 184.845 ;
        RECT 26.550 184.640 26.890 185.470 ;
        RECT 28.370 184.960 28.720 186.210 ;
        RECT 30.485 185.555 33.075 186.645 ;
        RECT 30.485 184.865 31.695 185.385 ;
        RECT 31.865 185.035 33.075 185.555 ;
        RECT 24.965 184.095 30.310 184.640 ;
        RECT 30.485 184.095 33.075 184.865 ;
        RECT 33.245 184.375 33.525 186.475 ;
        RECT 33.715 185.885 34.500 186.645 ;
        RECT 34.895 185.815 35.280 186.475 ;
        RECT 34.895 185.715 35.305 185.815 ;
        RECT 33.695 185.505 35.305 185.715 ;
        RECT 35.605 185.625 35.805 186.415 ;
        RECT 33.695 184.905 33.970 185.505 ;
        RECT 35.475 185.455 35.805 185.625 ;
        RECT 35.975 185.465 36.295 186.645 ;
        RECT 36.465 185.480 36.755 186.645 ;
        RECT 36.930 185.505 37.265 186.475 ;
        RECT 37.435 185.505 37.605 186.645 ;
        RECT 37.775 186.305 39.805 186.475 ;
        RECT 35.475 185.335 35.655 185.455 ;
        RECT 34.140 185.085 34.495 185.335 ;
        RECT 34.690 185.285 35.155 185.335 ;
        RECT 34.685 185.115 35.155 185.285 ;
        RECT 34.690 185.085 35.155 185.115 ;
        RECT 35.325 185.085 35.655 185.335 ;
        RECT 35.830 185.085 36.295 185.285 ;
        RECT 33.695 184.725 34.945 184.905 ;
        RECT 34.580 184.655 34.945 184.725 ;
        RECT 35.115 184.705 36.295 184.875 ;
        RECT 36.930 184.835 37.100 185.505 ;
        RECT 37.775 185.335 37.945 186.305 ;
        RECT 37.270 185.005 37.525 185.335 ;
        RECT 37.750 185.005 37.945 185.335 ;
        RECT 38.115 185.965 39.240 186.135 ;
        RECT 37.355 184.835 37.525 185.005 ;
        RECT 38.115 184.835 38.285 185.965 ;
        RECT 33.755 184.095 33.925 184.555 ;
        RECT 35.115 184.485 35.445 184.705 ;
        RECT 34.195 184.305 35.445 184.485 ;
        RECT 35.615 184.095 35.785 184.535 ;
        RECT 35.955 184.290 36.295 184.705 ;
        RECT 36.465 184.095 36.755 184.820 ;
        RECT 36.930 184.265 37.185 184.835 ;
        RECT 37.355 184.665 38.285 184.835 ;
        RECT 38.455 185.625 39.465 185.795 ;
        RECT 38.455 184.825 38.625 185.625 ;
        RECT 38.110 184.630 38.285 184.665 ;
        RECT 37.355 184.095 37.685 184.495 ;
        RECT 38.110 184.265 38.640 184.630 ;
        RECT 38.830 184.605 39.105 185.425 ;
        RECT 38.825 184.435 39.105 184.605 ;
        RECT 38.830 184.265 39.105 184.435 ;
        RECT 39.275 184.265 39.465 185.625 ;
        RECT 39.635 185.640 39.805 186.305 ;
        RECT 39.975 185.885 40.145 186.645 ;
        RECT 40.380 185.885 40.895 186.295 ;
        RECT 41.265 185.975 41.545 186.645 ;
        RECT 39.635 185.450 40.385 185.640 ;
        RECT 40.555 185.075 40.895 185.885 ;
        RECT 41.065 185.335 41.380 185.775 ;
        RECT 41.715 185.755 42.015 186.305 ;
        RECT 42.225 185.925 42.555 186.645 ;
        RECT 42.745 185.925 43.195 186.475 ;
        RECT 41.715 185.585 42.655 185.755 ;
        RECT 42.485 185.335 42.655 185.585 ;
        RECT 41.065 185.085 41.755 185.335 ;
        RECT 41.985 185.085 42.315 185.335 ;
        RECT 39.665 184.905 40.895 185.075 ;
        RECT 42.485 185.005 42.775 185.335 ;
        RECT 42.485 184.915 42.655 185.005 ;
        RECT 39.645 184.095 40.155 184.630 ;
        RECT 40.375 184.300 40.620 184.905 ;
        RECT 41.265 184.725 42.655 184.915 ;
        RECT 41.265 184.365 41.595 184.725 ;
        RECT 42.945 184.555 43.195 185.925 ;
        RECT 43.365 185.505 43.655 186.645 ;
        RECT 43.825 185.505 44.105 186.645 ;
        RECT 44.275 185.495 44.605 186.475 ;
        RECT 44.775 185.505 45.035 186.645 ;
        RECT 45.665 185.505 45.925 186.645 ;
        RECT 46.095 185.495 46.425 186.475 ;
        RECT 46.595 185.505 46.875 186.645 ;
        RECT 47.975 186.035 48.305 186.465 ;
        RECT 48.485 186.205 48.680 186.645 ;
        RECT 48.850 186.035 49.180 186.465 ;
        RECT 47.975 185.865 49.180 186.035 ;
        RECT 47.975 185.535 48.870 185.865 ;
        RECT 49.350 185.695 49.625 186.465 ;
        RECT 49.040 185.505 49.625 185.695 ;
        RECT 49.825 185.755 50.085 186.465 ;
        RECT 50.255 185.935 50.585 186.645 ;
        RECT 50.755 185.755 50.985 186.465 ;
        RECT 49.825 185.515 50.985 185.755 ;
        RECT 51.165 185.735 51.435 186.465 ;
        RECT 51.615 185.915 51.955 186.645 ;
        RECT 51.165 185.515 51.935 185.735 ;
        RECT 44.340 185.455 44.515 185.495 ;
        RECT 43.835 185.065 44.170 185.335 ;
        RECT 44.340 184.895 44.510 185.455 ;
        RECT 44.680 185.085 45.015 185.335 ;
        RECT 45.685 185.085 46.020 185.335 ;
        RECT 46.190 184.895 46.360 185.495 ;
        RECT 46.530 185.065 46.865 185.335 ;
        RECT 47.980 185.005 48.275 185.335 ;
        RECT 48.455 185.005 48.870 185.335 ;
        RECT 42.225 184.095 42.475 184.555 ;
        RECT 42.645 184.265 43.195 184.555 ;
        RECT 43.365 184.095 43.655 184.895 ;
        RECT 43.825 184.095 44.135 184.895 ;
        RECT 44.340 184.265 45.035 184.895 ;
        RECT 45.665 184.265 46.360 184.895 ;
        RECT 46.565 184.095 46.875 184.895 ;
        RECT 47.975 184.095 48.275 184.825 ;
        RECT 48.455 184.385 48.685 185.005 ;
        RECT 49.040 184.835 49.215 185.505 ;
        RECT 48.885 184.655 49.215 184.835 ;
        RECT 49.385 184.685 49.625 185.335 ;
        RECT 49.815 185.005 50.115 185.335 ;
        RECT 50.295 185.025 50.820 185.335 ;
        RECT 51.000 185.025 51.465 185.335 ;
        RECT 48.885 184.275 49.110 184.655 ;
        RECT 49.280 184.095 49.610 184.485 ;
        RECT 49.825 184.095 50.115 184.825 ;
        RECT 50.295 184.385 50.525 185.025 ;
        RECT 51.645 184.845 51.935 185.515 ;
        RECT 50.705 184.645 51.935 184.845 ;
        RECT 50.705 184.275 51.015 184.645 ;
        RECT 51.195 184.095 51.865 184.465 ;
        RECT 52.125 184.275 52.385 186.465 ;
        RECT 52.565 185.555 53.775 186.645 ;
        RECT 52.565 184.845 53.085 185.385 ;
        RECT 53.255 185.015 53.775 185.555 ;
        RECT 53.950 185.505 54.285 186.475 ;
        RECT 54.455 185.505 54.625 186.645 ;
        RECT 54.795 186.305 56.825 186.475 ;
        RECT 52.565 184.095 53.775 184.845 ;
        RECT 53.950 184.835 54.120 185.505 ;
        RECT 54.795 185.335 54.965 186.305 ;
        RECT 54.290 185.005 54.545 185.335 ;
        RECT 54.770 185.005 54.965 185.335 ;
        RECT 55.135 185.965 56.260 186.135 ;
        RECT 54.375 184.835 54.545 185.005 ;
        RECT 55.135 184.835 55.305 185.965 ;
        RECT 53.950 184.265 54.205 184.835 ;
        RECT 54.375 184.665 55.305 184.835 ;
        RECT 55.475 185.625 56.485 185.795 ;
        RECT 55.475 184.825 55.645 185.625 ;
        RECT 55.130 184.630 55.305 184.665 ;
        RECT 54.375 184.095 54.705 184.495 ;
        RECT 55.130 184.265 55.660 184.630 ;
        RECT 55.850 184.605 56.125 185.425 ;
        RECT 55.845 184.435 56.125 184.605 ;
        RECT 55.850 184.265 56.125 184.435 ;
        RECT 56.295 184.265 56.485 185.625 ;
        RECT 56.655 185.640 56.825 186.305 ;
        RECT 56.995 185.885 57.165 186.645 ;
        RECT 57.400 185.885 57.915 186.295 ;
        RECT 56.655 185.450 57.405 185.640 ;
        RECT 57.575 185.075 57.915 185.885 ;
        RECT 58.085 185.555 59.755 186.645 ;
        RECT 56.685 184.905 57.915 185.075 ;
        RECT 56.665 184.095 57.175 184.630 ;
        RECT 57.395 184.300 57.640 184.905 ;
        RECT 58.085 184.865 58.835 185.385 ;
        RECT 59.005 185.035 59.755 185.555 ;
        RECT 59.925 185.505 60.185 186.645 ;
        RECT 60.355 185.495 60.685 186.475 ;
        RECT 60.855 185.505 61.135 186.645 ;
        RECT 59.945 185.085 60.280 185.335 ;
        RECT 60.450 184.895 60.620 185.495 ;
        RECT 62.225 185.480 62.515 186.645 ;
        RECT 62.985 186.005 63.315 186.435 ;
        RECT 62.860 185.835 63.315 186.005 ;
        RECT 63.495 186.005 63.745 186.425 ;
        RECT 63.975 186.175 64.305 186.645 ;
        RECT 64.535 186.005 64.785 186.425 ;
        RECT 63.495 185.835 64.785 186.005 ;
        RECT 60.790 185.065 61.125 185.335 ;
        RECT 58.085 184.095 59.755 184.865 ;
        RECT 59.925 184.265 60.620 184.895 ;
        RECT 60.825 184.095 61.135 184.895 ;
        RECT 62.860 184.835 63.030 185.835 ;
        RECT 63.200 185.005 63.445 185.665 ;
        RECT 63.660 185.005 63.925 185.665 ;
        RECT 64.120 185.005 64.405 185.665 ;
        RECT 64.580 185.335 64.795 185.665 ;
        RECT 64.975 185.505 65.225 186.645 ;
        RECT 65.395 185.585 65.725 186.435 ;
        RECT 64.580 185.005 64.885 185.335 ;
        RECT 65.055 185.005 65.365 185.335 ;
        RECT 65.055 184.835 65.225 185.005 ;
        RECT 62.225 184.095 62.515 184.820 ;
        RECT 62.860 184.665 65.225 184.835 ;
        RECT 65.535 184.820 65.725 185.585 ;
        RECT 65.905 185.555 68.495 186.645 ;
        RECT 63.015 184.095 63.345 184.495 ;
        RECT 63.515 184.325 63.845 184.665 ;
        RECT 64.895 184.095 65.225 184.495 ;
        RECT 65.395 184.310 65.725 184.820 ;
        RECT 65.905 184.865 67.115 185.385 ;
        RECT 67.285 185.035 68.495 185.555 ;
        RECT 69.290 185.680 69.620 186.475 ;
        RECT 69.790 185.860 70.030 186.645 ;
        RECT 70.590 186.055 71.345 186.475 ;
        RECT 70.200 185.885 71.665 186.055 ;
        RECT 70.200 185.680 70.370 185.885 ;
        RECT 69.290 185.505 70.370 185.680 ;
        RECT 69.585 185.455 70.370 185.505 ;
        RECT 69.125 184.985 69.385 185.335 ;
        RECT 65.905 184.095 68.495 184.865 ;
        RECT 69.585 184.815 69.755 185.455 ;
        RECT 70.540 185.285 70.830 185.715 ;
        RECT 69.925 185.085 70.270 185.285 ;
        RECT 70.440 185.085 70.830 185.285 ;
        RECT 71.020 185.295 71.325 185.715 ;
        RECT 71.495 185.635 71.665 185.885 ;
        RECT 71.835 185.805 72.165 186.645 ;
        RECT 72.335 186.055 72.585 186.475 ;
        RECT 72.755 186.225 73.095 186.645 ;
        RECT 72.335 185.885 73.095 186.055 ;
        RECT 71.495 185.465 72.455 185.635 ;
        RECT 72.285 185.295 72.455 185.465 ;
        RECT 71.020 185.085 71.505 185.295 ;
        RECT 71.675 185.085 72.115 185.295 ;
        RECT 72.285 185.085 72.615 185.295 ;
        RECT 72.785 184.915 73.095 185.885 ;
        RECT 69.210 184.645 69.755 184.815 ;
        RECT 70.125 184.745 71.825 184.915 ;
        RECT 70.125 184.655 70.510 184.745 ;
        RECT 69.210 184.265 69.540 184.645 ;
        RECT 69.710 184.305 70.895 184.475 ;
        RECT 71.155 184.095 71.325 184.565 ;
        RECT 71.495 184.280 71.825 184.745 ;
        RECT 71.995 184.095 72.165 184.915 ;
        RECT 72.335 184.745 73.095 184.915 ;
        RECT 73.725 185.805 73.985 186.475 ;
        RECT 74.155 186.245 74.485 186.645 ;
        RECT 75.355 186.245 75.755 186.645 ;
        RECT 76.045 186.065 76.375 186.300 ;
        RECT 74.295 185.895 76.375 186.065 ;
        RECT 73.725 185.795 73.955 185.805 ;
        RECT 73.725 184.835 73.900 185.795 ;
        RECT 74.295 185.625 74.465 185.895 ;
        RECT 74.070 185.455 74.465 185.625 ;
        RECT 74.635 185.505 75.650 185.725 ;
        RECT 74.070 185.005 74.240 185.455 ;
        RECT 75.375 185.365 75.650 185.505 ;
        RECT 75.820 185.505 76.375 185.895 ;
        RECT 74.410 185.085 74.860 185.285 ;
        RECT 75.030 184.915 75.205 185.110 ;
        RECT 72.335 184.275 72.665 184.745 ;
        RECT 72.835 184.095 73.005 184.575 ;
        RECT 73.725 184.265 74.065 184.835 ;
        RECT 74.260 184.095 74.430 184.760 ;
        RECT 74.710 184.745 75.205 184.915 ;
        RECT 74.710 184.605 74.930 184.745 ;
        RECT 74.705 184.435 74.930 184.605 ;
        RECT 75.375 184.575 75.545 185.365 ;
        RECT 75.820 185.255 75.990 185.505 ;
        RECT 76.545 185.335 76.720 186.435 ;
        RECT 76.890 185.825 77.235 186.645 ;
        RECT 75.795 185.085 75.990 185.255 ;
        RECT 76.160 185.085 76.720 185.335 ;
        RECT 76.890 185.085 77.235 185.655 ;
        RECT 77.405 185.505 77.685 186.645 ;
        RECT 77.855 185.495 78.185 186.475 ;
        RECT 78.355 185.505 78.615 186.645 ;
        RECT 79.705 185.885 80.220 186.295 ;
        RECT 80.455 185.885 80.625 186.645 ;
        RECT 80.795 186.305 82.825 186.475 ;
        RECT 77.920 185.455 78.095 185.495 ;
        RECT 75.795 184.700 75.965 185.085 ;
        RECT 77.415 185.065 77.750 185.335 ;
        RECT 74.710 184.390 74.930 184.435 ;
        RECT 75.100 184.405 75.545 184.575 ;
        RECT 75.715 184.330 75.965 184.700 ;
        RECT 76.135 184.735 77.235 184.915 ;
        RECT 77.920 184.895 78.090 185.455 ;
        RECT 78.260 185.085 78.595 185.335 ;
        RECT 79.705 185.075 80.045 185.885 ;
        RECT 80.795 185.640 80.965 186.305 ;
        RECT 81.360 185.965 82.485 186.135 ;
        RECT 80.215 185.450 80.965 185.640 ;
        RECT 81.135 185.625 82.145 185.795 ;
        RECT 79.705 184.905 80.935 185.075 ;
        RECT 76.135 184.330 76.385 184.735 ;
        RECT 76.555 184.095 76.725 184.565 ;
        RECT 76.895 184.330 77.235 184.735 ;
        RECT 77.405 184.095 77.715 184.895 ;
        RECT 77.920 184.265 78.615 184.895 ;
        RECT 79.980 184.300 80.225 184.905 ;
        RECT 80.445 184.095 80.955 184.630 ;
        RECT 81.135 184.265 81.325 185.625 ;
        RECT 81.495 184.605 81.770 185.425 ;
        RECT 81.975 184.825 82.145 185.625 ;
        RECT 82.315 184.835 82.485 185.965 ;
        RECT 82.655 185.335 82.825 186.305 ;
        RECT 82.995 185.505 83.165 186.645 ;
        RECT 83.335 185.505 83.670 186.475 ;
        RECT 82.655 185.005 82.850 185.335 ;
        RECT 83.075 185.005 83.330 185.335 ;
        RECT 83.075 184.835 83.245 185.005 ;
        RECT 83.500 184.835 83.670 185.505 ;
        RECT 82.315 184.665 83.245 184.835 ;
        RECT 82.315 184.630 82.490 184.665 ;
        RECT 81.495 184.435 81.775 184.605 ;
        RECT 81.495 184.265 81.770 184.435 ;
        RECT 81.960 184.265 82.490 184.630 ;
        RECT 82.915 184.095 83.245 184.495 ;
        RECT 83.415 184.265 83.670 184.835 ;
        RECT 83.850 185.505 84.185 186.475 ;
        RECT 84.355 185.505 84.525 186.645 ;
        RECT 84.695 186.305 86.725 186.475 ;
        RECT 83.850 184.835 84.020 185.505 ;
        RECT 84.695 185.335 84.865 186.305 ;
        RECT 84.190 185.005 84.445 185.335 ;
        RECT 84.670 185.005 84.865 185.335 ;
        RECT 85.035 185.965 86.160 186.135 ;
        RECT 84.275 184.835 84.445 185.005 ;
        RECT 85.035 184.835 85.205 185.965 ;
        RECT 83.850 184.265 84.105 184.835 ;
        RECT 84.275 184.665 85.205 184.835 ;
        RECT 85.375 185.625 86.385 185.795 ;
        RECT 85.375 184.825 85.545 185.625 ;
        RECT 85.750 185.285 86.025 185.425 ;
        RECT 85.745 185.115 86.025 185.285 ;
        RECT 85.030 184.630 85.205 184.665 ;
        RECT 84.275 184.095 84.605 184.495 ;
        RECT 85.030 184.265 85.560 184.630 ;
        RECT 85.750 184.265 86.025 185.115 ;
        RECT 86.195 184.265 86.385 185.625 ;
        RECT 86.555 185.640 86.725 186.305 ;
        RECT 86.895 185.885 87.065 186.645 ;
        RECT 87.300 185.885 87.815 186.295 ;
        RECT 86.555 185.450 87.305 185.640 ;
        RECT 87.475 185.075 87.815 185.885 ;
        RECT 87.985 185.480 88.275 186.645 ;
        RECT 88.445 185.555 91.035 186.645 ;
        RECT 86.585 184.905 87.815 185.075 ;
        RECT 86.565 184.095 87.075 184.630 ;
        RECT 87.295 184.300 87.540 184.905 ;
        RECT 88.445 184.865 89.655 185.385 ;
        RECT 89.825 185.035 91.035 185.555 ;
        RECT 91.205 185.040 91.485 186.475 ;
        RECT 91.655 185.870 92.365 186.645 ;
        RECT 92.535 185.700 92.865 186.475 ;
        RECT 91.715 185.485 92.865 185.700 ;
        RECT 87.985 184.095 88.275 184.820 ;
        RECT 88.445 184.095 91.035 184.865 ;
        RECT 91.205 184.265 91.545 185.040 ;
        RECT 91.715 184.915 92.000 185.485 ;
        RECT 92.185 185.085 92.655 185.315 ;
        RECT 93.060 185.285 93.275 186.400 ;
        RECT 93.455 185.925 93.785 186.645 ;
        RECT 94.890 186.255 95.225 186.475 ;
        RECT 96.230 186.265 96.585 186.645 ;
        RECT 94.890 185.635 95.145 186.255 ;
        RECT 95.395 186.095 95.625 186.135 ;
        RECT 96.755 186.095 97.005 186.475 ;
        RECT 95.395 185.895 97.005 186.095 ;
        RECT 95.395 185.805 95.580 185.895 ;
        RECT 96.170 185.885 97.005 185.895 ;
        RECT 97.255 185.865 97.505 186.645 ;
        RECT 97.675 185.795 97.935 186.475 ;
        RECT 95.735 185.695 96.065 185.725 ;
        RECT 95.735 185.635 97.535 185.695 ;
        RECT 93.565 185.285 93.795 185.625 ;
        RECT 94.890 185.525 97.595 185.635 ;
        RECT 94.890 185.465 96.065 185.525 ;
        RECT 97.395 185.490 97.595 185.525 ;
        RECT 92.825 185.105 93.275 185.285 ;
        RECT 92.825 185.085 93.155 185.105 ;
        RECT 93.465 185.085 93.795 185.285 ;
        RECT 94.885 185.085 95.375 185.285 ;
        RECT 95.565 185.085 96.040 185.295 ;
        RECT 91.715 184.725 92.425 184.915 ;
        RECT 92.125 184.585 92.425 184.725 ;
        RECT 92.615 184.725 93.795 184.915 ;
        RECT 92.615 184.645 92.945 184.725 ;
        RECT 92.125 184.575 92.440 184.585 ;
        RECT 92.125 184.565 92.450 184.575 ;
        RECT 92.125 184.560 92.460 184.565 ;
        RECT 91.715 184.095 91.885 184.555 ;
        RECT 92.125 184.550 92.465 184.560 ;
        RECT 92.125 184.545 92.470 184.550 ;
        RECT 92.125 184.535 92.475 184.545 ;
        RECT 92.125 184.530 92.480 184.535 ;
        RECT 92.125 184.265 92.485 184.530 ;
        RECT 93.115 184.095 93.285 184.555 ;
        RECT 93.455 184.265 93.795 184.725 ;
        RECT 94.890 184.095 95.345 184.860 ;
        RECT 95.820 184.685 96.040 185.085 ;
        RECT 96.285 185.085 96.615 185.295 ;
        RECT 96.285 184.685 96.495 185.085 ;
        RECT 96.785 185.050 97.195 185.355 ;
        RECT 97.425 184.915 97.595 185.490 ;
        RECT 97.325 184.795 97.595 184.915 ;
        RECT 96.750 184.750 97.595 184.795 ;
        RECT 96.750 184.625 97.505 184.750 ;
        RECT 96.750 184.475 96.920 184.625 ;
        RECT 97.765 184.595 97.935 185.795 ;
        RECT 98.185 185.715 98.365 186.475 ;
        RECT 98.545 185.885 98.875 186.645 ;
        RECT 98.185 185.545 98.860 185.715 ;
        RECT 99.045 185.570 99.315 186.475 ;
        RECT 98.690 185.400 98.860 185.545 ;
        RECT 98.125 184.995 98.465 185.365 ;
        RECT 98.690 185.070 98.965 185.400 ;
        RECT 98.690 184.815 98.860 185.070 ;
        RECT 95.620 184.265 96.920 184.475 ;
        RECT 97.175 184.095 97.505 184.455 ;
        RECT 97.675 184.265 97.935 184.595 ;
        RECT 98.195 184.645 98.860 184.815 ;
        RECT 99.135 184.770 99.315 185.570 ;
        RECT 99.495 185.505 99.825 186.645 ;
        RECT 100.355 185.675 100.685 186.460 ;
        RECT 100.005 185.505 100.685 185.675 ;
        RECT 100.925 185.505 101.135 186.645 ;
        RECT 99.485 185.085 99.835 185.335 ;
        RECT 100.005 184.905 100.175 185.505 ;
        RECT 101.305 185.495 101.635 186.475 ;
        RECT 101.805 185.505 102.035 186.645 ;
        RECT 102.305 185.505 102.515 186.645 ;
        RECT 102.685 185.495 103.015 186.475 ;
        RECT 103.185 185.505 103.415 186.645 ;
        RECT 103.715 185.715 103.885 186.475 ;
        RECT 104.065 185.885 104.395 186.645 ;
        RECT 103.715 185.545 104.380 185.715 ;
        RECT 104.565 185.570 104.835 186.475 ;
        RECT 100.345 185.085 100.695 185.335 ;
        RECT 98.195 184.265 98.365 184.645 ;
        RECT 98.545 184.095 98.875 184.475 ;
        RECT 99.055 184.265 99.315 184.770 ;
        RECT 99.495 184.095 99.765 184.905 ;
        RECT 99.935 184.265 100.265 184.905 ;
        RECT 100.435 184.095 100.675 184.905 ;
        RECT 100.925 184.095 101.135 184.915 ;
        RECT 101.305 184.895 101.555 185.495 ;
        RECT 101.725 185.085 102.055 185.335 ;
        RECT 101.305 184.265 101.635 184.895 ;
        RECT 101.805 184.095 102.035 184.915 ;
        RECT 102.305 184.095 102.515 184.915 ;
        RECT 102.685 184.895 102.935 185.495 ;
        RECT 104.210 185.400 104.380 185.545 ;
        RECT 103.105 185.085 103.435 185.335 ;
        RECT 103.645 184.995 103.975 185.365 ;
        RECT 104.210 185.070 104.495 185.400 ;
        RECT 102.685 184.265 103.015 184.895 ;
        RECT 103.185 184.095 103.415 184.915 ;
        RECT 104.210 184.815 104.380 185.070 ;
        RECT 103.715 184.645 104.380 184.815 ;
        RECT 104.665 184.770 104.835 185.570 ;
        RECT 103.715 184.265 103.885 184.645 ;
        RECT 104.065 184.095 104.395 184.475 ;
        RECT 104.575 184.265 104.835 184.770 ;
        RECT 105.005 185.570 105.275 186.475 ;
        RECT 105.445 185.885 105.775 186.645 ;
        RECT 105.955 185.715 106.135 186.475 ;
        RECT 105.005 184.770 105.185 185.570 ;
        RECT 105.460 185.545 106.135 185.715 ;
        RECT 106.385 185.570 106.655 186.475 ;
        RECT 106.825 185.885 107.155 186.645 ;
        RECT 107.335 185.715 107.515 186.475 ;
        RECT 105.460 185.400 105.630 185.545 ;
        RECT 105.355 185.070 105.630 185.400 ;
        RECT 105.460 184.815 105.630 185.070 ;
        RECT 105.855 184.995 106.195 185.365 ;
        RECT 105.005 184.265 105.265 184.770 ;
        RECT 105.460 184.645 106.125 184.815 ;
        RECT 105.445 184.095 105.775 184.475 ;
        RECT 105.955 184.265 106.125 184.645 ;
        RECT 106.385 184.770 106.565 185.570 ;
        RECT 106.840 185.545 107.515 185.715 ;
        RECT 107.950 185.675 108.340 185.850 ;
        RECT 108.825 185.845 109.155 186.645 ;
        RECT 109.325 185.855 109.860 186.475 ;
        RECT 106.840 185.400 107.010 185.545 ;
        RECT 107.950 185.505 109.375 185.675 ;
        RECT 106.735 185.070 107.010 185.400 ;
        RECT 106.840 184.815 107.010 185.070 ;
        RECT 107.235 184.995 107.575 185.365 ;
        RECT 106.385 184.265 106.645 184.770 ;
        RECT 106.840 184.645 107.505 184.815 ;
        RECT 107.825 184.775 108.180 185.335 ;
        RECT 106.825 184.095 107.155 184.475 ;
        RECT 107.335 184.265 107.505 184.645 ;
        RECT 108.350 184.605 108.520 185.505 ;
        RECT 108.690 184.775 108.955 185.335 ;
        RECT 109.205 185.005 109.375 185.505 ;
        RECT 109.545 184.835 109.860 185.855 ;
        RECT 110.070 185.500 110.365 186.645 ;
        RECT 107.930 184.095 108.170 184.605 ;
        RECT 108.350 184.275 108.630 184.605 ;
        RECT 108.860 184.095 109.075 184.605 ;
        RECT 109.245 184.265 109.860 184.835 ;
        RECT 110.070 184.095 110.365 184.915 ;
        RECT 110.535 184.645 110.765 186.345 ;
        RECT 110.980 185.840 111.235 186.645 ;
        RECT 111.435 186.030 111.765 186.475 ;
        RECT 111.935 186.200 112.210 186.645 ;
        RECT 112.445 186.030 112.775 186.475 ;
        RECT 111.435 185.850 112.775 186.030 ;
        RECT 113.235 185.670 113.565 186.335 ;
        RECT 110.980 185.500 113.565 185.670 ;
        RECT 110.980 184.885 111.290 185.500 ;
        RECT 113.745 185.480 114.035 186.645 ;
        RECT 114.210 185.775 114.475 186.475 ;
        RECT 114.645 185.945 114.975 186.645 ;
        RECT 115.145 185.775 115.815 186.475 ;
        RECT 116.320 185.945 116.750 186.645 ;
        RECT 116.930 186.085 117.120 186.475 ;
        RECT 117.290 186.265 117.620 186.645 ;
        RECT 116.930 185.915 117.660 186.085 ;
        RECT 114.210 185.520 116.785 185.775 ;
        RECT 111.460 185.055 111.790 185.285 ;
        RECT 111.960 185.055 112.430 185.285 ;
        RECT 112.600 185.115 113.055 185.285 ;
        RECT 112.600 185.055 113.050 185.115 ;
        RECT 113.240 185.055 113.575 185.285 ;
        RECT 114.205 185.005 114.480 185.335 ;
        RECT 110.980 184.705 113.565 184.885 ;
        RECT 114.650 184.835 114.830 185.520 ;
        RECT 116.615 185.335 116.785 185.520 ;
        RECT 115.000 185.005 115.360 185.335 ;
        RECT 115.650 185.285 115.940 185.335 ;
        RECT 115.645 185.115 115.940 185.285 ;
        RECT 115.650 185.005 115.940 185.115 ;
        RECT 116.110 185.005 116.445 185.335 ;
        RECT 116.615 185.005 117.295 185.335 ;
        RECT 110.535 184.265 110.755 184.645 ;
        RECT 110.925 184.095 111.775 184.455 ;
        RECT 112.255 184.285 112.585 184.705 ;
        RECT 112.790 184.095 113.065 184.535 ;
        RECT 113.235 184.285 113.565 184.705 ;
        RECT 113.745 184.095 114.035 184.820 ;
        RECT 114.215 184.435 114.830 184.835 ;
        RECT 115.000 184.645 116.270 184.835 ;
        RECT 117.465 184.795 117.660 185.915 ;
        RECT 116.840 184.625 117.660 184.795 ;
        RECT 117.885 185.570 118.155 186.475 ;
        RECT 118.325 185.885 118.655 186.645 ;
        RECT 118.835 185.715 119.005 186.475 ;
        RECT 119.355 185.900 119.625 186.645 ;
        RECT 120.255 186.640 126.530 186.645 ;
        RECT 119.795 185.730 120.085 186.470 ;
        RECT 120.255 185.915 120.510 186.640 ;
        RECT 120.695 185.745 120.955 186.470 ;
        RECT 121.125 185.915 121.370 186.640 ;
        RECT 121.555 185.745 121.815 186.470 ;
        RECT 121.985 185.915 122.230 186.640 ;
        RECT 122.415 185.745 122.675 186.470 ;
        RECT 122.845 185.915 123.090 186.640 ;
        RECT 123.260 185.745 123.520 186.470 ;
        RECT 123.690 185.915 123.950 186.640 ;
        RECT 124.120 185.745 124.380 186.470 ;
        RECT 124.550 185.915 124.810 186.640 ;
        RECT 124.980 185.745 125.240 186.470 ;
        RECT 125.410 185.915 125.670 186.640 ;
        RECT 125.840 185.745 126.100 186.470 ;
        RECT 126.270 185.845 126.530 186.640 ;
        RECT 120.695 185.730 126.100 185.745 ;
        RECT 117.885 184.770 118.055 185.570 ;
        RECT 118.340 185.545 119.005 185.715 ;
        RECT 118.340 185.400 118.510 185.545 ;
        RECT 118.225 185.070 118.510 185.400 ;
        RECT 119.355 185.505 126.100 185.730 ;
        RECT 118.340 184.815 118.510 185.070 ;
        RECT 118.745 184.995 119.075 185.365 ;
        RECT 119.355 184.915 120.520 185.505 ;
        RECT 126.700 185.335 126.950 186.470 ;
        RECT 127.130 185.835 127.390 186.645 ;
        RECT 127.565 185.335 127.810 186.475 ;
        RECT 127.990 185.835 128.285 186.645 ;
        RECT 129.600 185.545 129.930 186.645 ;
        RECT 130.405 186.045 130.730 186.475 ;
        RECT 130.900 186.225 131.230 186.645 ;
        RECT 131.975 186.215 132.385 186.645 ;
        RECT 130.405 185.875 132.385 186.045 ;
        RECT 130.405 185.465 131.110 185.875 ;
        RECT 120.690 185.085 127.810 185.335 ;
        RECT 114.215 184.265 114.550 184.435 ;
        RECT 115.510 184.095 115.845 184.475 ;
        RECT 116.435 184.095 116.670 184.535 ;
        RECT 116.840 184.265 117.170 184.625 ;
        RECT 117.340 184.095 117.670 184.455 ;
        RECT 117.885 184.265 118.145 184.770 ;
        RECT 118.340 184.645 119.005 184.815 ;
        RECT 119.355 184.745 126.100 184.915 ;
        RECT 118.325 184.095 118.655 184.475 ;
        RECT 118.835 184.265 119.005 184.645 ;
        RECT 119.355 184.095 119.655 184.575 ;
        RECT 119.825 184.290 120.085 184.745 ;
        RECT 120.255 184.095 120.515 184.575 ;
        RECT 120.695 184.290 120.955 184.745 ;
        RECT 121.125 184.095 121.375 184.575 ;
        RECT 121.555 184.290 121.815 184.745 ;
        RECT 121.985 184.095 122.235 184.575 ;
        RECT 122.415 184.290 122.675 184.745 ;
        RECT 122.845 184.095 123.090 184.575 ;
        RECT 123.260 184.290 123.535 184.745 ;
        RECT 123.705 184.095 123.950 184.575 ;
        RECT 124.120 184.290 124.380 184.745 ;
        RECT 124.550 184.095 124.810 184.575 ;
        RECT 124.980 184.290 125.240 184.745 ;
        RECT 125.410 184.095 125.670 184.575 ;
        RECT 125.840 184.290 126.100 184.745 ;
        RECT 126.270 184.095 126.530 184.655 ;
        RECT 126.700 184.275 126.950 185.085 ;
        RECT 127.130 184.095 127.390 184.620 ;
        RECT 127.560 184.275 127.810 185.085 ;
        RECT 127.980 184.775 128.295 185.335 ;
        RECT 129.385 185.085 130.030 185.295 ;
        RECT 130.200 185.085 130.770 185.295 ;
        RECT 129.540 184.745 130.710 184.915 ;
        RECT 127.990 184.095 128.295 184.605 ;
        RECT 129.540 184.280 129.870 184.745 ;
        RECT 130.040 184.095 130.210 184.565 ;
        RECT 130.380 184.265 130.710 184.745 ;
        RECT 130.940 184.265 131.110 185.465 ;
        RECT 131.280 185.535 131.905 185.705 ;
        RECT 131.280 184.835 131.450 185.535 ;
        RECT 132.120 185.335 132.385 185.875 ;
        RECT 132.555 185.490 132.895 186.475 ;
        RECT 133.145 185.715 133.325 186.475 ;
        RECT 133.505 185.885 133.835 186.645 ;
        RECT 133.145 185.545 133.820 185.715 ;
        RECT 134.005 185.570 134.275 186.475 ;
        RECT 131.620 185.005 131.950 185.335 ;
        RECT 132.120 185.005 132.470 185.335 ;
        RECT 132.640 184.835 132.895 185.490 ;
        RECT 133.650 185.400 133.820 185.545 ;
        RECT 133.085 184.995 133.425 185.365 ;
        RECT 133.650 185.070 133.925 185.400 ;
        RECT 131.280 184.665 131.820 184.835 ;
        RECT 131.650 184.460 131.820 184.665 ;
        RECT 132.100 184.095 132.270 184.835 ;
        RECT 132.535 184.460 132.895 184.835 ;
        RECT 133.650 184.815 133.820 185.070 ;
        RECT 133.155 184.645 133.820 184.815 ;
        RECT 134.095 184.770 134.275 185.570 ;
        RECT 134.905 185.555 136.115 186.645 ;
        RECT 134.905 185.015 135.425 185.555 ;
        RECT 135.595 184.845 136.115 185.385 ;
        RECT 132.665 184.435 132.835 184.460 ;
        RECT 133.155 184.265 133.325 184.645 ;
        RECT 133.505 184.095 133.835 184.475 ;
        RECT 134.015 184.265 134.275 184.770 ;
        RECT 134.905 184.095 136.115 184.845 ;
        RECT 23.500 183.925 136.200 184.095 ;
        RECT 23.585 183.175 24.795 183.925 ;
        RECT 24.965 183.380 30.310 183.925 ;
        RECT 23.585 182.635 24.105 183.175 ;
        RECT 24.275 182.465 24.795 183.005 ;
        RECT 26.550 182.550 26.890 183.380 ;
        RECT 30.485 183.155 33.995 183.925 ;
        RECT 35.090 183.185 35.345 183.755 ;
        RECT 35.515 183.525 35.845 183.925 ;
        RECT 36.270 183.390 36.800 183.755 ;
        RECT 36.990 183.585 37.265 183.755 ;
        RECT 36.985 183.415 37.265 183.585 ;
        RECT 36.270 183.355 36.445 183.390 ;
        RECT 35.515 183.185 36.445 183.355 ;
        RECT 23.585 181.375 24.795 182.465 ;
        RECT 28.370 181.810 28.720 183.060 ;
        RECT 30.485 182.635 32.135 183.155 ;
        RECT 32.305 182.465 33.995 182.985 ;
        RECT 24.965 181.375 30.310 181.810 ;
        RECT 30.485 181.375 33.995 182.465 ;
        RECT 35.090 182.515 35.260 183.185 ;
        RECT 35.515 183.015 35.685 183.185 ;
        RECT 35.430 182.685 35.685 183.015 ;
        RECT 35.910 182.685 36.105 183.015 ;
        RECT 35.090 181.545 35.425 182.515 ;
        RECT 35.595 181.375 35.765 182.515 ;
        RECT 35.935 181.715 36.105 182.685 ;
        RECT 36.275 182.055 36.445 183.185 ;
        RECT 36.615 182.395 36.785 183.195 ;
        RECT 36.990 182.595 37.265 183.415 ;
        RECT 37.435 182.395 37.625 183.755 ;
        RECT 37.805 183.390 38.315 183.925 ;
        RECT 38.535 183.115 38.780 183.720 ;
        RECT 39.270 183.465 40.020 183.755 ;
        RECT 40.530 183.465 40.860 183.925 ;
        RECT 37.825 182.945 39.055 183.115 ;
        RECT 36.615 182.225 37.625 182.395 ;
        RECT 37.795 182.380 38.545 182.570 ;
        RECT 36.275 181.885 37.400 182.055 ;
        RECT 37.795 181.715 37.965 182.380 ;
        RECT 38.715 182.135 39.055 182.945 ;
        RECT 35.935 181.545 37.965 181.715 ;
        RECT 38.135 181.375 38.305 182.135 ;
        RECT 38.540 181.725 39.055 182.135 ;
        RECT 39.270 182.175 39.640 183.465 ;
        RECT 41.080 183.275 41.350 183.485 ;
        RECT 40.015 183.105 41.350 183.275 ;
        RECT 41.585 183.105 41.795 183.925 ;
        RECT 41.965 183.125 42.295 183.755 ;
        RECT 40.015 182.935 40.185 183.105 ;
        RECT 39.810 182.685 40.185 182.935 ;
        RECT 40.355 182.695 40.830 182.935 ;
        RECT 41.000 182.695 41.350 182.935 ;
        RECT 40.015 182.515 40.185 182.685 ;
        RECT 41.965 182.525 42.215 183.125 ;
        RECT 42.465 183.105 42.695 183.925 ;
        RECT 42.905 183.155 46.415 183.925 ;
        RECT 42.385 182.685 42.715 182.935 ;
        RECT 42.905 182.635 44.555 183.155 ;
        RECT 47.545 183.105 47.775 183.925 ;
        RECT 47.945 183.125 48.275 183.755 ;
        RECT 40.015 182.345 41.350 182.515 ;
        RECT 41.070 182.185 41.350 182.345 ;
        RECT 39.270 182.005 40.440 182.175 ;
        RECT 39.725 181.375 39.940 181.835 ;
        RECT 40.110 181.545 40.440 182.005 ;
        RECT 40.610 181.375 40.860 182.175 ;
        RECT 41.585 181.375 41.795 182.515 ;
        RECT 41.965 181.545 42.295 182.525 ;
        RECT 42.465 181.375 42.695 182.515 ;
        RECT 44.725 182.465 46.415 182.985 ;
        RECT 47.525 182.685 47.855 182.935 ;
        RECT 48.025 182.525 48.275 183.125 ;
        RECT 48.445 183.105 48.655 183.925 ;
        RECT 49.345 183.200 49.635 183.925 ;
        RECT 50.265 183.125 50.960 183.755 ;
        RECT 51.165 183.125 51.475 183.925 ;
        RECT 51.645 183.380 56.990 183.925 ;
        RECT 50.285 182.685 50.620 182.935 ;
        RECT 42.905 181.375 46.415 182.465 ;
        RECT 47.545 181.375 47.775 182.515 ;
        RECT 47.945 181.545 48.275 182.525 ;
        RECT 48.445 181.375 48.655 182.515 ;
        RECT 49.345 181.375 49.635 182.540 ;
        RECT 50.790 182.525 50.960 183.125 ;
        RECT 51.130 182.685 51.465 182.955 ;
        RECT 53.230 182.550 53.570 183.380 ;
        RECT 57.165 183.155 60.675 183.925 ;
        RECT 60.845 183.175 62.055 183.925 ;
        RECT 62.310 183.425 62.805 183.755 ;
        RECT 50.265 181.375 50.525 182.515 ;
        RECT 50.695 181.545 51.025 182.525 ;
        RECT 51.195 181.375 51.475 182.515 ;
        RECT 55.050 181.810 55.400 183.060 ;
        RECT 57.165 182.635 58.815 183.155 ;
        RECT 58.985 182.465 60.675 182.985 ;
        RECT 60.845 182.635 61.365 183.175 ;
        RECT 61.535 182.465 62.055 183.005 ;
        RECT 51.645 181.375 56.990 181.810 ;
        RECT 57.165 181.375 60.675 182.465 ;
        RECT 60.845 181.375 62.055 182.465 ;
        RECT 62.225 181.935 62.465 183.245 ;
        RECT 62.635 182.515 62.805 183.425 ;
        RECT 63.025 182.685 63.375 183.650 ;
        RECT 63.555 182.685 63.855 183.655 ;
        RECT 64.035 182.685 64.315 183.655 ;
        RECT 64.495 183.125 64.765 183.925 ;
        RECT 64.935 183.205 65.275 183.715 ;
        RECT 64.510 182.685 64.840 182.935 ;
        RECT 64.510 182.515 64.825 182.685 ;
        RECT 62.635 182.345 64.825 182.515 ;
        RECT 62.230 181.375 62.565 181.755 ;
        RECT 62.735 181.545 62.985 182.345 ;
        RECT 63.205 181.375 63.535 182.095 ;
        RECT 63.720 181.545 63.970 182.345 ;
        RECT 64.435 181.375 64.765 182.175 ;
        RECT 65.015 181.805 65.275 183.205 ;
        RECT 65.455 183.395 65.785 183.755 ;
        RECT 65.955 183.565 66.285 183.925 ;
        RECT 66.485 183.395 66.815 183.755 ;
        RECT 65.455 183.185 66.815 183.395 ;
        RECT 67.325 183.165 68.035 183.755 ;
        RECT 68.205 183.380 73.550 183.925 ;
        RECT 65.445 182.685 65.755 183.015 ;
        RECT 65.965 182.685 66.340 183.015 ;
        RECT 66.660 182.685 67.155 183.015 ;
        RECT 64.935 181.545 65.275 181.805 ;
        RECT 65.455 181.375 65.785 182.435 ;
        RECT 65.965 181.715 66.135 182.685 ;
        RECT 66.305 182.195 66.635 182.415 ;
        RECT 66.830 182.395 67.155 182.685 ;
        RECT 67.330 182.395 67.660 182.935 ;
        RECT 67.830 182.195 68.035 183.165 ;
        RECT 69.790 182.550 70.130 183.380 ;
        RECT 73.725 183.175 74.935 183.925 ;
        RECT 75.105 183.200 75.395 183.925 ;
        RECT 66.305 181.965 68.035 182.195 ;
        RECT 66.305 181.565 66.635 181.965 ;
        RECT 66.805 181.375 67.135 181.735 ;
        RECT 67.335 181.545 68.035 181.965 ;
        RECT 71.610 181.810 71.960 183.060 ;
        RECT 73.725 182.635 74.245 183.175 ;
        RECT 75.565 183.125 75.875 183.925 ;
        RECT 76.080 183.125 76.775 183.755 ;
        RECT 77.410 183.395 77.700 183.745 ;
        RECT 77.895 183.565 78.225 183.925 ;
        RECT 78.395 183.395 78.625 183.700 ;
        RECT 77.410 183.225 78.625 183.395 ;
        RECT 78.815 183.585 78.985 183.620 ;
        RECT 78.815 183.415 79.015 183.585 ;
        RECT 74.415 182.465 74.935 183.005 ;
        RECT 75.575 182.685 75.910 182.955 ;
        RECT 68.205 181.375 73.550 181.810 ;
        RECT 73.725 181.375 74.935 182.465 ;
        RECT 75.105 181.375 75.395 182.540 ;
        RECT 76.080 182.525 76.250 183.125 ;
        RECT 78.815 183.055 78.985 183.415 ;
        RECT 76.420 182.685 76.755 182.935 ;
        RECT 77.470 182.905 77.730 183.015 ;
        RECT 77.465 182.735 77.730 182.905 ;
        RECT 77.470 182.685 77.730 182.735 ;
        RECT 77.910 182.685 78.295 183.015 ;
        RECT 78.465 182.885 78.985 183.055 ;
        RECT 79.245 183.155 80.915 183.925 ;
        RECT 75.565 181.375 75.845 182.515 ;
        RECT 76.015 181.545 76.345 182.525 ;
        RECT 76.515 181.375 76.775 182.515 ;
        RECT 77.410 181.375 77.730 182.515 ;
        RECT 77.910 181.635 78.105 182.685 ;
        RECT 78.465 182.505 78.635 182.885 ;
        RECT 78.285 182.225 78.635 182.505 ;
        RECT 78.825 182.355 79.070 182.715 ;
        RECT 79.245 182.635 79.995 183.155 ;
        RECT 81.085 183.125 81.395 183.925 ;
        RECT 81.600 183.125 82.295 183.755 ;
        RECT 82.465 183.380 87.810 183.925 ;
        RECT 88.450 183.450 88.785 183.710 ;
        RECT 88.955 183.525 89.285 183.925 ;
        RECT 89.455 183.525 91.070 183.695 ;
        RECT 80.165 182.465 80.915 182.985 ;
        RECT 81.095 182.685 81.430 182.955 ;
        RECT 81.600 182.525 81.770 183.125 ;
        RECT 81.940 182.685 82.275 182.935 ;
        RECT 84.050 182.550 84.390 183.380 ;
        RECT 78.285 181.545 78.615 182.225 ;
        RECT 78.815 181.375 79.070 182.175 ;
        RECT 79.245 181.375 80.915 182.465 ;
        RECT 81.085 181.375 81.365 182.515 ;
        RECT 81.535 181.545 81.865 182.525 ;
        RECT 82.035 181.375 82.295 182.515 ;
        RECT 85.870 181.810 86.220 183.060 ;
        RECT 88.450 182.095 88.705 183.450 ;
        RECT 89.455 183.355 89.625 183.525 ;
        RECT 89.065 183.185 89.625 183.355 ;
        RECT 89.065 183.015 89.235 183.185 ;
        RECT 88.930 182.685 89.235 183.015 ;
        RECT 89.430 182.905 89.680 183.015 ;
        RECT 89.890 182.905 90.160 183.345 ;
        RECT 90.350 182.905 90.640 183.345 ;
        RECT 89.425 182.735 89.680 182.905 ;
        RECT 89.885 182.735 90.160 182.905 ;
        RECT 90.345 182.735 90.640 182.905 ;
        RECT 89.430 182.685 89.680 182.735 ;
        RECT 89.890 182.685 90.160 182.735 ;
        RECT 90.350 182.685 90.640 182.735 ;
        RECT 90.810 182.685 91.230 183.350 ;
        RECT 91.615 183.205 91.945 183.925 ;
        RECT 91.540 182.905 91.890 183.015 ;
        RECT 91.540 182.735 91.895 182.905 ;
        RECT 91.540 182.685 91.890 182.735 ;
        RECT 89.065 182.515 89.235 182.685 ;
        RECT 89.065 182.345 91.435 182.515 ;
        RECT 91.685 182.395 91.890 182.685 ;
        RECT 82.465 181.375 87.810 181.810 ;
        RECT 88.450 181.585 88.785 182.095 ;
        RECT 89.035 181.375 89.365 182.175 ;
        RECT 89.610 181.965 91.035 182.135 ;
        RECT 89.610 181.545 89.895 181.965 ;
        RECT 90.150 181.375 90.480 181.795 ;
        RECT 90.705 181.715 91.035 181.965 ;
        RECT 91.265 181.885 91.435 182.345 ;
        RECT 91.695 181.715 91.865 182.215 ;
        RECT 90.705 181.545 91.865 181.715 ;
        RECT 92.125 181.545 92.875 183.755 ;
        RECT 93.135 183.375 93.305 183.755 ;
        RECT 93.485 183.545 93.815 183.925 ;
        RECT 93.135 183.205 93.800 183.375 ;
        RECT 93.995 183.250 94.255 183.755 ;
        RECT 93.065 182.655 93.405 183.025 ;
        RECT 93.630 182.950 93.800 183.205 ;
        RECT 93.630 182.620 93.905 182.950 ;
        RECT 93.630 182.475 93.800 182.620 ;
        RECT 93.125 182.305 93.800 182.475 ;
        RECT 94.075 182.450 94.255 183.250 ;
        RECT 94.585 183.365 94.915 183.755 ;
        RECT 95.085 183.535 96.270 183.705 ;
        RECT 96.530 183.455 96.700 183.925 ;
        RECT 94.585 183.185 95.095 183.365 ;
        RECT 94.425 182.725 94.755 183.015 ;
        RECT 94.925 182.555 95.095 183.185 ;
        RECT 95.500 183.275 95.885 183.365 ;
        RECT 96.870 183.275 97.200 183.740 ;
        RECT 95.500 183.105 97.200 183.275 ;
        RECT 97.370 183.105 97.540 183.925 ;
        RECT 97.710 183.105 98.395 183.745 ;
        RECT 99.495 183.115 99.765 183.925 ;
        RECT 99.935 183.115 100.265 183.755 ;
        RECT 100.435 183.115 100.675 183.925 ;
        RECT 100.865 183.200 101.155 183.925 ;
        RECT 101.415 183.375 101.585 183.755 ;
        RECT 101.765 183.545 102.095 183.925 ;
        RECT 101.415 183.205 102.080 183.375 ;
        RECT 102.275 183.250 102.535 183.755 ;
        RECT 95.265 182.725 95.595 182.935 ;
        RECT 95.775 182.685 96.155 182.935 ;
        RECT 93.125 181.545 93.305 182.305 ;
        RECT 93.485 181.375 93.815 182.135 ;
        RECT 93.985 181.545 94.255 182.450 ;
        RECT 94.580 182.385 95.665 182.555 ;
        RECT 94.580 181.545 94.880 182.385 ;
        RECT 95.075 181.375 95.325 182.215 ;
        RECT 95.495 182.135 95.665 182.385 ;
        RECT 95.835 182.305 96.155 182.685 ;
        RECT 96.345 182.725 96.830 182.935 ;
        RECT 97.020 182.725 97.470 182.935 ;
        RECT 97.640 182.725 97.975 182.935 ;
        RECT 96.345 182.565 96.720 182.725 ;
        RECT 96.325 182.395 96.720 182.565 ;
        RECT 97.640 182.555 97.810 182.725 ;
        RECT 96.345 182.305 96.720 182.395 ;
        RECT 96.890 182.385 97.810 182.555 ;
        RECT 96.890 182.135 97.060 182.385 ;
        RECT 95.495 181.965 97.060 182.135 ;
        RECT 95.915 181.545 96.720 181.965 ;
        RECT 97.230 181.375 97.560 182.215 ;
        RECT 98.145 182.135 98.395 183.105 ;
        RECT 99.485 182.685 99.835 182.935 ;
        RECT 100.005 182.515 100.175 183.115 ;
        RECT 100.345 182.685 100.695 182.935 ;
        RECT 101.345 182.655 101.685 183.025 ;
        RECT 101.910 182.950 102.080 183.205 ;
        RECT 101.910 182.620 102.185 182.950 ;
        RECT 97.730 181.545 98.395 182.135 ;
        RECT 99.495 181.375 99.825 182.515 ;
        RECT 100.005 182.345 100.685 182.515 ;
        RECT 100.355 181.560 100.685 182.345 ;
        RECT 100.865 181.375 101.155 182.540 ;
        RECT 101.910 182.475 102.080 182.620 ;
        RECT 101.405 182.305 102.080 182.475 ;
        RECT 102.355 182.450 102.535 183.250 ;
        RECT 102.705 183.125 103.400 183.755 ;
        RECT 103.605 183.125 103.915 183.925 ;
        RECT 104.085 183.125 104.780 183.755 ;
        RECT 104.985 183.125 105.295 183.925 ;
        RECT 105.470 183.160 105.925 183.925 ;
        RECT 106.200 183.545 107.500 183.755 ;
        RECT 107.755 183.565 108.085 183.925 ;
        RECT 107.330 183.395 107.500 183.545 ;
        RECT 108.255 183.425 108.515 183.755 ;
        RECT 108.685 183.445 108.945 183.925 ;
        RECT 109.115 183.675 109.360 183.755 ;
        RECT 109.115 183.505 109.445 183.675 ;
        RECT 102.725 182.685 103.060 182.935 ;
        RECT 103.230 182.525 103.400 183.125 ;
        RECT 103.570 182.685 103.905 182.955 ;
        RECT 104.105 182.685 104.440 182.935 ;
        RECT 104.610 182.525 104.780 183.125 ;
        RECT 104.950 182.685 105.285 182.955 ;
        RECT 106.400 182.935 106.620 183.335 ;
        RECT 105.465 182.735 105.955 182.935 ;
        RECT 106.145 182.725 106.620 182.935 ;
        RECT 106.865 182.935 107.075 183.335 ;
        RECT 107.330 183.270 108.085 183.395 ;
        RECT 107.330 183.225 108.175 183.270 ;
        RECT 107.905 183.105 108.175 183.225 ;
        RECT 106.865 182.725 107.195 182.935 ;
        RECT 107.365 182.665 107.775 182.970 ;
        RECT 101.405 181.545 101.585 182.305 ;
        RECT 101.765 181.375 102.095 182.135 ;
        RECT 102.265 181.545 102.535 182.450 ;
        RECT 102.705 181.375 102.965 182.515 ;
        RECT 103.135 181.545 103.465 182.525 ;
        RECT 103.635 181.375 103.915 182.515 ;
        RECT 104.085 181.375 104.345 182.515 ;
        RECT 104.515 181.545 104.845 182.525 ;
        RECT 105.015 181.375 105.295 182.515 ;
        RECT 105.470 182.495 106.645 182.555 ;
        RECT 108.005 182.530 108.175 183.105 ;
        RECT 107.975 182.495 108.175 182.530 ;
        RECT 105.470 182.385 108.175 182.495 ;
        RECT 105.470 181.765 105.725 182.385 ;
        RECT 106.315 182.325 108.115 182.385 ;
        RECT 106.315 182.295 106.645 182.325 ;
        RECT 108.345 182.225 108.515 183.425 ;
        RECT 108.730 182.685 108.925 183.255 ;
        RECT 109.115 182.515 109.285 183.505 ;
        RECT 109.645 183.310 109.855 183.595 ;
        RECT 110.120 183.585 110.290 183.610 ;
        RECT 110.120 183.415 110.295 183.585 ;
        RECT 110.535 183.545 110.865 183.925 ;
        RECT 110.635 183.465 110.805 183.545 ;
        RECT 110.120 183.315 110.290 183.415 ;
        RECT 109.465 183.140 109.855 183.310 ;
        RECT 110.025 183.145 110.290 183.315 ;
        RECT 111.055 183.295 111.225 183.755 ;
        RECT 111.475 183.465 111.730 183.925 ;
        RECT 109.465 183.075 109.745 183.140 ;
        RECT 109.465 182.685 109.635 183.075 ;
        RECT 110.025 182.935 110.195 183.145 ;
        RECT 110.550 183.015 110.755 183.250 ;
        RECT 111.055 183.125 111.730 183.295 ;
        RECT 111.915 183.185 112.245 183.925 ;
        RECT 112.425 183.395 112.745 183.755 ;
        RECT 112.950 183.565 113.280 183.925 ;
        RECT 113.740 183.395 114.085 183.755 ;
        RECT 112.425 183.225 114.085 183.395 ;
        RECT 109.865 182.765 110.195 182.935 ;
        RECT 110.025 182.750 110.195 182.765 ;
        RECT 110.425 182.685 110.755 183.015 ;
        RECT 110.935 182.765 111.265 182.935 ;
        RECT 111.095 182.515 111.265 182.765 ;
        RECT 105.975 182.125 106.160 182.215 ;
        RECT 106.750 182.125 107.585 182.135 ;
        RECT 105.975 181.925 107.585 182.125 ;
        RECT 105.975 181.885 106.205 181.925 ;
        RECT 105.470 181.545 105.805 181.765 ;
        RECT 106.810 181.375 107.165 181.755 ;
        RECT 107.335 181.545 107.585 181.925 ;
        RECT 107.835 181.375 108.085 182.155 ;
        RECT 108.255 181.545 108.515 182.225 ;
        RECT 108.775 182.345 111.265 182.515 ;
        RECT 108.775 181.545 108.945 182.345 ;
        RECT 111.475 182.175 111.730 183.125 ;
        RECT 111.965 182.385 112.240 183.015 ;
        RECT 109.175 182.005 110.465 182.175 ;
        RECT 109.235 181.585 109.485 182.005 ;
        RECT 109.675 181.375 110.005 181.835 ;
        RECT 110.215 181.585 110.465 182.005 ;
        RECT 110.635 181.375 110.885 182.175 ;
        RECT 111.055 182.005 111.730 182.175 ;
        RECT 111.055 181.545 111.225 182.005 ;
        RECT 111.435 181.375 111.685 181.835 ;
        RECT 111.950 181.725 112.255 182.215 ;
        RECT 112.425 181.895 112.725 183.225 ;
        RECT 114.645 183.145 114.940 183.925 ;
        RECT 115.125 183.185 115.440 183.560 ;
        RECT 115.695 183.185 115.865 183.925 ;
        RECT 116.115 183.355 116.285 183.560 ;
        RECT 116.555 183.530 116.885 183.925 ;
        RECT 117.135 183.355 117.305 183.705 ;
        RECT 117.505 183.525 117.835 183.925 ;
        RECT 118.005 183.355 118.175 183.705 ;
        RECT 118.395 183.525 118.775 183.925 ;
        RECT 116.115 183.185 116.635 183.355 ;
        RECT 113.105 182.765 113.435 182.935 ;
        RECT 113.110 182.515 113.435 182.765 ;
        RECT 113.615 182.685 114.225 183.015 ;
        RECT 114.395 182.515 114.895 182.975 ;
        RECT 113.110 182.335 114.895 182.515 ;
        RECT 112.895 181.985 114.930 182.155 ;
        RECT 112.895 181.725 113.225 181.985 ;
        RECT 113.820 181.905 114.930 181.985 ;
        RECT 111.950 181.545 113.225 181.725 ;
        RECT 113.395 181.375 113.565 181.815 ;
        RECT 113.820 181.545 113.990 181.905 ;
        RECT 114.170 181.375 114.500 181.735 ;
        RECT 114.670 181.545 114.930 181.905 ;
        RECT 115.125 182.145 115.295 183.185 ;
        RECT 116.445 183.015 116.635 183.185 ;
        RECT 116.975 183.185 118.785 183.355 ;
        RECT 115.465 182.315 115.815 183.015 ;
        RECT 115.985 182.685 116.275 183.015 ;
        RECT 116.445 182.685 116.735 183.015 ;
        RECT 116.445 182.485 116.635 182.685 ;
        RECT 116.030 182.315 116.635 182.485 ;
        RECT 115.125 181.975 116.335 182.145 ;
        RECT 116.975 182.055 117.145 183.185 ;
        RECT 115.125 181.555 115.385 181.975 ;
        RECT 115.555 181.375 115.885 181.805 ;
        RECT 116.165 181.715 116.335 181.975 ;
        RECT 116.550 181.885 117.145 182.055 ;
        RECT 117.315 181.715 117.485 183.015 ;
        RECT 117.715 182.560 118.045 183.015 ;
        RECT 116.165 181.545 117.485 181.715 ;
        RECT 117.835 182.225 118.045 182.560 ;
        RECT 118.275 182.565 118.445 183.015 ;
        RECT 118.615 182.935 118.785 183.185 ;
        RECT 118.955 183.285 119.205 183.755 ;
        RECT 119.375 183.455 119.545 183.925 ;
        RECT 119.715 183.285 120.045 183.755 ;
        RECT 120.215 183.455 120.385 183.925 ;
        RECT 118.955 183.105 120.475 183.285 ;
        RECT 120.735 183.275 120.905 183.755 ;
        RECT 121.075 183.445 121.405 183.925 ;
        RECT 121.630 183.505 123.165 183.755 ;
        RECT 121.630 183.275 121.800 183.505 ;
        RECT 120.735 183.105 121.800 183.275 ;
        RECT 118.615 182.765 120.075 182.935 ;
        RECT 118.275 182.395 118.710 182.565 ;
        RECT 120.245 182.555 120.475 183.105 ;
        RECT 121.980 182.935 122.260 183.335 ;
        RECT 120.645 182.725 121.000 182.935 ;
        RECT 121.170 182.735 121.615 182.935 ;
        RECT 121.785 182.735 122.260 182.935 ;
        RECT 122.530 182.935 122.815 183.335 ;
        RECT 122.995 183.275 123.165 183.505 ;
        RECT 123.335 183.445 123.665 183.925 ;
        RECT 123.880 183.425 124.135 183.755 ;
        RECT 123.925 183.415 124.135 183.425 ;
        RECT 123.950 183.345 124.135 183.415 ;
        RECT 122.995 183.105 123.795 183.275 ;
        RECT 122.530 182.735 122.860 182.935 ;
        RECT 123.030 182.735 123.395 182.935 ;
        RECT 123.625 182.555 123.795 183.105 ;
        RECT 118.915 182.385 120.475 182.555 ;
        RECT 120.735 182.385 123.795 182.555 ;
        RECT 117.835 181.635 118.155 182.225 ;
        RECT 118.440 181.375 118.690 182.215 ;
        RECT 118.915 181.545 119.165 182.385 ;
        RECT 119.335 181.375 119.585 182.215 ;
        RECT 119.755 181.545 120.005 182.385 ;
        RECT 120.175 181.375 120.425 182.215 ;
        RECT 120.735 181.545 120.905 182.385 ;
        RECT 123.965 182.215 124.135 183.345 ;
        RECT 124.305 183.030 124.475 183.925 ;
        RECT 124.785 183.250 125.045 183.755 ;
        RECT 125.225 183.545 125.555 183.925 ;
        RECT 125.735 183.375 125.905 183.755 ;
        RECT 121.075 181.715 121.405 182.215 ;
        RECT 121.575 181.975 123.210 182.215 ;
        RECT 121.575 181.885 121.805 181.975 ;
        RECT 121.915 181.715 122.245 181.755 ;
        RECT 121.075 181.545 122.245 181.715 ;
        RECT 122.435 181.375 122.790 181.795 ;
        RECT 122.960 181.545 123.210 181.975 ;
        RECT 123.380 181.375 123.710 182.135 ;
        RECT 123.880 181.545 124.135 182.215 ;
        RECT 124.305 181.375 124.475 182.565 ;
        RECT 124.785 182.450 124.965 183.250 ;
        RECT 125.240 183.205 125.905 183.375 ;
        RECT 125.240 182.950 125.410 183.205 ;
        RECT 126.625 183.200 126.915 183.925 ;
        RECT 127.090 183.105 127.365 183.925 ;
        RECT 127.535 183.285 127.865 183.755 ;
        RECT 128.035 183.455 128.205 183.925 ;
        RECT 128.375 183.285 128.705 183.755 ;
        RECT 128.875 183.455 129.165 183.925 ;
        RECT 127.535 183.275 128.705 183.285 ;
        RECT 127.535 183.105 129.135 183.275 ;
        RECT 125.135 182.620 125.410 182.950 ;
        RECT 125.635 182.655 125.975 183.025 ;
        RECT 127.090 182.735 127.810 182.935 ;
        RECT 127.980 182.735 128.750 182.935 ;
        RECT 125.240 182.475 125.410 182.620 ;
        RECT 128.920 182.565 129.135 183.105 ;
        RECT 124.785 181.545 125.055 182.450 ;
        RECT 125.240 182.305 125.915 182.475 ;
        RECT 125.225 181.375 125.555 182.135 ;
        RECT 125.735 181.545 125.915 182.305 ;
        RECT 126.625 181.375 126.915 182.540 ;
        RECT 127.090 182.345 128.205 182.555 ;
        RECT 127.090 181.545 127.365 182.345 ;
        RECT 127.535 181.375 127.865 182.175 ;
        RECT 128.035 181.715 128.205 182.345 ;
        RECT 128.375 182.345 129.135 182.565 ;
        RECT 129.385 183.185 129.745 183.560 ;
        RECT 130.010 183.185 130.180 183.925 ;
        RECT 130.460 183.355 130.630 183.560 ;
        RECT 130.460 183.185 131.000 183.355 ;
        RECT 129.385 182.530 129.640 183.185 ;
        RECT 129.810 182.685 130.160 183.015 ;
        RECT 130.330 182.685 130.660 183.015 ;
        RECT 128.375 181.885 128.705 182.345 ;
        RECT 128.875 181.715 129.175 182.175 ;
        RECT 128.035 181.545 129.175 181.715 ;
        RECT 129.385 181.545 129.725 182.530 ;
        RECT 129.895 182.145 130.160 182.685 ;
        RECT 130.830 182.485 131.000 183.185 ;
        RECT 130.375 182.315 131.000 182.485 ;
        RECT 131.170 182.555 131.340 183.755 ;
        RECT 131.570 183.275 131.900 183.755 ;
        RECT 132.070 183.455 132.240 183.925 ;
        RECT 132.410 183.275 132.740 183.740 ;
        RECT 131.570 183.105 132.740 183.275 ;
        RECT 133.065 183.250 133.325 183.755 ;
        RECT 133.505 183.545 133.835 183.925 ;
        RECT 134.015 183.375 134.185 183.755 ;
        RECT 131.510 182.725 132.080 182.935 ;
        RECT 132.250 182.725 132.895 182.935 ;
        RECT 131.170 182.145 131.875 182.555 ;
        RECT 129.895 181.975 131.875 182.145 ;
        RECT 129.895 181.375 130.305 181.805 ;
        RECT 131.050 181.375 131.380 181.795 ;
        RECT 131.550 181.545 131.875 181.975 ;
        RECT 132.350 181.375 132.680 182.475 ;
        RECT 133.065 182.450 133.235 183.250 ;
        RECT 133.520 183.205 134.185 183.375 ;
        RECT 133.520 182.950 133.690 183.205 ;
        RECT 134.905 183.175 136.115 183.925 ;
        RECT 133.405 182.620 133.690 182.950 ;
        RECT 133.925 182.655 134.255 183.025 ;
        RECT 133.520 182.475 133.690 182.620 ;
        RECT 133.065 181.545 133.335 182.450 ;
        RECT 133.520 182.305 134.185 182.475 ;
        RECT 133.505 181.375 133.835 182.135 ;
        RECT 134.015 181.545 134.185 182.305 ;
        RECT 134.905 182.465 135.425 183.005 ;
        RECT 135.595 182.635 136.115 183.175 ;
        RECT 134.905 181.375 136.115 182.465 ;
        RECT 23.500 181.205 136.200 181.375 ;
        RECT 23.585 180.115 24.795 181.205 ;
        RECT 24.965 180.610 25.400 181.035 ;
        RECT 25.570 180.780 25.955 181.205 ;
        RECT 24.965 180.440 25.955 180.610 ;
        RECT 23.585 179.405 24.105 179.945 ;
        RECT 24.275 179.575 24.795 180.115 ;
        RECT 24.965 179.565 25.450 180.270 ;
        RECT 25.620 179.895 25.955 180.440 ;
        RECT 26.125 180.245 26.550 181.035 ;
        RECT 26.720 180.610 26.995 181.035 ;
        RECT 27.165 180.780 27.550 181.205 ;
        RECT 26.720 180.415 27.550 180.610 ;
        RECT 26.125 180.065 27.030 180.245 ;
        RECT 25.620 179.565 26.030 179.895 ;
        RECT 26.200 179.565 27.030 180.065 ;
        RECT 27.200 179.895 27.550 180.415 ;
        RECT 27.720 180.245 27.965 181.035 ;
        RECT 28.155 180.610 28.410 181.035 ;
        RECT 28.580 180.780 28.965 181.205 ;
        RECT 28.155 180.415 28.965 180.610 ;
        RECT 27.720 180.065 28.445 180.245 ;
        RECT 27.200 179.565 27.625 179.895 ;
        RECT 27.795 179.565 28.445 180.065 ;
        RECT 28.615 179.895 28.965 180.415 ;
        RECT 29.135 180.065 29.395 181.035 ;
        RECT 29.565 180.115 33.075 181.205 ;
        RECT 33.245 180.115 34.455 181.205 ;
        RECT 28.615 179.565 29.040 179.895 ;
        RECT 23.585 178.655 24.795 179.405 ;
        RECT 25.620 179.395 25.955 179.565 ;
        RECT 26.200 179.395 26.550 179.565 ;
        RECT 27.200 179.395 27.550 179.565 ;
        RECT 27.795 179.395 27.965 179.565 ;
        RECT 28.615 179.395 28.965 179.565 ;
        RECT 29.210 179.395 29.395 180.065 ;
        RECT 24.965 179.225 25.955 179.395 ;
        RECT 24.965 178.825 25.400 179.225 ;
        RECT 25.570 178.655 25.955 179.055 ;
        RECT 26.125 178.825 26.550 179.395 ;
        RECT 26.740 179.225 27.550 179.395 ;
        RECT 26.740 178.825 26.995 179.225 ;
        RECT 27.165 178.655 27.550 179.055 ;
        RECT 27.720 178.825 27.965 179.395 ;
        RECT 28.155 179.225 28.965 179.395 ;
        RECT 28.155 178.825 28.410 179.225 ;
        RECT 28.580 178.655 28.965 179.055 ;
        RECT 29.135 178.825 29.395 179.395 ;
        RECT 29.565 179.425 31.215 179.945 ;
        RECT 31.385 179.595 33.075 180.115 ;
        RECT 29.565 178.655 33.075 179.425 ;
        RECT 33.245 179.405 33.765 179.945 ;
        RECT 33.935 179.575 34.455 180.115 ;
        RECT 34.630 180.065 34.950 181.205 ;
        RECT 35.130 179.895 35.325 180.945 ;
        RECT 35.505 180.355 35.835 181.035 ;
        RECT 36.035 180.405 36.290 181.205 ;
        RECT 35.505 180.075 35.855 180.355 ;
        RECT 34.690 179.845 34.950 179.895 ;
        RECT 34.685 179.675 34.950 179.845 ;
        RECT 34.690 179.565 34.950 179.675 ;
        RECT 35.130 179.565 35.515 179.895 ;
        RECT 35.685 179.695 35.855 180.075 ;
        RECT 36.045 179.865 36.290 180.225 ;
        RECT 36.465 180.040 36.755 181.205 ;
        RECT 37.015 180.275 37.185 181.035 ;
        RECT 37.400 180.445 37.730 181.205 ;
        RECT 37.015 180.105 37.730 180.275 ;
        RECT 37.900 180.130 38.155 181.035 ;
        RECT 35.685 179.525 36.205 179.695 ;
        RECT 36.925 179.555 37.280 179.925 ;
        RECT 37.560 179.895 37.730 180.105 ;
        RECT 37.560 179.565 37.815 179.895 ;
        RECT 33.245 178.655 34.455 179.405 ;
        RECT 34.630 179.185 35.845 179.355 ;
        RECT 34.630 178.835 34.920 179.185 ;
        RECT 35.115 178.655 35.445 179.015 ;
        RECT 35.615 178.880 35.845 179.185 ;
        RECT 36.035 178.960 36.205 179.525 ;
        RECT 36.465 178.655 36.755 179.380 ;
        RECT 37.560 179.375 37.730 179.565 ;
        RECT 37.985 179.400 38.155 180.130 ;
        RECT 38.330 180.055 38.590 181.205 ;
        RECT 38.770 180.065 39.090 181.205 ;
        RECT 39.270 179.895 39.465 180.945 ;
        RECT 39.645 180.355 39.975 181.035 ;
        RECT 40.175 180.405 40.430 181.205 ;
        RECT 39.645 180.075 39.995 180.355 ;
        RECT 38.830 179.845 39.090 179.895 ;
        RECT 38.825 179.675 39.090 179.845 ;
        RECT 38.830 179.565 39.090 179.675 ;
        RECT 39.270 179.565 39.655 179.895 ;
        RECT 39.825 179.695 39.995 180.075 ;
        RECT 40.185 179.865 40.430 180.225 ;
        RECT 40.645 180.065 40.875 181.205 ;
        RECT 41.045 180.055 41.375 181.035 ;
        RECT 41.545 180.065 41.755 181.205 ;
        RECT 41.985 180.115 44.575 181.205 ;
        RECT 39.825 179.525 40.345 179.695 ;
        RECT 40.625 179.645 40.955 179.895 ;
        RECT 37.015 179.205 37.730 179.375 ;
        RECT 37.015 178.825 37.185 179.205 ;
        RECT 37.400 178.655 37.730 179.035 ;
        RECT 37.900 178.825 38.155 179.400 ;
        RECT 38.330 178.655 38.590 179.495 ;
        RECT 38.770 179.185 39.985 179.355 ;
        RECT 38.770 178.835 39.060 179.185 ;
        RECT 39.255 178.655 39.585 179.015 ;
        RECT 39.755 178.880 39.985 179.185 ;
        RECT 40.175 178.960 40.345 179.525 ;
        RECT 40.645 178.655 40.875 179.475 ;
        RECT 41.125 179.455 41.375 180.055 ;
        RECT 41.045 178.825 41.375 179.455 ;
        RECT 41.545 178.655 41.755 179.475 ;
        RECT 41.985 179.425 43.195 179.945 ;
        RECT 43.365 179.595 44.575 180.115 ;
        RECT 44.775 180.015 45.025 181.205 ;
        RECT 41.985 178.655 44.575 179.425 ;
        RECT 44.845 178.655 45.015 179.455 ;
        RECT 45.250 178.935 45.465 181.035 ;
        RECT 45.655 180.445 46.455 181.205 ;
        RECT 46.850 180.275 47.235 181.035 ;
        RECT 45.635 180.065 47.235 180.275 ;
        RECT 47.560 180.185 47.760 180.975 ;
        RECT 47.930 180.365 48.250 181.205 ;
        RECT 45.635 179.465 45.915 180.065 ;
        RECT 47.405 180.015 47.760 180.185 ;
        RECT 47.405 179.895 47.585 180.015 ;
        RECT 46.095 179.645 46.450 179.895 ;
        RECT 46.620 179.645 47.085 179.895 ;
        RECT 47.255 179.645 47.585 179.895 ;
        RECT 47.930 179.845 48.250 180.185 ;
        RECT 47.755 179.645 48.250 179.845 ;
        RECT 48.425 180.065 48.810 181.025 ;
        RECT 49.025 180.405 49.315 181.205 ;
        RECT 49.485 180.865 50.850 181.035 ;
        RECT 49.485 180.235 49.655 180.865 ;
        RECT 48.980 180.065 49.655 180.235 ;
        RECT 45.635 179.285 46.875 179.465 ;
        RECT 47.220 179.395 48.250 179.435 ;
        RECT 46.510 179.215 46.875 179.285 ;
        RECT 47.050 179.265 48.250 179.395 ;
        RECT 45.685 178.655 45.865 179.115 ;
        RECT 47.050 179.045 47.390 179.265 ;
        RECT 46.125 178.865 47.390 179.045 ;
        RECT 47.575 178.655 47.745 179.095 ;
        RECT 47.915 178.850 48.250 179.265 ;
        RECT 48.425 179.395 48.600 180.065 ;
        RECT 48.980 179.895 49.150 180.065 ;
        RECT 49.825 179.895 50.150 180.695 ;
        RECT 50.520 180.655 50.850 180.865 ;
        RECT 50.520 180.405 51.475 180.655 ;
        RECT 48.785 179.645 49.150 179.895 ;
        RECT 49.345 179.645 49.595 179.895 ;
        RECT 48.785 179.565 48.975 179.645 ;
        RECT 49.345 179.565 49.515 179.645 ;
        RECT 49.805 179.565 50.150 179.895 ;
        RECT 50.320 179.565 50.595 180.230 ;
        RECT 50.780 179.565 51.135 180.230 ;
        RECT 51.305 179.395 51.475 180.405 ;
        RECT 51.645 180.065 51.935 181.205 ;
        RECT 52.105 180.065 52.365 181.205 ;
        RECT 52.535 180.055 52.865 181.035 ;
        RECT 53.035 180.065 53.315 181.205 ;
        RECT 53.945 180.485 54.405 181.035 ;
        RECT 54.595 180.485 54.925 181.205 ;
        RECT 51.660 179.565 51.935 179.895 ;
        RECT 52.125 179.645 52.460 179.895 ;
        RECT 52.630 179.455 52.800 180.055 ;
        RECT 52.970 179.625 53.305 179.895 ;
        RECT 48.425 178.825 48.935 179.395 ;
        RECT 49.480 179.225 50.880 179.395 ;
        RECT 49.105 178.655 49.275 179.215 ;
        RECT 49.480 178.825 49.810 179.225 ;
        RECT 49.985 178.655 50.315 179.055 ;
        RECT 50.550 179.035 50.880 179.225 ;
        RECT 51.050 179.205 51.475 179.395 ;
        RECT 51.645 179.035 51.935 179.305 ;
        RECT 50.550 178.825 51.935 179.035 ;
        RECT 52.105 178.825 52.800 179.455 ;
        RECT 53.005 178.655 53.315 179.455 ;
        RECT 53.945 179.115 54.195 180.485 ;
        RECT 55.125 180.315 55.425 180.865 ;
        RECT 55.595 180.535 55.875 181.205 ;
        RECT 54.485 180.145 55.425 180.315 ;
        RECT 54.485 179.895 54.655 180.145 ;
        RECT 55.795 179.895 56.060 180.255 ;
        RECT 56.250 180.065 56.570 181.205 ;
        RECT 56.750 179.895 56.945 180.945 ;
        RECT 57.125 180.355 57.455 181.035 ;
        RECT 57.655 180.405 57.910 181.205 ;
        RECT 58.190 180.745 58.360 181.205 ;
        RECT 58.530 180.575 58.860 181.035 ;
        RECT 58.085 180.405 58.860 180.575 ;
        RECT 59.030 180.405 59.200 181.205 ;
        RECT 60.395 180.595 60.725 181.025 ;
        RECT 60.905 180.765 61.100 181.205 ;
        RECT 61.270 180.595 61.600 181.025 ;
        RECT 60.395 180.425 61.600 180.595 ;
        RECT 57.125 180.075 57.475 180.355 ;
        RECT 54.365 179.565 54.655 179.895 ;
        RECT 54.825 179.645 55.165 179.895 ;
        RECT 55.385 179.645 56.060 179.895 ;
        RECT 56.310 179.845 56.570 179.895 ;
        RECT 56.305 179.675 56.570 179.845 ;
        RECT 56.310 179.565 56.570 179.675 ;
        RECT 56.750 179.565 57.135 179.895 ;
        RECT 57.305 179.695 57.475 180.075 ;
        RECT 57.665 179.865 57.910 180.225 ;
        RECT 54.485 179.475 54.655 179.565 ;
        RECT 57.305 179.525 57.825 179.695 ;
        RECT 54.485 179.285 55.875 179.475 ;
        RECT 53.945 178.825 54.505 179.115 ;
        RECT 54.675 178.655 54.925 179.115 ;
        RECT 55.545 178.925 55.875 179.285 ;
        RECT 56.250 179.185 57.465 179.355 ;
        RECT 56.250 178.835 56.540 179.185 ;
        RECT 56.735 178.655 57.065 179.015 ;
        RECT 57.235 178.880 57.465 179.185 ;
        RECT 57.655 178.960 57.825 179.525 ;
        RECT 58.085 179.395 58.515 180.405 ;
        RECT 59.785 180.235 60.145 180.410 ;
        RECT 58.685 180.065 60.145 180.235 ;
        RECT 60.395 180.095 61.290 180.425 ;
        RECT 61.770 180.255 62.045 181.025 ;
        RECT 61.460 180.065 62.045 180.255 ;
        RECT 58.685 179.565 58.855 180.065 ;
        RECT 58.085 179.225 58.780 179.395 ;
        RECT 59.025 179.335 59.435 179.895 ;
        RECT 58.110 178.655 58.440 179.055 ;
        RECT 58.610 178.955 58.780 179.225 ;
        RECT 59.605 179.165 59.785 180.065 ;
        RECT 59.955 179.505 60.150 179.895 ;
        RECT 60.400 179.565 60.695 179.895 ;
        RECT 60.875 179.565 61.290 179.895 ;
        RECT 59.955 179.335 60.155 179.505 ;
        RECT 58.950 178.655 59.265 179.165 ;
        RECT 59.495 178.825 59.785 179.165 ;
        RECT 59.955 178.655 60.195 179.165 ;
        RECT 60.395 178.655 60.695 179.385 ;
        RECT 60.875 178.945 61.105 179.565 ;
        RECT 61.460 179.395 61.635 180.065 ;
        RECT 62.225 180.040 62.515 181.205 ;
        RECT 62.690 180.485 63.025 180.995 ;
        RECT 61.305 179.215 61.635 179.395 ;
        RECT 61.805 179.245 62.045 179.895 ;
        RECT 61.305 178.835 61.530 179.215 ;
        RECT 61.700 178.655 62.030 179.045 ;
        RECT 62.225 178.655 62.515 179.380 ;
        RECT 62.690 179.130 62.945 180.485 ;
        RECT 63.275 180.405 63.605 181.205 ;
        RECT 63.850 180.615 64.135 181.035 ;
        RECT 64.390 180.785 64.720 181.205 ;
        RECT 64.945 180.865 66.105 181.035 ;
        RECT 64.945 180.615 65.275 180.865 ;
        RECT 63.850 180.445 65.275 180.615 ;
        RECT 65.505 180.235 65.675 180.695 ;
        RECT 65.935 180.365 66.105 180.865 ;
        RECT 66.385 180.365 66.640 181.035 ;
        RECT 66.810 180.445 67.140 181.205 ;
        RECT 67.310 180.605 67.560 181.035 ;
        RECT 67.730 180.785 68.085 181.205 ;
        RECT 68.275 180.865 69.445 181.035 ;
        RECT 68.275 180.825 68.605 180.865 ;
        RECT 68.715 180.605 68.945 180.695 ;
        RECT 67.310 180.365 68.945 180.605 ;
        RECT 69.115 180.365 69.445 180.865 ;
        RECT 63.305 180.065 65.675 180.235 ;
        RECT 63.305 179.895 63.475 180.065 ;
        RECT 65.925 180.015 66.135 180.185 ;
        RECT 65.925 179.895 66.130 180.015 ;
        RECT 63.170 179.565 63.475 179.895 ;
        RECT 63.670 179.845 63.920 179.895 ;
        RECT 63.665 179.675 63.920 179.845 ;
        RECT 63.670 179.565 63.920 179.675 ;
        RECT 63.305 179.395 63.475 179.565 ;
        RECT 64.130 179.505 64.400 179.895 ;
        RECT 63.305 179.225 63.865 179.395 ;
        RECT 64.125 179.335 64.400 179.505 ;
        RECT 64.130 179.235 64.400 179.335 ;
        RECT 64.590 179.235 64.880 179.895 ;
        RECT 65.050 179.230 65.470 179.895 ;
        RECT 65.780 179.565 66.130 179.895 ;
        RECT 62.690 178.870 63.025 179.130 ;
        RECT 63.695 179.055 63.865 179.225 ;
        RECT 63.195 178.655 63.525 179.055 ;
        RECT 63.695 178.885 65.310 179.055 ;
        RECT 65.855 178.655 66.185 179.375 ;
        RECT 66.385 179.235 66.555 180.365 ;
        RECT 69.615 180.195 69.785 181.035 ;
        RECT 70.045 180.770 75.390 181.205 ;
        RECT 66.725 180.025 69.785 180.195 ;
        RECT 66.725 179.475 66.895 180.025 ;
        RECT 67.125 179.645 67.490 179.845 ;
        RECT 67.660 179.645 67.990 179.845 ;
        RECT 66.725 179.305 67.525 179.475 ;
        RECT 66.385 179.165 66.570 179.235 ;
        RECT 66.385 179.155 66.595 179.165 ;
        RECT 66.385 178.825 66.640 179.155 ;
        RECT 66.855 178.655 67.185 179.135 ;
        RECT 67.355 179.075 67.525 179.305 ;
        RECT 67.705 179.245 67.990 179.645 ;
        RECT 68.260 179.645 68.735 179.845 ;
        RECT 68.905 179.645 69.350 179.845 ;
        RECT 69.520 179.645 69.870 179.855 ;
        RECT 68.260 179.245 68.540 179.645 ;
        RECT 68.720 179.305 69.785 179.475 ;
        RECT 68.720 179.075 68.890 179.305 ;
        RECT 67.355 178.825 68.890 179.075 ;
        RECT 69.115 178.655 69.445 179.135 ;
        RECT 69.615 178.825 69.785 179.305 ;
        RECT 71.630 179.200 71.970 180.030 ;
        RECT 73.450 179.520 73.800 180.770 ;
        RECT 75.565 180.115 77.235 181.205 ;
        RECT 75.565 179.425 76.315 179.945 ;
        RECT 76.485 179.595 77.235 180.115 ;
        RECT 77.410 180.065 77.730 181.205 ;
        RECT 77.910 179.895 78.105 180.945 ;
        RECT 78.285 180.355 78.615 181.035 ;
        RECT 78.815 180.405 79.070 181.205 ;
        RECT 79.245 180.405 79.685 181.035 ;
        RECT 78.285 180.075 78.635 180.355 ;
        RECT 77.470 179.845 77.730 179.895 ;
        RECT 77.465 179.675 77.730 179.845 ;
        RECT 77.470 179.565 77.730 179.675 ;
        RECT 77.910 179.565 78.295 179.895 ;
        RECT 78.465 179.695 78.635 180.075 ;
        RECT 78.825 179.865 79.070 180.225 ;
        RECT 78.465 179.525 78.985 179.695 ;
        RECT 70.045 178.655 75.390 179.200 ;
        RECT 75.565 178.655 77.235 179.425 ;
        RECT 77.410 179.185 78.625 179.355 ;
        RECT 77.410 178.835 77.700 179.185 ;
        RECT 77.895 178.655 78.225 179.015 ;
        RECT 78.395 178.880 78.625 179.185 ;
        RECT 78.815 178.960 78.985 179.525 ;
        RECT 79.245 179.395 79.555 180.405 ;
        RECT 79.860 180.355 80.175 181.205 ;
        RECT 80.345 180.865 81.775 181.035 ;
        RECT 80.345 180.185 80.515 180.865 ;
        RECT 79.725 180.015 80.515 180.185 ;
        RECT 79.725 179.565 79.895 180.015 ;
        RECT 80.685 179.895 80.885 180.695 ;
        RECT 80.065 179.565 80.455 179.845 ;
        RECT 80.640 179.565 80.885 179.895 ;
        RECT 81.085 179.565 81.335 180.695 ;
        RECT 81.525 180.235 81.775 180.865 ;
        RECT 81.955 180.405 82.285 181.205 ;
        RECT 82.465 180.405 82.905 181.035 ;
        RECT 81.525 180.065 82.295 180.235 ;
        RECT 81.550 179.565 81.955 179.895 ;
        RECT 82.125 179.395 82.295 180.065 ;
        RECT 79.245 178.835 79.685 179.395 ;
        RECT 79.855 178.655 80.305 179.395 ;
        RECT 80.475 179.225 81.635 179.395 ;
        RECT 80.475 178.825 80.645 179.225 ;
        RECT 80.815 178.655 81.235 179.055 ;
        RECT 81.405 178.825 81.635 179.225 ;
        RECT 81.805 178.825 82.295 179.395 ;
        RECT 82.465 179.395 82.775 180.405 ;
        RECT 83.080 180.355 83.395 181.205 ;
        RECT 83.565 180.865 84.995 181.035 ;
        RECT 83.565 180.185 83.735 180.865 ;
        RECT 82.945 180.015 83.735 180.185 ;
        RECT 82.945 179.565 83.115 180.015 ;
        RECT 83.905 179.895 84.105 180.695 ;
        RECT 83.285 179.565 83.675 179.845 ;
        RECT 83.860 179.565 84.105 179.895 ;
        RECT 84.305 179.565 84.555 180.695 ;
        RECT 84.745 180.235 84.995 180.865 ;
        RECT 85.175 180.405 85.505 181.205 ;
        RECT 84.745 180.065 85.515 180.235 ;
        RECT 85.685 180.065 85.945 181.205 ;
        RECT 84.770 179.565 85.175 179.895 ;
        RECT 85.345 179.395 85.515 180.065 ;
        RECT 86.115 180.055 86.445 181.035 ;
        RECT 86.615 180.065 86.895 181.205 ;
        RECT 86.205 180.015 86.380 180.055 ;
        RECT 87.985 180.040 88.275 181.205 ;
        RECT 88.450 180.485 88.785 180.995 ;
        RECT 85.705 179.645 86.040 179.895 ;
        RECT 86.210 179.455 86.380 180.015 ;
        RECT 86.550 179.625 86.885 179.895 ;
        RECT 82.465 178.835 82.905 179.395 ;
        RECT 83.075 178.655 83.525 179.395 ;
        RECT 83.695 179.225 84.855 179.395 ;
        RECT 83.695 178.825 83.865 179.225 ;
        RECT 84.035 178.655 84.455 179.055 ;
        RECT 84.625 178.825 84.855 179.225 ;
        RECT 85.025 178.825 85.515 179.395 ;
        RECT 85.685 178.825 86.380 179.455 ;
        RECT 86.585 178.655 86.895 179.455 ;
        RECT 87.985 178.655 88.275 179.380 ;
        RECT 88.450 179.130 88.705 180.485 ;
        RECT 89.035 180.405 89.365 181.205 ;
        RECT 89.610 180.615 89.895 181.035 ;
        RECT 90.150 180.785 90.480 181.205 ;
        RECT 90.705 180.865 91.865 181.035 ;
        RECT 90.705 180.615 91.035 180.865 ;
        RECT 89.610 180.445 91.035 180.615 ;
        RECT 91.265 180.235 91.435 180.695 ;
        RECT 91.695 180.365 91.865 180.865 ;
        RECT 89.065 180.065 91.435 180.235 ;
        RECT 89.065 179.895 89.235 180.065 ;
        RECT 91.685 180.015 91.895 180.185 ;
        RECT 91.685 179.895 91.890 180.015 ;
        RECT 88.930 179.565 89.235 179.895 ;
        RECT 89.430 179.845 89.680 179.895 ;
        RECT 89.425 179.675 89.680 179.845 ;
        RECT 89.430 179.565 89.680 179.675 ;
        RECT 89.065 179.395 89.235 179.565 ;
        RECT 89.890 179.505 90.160 179.895 ;
        RECT 90.350 179.845 90.640 179.895 ;
        RECT 90.345 179.675 90.640 179.845 ;
        RECT 89.065 179.225 89.625 179.395 ;
        RECT 89.885 179.335 90.160 179.505 ;
        RECT 89.890 179.235 90.160 179.335 ;
        RECT 90.350 179.235 90.640 179.675 ;
        RECT 90.810 179.230 91.230 179.895 ;
        RECT 91.540 179.565 91.890 179.895 ;
        RECT 88.450 178.870 88.785 179.130 ;
        RECT 89.455 179.055 89.625 179.225 ;
        RECT 88.955 178.655 89.285 179.055 ;
        RECT 89.455 178.885 91.070 179.055 ;
        RECT 91.615 178.655 91.945 179.375 ;
        RECT 92.125 178.825 92.875 181.035 ;
        RECT 93.135 180.275 93.305 181.035 ;
        RECT 93.485 180.445 93.815 181.205 ;
        RECT 93.135 180.105 93.800 180.275 ;
        RECT 93.985 180.130 94.255 181.035 ;
        RECT 94.425 180.195 94.690 181.205 ;
        RECT 94.860 180.365 95.145 181.035 ;
        RECT 93.630 179.960 93.800 180.105 ;
        RECT 93.065 179.555 93.395 179.925 ;
        RECT 93.630 179.630 93.915 179.960 ;
        RECT 93.630 179.375 93.800 179.630 ;
        RECT 93.135 179.205 93.800 179.375 ;
        RECT 94.085 179.330 94.255 180.130 ;
        RECT 94.860 180.015 95.030 180.365 ;
        RECT 95.345 180.360 95.560 181.205 ;
        RECT 95.730 180.695 96.205 181.035 ;
        RECT 96.375 180.700 96.990 181.205 ;
        RECT 96.375 180.525 96.565 180.700 ;
        RECT 95.820 180.165 96.010 180.460 ;
        RECT 96.235 180.335 96.565 180.525 ;
        RECT 96.735 180.165 96.970 180.530 ;
        RECT 94.425 179.495 95.030 180.015 ;
        RECT 95.200 179.995 96.970 180.165 ;
        RECT 95.200 179.565 95.430 179.995 ;
        RECT 93.135 178.825 93.305 179.205 ;
        RECT 93.485 178.655 93.815 179.035 ;
        RECT 93.995 178.825 94.255 179.330 ;
        RECT 94.425 178.655 94.690 179.315 ;
        RECT 94.860 179.285 95.030 179.495 ;
        RECT 95.600 179.335 96.010 179.815 ;
        RECT 94.860 178.825 95.105 179.285 ;
        RECT 95.280 178.655 95.610 179.150 ;
        RECT 95.800 178.875 96.010 179.335 ;
        RECT 96.180 179.140 96.435 179.995 ;
        RECT 97.165 179.815 97.440 180.475 ;
        RECT 97.620 180.145 97.935 181.205 ;
        RECT 98.105 180.485 98.565 181.035 ;
        RECT 98.755 180.485 99.085 181.205 ;
        RECT 96.605 179.585 97.440 179.815 ;
        RECT 96.180 178.875 96.965 179.140 ;
        RECT 97.165 178.875 97.440 179.585 ;
        RECT 97.610 179.315 97.875 179.895 ;
        RECT 97.665 178.655 97.935 179.145 ;
        RECT 98.105 179.115 98.355 180.485 ;
        RECT 99.285 180.315 99.585 180.865 ;
        RECT 99.755 180.535 100.035 181.205 ;
        RECT 98.645 180.145 99.585 180.315 ;
        RECT 98.645 179.895 98.815 180.145 ;
        RECT 99.955 179.895 100.220 180.255 ;
        RECT 98.525 179.565 98.815 179.895 ;
        RECT 98.985 179.645 99.325 179.895 ;
        RECT 99.545 179.645 100.220 179.895 ;
        RECT 101.325 179.915 101.595 181.015 ;
        RECT 101.765 180.275 102.040 180.780 ;
        RECT 102.210 180.445 102.540 181.205 ;
        RECT 101.765 180.105 102.255 180.275 ;
        RECT 102.710 180.195 103.035 181.035 ;
        RECT 101.325 179.565 101.775 179.915 ;
        RECT 101.960 179.565 102.255 180.105 ;
        RECT 102.425 180.025 103.035 180.195 ;
        RECT 103.510 180.105 103.885 181.205 ;
        RECT 104.140 180.335 104.425 181.205 ;
        RECT 104.595 180.575 104.855 181.035 ;
        RECT 105.030 180.745 105.285 181.205 ;
        RECT 105.455 180.575 105.715 181.035 ;
        RECT 104.595 180.405 105.715 180.575 ;
        RECT 105.885 180.405 106.195 181.205 ;
        RECT 104.595 180.155 104.855 180.405 ;
        RECT 106.365 180.235 106.675 181.035 ;
        RECT 98.645 179.475 98.815 179.565 ;
        RECT 98.645 179.285 100.035 179.475 ;
        RECT 101.960 179.395 102.130 179.565 ;
        RECT 102.425 179.395 102.595 180.025 ;
        RECT 104.100 179.985 104.855 180.155 ;
        RECT 105.645 180.065 106.675 180.235 ;
        RECT 102.765 179.645 103.265 179.855 ;
        RECT 103.435 179.645 103.915 179.855 ;
        RECT 104.100 179.475 104.505 179.985 ;
        RECT 105.645 179.815 105.815 180.065 ;
        RECT 104.675 179.645 105.815 179.815 ;
        RECT 98.105 178.825 98.665 179.115 ;
        RECT 98.835 178.655 99.085 179.115 ;
        RECT 99.705 178.925 100.035 179.285 ;
        RECT 101.325 178.655 101.600 179.395 ;
        RECT 101.820 179.225 102.130 179.395 ;
        RECT 101.820 179.065 102.010 179.225 ;
        RECT 102.355 179.215 102.595 179.395 ;
        RECT 102.810 179.305 103.905 179.475 ;
        RECT 104.100 179.305 105.750 179.475 ;
        RECT 105.985 179.325 106.335 179.895 ;
        RECT 102.355 179.165 102.525 179.215 ;
        RECT 102.305 178.995 102.525 179.165 ;
        RECT 102.810 179.055 102.980 179.305 ;
        RECT 102.355 178.825 102.525 178.995 ;
        RECT 102.730 178.825 103.060 179.055 ;
        RECT 103.235 178.655 103.405 179.125 ;
        RECT 103.575 178.840 103.905 179.305 ;
        RECT 104.145 178.655 104.425 179.135 ;
        RECT 104.595 178.915 104.855 179.305 ;
        RECT 105.030 178.655 105.285 179.135 ;
        RECT 105.455 178.915 105.750 179.305 ;
        RECT 106.505 179.155 106.675 180.065 ;
        RECT 106.850 180.815 107.185 181.035 ;
        RECT 108.190 180.825 108.545 181.205 ;
        RECT 106.850 180.195 107.105 180.815 ;
        RECT 107.355 180.655 107.585 180.695 ;
        RECT 108.715 180.655 108.965 181.035 ;
        RECT 107.355 180.455 108.965 180.655 ;
        RECT 107.355 180.365 107.540 180.455 ;
        RECT 108.130 180.445 108.965 180.455 ;
        RECT 109.215 180.425 109.465 181.205 ;
        RECT 109.635 180.355 109.895 181.035 ;
        RECT 110.075 180.825 110.405 181.205 ;
        RECT 107.695 180.255 108.025 180.285 ;
        RECT 107.695 180.195 109.495 180.255 ;
        RECT 106.850 180.085 109.555 180.195 ;
        RECT 106.850 180.025 108.025 180.085 ;
        RECT 109.355 180.050 109.555 180.085 ;
        RECT 106.845 179.645 107.335 179.845 ;
        RECT 107.525 179.645 108.000 179.855 ;
        RECT 105.930 178.655 106.205 179.135 ;
        RECT 106.375 178.825 106.675 179.155 ;
        RECT 106.850 178.655 107.305 179.420 ;
        RECT 107.780 179.245 108.000 179.645 ;
        RECT 108.245 179.645 108.575 179.855 ;
        RECT 108.245 179.245 108.455 179.645 ;
        RECT 108.745 179.610 109.155 179.915 ;
        RECT 109.385 179.475 109.555 180.050 ;
        RECT 109.285 179.355 109.555 179.475 ;
        RECT 108.710 179.310 109.555 179.355 ;
        RECT 108.710 179.185 109.465 179.310 ;
        RECT 108.710 179.035 108.880 179.185 ;
        RECT 109.725 179.165 109.895 180.355 ;
        RECT 110.105 179.325 110.310 180.645 ;
        RECT 110.580 180.235 110.830 181.035 ;
        RECT 111.050 180.485 111.380 181.205 ;
        RECT 111.565 180.235 111.815 181.035 ;
        RECT 112.215 180.405 112.545 181.205 ;
        RECT 112.715 180.865 113.050 181.035 ;
        RECT 112.715 180.695 113.055 180.865 ;
        RECT 110.480 180.065 112.535 180.235 ;
        RECT 112.715 180.065 113.050 180.695 ;
        RECT 113.225 180.405 113.555 181.205 ;
        RECT 109.665 179.155 109.895 179.165 ;
        RECT 110.480 179.155 110.650 180.065 ;
        RECT 107.580 178.825 108.880 179.035 ;
        RECT 109.135 178.655 109.465 179.015 ;
        RECT 109.635 178.825 109.895 179.155 ;
        RECT 110.155 178.825 110.650 179.155 ;
        RECT 110.870 178.990 111.225 179.895 ;
        RECT 111.400 179.875 111.570 179.895 ;
        RECT 111.400 178.985 111.700 179.875 ;
        RECT 111.880 178.985 112.140 179.895 ;
        RECT 112.310 179.885 112.535 180.065 ;
        RECT 112.310 179.645 112.705 179.885 ;
        RECT 112.310 178.655 112.545 179.460 ;
        RECT 112.875 179.375 113.050 180.065 ;
        RECT 113.745 180.040 114.035 181.205 ;
        RECT 114.295 180.460 114.565 181.205 ;
        RECT 115.195 181.200 121.470 181.205 ;
        RECT 114.735 180.290 115.025 181.030 ;
        RECT 115.195 180.475 115.450 181.200 ;
        RECT 115.635 180.305 115.895 181.030 ;
        RECT 116.065 180.475 116.310 181.200 ;
        RECT 116.495 180.305 116.755 181.030 ;
        RECT 116.925 180.475 117.170 181.200 ;
        RECT 117.355 180.305 117.615 181.030 ;
        RECT 117.785 180.475 118.030 181.200 ;
        RECT 118.200 180.305 118.460 181.030 ;
        RECT 118.630 180.475 118.890 181.200 ;
        RECT 119.060 180.305 119.320 181.030 ;
        RECT 119.490 180.475 119.750 181.200 ;
        RECT 119.920 180.305 120.180 181.030 ;
        RECT 120.350 180.475 120.610 181.200 ;
        RECT 120.780 180.305 121.040 181.030 ;
        RECT 121.210 180.405 121.470 181.200 ;
        RECT 115.635 180.290 121.040 180.305 ;
        RECT 114.295 180.065 121.040 180.290 ;
        RECT 114.295 179.475 115.460 180.065 ;
        RECT 121.640 179.895 121.890 181.030 ;
        RECT 122.070 180.395 122.330 181.205 ;
        RECT 122.505 179.895 122.750 181.035 ;
        RECT 122.930 180.395 123.225 181.205 ;
        RECT 123.415 180.395 123.710 181.205 ;
        RECT 123.890 179.895 124.135 181.035 ;
        RECT 124.310 180.395 124.570 181.205 ;
        RECT 125.170 181.200 131.445 181.205 ;
        RECT 124.750 179.895 125.000 181.030 ;
        RECT 125.170 180.405 125.430 181.200 ;
        RECT 125.600 180.305 125.860 181.030 ;
        RECT 126.030 180.475 126.290 181.200 ;
        RECT 126.460 180.305 126.720 181.030 ;
        RECT 126.890 180.475 127.150 181.200 ;
        RECT 127.320 180.305 127.580 181.030 ;
        RECT 127.750 180.475 128.010 181.200 ;
        RECT 128.180 180.305 128.440 181.030 ;
        RECT 128.610 180.475 128.855 181.200 ;
        RECT 129.025 180.305 129.285 181.030 ;
        RECT 129.470 180.475 129.715 181.200 ;
        RECT 129.885 180.305 130.145 181.030 ;
        RECT 130.330 180.475 130.575 181.200 ;
        RECT 130.745 180.305 131.005 181.030 ;
        RECT 131.190 180.475 131.445 181.200 ;
        RECT 125.600 180.290 131.005 180.305 ;
        RECT 131.615 180.290 131.905 181.030 ;
        RECT 132.075 180.460 132.345 181.205 ;
        RECT 125.600 180.065 132.345 180.290 ;
        RECT 115.630 179.645 122.750 179.895 ;
        RECT 112.715 178.910 113.050 179.375 ;
        RECT 112.715 178.865 113.045 178.910 ;
        RECT 113.235 178.655 113.565 179.380 ;
        RECT 113.745 178.655 114.035 179.380 ;
        RECT 114.295 179.305 121.040 179.475 ;
        RECT 114.295 178.655 114.595 179.135 ;
        RECT 114.765 178.850 115.025 179.305 ;
        RECT 115.195 178.655 115.455 179.135 ;
        RECT 115.635 178.850 115.895 179.305 ;
        RECT 116.065 178.655 116.315 179.135 ;
        RECT 116.495 178.850 116.755 179.305 ;
        RECT 116.925 178.655 117.175 179.135 ;
        RECT 117.355 178.850 117.615 179.305 ;
        RECT 117.785 178.655 118.030 179.135 ;
        RECT 118.200 178.850 118.475 179.305 ;
        RECT 118.645 178.655 118.890 179.135 ;
        RECT 119.060 178.850 119.320 179.305 ;
        RECT 119.490 178.655 119.750 179.135 ;
        RECT 119.920 178.850 120.180 179.305 ;
        RECT 120.350 178.655 120.610 179.135 ;
        RECT 120.780 178.850 121.040 179.305 ;
        RECT 121.210 178.655 121.470 179.215 ;
        RECT 121.640 178.835 121.890 179.645 ;
        RECT 122.070 178.655 122.330 179.180 ;
        RECT 122.500 178.835 122.750 179.645 ;
        RECT 122.920 179.335 123.235 179.895 ;
        RECT 123.405 179.335 123.720 179.895 ;
        RECT 123.890 179.645 131.010 179.895 ;
        RECT 122.930 178.655 123.235 179.165 ;
        RECT 123.405 178.655 123.710 179.165 ;
        RECT 123.890 178.835 124.140 179.645 ;
        RECT 124.310 178.655 124.570 179.180 ;
        RECT 124.750 178.835 125.000 179.645 ;
        RECT 131.180 179.475 132.345 180.065 ;
        RECT 125.600 179.305 132.345 179.475 ;
        RECT 133.065 180.130 133.335 181.035 ;
        RECT 133.505 180.445 133.835 181.205 ;
        RECT 134.015 180.275 134.185 181.035 ;
        RECT 133.065 179.330 133.235 180.130 ;
        RECT 133.520 180.105 134.185 180.275 ;
        RECT 134.905 180.115 136.115 181.205 ;
        RECT 133.520 179.960 133.690 180.105 ;
        RECT 133.405 179.630 133.690 179.960 ;
        RECT 133.520 179.375 133.690 179.630 ;
        RECT 133.925 179.555 134.255 179.925 ;
        RECT 134.905 179.575 135.425 180.115 ;
        RECT 135.595 179.405 136.115 179.945 ;
        RECT 125.170 178.655 125.430 179.215 ;
        RECT 125.600 178.850 125.860 179.305 ;
        RECT 126.030 178.655 126.290 179.135 ;
        RECT 126.460 178.850 126.720 179.305 ;
        RECT 126.890 178.655 127.150 179.135 ;
        RECT 127.320 178.850 127.580 179.305 ;
        RECT 127.750 178.655 127.995 179.135 ;
        RECT 128.165 178.850 128.440 179.305 ;
        RECT 128.610 178.655 128.855 179.135 ;
        RECT 129.025 178.850 129.285 179.305 ;
        RECT 129.465 178.655 129.715 179.135 ;
        RECT 129.885 178.850 130.145 179.305 ;
        RECT 130.325 178.655 130.575 179.135 ;
        RECT 130.745 178.850 131.005 179.305 ;
        RECT 131.185 178.655 131.445 179.135 ;
        RECT 131.615 178.850 131.875 179.305 ;
        RECT 132.045 178.655 132.345 179.135 ;
        RECT 133.065 178.825 133.325 179.330 ;
        RECT 133.520 179.205 134.185 179.375 ;
        RECT 133.505 178.655 133.835 179.035 ;
        RECT 134.015 178.825 134.185 179.205 ;
        RECT 134.905 178.655 136.115 179.405 ;
        RECT 23.500 178.485 136.200 178.655 ;
        RECT 23.585 177.735 24.795 178.485 ;
        RECT 23.585 177.195 24.105 177.735 ;
        RECT 24.970 177.645 25.230 178.485 ;
        RECT 25.405 177.740 25.660 178.315 ;
        RECT 25.830 178.105 26.160 178.485 ;
        RECT 26.375 177.935 26.545 178.315 ;
        RECT 26.805 177.940 32.150 178.485 ;
        RECT 25.830 177.765 26.545 177.935 ;
        RECT 24.275 177.025 24.795 177.565 ;
        RECT 23.585 175.935 24.795 177.025 ;
        RECT 24.970 175.935 25.230 177.085 ;
        RECT 25.405 177.010 25.575 177.740 ;
        RECT 25.830 177.575 26.000 177.765 ;
        RECT 25.745 177.245 26.000 177.575 ;
        RECT 25.830 177.035 26.000 177.245 ;
        RECT 26.280 177.215 26.635 177.585 ;
        RECT 28.390 177.110 28.730 177.940 ;
        RECT 32.325 177.715 35.835 178.485 ;
        RECT 25.405 176.105 25.660 177.010 ;
        RECT 25.830 176.865 26.545 177.035 ;
        RECT 25.830 175.935 26.160 176.695 ;
        RECT 26.375 176.105 26.545 176.865 ;
        RECT 30.210 176.370 30.560 177.620 ;
        RECT 32.325 177.195 33.975 177.715 ;
        RECT 36.005 177.665 36.265 178.485 ;
        RECT 36.435 177.665 36.765 178.085 ;
        RECT 36.945 178.000 37.735 178.265 ;
        RECT 36.515 177.575 36.765 177.665 ;
        RECT 34.145 177.025 35.835 177.545 ;
        RECT 26.805 175.935 32.150 176.370 ;
        RECT 32.325 175.935 35.835 177.025 ;
        RECT 36.005 176.615 36.345 177.495 ;
        RECT 36.515 177.325 37.310 177.575 ;
        RECT 36.005 175.935 36.265 176.445 ;
        RECT 36.515 176.105 36.685 177.325 ;
        RECT 37.480 177.145 37.735 178.000 ;
        RECT 37.905 177.845 38.105 178.265 ;
        RECT 38.295 178.025 38.625 178.485 ;
        RECT 37.905 177.325 38.315 177.845 ;
        RECT 38.795 177.835 39.055 178.315 ;
        RECT 38.485 177.145 38.715 177.575 ;
        RECT 36.925 176.975 38.715 177.145 ;
        RECT 36.925 176.610 37.175 176.975 ;
        RECT 37.345 176.615 37.675 176.805 ;
        RECT 37.895 176.680 38.610 176.975 ;
        RECT 38.885 176.805 39.055 177.835 ;
        RECT 39.235 177.675 39.505 178.485 ;
        RECT 39.675 177.675 40.005 178.315 ;
        RECT 40.175 177.675 40.415 178.485 ;
        RECT 40.605 177.715 43.195 178.485 ;
        RECT 43.375 177.755 43.675 178.485 ;
        RECT 39.225 177.245 39.575 177.495 ;
        RECT 39.745 177.075 39.915 177.675 ;
        RECT 40.085 177.245 40.435 177.495 ;
        RECT 40.605 177.195 41.815 177.715 ;
        RECT 43.855 177.575 44.085 178.195 ;
        RECT 44.285 177.925 44.510 178.305 ;
        RECT 44.680 178.095 45.010 178.485 ;
        RECT 44.285 177.745 44.615 177.925 ;
        RECT 37.345 176.440 37.540 176.615 ;
        RECT 36.925 175.935 37.540 176.440 ;
        RECT 37.710 176.105 38.185 176.445 ;
        RECT 38.355 175.935 38.570 176.480 ;
        RECT 38.780 176.105 39.055 176.805 ;
        RECT 39.235 175.935 39.565 177.075 ;
        RECT 39.745 176.905 40.425 177.075 ;
        RECT 41.985 177.025 43.195 177.545 ;
        RECT 43.380 177.245 43.675 177.575 ;
        RECT 43.855 177.245 44.270 177.575 ;
        RECT 44.440 177.075 44.615 177.745 ;
        RECT 44.785 177.245 45.025 177.895 ;
        RECT 45.305 177.810 45.545 178.485 ;
        RECT 45.720 177.725 46.275 178.285 ;
        RECT 46.455 177.915 46.660 178.310 ;
        RECT 46.830 178.085 47.175 178.485 ;
        RECT 47.345 177.920 47.675 178.310 ;
        RECT 47.950 178.100 48.625 178.485 ;
        RECT 47.345 177.915 48.565 177.920 ;
        RECT 46.455 177.745 48.565 177.915 ;
        RECT 45.970 177.575 46.275 177.725 ;
        RECT 45.250 177.280 45.750 177.545 ;
        RECT 45.970 177.245 46.355 177.575 ;
        RECT 40.095 176.120 40.425 176.905 ;
        RECT 40.605 175.935 43.195 177.025 ;
        RECT 43.375 176.715 44.270 177.045 ;
        RECT 44.440 176.885 45.025 177.075 ;
        RECT 43.375 176.545 44.580 176.715 ;
        RECT 43.375 176.115 43.705 176.545 ;
        RECT 43.885 175.935 44.080 176.375 ;
        RECT 44.250 176.115 44.580 176.545 ;
        RECT 44.750 176.115 45.025 176.885 ;
        RECT 45.270 176.905 46.400 177.075 ;
        RECT 45.270 176.110 45.540 176.905 ;
        RECT 45.720 175.935 45.935 176.735 ;
        RECT 46.115 176.110 46.400 176.905 ;
        RECT 46.580 176.105 46.860 177.575 ;
        RECT 47.040 176.105 47.370 177.520 ;
        RECT 47.540 177.280 47.970 177.520 ;
        RECT 47.540 176.105 47.745 177.280 ;
        RECT 48.345 177.105 48.565 177.745 ;
        RECT 47.915 176.925 48.565 177.105 ;
        RECT 48.795 176.950 49.125 178.315 ;
        RECT 49.345 177.760 49.635 178.485 ;
        RECT 49.830 178.095 50.160 178.485 ;
        RECT 50.330 177.925 50.555 178.305 ;
        RECT 49.815 177.245 50.055 177.895 ;
        RECT 50.225 177.745 50.555 177.925 ;
        RECT 47.915 176.110 48.125 176.925 ;
        RECT 48.365 175.935 48.695 176.755 ;
        RECT 48.870 176.110 49.125 176.950 ;
        RECT 49.345 175.935 49.635 177.100 ;
        RECT 50.225 177.075 50.400 177.745 ;
        RECT 50.755 177.575 50.985 178.195 ;
        RECT 51.165 177.755 51.465 178.485 ;
        RECT 51.665 177.675 51.905 178.485 ;
        RECT 52.075 177.675 52.405 178.315 ;
        RECT 52.575 177.675 52.845 178.485 ;
        RECT 53.025 177.940 58.370 178.485 ;
        RECT 50.570 177.245 50.985 177.575 ;
        RECT 51.165 177.245 51.460 177.575 ;
        RECT 51.645 177.245 51.995 177.495 ;
        RECT 52.165 177.075 52.335 177.675 ;
        RECT 52.505 177.245 52.855 177.495 ;
        RECT 54.610 177.110 54.950 177.940 ;
        RECT 58.545 177.715 60.215 178.485 ;
        RECT 60.850 177.980 61.185 178.485 ;
        RECT 61.355 177.915 61.595 178.290 ;
        RECT 61.875 178.155 62.045 178.300 ;
        RECT 61.875 177.960 62.250 178.155 ;
        RECT 62.610 177.990 63.005 178.485 ;
        RECT 49.815 176.885 50.400 177.075 ;
        RECT 49.815 176.115 50.090 176.885 ;
        RECT 50.570 176.715 51.465 177.045 ;
        RECT 50.260 176.545 51.465 176.715 ;
        RECT 50.260 176.115 50.590 176.545 ;
        RECT 50.760 175.935 50.955 176.375 ;
        RECT 51.135 176.115 51.465 176.545 ;
        RECT 51.655 176.905 52.335 177.075 ;
        RECT 51.655 176.120 51.985 176.905 ;
        RECT 52.515 175.935 52.845 177.075 ;
        RECT 56.430 176.370 56.780 177.620 ;
        RECT 58.545 177.195 59.295 177.715 ;
        RECT 59.465 177.025 60.215 177.545 ;
        RECT 53.025 175.935 58.370 176.370 ;
        RECT 58.545 175.935 60.215 177.025 ;
        RECT 60.905 176.955 61.205 177.805 ;
        RECT 61.375 177.765 61.595 177.915 ;
        RECT 61.375 177.435 61.910 177.765 ;
        RECT 62.080 177.625 62.250 177.960 ;
        RECT 63.175 177.795 63.415 178.315 ;
        RECT 61.375 176.785 61.610 177.435 ;
        RECT 62.080 177.265 63.065 177.625 ;
        RECT 60.935 176.555 61.610 176.785 ;
        RECT 61.780 177.245 63.065 177.265 ;
        RECT 61.780 177.095 62.640 177.245 ;
        RECT 60.935 176.125 61.105 176.555 ;
        RECT 61.275 175.935 61.605 176.385 ;
        RECT 61.780 176.150 62.065 177.095 ;
        RECT 63.240 176.990 63.415 177.795 ;
        RECT 62.240 176.615 62.935 176.925 ;
        RECT 62.245 175.935 62.930 176.405 ;
        RECT 63.110 176.205 63.415 176.990 ;
        RECT 63.605 177.760 63.865 178.315 ;
        RECT 64.035 178.040 64.465 178.485 ;
        RECT 64.700 177.915 64.870 178.315 ;
        RECT 65.040 178.085 65.760 178.485 ;
        RECT 63.605 177.045 63.780 177.760 ;
        RECT 64.700 177.745 65.580 177.915 ;
        RECT 65.930 177.870 66.100 178.315 ;
        RECT 66.675 177.975 67.075 178.485 ;
        RECT 67.285 177.940 72.630 178.485 ;
        RECT 63.950 177.245 64.205 177.575 ;
        RECT 63.605 176.105 63.865 177.045 ;
        RECT 64.035 176.765 64.205 177.245 ;
        RECT 64.430 176.955 64.760 177.575 ;
        RECT 64.930 177.195 65.220 177.575 ;
        RECT 65.410 177.025 65.580 177.745 ;
        RECT 65.060 176.855 65.580 177.025 ;
        RECT 65.750 177.700 66.100 177.870 ;
        RECT 64.035 176.595 64.795 176.765 ;
        RECT 65.060 176.665 65.230 176.855 ;
        RECT 65.750 176.675 65.920 177.700 ;
        RECT 66.340 177.215 66.600 177.805 ;
        RECT 66.120 176.915 66.600 177.215 ;
        RECT 66.800 176.915 67.060 177.805 ;
        RECT 68.870 177.110 69.210 177.940 ;
        RECT 72.805 177.715 74.475 178.485 ;
        RECT 75.105 177.760 75.395 178.485 ;
        RECT 75.565 177.715 79.075 178.485 ;
        RECT 80.625 178.105 80.955 178.485 ;
        RECT 80.180 177.935 80.455 178.075 ;
        RECT 81.125 177.935 81.335 178.105 ;
        RECT 80.180 177.745 81.335 177.935 ;
        RECT 81.505 177.935 81.835 178.315 ;
        RECT 82.025 178.105 82.355 178.485 ;
        RECT 81.505 177.730 82.355 177.935 ;
        RECT 64.625 176.370 64.795 176.595 ;
        RECT 65.510 176.505 65.920 176.675 ;
        RECT 66.095 176.565 67.035 176.735 ;
        RECT 65.510 176.370 65.765 176.505 ;
        RECT 64.035 175.935 64.365 176.335 ;
        RECT 64.625 176.200 65.765 176.370 ;
        RECT 66.095 176.315 66.265 176.565 ;
        RECT 65.510 176.105 65.765 176.200 ;
        RECT 65.935 176.145 66.265 176.315 ;
        RECT 66.435 175.935 66.685 176.395 ;
        RECT 66.855 176.105 67.035 176.565 ;
        RECT 70.690 176.370 71.040 177.620 ;
        RECT 72.805 177.195 73.555 177.715 ;
        RECT 73.725 177.025 74.475 177.545 ;
        RECT 75.565 177.195 77.215 177.715 ;
        RECT 67.285 175.935 72.630 176.370 ;
        RECT 72.805 175.935 74.475 177.025 ;
        RECT 75.105 175.935 75.395 177.100 ;
        RECT 77.385 177.025 79.075 177.545 ;
        RECT 80.175 177.120 80.435 177.575 ;
        RECT 80.690 177.170 81.275 177.545 ;
        RECT 75.565 175.935 79.075 177.025 ;
        RECT 80.180 175.935 80.505 176.920 ;
        RECT 80.690 176.785 80.895 177.170 ;
        RECT 81.445 176.955 81.855 177.560 ;
        RECT 82.025 177.240 82.355 177.730 ;
        RECT 82.025 176.785 82.195 177.240 ;
        RECT 80.685 176.615 80.895 176.785 ;
        RECT 80.690 176.585 80.895 176.615 ;
        RECT 81.075 176.565 82.195 176.785 ;
        RECT 81.075 176.105 81.335 176.565 ;
        RECT 81.505 175.935 82.355 176.385 ;
        RECT 82.525 176.105 82.770 178.315 ;
        RECT 82.955 177.685 83.195 178.485 ;
        RECT 83.475 178.005 83.775 178.485 ;
        RECT 83.945 177.835 84.205 178.290 ;
        RECT 84.375 178.005 84.635 178.485 ;
        RECT 84.815 177.835 85.075 178.290 ;
        RECT 85.245 178.005 85.495 178.485 ;
        RECT 85.675 177.835 85.935 178.290 ;
        RECT 86.105 178.005 86.355 178.485 ;
        RECT 86.535 177.835 86.795 178.290 ;
        RECT 86.965 178.005 87.210 178.485 ;
        RECT 87.380 177.835 87.655 178.290 ;
        RECT 87.825 178.005 88.070 178.485 ;
        RECT 88.240 177.835 88.500 178.290 ;
        RECT 88.670 178.005 88.930 178.485 ;
        RECT 89.100 177.835 89.360 178.290 ;
        RECT 89.530 178.005 89.790 178.485 ;
        RECT 89.960 177.835 90.220 178.290 ;
        RECT 90.390 177.925 90.650 178.485 ;
        RECT 83.475 177.805 90.220 177.835 ;
        RECT 83.445 177.665 90.220 177.805 ;
        RECT 83.445 177.635 84.640 177.665 ;
        RECT 83.475 177.075 84.640 177.635 ;
        RECT 90.820 177.495 91.070 178.305 ;
        RECT 91.250 177.960 91.510 178.485 ;
        RECT 91.680 177.495 91.930 178.305 ;
        RECT 92.110 177.975 92.415 178.485 ;
        RECT 92.585 177.985 92.845 178.315 ;
        RECT 93.015 178.125 93.345 178.485 ;
        RECT 93.600 178.105 94.900 178.315 ;
        RECT 92.585 177.975 92.815 177.985 ;
        RECT 84.810 177.245 91.930 177.495 ;
        RECT 92.100 177.245 92.415 177.805 ;
        RECT 82.955 175.935 83.210 176.935 ;
        RECT 83.475 176.850 90.220 177.075 ;
        RECT 83.475 175.935 83.745 176.680 ;
        RECT 83.915 176.110 84.205 176.850 ;
        RECT 84.815 176.835 90.220 176.850 ;
        RECT 84.375 175.940 84.630 176.665 ;
        RECT 84.815 176.110 85.075 176.835 ;
        RECT 85.245 175.940 85.490 176.665 ;
        RECT 85.675 176.110 85.935 176.835 ;
        RECT 86.105 175.940 86.350 176.665 ;
        RECT 86.535 176.110 86.795 176.835 ;
        RECT 86.965 175.940 87.210 176.665 ;
        RECT 87.380 176.110 87.640 176.835 ;
        RECT 87.810 175.940 88.070 176.665 ;
        RECT 88.240 176.110 88.500 176.835 ;
        RECT 88.670 175.940 88.930 176.665 ;
        RECT 89.100 176.110 89.360 176.835 ;
        RECT 89.530 175.940 89.790 176.665 ;
        RECT 89.960 176.110 90.220 176.835 ;
        RECT 90.390 175.940 90.650 176.735 ;
        RECT 90.820 176.110 91.070 177.245 ;
        RECT 84.375 175.935 90.650 175.940 ;
        RECT 91.250 175.935 91.510 176.745 ;
        RECT 91.685 176.105 91.930 177.245 ;
        RECT 92.585 176.785 92.755 177.975 ;
        RECT 93.600 177.955 93.770 178.105 ;
        RECT 93.015 177.830 93.770 177.955 ;
        RECT 92.925 177.785 93.770 177.830 ;
        RECT 92.925 177.665 93.195 177.785 ;
        RECT 92.925 177.090 93.095 177.665 ;
        RECT 93.325 177.225 93.735 177.530 ;
        RECT 94.025 177.495 94.235 177.895 ;
        RECT 93.905 177.285 94.235 177.495 ;
        RECT 94.480 177.495 94.700 177.895 ;
        RECT 95.175 177.720 95.630 178.485 ;
        RECT 95.840 177.745 96.455 178.315 ;
        RECT 96.625 177.975 96.840 178.485 ;
        RECT 97.070 177.975 97.350 178.305 ;
        RECT 97.530 177.975 97.770 178.485 ;
        RECT 94.480 177.285 94.955 177.495 ;
        RECT 95.145 177.295 95.635 177.495 ;
        RECT 92.925 177.055 93.125 177.090 ;
        RECT 94.455 177.055 95.630 177.115 ;
        RECT 92.925 176.945 95.630 177.055 ;
        RECT 92.985 176.885 94.785 176.945 ;
        RECT 94.455 176.855 94.785 176.885 ;
        RECT 92.110 175.935 92.405 176.745 ;
        RECT 92.585 176.105 92.845 176.785 ;
        RECT 93.015 175.935 93.265 176.715 ;
        RECT 93.515 176.685 94.350 176.695 ;
        RECT 94.940 176.685 95.125 176.775 ;
        RECT 93.515 176.485 95.125 176.685 ;
        RECT 93.515 176.105 93.765 176.485 ;
        RECT 94.895 176.445 95.125 176.485 ;
        RECT 95.375 176.325 95.630 176.945 ;
        RECT 93.935 175.935 94.290 176.315 ;
        RECT 95.295 176.105 95.630 176.325 ;
        RECT 95.840 176.725 96.155 177.745 ;
        RECT 96.325 177.075 96.495 177.575 ;
        RECT 96.745 177.245 97.010 177.805 ;
        RECT 97.180 177.075 97.350 177.975 ;
        RECT 98.105 177.810 98.365 178.315 ;
        RECT 98.545 178.105 98.875 178.485 ;
        RECT 99.055 177.935 99.225 178.315 ;
        RECT 97.520 177.245 97.875 177.805 ;
        RECT 96.325 176.905 97.750 177.075 ;
        RECT 95.840 176.105 96.375 176.725 ;
        RECT 96.545 175.935 96.875 176.735 ;
        RECT 97.360 176.730 97.750 176.905 ;
        RECT 98.105 177.010 98.285 177.810 ;
        RECT 98.560 177.765 99.225 177.935 ;
        RECT 98.560 177.510 98.730 177.765 ;
        RECT 99.545 177.665 99.755 178.485 ;
        RECT 99.925 177.685 100.255 178.315 ;
        RECT 98.455 177.180 98.730 177.510 ;
        RECT 98.955 177.215 99.295 177.585 ;
        RECT 98.560 177.035 98.730 177.180 ;
        RECT 99.925 177.085 100.175 177.685 ;
        RECT 100.425 177.665 100.655 178.485 ;
        RECT 100.865 177.760 101.155 178.485 ;
        RECT 101.330 178.085 101.665 178.485 ;
        RECT 101.835 177.915 102.040 178.315 ;
        RECT 102.250 178.005 102.525 178.485 ;
        RECT 102.735 177.985 102.995 178.315 ;
        RECT 101.355 177.745 102.040 177.915 ;
        RECT 100.345 177.245 100.675 177.495 ;
        RECT 98.105 176.105 98.375 177.010 ;
        RECT 98.560 176.865 99.235 177.035 ;
        RECT 98.545 175.935 98.875 176.695 ;
        RECT 99.055 176.105 99.235 176.865 ;
        RECT 99.545 175.935 99.755 177.075 ;
        RECT 99.925 176.105 100.255 177.085 ;
        RECT 100.425 175.935 100.655 177.075 ;
        RECT 100.865 175.935 101.155 177.100 ;
        RECT 101.355 176.715 101.695 177.745 ;
        RECT 101.865 177.075 102.115 177.575 ;
        RECT 102.295 177.245 102.655 177.825 ;
        RECT 102.825 177.075 102.995 177.985 ;
        RECT 103.165 177.875 103.505 178.290 ;
        RECT 103.675 178.045 103.845 178.485 ;
        RECT 104.015 178.095 105.265 178.275 ;
        RECT 104.015 177.875 104.345 178.095 ;
        RECT 105.535 178.025 105.705 178.485 ;
        RECT 103.165 177.705 104.345 177.875 ;
        RECT 104.515 177.855 104.880 177.925 ;
        RECT 104.515 177.675 105.765 177.855 ;
        RECT 103.165 177.295 103.630 177.495 ;
        RECT 103.805 177.245 104.135 177.495 ;
        RECT 104.305 177.465 104.770 177.495 ;
        RECT 104.305 177.295 104.775 177.465 ;
        RECT 104.305 177.245 104.770 177.295 ;
        RECT 104.965 177.245 105.320 177.495 ;
        RECT 103.805 177.125 103.985 177.245 ;
        RECT 101.865 176.905 102.995 177.075 ;
        RECT 101.355 176.540 102.020 176.715 ;
        RECT 101.330 175.935 101.665 176.360 ;
        RECT 101.835 176.135 102.020 176.540 ;
        RECT 102.225 175.935 102.555 176.715 ;
        RECT 102.725 176.135 102.995 176.905 ;
        RECT 103.165 175.935 103.485 177.115 ;
        RECT 103.655 176.955 103.985 177.125 ;
        RECT 105.490 177.075 105.765 177.675 ;
        RECT 103.655 176.165 103.855 176.955 ;
        RECT 104.155 176.865 105.765 177.075 ;
        RECT 104.155 176.765 104.565 176.865 ;
        RECT 104.180 176.105 104.565 176.765 ;
        RECT 104.960 175.935 105.745 176.695 ;
        RECT 105.935 176.105 106.215 178.205 ;
        RECT 106.385 177.975 106.690 178.485 ;
        RECT 106.385 177.245 106.700 177.805 ;
        RECT 106.870 177.495 107.120 178.305 ;
        RECT 107.290 177.960 107.550 178.485 ;
        RECT 107.730 177.495 107.980 178.305 ;
        RECT 108.150 177.925 108.410 178.485 ;
        RECT 108.580 177.835 108.840 178.290 ;
        RECT 109.010 178.005 109.270 178.485 ;
        RECT 109.440 177.835 109.700 178.290 ;
        RECT 109.870 178.005 110.130 178.485 ;
        RECT 110.300 177.835 110.560 178.290 ;
        RECT 110.730 178.005 110.975 178.485 ;
        RECT 111.145 177.835 111.420 178.290 ;
        RECT 111.590 178.005 111.835 178.485 ;
        RECT 112.005 177.835 112.265 178.290 ;
        RECT 112.445 178.005 112.695 178.485 ;
        RECT 112.865 177.835 113.125 178.290 ;
        RECT 113.305 178.005 113.555 178.485 ;
        RECT 113.725 177.835 113.985 178.290 ;
        RECT 114.165 178.005 114.425 178.485 ;
        RECT 114.595 177.835 114.855 178.290 ;
        RECT 115.025 178.005 115.325 178.485 ;
        RECT 108.580 177.665 115.325 177.835 ;
        RECT 115.595 177.675 115.865 178.485 ;
        RECT 116.035 177.675 116.365 178.315 ;
        RECT 116.535 177.675 116.775 178.485 ;
        RECT 116.965 177.715 120.475 178.485 ;
        RECT 106.870 177.245 113.990 177.495 ;
        RECT 106.395 175.935 106.690 176.745 ;
        RECT 106.870 176.105 107.115 177.245 ;
        RECT 107.290 175.935 107.550 176.745 ;
        RECT 107.730 176.110 107.980 177.245 ;
        RECT 114.160 177.075 115.325 177.665 ;
        RECT 115.585 177.245 115.935 177.495 ;
        RECT 116.105 177.075 116.275 177.675 ;
        RECT 116.445 177.245 116.795 177.495 ;
        RECT 116.965 177.195 118.615 177.715 ;
        RECT 121.105 177.685 121.415 178.485 ;
        RECT 121.620 177.685 122.315 178.315 ;
        RECT 122.575 177.935 122.745 178.315 ;
        RECT 122.925 178.105 123.255 178.485 ;
        RECT 122.575 177.765 123.240 177.935 ;
        RECT 123.435 177.810 123.695 178.315 ;
        RECT 108.580 176.850 115.325 177.075 ;
        RECT 108.580 176.835 113.985 176.850 ;
        RECT 108.150 175.940 108.410 176.735 ;
        RECT 108.580 176.110 108.840 176.835 ;
        RECT 109.010 175.940 109.270 176.665 ;
        RECT 109.440 176.110 109.700 176.835 ;
        RECT 109.870 175.940 110.130 176.665 ;
        RECT 110.300 176.110 110.560 176.835 ;
        RECT 110.730 175.940 110.990 176.665 ;
        RECT 111.160 176.110 111.420 176.835 ;
        RECT 111.590 175.940 111.835 176.665 ;
        RECT 112.005 176.110 112.265 176.835 ;
        RECT 112.450 175.940 112.695 176.665 ;
        RECT 112.865 176.110 113.125 176.835 ;
        RECT 113.310 175.940 113.555 176.665 ;
        RECT 113.725 176.110 113.985 176.835 ;
        RECT 114.170 175.940 114.425 176.665 ;
        RECT 114.595 176.110 114.885 176.850 ;
        RECT 108.150 175.935 114.425 175.940 ;
        RECT 115.055 175.935 115.325 176.680 ;
        RECT 115.595 175.935 115.925 177.075 ;
        RECT 116.105 176.905 116.785 177.075 ;
        RECT 118.785 177.025 120.475 177.545 ;
        RECT 121.115 177.245 121.450 177.515 ;
        RECT 121.620 177.085 121.790 177.685 ;
        RECT 121.960 177.245 122.295 177.495 ;
        RECT 122.505 177.215 122.835 177.585 ;
        RECT 123.070 177.510 123.240 177.765 ;
        RECT 123.070 177.180 123.355 177.510 ;
        RECT 116.455 176.120 116.785 176.905 ;
        RECT 116.965 175.935 120.475 177.025 ;
        RECT 121.105 175.935 121.385 177.075 ;
        RECT 121.555 176.105 121.885 177.085 ;
        RECT 122.055 175.935 122.315 177.075 ;
        RECT 123.070 177.035 123.240 177.180 ;
        RECT 122.575 176.865 123.240 177.035 ;
        RECT 123.525 177.010 123.695 177.810 ;
        RECT 122.575 176.105 122.745 176.865 ;
        RECT 122.925 175.935 123.255 176.695 ;
        RECT 123.425 176.105 123.695 177.010 ;
        RECT 123.865 177.985 124.165 178.315 ;
        RECT 124.335 178.005 124.610 178.485 ;
        RECT 123.865 177.075 124.035 177.985 ;
        RECT 124.790 177.835 125.085 178.225 ;
        RECT 125.255 178.005 125.510 178.485 ;
        RECT 125.685 177.835 125.945 178.225 ;
        RECT 126.115 178.005 126.395 178.485 ;
        RECT 124.205 177.245 124.555 177.815 ;
        RECT 124.790 177.665 126.440 177.835 ;
        RECT 126.625 177.760 126.915 178.485 ;
        RECT 127.090 177.685 127.345 178.485 ;
        RECT 124.725 177.325 125.865 177.495 ;
        RECT 124.725 177.075 124.895 177.325 ;
        RECT 126.035 177.155 126.440 177.665 ;
        RECT 123.865 176.905 124.895 177.075 ;
        RECT 125.685 176.985 126.440 177.155 ;
        RECT 123.865 176.105 124.175 176.905 ;
        RECT 125.685 176.735 125.945 176.985 ;
        RECT 124.345 175.935 124.655 176.735 ;
        RECT 124.825 176.565 125.945 176.735 ;
        RECT 124.825 176.105 125.085 176.565 ;
        RECT 125.255 175.935 125.510 176.395 ;
        RECT 125.685 176.105 125.945 176.565 ;
        RECT 126.115 175.935 126.400 176.805 ;
        RECT 126.625 175.935 126.915 177.100 ;
        RECT 127.090 175.935 127.345 177.075 ;
        RECT 127.515 176.145 127.845 178.275 ;
        RECT 128.015 178.105 128.345 178.485 ;
        RECT 128.525 178.145 129.960 178.315 ;
        RECT 128.525 177.915 128.695 178.145 ;
        RECT 128.015 177.745 128.695 177.915 ;
        RECT 128.015 177.075 128.185 177.745 ;
        RECT 128.495 177.245 128.710 177.575 ;
        RECT 128.895 177.245 129.165 177.965 ;
        RECT 129.440 177.575 129.620 177.965 ;
        RECT 129.790 177.915 129.960 178.145 ;
        RECT 130.220 178.085 130.550 178.485 ;
        RECT 130.795 177.915 130.965 178.315 ;
        RECT 129.790 177.745 130.965 177.915 ;
        RECT 131.225 177.745 131.710 178.315 ;
        RECT 131.880 177.915 132.110 178.315 ;
        RECT 132.280 178.085 132.700 178.485 ;
        RECT 132.870 177.915 133.040 178.315 ;
        RECT 131.880 177.745 133.040 177.915 ;
        RECT 133.210 177.745 133.660 178.485 ;
        RECT 133.830 177.745 134.270 178.305 ;
        RECT 129.440 177.245 129.675 177.575 ;
        RECT 129.895 177.245 130.235 177.575 ;
        RECT 130.695 177.245 131.005 177.575 ;
        RECT 131.225 177.075 131.395 177.745 ;
        RECT 131.565 177.245 131.965 177.575 ;
        RECT 128.015 176.905 130.965 177.075 ;
        RECT 131.225 176.905 131.990 177.075 ;
        RECT 128.160 175.935 128.380 176.735 ;
        RECT 128.590 176.565 130.025 176.735 ;
        RECT 128.590 176.105 128.840 176.565 ;
        RECT 129.125 175.935 129.455 176.315 ;
        RECT 129.715 176.105 130.025 176.565 ;
        RECT 130.795 176.105 130.965 176.905 ;
        RECT 131.230 175.935 131.565 176.735 ;
        RECT 131.740 176.275 131.990 176.905 ;
        RECT 132.180 176.445 132.430 177.575 ;
        RECT 132.630 177.245 132.875 177.575 ;
        RECT 133.060 177.295 133.450 177.575 ;
        RECT 132.630 176.445 132.830 177.245 ;
        RECT 133.620 177.125 133.790 177.575 ;
        RECT 133.000 176.955 133.790 177.125 ;
        RECT 133.960 177.495 134.270 177.745 ;
        RECT 134.440 177.665 134.735 178.485 ;
        RECT 134.905 177.735 136.115 178.485 ;
        RECT 133.960 177.275 134.735 177.495 ;
        RECT 133.000 176.275 133.170 176.955 ;
        RECT 131.740 176.105 133.170 176.275 ;
        RECT 133.340 175.935 133.655 176.785 ;
        RECT 133.960 176.735 134.270 177.275 ;
        RECT 133.830 176.105 134.270 176.735 ;
        RECT 134.440 175.935 134.735 177.105 ;
        RECT 134.905 177.025 135.425 177.565 ;
        RECT 135.595 177.195 136.115 177.735 ;
        RECT 134.905 175.935 136.115 177.025 ;
        RECT 23.500 175.765 136.200 175.935 ;
        RECT 23.585 174.675 24.795 175.765 ;
        RECT 24.965 174.675 26.175 175.765 ;
        RECT 23.585 173.965 24.105 174.505 ;
        RECT 24.275 174.135 24.795 174.675 ;
        RECT 24.965 173.965 25.485 174.505 ;
        RECT 25.655 174.135 26.175 174.675 ;
        RECT 26.385 174.625 26.615 175.765 ;
        RECT 26.785 174.615 27.115 175.595 ;
        RECT 27.285 174.625 27.495 175.765 ;
        RECT 27.815 175.145 27.985 175.575 ;
        RECT 28.155 175.315 28.485 175.765 ;
        RECT 27.815 174.915 28.495 175.145 ;
        RECT 26.365 174.205 26.695 174.455 ;
        RECT 23.585 173.215 24.795 173.965 ;
        RECT 24.965 173.215 26.175 173.965 ;
        RECT 26.385 173.215 26.615 174.035 ;
        RECT 26.865 174.015 27.115 174.615 ;
        RECT 27.785 174.575 28.090 174.745 ;
        RECT 26.785 173.385 27.115 174.015 ;
        RECT 27.285 173.215 27.495 174.035 ;
        RECT 27.790 173.895 28.090 174.575 ;
        RECT 28.260 174.265 28.495 174.915 ;
        RECT 28.685 174.605 28.970 175.550 ;
        RECT 29.150 175.295 29.835 175.765 ;
        RECT 29.145 174.775 29.840 175.085 ;
        RECT 30.015 174.710 30.320 175.495 ;
        RECT 30.505 174.810 30.775 175.765 ;
        RECT 31.035 175.145 31.205 175.575 ;
        RECT 31.375 175.315 31.705 175.765 ;
        RECT 31.035 174.915 31.710 175.145 ;
        RECT 28.685 174.455 29.545 174.605 ;
        RECT 28.685 174.435 29.975 174.455 ;
        RECT 28.260 173.935 28.815 174.265 ;
        RECT 28.985 174.075 29.975 174.435 ;
        RECT 28.260 173.785 28.475 173.935 ;
        RECT 27.735 173.215 28.065 173.720 ;
        RECT 28.235 173.410 28.475 173.785 ;
        RECT 28.985 173.740 29.155 174.075 ;
        RECT 30.145 173.905 30.320 174.710 ;
        RECT 28.755 173.545 29.155 173.740 ;
        RECT 28.755 173.400 28.925 173.545 ;
        RECT 29.515 173.215 29.915 173.710 ;
        RECT 30.085 173.385 30.320 173.905 ;
        RECT 31.005 173.895 31.305 174.745 ;
        RECT 31.475 174.265 31.710 174.915 ;
        RECT 31.880 174.605 32.165 175.550 ;
        RECT 32.345 175.295 33.030 175.765 ;
        RECT 32.340 174.775 33.035 175.085 ;
        RECT 33.210 174.710 33.515 175.495 ;
        RECT 33.905 175.095 34.185 175.765 ;
        RECT 31.880 174.455 32.740 174.605 ;
        RECT 31.880 174.435 33.165 174.455 ;
        RECT 31.475 173.935 32.010 174.265 ;
        RECT 32.180 174.075 33.165 174.435 ;
        RECT 30.505 173.215 30.775 173.850 ;
        RECT 31.475 173.785 31.695 173.935 ;
        RECT 30.950 173.215 31.285 173.720 ;
        RECT 31.455 173.410 31.695 173.785 ;
        RECT 32.180 173.740 32.350 174.075 ;
        RECT 33.340 173.905 33.515 174.710 ;
        RECT 33.705 174.455 34.020 174.895 ;
        RECT 34.355 174.875 34.655 175.425 ;
        RECT 34.865 175.045 35.195 175.765 ;
        RECT 35.385 175.045 35.835 175.595 ;
        RECT 34.355 174.705 35.295 174.875 ;
        RECT 35.125 174.455 35.295 174.705 ;
        RECT 33.705 174.205 34.395 174.455 ;
        RECT 34.625 174.205 34.955 174.455 ;
        RECT 35.125 174.125 35.415 174.455 ;
        RECT 35.125 174.035 35.295 174.125 ;
        RECT 31.975 173.545 32.350 173.740 ;
        RECT 31.975 173.400 32.145 173.545 ;
        RECT 32.710 173.215 33.105 173.710 ;
        RECT 33.275 173.385 33.515 173.905 ;
        RECT 33.905 173.845 35.295 174.035 ;
        RECT 33.905 173.485 34.235 173.845 ;
        RECT 35.585 173.675 35.835 175.045 ;
        RECT 36.005 174.625 36.295 175.765 ;
        RECT 36.465 174.600 36.755 175.765 ;
        RECT 37.010 175.145 37.185 175.595 ;
        RECT 37.355 175.325 37.685 175.765 ;
        RECT 37.990 175.175 38.160 175.595 ;
        RECT 38.395 175.355 39.065 175.765 ;
        RECT 39.280 175.175 39.450 175.595 ;
        RECT 39.650 175.355 39.980 175.765 ;
        RECT 37.010 174.975 37.640 175.145 ;
        RECT 36.925 174.125 37.290 174.805 ;
        RECT 37.470 174.455 37.640 174.975 ;
        RECT 37.990 175.005 40.005 175.175 ;
        RECT 37.470 174.125 37.820 174.455 ;
        RECT 34.865 173.215 35.115 173.675 ;
        RECT 35.285 173.385 35.835 173.675 ;
        RECT 36.005 173.215 36.295 174.015 ;
        RECT 37.470 173.955 37.640 174.125 ;
        RECT 36.465 173.215 36.755 173.940 ;
        RECT 37.010 173.785 37.640 173.955 ;
        RECT 37.010 173.385 37.185 173.785 ;
        RECT 37.990 173.715 38.160 175.005 ;
        RECT 37.355 173.215 37.685 173.595 ;
        RECT 37.930 173.385 38.160 173.715 ;
        RECT 38.360 173.550 38.640 174.825 ;
        RECT 38.865 173.725 39.135 174.825 ;
        RECT 39.325 173.795 39.665 174.825 ;
        RECT 39.835 174.455 40.005 175.005 ;
        RECT 40.175 174.625 40.435 175.595 ;
        RECT 40.605 174.675 44.115 175.765 ;
        RECT 39.835 174.125 40.095 174.455 ;
        RECT 40.265 173.935 40.435 174.625 ;
        RECT 38.825 173.555 39.135 173.725 ;
        RECT 38.865 173.550 39.135 173.555 ;
        RECT 39.595 173.215 39.925 173.595 ;
        RECT 40.095 173.470 40.435 173.935 ;
        RECT 40.605 173.985 42.255 174.505 ;
        RECT 42.425 174.155 44.115 174.675 ;
        RECT 44.500 174.665 44.830 175.765 ;
        RECT 45.305 175.165 45.630 175.595 ;
        RECT 45.800 175.345 46.130 175.765 ;
        RECT 46.875 175.335 47.285 175.765 ;
        RECT 45.305 174.995 47.285 175.165 ;
        RECT 45.305 174.585 46.010 174.995 ;
        RECT 44.285 174.205 44.930 174.415 ;
        RECT 45.100 174.205 45.670 174.415 ;
        RECT 40.095 173.425 40.430 173.470 ;
        RECT 40.605 173.215 44.115 173.985 ;
        RECT 44.440 173.865 45.610 174.035 ;
        RECT 44.440 173.400 44.770 173.865 ;
        RECT 44.940 173.215 45.110 173.685 ;
        RECT 45.280 173.385 45.610 173.865 ;
        RECT 45.840 173.385 46.010 174.585 ;
        RECT 46.180 174.655 46.805 174.825 ;
        RECT 46.180 173.955 46.350 174.655 ;
        RECT 47.020 174.455 47.285 174.995 ;
        RECT 47.455 174.610 47.795 175.595 ;
        RECT 48.895 175.155 49.225 175.585 ;
        RECT 49.405 175.325 49.600 175.765 ;
        RECT 49.770 175.155 50.100 175.585 ;
        RECT 48.895 174.985 50.100 175.155 ;
        RECT 48.895 174.655 49.790 174.985 ;
        RECT 50.270 174.815 50.545 175.585 ;
        RECT 50.725 175.330 56.070 175.765 ;
        RECT 46.520 174.125 46.850 174.455 ;
        RECT 47.020 174.125 47.370 174.455 ;
        RECT 47.540 173.955 47.795 174.610 ;
        RECT 49.960 174.625 50.545 174.815 ;
        RECT 48.900 174.125 49.195 174.455 ;
        RECT 49.375 174.125 49.790 174.455 ;
        RECT 46.180 173.785 46.720 173.955 ;
        RECT 46.550 173.580 46.720 173.785 ;
        RECT 47.000 173.215 47.170 173.955 ;
        RECT 47.435 173.580 47.795 173.955 ;
        RECT 48.895 173.215 49.195 173.945 ;
        RECT 49.375 173.505 49.605 174.125 ;
        RECT 49.960 173.955 50.135 174.625 ;
        RECT 49.805 173.775 50.135 173.955 ;
        RECT 50.305 173.805 50.545 174.455 ;
        RECT 49.805 173.395 50.030 173.775 ;
        RECT 52.310 173.760 52.650 174.590 ;
        RECT 54.130 174.080 54.480 175.330 ;
        RECT 56.745 174.625 56.975 175.765 ;
        RECT 57.145 174.615 57.475 175.595 ;
        RECT 57.645 174.625 57.855 175.765 ;
        RECT 58.085 174.675 61.595 175.765 ;
        RECT 56.725 174.205 57.055 174.455 ;
        RECT 50.200 173.215 50.530 173.605 ;
        RECT 50.725 173.215 56.070 173.760 ;
        RECT 56.745 173.215 56.975 174.035 ;
        RECT 57.225 174.015 57.475 174.615 ;
        RECT 57.145 173.385 57.475 174.015 ;
        RECT 57.645 173.215 57.855 174.035 ;
        RECT 58.085 173.985 59.735 174.505 ;
        RECT 59.905 174.155 61.595 174.675 ;
        RECT 62.225 174.600 62.515 175.765 ;
        RECT 62.775 175.145 62.945 175.575 ;
        RECT 63.115 175.315 63.445 175.765 ;
        RECT 62.775 174.915 63.450 175.145 ;
        RECT 58.085 173.215 61.595 173.985 ;
        RECT 62.225 173.215 62.515 173.940 ;
        RECT 62.745 173.895 63.045 174.745 ;
        RECT 63.215 174.265 63.450 174.915 ;
        RECT 63.620 174.605 63.905 175.550 ;
        RECT 64.085 175.295 64.770 175.765 ;
        RECT 64.080 174.775 64.775 175.085 ;
        RECT 64.950 174.710 65.255 175.495 ;
        RECT 63.620 174.455 64.480 174.605 ;
        RECT 63.620 174.435 64.905 174.455 ;
        RECT 63.215 173.935 63.750 174.265 ;
        RECT 63.920 174.075 64.905 174.435 ;
        RECT 63.215 173.785 63.435 173.935 ;
        RECT 62.690 173.215 63.025 173.720 ;
        RECT 63.195 173.410 63.435 173.785 ;
        RECT 63.920 173.740 64.090 174.075 ;
        RECT 65.080 173.905 65.255 174.710 ;
        RECT 66.365 174.625 66.625 175.765 ;
        RECT 66.865 175.255 68.480 175.585 ;
        RECT 66.875 174.455 67.045 175.015 ;
        RECT 67.305 174.915 68.480 175.085 ;
        RECT 68.650 174.965 68.930 175.765 ;
        RECT 67.305 174.625 67.635 174.915 ;
        RECT 68.310 174.795 68.480 174.915 ;
        RECT 67.805 174.455 68.050 174.745 ;
        RECT 68.310 174.625 68.970 174.795 ;
        RECT 69.140 174.625 69.415 175.595 ;
        RECT 69.605 174.875 69.865 175.585 ;
        RECT 70.035 175.055 70.365 175.765 ;
        RECT 70.535 174.875 70.765 175.585 ;
        RECT 69.605 174.635 70.765 174.875 ;
        RECT 70.945 174.855 71.215 175.585 ;
        RECT 71.395 175.035 71.735 175.765 ;
        RECT 70.945 174.635 71.715 174.855 ;
        RECT 68.800 174.455 68.970 174.625 ;
        RECT 66.370 174.205 66.705 174.455 ;
        RECT 66.875 174.125 67.590 174.455 ;
        RECT 67.805 174.125 68.630 174.455 ;
        RECT 68.800 174.125 69.075 174.455 ;
        RECT 66.875 174.035 67.125 174.125 ;
        RECT 63.715 173.545 64.090 173.740 ;
        RECT 63.715 173.400 63.885 173.545 ;
        RECT 64.450 173.215 64.845 173.710 ;
        RECT 65.015 173.385 65.255 173.905 ;
        RECT 66.365 173.215 66.625 174.035 ;
        RECT 66.795 173.615 67.125 174.035 ;
        RECT 68.800 173.955 68.970 174.125 ;
        RECT 67.305 173.785 68.970 173.955 ;
        RECT 69.245 173.890 69.415 174.625 ;
        RECT 69.595 174.125 69.895 174.455 ;
        RECT 70.075 174.145 70.600 174.455 ;
        RECT 70.780 174.145 71.245 174.455 ;
        RECT 67.305 173.385 67.565 173.785 ;
        RECT 67.735 173.215 68.065 173.615 ;
        RECT 68.235 173.435 68.405 173.785 ;
        RECT 68.575 173.215 68.950 173.615 ;
        RECT 69.140 173.545 69.415 173.890 ;
        RECT 69.605 173.215 69.895 173.945 ;
        RECT 70.075 173.505 70.305 174.145 ;
        RECT 71.425 173.965 71.715 174.635 ;
        RECT 70.485 173.765 71.715 173.965 ;
        RECT 70.485 173.395 70.795 173.765 ;
        RECT 70.975 173.215 71.645 173.585 ;
        RECT 71.905 173.395 72.165 175.585 ;
        RECT 72.345 174.625 72.605 175.765 ;
        RECT 72.775 174.615 73.105 175.595 ;
        RECT 73.275 174.625 73.555 175.765 ;
        RECT 73.725 174.675 75.395 175.765 ;
        RECT 72.365 174.205 72.700 174.455 ;
        RECT 72.870 174.015 73.040 174.615 ;
        RECT 73.210 174.185 73.545 174.455 ;
        RECT 72.345 173.385 73.040 174.015 ;
        RECT 73.245 173.215 73.555 174.015 ;
        RECT 73.725 173.985 74.475 174.505 ;
        RECT 74.645 174.155 75.395 174.675 ;
        RECT 75.565 174.585 75.885 175.765 ;
        RECT 76.055 174.745 76.255 175.535 ;
        RECT 76.580 174.935 76.965 175.595 ;
        RECT 77.360 175.005 78.145 175.765 ;
        RECT 76.555 174.835 76.965 174.935 ;
        RECT 76.055 174.575 76.385 174.745 ;
        RECT 76.555 174.625 78.165 174.835 ;
        RECT 76.205 174.455 76.385 174.575 ;
        RECT 75.565 174.205 76.030 174.405 ;
        RECT 76.205 174.205 76.535 174.455 ;
        RECT 76.705 174.405 77.170 174.455 ;
        RECT 76.705 174.235 77.175 174.405 ;
        RECT 76.705 174.205 77.170 174.235 ;
        RECT 77.365 174.205 77.720 174.455 ;
        RECT 77.890 174.025 78.165 174.625 ;
        RECT 73.725 173.215 75.395 173.985 ;
        RECT 75.565 173.825 76.745 173.995 ;
        RECT 75.565 173.410 75.905 173.825 ;
        RECT 76.075 173.215 76.245 173.655 ;
        RECT 76.415 173.605 76.745 173.825 ;
        RECT 76.915 173.845 78.165 174.025 ;
        RECT 76.915 173.775 77.280 173.845 ;
        RECT 76.415 173.425 77.665 173.605 ;
        RECT 77.935 173.215 78.105 173.675 ;
        RECT 78.335 173.495 78.615 175.595 ;
        RECT 78.785 175.345 79.125 175.765 ;
        RECT 79.295 175.175 79.545 175.595 ;
        RECT 78.785 175.005 79.545 175.175 ;
        RECT 78.785 174.035 79.095 175.005 ;
        RECT 79.715 174.925 80.045 175.765 ;
        RECT 80.535 175.175 81.290 175.595 ;
        RECT 80.215 175.005 81.680 175.175 ;
        RECT 80.215 174.755 80.385 175.005 ;
        RECT 79.425 174.585 80.385 174.755 ;
        RECT 79.425 174.415 79.595 174.585 ;
        RECT 80.555 174.415 80.860 174.835 ;
        RECT 79.265 174.205 79.595 174.415 ;
        RECT 79.765 174.205 80.205 174.415 ;
        RECT 80.375 174.205 80.860 174.415 ;
        RECT 81.050 174.405 81.340 174.835 ;
        RECT 81.510 174.800 81.680 175.005 ;
        RECT 81.850 174.980 82.090 175.765 ;
        RECT 82.260 174.800 82.590 175.595 ;
        RECT 81.510 174.625 82.590 174.800 ;
        RECT 82.935 174.815 83.210 175.585 ;
        RECT 83.380 175.155 83.710 175.585 ;
        RECT 83.880 175.325 84.075 175.765 ;
        RECT 84.255 175.155 84.585 175.585 ;
        RECT 83.380 174.985 84.585 175.155 ;
        RECT 82.935 174.625 83.520 174.815 ;
        RECT 83.690 174.655 84.585 174.985 ;
        RECT 81.510 174.575 82.295 174.625 ;
        RECT 81.050 174.205 81.440 174.405 ;
        RECT 81.610 174.205 81.955 174.405 ;
        RECT 78.785 173.865 79.545 174.035 ;
        RECT 78.875 173.215 79.045 173.695 ;
        RECT 79.215 173.395 79.545 173.865 ;
        RECT 79.715 173.215 79.885 174.035 ;
        RECT 80.055 173.865 81.755 174.035 ;
        RECT 80.055 173.400 80.385 173.865 ;
        RECT 81.370 173.775 81.755 173.865 ;
        RECT 82.125 173.935 82.295 174.575 ;
        RECT 82.495 174.105 82.755 174.455 ;
        RECT 82.125 173.765 82.670 173.935 ;
        RECT 82.935 173.805 83.175 174.455 ;
        RECT 83.345 173.955 83.520 174.625 ;
        RECT 83.690 174.125 84.105 174.455 ;
        RECT 84.285 174.125 84.580 174.455 ;
        RECT 83.345 173.775 83.675 173.955 ;
        RECT 80.555 173.215 80.725 173.685 ;
        RECT 80.985 173.425 82.170 173.595 ;
        RECT 82.340 173.385 82.670 173.765 ;
        RECT 82.950 173.215 83.280 173.605 ;
        RECT 83.450 173.395 83.675 173.775 ;
        RECT 83.875 173.505 84.105 174.125 ;
        RECT 84.285 173.215 84.585 173.945 ;
        RECT 85.685 173.385 86.435 175.595 ;
        RECT 86.695 174.835 86.865 175.595 ;
        RECT 87.045 175.005 87.375 175.765 ;
        RECT 86.695 174.665 87.360 174.835 ;
        RECT 87.545 174.690 87.815 175.595 ;
        RECT 87.190 174.520 87.360 174.665 ;
        RECT 86.625 174.115 86.955 174.485 ;
        RECT 87.190 174.190 87.475 174.520 ;
        RECT 87.190 173.935 87.360 174.190 ;
        RECT 86.695 173.765 87.360 173.935 ;
        RECT 87.645 173.890 87.815 174.690 ;
        RECT 87.985 174.600 88.275 175.765 ;
        RECT 89.375 174.625 89.705 175.765 ;
        RECT 90.235 174.795 90.565 175.580 ;
        RECT 89.885 174.625 90.565 174.795 ;
        RECT 90.745 174.915 91.005 175.595 ;
        RECT 91.175 174.985 91.425 175.765 ;
        RECT 91.675 175.215 91.925 175.595 ;
        RECT 92.095 175.385 92.450 175.765 ;
        RECT 93.455 175.375 93.790 175.595 ;
        RECT 93.055 175.215 93.285 175.255 ;
        RECT 91.675 175.015 93.285 175.215 ;
        RECT 91.675 175.005 92.510 175.015 ;
        RECT 93.100 174.925 93.285 175.015 ;
        RECT 89.365 174.205 89.715 174.455 ;
        RECT 89.885 174.025 90.055 174.625 ;
        RECT 90.225 174.205 90.575 174.455 ;
        RECT 86.695 173.385 86.865 173.765 ;
        RECT 87.045 173.215 87.375 173.595 ;
        RECT 87.555 173.385 87.815 173.890 ;
        RECT 87.985 173.215 88.275 173.940 ;
        RECT 89.375 173.215 89.645 174.025 ;
        RECT 89.815 173.385 90.145 174.025 ;
        RECT 90.315 173.215 90.555 174.025 ;
        RECT 90.745 173.725 90.915 174.915 ;
        RECT 92.615 174.815 92.945 174.845 ;
        RECT 91.145 174.755 92.945 174.815 ;
        RECT 93.535 174.755 93.790 175.375 ;
        RECT 94.055 175.020 94.325 175.765 ;
        RECT 94.955 175.760 101.230 175.765 ;
        RECT 94.495 174.850 94.785 175.590 ;
        RECT 94.955 175.035 95.210 175.760 ;
        RECT 95.395 174.865 95.655 175.590 ;
        RECT 95.825 175.035 96.070 175.760 ;
        RECT 96.255 174.865 96.515 175.590 ;
        RECT 96.685 175.035 96.930 175.760 ;
        RECT 97.115 174.865 97.375 175.590 ;
        RECT 97.545 175.035 97.790 175.760 ;
        RECT 97.960 174.865 98.220 175.590 ;
        RECT 98.390 175.035 98.650 175.760 ;
        RECT 98.820 174.865 99.080 175.590 ;
        RECT 99.250 175.035 99.510 175.760 ;
        RECT 99.680 174.865 99.940 175.590 ;
        RECT 100.110 175.035 100.370 175.760 ;
        RECT 100.540 174.865 100.800 175.590 ;
        RECT 100.970 174.965 101.230 175.760 ;
        RECT 95.395 174.850 100.800 174.865 ;
        RECT 91.085 174.645 93.790 174.755 ;
        RECT 91.085 174.610 91.285 174.645 ;
        RECT 91.085 174.035 91.255 174.610 ;
        RECT 92.615 174.585 93.790 174.645 ;
        RECT 94.055 174.625 100.800 174.850 ;
        RECT 91.485 174.170 91.895 174.475 ;
        RECT 92.065 174.205 92.395 174.415 ;
        RECT 91.085 173.915 91.355 174.035 ;
        RECT 91.085 173.870 91.930 173.915 ;
        RECT 91.175 173.745 91.930 173.870 ;
        RECT 92.185 173.805 92.395 174.205 ;
        RECT 92.640 174.205 93.115 174.415 ;
        RECT 93.305 174.205 93.795 174.405 ;
        RECT 92.640 173.805 92.860 174.205 ;
        RECT 94.055 174.035 95.220 174.625 ;
        RECT 101.400 174.455 101.650 175.590 ;
        RECT 101.830 174.955 102.090 175.765 ;
        RECT 102.265 174.455 102.510 175.595 ;
        RECT 102.690 174.955 102.985 175.765 ;
        RECT 103.175 174.625 103.505 175.765 ;
        RECT 104.035 174.795 104.365 175.580 ;
        RECT 103.685 174.625 104.365 174.795 ;
        RECT 104.545 174.675 108.055 175.765 ;
        RECT 95.390 174.205 102.510 174.455 ;
        RECT 90.745 173.715 90.975 173.725 ;
        RECT 90.745 173.385 91.005 173.715 ;
        RECT 91.760 173.595 91.930 173.745 ;
        RECT 91.175 173.215 91.505 173.575 ;
        RECT 91.760 173.385 93.060 173.595 ;
        RECT 93.335 173.215 93.790 173.980 ;
        RECT 94.055 173.865 100.800 174.035 ;
        RECT 94.055 173.215 94.355 173.695 ;
        RECT 94.525 173.410 94.785 173.865 ;
        RECT 94.955 173.215 95.215 173.695 ;
        RECT 95.395 173.410 95.655 173.865 ;
        RECT 95.825 173.215 96.075 173.695 ;
        RECT 96.255 173.410 96.515 173.865 ;
        RECT 96.685 173.215 96.935 173.695 ;
        RECT 97.115 173.410 97.375 173.865 ;
        RECT 97.545 173.215 97.790 173.695 ;
        RECT 97.960 173.410 98.235 173.865 ;
        RECT 98.405 173.215 98.650 173.695 ;
        RECT 98.820 173.410 99.080 173.865 ;
        RECT 99.250 173.215 99.510 173.695 ;
        RECT 99.680 173.410 99.940 173.865 ;
        RECT 100.110 173.215 100.370 173.695 ;
        RECT 100.540 173.410 100.800 173.865 ;
        RECT 100.970 173.215 101.230 173.775 ;
        RECT 101.400 173.395 101.650 174.205 ;
        RECT 101.830 173.215 102.090 173.740 ;
        RECT 102.260 173.395 102.510 174.205 ;
        RECT 102.680 173.895 102.995 174.455 ;
        RECT 103.165 174.205 103.515 174.455 ;
        RECT 103.685 174.025 103.855 174.625 ;
        RECT 104.025 174.205 104.375 174.455 ;
        RECT 102.690 173.215 102.995 173.725 ;
        RECT 103.175 173.215 103.445 174.025 ;
        RECT 103.615 173.385 103.945 174.025 ;
        RECT 104.115 173.215 104.355 174.025 ;
        RECT 104.545 173.985 106.195 174.505 ;
        RECT 106.365 174.155 108.055 174.675 ;
        RECT 108.225 174.625 108.585 175.765 ;
        RECT 109.255 175.085 109.585 175.595 ;
        RECT 110.755 175.255 111.265 175.765 ;
        RECT 108.755 174.915 111.265 175.085 ;
        RECT 108.225 174.375 108.555 174.455 ;
        RECT 108.225 174.205 108.585 174.375 ;
        RECT 104.545 173.215 108.055 173.985 ;
        RECT 108.225 173.555 108.585 174.035 ;
        RECT 108.755 173.955 108.955 174.915 ;
        RECT 109.125 174.575 109.375 174.745 ;
        RECT 109.125 174.125 109.370 174.575 ;
        RECT 109.645 174.125 109.865 174.745 ;
        RECT 110.120 174.125 110.295 174.745 ;
        RECT 110.565 174.125 110.785 174.745 ;
        RECT 110.955 174.125 111.265 174.915 ;
        RECT 108.755 173.725 109.085 173.955 ;
        RECT 109.255 173.785 110.585 173.955 ;
        RECT 109.255 173.555 109.585 173.785 ;
        RECT 108.225 173.385 109.585 173.555 ;
        RECT 109.755 173.215 110.085 173.615 ;
        RECT 110.255 173.385 110.585 173.785 ;
        RECT 110.855 173.215 111.185 173.955 ;
        RECT 111.435 173.385 111.765 175.595 ;
        RECT 111.935 174.625 112.195 175.765 ;
        RECT 112.365 174.625 112.645 175.765 ;
        RECT 112.815 174.615 113.145 175.595 ;
        RECT 113.315 174.625 113.575 175.765 ;
        RECT 112.375 174.185 112.710 174.455 ;
        RECT 112.880 174.015 113.050 174.615 ;
        RECT 113.745 174.600 114.035 175.765 ;
        RECT 114.215 174.955 114.510 175.765 ;
        RECT 114.690 174.455 114.935 175.595 ;
        RECT 115.110 174.955 115.370 175.765 ;
        RECT 115.970 175.760 122.245 175.765 ;
        RECT 115.550 174.455 115.800 175.590 ;
        RECT 115.970 174.965 116.230 175.760 ;
        RECT 116.400 174.865 116.660 175.590 ;
        RECT 116.830 175.035 117.090 175.760 ;
        RECT 117.260 174.865 117.520 175.590 ;
        RECT 117.690 175.035 117.950 175.760 ;
        RECT 118.120 174.865 118.380 175.590 ;
        RECT 118.550 175.035 118.810 175.760 ;
        RECT 118.980 174.865 119.240 175.590 ;
        RECT 119.410 175.035 119.655 175.760 ;
        RECT 119.825 174.865 120.085 175.590 ;
        RECT 120.270 175.035 120.515 175.760 ;
        RECT 120.685 174.865 120.945 175.590 ;
        RECT 121.130 175.035 121.375 175.760 ;
        RECT 121.545 174.865 121.805 175.590 ;
        RECT 121.990 175.035 122.245 175.760 ;
        RECT 116.400 174.850 121.805 174.865 ;
        RECT 122.415 174.850 122.705 175.590 ;
        RECT 122.875 175.020 123.145 175.765 ;
        RECT 123.415 174.955 123.710 175.765 ;
        RECT 116.400 174.625 123.145 174.850 ;
        RECT 113.220 174.205 113.555 174.455 ;
        RECT 111.935 173.215 112.195 174.015 ;
        RECT 112.365 173.215 112.675 174.015 ;
        RECT 112.880 173.385 113.575 174.015 ;
        RECT 113.745 173.215 114.035 173.940 ;
        RECT 114.205 173.895 114.520 174.455 ;
        RECT 114.690 174.205 121.810 174.455 ;
        RECT 114.205 173.215 114.510 173.725 ;
        RECT 114.690 173.395 114.940 174.205 ;
        RECT 115.110 173.215 115.370 173.740 ;
        RECT 115.550 173.395 115.800 174.205 ;
        RECT 121.980 174.035 123.145 174.625 ;
        RECT 123.890 174.455 124.135 175.595 ;
        RECT 124.310 174.955 124.570 175.765 ;
        RECT 125.170 175.760 131.445 175.765 ;
        RECT 124.750 174.455 125.000 175.590 ;
        RECT 125.170 174.965 125.430 175.760 ;
        RECT 125.600 174.865 125.860 175.590 ;
        RECT 126.030 175.035 126.290 175.760 ;
        RECT 126.460 174.865 126.720 175.590 ;
        RECT 126.890 175.035 127.150 175.760 ;
        RECT 127.320 174.865 127.580 175.590 ;
        RECT 127.750 175.035 128.010 175.760 ;
        RECT 128.180 174.865 128.440 175.590 ;
        RECT 128.610 175.035 128.855 175.760 ;
        RECT 129.025 174.865 129.285 175.590 ;
        RECT 129.470 175.035 129.715 175.760 ;
        RECT 129.885 174.865 130.145 175.590 ;
        RECT 130.330 175.035 130.575 175.760 ;
        RECT 130.745 174.865 131.005 175.590 ;
        RECT 131.190 175.035 131.445 175.760 ;
        RECT 125.600 174.850 131.005 174.865 ;
        RECT 131.615 174.850 131.905 175.590 ;
        RECT 132.075 175.020 132.345 175.765 ;
        RECT 125.600 174.625 132.345 174.850 ;
        RECT 133.155 174.835 133.325 175.595 ;
        RECT 133.540 175.005 133.870 175.765 ;
        RECT 133.155 174.665 133.870 174.835 ;
        RECT 134.040 174.690 134.295 175.595 ;
        RECT 116.400 173.865 123.145 174.035 ;
        RECT 123.405 173.895 123.720 174.455 ;
        RECT 123.890 174.205 131.010 174.455 ;
        RECT 115.970 173.215 116.230 173.775 ;
        RECT 116.400 173.410 116.660 173.865 ;
        RECT 116.830 173.215 117.090 173.695 ;
        RECT 117.260 173.410 117.520 173.865 ;
        RECT 117.690 173.215 117.950 173.695 ;
        RECT 118.120 173.410 118.380 173.865 ;
        RECT 118.550 173.215 118.795 173.695 ;
        RECT 118.965 173.410 119.240 173.865 ;
        RECT 119.410 173.215 119.655 173.695 ;
        RECT 119.825 173.410 120.085 173.865 ;
        RECT 120.265 173.215 120.515 173.695 ;
        RECT 120.685 173.410 120.945 173.865 ;
        RECT 121.125 173.215 121.375 173.695 ;
        RECT 121.545 173.410 121.805 173.865 ;
        RECT 121.985 173.215 122.245 173.695 ;
        RECT 122.415 173.410 122.675 173.865 ;
        RECT 122.845 173.215 123.145 173.695 ;
        RECT 123.405 173.215 123.710 173.725 ;
        RECT 123.890 173.395 124.140 174.205 ;
        RECT 124.310 173.215 124.570 173.740 ;
        RECT 124.750 173.395 125.000 174.205 ;
        RECT 131.180 174.035 132.345 174.625 ;
        RECT 133.065 174.115 133.420 174.485 ;
        RECT 133.700 174.455 133.870 174.665 ;
        RECT 133.700 174.125 133.955 174.455 ;
        RECT 125.600 173.865 132.345 174.035 ;
        RECT 133.700 173.935 133.870 174.125 ;
        RECT 134.125 173.960 134.295 174.690 ;
        RECT 134.470 174.615 134.730 175.765 ;
        RECT 134.905 174.675 136.115 175.765 ;
        RECT 134.905 174.135 135.425 174.675 ;
        RECT 125.170 173.215 125.430 173.775 ;
        RECT 125.600 173.410 125.860 173.865 ;
        RECT 126.030 173.215 126.290 173.695 ;
        RECT 126.460 173.410 126.720 173.865 ;
        RECT 126.890 173.215 127.150 173.695 ;
        RECT 127.320 173.410 127.580 173.865 ;
        RECT 127.750 173.215 127.995 173.695 ;
        RECT 128.165 173.410 128.440 173.865 ;
        RECT 128.610 173.215 128.855 173.695 ;
        RECT 129.025 173.410 129.285 173.865 ;
        RECT 129.465 173.215 129.715 173.695 ;
        RECT 129.885 173.410 130.145 173.865 ;
        RECT 130.325 173.215 130.575 173.695 ;
        RECT 130.745 173.410 131.005 173.865 ;
        RECT 131.185 173.215 131.445 173.695 ;
        RECT 131.615 173.410 131.875 173.865 ;
        RECT 133.155 173.765 133.870 173.935 ;
        RECT 132.045 173.215 132.345 173.695 ;
        RECT 133.155 173.385 133.325 173.765 ;
        RECT 133.540 173.215 133.870 173.595 ;
        RECT 134.040 173.385 134.295 173.960 ;
        RECT 134.470 173.215 134.730 174.055 ;
        RECT 135.595 173.965 136.115 174.505 ;
        RECT 134.905 173.215 136.115 173.965 ;
        RECT 23.500 173.045 136.200 173.215 ;
        RECT 23.585 172.295 24.795 173.045 ;
        RECT 24.965 172.545 25.225 172.875 ;
        RECT 25.435 172.565 25.710 173.045 ;
        RECT 23.585 171.755 24.105 172.295 ;
        RECT 24.275 171.585 24.795 172.125 ;
        RECT 23.585 170.495 24.795 171.585 ;
        RECT 24.965 171.635 25.135 172.545 ;
        RECT 25.920 172.475 26.125 172.875 ;
        RECT 26.295 172.645 26.630 173.045 ;
        RECT 25.305 171.805 25.665 172.385 ;
        RECT 25.920 172.305 26.605 172.475 ;
        RECT 25.845 171.635 26.095 172.135 ;
        RECT 24.965 171.465 26.095 171.635 ;
        RECT 24.965 170.695 25.235 171.465 ;
        RECT 26.265 171.275 26.605 172.305 ;
        RECT 25.405 170.495 25.735 171.275 ;
        RECT 25.940 171.100 26.605 171.275 ;
        RECT 27.725 172.370 27.985 172.875 ;
        RECT 28.165 172.665 28.495 173.045 ;
        RECT 28.675 172.495 28.845 172.875 ;
        RECT 29.105 172.500 34.450 173.045 ;
        RECT 27.725 171.570 27.895 172.370 ;
        RECT 28.180 172.325 28.845 172.495 ;
        RECT 28.180 172.070 28.350 172.325 ;
        RECT 28.065 171.740 28.350 172.070 ;
        RECT 28.585 171.775 28.915 172.145 ;
        RECT 28.180 171.595 28.350 171.740 ;
        RECT 30.690 171.670 31.030 172.500 ;
        RECT 35.175 172.495 35.345 172.875 ;
        RECT 35.515 172.665 35.845 173.045 ;
        RECT 35.175 172.325 35.670 172.495 ;
        RECT 25.940 170.695 26.125 171.100 ;
        RECT 26.295 170.495 26.630 170.920 ;
        RECT 27.725 170.665 27.995 171.570 ;
        RECT 28.180 171.425 28.845 171.595 ;
        RECT 28.165 170.495 28.495 171.255 ;
        RECT 28.675 170.665 28.845 171.425 ;
        RECT 32.510 170.930 32.860 172.180 ;
        RECT 35.150 172.025 35.330 172.135 ;
        RECT 35.145 171.855 35.330 172.025 ;
        RECT 35.150 171.495 35.330 171.855 ;
        RECT 35.500 171.245 35.670 172.325 ;
        RECT 36.015 171.585 36.240 172.875 ;
        RECT 36.410 172.665 36.740 173.045 ;
        RECT 37.010 172.495 37.180 172.875 ;
        RECT 36.415 172.325 37.405 172.495 ;
        RECT 36.415 171.805 36.585 172.325 ;
        RECT 36.755 171.805 37.065 172.135 ;
        RECT 35.990 171.415 36.320 171.585 ;
        RECT 36.755 171.245 36.925 171.805 ;
        RECT 35.175 171.075 36.925 171.245 ;
        RECT 37.235 171.215 37.405 172.325 ;
        RECT 37.910 172.025 38.175 172.710 ;
        RECT 37.905 171.855 38.175 172.025 ;
        RECT 37.575 171.555 37.745 171.730 ;
        RECT 38.350 171.725 38.655 172.705 ;
        RECT 38.835 172.545 39.085 173.045 ;
        RECT 39.255 172.545 39.515 172.875 ;
        RECT 38.825 171.825 39.175 172.365 ;
        RECT 37.575 171.385 38.755 171.555 ;
        RECT 38.585 171.215 38.755 171.385 ;
        RECT 39.345 171.215 39.515 172.545 ;
        RECT 29.105 170.495 34.450 170.930 ;
        RECT 35.175 170.665 35.345 171.075 ;
        RECT 37.235 171.045 38.415 171.215 ;
        RECT 38.585 171.045 39.515 171.215 ;
        RECT 35.515 170.495 35.845 170.875 ;
        RECT 36.490 170.495 37.160 170.875 ;
        RECT 37.395 170.665 37.565 171.045 ;
        RECT 37.735 170.495 38.075 170.875 ;
        RECT 38.245 170.665 38.415 171.045 ;
        RECT 38.755 170.495 39.085 170.875 ;
        RECT 39.255 170.665 39.515 171.045 ;
        RECT 39.685 172.395 39.945 172.875 ;
        RECT 40.115 172.585 40.445 173.045 ;
        RECT 40.635 172.405 40.835 172.825 ;
        RECT 39.685 171.365 39.855 172.395 ;
        RECT 40.025 171.705 40.255 172.135 ;
        RECT 40.425 171.885 40.835 172.405 ;
        RECT 41.005 172.560 41.795 172.825 ;
        RECT 41.005 171.705 41.260 172.560 ;
        RECT 41.975 172.225 42.305 172.645 ;
        RECT 42.475 172.225 42.735 173.045 ;
        RECT 43.105 172.415 43.435 172.775 ;
        RECT 44.055 172.585 44.305 173.045 ;
        RECT 44.475 172.585 45.035 172.875 ;
        RECT 43.105 172.225 44.495 172.415 ;
        RECT 41.975 172.135 42.225 172.225 ;
        RECT 41.430 171.885 42.225 172.135 ;
        RECT 44.325 172.135 44.495 172.225 ;
        RECT 40.025 171.535 41.815 171.705 ;
        RECT 39.685 170.665 39.960 171.365 ;
        RECT 40.130 171.240 40.845 171.535 ;
        RECT 41.065 171.175 41.395 171.365 ;
        RECT 40.170 170.495 40.385 171.040 ;
        RECT 40.555 170.665 41.030 171.005 ;
        RECT 41.200 171.000 41.395 171.175 ;
        RECT 41.565 171.170 41.815 171.535 ;
        RECT 41.200 170.495 41.815 171.000 ;
        RECT 42.055 170.665 42.225 171.885 ;
        RECT 42.395 171.175 42.735 172.055 ;
        RECT 42.920 171.805 43.595 172.055 ;
        RECT 43.815 171.805 44.155 172.055 ;
        RECT 44.325 171.805 44.615 172.135 ;
        RECT 42.920 171.445 43.185 171.805 ;
        RECT 44.325 171.555 44.495 171.805 ;
        RECT 43.555 171.385 44.495 171.555 ;
        RECT 42.475 170.495 42.735 171.005 ;
        RECT 43.105 170.495 43.385 171.165 ;
        RECT 43.555 170.835 43.855 171.385 ;
        RECT 44.785 171.215 45.035 172.585 ;
        RECT 45.205 172.275 48.715 173.045 ;
        RECT 49.345 172.320 49.635 173.045 ;
        RECT 49.805 172.500 55.150 173.045 ;
        RECT 55.325 172.500 60.670 173.045 ;
        RECT 45.205 171.755 46.855 172.275 ;
        RECT 47.025 171.585 48.715 172.105 ;
        RECT 51.390 171.670 51.730 172.500 ;
        RECT 44.055 170.495 44.385 171.215 ;
        RECT 44.575 170.665 45.035 171.215 ;
        RECT 45.205 170.495 48.715 171.585 ;
        RECT 49.345 170.495 49.635 171.660 ;
        RECT 53.210 170.930 53.560 172.180 ;
        RECT 56.910 171.670 57.250 172.500 ;
        RECT 60.845 172.275 63.435 173.045 ;
        RECT 63.605 172.405 63.945 172.810 ;
        RECT 64.115 172.575 64.285 173.045 ;
        RECT 64.455 172.405 64.705 172.810 ;
        RECT 58.730 170.930 59.080 172.180 ;
        RECT 60.845 171.755 62.055 172.275 ;
        RECT 63.605 172.225 64.705 172.405 ;
        RECT 64.875 172.440 65.125 172.810 ;
        RECT 65.295 172.565 65.740 172.735 ;
        RECT 65.910 172.705 66.130 172.750 ;
        RECT 62.225 171.585 63.435 172.105 ;
        RECT 64.875 172.055 65.045 172.440 ;
        RECT 49.805 170.495 55.150 170.930 ;
        RECT 55.325 170.495 60.670 170.930 ;
        RECT 60.845 170.495 63.435 171.585 ;
        RECT 63.605 171.485 63.950 172.055 ;
        RECT 64.120 171.805 64.680 172.055 ;
        RECT 64.850 171.885 65.045 172.055 ;
        RECT 63.605 170.495 63.950 171.315 ;
        RECT 64.120 170.705 64.295 171.805 ;
        RECT 64.850 171.635 65.020 171.885 ;
        RECT 65.295 171.775 65.465 172.565 ;
        RECT 65.910 172.535 66.135 172.705 ;
        RECT 65.910 172.395 66.130 172.535 ;
        RECT 65.635 172.225 66.130 172.395 ;
        RECT 66.410 172.380 66.580 173.045 ;
        RECT 66.775 172.305 67.115 172.875 ;
        RECT 65.635 172.030 65.810 172.225 ;
        RECT 65.980 171.855 66.430 172.055 ;
        RECT 64.465 171.245 65.020 171.635 ;
        RECT 65.190 171.635 65.465 171.775 ;
        RECT 66.600 171.685 66.770 172.135 ;
        RECT 65.190 171.415 66.205 171.635 ;
        RECT 66.375 171.515 66.770 171.685 ;
        RECT 66.375 171.245 66.545 171.515 ;
        RECT 66.940 171.335 67.115 172.305 ;
        RECT 67.745 172.225 68.005 173.045 ;
        RECT 68.175 172.225 68.505 172.645 ;
        RECT 68.685 172.475 68.945 172.875 ;
        RECT 69.115 172.645 69.445 173.045 ;
        RECT 69.615 172.475 69.785 172.825 ;
        RECT 69.955 172.645 70.330 173.045 ;
        RECT 68.685 172.305 70.350 172.475 ;
        RECT 70.520 172.370 70.795 172.715 ;
        RECT 68.255 172.135 68.505 172.225 ;
        RECT 70.180 172.135 70.350 172.305 ;
        RECT 67.750 171.805 68.085 172.055 ;
        RECT 68.255 171.805 68.970 172.135 ;
        RECT 69.185 171.805 70.010 172.135 ;
        RECT 70.180 171.805 70.455 172.135 ;
        RECT 64.465 171.075 66.545 171.245 ;
        RECT 64.465 170.840 64.795 171.075 ;
        RECT 65.085 170.495 65.485 170.895 ;
        RECT 66.355 170.495 66.685 170.895 ;
        RECT 66.855 170.665 67.115 171.335 ;
        RECT 67.745 170.495 68.005 171.635 ;
        RECT 68.255 171.245 68.425 171.805 ;
        RECT 68.685 171.345 69.015 171.635 ;
        RECT 69.185 171.515 69.430 171.805 ;
        RECT 70.180 171.635 70.350 171.805 ;
        RECT 70.625 171.635 70.795 172.370 ;
        RECT 69.690 171.465 70.350 171.635 ;
        RECT 69.690 171.345 69.860 171.465 ;
        RECT 68.685 171.175 69.860 171.345 ;
        RECT 68.245 170.675 69.860 171.005 ;
        RECT 70.030 170.495 70.310 171.295 ;
        RECT 70.520 170.665 70.795 171.635 ;
        RECT 70.975 172.320 71.305 172.830 ;
        RECT 71.475 172.645 71.805 173.045 ;
        RECT 72.855 172.475 73.185 172.815 ;
        RECT 73.355 172.645 73.685 173.045 ;
        RECT 70.975 171.555 71.165 172.320 ;
        RECT 71.475 172.305 73.840 172.475 ;
        RECT 75.105 172.320 75.395 173.045 ;
        RECT 76.495 172.315 76.795 173.045 ;
        RECT 71.475 172.135 71.645 172.305 ;
        RECT 71.335 171.805 71.645 172.135 ;
        RECT 71.815 171.805 72.120 172.135 ;
        RECT 70.975 170.705 71.305 171.555 ;
        RECT 71.475 170.495 71.725 171.635 ;
        RECT 71.905 171.475 72.120 171.805 ;
        RECT 72.295 171.475 72.580 172.135 ;
        RECT 72.775 171.475 73.040 172.135 ;
        RECT 73.255 171.475 73.500 172.135 ;
        RECT 73.670 171.305 73.840 172.305 ;
        RECT 76.975 172.135 77.205 172.755 ;
        RECT 77.405 172.485 77.630 172.865 ;
        RECT 77.800 172.655 78.130 173.045 ;
        RECT 78.335 172.705 78.670 172.875 ;
        RECT 77.405 172.305 77.735 172.485 ;
        RECT 76.500 171.805 76.795 172.135 ;
        RECT 76.975 171.805 77.390 172.135 ;
        RECT 71.915 171.135 73.205 171.305 ;
        RECT 71.915 170.715 72.165 171.135 ;
        RECT 72.395 170.495 72.725 170.965 ;
        RECT 72.955 170.715 73.205 171.135 ;
        RECT 73.385 171.135 73.840 171.305 ;
        RECT 73.385 170.705 73.715 171.135 ;
        RECT 75.105 170.495 75.395 171.660 ;
        RECT 77.560 171.635 77.735 172.305 ;
        RECT 77.905 171.805 78.145 172.455 ;
        RECT 78.335 172.305 78.950 172.705 ;
        RECT 79.630 172.665 79.965 173.045 ;
        RECT 80.555 172.605 80.790 173.045 ;
        RECT 80.960 172.515 81.290 172.875 ;
        RECT 81.460 172.685 81.790 173.045 ;
        RECT 79.120 172.305 80.390 172.495 ;
        RECT 80.960 172.345 81.780 172.515 ;
        RECT 78.325 171.805 78.600 172.135 ;
        RECT 76.495 171.275 77.390 171.605 ;
        RECT 77.560 171.445 78.145 171.635 ;
        RECT 78.770 171.620 78.950 172.305 ;
        RECT 79.120 171.805 79.480 172.135 ;
        RECT 79.770 172.025 80.060 172.135 ;
        RECT 79.765 171.855 80.060 172.025 ;
        RECT 79.770 171.805 80.060 171.855 ;
        RECT 80.230 171.805 80.565 172.135 ;
        RECT 80.735 171.805 81.415 172.135 ;
        RECT 80.735 171.620 80.905 171.805 ;
        RECT 76.495 171.105 77.700 171.275 ;
        RECT 76.495 170.675 76.825 171.105 ;
        RECT 77.005 170.495 77.200 170.935 ;
        RECT 77.370 170.675 77.700 171.105 ;
        RECT 77.870 170.675 78.145 171.445 ;
        RECT 78.330 171.365 80.905 171.620 ;
        RECT 78.330 170.665 78.595 171.365 ;
        RECT 78.765 170.495 79.095 171.195 ;
        RECT 79.265 170.665 79.935 171.365 ;
        RECT 81.585 171.225 81.780 172.345 ;
        RECT 82.945 171.465 83.175 172.805 ;
        RECT 83.355 171.965 83.585 172.865 ;
        RECT 83.785 172.265 84.030 173.045 ;
        RECT 84.200 172.505 84.630 172.865 ;
        RECT 85.210 172.675 85.940 173.045 ;
        RECT 84.200 172.315 85.940 172.505 ;
        RECT 84.200 172.085 84.420 172.315 ;
        RECT 83.355 171.285 83.695 171.965 ;
        RECT 80.440 170.495 80.870 171.195 ;
        RECT 81.050 171.055 81.780 171.225 ;
        RECT 82.945 171.085 83.695 171.285 ;
        RECT 83.875 171.785 84.420 172.085 ;
        RECT 81.050 170.665 81.240 171.055 ;
        RECT 81.410 170.495 81.740 170.875 ;
        RECT 82.945 170.695 83.185 171.085 ;
        RECT 83.355 170.495 83.705 170.905 ;
        RECT 83.875 170.675 84.205 171.785 ;
        RECT 84.590 171.515 85.015 172.135 ;
        RECT 85.210 171.515 85.470 172.135 ;
        RECT 85.680 171.805 85.940 172.315 ;
        RECT 84.375 171.145 85.400 171.345 ;
        RECT 84.375 170.675 84.555 171.145 ;
        RECT 84.725 170.495 85.055 170.975 ;
        RECT 85.230 170.675 85.400 171.145 ;
        RECT 85.665 170.495 85.950 171.635 ;
        RECT 86.140 170.675 86.420 172.865 ;
        RECT 86.625 171.465 86.855 172.805 ;
        RECT 87.035 171.965 87.265 172.865 ;
        RECT 87.465 172.265 87.710 173.045 ;
        RECT 87.880 172.505 88.310 172.865 ;
        RECT 88.890 172.675 89.620 173.045 ;
        RECT 87.880 172.315 89.620 172.505 ;
        RECT 87.880 172.085 88.100 172.315 ;
        RECT 87.035 171.285 87.375 171.965 ;
        RECT 86.625 171.085 87.375 171.285 ;
        RECT 87.555 171.785 88.100 172.085 ;
        RECT 86.625 170.695 86.865 171.085 ;
        RECT 87.035 170.495 87.385 170.905 ;
        RECT 87.555 170.675 87.885 171.785 ;
        RECT 88.270 171.515 88.695 172.135 ;
        RECT 88.890 171.515 89.150 172.135 ;
        RECT 89.360 171.805 89.620 172.315 ;
        RECT 88.055 171.145 89.080 171.345 ;
        RECT 88.055 170.675 88.235 171.145 ;
        RECT 88.405 170.495 88.735 170.975 ;
        RECT 88.910 170.675 89.080 171.145 ;
        RECT 89.345 170.495 89.630 171.635 ;
        RECT 89.820 170.675 90.100 172.865 ;
        RECT 90.745 172.245 91.440 172.875 ;
        RECT 91.645 172.245 91.955 173.045 ;
        RECT 92.165 172.645 92.495 173.045 ;
        RECT 92.675 172.625 93.980 172.875 ;
        RECT 92.675 172.475 92.855 172.625 ;
        RECT 94.255 172.535 94.705 173.045 ;
        RECT 92.125 172.305 92.855 172.475 ;
        RECT 95.505 172.485 95.835 172.875 ;
        RECT 96.005 172.655 97.190 172.825 ;
        RECT 97.450 172.575 97.620 173.045 ;
        RECT 90.765 171.805 91.100 172.055 ;
        RECT 91.270 171.645 91.440 172.245 ;
        RECT 91.610 171.805 91.945 172.075 ;
        RECT 90.745 170.495 91.005 171.635 ;
        RECT 91.175 170.665 91.505 171.645 ;
        RECT 92.125 171.635 92.295 172.305 ;
        RECT 92.465 171.805 92.790 172.135 ;
        RECT 93.100 172.055 93.310 172.455 ;
        RECT 92.960 171.855 93.310 172.055 ;
        RECT 93.560 172.055 93.810 172.455 ;
        RECT 93.560 171.855 94.035 172.055 ;
        RECT 94.225 171.855 94.675 172.365 ;
        RECT 95.505 172.305 96.015 172.485 ;
        RECT 95.345 171.845 95.675 172.135 ;
        RECT 92.960 171.635 94.705 171.685 ;
        RECT 95.845 171.675 96.015 172.305 ;
        RECT 96.420 172.395 96.805 172.485 ;
        RECT 97.790 172.395 98.120 172.860 ;
        RECT 96.420 172.225 98.120 172.395 ;
        RECT 98.290 172.225 98.460 173.045 ;
        RECT 98.630 172.225 99.315 172.865 ;
        RECT 99.495 172.235 99.765 173.045 ;
        RECT 99.935 172.235 100.265 172.875 ;
        RECT 100.435 172.235 100.675 173.045 ;
        RECT 100.865 172.320 101.155 173.045 ;
        RECT 96.185 171.845 96.515 172.055 ;
        RECT 96.695 171.805 97.075 172.055 ;
        RECT 91.675 170.495 91.955 171.635 ;
        RECT 92.125 171.505 94.705 171.635 ;
        RECT 92.125 171.465 93.185 171.505 ;
        RECT 93.325 171.295 94.205 171.335 ;
        RECT 92.175 170.495 92.440 171.275 ;
        RECT 92.675 171.095 94.205 171.295 ;
        RECT 92.675 170.965 92.845 171.095 ;
        RECT 93.590 171.045 94.205 171.095 ;
        RECT 93.975 171.005 94.205 171.045 ;
        RECT 92.990 170.495 93.365 170.875 ;
        RECT 93.535 170.835 93.865 170.875 ;
        RECT 94.375 170.835 94.705 171.505 ;
        RECT 93.535 170.665 94.705 170.835 ;
        RECT 95.500 171.505 96.585 171.675 ;
        RECT 95.500 170.665 95.800 171.505 ;
        RECT 95.995 170.495 96.245 171.335 ;
        RECT 96.415 171.255 96.585 171.505 ;
        RECT 96.755 171.425 97.075 171.805 ;
        RECT 97.265 171.845 97.750 172.055 ;
        RECT 97.940 171.845 98.390 172.055 ;
        RECT 98.560 171.845 98.895 172.055 ;
        RECT 97.265 171.685 97.640 171.845 ;
        RECT 97.245 171.515 97.640 171.685 ;
        RECT 98.560 171.675 98.730 171.845 ;
        RECT 97.265 171.425 97.640 171.515 ;
        RECT 97.810 171.505 98.730 171.675 ;
        RECT 97.810 171.255 97.980 171.505 ;
        RECT 96.415 171.085 97.980 171.255 ;
        RECT 96.835 170.665 97.640 171.085 ;
        RECT 98.150 170.495 98.480 171.335 ;
        RECT 99.065 171.255 99.315 172.225 ;
        RECT 99.485 171.805 99.835 172.055 ;
        RECT 100.005 171.635 100.175 172.235 ;
        RECT 101.385 172.225 101.595 173.045 ;
        RECT 101.765 172.245 102.095 172.875 ;
        RECT 100.345 171.805 100.695 172.055 ;
        RECT 98.650 170.665 99.315 171.255 ;
        RECT 99.495 170.495 99.825 171.635 ;
        RECT 100.005 171.465 100.685 171.635 ;
        RECT 100.355 170.680 100.685 171.465 ;
        RECT 100.865 170.495 101.155 171.660 ;
        RECT 101.765 171.645 102.015 172.245 ;
        RECT 102.265 172.225 102.495 173.045 ;
        RECT 103.165 172.665 103.495 173.045 ;
        RECT 102.720 172.495 102.995 172.635 ;
        RECT 103.665 172.495 103.875 172.665 ;
        RECT 102.720 172.305 103.875 172.495 ;
        RECT 104.045 172.495 104.375 172.875 ;
        RECT 104.565 172.665 104.895 173.045 ;
        RECT 104.045 172.290 104.895 172.495 ;
        RECT 102.185 171.805 102.515 172.055 ;
        RECT 102.715 171.680 102.975 172.135 ;
        RECT 103.230 172.025 103.815 172.105 ;
        RECT 103.225 171.855 103.815 172.025 ;
        RECT 103.230 171.730 103.815 171.855 ;
        RECT 101.385 170.495 101.595 171.635 ;
        RECT 101.765 170.665 102.095 171.645 ;
        RECT 102.265 170.495 102.495 171.635 ;
        RECT 102.720 170.495 103.045 171.480 ;
        RECT 103.230 171.145 103.435 171.730 ;
        RECT 103.985 171.515 104.395 172.120 ;
        RECT 104.565 171.800 104.895 172.290 ;
        RECT 104.565 171.345 104.735 171.800 ;
        RECT 103.615 171.125 104.735 171.345 ;
        RECT 103.615 170.665 103.875 171.125 ;
        RECT 104.045 170.495 104.895 170.945 ;
        RECT 105.065 170.665 105.310 172.875 ;
        RECT 105.495 172.245 105.735 173.045 ;
        RECT 106.015 172.565 106.315 173.045 ;
        RECT 106.485 172.395 106.745 172.850 ;
        RECT 106.915 172.565 107.175 173.045 ;
        RECT 107.355 172.395 107.615 172.850 ;
        RECT 107.785 172.565 108.035 173.045 ;
        RECT 108.215 172.395 108.475 172.850 ;
        RECT 108.645 172.565 108.895 173.045 ;
        RECT 109.075 172.395 109.335 172.850 ;
        RECT 109.505 172.565 109.750 173.045 ;
        RECT 109.920 172.395 110.195 172.850 ;
        RECT 110.365 172.565 110.610 173.045 ;
        RECT 110.780 172.395 111.040 172.850 ;
        RECT 111.210 172.565 111.470 173.045 ;
        RECT 111.640 172.395 111.900 172.850 ;
        RECT 112.070 172.565 112.330 173.045 ;
        RECT 112.500 172.395 112.760 172.850 ;
        RECT 112.930 172.485 113.190 173.045 ;
        RECT 106.015 172.225 112.760 172.395 ;
        RECT 106.015 171.635 107.180 172.225 ;
        RECT 113.360 172.055 113.610 172.865 ;
        RECT 113.790 172.520 114.050 173.045 ;
        RECT 114.220 172.055 114.470 172.865 ;
        RECT 114.650 172.535 114.955 173.045 ;
        RECT 107.350 171.805 114.470 172.055 ;
        RECT 114.640 171.805 114.955 172.365 ;
        RECT 115.125 172.275 117.715 173.045 ;
        RECT 118.530 172.565 118.700 173.045 ;
        RECT 118.870 172.395 119.200 172.865 ;
        RECT 119.370 172.565 119.540 173.045 ;
        RECT 119.710 172.395 120.040 172.865 ;
        RECT 105.495 170.495 105.750 171.495 ;
        RECT 106.015 171.410 112.760 171.635 ;
        RECT 106.015 170.495 106.285 171.240 ;
        RECT 106.455 170.670 106.745 171.410 ;
        RECT 107.355 171.395 112.760 171.410 ;
        RECT 106.915 170.500 107.170 171.225 ;
        RECT 107.355 170.670 107.615 171.395 ;
        RECT 107.785 170.500 108.030 171.225 ;
        RECT 108.215 170.670 108.475 171.395 ;
        RECT 108.645 170.500 108.890 171.225 ;
        RECT 109.075 170.670 109.335 171.395 ;
        RECT 109.505 170.500 109.750 171.225 ;
        RECT 109.920 170.670 110.180 171.395 ;
        RECT 110.350 170.500 110.610 171.225 ;
        RECT 110.780 170.670 111.040 171.395 ;
        RECT 111.210 170.500 111.470 171.225 ;
        RECT 111.640 170.670 111.900 171.395 ;
        RECT 112.070 170.500 112.330 171.225 ;
        RECT 112.500 170.670 112.760 171.395 ;
        RECT 112.930 170.500 113.190 171.295 ;
        RECT 113.360 170.670 113.610 171.805 ;
        RECT 106.915 170.495 113.190 170.500 ;
        RECT 113.790 170.495 114.050 171.305 ;
        RECT 114.225 170.665 114.470 171.805 ;
        RECT 115.125 171.755 116.335 172.275 ;
        RECT 118.345 172.225 120.040 172.395 ;
        RECT 120.250 172.305 120.420 173.045 ;
        RECT 120.635 172.305 120.965 172.840 ;
        RECT 121.135 172.535 121.375 173.045 ;
        RECT 121.835 172.665 123.845 172.875 ;
        RECT 116.505 171.585 117.715 172.105 ;
        RECT 114.650 170.495 114.945 171.305 ;
        RECT 115.125 170.495 117.715 171.585 ;
        RECT 118.345 171.635 118.690 172.225 ;
        RECT 118.860 171.885 120.070 172.055 ;
        RECT 119.865 171.635 120.070 171.885 ;
        RECT 120.240 171.805 120.615 172.135 ;
        RECT 120.785 171.635 120.965 172.305 ;
        RECT 121.135 171.805 121.390 172.365 ;
        RECT 121.835 172.245 122.085 172.665 ;
        RECT 122.255 172.325 123.425 172.495 ;
        RECT 123.175 172.055 123.425 172.325 ;
        RECT 123.595 172.415 123.845 172.665 ;
        RECT 124.015 172.585 124.185 173.045 ;
        RECT 124.355 172.415 124.685 172.875 ;
        RECT 124.855 172.585 125.025 173.045 ;
        RECT 125.195 172.415 125.530 172.875 ;
        RECT 123.595 172.225 125.530 172.415 ;
        RECT 126.625 172.320 126.915 173.045 ;
        RECT 127.135 172.535 127.535 173.045 ;
        RECT 128.110 172.430 128.280 172.875 ;
        RECT 128.450 172.645 129.185 173.045 ;
        RECT 129.355 172.475 129.525 172.875 ;
        RECT 129.760 172.600 130.190 173.045 ;
        RECT 127.145 172.195 127.410 172.365 ;
        RECT 127.605 172.195 127.870 172.365 ;
        RECT 128.110 172.260 128.460 172.430 ;
        RECT 121.565 171.805 123.005 172.055 ;
        RECT 123.175 171.635 123.710 172.055 ;
        RECT 123.890 171.805 125.510 172.055 ;
        RECT 118.345 171.465 119.200 171.635 ;
        RECT 119.865 171.465 121.325 171.635 ;
        RECT 118.870 171.295 119.200 171.465 ;
        RECT 118.530 170.495 118.700 171.295 ;
        RECT 118.870 171.125 120.040 171.295 ;
        RECT 118.870 170.665 119.200 171.125 ;
        RECT 119.370 170.495 119.540 170.955 ;
        RECT 119.710 170.665 120.040 171.125 ;
        RECT 120.250 170.495 120.420 171.295 ;
        RECT 120.965 170.665 121.325 171.465 ;
        RECT 122.255 171.465 125.105 171.635 ;
        RECT 121.835 170.495 122.085 171.295 ;
        RECT 122.255 170.665 122.585 171.465 ;
        RECT 122.755 170.495 122.925 171.295 ;
        RECT 123.095 170.665 123.425 171.465 ;
        RECT 123.595 170.495 123.765 171.295 ;
        RECT 123.935 170.665 124.265 171.465 ;
        RECT 124.435 170.495 124.605 171.295 ;
        RECT 124.775 170.665 125.105 171.465 ;
        RECT 125.275 170.495 125.530 171.635 ;
        RECT 126.625 170.495 126.915 171.660 ;
        RECT 127.150 171.475 127.410 172.195 ;
        RECT 127.610 171.775 127.870 172.195 ;
        RECT 127.610 171.475 128.090 171.775 ;
        RECT 127.175 171.125 128.105 171.295 ;
        RECT 127.175 170.665 127.345 171.125 ;
        RECT 127.515 170.495 127.765 170.955 ;
        RECT 127.935 170.875 128.105 171.125 ;
        RECT 128.290 171.235 128.460 172.260 ;
        RECT 128.630 172.305 129.525 172.475 ;
        RECT 130.360 172.320 130.615 172.875 ;
        RECT 128.630 171.585 128.800 172.305 ;
        RECT 129.005 172.025 129.295 172.135 ;
        RECT 128.985 171.855 129.295 172.025 ;
        RECT 129.005 171.755 129.295 171.855 ;
        RECT 128.630 171.415 129.165 171.585 ;
        RECT 129.465 171.515 129.795 172.135 ;
        RECT 130.020 171.805 130.275 172.135 ;
        RECT 128.290 171.065 128.700 171.235 ;
        RECT 128.995 171.225 129.165 171.415 ;
        RECT 130.020 171.325 130.190 171.805 ;
        RECT 130.445 171.605 130.615 172.320 ;
        RECT 130.785 172.200 130.955 173.045 ;
        RECT 131.235 172.435 131.565 172.855 ;
        RECT 131.735 172.605 132.010 173.045 ;
        RECT 132.215 172.435 132.545 172.855 ;
        RECT 133.025 172.685 133.875 173.045 ;
        RECT 134.045 172.495 134.265 172.875 ;
        RECT 131.235 172.255 133.820 172.435 ;
        RECT 131.225 171.855 131.560 172.085 ;
        RECT 131.750 172.025 132.200 172.085 ;
        RECT 131.745 171.855 132.200 172.025 ;
        RECT 132.370 171.855 132.840 172.085 ;
        RECT 133.010 171.855 133.340 172.085 ;
        RECT 128.470 170.930 128.700 171.065 ;
        RECT 129.430 171.155 130.190 171.325 ;
        RECT 129.430 170.930 129.600 171.155 ;
        RECT 127.935 170.705 128.265 170.875 ;
        RECT 128.470 170.760 129.600 170.930 ;
        RECT 128.470 170.665 128.640 170.760 ;
        RECT 129.860 170.495 130.190 170.895 ;
        RECT 130.360 170.665 130.615 171.605 ;
        RECT 130.785 170.495 130.955 171.685 ;
        RECT 133.510 171.640 133.820 172.255 ;
        RECT 131.235 171.470 133.820 171.640 ;
        RECT 131.235 170.805 131.565 171.470 ;
        RECT 132.025 171.110 133.365 171.290 ;
        RECT 132.025 170.665 132.355 171.110 ;
        RECT 132.590 170.495 132.865 170.940 ;
        RECT 133.035 170.665 133.365 171.110 ;
        RECT 133.565 170.495 133.820 171.300 ;
        RECT 134.035 170.795 134.265 172.495 ;
        RECT 134.435 172.225 134.730 173.045 ;
        RECT 134.905 172.295 136.115 173.045 ;
        RECT 134.435 170.495 134.730 171.640 ;
        RECT 134.905 171.585 135.425 172.125 ;
        RECT 135.595 171.755 136.115 172.295 ;
        RECT 134.905 170.495 136.115 171.585 ;
        RECT 23.500 170.325 136.200 170.495 ;
        RECT 23.585 169.235 24.795 170.325 ;
        RECT 23.585 168.525 24.105 169.065 ;
        RECT 24.275 168.695 24.795 169.235 ;
        RECT 24.970 169.175 25.230 170.325 ;
        RECT 25.405 169.250 25.660 170.155 ;
        RECT 25.830 169.565 26.160 170.325 ;
        RECT 26.375 169.395 26.545 170.155 ;
        RECT 23.585 167.775 24.795 168.525 ;
        RECT 24.970 167.775 25.230 168.615 ;
        RECT 25.405 168.520 25.575 169.250 ;
        RECT 25.830 169.225 26.545 169.395 ;
        RECT 27.725 169.250 27.995 170.155 ;
        RECT 28.165 169.565 28.495 170.325 ;
        RECT 28.675 169.395 28.845 170.155 ;
        RECT 29.105 169.890 34.450 170.325 ;
        RECT 25.830 169.015 26.000 169.225 ;
        RECT 25.745 168.685 26.000 169.015 ;
        RECT 25.405 167.945 25.660 168.520 ;
        RECT 25.830 168.495 26.000 168.685 ;
        RECT 26.280 168.675 26.635 169.045 ;
        RECT 25.830 168.325 26.545 168.495 ;
        RECT 25.830 167.775 26.160 168.155 ;
        RECT 26.375 167.945 26.545 168.325 ;
        RECT 27.725 168.450 27.895 169.250 ;
        RECT 28.180 169.225 28.845 169.395 ;
        RECT 28.180 169.080 28.350 169.225 ;
        RECT 28.065 168.750 28.350 169.080 ;
        RECT 28.180 168.495 28.350 168.750 ;
        RECT 28.585 168.675 28.915 169.045 ;
        RECT 27.725 167.945 27.985 168.450 ;
        RECT 28.180 168.325 28.845 168.495 ;
        RECT 28.165 167.775 28.495 168.155 ;
        RECT 28.675 167.945 28.845 168.325 ;
        RECT 30.690 168.320 31.030 169.150 ;
        RECT 32.510 168.640 32.860 169.890 ;
        RECT 34.625 169.235 36.295 170.325 ;
        RECT 34.625 168.545 35.375 169.065 ;
        RECT 35.545 168.715 36.295 169.235 ;
        RECT 36.465 169.160 36.755 170.325 ;
        RECT 36.925 169.235 38.595 170.325 ;
        RECT 38.965 169.655 39.245 170.325 ;
        RECT 39.415 169.435 39.715 169.985 ;
        RECT 39.915 169.605 40.245 170.325 ;
        RECT 40.435 169.605 40.895 170.155 ;
        RECT 36.925 168.545 37.675 169.065 ;
        RECT 37.845 168.715 38.595 169.235 ;
        RECT 38.780 169.015 39.045 169.375 ;
        RECT 39.415 169.265 40.355 169.435 ;
        RECT 40.185 169.015 40.355 169.265 ;
        RECT 38.780 168.765 39.455 169.015 ;
        RECT 39.675 168.765 40.015 169.015 ;
        RECT 40.185 168.685 40.475 169.015 ;
        RECT 40.185 168.595 40.355 168.685 ;
        RECT 29.105 167.775 34.450 168.320 ;
        RECT 34.625 167.775 36.295 168.545 ;
        RECT 36.465 167.775 36.755 168.500 ;
        RECT 36.925 167.775 38.595 168.545 ;
        RECT 38.965 168.405 40.355 168.595 ;
        RECT 38.965 168.045 39.295 168.405 ;
        RECT 40.645 168.235 40.895 169.605 ;
        RECT 39.915 167.775 40.165 168.235 ;
        RECT 40.335 167.945 40.895 168.235 ;
        RECT 41.065 168.720 41.345 170.155 ;
        RECT 41.515 169.550 42.225 170.325 ;
        RECT 42.395 169.380 42.725 170.155 ;
        RECT 41.575 169.165 42.725 169.380 ;
        RECT 41.065 167.945 41.405 168.720 ;
        RECT 41.575 168.595 41.860 169.165 ;
        RECT 42.045 168.765 42.515 168.995 ;
        RECT 42.920 168.965 43.135 170.080 ;
        RECT 43.315 169.605 43.645 170.325 ;
        RECT 43.915 169.395 44.085 170.155 ;
        RECT 44.300 169.565 44.630 170.325 ;
        RECT 43.425 168.965 43.655 169.305 ;
        RECT 43.915 169.225 44.630 169.395 ;
        RECT 44.800 169.250 45.055 170.155 ;
        RECT 42.685 168.785 43.135 168.965 ;
        RECT 42.685 168.765 43.015 168.785 ;
        RECT 43.325 168.765 43.655 168.965 ;
        RECT 43.825 168.675 44.180 169.045 ;
        RECT 44.460 169.015 44.630 169.225 ;
        RECT 44.460 168.685 44.715 169.015 ;
        RECT 41.575 168.405 42.285 168.595 ;
        RECT 41.985 168.265 42.285 168.405 ;
        RECT 42.475 168.405 43.655 168.595 ;
        RECT 44.460 168.495 44.630 168.685 ;
        RECT 44.885 168.520 45.055 169.250 ;
        RECT 45.230 169.175 45.490 170.325 ;
        RECT 45.850 169.355 46.240 169.530 ;
        RECT 46.725 169.525 47.055 170.325 ;
        RECT 47.225 169.535 47.760 170.155 ;
        RECT 47.965 169.890 53.310 170.325 ;
        RECT 45.850 169.185 47.275 169.355 ;
        RECT 42.475 168.325 42.805 168.405 ;
        RECT 41.985 168.255 42.300 168.265 ;
        RECT 41.985 168.245 42.310 168.255 ;
        RECT 41.985 168.240 42.320 168.245 ;
        RECT 41.575 167.775 41.745 168.235 ;
        RECT 41.985 168.230 42.325 168.240 ;
        RECT 41.985 168.225 42.330 168.230 ;
        RECT 41.985 168.215 42.335 168.225 ;
        RECT 41.985 168.210 42.340 168.215 ;
        RECT 41.985 167.945 42.345 168.210 ;
        RECT 42.975 167.775 43.145 168.235 ;
        RECT 43.315 167.945 43.655 168.405 ;
        RECT 43.915 168.325 44.630 168.495 ;
        RECT 43.915 167.945 44.085 168.325 ;
        RECT 44.300 167.775 44.630 168.155 ;
        RECT 44.800 167.945 45.055 168.520 ;
        RECT 45.230 167.775 45.490 168.615 ;
        RECT 45.725 168.455 46.080 169.015 ;
        RECT 46.250 168.285 46.420 169.185 ;
        RECT 46.590 168.455 46.855 169.015 ;
        RECT 47.105 168.685 47.275 169.185 ;
        RECT 47.445 168.515 47.760 169.535 ;
        RECT 45.830 167.775 46.070 168.285 ;
        RECT 46.250 167.955 46.530 168.285 ;
        RECT 46.760 167.775 46.975 168.285 ;
        RECT 47.145 167.945 47.760 168.515 ;
        RECT 49.550 168.320 49.890 169.150 ;
        RECT 51.370 168.640 51.720 169.890 ;
        RECT 53.485 169.235 55.155 170.325 ;
        RECT 53.485 168.545 54.235 169.065 ;
        RECT 54.405 168.715 55.155 169.235 ;
        RECT 55.810 169.355 56.110 169.550 ;
        RECT 56.280 169.525 56.535 170.325 ;
        RECT 56.735 169.695 57.065 170.155 ;
        RECT 57.235 169.865 57.810 170.325 ;
        RECT 57.980 169.695 58.335 170.155 ;
        RECT 56.735 169.525 58.335 169.695 ;
        RECT 55.810 169.185 57.060 169.355 ;
        RECT 47.965 167.775 53.310 168.320 ;
        RECT 53.485 167.775 55.155 168.545 ;
        RECT 55.810 168.530 55.980 169.185 ;
        RECT 56.155 168.685 56.500 169.015 ;
        RECT 56.730 168.765 57.060 169.185 ;
        RECT 57.230 168.595 57.510 169.525 ;
        RECT 57.690 168.965 57.880 169.345 ;
        RECT 58.060 169.185 58.335 169.525 ;
        RECT 58.505 169.185 58.835 170.325 ;
        RECT 59.465 169.185 59.745 170.325 ;
        RECT 59.915 169.175 60.245 170.155 ;
        RECT 60.415 169.185 60.675 170.325 ;
        RECT 60.845 169.235 62.055 170.325 ;
        RECT 57.685 168.795 58.835 168.965 ;
        RECT 57.690 168.765 58.835 168.795 ;
        RECT 59.475 168.745 59.810 169.015 ;
        RECT 55.810 168.200 56.045 168.530 ;
        RECT 56.215 167.775 56.545 168.515 ;
        RECT 56.780 168.155 57.055 168.595 ;
        RECT 57.230 168.495 57.555 168.595 ;
        RECT 57.225 168.325 57.555 168.495 ;
        RECT 57.725 168.385 58.835 168.595 ;
        RECT 59.980 168.575 60.150 169.175 ;
        RECT 60.320 168.765 60.655 169.015 ;
        RECT 57.725 168.155 57.975 168.385 ;
        RECT 56.780 167.945 57.975 168.155 ;
        RECT 58.145 167.775 58.315 168.215 ;
        RECT 58.485 167.945 58.835 168.385 ;
        RECT 59.465 167.775 59.775 168.575 ;
        RECT 59.980 167.945 60.675 168.575 ;
        RECT 60.845 168.525 61.365 169.065 ;
        RECT 61.535 168.695 62.055 169.235 ;
        RECT 62.225 169.160 62.515 170.325 ;
        RECT 62.685 169.235 65.275 170.325 ;
        RECT 62.685 168.545 63.895 169.065 ;
        RECT 64.065 168.715 65.275 169.235 ;
        RECT 65.905 169.185 66.245 170.155 ;
        RECT 66.415 169.185 66.585 170.325 ;
        RECT 66.855 169.525 67.105 170.325 ;
        RECT 67.750 169.355 68.080 170.155 ;
        RECT 68.380 169.525 68.710 170.325 ;
        RECT 68.880 169.355 69.210 170.155 ;
        RECT 69.585 169.945 70.845 170.155 ;
        RECT 69.585 169.525 69.845 169.945 ;
        RECT 66.775 169.185 69.210 169.355 ;
        RECT 70.015 169.475 70.365 169.775 ;
        RECT 70.595 169.645 70.845 169.945 ;
        RECT 71.055 169.825 71.305 170.325 ;
        RECT 71.515 169.645 71.685 170.155 ;
        RECT 70.595 169.475 71.685 169.645 ;
        RECT 65.905 168.575 66.080 169.185 ;
        RECT 66.775 168.935 66.945 169.185 ;
        RECT 66.250 168.765 66.945 168.935 ;
        RECT 67.120 168.765 67.540 168.965 ;
        RECT 67.710 168.765 68.040 168.965 ;
        RECT 68.210 168.765 68.540 168.965 ;
        RECT 60.845 167.775 62.055 168.525 ;
        RECT 62.225 167.775 62.515 168.500 ;
        RECT 62.685 167.775 65.275 168.545 ;
        RECT 65.905 167.945 66.245 168.575 ;
        RECT 66.415 167.775 66.665 168.575 ;
        RECT 66.855 168.425 68.080 168.595 ;
        RECT 66.855 167.945 67.185 168.425 ;
        RECT 67.355 167.775 67.580 168.235 ;
        RECT 67.750 167.945 68.080 168.425 ;
        RECT 68.710 168.555 68.880 169.185 ;
        RECT 69.065 168.765 69.415 169.015 ;
        RECT 69.585 168.685 69.845 169.015 ;
        RECT 68.710 167.945 69.210 168.555 ;
        RECT 70.015 168.495 70.185 169.475 ;
        RECT 71.515 169.435 71.685 169.475 ;
        RECT 70.355 169.115 70.755 169.305 ;
        RECT 71.855 169.185 72.195 170.325 ;
        RECT 72.990 169.355 73.380 169.530 ;
        RECT 73.865 169.525 74.195 170.325 ;
        RECT 74.365 169.535 74.900 170.155 ;
        RECT 72.990 169.185 74.415 169.355 ;
        RECT 70.355 168.685 70.525 169.115 ;
        RECT 70.730 168.765 71.095 168.945 ;
        RECT 70.015 168.325 70.665 168.495 ;
        RECT 69.595 167.775 69.925 168.155 ;
        RECT 70.415 167.985 70.665 168.325 ;
        RECT 70.905 168.455 71.095 168.765 ;
        RECT 71.305 168.685 71.665 169.015 ;
        RECT 71.835 168.705 72.250 169.015 ;
        RECT 70.905 168.035 71.205 168.455 ;
        RECT 71.465 168.105 71.665 168.685 ;
        RECT 71.855 167.775 72.195 168.495 ;
        RECT 72.865 168.455 73.220 169.015 ;
        RECT 73.390 168.285 73.560 169.185 ;
        RECT 73.730 168.455 73.995 169.015 ;
        RECT 74.245 168.685 74.415 169.185 ;
        RECT 74.585 168.515 74.900 169.535 ;
        RECT 75.105 169.235 78.615 170.325 ;
        RECT 72.970 167.775 73.210 168.285 ;
        RECT 73.390 167.955 73.670 168.285 ;
        RECT 73.900 167.775 74.115 168.285 ;
        RECT 74.285 167.945 74.900 168.515 ;
        RECT 75.105 168.545 76.755 169.065 ;
        RECT 76.925 168.715 78.615 169.235 ;
        RECT 79.715 169.375 79.990 170.145 ;
        RECT 80.160 169.715 80.490 170.145 ;
        RECT 80.660 169.885 80.855 170.325 ;
        RECT 81.035 169.715 81.365 170.145 ;
        RECT 80.160 169.545 81.365 169.715 ;
        RECT 79.715 169.185 80.300 169.375 ;
        RECT 80.470 169.215 81.365 169.545 ;
        RECT 82.015 169.715 82.345 170.145 ;
        RECT 82.525 169.885 82.720 170.325 ;
        RECT 82.890 169.715 83.220 170.145 ;
        RECT 82.015 169.545 83.220 169.715 ;
        RECT 82.015 169.215 82.910 169.545 ;
        RECT 83.390 169.375 83.665 170.145 ;
        RECT 75.105 167.775 78.615 168.545 ;
        RECT 79.715 168.365 79.955 169.015 ;
        RECT 80.125 168.515 80.300 169.185 ;
        RECT 83.080 169.185 83.665 169.375 ;
        RECT 80.470 168.685 80.885 169.015 ;
        RECT 81.065 168.685 81.360 169.015 ;
        RECT 82.020 168.685 82.315 169.015 ;
        RECT 82.495 168.685 82.910 169.015 ;
        RECT 80.125 168.335 80.455 168.515 ;
        RECT 79.730 167.775 80.060 168.165 ;
        RECT 80.230 167.955 80.455 168.335 ;
        RECT 80.655 168.065 80.885 168.685 ;
        RECT 81.065 167.775 81.365 168.505 ;
        RECT 82.015 167.775 82.315 168.505 ;
        RECT 82.495 168.065 82.725 168.685 ;
        RECT 83.080 168.515 83.255 169.185 ;
        RECT 82.925 168.335 83.255 168.515 ;
        RECT 83.425 168.365 83.665 169.015 ;
        RECT 82.925 167.955 83.150 168.335 ;
        RECT 83.320 167.775 83.650 168.165 ;
        RECT 83.845 167.945 84.595 170.155 ;
        RECT 85.230 169.815 86.885 170.105 ;
        RECT 85.230 169.475 86.820 169.645 ;
        RECT 87.055 169.525 87.335 170.325 ;
        RECT 85.230 169.185 85.550 169.475 ;
        RECT 86.650 169.355 86.820 169.475 ;
        RECT 85.230 168.445 85.580 169.015 ;
        RECT 85.750 168.685 86.460 169.305 ;
        RECT 86.650 169.185 87.375 169.355 ;
        RECT 87.545 169.185 87.815 170.155 ;
        RECT 87.205 169.015 87.375 169.185 ;
        RECT 86.630 168.685 87.035 169.015 ;
        RECT 87.205 168.685 87.475 169.015 ;
        RECT 87.205 168.515 87.375 168.685 ;
        RECT 85.765 168.345 87.375 168.515 ;
        RECT 87.645 168.450 87.815 169.185 ;
        RECT 87.985 169.160 88.275 170.325 ;
        RECT 88.495 169.545 88.760 170.325 ;
        RECT 89.310 169.945 89.685 170.325 ;
        RECT 89.855 169.985 91.025 170.155 ;
        RECT 89.855 169.945 90.185 169.985 ;
        RECT 88.995 169.725 89.165 169.855 ;
        RECT 90.295 169.775 90.525 169.815 ;
        RECT 89.910 169.725 90.525 169.775 ;
        RECT 88.995 169.525 90.525 169.725 ;
        RECT 89.645 169.485 90.525 169.525 ;
        RECT 88.445 169.315 89.505 169.355 ;
        RECT 90.695 169.315 91.025 169.985 ;
        RECT 88.445 169.185 91.025 169.315 ;
        RECT 88.445 168.515 88.615 169.185 ;
        RECT 89.280 169.135 91.025 169.185 ;
        RECT 91.205 169.475 91.465 170.155 ;
        RECT 91.635 169.545 91.885 170.325 ;
        RECT 92.135 169.775 92.385 170.155 ;
        RECT 92.555 169.945 92.910 170.325 ;
        RECT 93.915 169.935 94.250 170.155 ;
        RECT 93.515 169.775 93.745 169.815 ;
        RECT 92.135 169.575 93.745 169.775 ;
        RECT 92.135 169.565 92.970 169.575 ;
        RECT 93.560 169.485 93.745 169.575 ;
        RECT 88.785 168.685 89.110 169.015 ;
        RECT 89.280 168.765 89.630 168.965 ;
        RECT 85.235 167.775 85.565 168.275 ;
        RECT 85.765 167.995 85.935 168.345 ;
        RECT 86.135 167.775 86.465 168.175 ;
        RECT 86.635 167.995 86.805 168.345 ;
        RECT 86.975 167.775 87.355 168.175 ;
        RECT 87.545 168.105 87.815 168.450 ;
        RECT 87.985 167.775 88.275 168.500 ;
        RECT 88.445 168.345 89.175 168.515 ;
        RECT 89.420 168.365 89.630 168.765 ;
        RECT 89.880 168.765 90.355 168.965 ;
        RECT 89.880 168.365 90.130 168.765 ;
        RECT 90.545 168.455 90.995 168.965 ;
        RECT 88.995 168.195 89.175 168.345 ;
        RECT 88.485 167.775 88.815 168.175 ;
        RECT 88.995 167.945 90.300 168.195 ;
        RECT 90.575 167.775 91.025 168.285 ;
        RECT 91.205 168.275 91.375 169.475 ;
        RECT 93.075 169.375 93.405 169.405 ;
        RECT 91.605 169.315 93.405 169.375 ;
        RECT 93.995 169.315 94.250 169.935 ;
        RECT 91.545 169.205 94.250 169.315 ;
        RECT 91.545 169.170 91.745 169.205 ;
        RECT 91.545 168.595 91.715 169.170 ;
        RECT 93.075 169.145 94.250 169.205 ;
        RECT 94.425 169.215 94.685 170.155 ;
        RECT 94.855 169.925 95.185 170.325 ;
        RECT 96.330 170.060 96.585 170.155 ;
        RECT 95.445 169.890 96.585 170.060 ;
        RECT 96.755 169.945 97.085 170.115 ;
        RECT 95.445 169.665 95.615 169.890 ;
        RECT 94.855 169.495 95.615 169.665 ;
        RECT 96.330 169.755 96.585 169.890 ;
        RECT 91.945 168.730 92.355 169.035 ;
        RECT 92.525 168.765 92.855 168.975 ;
        RECT 91.545 168.475 91.815 168.595 ;
        RECT 91.545 168.430 92.390 168.475 ;
        RECT 91.635 168.305 92.390 168.430 ;
        RECT 92.645 168.365 92.855 168.765 ;
        RECT 93.100 168.765 93.575 168.975 ;
        RECT 93.765 168.765 94.255 168.965 ;
        RECT 93.100 168.365 93.320 168.765 ;
        RECT 91.205 167.945 91.465 168.275 ;
        RECT 92.220 168.155 92.390 168.305 ;
        RECT 91.635 167.775 91.965 168.135 ;
        RECT 92.220 167.945 93.520 168.155 ;
        RECT 93.795 167.775 94.250 168.540 ;
        RECT 94.425 168.500 94.600 169.215 ;
        RECT 94.855 169.015 95.025 169.495 ;
        RECT 95.880 169.405 96.050 169.595 ;
        RECT 96.330 169.585 96.740 169.755 ;
        RECT 94.770 168.685 95.025 169.015 ;
        RECT 95.250 168.685 95.580 169.305 ;
        RECT 95.880 169.235 96.400 169.405 ;
        RECT 95.750 168.685 96.040 169.065 ;
        RECT 96.230 168.515 96.400 169.235 ;
        RECT 94.425 167.945 94.685 168.500 ;
        RECT 95.520 168.345 96.400 168.515 ;
        RECT 96.570 168.560 96.740 169.585 ;
        RECT 96.915 169.695 97.085 169.945 ;
        RECT 97.255 169.865 97.505 170.325 ;
        RECT 97.675 169.695 97.855 170.155 ;
        RECT 96.915 169.525 97.855 169.695 ;
        RECT 98.575 169.715 98.905 170.145 ;
        RECT 99.085 169.885 99.280 170.325 ;
        RECT 99.450 169.715 99.780 170.145 ;
        RECT 98.575 169.545 99.780 169.715 ;
        RECT 96.940 169.045 97.420 169.345 ;
        RECT 96.570 168.390 96.920 168.560 ;
        RECT 97.160 168.455 97.420 169.045 ;
        RECT 97.620 168.455 97.880 169.345 ;
        RECT 98.575 169.215 99.470 169.545 ;
        RECT 99.950 169.375 100.225 170.145 ;
        RECT 99.640 169.185 100.225 169.375 ;
        RECT 100.405 169.185 100.745 170.155 ;
        RECT 100.915 169.185 101.085 170.325 ;
        RECT 101.355 169.525 101.605 170.325 ;
        RECT 102.250 169.355 102.580 170.155 ;
        RECT 102.880 169.525 103.210 170.325 ;
        RECT 103.380 169.355 103.710 170.155 ;
        RECT 105.060 169.485 105.265 170.325 ;
        RECT 105.475 169.985 106.565 170.155 ;
        RECT 105.475 169.475 105.725 169.985 ;
        RECT 106.315 169.815 106.565 169.985 ;
        RECT 106.735 169.815 106.985 170.325 ;
        RECT 105.895 169.645 106.145 169.815 ;
        RECT 107.155 169.655 107.445 170.155 ;
        RECT 107.615 169.825 108.345 170.325 ;
        RECT 108.935 169.825 109.185 170.325 ;
        RECT 108.515 169.655 108.765 169.815 ;
        RECT 109.355 169.655 109.605 170.155 ;
        RECT 107.155 169.645 107.535 169.655 ;
        RECT 105.895 169.475 107.535 169.645 ;
        RECT 101.275 169.185 103.710 169.355 ;
        RECT 98.580 168.685 98.875 169.015 ;
        RECT 99.055 168.685 99.470 169.015 ;
        RECT 94.855 167.775 95.285 168.220 ;
        RECT 95.520 167.945 95.690 168.345 ;
        RECT 95.860 167.775 96.580 168.175 ;
        RECT 96.750 167.945 96.920 168.390 ;
        RECT 97.495 167.775 97.895 168.285 ;
        RECT 98.575 167.775 98.875 168.505 ;
        RECT 99.055 168.065 99.285 168.685 ;
        RECT 99.640 168.515 99.815 169.185 ;
        RECT 99.485 168.335 99.815 168.515 ;
        RECT 99.985 168.365 100.225 169.015 ;
        RECT 100.405 168.575 100.580 169.185 ;
        RECT 101.275 168.935 101.445 169.185 ;
        RECT 100.750 168.765 101.445 168.935 ;
        RECT 101.620 168.765 102.040 168.965 ;
        RECT 102.210 168.765 102.540 168.965 ;
        RECT 102.710 168.765 103.040 168.965 ;
        RECT 99.485 167.955 99.710 168.335 ;
        RECT 99.880 167.775 100.210 168.165 ;
        RECT 100.405 167.945 100.745 168.575 ;
        RECT 100.915 167.775 101.165 168.575 ;
        RECT 101.355 168.425 102.580 168.595 ;
        RECT 101.355 167.945 101.685 168.425 ;
        RECT 101.855 167.775 102.080 168.235 ;
        RECT 102.250 167.945 102.580 168.425 ;
        RECT 103.210 168.555 103.380 169.185 ;
        RECT 105.005 169.135 106.815 169.305 ;
        RECT 103.565 168.765 103.915 169.015 ;
        RECT 105.005 168.765 105.495 169.135 ;
        RECT 105.725 168.765 106.265 168.965 ;
        RECT 106.485 168.765 106.815 169.135 ;
        RECT 106.985 169.105 107.535 169.475 ;
        RECT 107.875 169.475 109.605 169.655 ;
        RECT 109.775 169.485 110.025 170.325 ;
        RECT 110.195 169.645 110.445 170.155 ;
        RECT 110.615 169.855 110.865 170.325 ;
        RECT 111.035 169.645 111.285 170.155 ;
        RECT 110.195 169.475 111.285 169.645 ;
        RECT 111.455 169.515 111.705 170.325 ;
        RECT 106.985 168.765 107.365 169.105 ;
        RECT 107.875 168.935 108.065 169.475 ;
        RECT 111.035 169.345 111.285 169.475 ;
        RECT 107.535 168.765 108.065 168.935 ;
        RECT 108.235 169.135 109.885 169.305 ;
        RECT 108.235 168.765 108.565 169.135 ;
        RECT 108.735 168.765 109.355 168.965 ;
        RECT 109.525 168.765 109.885 169.135 ;
        RECT 110.085 168.935 110.375 169.305 ;
        RECT 111.035 169.105 111.830 169.345 ;
        RECT 112.405 169.185 112.635 170.325 ;
        RECT 112.805 169.175 113.135 170.155 ;
        RECT 113.305 169.185 113.515 170.325 ;
        RECT 110.085 168.765 111.355 168.935 ;
        RECT 103.210 167.945 103.710 168.555 ;
        RECT 105.015 168.425 106.945 168.595 ;
        RECT 105.015 168.415 106.185 168.425 ;
        RECT 105.015 167.945 105.345 168.415 ;
        RECT 105.515 167.775 105.685 168.245 ;
        RECT 105.855 167.945 106.185 168.415 ;
        RECT 106.355 167.775 106.525 168.245 ;
        RECT 106.695 168.165 106.945 168.425 ;
        RECT 107.115 168.505 107.365 168.765 ;
        RECT 107.875 168.595 108.065 168.765 ;
        RECT 111.525 168.595 111.830 169.105 ;
        RECT 112.385 168.765 112.715 169.015 ;
        RECT 107.115 168.335 107.445 168.505 ;
        RECT 107.875 168.415 109.225 168.595 ;
        RECT 108.895 168.335 109.225 168.415 ;
        RECT 106.695 167.945 107.865 168.165 ;
        RECT 108.135 167.775 108.305 168.245 ;
        RECT 109.395 168.165 109.645 168.585 ;
        RECT 108.475 167.995 109.645 168.165 ;
        RECT 109.815 167.775 109.985 168.585 ;
        RECT 110.155 168.415 111.830 168.595 ;
        RECT 110.155 167.965 110.485 168.415 ;
        RECT 110.655 167.775 110.825 168.245 ;
        RECT 110.995 167.965 111.325 168.415 ;
        RECT 111.495 167.775 111.665 168.245 ;
        RECT 112.405 167.775 112.635 168.595 ;
        RECT 112.885 168.575 113.135 169.175 ;
        RECT 113.745 169.160 114.035 170.325 ;
        RECT 114.215 169.515 114.510 170.325 ;
        RECT 114.690 169.015 114.935 170.155 ;
        RECT 115.110 169.515 115.370 170.325 ;
        RECT 115.970 170.320 122.245 170.325 ;
        RECT 115.550 169.015 115.800 170.150 ;
        RECT 115.970 169.525 116.230 170.320 ;
        RECT 116.400 169.425 116.660 170.150 ;
        RECT 116.830 169.595 117.090 170.320 ;
        RECT 117.260 169.425 117.520 170.150 ;
        RECT 117.690 169.595 117.950 170.320 ;
        RECT 118.120 169.425 118.380 170.150 ;
        RECT 118.550 169.595 118.810 170.320 ;
        RECT 118.980 169.425 119.240 170.150 ;
        RECT 119.410 169.595 119.655 170.320 ;
        RECT 119.825 169.425 120.085 170.150 ;
        RECT 120.270 169.595 120.515 170.320 ;
        RECT 120.685 169.425 120.945 170.150 ;
        RECT 121.130 169.595 121.375 170.320 ;
        RECT 121.545 169.425 121.805 170.150 ;
        RECT 121.990 169.595 122.245 170.320 ;
        RECT 116.400 169.410 121.805 169.425 ;
        RECT 122.415 169.410 122.705 170.150 ;
        RECT 122.875 169.580 123.145 170.325 ;
        RECT 116.400 169.185 123.145 169.410 ;
        RECT 124.385 169.185 124.595 170.325 ;
        RECT 112.805 167.945 113.135 168.575 ;
        RECT 113.305 167.775 113.515 168.595 ;
        RECT 113.745 167.775 114.035 168.500 ;
        RECT 114.205 168.455 114.520 169.015 ;
        RECT 114.690 168.765 121.810 169.015 ;
        RECT 114.205 167.775 114.510 168.285 ;
        RECT 114.690 167.955 114.940 168.765 ;
        RECT 115.110 167.775 115.370 168.300 ;
        RECT 115.550 167.955 115.800 168.765 ;
        RECT 121.980 168.595 123.145 169.185 ;
        RECT 124.765 169.175 125.095 170.155 ;
        RECT 125.265 169.185 125.495 170.325 ;
        RECT 125.715 169.515 126.010 170.325 ;
        RECT 116.400 168.425 123.145 168.595 ;
        RECT 115.970 167.775 116.230 168.335 ;
        RECT 116.400 167.970 116.660 168.425 ;
        RECT 116.830 167.775 117.090 168.255 ;
        RECT 117.260 167.970 117.520 168.425 ;
        RECT 117.690 167.775 117.950 168.255 ;
        RECT 118.120 167.970 118.380 168.425 ;
        RECT 118.550 167.775 118.795 168.255 ;
        RECT 118.965 167.970 119.240 168.425 ;
        RECT 119.410 167.775 119.655 168.255 ;
        RECT 119.825 167.970 120.085 168.425 ;
        RECT 120.265 167.775 120.515 168.255 ;
        RECT 120.685 167.970 120.945 168.425 ;
        RECT 121.125 167.775 121.375 168.255 ;
        RECT 121.545 167.970 121.805 168.425 ;
        RECT 121.985 167.775 122.245 168.255 ;
        RECT 122.415 167.970 122.675 168.425 ;
        RECT 122.845 167.775 123.145 168.255 ;
        RECT 124.385 167.775 124.595 168.595 ;
        RECT 124.765 168.575 125.015 169.175 ;
        RECT 126.190 169.015 126.435 170.155 ;
        RECT 126.610 169.515 126.870 170.325 ;
        RECT 127.470 170.320 133.745 170.325 ;
        RECT 127.050 169.015 127.300 170.150 ;
        RECT 127.470 169.525 127.730 170.320 ;
        RECT 127.900 169.425 128.160 170.150 ;
        RECT 128.330 169.595 128.590 170.320 ;
        RECT 128.760 169.425 129.020 170.150 ;
        RECT 129.190 169.595 129.450 170.320 ;
        RECT 129.620 169.425 129.880 170.150 ;
        RECT 130.050 169.595 130.310 170.320 ;
        RECT 130.480 169.425 130.740 170.150 ;
        RECT 130.910 169.595 131.155 170.320 ;
        RECT 131.325 169.425 131.585 170.150 ;
        RECT 131.770 169.595 132.015 170.320 ;
        RECT 132.185 169.425 132.445 170.150 ;
        RECT 132.630 169.595 132.875 170.320 ;
        RECT 133.045 169.425 133.305 170.150 ;
        RECT 133.490 169.595 133.745 170.320 ;
        RECT 127.900 169.410 133.305 169.425 ;
        RECT 133.915 169.410 134.205 170.150 ;
        RECT 134.375 169.580 134.645 170.325 ;
        RECT 127.900 169.185 134.645 169.410 ;
        RECT 125.185 168.765 125.515 169.015 ;
        RECT 124.765 167.945 125.095 168.575 ;
        RECT 125.265 167.775 125.495 168.595 ;
        RECT 125.705 168.455 126.020 169.015 ;
        RECT 126.190 168.765 133.310 169.015 ;
        RECT 125.705 167.775 126.010 168.285 ;
        RECT 126.190 167.955 126.440 168.765 ;
        RECT 126.610 167.775 126.870 168.300 ;
        RECT 127.050 167.955 127.300 168.765 ;
        RECT 133.480 168.595 134.645 169.185 ;
        RECT 134.905 169.235 136.115 170.325 ;
        RECT 134.905 168.695 135.425 169.235 ;
        RECT 127.900 168.425 134.645 168.595 ;
        RECT 135.595 168.525 136.115 169.065 ;
        RECT 127.470 167.775 127.730 168.335 ;
        RECT 127.900 167.970 128.160 168.425 ;
        RECT 128.330 167.775 128.590 168.255 ;
        RECT 128.760 167.970 129.020 168.425 ;
        RECT 129.190 167.775 129.450 168.255 ;
        RECT 129.620 167.970 129.880 168.425 ;
        RECT 130.050 167.775 130.295 168.255 ;
        RECT 130.465 167.970 130.740 168.425 ;
        RECT 130.910 167.775 131.155 168.255 ;
        RECT 131.325 167.970 131.585 168.425 ;
        RECT 131.765 167.775 132.015 168.255 ;
        RECT 132.185 167.970 132.445 168.425 ;
        RECT 132.625 167.775 132.875 168.255 ;
        RECT 133.045 167.970 133.305 168.425 ;
        RECT 133.485 167.775 133.745 168.255 ;
        RECT 133.915 167.970 134.175 168.425 ;
        RECT 134.345 167.775 134.645 168.255 ;
        RECT 134.905 167.775 136.115 168.525 ;
        RECT 23.500 167.605 136.200 167.775 ;
        RECT 23.585 166.855 24.795 167.605 ;
        RECT 24.965 167.105 25.225 167.435 ;
        RECT 25.435 167.125 25.710 167.605 ;
        RECT 23.585 166.315 24.105 166.855 ;
        RECT 24.275 166.145 24.795 166.685 ;
        RECT 23.585 165.055 24.795 166.145 ;
        RECT 24.965 166.195 25.135 167.105 ;
        RECT 25.920 167.035 26.125 167.435 ;
        RECT 26.295 167.205 26.630 167.605 ;
        RECT 26.805 167.060 32.150 167.605 ;
        RECT 25.305 166.365 25.665 166.945 ;
        RECT 25.920 166.865 26.605 167.035 ;
        RECT 25.845 166.195 26.095 166.695 ;
        RECT 24.965 166.025 26.095 166.195 ;
        RECT 24.965 165.255 25.235 166.025 ;
        RECT 26.265 165.835 26.605 166.865 ;
        RECT 28.390 166.230 28.730 167.060 ;
        RECT 32.325 166.835 35.835 167.605 ;
        RECT 36.005 166.855 37.215 167.605 ;
        RECT 37.405 166.875 37.695 167.605 ;
        RECT 25.405 165.055 25.735 165.835 ;
        RECT 25.940 165.660 26.605 165.835 ;
        RECT 25.940 165.255 26.125 165.660 ;
        RECT 30.210 165.490 30.560 166.740 ;
        RECT 32.325 166.315 33.975 166.835 ;
        RECT 34.145 166.145 35.835 166.665 ;
        RECT 36.005 166.315 36.525 166.855 ;
        RECT 36.695 166.145 37.215 166.685 ;
        RECT 37.395 166.365 37.695 166.695 ;
        RECT 37.875 166.675 38.105 167.315 ;
        RECT 38.285 167.055 38.595 167.425 ;
        RECT 38.775 167.235 39.445 167.605 ;
        RECT 38.285 166.855 39.515 167.055 ;
        RECT 37.875 166.365 38.400 166.675 ;
        RECT 38.580 166.365 39.045 166.675 ;
        RECT 39.225 166.185 39.515 166.855 ;
        RECT 26.295 165.055 26.630 165.480 ;
        RECT 26.805 165.055 32.150 165.490 ;
        RECT 32.325 165.055 35.835 166.145 ;
        RECT 36.005 165.055 37.215 166.145 ;
        RECT 37.405 165.945 38.565 166.185 ;
        RECT 37.405 165.235 37.665 165.945 ;
        RECT 37.835 165.055 38.165 165.765 ;
        RECT 38.335 165.235 38.565 165.945 ;
        RECT 38.745 165.965 39.515 166.185 ;
        RECT 38.745 165.235 39.015 165.965 ;
        RECT 39.195 165.055 39.535 165.785 ;
        RECT 39.705 165.235 39.965 167.425 ;
        RECT 40.195 167.065 40.420 167.425 ;
        RECT 40.600 167.235 40.930 167.605 ;
        RECT 41.110 167.065 41.365 167.425 ;
        RECT 41.930 167.235 42.675 167.605 ;
        RECT 40.195 166.875 42.680 167.065 ;
        RECT 40.155 166.365 40.425 166.695 ;
        RECT 40.605 166.365 41.040 166.695 ;
        RECT 41.220 166.365 41.795 166.695 ;
        RECT 41.975 166.365 42.255 166.695 ;
        RECT 42.455 166.185 42.680 166.875 ;
        RECT 40.185 166.005 42.680 166.185 ;
        RECT 42.855 166.005 43.190 167.425 ;
        RECT 44.445 167.045 44.775 167.435 ;
        RECT 44.945 167.215 46.130 167.385 ;
        RECT 46.390 167.135 46.560 167.605 ;
        RECT 44.445 166.865 44.955 167.045 ;
        RECT 44.285 166.405 44.615 166.695 ;
        RECT 44.785 166.235 44.955 166.865 ;
        RECT 45.360 166.955 45.745 167.045 ;
        RECT 46.730 166.955 47.060 167.420 ;
        RECT 45.360 166.785 47.060 166.955 ;
        RECT 47.230 166.785 47.400 167.605 ;
        RECT 47.570 166.785 48.255 167.425 ;
        RECT 49.345 166.880 49.635 167.605 ;
        RECT 49.810 167.130 50.145 167.390 ;
        RECT 50.315 167.205 50.645 167.605 ;
        RECT 50.815 167.205 52.430 167.375 ;
        RECT 45.125 166.405 45.455 166.615 ;
        RECT 45.635 166.365 46.015 166.615 ;
        RECT 46.205 166.585 46.690 166.615 ;
        RECT 46.185 166.415 46.690 166.585 ;
        RECT 40.185 165.235 40.475 166.005 ;
        RECT 41.045 165.595 42.235 165.825 ;
        RECT 41.045 165.235 41.305 165.595 ;
        RECT 41.475 165.055 41.805 165.425 ;
        RECT 41.975 165.235 42.235 165.595 ;
        RECT 42.425 165.055 42.755 165.775 ;
        RECT 42.925 165.235 43.190 166.005 ;
        RECT 44.440 166.065 45.525 166.235 ;
        RECT 44.440 165.225 44.740 166.065 ;
        RECT 44.935 165.055 45.185 165.895 ;
        RECT 45.355 165.815 45.525 166.065 ;
        RECT 45.695 165.985 46.015 166.365 ;
        RECT 46.205 166.405 46.690 166.415 ;
        RECT 46.880 166.405 47.330 166.615 ;
        RECT 47.500 166.405 47.835 166.615 ;
        RECT 46.205 165.985 46.580 166.405 ;
        RECT 47.500 166.235 47.670 166.405 ;
        RECT 46.750 166.065 47.670 166.235 ;
        RECT 46.750 165.815 46.920 166.065 ;
        RECT 45.355 165.645 46.920 165.815 ;
        RECT 45.775 165.225 46.580 165.645 ;
        RECT 47.090 165.055 47.420 165.895 ;
        RECT 48.005 165.815 48.255 166.785 ;
        RECT 47.590 165.225 48.255 165.815 ;
        RECT 49.345 165.055 49.635 166.220 ;
        RECT 49.810 165.775 50.065 167.130 ;
        RECT 50.815 167.035 50.985 167.205 ;
        RECT 50.425 166.865 50.985 167.035 ;
        RECT 51.250 166.925 51.520 167.025 ;
        RECT 51.710 166.925 52.000 167.025 ;
        RECT 50.425 166.695 50.595 166.865 ;
        RECT 51.245 166.755 51.520 166.925 ;
        RECT 51.705 166.755 52.000 166.925 ;
        RECT 50.290 166.365 50.595 166.695 ;
        RECT 50.790 166.585 51.040 166.695 ;
        RECT 50.785 166.415 51.040 166.585 ;
        RECT 50.790 166.365 51.040 166.415 ;
        RECT 51.250 166.365 51.520 166.755 ;
        RECT 51.710 166.365 52.000 166.755 ;
        RECT 52.170 166.365 52.590 167.030 ;
        RECT 52.975 166.885 53.305 167.605 ;
        RECT 53.485 167.105 53.745 167.435 ;
        RECT 53.915 167.245 54.245 167.605 ;
        RECT 54.500 167.225 55.800 167.435 ;
        RECT 53.485 167.095 53.715 167.105 ;
        RECT 52.900 166.585 53.250 166.695 ;
        RECT 52.900 166.415 53.255 166.585 ;
        RECT 52.900 166.365 53.250 166.415 ;
        RECT 50.425 166.195 50.595 166.365 ;
        RECT 50.425 166.025 52.795 166.195 ;
        RECT 53.045 166.075 53.250 166.365 ;
        RECT 49.810 165.265 50.145 165.775 ;
        RECT 50.395 165.055 50.725 165.855 ;
        RECT 50.970 165.645 52.395 165.815 ;
        RECT 50.970 165.225 51.255 165.645 ;
        RECT 51.510 165.055 51.840 165.475 ;
        RECT 52.065 165.395 52.395 165.645 ;
        RECT 52.625 165.565 52.795 166.025 ;
        RECT 53.485 165.905 53.655 167.095 ;
        RECT 54.500 167.075 54.670 167.225 ;
        RECT 53.915 166.950 54.670 167.075 ;
        RECT 53.825 166.905 54.670 166.950 ;
        RECT 53.825 166.785 54.095 166.905 ;
        RECT 53.825 166.210 53.995 166.785 ;
        RECT 54.225 166.345 54.635 166.650 ;
        RECT 54.925 166.615 55.135 167.015 ;
        RECT 54.805 166.405 55.135 166.615 ;
        RECT 55.380 166.615 55.600 167.015 ;
        RECT 56.075 166.840 56.530 167.605 ;
        RECT 56.705 166.970 56.975 167.605 ;
        RECT 57.160 166.915 57.395 167.435 ;
        RECT 57.565 167.110 57.965 167.605 ;
        RECT 58.555 167.275 58.725 167.420 ;
        RECT 58.325 167.080 58.725 167.275 ;
        RECT 55.380 166.405 55.855 166.615 ;
        RECT 56.045 166.415 56.535 166.615 ;
        RECT 53.825 166.175 54.025 166.210 ;
        RECT 55.355 166.175 56.530 166.235 ;
        RECT 53.825 166.065 56.530 166.175 ;
        RECT 53.885 166.005 55.685 166.065 ;
        RECT 55.355 165.975 55.685 166.005 ;
        RECT 53.055 165.395 53.225 165.895 ;
        RECT 52.065 165.225 53.225 165.395 ;
        RECT 53.485 165.225 53.745 165.905 ;
        RECT 53.915 165.055 54.165 165.835 ;
        RECT 54.415 165.805 55.250 165.815 ;
        RECT 55.840 165.805 56.025 165.895 ;
        RECT 54.415 165.605 56.025 165.805 ;
        RECT 54.415 165.225 54.665 165.605 ;
        RECT 55.795 165.565 56.025 165.605 ;
        RECT 56.275 165.445 56.530 166.065 ;
        RECT 57.160 166.110 57.335 166.915 ;
        RECT 58.325 166.745 58.495 167.080 ;
        RECT 59.005 167.035 59.245 167.410 ;
        RECT 59.415 167.100 59.745 167.605 ;
        RECT 59.005 166.885 59.220 167.035 ;
        RECT 57.505 166.385 58.495 166.745 ;
        RECT 58.665 166.555 59.220 166.885 ;
        RECT 57.505 166.365 58.795 166.385 ;
        RECT 57.935 166.215 58.795 166.365 ;
        RECT 54.835 165.055 55.190 165.435 ;
        RECT 56.195 165.225 56.530 165.445 ;
        RECT 56.705 165.055 56.975 166.010 ;
        RECT 57.160 165.325 57.465 166.110 ;
        RECT 57.640 165.735 58.335 166.045 ;
        RECT 57.645 165.055 58.330 165.525 ;
        RECT 58.510 165.270 58.795 166.215 ;
        RECT 58.985 165.905 59.220 166.555 ;
        RECT 59.390 166.585 59.690 166.925 ;
        RECT 59.945 166.795 60.185 167.605 ;
        RECT 60.355 166.795 60.685 167.435 ;
        RECT 60.855 166.795 61.125 167.605 ;
        RECT 61.305 167.060 66.650 167.605 ;
        RECT 66.825 167.060 72.170 167.605 ;
        RECT 73.265 167.105 73.525 167.435 ;
        RECT 73.735 167.125 74.010 167.605 ;
        RECT 59.390 166.415 59.695 166.585 ;
        RECT 59.390 166.075 59.690 166.415 ;
        RECT 59.925 166.365 60.275 166.615 ;
        RECT 60.445 166.195 60.615 166.795 ;
        RECT 60.785 166.365 61.135 166.615 ;
        RECT 62.890 166.230 63.230 167.060 ;
        RECT 59.935 166.025 60.615 166.195 ;
        RECT 58.985 165.675 59.665 165.905 ;
        RECT 58.995 165.055 59.325 165.505 ;
        RECT 59.495 165.245 59.665 165.675 ;
        RECT 59.935 165.240 60.265 166.025 ;
        RECT 60.795 165.055 61.125 166.195 ;
        RECT 64.710 165.490 65.060 166.740 ;
        RECT 68.410 166.230 68.750 167.060 ;
        RECT 70.230 165.490 70.580 166.740 ;
        RECT 73.265 166.195 73.435 167.105 ;
        RECT 74.220 167.035 74.425 167.435 ;
        RECT 74.595 167.205 74.930 167.605 ;
        RECT 73.605 166.365 73.965 166.945 ;
        RECT 74.220 166.865 74.905 167.035 ;
        RECT 75.105 166.880 75.395 167.605 ;
        RECT 75.575 167.010 75.825 167.435 ;
        RECT 75.995 167.180 76.325 167.605 ;
        RECT 76.495 167.185 77.585 167.435 ;
        RECT 77.775 167.185 78.865 167.435 ;
        RECT 76.495 167.010 76.665 167.185 ;
        RECT 74.145 166.195 74.395 166.695 ;
        RECT 73.265 166.025 74.395 166.195 ;
        RECT 61.305 165.055 66.650 165.490 ;
        RECT 66.825 165.055 72.170 165.490 ;
        RECT 73.265 165.255 73.535 166.025 ;
        RECT 74.565 165.835 74.905 166.865 ;
        RECT 75.575 166.840 76.665 167.010 ;
        RECT 76.835 166.845 78.525 167.015 ;
        RECT 78.695 167.010 78.865 167.185 ;
        RECT 79.035 167.180 79.365 167.605 ;
        RECT 79.535 167.010 79.855 167.435 ;
        RECT 75.630 166.585 76.260 166.615 ;
        RECT 76.550 166.585 77.180 166.615 ;
        RECT 75.625 166.415 76.260 166.585 ;
        RECT 76.545 166.415 77.180 166.585 ;
        RECT 73.705 165.055 74.035 165.835 ;
        RECT 74.240 165.660 74.905 165.835 ;
        RECT 74.240 165.255 74.425 165.660 ;
        RECT 74.595 165.055 74.930 165.480 ;
        RECT 75.105 165.055 75.395 166.220 ;
        RECT 77.350 166.205 77.640 166.845 ;
        RECT 78.695 166.840 79.855 167.010 ;
        RECT 81.085 167.105 81.345 167.435 ;
        RECT 81.555 167.125 81.830 167.605 ;
        RECT 77.925 166.415 78.580 166.615 ;
        RECT 78.870 166.585 79.980 166.615 ;
        RECT 78.845 166.415 79.980 166.585 ;
        RECT 75.575 166.035 77.640 166.205 ;
        RECT 75.575 165.225 75.825 166.035 ;
        RECT 75.995 165.395 76.245 165.865 ;
        RECT 76.415 165.565 76.745 166.035 ;
        RECT 76.915 165.395 77.085 165.865 ;
        RECT 77.255 165.565 77.640 166.035 ;
        RECT 77.855 166.035 79.785 166.205 ;
        RECT 77.855 165.395 78.105 166.035 ;
        RECT 75.995 165.225 78.105 165.395 ;
        RECT 78.275 165.055 78.445 165.865 ;
        RECT 78.615 165.225 78.945 166.035 ;
        RECT 79.115 165.055 79.285 165.865 ;
        RECT 79.455 165.225 79.785 166.035 ;
        RECT 81.085 166.195 81.255 167.105 ;
        RECT 82.040 167.035 82.245 167.435 ;
        RECT 82.415 167.205 82.750 167.605 ;
        RECT 83.015 167.055 83.185 167.435 ;
        RECT 83.365 167.225 83.695 167.605 ;
        RECT 81.425 166.365 81.785 166.945 ;
        RECT 82.040 166.865 82.725 167.035 ;
        RECT 83.015 166.885 83.680 167.055 ;
        RECT 83.875 166.930 84.135 167.435 ;
        RECT 81.965 166.195 82.215 166.695 ;
        RECT 81.085 166.025 82.215 166.195 ;
        RECT 81.085 165.255 81.355 166.025 ;
        RECT 82.385 165.835 82.725 166.865 ;
        RECT 82.945 166.335 83.285 166.705 ;
        RECT 83.510 166.630 83.680 166.885 ;
        RECT 83.510 166.300 83.785 166.630 ;
        RECT 83.510 166.155 83.680 166.300 ;
        RECT 81.525 165.055 81.855 165.835 ;
        RECT 82.060 165.660 82.725 165.835 ;
        RECT 83.005 165.985 83.680 166.155 ;
        RECT 83.955 166.130 84.135 166.930 ;
        RECT 84.855 167.055 85.025 167.435 ;
        RECT 85.205 167.225 85.535 167.605 ;
        RECT 84.855 166.885 85.520 167.055 ;
        RECT 85.715 166.930 85.975 167.435 ;
        RECT 84.785 166.335 85.125 166.705 ;
        RECT 85.350 166.630 85.520 166.885 ;
        RECT 85.350 166.300 85.625 166.630 ;
        RECT 85.350 166.155 85.520 166.300 ;
        RECT 82.060 165.255 82.245 165.660 ;
        RECT 82.415 165.055 82.750 165.480 ;
        RECT 83.005 165.225 83.185 165.985 ;
        RECT 83.365 165.055 83.695 165.815 ;
        RECT 83.865 165.225 84.135 166.130 ;
        RECT 84.845 165.985 85.520 166.155 ;
        RECT 85.795 166.130 85.975 166.930 ;
        RECT 86.235 167.055 86.405 167.435 ;
        RECT 86.585 167.225 86.915 167.605 ;
        RECT 86.235 166.885 86.900 167.055 ;
        RECT 87.095 166.930 87.355 167.435 ;
        RECT 86.165 166.335 86.505 166.705 ;
        RECT 86.730 166.630 86.900 166.885 ;
        RECT 86.730 166.300 87.005 166.630 ;
        RECT 86.730 166.155 86.900 166.300 ;
        RECT 84.845 165.225 85.025 165.985 ;
        RECT 85.205 165.055 85.535 165.815 ;
        RECT 85.705 165.225 85.975 166.130 ;
        RECT 86.225 165.985 86.900 166.155 ;
        RECT 87.175 166.130 87.355 166.930 ;
        RECT 87.615 167.055 87.785 167.435 ;
        RECT 87.965 167.225 88.295 167.605 ;
        RECT 87.615 166.885 88.280 167.055 ;
        RECT 88.475 166.930 88.735 167.435 ;
        RECT 87.545 166.335 87.875 166.705 ;
        RECT 88.110 166.630 88.280 166.885 ;
        RECT 88.110 166.300 88.395 166.630 ;
        RECT 88.110 166.155 88.280 166.300 ;
        RECT 86.225 165.225 86.405 165.985 ;
        RECT 86.585 165.055 86.915 165.815 ;
        RECT 87.085 165.225 87.355 166.130 ;
        RECT 87.615 165.985 88.280 166.155 ;
        RECT 88.565 166.130 88.735 166.930 ;
        RECT 88.910 166.765 89.170 167.605 ;
        RECT 89.345 166.860 89.600 167.435 ;
        RECT 89.770 167.225 90.100 167.605 ;
        RECT 90.315 167.055 90.485 167.435 ;
        RECT 89.770 166.885 90.485 167.055 ;
        RECT 87.615 165.225 87.785 165.985 ;
        RECT 87.965 165.055 88.295 165.815 ;
        RECT 88.465 165.225 88.735 166.130 ;
        RECT 88.910 165.055 89.170 166.205 ;
        RECT 89.345 166.130 89.515 166.860 ;
        RECT 89.770 166.695 89.940 166.885 ;
        RECT 89.685 166.365 89.940 166.695 ;
        RECT 89.770 166.155 89.940 166.365 ;
        RECT 90.220 166.335 90.575 166.705 ;
        RECT 89.345 165.225 89.600 166.130 ;
        RECT 89.770 165.985 90.485 166.155 ;
        RECT 89.770 165.055 90.100 165.815 ;
        RECT 90.315 165.225 90.485 165.985 ;
        RECT 90.745 165.225 91.495 167.435 ;
        RECT 91.665 167.105 91.925 167.435 ;
        RECT 92.095 167.245 92.425 167.605 ;
        RECT 92.680 167.225 93.980 167.435 ;
        RECT 91.665 165.905 91.835 167.105 ;
        RECT 92.680 167.075 92.850 167.225 ;
        RECT 92.095 166.950 92.850 167.075 ;
        RECT 92.005 166.905 92.850 166.950 ;
        RECT 92.005 166.785 92.275 166.905 ;
        RECT 92.005 166.210 92.175 166.785 ;
        RECT 92.405 166.345 92.815 166.650 ;
        RECT 93.105 166.615 93.315 167.015 ;
        RECT 92.985 166.405 93.315 166.615 ;
        RECT 93.560 166.615 93.780 167.015 ;
        RECT 94.255 166.840 94.710 167.605 ;
        RECT 94.945 166.785 95.155 167.605 ;
        RECT 95.325 166.805 95.655 167.435 ;
        RECT 93.560 166.405 94.035 166.615 ;
        RECT 94.225 166.415 94.715 166.615 ;
        RECT 92.005 166.175 92.205 166.210 ;
        RECT 93.535 166.175 94.710 166.235 ;
        RECT 95.325 166.205 95.575 166.805 ;
        RECT 95.825 166.785 96.055 167.605 ;
        RECT 96.265 167.105 96.525 167.435 ;
        RECT 96.695 167.245 97.025 167.605 ;
        RECT 97.280 167.225 98.580 167.435 ;
        RECT 96.265 167.095 96.495 167.105 ;
        RECT 95.745 166.365 96.075 166.615 ;
        RECT 92.005 166.065 94.710 166.175 ;
        RECT 92.065 166.005 93.865 166.065 ;
        RECT 93.535 165.975 93.865 166.005 ;
        RECT 91.665 165.225 91.925 165.905 ;
        RECT 92.095 165.055 92.345 165.835 ;
        RECT 92.595 165.805 93.430 165.815 ;
        RECT 94.020 165.805 94.205 165.895 ;
        RECT 92.595 165.605 94.205 165.805 ;
        RECT 92.595 165.225 92.845 165.605 ;
        RECT 93.975 165.565 94.205 165.605 ;
        RECT 94.455 165.445 94.710 166.065 ;
        RECT 93.015 165.055 93.370 165.435 ;
        RECT 94.375 165.225 94.710 165.445 ;
        RECT 94.945 165.055 95.155 166.195 ;
        RECT 95.325 165.225 95.655 166.205 ;
        RECT 95.825 165.055 96.055 166.195 ;
        RECT 96.265 165.905 96.435 167.095 ;
        RECT 97.280 167.075 97.450 167.225 ;
        RECT 96.695 166.950 97.450 167.075 ;
        RECT 96.605 166.905 97.450 166.950 ;
        RECT 96.605 166.785 96.875 166.905 ;
        RECT 96.605 166.210 96.775 166.785 ;
        RECT 97.005 166.345 97.415 166.650 ;
        RECT 97.705 166.615 97.915 167.015 ;
        RECT 97.585 166.405 97.915 166.615 ;
        RECT 98.160 166.615 98.380 167.015 ;
        RECT 98.855 166.840 99.310 167.605 ;
        RECT 99.485 166.930 99.745 167.435 ;
        RECT 99.925 167.225 100.255 167.605 ;
        RECT 100.435 167.055 100.605 167.435 ;
        RECT 98.160 166.405 98.635 166.615 ;
        RECT 98.825 166.415 99.315 166.615 ;
        RECT 96.605 166.175 96.805 166.210 ;
        RECT 98.135 166.175 99.310 166.235 ;
        RECT 96.605 166.065 99.310 166.175 ;
        RECT 96.665 166.005 98.465 166.065 ;
        RECT 98.135 165.975 98.465 166.005 ;
        RECT 96.265 165.225 96.525 165.905 ;
        RECT 96.695 165.055 96.945 165.835 ;
        RECT 97.195 165.805 98.030 165.815 ;
        RECT 98.620 165.805 98.805 165.895 ;
        RECT 97.195 165.605 98.805 165.805 ;
        RECT 97.195 165.225 97.445 165.605 ;
        RECT 98.575 165.565 98.805 165.605 ;
        RECT 99.055 165.445 99.310 166.065 ;
        RECT 97.615 165.055 97.970 165.435 ;
        RECT 98.975 165.225 99.310 165.445 ;
        RECT 99.485 166.130 99.655 166.930 ;
        RECT 99.940 166.885 100.605 167.055 ;
        RECT 99.940 166.630 100.110 166.885 ;
        RECT 100.865 166.880 101.155 167.605 ;
        RECT 101.325 166.945 101.600 167.605 ;
        RECT 101.770 166.975 102.020 167.435 ;
        RECT 102.195 167.110 102.525 167.605 ;
        RECT 101.770 166.765 101.940 166.975 ;
        RECT 102.705 166.940 102.935 167.385 ;
        RECT 99.825 166.300 100.110 166.630 ;
        RECT 100.345 166.335 100.675 166.705 ;
        RECT 99.940 166.155 100.110 166.300 ;
        RECT 101.325 166.245 101.940 166.765 ;
        RECT 102.110 166.265 102.340 166.695 ;
        RECT 102.525 166.445 102.935 166.940 ;
        RECT 103.105 167.120 103.895 167.385 ;
        RECT 103.105 166.265 103.360 167.120 ;
        RECT 104.170 167.055 104.500 167.435 ;
        RECT 104.670 167.225 105.855 167.395 ;
        RECT 106.115 167.135 106.285 167.605 ;
        RECT 103.530 166.445 103.915 166.925 ;
        RECT 104.170 166.885 104.715 167.055 ;
        RECT 104.085 166.365 104.345 166.715 ;
        RECT 99.485 165.225 99.755 166.130 ;
        RECT 99.940 165.985 100.605 166.155 ;
        RECT 99.925 165.055 100.255 165.815 ;
        RECT 100.435 165.225 100.605 165.985 ;
        RECT 100.865 165.055 101.155 166.220 ;
        RECT 101.325 165.055 101.585 166.065 ;
        RECT 101.755 165.895 101.925 166.245 ;
        RECT 102.110 166.095 103.900 166.265 ;
        RECT 104.545 166.245 104.715 166.885 ;
        RECT 105.085 166.955 105.470 167.045 ;
        RECT 106.455 166.955 106.785 167.420 ;
        RECT 105.085 166.785 106.785 166.955 ;
        RECT 106.955 166.785 107.125 167.605 ;
        RECT 107.295 166.955 107.625 167.425 ;
        RECT 107.795 167.125 107.965 167.605 ;
        RECT 107.295 166.785 108.055 166.955 ;
        RECT 108.225 166.805 108.920 167.435 ;
        RECT 109.125 166.805 109.435 167.605 ;
        RECT 109.605 167.095 109.910 167.605 ;
        RECT 104.885 166.415 105.230 166.615 ;
        RECT 105.400 166.415 105.790 166.615 ;
        RECT 104.545 166.195 105.330 166.245 ;
        RECT 101.755 165.225 102.030 165.895 ;
        RECT 102.230 165.055 102.445 165.900 ;
        RECT 102.670 165.800 102.920 166.095 ;
        RECT 103.145 165.735 103.475 165.925 ;
        RECT 102.630 165.225 103.105 165.565 ;
        RECT 103.285 165.560 103.475 165.735 ;
        RECT 103.645 165.730 103.900 166.095 ;
        RECT 104.250 166.020 105.330 166.195 ;
        RECT 103.285 165.055 103.915 165.560 ;
        RECT 104.250 165.225 104.580 166.020 ;
        RECT 104.750 165.055 104.990 165.840 ;
        RECT 105.160 165.815 105.330 166.020 ;
        RECT 105.500 165.985 105.790 166.415 ;
        RECT 105.980 166.405 106.465 166.615 ;
        RECT 106.635 166.405 107.075 166.615 ;
        RECT 107.245 166.405 107.575 166.615 ;
        RECT 105.980 165.985 106.285 166.405 ;
        RECT 107.245 166.235 107.415 166.405 ;
        RECT 106.455 166.065 107.415 166.235 ;
        RECT 106.455 165.815 106.625 166.065 ;
        RECT 105.160 165.645 106.625 165.815 ;
        RECT 105.550 165.225 106.305 165.645 ;
        RECT 106.795 165.055 107.125 165.895 ;
        RECT 107.745 165.815 108.055 166.785 ;
        RECT 108.245 166.365 108.580 166.615 ;
        RECT 108.750 166.245 108.920 166.805 ;
        RECT 109.090 166.365 109.425 166.635 ;
        RECT 109.605 166.365 109.920 166.925 ;
        RECT 110.090 166.615 110.340 167.425 ;
        RECT 110.510 167.080 110.770 167.605 ;
        RECT 110.950 166.615 111.200 167.425 ;
        RECT 111.370 167.045 111.630 167.605 ;
        RECT 111.800 166.955 112.060 167.410 ;
        RECT 112.230 167.125 112.490 167.605 ;
        RECT 112.660 166.955 112.920 167.410 ;
        RECT 113.090 167.125 113.350 167.605 ;
        RECT 113.520 166.955 113.780 167.410 ;
        RECT 113.950 167.125 114.195 167.605 ;
        RECT 114.365 166.955 114.640 167.410 ;
        RECT 114.810 167.125 115.055 167.605 ;
        RECT 115.225 166.955 115.485 167.410 ;
        RECT 115.665 167.125 115.915 167.605 ;
        RECT 116.085 166.955 116.345 167.410 ;
        RECT 116.525 167.125 116.775 167.605 ;
        RECT 116.945 166.955 117.205 167.410 ;
        RECT 117.385 167.125 117.645 167.605 ;
        RECT 117.815 166.955 118.075 167.410 ;
        RECT 118.245 167.125 118.545 167.605 ;
        RECT 118.865 167.145 119.110 167.605 ;
        RECT 111.800 166.785 118.545 166.955 ;
        RECT 110.090 166.365 117.210 166.615 ;
        RECT 108.745 166.205 108.920 166.245 ;
        RECT 107.295 165.645 108.055 165.815 ;
        RECT 107.295 165.225 107.545 165.645 ;
        RECT 107.715 165.055 108.055 165.475 ;
        RECT 108.225 165.055 108.485 166.195 ;
        RECT 108.655 165.225 108.985 166.205 ;
        RECT 109.155 165.055 109.435 166.195 ;
        RECT 109.615 165.055 109.910 165.865 ;
        RECT 110.090 165.225 110.335 166.365 ;
        RECT 110.510 165.055 110.770 165.865 ;
        RECT 110.950 165.230 111.200 166.365 ;
        RECT 117.380 166.195 118.545 166.785 ;
        RECT 118.805 166.365 119.120 166.975 ;
        RECT 119.290 166.615 119.540 167.425 ;
        RECT 119.710 167.080 119.970 167.605 ;
        RECT 120.140 166.955 120.400 167.410 ;
        RECT 120.570 167.125 120.830 167.605 ;
        RECT 121.000 166.955 121.260 167.410 ;
        RECT 121.430 167.125 121.690 167.605 ;
        RECT 121.860 166.955 122.120 167.410 ;
        RECT 122.290 167.125 122.550 167.605 ;
        RECT 122.720 166.955 122.980 167.410 ;
        RECT 123.150 167.125 123.450 167.605 ;
        RECT 120.140 166.785 123.450 166.955 ;
        RECT 119.290 166.365 122.310 166.615 ;
        RECT 111.800 165.970 118.545 166.195 ;
        RECT 111.800 165.955 117.205 165.970 ;
        RECT 111.370 165.060 111.630 165.855 ;
        RECT 111.800 165.230 112.060 165.955 ;
        RECT 112.230 165.060 112.490 165.785 ;
        RECT 112.660 165.230 112.920 165.955 ;
        RECT 113.090 165.060 113.350 165.785 ;
        RECT 113.520 165.230 113.780 165.955 ;
        RECT 113.950 165.060 114.210 165.785 ;
        RECT 114.380 165.230 114.640 165.955 ;
        RECT 114.810 165.060 115.055 165.785 ;
        RECT 115.225 165.230 115.485 165.955 ;
        RECT 115.670 165.060 115.915 165.785 ;
        RECT 116.085 165.230 116.345 165.955 ;
        RECT 116.530 165.060 116.775 165.785 ;
        RECT 116.945 165.230 117.205 165.955 ;
        RECT 117.390 165.060 117.645 165.785 ;
        RECT 117.815 165.230 118.105 165.970 ;
        RECT 111.370 165.055 117.645 165.060 ;
        RECT 118.275 165.055 118.545 165.800 ;
        RECT 118.815 165.055 119.110 166.165 ;
        RECT 119.290 165.230 119.540 166.365 ;
        RECT 122.480 166.195 123.450 166.785 ;
        RECT 119.710 165.055 119.970 166.165 ;
        RECT 120.140 165.955 123.450 166.195 ;
        RECT 123.865 166.930 124.135 167.275 ;
        RECT 124.325 167.205 124.705 167.605 ;
        RECT 124.875 167.035 125.045 167.385 ;
        RECT 125.215 167.205 125.545 167.605 ;
        RECT 125.745 167.035 125.915 167.385 ;
        RECT 126.115 167.105 126.445 167.605 ;
        RECT 123.865 166.195 124.035 166.930 ;
        RECT 124.305 166.865 125.915 167.035 ;
        RECT 124.305 166.695 124.475 166.865 ;
        RECT 124.205 166.365 124.475 166.695 ;
        RECT 124.645 166.365 125.050 166.695 ;
        RECT 124.305 166.195 124.475 166.365 ;
        RECT 125.220 166.245 125.930 166.695 ;
        RECT 126.100 166.365 126.450 166.935 ;
        RECT 126.625 166.880 126.915 167.605 ;
        RECT 127.085 166.865 127.345 167.605 ;
        RECT 127.595 166.785 127.785 167.255 ;
        RECT 128.035 167.105 128.285 167.605 ;
        RECT 128.615 167.035 128.785 167.385 ;
        RECT 128.985 167.205 129.315 167.605 ;
        RECT 129.485 167.035 129.655 167.385 ;
        RECT 129.875 167.205 130.255 167.605 ;
        RECT 127.615 166.695 127.785 166.785 ;
        RECT 128.455 166.865 130.265 167.035 ;
        RECT 120.140 165.230 120.400 165.955 ;
        RECT 120.570 165.055 120.830 165.785 ;
        RECT 121.000 165.230 121.260 165.955 ;
        RECT 121.430 165.055 121.690 165.785 ;
        RECT 121.860 165.230 122.120 165.955 ;
        RECT 122.290 165.055 122.550 165.785 ;
        RECT 122.720 165.230 122.980 165.955 ;
        RECT 123.150 165.055 123.445 165.785 ;
        RECT 123.865 165.225 124.135 166.195 ;
        RECT 124.305 166.025 125.030 166.195 ;
        RECT 125.220 166.075 125.935 166.245 ;
        RECT 124.860 165.905 125.030 166.025 ;
        RECT 126.130 165.905 126.450 166.195 ;
        RECT 124.345 165.055 124.625 165.855 ;
        RECT 124.860 165.735 126.450 165.905 ;
        RECT 124.795 165.275 126.450 165.565 ;
        RECT 126.625 165.055 126.915 166.220 ;
        RECT 127.105 165.735 127.445 166.695 ;
        RECT 127.615 166.365 128.215 166.695 ;
        RECT 127.615 165.625 127.785 166.365 ;
        RECT 128.455 166.115 128.625 166.865 ;
        RECT 127.085 165.055 127.365 165.555 ;
        RECT 127.595 165.235 127.785 165.625 ;
        RECT 128.035 165.945 128.625 166.115 ;
        RECT 128.795 166.070 128.965 166.695 ;
        RECT 129.195 166.240 129.525 166.695 ;
        RECT 128.035 165.240 128.365 165.945 ;
        RECT 128.795 165.315 129.155 166.070 ;
        RECT 129.335 165.905 129.525 166.240 ;
        RECT 129.755 166.245 129.925 166.695 ;
        RECT 130.095 166.615 130.265 166.865 ;
        RECT 130.435 166.965 130.685 167.435 ;
        RECT 130.855 167.135 131.025 167.605 ;
        RECT 131.195 166.965 131.525 167.435 ;
        RECT 131.695 167.135 131.865 167.605 ;
        RECT 130.435 166.785 131.965 166.965 ;
        RECT 132.155 166.955 132.485 167.420 ;
        RECT 132.655 167.135 132.825 167.605 ;
        RECT 133.000 167.205 133.330 167.435 ;
        RECT 133.535 167.265 133.705 167.435 ;
        RECT 133.080 166.955 133.250 167.205 ;
        RECT 133.535 167.095 133.755 167.265 ;
        RECT 133.535 167.045 133.705 167.095 ;
        RECT 132.155 166.785 133.250 166.955 ;
        RECT 133.465 166.865 133.705 167.045 ;
        RECT 134.050 167.035 134.240 167.195 ;
        RECT 133.930 166.865 134.240 167.035 ;
        RECT 134.460 166.865 134.735 167.605 ;
        RECT 130.095 166.445 131.555 166.615 ;
        RECT 129.755 166.075 130.190 166.245 ;
        RECT 131.725 166.235 131.965 166.785 ;
        RECT 132.145 166.405 132.625 166.615 ;
        RECT 132.795 166.405 133.295 166.615 ;
        RECT 133.465 166.235 133.635 166.865 ;
        RECT 133.930 166.695 134.100 166.865 ;
        RECT 134.905 166.855 136.115 167.605 ;
        RECT 130.395 166.065 131.965 166.235 ;
        RECT 129.335 165.315 129.635 165.905 ;
        RECT 129.920 165.055 130.170 165.895 ;
        RECT 130.395 165.225 130.645 166.065 ;
        RECT 130.815 165.055 131.065 165.895 ;
        RECT 131.235 165.225 131.485 166.065 ;
        RECT 131.655 165.055 131.905 165.895 ;
        RECT 132.175 165.055 132.550 166.155 ;
        RECT 133.025 166.065 133.635 166.235 ;
        RECT 133.805 166.155 134.100 166.695 ;
        RECT 134.285 166.345 134.735 166.695 ;
        RECT 133.025 165.225 133.350 166.065 ;
        RECT 133.805 165.985 134.295 166.155 ;
        RECT 133.520 165.055 133.850 165.815 ;
        RECT 134.020 165.480 134.295 165.985 ;
        RECT 134.465 165.245 134.735 166.345 ;
        RECT 134.905 166.145 135.425 166.685 ;
        RECT 135.595 166.315 136.115 166.855 ;
        RECT 134.905 165.055 136.115 166.145 ;
        RECT 23.500 164.885 136.200 165.055 ;
        RECT 23.585 163.795 24.795 164.885 ;
        RECT 24.965 164.450 30.310 164.885 ;
        RECT 30.485 164.450 35.830 164.885 ;
        RECT 23.585 163.085 24.105 163.625 ;
        RECT 24.275 163.255 24.795 163.795 ;
        RECT 23.585 162.335 24.795 163.085 ;
        RECT 26.550 162.880 26.890 163.710 ;
        RECT 28.370 163.200 28.720 164.450 ;
        RECT 32.070 162.880 32.410 163.710 ;
        RECT 33.890 163.200 34.240 164.450 ;
        RECT 36.465 163.720 36.755 164.885 ;
        RECT 36.925 163.795 38.135 164.885 ;
        RECT 38.395 164.265 38.565 164.695 ;
        RECT 38.735 164.435 39.065 164.885 ;
        RECT 38.395 164.035 39.075 164.265 ;
        RECT 36.925 163.085 37.445 163.625 ;
        RECT 37.615 163.255 38.135 163.795 ;
        RECT 38.370 163.185 38.670 163.865 ;
        RECT 24.965 162.335 30.310 162.880 ;
        RECT 30.485 162.335 35.830 162.880 ;
        RECT 36.465 162.335 36.755 163.060 ;
        RECT 36.925 162.335 38.135 163.085 ;
        RECT 38.365 163.015 38.670 163.185 ;
        RECT 38.840 163.385 39.075 164.035 ;
        RECT 39.265 163.725 39.550 164.670 ;
        RECT 39.730 164.415 40.415 164.885 ;
        RECT 39.725 163.895 40.420 164.205 ;
        RECT 40.595 163.830 40.900 164.615 ;
        RECT 41.085 163.930 41.355 164.885 ;
        RECT 41.615 164.265 41.785 164.695 ;
        RECT 41.955 164.435 42.285 164.885 ;
        RECT 41.615 164.035 42.290 164.265 ;
        RECT 39.265 163.575 40.125 163.725 ;
        RECT 39.265 163.555 40.555 163.575 ;
        RECT 38.840 163.055 39.395 163.385 ;
        RECT 39.565 163.195 40.555 163.555 ;
        RECT 38.840 162.905 39.055 163.055 ;
        RECT 38.315 162.335 38.645 162.840 ;
        RECT 38.815 162.530 39.055 162.905 ;
        RECT 39.565 162.860 39.735 163.195 ;
        RECT 40.725 163.025 40.900 163.830 ;
        RECT 39.335 162.665 39.735 162.860 ;
        RECT 39.335 162.520 39.505 162.665 ;
        RECT 40.095 162.335 40.495 162.830 ;
        RECT 40.665 162.505 40.900 163.025 ;
        RECT 41.585 163.015 41.885 163.865 ;
        RECT 42.055 163.385 42.290 164.035 ;
        RECT 42.460 163.725 42.745 164.670 ;
        RECT 42.925 164.415 43.610 164.885 ;
        RECT 42.920 163.895 43.615 164.205 ;
        RECT 43.790 163.830 44.095 164.615 ;
        RECT 42.460 163.575 43.320 163.725 ;
        RECT 43.885 163.695 44.095 163.830 ;
        RECT 44.285 163.795 46.875 164.885 ;
        RECT 42.460 163.555 43.745 163.575 ;
        RECT 42.055 163.055 42.590 163.385 ;
        RECT 42.760 163.195 43.745 163.555 ;
        RECT 41.085 162.335 41.355 162.970 ;
        RECT 42.055 162.905 42.275 163.055 ;
        RECT 41.530 162.335 41.865 162.840 ;
        RECT 42.035 162.530 42.275 162.905 ;
        RECT 42.760 162.860 42.930 163.195 ;
        RECT 43.920 163.025 44.095 163.695 ;
        RECT 42.555 162.665 42.930 162.860 ;
        RECT 42.555 162.520 42.725 162.665 ;
        RECT 43.290 162.335 43.685 162.830 ;
        RECT 43.855 162.505 44.095 163.025 ;
        RECT 44.285 163.105 45.495 163.625 ;
        RECT 45.665 163.275 46.875 163.795 ;
        RECT 47.545 163.935 47.835 164.705 ;
        RECT 48.405 164.345 48.665 164.705 ;
        RECT 48.835 164.515 49.165 164.885 ;
        RECT 49.335 164.345 49.595 164.705 ;
        RECT 48.405 164.115 49.595 164.345 ;
        RECT 49.785 164.165 50.115 164.885 ;
        RECT 50.285 163.935 50.550 164.705 ;
        RECT 47.545 163.755 50.040 163.935 ;
        RECT 47.515 163.245 47.785 163.575 ;
        RECT 47.965 163.245 48.400 163.575 ;
        RECT 48.580 163.245 49.155 163.575 ;
        RECT 49.335 163.245 49.615 163.575 ;
        RECT 44.285 162.335 46.875 163.105 ;
        RECT 49.815 163.065 50.040 163.755 ;
        RECT 47.555 162.875 50.040 163.065 ;
        RECT 47.555 162.515 47.780 162.875 ;
        RECT 47.960 162.335 48.290 162.705 ;
        RECT 48.470 162.515 48.725 162.875 ;
        RECT 49.290 162.335 50.035 162.705 ;
        RECT 50.215 162.515 50.550 163.935 ;
        RECT 50.725 163.795 53.315 164.885 ;
        RECT 50.725 163.105 51.935 163.625 ;
        RECT 52.105 163.275 53.315 163.795 ;
        RECT 53.955 163.745 54.285 164.885 ;
        RECT 54.815 163.915 55.145 164.700 ;
        RECT 55.820 164.085 56.070 164.885 ;
        RECT 56.240 164.255 56.570 164.715 ;
        RECT 56.740 164.425 56.955 164.885 ;
        RECT 56.240 164.085 57.410 164.255 ;
        RECT 54.465 163.745 55.145 163.915 ;
        RECT 55.330 163.915 55.610 164.075 ;
        RECT 55.330 163.745 56.665 163.915 ;
        RECT 53.945 163.325 54.295 163.575 ;
        RECT 54.465 163.145 54.635 163.745 ;
        RECT 56.495 163.575 56.665 163.745 ;
        RECT 54.805 163.325 55.155 163.575 ;
        RECT 55.330 163.325 55.680 163.565 ;
        RECT 55.850 163.325 56.325 163.565 ;
        RECT 56.495 163.325 56.870 163.575 ;
        RECT 56.495 163.155 56.665 163.325 ;
        RECT 50.725 162.335 53.315 163.105 ;
        RECT 53.955 162.335 54.225 163.145 ;
        RECT 54.395 162.505 54.725 163.145 ;
        RECT 54.895 162.335 55.135 163.145 ;
        RECT 55.330 162.985 56.665 163.155 ;
        RECT 55.330 162.775 55.600 162.985 ;
        RECT 57.040 162.795 57.410 164.085 ;
        RECT 58.175 163.915 58.345 164.715 ;
        RECT 59.105 164.255 59.355 164.715 ;
        RECT 59.555 164.505 60.225 164.885 ;
        RECT 60.415 164.255 60.665 164.715 ;
        RECT 60.840 164.425 61.085 164.885 ;
        RECT 59.105 164.085 60.665 164.255 ;
        RECT 61.255 164.035 61.595 164.675 ;
        RECT 58.175 163.745 61.115 163.915 ;
        RECT 60.945 163.575 61.115 163.745 ;
        RECT 58.145 163.245 58.330 163.575 ;
        RECT 58.585 163.245 59.060 163.575 ;
        RECT 59.370 163.245 59.715 163.575 ;
        RECT 55.820 162.335 56.150 162.795 ;
        RECT 56.660 162.505 57.410 162.795 ;
        RECT 58.175 162.905 59.355 163.075 ;
        RECT 59.525 163.015 59.715 163.245 ;
        RECT 59.975 163.000 60.170 163.575 ;
        RECT 60.440 163.245 60.775 163.575 ;
        RECT 60.945 163.245 61.255 163.575 ;
        RECT 60.945 163.075 61.115 163.245 ;
        RECT 58.175 162.505 58.345 162.905 ;
        RECT 58.585 162.335 58.915 162.735 ;
        RECT 59.185 162.675 59.355 162.905 ;
        RECT 60.420 162.905 61.115 163.075 ;
        RECT 61.425 162.920 61.595 164.035 ;
        RECT 62.225 163.720 62.515 164.885 ;
        RECT 62.690 163.735 62.950 164.885 ;
        RECT 63.125 163.810 63.380 164.715 ;
        RECT 63.550 164.125 63.880 164.885 ;
        RECT 64.095 163.955 64.265 164.715 ;
        RECT 64.525 164.450 69.870 164.885 ;
        RECT 60.420 162.675 60.590 162.905 ;
        RECT 59.185 162.505 60.590 162.675 ;
        RECT 60.760 162.335 61.090 162.715 ;
        RECT 61.285 162.505 61.595 162.920 ;
        RECT 62.225 162.335 62.515 163.060 ;
        RECT 62.690 162.335 62.950 163.175 ;
        RECT 63.125 163.080 63.295 163.810 ;
        RECT 63.550 163.785 64.265 163.955 ;
        RECT 63.550 163.575 63.720 163.785 ;
        RECT 63.465 163.245 63.720 163.575 ;
        RECT 63.125 162.505 63.380 163.080 ;
        RECT 63.550 163.055 63.720 163.245 ;
        RECT 64.000 163.235 64.355 163.605 ;
        RECT 63.550 162.885 64.265 163.055 ;
        RECT 63.550 162.335 63.880 162.715 ;
        RECT 64.095 162.505 64.265 162.885 ;
        RECT 66.110 162.880 66.450 163.710 ;
        RECT 67.930 163.200 68.280 164.450 ;
        RECT 70.045 163.795 71.255 164.885 ;
        RECT 70.045 163.085 70.565 163.625 ;
        RECT 70.735 163.255 71.255 163.795 ;
        RECT 64.525 162.335 69.870 162.880 ;
        RECT 70.045 162.335 71.255 163.085 ;
        RECT 71.435 162.515 71.695 164.705 ;
        RECT 71.865 164.155 72.205 164.885 ;
        RECT 72.385 163.975 72.655 164.705 ;
        RECT 71.885 163.755 72.655 163.975 ;
        RECT 72.835 163.995 73.065 164.705 ;
        RECT 73.235 164.175 73.565 164.885 ;
        RECT 73.735 163.995 73.995 164.705 ;
        RECT 72.835 163.755 73.995 163.995 ;
        RECT 74.195 163.935 74.470 164.705 ;
        RECT 74.640 164.275 74.970 164.705 ;
        RECT 75.140 164.445 75.335 164.885 ;
        RECT 75.515 164.275 75.845 164.705 ;
        RECT 74.640 164.105 75.845 164.275 ;
        RECT 71.885 163.085 72.175 163.755 ;
        RECT 74.195 163.745 74.780 163.935 ;
        RECT 74.950 163.775 75.845 164.105 ;
        RECT 77.035 163.955 77.205 164.715 ;
        RECT 77.385 164.125 77.715 164.885 ;
        RECT 77.035 163.785 77.700 163.955 ;
        RECT 77.885 163.810 78.155 164.715 ;
        RECT 72.355 163.265 72.820 163.575 ;
        RECT 73.000 163.265 73.525 163.575 ;
        RECT 71.885 162.885 73.115 163.085 ;
        RECT 71.955 162.335 72.625 162.705 ;
        RECT 72.805 162.515 73.115 162.885 ;
        RECT 73.295 162.625 73.525 163.265 ;
        RECT 73.705 163.245 74.005 163.575 ;
        RECT 73.705 162.335 73.995 163.065 ;
        RECT 74.195 162.925 74.435 163.575 ;
        RECT 74.605 163.075 74.780 163.745 ;
        RECT 77.530 163.640 77.700 163.785 ;
        RECT 74.950 163.245 75.365 163.575 ;
        RECT 75.545 163.245 75.840 163.575 ;
        RECT 74.605 162.895 74.935 163.075 ;
        RECT 74.210 162.335 74.540 162.725 ;
        RECT 74.710 162.515 74.935 162.895 ;
        RECT 75.135 162.625 75.365 163.245 ;
        RECT 76.965 163.235 77.295 163.605 ;
        RECT 77.530 163.310 77.815 163.640 ;
        RECT 75.545 162.335 75.845 163.065 ;
        RECT 77.530 163.055 77.700 163.310 ;
        RECT 77.035 162.885 77.700 163.055 ;
        RECT 77.985 163.010 78.155 163.810 ;
        RECT 78.385 163.745 78.595 164.885 ;
        RECT 78.765 163.735 79.095 164.715 ;
        RECT 79.265 163.745 79.495 164.885 ;
        RECT 79.795 163.875 79.965 164.715 ;
        RECT 80.135 164.545 81.305 164.715 ;
        RECT 80.135 164.045 80.465 164.545 ;
        RECT 80.975 164.505 81.305 164.545 ;
        RECT 81.495 164.465 81.850 164.885 ;
        RECT 80.635 164.285 80.865 164.375 ;
        RECT 82.020 164.285 82.270 164.715 ;
        RECT 80.635 164.045 82.270 164.285 ;
        RECT 82.440 164.125 82.770 164.885 ;
        RECT 82.940 164.045 83.195 164.715 ;
        RECT 77.035 162.505 77.205 162.885 ;
        RECT 77.385 162.335 77.715 162.715 ;
        RECT 77.895 162.505 78.155 163.010 ;
        RECT 78.385 162.335 78.595 163.155 ;
        RECT 78.765 163.135 79.015 163.735 ;
        RECT 79.795 163.705 82.855 163.875 ;
        RECT 79.185 163.325 79.515 163.575 ;
        RECT 79.710 163.325 80.060 163.535 ;
        RECT 80.230 163.325 80.675 163.525 ;
        RECT 80.845 163.325 81.320 163.525 ;
        RECT 78.765 162.505 79.095 163.135 ;
        RECT 79.265 162.335 79.495 163.155 ;
        RECT 79.795 162.985 80.860 163.155 ;
        RECT 79.795 162.505 79.965 162.985 ;
        RECT 80.135 162.335 80.465 162.815 ;
        RECT 80.690 162.755 80.860 162.985 ;
        RECT 81.040 162.925 81.320 163.325 ;
        RECT 81.590 163.325 81.920 163.525 ;
        RECT 82.090 163.325 82.455 163.525 ;
        RECT 81.590 162.925 81.875 163.325 ;
        RECT 82.685 163.155 82.855 163.705 ;
        RECT 82.055 162.985 82.855 163.155 ;
        RECT 82.055 162.755 82.225 162.985 ;
        RECT 83.025 162.915 83.195 164.045 ;
        RECT 83.855 164.275 84.185 164.705 ;
        RECT 84.365 164.445 84.560 164.885 ;
        RECT 84.730 164.275 85.060 164.705 ;
        RECT 83.855 164.105 85.060 164.275 ;
        RECT 83.855 163.775 84.750 164.105 ;
        RECT 85.230 163.935 85.505 164.705 ;
        RECT 84.920 163.745 85.505 163.935 ;
        RECT 83.860 163.245 84.155 163.575 ;
        RECT 84.335 163.245 84.750 163.575 ;
        RECT 83.010 162.835 83.195 162.915 ;
        RECT 80.690 162.505 82.225 162.755 ;
        RECT 82.395 162.335 82.725 162.815 ;
        RECT 82.940 162.505 83.195 162.835 ;
        RECT 83.855 162.335 84.155 163.065 ;
        RECT 84.335 162.625 84.565 163.245 ;
        RECT 84.920 163.075 85.095 163.745 ;
        RECT 84.765 162.895 85.095 163.075 ;
        RECT 85.265 162.925 85.505 163.575 ;
        RECT 84.765 162.515 84.990 162.895 ;
        RECT 85.160 162.335 85.490 162.725 ;
        RECT 85.685 162.505 86.435 164.715 ;
        RECT 86.695 163.955 86.865 164.715 ;
        RECT 87.045 164.125 87.375 164.885 ;
        RECT 86.695 163.785 87.360 163.955 ;
        RECT 87.545 163.810 87.815 164.715 ;
        RECT 87.190 163.640 87.360 163.785 ;
        RECT 86.625 163.235 86.955 163.605 ;
        RECT 87.190 163.310 87.475 163.640 ;
        RECT 87.190 163.055 87.360 163.310 ;
        RECT 86.695 162.885 87.360 163.055 ;
        RECT 87.645 163.010 87.815 163.810 ;
        RECT 87.985 163.720 88.275 164.885 ;
        RECT 89.860 164.085 90.110 164.885 ;
        RECT 90.280 164.255 90.610 164.715 ;
        RECT 90.780 164.425 90.995 164.885 ;
        RECT 92.625 164.545 93.765 164.715 ;
        RECT 90.280 164.085 91.450 164.255 ;
        RECT 92.625 164.085 92.925 164.545 ;
        RECT 89.370 163.915 89.650 164.075 ;
        RECT 89.370 163.745 90.705 163.915 ;
        RECT 90.535 163.575 90.705 163.745 ;
        RECT 89.370 163.325 89.720 163.565 ;
        RECT 89.890 163.325 90.365 163.565 ;
        RECT 90.535 163.325 90.910 163.575 ;
        RECT 90.535 163.155 90.705 163.325 ;
        RECT 86.695 162.505 86.865 162.885 ;
        RECT 87.045 162.335 87.375 162.715 ;
        RECT 87.555 162.505 87.815 163.010 ;
        RECT 87.985 162.335 88.275 163.060 ;
        RECT 89.370 162.985 90.705 163.155 ;
        RECT 89.370 162.775 89.640 162.985 ;
        RECT 91.080 162.795 91.450 164.085 ;
        RECT 93.095 163.915 93.425 164.375 ;
        RECT 92.665 163.695 93.425 163.915 ;
        RECT 93.595 163.915 93.765 164.545 ;
        RECT 93.935 164.085 94.265 164.885 ;
        RECT 94.435 163.915 94.710 164.715 ;
        RECT 94.940 164.015 95.225 164.885 ;
        RECT 95.395 164.255 95.655 164.715 ;
        RECT 95.830 164.425 96.085 164.885 ;
        RECT 96.255 164.255 96.515 164.715 ;
        RECT 95.395 164.085 96.515 164.255 ;
        RECT 96.685 164.085 96.995 164.885 ;
        RECT 93.595 163.705 94.710 163.915 ;
        RECT 95.395 163.835 95.655 164.085 ;
        RECT 97.165 163.915 97.475 164.715 ;
        RECT 92.665 163.185 92.880 163.695 ;
        RECT 94.900 163.665 95.655 163.835 ;
        RECT 96.445 163.745 97.475 163.915 ;
        RECT 97.650 163.885 97.905 164.885 ;
        RECT 93.050 163.325 93.820 163.525 ;
        RECT 93.990 163.325 94.710 163.525 ;
        RECT 92.645 163.155 92.880 163.185 ;
        RECT 94.900 163.155 95.305 163.665 ;
        RECT 96.445 163.495 96.615 163.745 ;
        RECT 95.475 163.325 96.615 163.495 ;
        RECT 92.645 163.015 94.265 163.155 ;
        RECT 92.665 162.985 94.265 163.015 ;
        RECT 93.095 162.975 94.265 162.985 ;
        RECT 89.860 162.335 90.190 162.795 ;
        RECT 90.700 162.505 91.450 162.795 ;
        RECT 92.635 162.335 92.925 162.805 ;
        RECT 93.095 162.505 93.425 162.975 ;
        RECT 93.595 162.335 93.765 162.805 ;
        RECT 93.935 162.505 94.265 162.975 ;
        RECT 94.435 162.335 94.710 163.155 ;
        RECT 94.900 162.985 96.550 163.155 ;
        RECT 96.785 163.005 97.135 163.575 ;
        RECT 94.945 162.335 95.225 162.815 ;
        RECT 95.395 162.595 95.655 162.985 ;
        RECT 95.830 162.335 96.085 162.815 ;
        RECT 96.255 162.595 96.550 162.985 ;
        RECT 97.305 162.835 97.475 163.745 ;
        RECT 96.730 162.335 97.005 162.815 ;
        RECT 97.175 162.505 97.475 162.835 ;
        RECT 97.665 162.335 97.905 163.135 ;
        RECT 98.090 162.505 98.335 164.715 ;
        RECT 98.505 164.435 99.355 164.885 ;
        RECT 99.525 164.255 99.785 164.715 ;
        RECT 98.665 164.035 99.785 164.255 ;
        RECT 98.665 163.580 98.835 164.035 ;
        RECT 98.505 163.090 98.835 163.580 ;
        RECT 99.005 163.260 99.415 163.865 ;
        RECT 99.965 163.650 100.170 164.235 ;
        RECT 100.355 163.900 100.680 164.885 ;
        RECT 100.885 164.295 101.125 164.685 ;
        RECT 101.295 164.475 101.645 164.885 ;
        RECT 100.885 164.095 101.635 164.295 ;
        RECT 99.585 163.525 100.170 163.650 ;
        RECT 99.585 163.355 100.175 163.525 ;
        RECT 99.585 163.275 100.170 163.355 ;
        RECT 100.425 163.245 100.685 163.700 ;
        RECT 98.505 162.885 99.355 163.090 ;
        RECT 98.505 162.335 98.835 162.715 ;
        RECT 99.025 162.505 99.355 162.885 ;
        RECT 99.525 162.885 100.680 163.075 ;
        RECT 99.525 162.715 99.735 162.885 ;
        RECT 100.405 162.745 100.680 162.885 ;
        RECT 99.905 162.335 100.235 162.715 ;
        RECT 100.885 162.575 101.115 163.915 ;
        RECT 101.295 163.415 101.635 164.095 ;
        RECT 101.815 163.595 102.145 164.705 ;
        RECT 102.315 164.235 102.495 164.705 ;
        RECT 102.665 164.405 102.995 164.885 ;
        RECT 103.170 164.235 103.340 164.705 ;
        RECT 102.315 164.035 103.340 164.235 ;
        RECT 101.295 162.515 101.525 163.415 ;
        RECT 101.815 163.295 102.360 163.595 ;
        RECT 101.725 162.335 101.970 163.115 ;
        RECT 102.140 163.065 102.360 163.295 ;
        RECT 102.530 163.245 102.955 163.865 ;
        RECT 103.150 163.245 103.410 163.865 ;
        RECT 103.605 163.745 103.890 164.885 ;
        RECT 103.620 163.065 103.880 163.575 ;
        RECT 102.140 162.875 103.880 163.065 ;
        RECT 102.140 162.515 102.570 162.875 ;
        RECT 103.150 162.335 103.880 162.705 ;
        RECT 104.080 162.515 104.360 164.705 ;
        RECT 104.635 164.140 104.905 164.885 ;
        RECT 105.535 164.880 111.810 164.885 ;
        RECT 105.075 163.970 105.365 164.710 ;
        RECT 105.535 164.155 105.790 164.880 ;
        RECT 105.975 163.985 106.235 164.710 ;
        RECT 106.405 164.155 106.650 164.880 ;
        RECT 106.835 163.985 107.095 164.710 ;
        RECT 107.265 164.155 107.510 164.880 ;
        RECT 107.695 163.985 107.955 164.710 ;
        RECT 108.125 164.155 108.370 164.880 ;
        RECT 108.540 163.985 108.800 164.710 ;
        RECT 108.970 164.155 109.230 164.880 ;
        RECT 109.400 163.985 109.660 164.710 ;
        RECT 109.830 164.155 110.090 164.880 ;
        RECT 110.260 163.985 110.520 164.710 ;
        RECT 110.690 164.155 110.950 164.880 ;
        RECT 111.120 163.985 111.380 164.710 ;
        RECT 111.550 164.085 111.810 164.880 ;
        RECT 105.975 163.970 111.380 163.985 ;
        RECT 104.635 163.745 111.380 163.970 ;
        RECT 104.635 163.155 105.800 163.745 ;
        RECT 111.980 163.575 112.230 164.710 ;
        RECT 112.410 164.075 112.670 164.885 ;
        RECT 112.845 163.575 113.090 164.715 ;
        RECT 113.270 164.075 113.565 164.885 ;
        RECT 113.745 163.720 114.035 164.885 ;
        RECT 114.215 164.075 114.510 164.885 ;
        RECT 114.690 163.575 114.935 164.715 ;
        RECT 115.110 164.075 115.370 164.885 ;
        RECT 115.970 164.880 122.245 164.885 ;
        RECT 115.550 163.575 115.800 164.710 ;
        RECT 115.970 164.085 116.230 164.880 ;
        RECT 116.400 163.985 116.660 164.710 ;
        RECT 116.830 164.155 117.090 164.880 ;
        RECT 117.260 163.985 117.520 164.710 ;
        RECT 117.690 164.155 117.950 164.880 ;
        RECT 118.120 163.985 118.380 164.710 ;
        RECT 118.550 164.155 118.810 164.880 ;
        RECT 118.980 163.985 119.240 164.710 ;
        RECT 119.410 164.155 119.655 164.880 ;
        RECT 119.825 163.985 120.085 164.710 ;
        RECT 120.270 164.155 120.515 164.880 ;
        RECT 120.685 163.985 120.945 164.710 ;
        RECT 121.130 164.155 121.375 164.880 ;
        RECT 121.545 163.985 121.805 164.710 ;
        RECT 121.990 164.155 122.245 164.880 ;
        RECT 116.400 163.970 121.805 163.985 ;
        RECT 122.415 163.970 122.705 164.710 ;
        RECT 122.875 164.140 123.145 164.885 ;
        RECT 123.495 164.140 123.765 164.885 ;
        RECT 124.395 164.880 130.670 164.885 ;
        RECT 123.935 163.970 124.225 164.710 ;
        RECT 124.395 164.155 124.650 164.880 ;
        RECT 124.835 163.985 125.095 164.710 ;
        RECT 125.265 164.155 125.510 164.880 ;
        RECT 125.695 163.985 125.955 164.710 ;
        RECT 126.125 164.155 126.370 164.880 ;
        RECT 126.555 163.985 126.815 164.710 ;
        RECT 126.985 164.155 127.230 164.880 ;
        RECT 127.400 163.985 127.660 164.710 ;
        RECT 127.830 164.155 128.090 164.880 ;
        RECT 128.260 163.985 128.520 164.710 ;
        RECT 128.690 164.155 128.950 164.880 ;
        RECT 129.120 163.985 129.380 164.710 ;
        RECT 129.550 164.155 129.810 164.880 ;
        RECT 129.980 163.985 130.240 164.710 ;
        RECT 130.410 164.085 130.670 164.880 ;
        RECT 124.835 163.970 130.240 163.985 ;
        RECT 116.400 163.745 123.145 163.970 ;
        RECT 105.970 163.325 113.090 163.575 ;
        RECT 104.635 162.985 111.380 163.155 ;
        RECT 104.635 162.335 104.935 162.815 ;
        RECT 105.105 162.530 105.365 162.985 ;
        RECT 105.535 162.335 105.795 162.815 ;
        RECT 105.975 162.530 106.235 162.985 ;
        RECT 106.405 162.335 106.655 162.815 ;
        RECT 106.835 162.530 107.095 162.985 ;
        RECT 107.265 162.335 107.515 162.815 ;
        RECT 107.695 162.530 107.955 162.985 ;
        RECT 108.125 162.335 108.370 162.815 ;
        RECT 108.540 162.530 108.815 162.985 ;
        RECT 108.985 162.335 109.230 162.815 ;
        RECT 109.400 162.530 109.660 162.985 ;
        RECT 109.830 162.335 110.090 162.815 ;
        RECT 110.260 162.530 110.520 162.985 ;
        RECT 110.690 162.335 110.950 162.815 ;
        RECT 111.120 162.530 111.380 162.985 ;
        RECT 111.550 162.335 111.810 162.895 ;
        RECT 111.980 162.515 112.230 163.325 ;
        RECT 112.410 162.335 112.670 162.860 ;
        RECT 112.840 162.515 113.090 163.325 ;
        RECT 113.260 163.015 113.575 163.575 ;
        RECT 113.270 162.335 113.575 162.845 ;
        RECT 113.745 162.335 114.035 163.060 ;
        RECT 114.205 163.015 114.520 163.575 ;
        RECT 114.690 163.325 121.810 163.575 ;
        RECT 114.205 162.335 114.510 162.845 ;
        RECT 114.690 162.515 114.940 163.325 ;
        RECT 115.110 162.335 115.370 162.860 ;
        RECT 115.550 162.515 115.800 163.325 ;
        RECT 121.980 163.155 123.145 163.745 ;
        RECT 116.400 162.985 123.145 163.155 ;
        RECT 123.495 163.745 130.240 163.970 ;
        RECT 123.495 163.155 124.660 163.745 ;
        RECT 130.840 163.575 131.090 164.710 ;
        RECT 131.270 164.075 131.530 164.885 ;
        RECT 131.705 163.575 131.950 164.715 ;
        RECT 132.130 164.075 132.425 164.885 ;
        RECT 133.155 163.955 133.325 164.715 ;
        RECT 133.540 164.125 133.870 164.885 ;
        RECT 133.155 163.785 133.870 163.955 ;
        RECT 134.040 163.810 134.295 164.715 ;
        RECT 124.830 163.325 131.950 163.575 ;
        RECT 123.495 162.985 130.240 163.155 ;
        RECT 115.970 162.335 116.230 162.895 ;
        RECT 116.400 162.530 116.660 162.985 ;
        RECT 116.830 162.335 117.090 162.815 ;
        RECT 117.260 162.530 117.520 162.985 ;
        RECT 117.690 162.335 117.950 162.815 ;
        RECT 118.120 162.530 118.380 162.985 ;
        RECT 118.550 162.335 118.795 162.815 ;
        RECT 118.965 162.530 119.240 162.985 ;
        RECT 119.410 162.335 119.655 162.815 ;
        RECT 119.825 162.530 120.085 162.985 ;
        RECT 120.265 162.335 120.515 162.815 ;
        RECT 120.685 162.530 120.945 162.985 ;
        RECT 121.125 162.335 121.375 162.815 ;
        RECT 121.545 162.530 121.805 162.985 ;
        RECT 121.985 162.335 122.245 162.815 ;
        RECT 122.415 162.530 122.675 162.985 ;
        RECT 122.845 162.335 123.145 162.815 ;
        RECT 123.495 162.335 123.795 162.815 ;
        RECT 123.965 162.530 124.225 162.985 ;
        RECT 124.395 162.335 124.655 162.815 ;
        RECT 124.835 162.530 125.095 162.985 ;
        RECT 125.265 162.335 125.515 162.815 ;
        RECT 125.695 162.530 125.955 162.985 ;
        RECT 126.125 162.335 126.375 162.815 ;
        RECT 126.555 162.530 126.815 162.985 ;
        RECT 126.985 162.335 127.230 162.815 ;
        RECT 127.400 162.530 127.675 162.985 ;
        RECT 127.845 162.335 128.090 162.815 ;
        RECT 128.260 162.530 128.520 162.985 ;
        RECT 128.690 162.335 128.950 162.815 ;
        RECT 129.120 162.530 129.380 162.985 ;
        RECT 129.550 162.335 129.810 162.815 ;
        RECT 129.980 162.530 130.240 162.985 ;
        RECT 130.410 162.335 130.670 162.895 ;
        RECT 130.840 162.515 131.090 163.325 ;
        RECT 131.270 162.335 131.530 162.860 ;
        RECT 131.700 162.515 131.950 163.325 ;
        RECT 132.120 163.015 132.435 163.575 ;
        RECT 133.065 163.235 133.420 163.605 ;
        RECT 133.700 163.575 133.870 163.785 ;
        RECT 133.700 163.245 133.955 163.575 ;
        RECT 133.700 163.055 133.870 163.245 ;
        RECT 134.125 163.080 134.295 163.810 ;
        RECT 134.470 163.735 134.730 164.885 ;
        RECT 134.905 163.795 136.115 164.885 ;
        RECT 134.905 163.255 135.425 163.795 ;
        RECT 133.155 162.885 133.870 163.055 ;
        RECT 132.130 162.335 132.435 162.845 ;
        RECT 133.155 162.505 133.325 162.885 ;
        RECT 133.540 162.335 133.870 162.715 ;
        RECT 134.040 162.505 134.295 163.080 ;
        RECT 134.470 162.335 134.730 163.175 ;
        RECT 135.595 163.085 136.115 163.625 ;
        RECT 134.905 162.335 136.115 163.085 ;
        RECT 23.500 162.165 136.200 162.335 ;
        RECT 23.585 161.415 24.795 162.165 ;
        RECT 24.965 161.620 30.310 162.165 ;
        RECT 30.485 161.620 35.830 162.165 ;
        RECT 23.585 160.875 24.105 161.415 ;
        RECT 24.275 160.705 24.795 161.245 ;
        RECT 26.550 160.790 26.890 161.620 ;
        RECT 23.585 159.615 24.795 160.705 ;
        RECT 28.370 160.050 28.720 161.300 ;
        RECT 32.070 160.790 32.410 161.620 ;
        RECT 36.005 161.395 37.675 162.165 ;
        RECT 38.310 161.765 38.645 162.165 ;
        RECT 38.815 161.595 39.020 161.995 ;
        RECT 39.230 161.685 39.505 162.165 ;
        RECT 39.715 161.665 39.975 161.995 ;
        RECT 38.335 161.425 39.020 161.595 ;
        RECT 33.890 160.050 34.240 161.300 ;
        RECT 36.005 160.875 36.755 161.395 ;
        RECT 36.925 160.705 37.675 161.225 ;
        RECT 24.965 159.615 30.310 160.050 ;
        RECT 30.485 159.615 35.830 160.050 ;
        RECT 36.005 159.615 37.675 160.705 ;
        RECT 38.335 160.395 38.675 161.425 ;
        RECT 38.845 160.755 39.095 161.255 ;
        RECT 39.275 160.925 39.635 161.505 ;
        RECT 39.805 160.755 39.975 161.665 ;
        RECT 40.145 161.395 42.735 162.165 ;
        RECT 42.905 161.705 43.465 161.995 ;
        RECT 43.635 161.705 43.885 162.165 ;
        RECT 40.145 160.875 41.355 161.395 ;
        RECT 38.845 160.585 39.975 160.755 ;
        RECT 41.525 160.705 42.735 161.225 ;
        RECT 38.335 160.220 39.000 160.395 ;
        RECT 38.310 159.615 38.645 160.040 ;
        RECT 38.815 159.815 39.000 160.220 ;
        RECT 39.205 159.615 39.535 160.395 ;
        RECT 39.705 159.815 39.975 160.585 ;
        RECT 40.145 159.615 42.735 160.705 ;
        RECT 42.905 160.335 43.155 161.705 ;
        RECT 44.505 161.535 44.835 161.895 ;
        RECT 45.210 161.765 45.545 162.165 ;
        RECT 45.715 161.595 45.920 161.995 ;
        RECT 46.130 161.685 46.405 162.165 ;
        RECT 46.615 161.665 46.875 161.995 ;
        RECT 43.445 161.345 44.835 161.535 ;
        RECT 45.235 161.425 45.920 161.595 ;
        RECT 43.445 161.255 43.615 161.345 ;
        RECT 43.325 160.925 43.615 161.255 ;
        RECT 43.785 160.925 44.125 161.175 ;
        RECT 44.345 160.925 45.020 161.175 ;
        RECT 43.445 160.675 43.615 160.925 ;
        RECT 43.445 160.505 44.385 160.675 ;
        RECT 44.755 160.565 45.020 160.925 ;
        RECT 42.905 159.785 43.365 160.335 ;
        RECT 43.555 159.615 43.885 160.335 ;
        RECT 44.085 159.955 44.385 160.505 ;
        RECT 45.235 160.395 45.575 161.425 ;
        RECT 45.745 160.755 45.995 161.255 ;
        RECT 46.175 160.925 46.535 161.505 ;
        RECT 46.705 160.755 46.875 161.665 ;
        RECT 47.045 161.395 48.715 162.165 ;
        RECT 49.345 161.440 49.635 162.165 ;
        RECT 49.805 161.620 55.150 162.165 ;
        RECT 47.045 160.875 47.795 161.395 ;
        RECT 45.745 160.585 46.875 160.755 ;
        RECT 47.965 160.705 48.715 161.225 ;
        RECT 51.390 160.790 51.730 161.620 ;
        RECT 55.785 161.365 56.480 161.995 ;
        RECT 56.685 161.365 56.995 162.165 ;
        RECT 57.625 161.580 57.935 161.995 ;
        RECT 58.130 161.785 58.460 162.165 ;
        RECT 58.630 161.825 60.035 161.995 ;
        RECT 58.630 161.595 58.800 161.825 ;
        RECT 44.555 159.615 44.835 160.285 ;
        RECT 45.235 160.220 45.900 160.395 ;
        RECT 45.210 159.615 45.545 160.040 ;
        RECT 45.715 159.815 45.900 160.220 ;
        RECT 46.105 159.615 46.435 160.395 ;
        RECT 46.605 159.815 46.875 160.585 ;
        RECT 47.045 159.615 48.715 160.705 ;
        RECT 49.345 159.615 49.635 160.780 ;
        RECT 53.210 160.050 53.560 161.300 ;
        RECT 55.805 160.925 56.140 161.175 ;
        RECT 56.310 160.805 56.480 161.365 ;
        RECT 56.650 160.925 56.985 161.195 ;
        RECT 56.305 160.765 56.480 160.805 ;
        RECT 49.805 159.615 55.150 160.050 ;
        RECT 55.785 159.615 56.045 160.755 ;
        RECT 56.215 159.785 56.545 160.765 ;
        RECT 56.715 159.615 56.995 160.755 ;
        RECT 57.625 160.465 57.795 161.580 ;
        RECT 58.105 161.425 58.800 161.595 ;
        RECT 59.865 161.595 60.035 161.825 ;
        RECT 60.305 161.765 60.635 162.165 ;
        RECT 60.875 161.595 61.045 161.995 ;
        RECT 58.105 161.255 58.275 161.425 ;
        RECT 57.965 160.925 58.275 161.255 ;
        RECT 58.445 160.925 58.780 161.255 ;
        RECT 59.050 160.925 59.245 161.500 ;
        RECT 59.505 161.255 59.695 161.485 ;
        RECT 59.865 161.425 61.045 161.595 ;
        RECT 61.340 161.425 61.955 161.995 ;
        RECT 62.125 161.655 62.340 162.165 ;
        RECT 62.570 161.655 62.850 161.985 ;
        RECT 63.030 161.655 63.270 162.165 ;
        RECT 63.630 161.775 63.960 162.165 ;
        RECT 59.505 160.925 59.850 161.255 ;
        RECT 60.160 160.925 60.635 161.255 ;
        RECT 60.890 160.925 61.075 161.255 ;
        RECT 58.105 160.755 58.275 160.925 ;
        RECT 58.105 160.585 61.045 160.755 ;
        RECT 57.625 159.825 57.965 160.465 ;
        RECT 58.555 160.245 60.115 160.415 ;
        RECT 58.135 159.615 58.380 160.075 ;
        RECT 58.555 159.785 58.805 160.245 ;
        RECT 58.995 159.615 59.665 159.995 ;
        RECT 59.865 159.785 60.115 160.245 ;
        RECT 60.875 159.785 61.045 160.585 ;
        RECT 61.340 160.405 61.655 161.425 ;
        RECT 61.825 160.755 61.995 161.255 ;
        RECT 62.245 160.925 62.510 161.485 ;
        RECT 62.680 160.755 62.850 161.655 ;
        RECT 64.130 161.605 64.355 161.985 ;
        RECT 63.020 160.925 63.375 161.485 ;
        RECT 63.615 160.925 63.855 161.575 ;
        RECT 64.025 161.425 64.355 161.605 ;
        RECT 64.025 160.755 64.200 161.425 ;
        RECT 64.555 161.255 64.785 161.875 ;
        RECT 64.965 161.435 65.265 162.165 ;
        RECT 65.445 161.365 65.755 162.165 ;
        RECT 65.960 161.365 66.655 161.995 ;
        RECT 66.825 161.620 72.170 162.165 ;
        RECT 72.355 161.665 72.685 162.165 ;
        RECT 65.960 161.315 66.135 161.365 ;
        RECT 64.370 160.925 64.785 161.255 ;
        RECT 64.965 160.925 65.260 161.255 ;
        RECT 65.455 160.925 65.790 161.195 ;
        RECT 65.960 160.765 66.130 161.315 ;
        RECT 66.300 160.925 66.635 161.175 ;
        RECT 68.410 160.790 68.750 161.620 ;
        RECT 72.885 161.595 73.055 161.945 ;
        RECT 73.255 161.765 73.585 162.165 ;
        RECT 73.755 161.595 73.925 161.945 ;
        RECT 74.095 161.765 74.475 162.165 ;
        RECT 61.825 160.585 63.250 160.755 ;
        RECT 61.340 159.785 61.875 160.405 ;
        RECT 62.045 159.615 62.375 160.415 ;
        RECT 62.860 160.410 63.250 160.585 ;
        RECT 63.615 160.565 64.200 160.755 ;
        RECT 63.615 159.795 63.890 160.565 ;
        RECT 64.370 160.395 65.265 160.725 ;
        RECT 64.060 160.225 65.265 160.395 ;
        RECT 64.060 159.795 64.390 160.225 ;
        RECT 64.560 159.615 64.755 160.055 ;
        RECT 64.935 159.795 65.265 160.225 ;
        RECT 65.445 159.615 65.725 160.755 ;
        RECT 65.895 159.785 66.225 160.765 ;
        RECT 66.395 159.615 66.655 160.755 ;
        RECT 70.230 160.050 70.580 161.300 ;
        RECT 72.350 160.925 72.700 161.495 ;
        RECT 72.885 161.425 74.495 161.595 ;
        RECT 74.665 161.490 74.935 161.835 ;
        RECT 74.325 161.255 74.495 161.425 ;
        RECT 72.350 160.465 72.670 160.755 ;
        RECT 72.870 160.635 73.580 161.255 ;
        RECT 73.750 160.925 74.155 161.255 ;
        RECT 74.325 160.925 74.595 161.255 ;
        RECT 74.325 160.755 74.495 160.925 ;
        RECT 74.765 160.755 74.935 161.490 ;
        RECT 75.105 161.440 75.395 162.165 ;
        RECT 75.565 161.785 76.455 161.955 ;
        RECT 75.565 161.230 76.115 161.615 ;
        RECT 76.285 161.060 76.455 161.785 ;
        RECT 75.565 160.990 76.455 161.060 ;
        RECT 76.625 161.460 76.845 161.945 ;
        RECT 77.015 161.625 77.265 162.165 ;
        RECT 77.435 161.515 77.695 161.995 ;
        RECT 77.865 161.785 78.755 161.955 ;
        RECT 76.625 161.035 76.955 161.460 ;
        RECT 75.565 160.965 76.460 160.990 ;
        RECT 75.565 160.950 76.470 160.965 ;
        RECT 75.565 160.935 76.475 160.950 ;
        RECT 75.565 160.930 76.485 160.935 ;
        RECT 75.565 160.920 76.490 160.930 ;
        RECT 75.565 160.910 76.495 160.920 ;
        RECT 75.565 160.905 76.505 160.910 ;
        RECT 75.565 160.895 76.515 160.905 ;
        RECT 75.565 160.890 76.525 160.895 ;
        RECT 73.770 160.585 74.495 160.755 ;
        RECT 73.770 160.465 73.940 160.585 ;
        RECT 72.350 160.295 73.940 160.465 ;
        RECT 66.825 159.615 72.170 160.050 ;
        RECT 72.350 159.835 74.005 160.125 ;
        RECT 74.175 159.615 74.455 160.415 ;
        RECT 74.665 159.785 74.935 160.755 ;
        RECT 75.105 159.615 75.395 160.780 ;
        RECT 75.565 160.440 75.825 160.890 ;
        RECT 76.190 160.885 76.525 160.890 ;
        RECT 76.190 160.880 76.540 160.885 ;
        RECT 76.190 160.870 76.555 160.880 ;
        RECT 76.190 160.865 76.580 160.870 ;
        RECT 77.125 160.865 77.355 161.260 ;
        RECT 76.190 160.860 77.355 160.865 ;
        RECT 76.220 160.825 77.355 160.860 ;
        RECT 76.255 160.800 77.355 160.825 ;
        RECT 76.285 160.770 77.355 160.800 ;
        RECT 76.305 160.740 77.355 160.770 ;
        RECT 76.325 160.710 77.355 160.740 ;
        RECT 76.395 160.700 77.355 160.710 ;
        RECT 76.420 160.690 77.355 160.700 ;
        RECT 76.440 160.675 77.355 160.690 ;
        RECT 76.460 160.660 77.355 160.675 ;
        RECT 76.465 160.650 77.250 160.660 ;
        RECT 76.480 160.615 77.250 160.650 ;
        RECT 75.995 160.295 76.325 160.540 ;
        RECT 76.495 160.365 77.250 160.615 ;
        RECT 77.525 160.485 77.695 161.515 ;
        RECT 77.865 161.230 78.415 161.615 ;
        RECT 78.585 161.060 78.755 161.785 ;
        RECT 75.995 160.270 76.180 160.295 ;
        RECT 75.565 160.170 76.180 160.270 ;
        RECT 75.565 159.615 76.170 160.170 ;
        RECT 76.345 159.785 76.825 160.125 ;
        RECT 76.995 159.615 77.250 160.160 ;
        RECT 77.420 159.785 77.695 160.485 ;
        RECT 77.865 160.990 78.755 161.060 ;
        RECT 78.925 161.460 79.145 161.945 ;
        RECT 79.315 161.625 79.565 162.165 ;
        RECT 79.735 161.515 79.995 161.995 ;
        RECT 78.925 161.035 79.255 161.460 ;
        RECT 77.865 160.965 78.760 160.990 ;
        RECT 77.865 160.950 78.770 160.965 ;
        RECT 77.865 160.935 78.775 160.950 ;
        RECT 77.865 160.930 78.785 160.935 ;
        RECT 77.865 160.920 78.790 160.930 ;
        RECT 77.865 160.910 78.795 160.920 ;
        RECT 77.865 160.905 78.805 160.910 ;
        RECT 77.865 160.895 78.815 160.905 ;
        RECT 77.865 160.890 78.825 160.895 ;
        RECT 77.865 160.440 78.125 160.890 ;
        RECT 78.490 160.885 78.825 160.890 ;
        RECT 78.490 160.880 78.840 160.885 ;
        RECT 78.490 160.870 78.855 160.880 ;
        RECT 78.490 160.865 78.880 160.870 ;
        RECT 79.425 160.865 79.655 161.260 ;
        RECT 78.490 160.860 79.655 160.865 ;
        RECT 78.520 160.825 79.655 160.860 ;
        RECT 78.555 160.800 79.655 160.825 ;
        RECT 78.585 160.770 79.655 160.800 ;
        RECT 78.605 160.740 79.655 160.770 ;
        RECT 78.625 160.710 79.655 160.740 ;
        RECT 78.695 160.700 79.655 160.710 ;
        RECT 78.720 160.690 79.655 160.700 ;
        RECT 78.740 160.675 79.655 160.690 ;
        RECT 78.760 160.660 79.655 160.675 ;
        RECT 78.765 160.650 79.550 160.660 ;
        RECT 78.780 160.615 79.550 160.650 ;
        RECT 78.295 160.295 78.625 160.540 ;
        RECT 78.795 160.365 79.550 160.615 ;
        RECT 79.825 160.485 79.995 161.515 ;
        RECT 80.165 161.415 81.375 162.165 ;
        RECT 81.555 161.435 81.855 162.165 ;
        RECT 80.165 160.875 80.685 161.415 ;
        RECT 82.035 161.255 82.265 161.875 ;
        RECT 82.465 161.605 82.690 161.985 ;
        RECT 82.860 161.775 83.190 162.165 ;
        RECT 82.465 161.425 82.795 161.605 ;
        RECT 80.855 160.705 81.375 161.245 ;
        RECT 81.560 160.925 81.855 161.255 ;
        RECT 82.035 160.925 82.450 161.255 ;
        RECT 82.620 160.755 82.795 161.425 ;
        RECT 82.965 160.925 83.205 161.575 ;
        RECT 78.295 160.270 78.480 160.295 ;
        RECT 77.865 160.170 78.480 160.270 ;
        RECT 77.865 159.615 78.470 160.170 ;
        RECT 78.645 159.785 79.125 160.125 ;
        RECT 79.295 159.615 79.550 160.160 ;
        RECT 79.720 159.785 79.995 160.485 ;
        RECT 80.165 159.615 81.375 160.705 ;
        RECT 81.555 160.395 82.450 160.725 ;
        RECT 82.620 160.565 83.205 160.755 ;
        RECT 81.555 160.225 82.760 160.395 ;
        RECT 81.555 159.795 81.885 160.225 ;
        RECT 82.065 159.615 82.260 160.055 ;
        RECT 82.430 159.795 82.760 160.225 ;
        RECT 82.930 159.795 83.205 160.565 ;
        RECT 83.390 160.565 83.725 161.985 ;
        RECT 83.905 161.795 84.650 162.165 ;
        RECT 85.215 161.625 85.470 161.985 ;
        RECT 85.650 161.795 85.980 162.165 ;
        RECT 86.160 161.625 86.385 161.985 ;
        RECT 83.900 161.435 86.385 161.625 ;
        RECT 83.900 160.745 84.125 161.435 ;
        RECT 86.605 161.415 87.815 162.165 ;
        RECT 87.990 161.660 88.325 162.165 ;
        RECT 88.495 161.595 88.735 161.970 ;
        RECT 89.015 161.835 89.185 161.980 ;
        RECT 89.015 161.640 89.390 161.835 ;
        RECT 89.750 161.670 90.145 162.165 ;
        RECT 84.325 160.925 84.605 161.255 ;
        RECT 84.785 160.925 85.360 161.255 ;
        RECT 85.540 160.925 85.975 161.255 ;
        RECT 86.155 160.925 86.425 161.255 ;
        RECT 86.605 160.875 87.125 161.415 ;
        RECT 83.900 160.565 86.395 160.745 ;
        RECT 87.295 160.705 87.815 161.245 ;
        RECT 83.390 159.795 83.655 160.565 ;
        RECT 83.825 159.615 84.155 160.335 ;
        RECT 84.345 160.155 85.535 160.385 ;
        RECT 84.345 159.795 84.605 160.155 ;
        RECT 84.775 159.615 85.105 159.985 ;
        RECT 85.275 159.795 85.535 160.155 ;
        RECT 86.105 159.795 86.395 160.565 ;
        RECT 86.605 159.615 87.815 160.705 ;
        RECT 88.045 160.635 88.345 161.485 ;
        RECT 88.515 161.445 88.735 161.595 ;
        RECT 88.515 161.115 89.050 161.445 ;
        RECT 89.220 161.305 89.390 161.640 ;
        RECT 90.315 161.475 90.555 161.995 ;
        RECT 88.515 160.465 88.750 161.115 ;
        RECT 89.220 160.945 90.205 161.305 ;
        RECT 88.075 160.235 88.750 160.465 ;
        RECT 88.920 160.925 90.205 160.945 ;
        RECT 88.920 160.775 89.780 160.925 ;
        RECT 88.075 159.805 88.245 160.235 ;
        RECT 88.415 159.615 88.745 160.065 ;
        RECT 88.920 159.830 89.205 160.775 ;
        RECT 90.380 160.670 90.555 161.475 ;
        RECT 89.380 160.295 90.075 160.605 ;
        RECT 89.385 159.615 90.070 160.085 ;
        RECT 90.250 159.885 90.555 160.670 ;
        RECT 90.770 161.410 91.005 161.740 ;
        RECT 91.175 161.425 91.505 162.165 ;
        RECT 91.740 161.785 92.935 161.995 ;
        RECT 90.770 160.755 90.940 161.410 ;
        RECT 91.740 161.345 92.015 161.785 ;
        RECT 92.185 161.345 92.515 161.615 ;
        RECT 92.685 161.555 92.935 161.785 ;
        RECT 93.105 161.725 93.275 162.165 ;
        RECT 93.445 161.555 93.795 161.995 ;
        RECT 92.685 161.345 93.795 161.555 ;
        RECT 93.985 161.475 94.225 161.995 ;
        RECT 94.395 161.670 94.790 162.165 ;
        RECT 95.355 161.835 95.525 161.980 ;
        RECT 95.150 161.640 95.525 161.835 ;
        RECT 92.185 161.315 92.470 161.345 ;
        RECT 91.115 160.925 91.460 161.255 ;
        RECT 91.690 160.755 92.020 161.175 ;
        RECT 90.770 160.585 92.020 160.755 ;
        RECT 90.770 160.390 91.070 160.585 ;
        RECT 92.190 160.415 92.470 161.315 ;
        RECT 92.650 160.975 93.795 161.175 ;
        RECT 92.650 160.805 92.840 160.975 ;
        RECT 92.645 160.635 92.840 160.805 ;
        RECT 92.650 160.595 92.840 160.635 ;
        RECT 93.020 160.415 93.295 160.755 ;
        RECT 91.240 159.615 91.495 160.415 ;
        RECT 91.695 160.245 93.295 160.415 ;
        RECT 91.695 159.785 92.025 160.245 ;
        RECT 92.195 159.615 92.770 160.075 ;
        RECT 92.940 159.785 93.295 160.245 ;
        RECT 93.465 159.615 93.795 160.755 ;
        RECT 93.985 160.670 94.160 161.475 ;
        RECT 95.150 161.305 95.320 161.640 ;
        RECT 95.805 161.595 96.045 161.970 ;
        RECT 96.215 161.660 96.550 162.165 ;
        RECT 95.805 161.445 96.025 161.595 ;
        RECT 94.335 160.945 95.320 161.305 ;
        RECT 95.490 161.115 96.025 161.445 ;
        RECT 94.335 160.925 95.620 160.945 ;
        RECT 94.760 160.775 95.620 160.925 ;
        RECT 93.985 159.885 94.290 160.670 ;
        RECT 94.465 160.295 95.160 160.605 ;
        RECT 94.470 159.615 95.155 160.085 ;
        RECT 95.335 159.830 95.620 160.775 ;
        RECT 95.790 160.465 96.025 161.115 ;
        RECT 96.195 160.635 96.495 161.485 ;
        RECT 96.725 161.365 96.985 162.165 ;
        RECT 95.790 160.235 96.465 160.465 ;
        RECT 95.795 159.615 96.125 160.065 ;
        RECT 96.295 159.805 96.465 160.235 ;
        RECT 96.725 159.615 96.985 160.755 ;
        RECT 97.155 159.785 97.485 161.995 ;
        RECT 97.735 161.425 98.065 162.165 ;
        RECT 98.335 161.595 98.665 161.995 ;
        RECT 98.835 161.765 99.165 162.165 ;
        RECT 99.335 161.825 100.695 161.995 ;
        RECT 99.335 161.595 99.665 161.825 ;
        RECT 98.335 161.425 99.665 161.595 ;
        RECT 99.835 161.425 100.165 161.655 ;
        RECT 97.655 160.465 97.965 161.255 ;
        RECT 98.135 160.635 98.355 161.255 ;
        RECT 98.625 160.635 98.800 161.255 ;
        RECT 99.055 160.635 99.275 161.255 ;
        RECT 99.550 160.805 99.795 161.255 ;
        RECT 99.545 160.635 99.795 160.805 ;
        RECT 99.965 160.465 100.165 161.425 ;
        RECT 100.335 161.345 100.695 161.825 ;
        RECT 100.865 161.440 101.155 162.165 ;
        RECT 101.330 161.535 101.665 161.995 ;
        RECT 101.835 161.705 102.030 162.165 ;
        RECT 102.275 161.785 104.300 161.995 ;
        RECT 101.330 161.345 102.020 161.535 ;
        RECT 102.275 161.345 102.525 161.785 ;
        RECT 102.695 161.345 103.880 161.615 ;
        RECT 104.050 161.535 104.300 161.785 ;
        RECT 104.470 161.705 104.640 162.165 ;
        RECT 104.810 161.535 105.140 161.995 ;
        RECT 105.310 161.705 105.550 162.165 ;
        RECT 105.760 161.535 106.090 161.995 ;
        RECT 104.050 161.345 106.090 161.535 ;
        RECT 106.410 161.410 106.645 161.740 ;
        RECT 106.815 161.425 107.145 162.165 ;
        RECT 107.380 161.785 108.575 161.995 ;
        RECT 101.850 161.175 102.020 161.345 ;
        RECT 100.335 161.005 100.695 161.175 ;
        RECT 100.365 160.925 100.695 161.005 ;
        RECT 101.350 160.975 101.680 161.175 ;
        RECT 101.850 160.975 103.445 161.175 ;
        RECT 101.850 160.805 102.020 160.975 ;
        RECT 103.615 160.805 103.880 161.345 ;
        RECT 104.395 160.975 106.180 161.175 ;
        RECT 97.655 160.295 100.165 160.465 ;
        RECT 97.655 159.615 98.165 160.125 ;
        RECT 99.335 159.785 99.665 160.295 ;
        RECT 100.335 159.615 100.695 160.755 ;
        RECT 100.865 159.615 101.155 160.780 ;
        RECT 101.330 160.585 102.020 160.805 ;
        RECT 101.330 159.785 101.665 160.585 ;
        RECT 102.210 160.415 102.525 160.805 ;
        RECT 101.835 159.615 102.525 160.415 ;
        RECT 102.695 160.585 105.560 160.805 ;
        RECT 106.410 160.755 106.580 161.410 ;
        RECT 107.380 161.345 107.655 161.785 ;
        RECT 107.825 161.445 108.155 161.615 ;
        RECT 107.830 161.345 108.155 161.445 ;
        RECT 108.325 161.555 108.575 161.785 ;
        RECT 108.745 161.725 108.915 162.165 ;
        RECT 109.085 161.555 109.435 161.995 ;
        RECT 109.605 161.655 109.910 162.165 ;
        RECT 108.325 161.345 109.435 161.555 ;
        RECT 106.755 160.925 107.100 161.255 ;
        RECT 107.330 160.755 107.660 161.175 ;
        RECT 102.695 159.785 103.025 160.585 ;
        RECT 103.195 159.615 103.365 160.415 ;
        RECT 103.535 159.785 103.880 160.585 ;
        RECT 104.050 159.615 104.220 160.415 ;
        RECT 104.390 159.785 104.720 160.585 ;
        RECT 104.890 159.615 105.060 160.415 ;
        RECT 105.230 159.785 105.560 160.585 ;
        RECT 105.760 159.615 106.090 160.755 ;
        RECT 106.410 160.585 107.660 160.755 ;
        RECT 106.410 160.390 106.710 160.585 ;
        RECT 107.830 160.415 108.110 161.345 ;
        RECT 108.290 160.975 109.435 161.175 ;
        RECT 108.290 160.805 108.480 160.975 ;
        RECT 109.605 160.925 109.920 161.485 ;
        RECT 110.090 161.175 110.340 161.985 ;
        RECT 110.510 161.640 110.770 162.165 ;
        RECT 110.950 161.175 111.200 161.985 ;
        RECT 111.370 161.605 111.630 162.165 ;
        RECT 111.800 161.515 112.060 161.970 ;
        RECT 112.230 161.685 112.490 162.165 ;
        RECT 112.660 161.515 112.920 161.970 ;
        RECT 113.090 161.685 113.350 162.165 ;
        RECT 113.520 161.515 113.780 161.970 ;
        RECT 113.950 161.685 114.195 162.165 ;
        RECT 114.365 161.515 114.640 161.970 ;
        RECT 114.810 161.685 115.055 162.165 ;
        RECT 115.225 161.515 115.485 161.970 ;
        RECT 115.665 161.685 115.915 162.165 ;
        RECT 116.085 161.515 116.345 161.970 ;
        RECT 116.525 161.685 116.775 162.165 ;
        RECT 116.945 161.515 117.205 161.970 ;
        RECT 117.385 161.685 117.645 162.165 ;
        RECT 117.815 161.515 118.075 161.970 ;
        RECT 118.245 161.685 118.545 162.165 ;
        RECT 111.800 161.345 118.545 161.515 ;
        RECT 118.815 161.445 119.145 162.165 ;
        RECT 119.315 161.495 119.485 161.955 ;
        RECT 119.655 161.785 119.985 162.165 ;
        RECT 120.215 161.615 120.425 161.995 ;
        RECT 120.595 161.785 120.925 162.165 ;
        RECT 121.095 161.785 122.765 161.955 ;
        RECT 121.095 161.615 121.265 161.785 ;
        RECT 110.090 160.925 117.210 161.175 ;
        RECT 108.285 160.635 108.480 160.805 ;
        RECT 108.745 160.755 108.915 160.805 ;
        RECT 108.290 160.595 108.480 160.635 ;
        RECT 108.660 160.415 108.935 160.755 ;
        RECT 106.880 159.615 107.135 160.415 ;
        RECT 107.335 160.245 108.935 160.415 ;
        RECT 107.335 159.785 107.665 160.245 ;
        RECT 107.835 159.615 108.410 160.075 ;
        RECT 108.580 159.785 108.935 160.245 ;
        RECT 109.105 159.615 109.435 160.755 ;
        RECT 109.615 159.615 109.910 160.425 ;
        RECT 110.090 159.785 110.335 160.925 ;
        RECT 110.510 159.615 110.770 160.425 ;
        RECT 110.950 159.790 111.200 160.925 ;
        RECT 117.380 160.755 118.545 161.345 ;
        RECT 111.800 160.530 118.545 160.755 ;
        RECT 111.800 160.515 117.205 160.530 ;
        RECT 111.370 159.620 111.630 160.415 ;
        RECT 111.800 159.790 112.060 160.515 ;
        RECT 112.230 159.620 112.490 160.345 ;
        RECT 112.660 159.790 112.920 160.515 ;
        RECT 113.090 159.620 113.350 160.345 ;
        RECT 113.520 159.790 113.780 160.515 ;
        RECT 113.950 159.620 114.210 160.345 ;
        RECT 114.380 159.790 114.640 160.515 ;
        RECT 114.810 159.620 115.055 160.345 ;
        RECT 115.225 159.790 115.485 160.515 ;
        RECT 115.670 159.620 115.915 160.345 ;
        RECT 116.085 159.790 116.345 160.515 ;
        RECT 116.530 159.620 116.775 160.345 ;
        RECT 116.945 159.790 117.205 160.515 ;
        RECT 117.390 159.620 117.645 160.345 ;
        RECT 117.815 159.790 118.105 160.530 ;
        RECT 111.370 159.615 117.645 159.620 ;
        RECT 118.275 159.615 118.545 160.360 ;
        RECT 118.815 159.615 119.145 160.755 ;
        RECT 119.315 159.785 119.505 161.495 ;
        RECT 119.700 161.445 121.265 161.615 ;
        RECT 119.700 160.755 119.870 161.445 ;
        RECT 120.120 160.955 120.450 161.175 ;
        RECT 120.720 161.145 121.055 161.255 ;
        RECT 120.705 160.975 121.055 161.145 ;
        RECT 119.700 160.585 120.505 160.755 ;
        RECT 120.720 160.625 121.055 160.975 ;
        RECT 121.405 160.815 121.575 161.255 ;
        RECT 122.055 161.175 122.270 161.505 ;
        RECT 121.805 161.005 122.270 161.175 ;
        RECT 121.405 160.625 121.810 160.815 ;
        RECT 122.055 160.625 122.270 161.005 ;
        RECT 122.505 160.625 122.725 161.520 ;
        RECT 122.955 161.400 123.405 162.165 ;
        RECT 123.680 161.745 125.005 161.995 ;
        RECT 123.880 161.175 124.100 161.575 ;
        RECT 122.950 160.975 123.435 161.175 ;
        RECT 123.625 160.965 124.100 161.175 ;
        RECT 124.370 161.175 124.580 161.575 ;
        RECT 124.835 161.515 125.005 161.745 ;
        RECT 125.215 161.685 125.545 162.165 ;
        RECT 125.760 161.665 126.020 161.995 ;
        RECT 124.835 161.345 125.675 161.515 ;
        RECT 124.370 160.965 124.700 161.175 ;
        RECT 124.870 160.975 125.275 161.175 ;
        RECT 125.505 160.795 125.675 161.345 ;
        RECT 122.955 160.625 125.675 160.795 ;
        RECT 119.735 159.615 119.985 160.415 ;
        RECT 120.175 159.825 120.505 160.585 ;
        RECT 120.675 160.285 122.685 160.455 ;
        RECT 120.675 159.785 120.845 160.285 ;
        RECT 121.055 159.615 121.305 160.075 ;
        RECT 121.515 159.785 121.685 160.285 ;
        RECT 122.055 159.615 122.305 160.075 ;
        RECT 122.515 159.785 122.685 160.285 ;
        RECT 122.955 159.955 123.285 160.625 ;
        RECT 125.850 160.465 126.020 161.665 ;
        RECT 126.190 161.265 126.360 162.165 ;
        RECT 126.625 161.440 126.915 162.165 ;
        RECT 128.025 161.805 128.365 162.165 ;
        RECT 128.895 161.805 129.225 162.165 ;
        RECT 129.830 161.805 130.605 162.165 ;
        RECT 130.795 161.635 130.965 161.995 ;
        RECT 131.175 161.805 131.505 162.165 ;
        RECT 128.065 161.465 129.655 161.635 ;
        RECT 129.955 161.580 130.965 161.635 ;
        RECT 132.005 161.580 132.285 161.845 ;
        RECT 129.955 161.465 132.285 161.580 ;
        RECT 123.455 160.215 125.090 160.455 ;
        RECT 123.455 160.125 123.685 160.215 ;
        RECT 123.795 159.955 124.125 159.995 ;
        RECT 122.955 159.785 124.125 159.955 ;
        RECT 124.315 159.615 124.670 160.035 ;
        RECT 124.840 159.785 125.090 160.215 ;
        RECT 125.260 159.615 125.590 160.375 ;
        RECT 125.760 159.785 126.020 160.465 ;
        RECT 126.190 159.615 126.360 160.805 ;
        RECT 126.625 159.615 126.915 160.780 ;
        RECT 128.065 160.665 128.550 161.465 ;
        RECT 129.955 161.255 130.125 161.465 ;
        RECT 130.795 161.410 132.285 161.465 ;
        RECT 128.720 160.925 130.125 161.255 ;
        RECT 128.065 160.495 129.655 160.665 ;
        RECT 128.035 159.615 128.365 160.315 ;
        RECT 128.545 160.065 128.715 160.495 ;
        RECT 128.895 159.615 129.225 160.315 ;
        RECT 129.405 160.065 129.655 160.495 ;
        RECT 129.835 159.615 130.085 160.735 ;
        RECT 130.315 160.725 130.625 161.255 ;
        RECT 130.375 159.955 130.545 160.555 ;
        RECT 130.795 160.125 130.965 161.410 ;
        RECT 132.865 161.365 133.145 162.165 ;
        RECT 133.565 161.345 133.795 162.165 ;
        RECT 133.965 161.365 134.295 161.995 ;
        RECT 131.345 161.145 131.740 161.240 ;
        RECT 131.285 160.975 131.740 161.145 ;
        RECT 131.910 160.975 132.435 161.240 ;
        RECT 131.205 160.400 131.385 160.805 ;
        RECT 131.565 160.740 131.740 160.975 ;
        RECT 132.605 160.960 133.020 161.195 ;
        RECT 132.605 160.740 132.855 160.960 ;
        RECT 133.545 160.925 133.875 161.175 ;
        RECT 131.565 160.570 132.855 160.740 ;
        RECT 133.025 160.400 133.280 160.790 ;
        RECT 134.045 160.765 134.295 161.365 ;
        RECT 134.465 161.345 134.675 162.165 ;
        RECT 134.905 161.415 136.115 162.165 ;
        RECT 131.205 160.230 133.280 160.400 ;
        RECT 131.205 159.955 131.385 160.230 ;
        RECT 130.375 159.785 131.385 159.955 ;
        RECT 131.555 159.615 131.885 159.975 ;
        RECT 132.055 159.785 132.225 160.230 ;
        RECT 132.395 159.615 132.725 159.975 ;
        RECT 132.950 159.855 133.280 160.230 ;
        RECT 133.565 159.615 133.795 160.755 ;
        RECT 133.965 159.785 134.295 160.765 ;
        RECT 134.465 159.615 134.675 160.755 ;
        RECT 134.905 160.705 135.425 161.245 ;
        RECT 135.595 160.875 136.115 161.415 ;
        RECT 134.905 159.615 136.115 160.705 ;
        RECT 23.500 159.445 136.200 159.615 ;
        RECT 23.585 158.355 24.795 159.445 ;
        RECT 24.965 159.010 30.310 159.445 ;
        RECT 30.485 159.010 35.830 159.445 ;
        RECT 23.585 157.645 24.105 158.185 ;
        RECT 24.275 157.815 24.795 158.355 ;
        RECT 23.585 156.895 24.795 157.645 ;
        RECT 26.550 157.440 26.890 158.270 ;
        RECT 28.370 157.760 28.720 159.010 ;
        RECT 32.070 157.440 32.410 158.270 ;
        RECT 33.890 157.760 34.240 159.010 ;
        RECT 36.465 158.280 36.755 159.445 ;
        RECT 36.925 159.010 42.270 159.445 ;
        RECT 42.445 159.010 47.790 159.445 ;
        RECT 47.965 159.010 53.310 159.445 ;
        RECT 24.965 156.895 30.310 157.440 ;
        RECT 30.485 156.895 35.830 157.440 ;
        RECT 36.465 156.895 36.755 157.620 ;
        RECT 38.510 157.440 38.850 158.270 ;
        RECT 40.330 157.760 40.680 159.010 ;
        RECT 44.030 157.440 44.370 158.270 ;
        RECT 45.850 157.760 46.200 159.010 ;
        RECT 49.550 157.440 49.890 158.270 ;
        RECT 51.370 157.760 51.720 159.010 ;
        RECT 53.495 158.835 53.825 159.265 ;
        RECT 54.005 159.005 54.200 159.445 ;
        RECT 54.370 158.835 54.700 159.265 ;
        RECT 53.495 158.665 54.700 158.835 ;
        RECT 53.495 158.335 54.390 158.665 ;
        RECT 54.870 158.495 55.145 159.265 ;
        RECT 54.560 158.305 55.145 158.495 ;
        RECT 55.345 158.555 55.605 159.265 ;
        RECT 55.775 158.735 56.105 159.445 ;
        RECT 56.275 158.555 56.505 159.265 ;
        RECT 55.345 158.315 56.505 158.555 ;
        RECT 56.685 158.535 56.955 159.265 ;
        RECT 57.135 158.715 57.475 159.445 ;
        RECT 56.685 158.315 57.455 158.535 ;
        RECT 53.500 157.805 53.795 158.135 ;
        RECT 53.975 157.805 54.390 158.135 ;
        RECT 36.925 156.895 42.270 157.440 ;
        RECT 42.445 156.895 47.790 157.440 ;
        RECT 47.965 156.895 53.310 157.440 ;
        RECT 53.495 156.895 53.795 157.625 ;
        RECT 53.975 157.185 54.205 157.805 ;
        RECT 54.560 157.635 54.735 158.305 ;
        RECT 54.405 157.455 54.735 157.635 ;
        RECT 54.905 157.485 55.145 158.135 ;
        RECT 55.335 157.805 55.635 158.135 ;
        RECT 55.815 157.825 56.340 158.135 ;
        RECT 56.520 157.825 56.985 158.135 ;
        RECT 54.405 157.075 54.630 157.455 ;
        RECT 54.800 156.895 55.130 157.285 ;
        RECT 55.345 156.895 55.635 157.625 ;
        RECT 55.815 157.185 56.045 157.825 ;
        RECT 57.165 157.645 57.455 158.315 ;
        RECT 56.225 157.445 57.455 157.645 ;
        RECT 56.225 157.075 56.535 157.445 ;
        RECT 56.715 156.895 57.385 157.265 ;
        RECT 57.645 157.075 57.905 159.265 ;
        RECT 59.005 158.265 59.325 159.445 ;
        RECT 59.495 158.425 59.695 159.215 ;
        RECT 60.020 158.615 60.405 159.275 ;
        RECT 60.800 158.685 61.585 159.445 ;
        RECT 59.995 158.515 60.405 158.615 ;
        RECT 59.495 158.255 59.825 158.425 ;
        RECT 59.995 158.305 61.605 158.515 ;
        RECT 59.645 158.135 59.825 158.255 ;
        RECT 59.005 157.885 59.470 158.085 ;
        RECT 59.645 157.885 59.975 158.135 ;
        RECT 60.145 158.085 60.610 158.135 ;
        RECT 60.145 157.915 60.615 158.085 ;
        RECT 60.145 157.885 60.610 157.915 ;
        RECT 60.805 157.885 61.160 158.135 ;
        RECT 61.330 157.705 61.605 158.305 ;
        RECT 59.005 157.505 60.185 157.675 ;
        RECT 59.005 157.090 59.345 157.505 ;
        RECT 59.515 156.895 59.685 157.335 ;
        RECT 59.855 157.285 60.185 157.505 ;
        RECT 60.355 157.525 61.605 157.705 ;
        RECT 60.355 157.455 60.720 157.525 ;
        RECT 59.855 157.105 61.105 157.285 ;
        RECT 61.375 156.895 61.545 157.355 ;
        RECT 61.775 157.175 62.055 159.275 ;
        RECT 62.225 158.280 62.515 159.445 ;
        RECT 62.685 158.265 63.005 159.445 ;
        RECT 63.175 158.425 63.375 159.215 ;
        RECT 63.700 158.615 64.085 159.275 ;
        RECT 64.480 158.685 65.265 159.445 ;
        RECT 63.675 158.515 64.085 158.615 ;
        RECT 63.175 158.255 63.505 158.425 ;
        RECT 63.675 158.305 65.285 158.515 ;
        RECT 63.325 158.135 63.505 158.255 ;
        RECT 62.685 157.885 63.150 158.085 ;
        RECT 63.325 157.885 63.655 158.135 ;
        RECT 63.825 158.085 64.290 158.135 ;
        RECT 63.825 157.915 64.295 158.085 ;
        RECT 63.825 157.885 64.290 157.915 ;
        RECT 64.485 157.885 64.840 158.135 ;
        RECT 65.010 157.705 65.285 158.305 ;
        RECT 62.225 156.895 62.515 157.620 ;
        RECT 62.685 157.505 63.865 157.675 ;
        RECT 62.685 157.090 63.025 157.505 ;
        RECT 63.195 156.895 63.365 157.335 ;
        RECT 63.535 157.285 63.865 157.505 ;
        RECT 64.035 157.525 65.285 157.705 ;
        RECT 64.035 157.455 64.400 157.525 ;
        RECT 63.535 157.105 64.785 157.285 ;
        RECT 65.055 156.895 65.225 157.355 ;
        RECT 65.455 157.175 65.735 159.275 ;
        RECT 65.925 158.555 66.185 159.265 ;
        RECT 66.355 158.735 66.685 159.445 ;
        RECT 66.855 158.555 67.085 159.265 ;
        RECT 65.925 158.315 67.085 158.555 ;
        RECT 67.265 158.535 67.535 159.265 ;
        RECT 67.715 158.715 68.055 159.445 ;
        RECT 67.265 158.315 68.035 158.535 ;
        RECT 65.915 157.805 66.215 158.135 ;
        RECT 66.395 157.825 66.920 158.135 ;
        RECT 67.100 157.825 67.565 158.135 ;
        RECT 65.925 156.895 66.215 157.625 ;
        RECT 66.395 157.185 66.625 157.825 ;
        RECT 67.745 157.645 68.035 158.315 ;
        RECT 66.805 157.445 68.035 157.645 ;
        RECT 66.805 157.075 67.115 157.445 ;
        RECT 67.295 156.895 67.965 157.265 ;
        RECT 68.225 157.075 68.485 159.265 ;
        RECT 68.705 158.305 68.935 159.445 ;
        RECT 69.105 158.295 69.435 159.275 ;
        RECT 69.605 158.305 69.815 159.445 ;
        RECT 70.045 158.890 70.650 159.445 ;
        RECT 70.825 158.935 71.305 159.275 ;
        RECT 71.475 158.900 71.730 159.445 ;
        RECT 70.045 158.790 70.660 158.890 ;
        RECT 70.475 158.765 70.660 158.790 ;
        RECT 68.685 157.885 69.015 158.135 ;
        RECT 68.705 156.895 68.935 157.715 ;
        RECT 69.185 157.695 69.435 158.295 ;
        RECT 70.045 158.170 70.305 158.620 ;
        RECT 70.475 158.520 70.805 158.765 ;
        RECT 70.975 158.445 71.730 158.695 ;
        RECT 71.900 158.575 72.175 159.275 ;
        RECT 70.960 158.410 71.730 158.445 ;
        RECT 70.945 158.400 71.730 158.410 ;
        RECT 70.940 158.385 71.835 158.400 ;
        RECT 70.920 158.370 71.835 158.385 ;
        RECT 70.900 158.360 71.835 158.370 ;
        RECT 70.875 158.350 71.835 158.360 ;
        RECT 70.805 158.320 71.835 158.350 ;
        RECT 70.785 158.290 71.835 158.320 ;
        RECT 70.765 158.260 71.835 158.290 ;
        RECT 70.735 158.235 71.835 158.260 ;
        RECT 70.700 158.200 71.835 158.235 ;
        RECT 70.670 158.195 71.835 158.200 ;
        RECT 70.670 158.190 71.060 158.195 ;
        RECT 70.670 158.180 71.035 158.190 ;
        RECT 70.670 158.175 71.020 158.180 ;
        RECT 70.670 158.170 71.005 158.175 ;
        RECT 70.045 158.165 71.005 158.170 ;
        RECT 70.045 158.155 70.995 158.165 ;
        RECT 70.045 158.150 70.985 158.155 ;
        RECT 70.045 158.140 70.975 158.150 ;
        RECT 70.045 158.130 70.970 158.140 ;
        RECT 70.045 158.125 70.965 158.130 ;
        RECT 70.045 158.110 70.955 158.125 ;
        RECT 70.045 158.095 70.950 158.110 ;
        RECT 70.045 158.070 70.940 158.095 ;
        RECT 70.045 158.000 70.935 158.070 ;
        RECT 69.105 157.065 69.435 157.695 ;
        RECT 69.605 156.895 69.815 157.715 ;
        RECT 70.045 157.445 70.595 157.830 ;
        RECT 70.765 157.275 70.935 158.000 ;
        RECT 70.045 157.105 70.935 157.275 ;
        RECT 71.105 157.600 71.435 158.025 ;
        RECT 71.605 157.800 71.835 158.195 ;
        RECT 71.105 157.575 71.355 157.600 ;
        RECT 71.105 157.115 71.325 157.575 ;
        RECT 72.005 157.545 72.175 158.575 ;
        RECT 72.345 158.265 72.665 159.445 ;
        RECT 72.835 158.425 73.035 159.215 ;
        RECT 73.360 158.615 73.745 159.275 ;
        RECT 74.140 158.685 74.925 159.445 ;
        RECT 73.335 158.515 73.745 158.615 ;
        RECT 72.835 158.255 73.165 158.425 ;
        RECT 73.335 158.305 74.945 158.515 ;
        RECT 72.985 158.135 73.165 158.255 ;
        RECT 72.345 157.885 72.810 158.085 ;
        RECT 72.985 157.885 73.315 158.135 ;
        RECT 73.485 158.085 73.950 158.135 ;
        RECT 73.485 157.915 73.955 158.085 ;
        RECT 73.485 157.885 73.950 157.915 ;
        RECT 74.145 157.885 74.500 158.135 ;
        RECT 74.670 157.705 74.945 158.305 ;
        RECT 71.495 156.895 71.745 157.435 ;
        RECT 71.915 157.065 72.175 157.545 ;
        RECT 72.345 157.505 73.525 157.675 ;
        RECT 72.345 157.090 72.685 157.505 ;
        RECT 72.855 156.895 73.025 157.335 ;
        RECT 73.195 157.285 73.525 157.505 ;
        RECT 73.695 157.525 74.945 157.705 ;
        RECT 73.695 157.455 74.060 157.525 ;
        RECT 73.195 157.105 74.445 157.285 ;
        RECT 74.715 156.895 74.885 157.355 ;
        RECT 75.115 157.175 75.395 159.275 ;
        RECT 75.565 158.890 76.170 159.445 ;
        RECT 76.345 158.935 76.825 159.275 ;
        RECT 76.995 158.900 77.250 159.445 ;
        RECT 75.565 158.790 76.180 158.890 ;
        RECT 75.995 158.765 76.180 158.790 ;
        RECT 75.565 158.170 75.825 158.620 ;
        RECT 75.995 158.520 76.325 158.765 ;
        RECT 76.495 158.445 77.250 158.695 ;
        RECT 77.420 158.575 77.695 159.275 ;
        RECT 77.865 158.935 79.055 159.225 ;
        RECT 76.480 158.410 77.250 158.445 ;
        RECT 76.465 158.400 77.250 158.410 ;
        RECT 76.460 158.385 77.355 158.400 ;
        RECT 76.440 158.370 77.355 158.385 ;
        RECT 76.420 158.360 77.355 158.370 ;
        RECT 76.395 158.350 77.355 158.360 ;
        RECT 76.325 158.320 77.355 158.350 ;
        RECT 76.305 158.290 77.355 158.320 ;
        RECT 76.285 158.260 77.355 158.290 ;
        RECT 76.255 158.235 77.355 158.260 ;
        RECT 76.220 158.200 77.355 158.235 ;
        RECT 76.190 158.195 77.355 158.200 ;
        RECT 76.190 158.190 76.580 158.195 ;
        RECT 76.190 158.180 76.555 158.190 ;
        RECT 76.190 158.175 76.540 158.180 ;
        RECT 76.190 158.170 76.525 158.175 ;
        RECT 75.565 158.165 76.525 158.170 ;
        RECT 75.565 158.155 76.515 158.165 ;
        RECT 75.565 158.150 76.505 158.155 ;
        RECT 75.565 158.140 76.495 158.150 ;
        RECT 75.565 158.130 76.490 158.140 ;
        RECT 75.565 158.125 76.485 158.130 ;
        RECT 75.565 158.110 76.475 158.125 ;
        RECT 75.565 158.095 76.470 158.110 ;
        RECT 75.565 158.070 76.460 158.095 ;
        RECT 75.565 158.000 76.455 158.070 ;
        RECT 75.565 157.445 76.115 157.830 ;
        RECT 76.285 157.275 76.455 158.000 ;
        RECT 75.565 157.105 76.455 157.275 ;
        RECT 76.625 157.600 76.955 158.025 ;
        RECT 77.125 157.800 77.355 158.195 ;
        RECT 76.625 157.115 76.845 157.600 ;
        RECT 77.525 157.545 77.695 158.575 ;
        RECT 77.885 158.595 79.055 158.765 ;
        RECT 79.225 158.645 79.505 159.445 ;
        RECT 77.885 158.305 78.210 158.595 ;
        RECT 78.885 158.475 79.055 158.595 ;
        RECT 78.380 158.135 78.575 158.425 ;
        RECT 78.885 158.305 79.545 158.475 ;
        RECT 79.715 158.305 79.990 159.275 ;
        RECT 80.380 158.345 80.710 159.445 ;
        RECT 81.185 158.845 81.510 159.275 ;
        RECT 81.680 159.025 82.010 159.445 ;
        RECT 82.755 159.015 83.165 159.445 ;
        RECT 81.185 158.675 83.165 158.845 ;
        RECT 79.375 158.135 79.545 158.305 ;
        RECT 77.865 157.805 78.210 158.135 ;
        RECT 78.380 157.805 79.205 158.135 ;
        RECT 79.375 157.805 79.650 158.135 ;
        RECT 79.375 157.635 79.545 157.805 ;
        RECT 77.015 156.895 77.265 157.435 ;
        RECT 77.435 157.065 77.695 157.545 ;
        RECT 77.880 157.465 79.545 157.635 ;
        RECT 79.820 157.570 79.990 158.305 ;
        RECT 81.185 158.265 81.890 158.675 ;
        RECT 80.165 157.885 80.810 158.095 ;
        RECT 80.980 157.885 81.550 158.095 ;
        RECT 77.880 157.115 78.135 157.465 ;
        RECT 78.305 156.895 78.635 157.295 ;
        RECT 78.805 157.115 78.975 157.465 ;
        RECT 79.145 156.895 79.525 157.295 ;
        RECT 79.715 157.225 79.990 157.570 ;
        RECT 80.320 157.545 81.490 157.715 ;
        RECT 80.320 157.080 80.650 157.545 ;
        RECT 80.820 156.895 80.990 157.365 ;
        RECT 81.160 157.065 81.490 157.545 ;
        RECT 81.720 157.065 81.890 158.265 ;
        RECT 82.060 158.335 82.685 158.505 ;
        RECT 82.060 157.635 82.230 158.335 ;
        RECT 82.900 158.135 83.165 158.675 ;
        RECT 83.335 158.290 83.675 159.275 ;
        RECT 83.855 158.645 84.185 159.445 ;
        RECT 84.365 159.105 85.795 159.275 ;
        RECT 84.365 158.475 84.615 159.105 ;
        RECT 82.400 157.805 82.730 158.135 ;
        RECT 82.900 157.805 83.250 158.135 ;
        RECT 83.420 157.635 83.675 158.290 ;
        RECT 82.060 157.465 82.600 157.635 ;
        RECT 82.430 157.260 82.600 157.465 ;
        RECT 82.880 156.895 83.050 157.635 ;
        RECT 83.315 157.260 83.675 157.635 ;
        RECT 83.845 158.305 84.615 158.475 ;
        RECT 83.845 157.635 84.015 158.305 ;
        RECT 84.185 157.805 84.590 158.135 ;
        RECT 84.805 157.805 85.055 158.935 ;
        RECT 85.255 158.135 85.455 158.935 ;
        RECT 85.625 158.425 85.795 159.105 ;
        RECT 85.965 158.595 86.280 159.445 ;
        RECT 86.455 158.645 86.895 159.275 ;
        RECT 85.625 158.255 86.415 158.425 ;
        RECT 85.255 157.805 85.500 158.135 ;
        RECT 85.685 157.805 86.075 158.085 ;
        RECT 86.245 157.805 86.415 158.255 ;
        RECT 86.585 157.635 86.895 158.645 ;
        RECT 87.985 158.280 88.275 159.445 ;
        RECT 88.465 158.605 88.795 159.445 ;
        RECT 88.965 158.425 89.310 159.180 ;
        RECT 89.485 158.835 89.830 159.275 ;
        RECT 90.040 159.065 90.370 159.445 ;
        RECT 90.555 158.835 90.790 159.275 ;
        RECT 90.960 159.005 91.290 159.445 ;
        RECT 89.485 158.595 91.495 158.835 ;
        RECT 88.465 157.815 88.795 158.425 ;
        RECT 88.965 157.805 89.595 158.425 ;
        RECT 89.765 157.805 90.055 158.425 ;
        RECT 83.445 157.235 83.615 157.260 ;
        RECT 83.845 157.065 84.335 157.635 ;
        RECT 84.505 157.465 85.665 157.635 ;
        RECT 84.505 157.065 84.735 157.465 ;
        RECT 84.905 156.895 85.325 157.295 ;
        RECT 85.495 157.065 85.665 157.465 ;
        RECT 85.835 156.895 86.285 157.635 ;
        RECT 86.455 157.075 86.895 157.635 ;
        RECT 87.985 156.895 88.275 157.620 ;
        RECT 88.465 157.435 89.830 157.635 ;
        RECT 88.465 157.065 88.795 157.435 ;
        RECT 88.965 156.895 89.295 157.265 ;
        RECT 89.485 157.065 89.830 157.435 ;
        RECT 90.225 157.065 90.555 158.425 ;
        RECT 90.765 157.885 91.095 158.425 ;
        RECT 91.265 157.695 91.495 158.595 ;
        RECT 90.890 157.065 91.495 157.695 ;
        RECT 92.150 158.475 92.450 158.670 ;
        RECT 92.620 158.645 92.875 159.445 ;
        RECT 93.075 158.815 93.405 159.275 ;
        RECT 93.575 158.985 94.150 159.445 ;
        RECT 94.320 158.815 94.675 159.275 ;
        RECT 93.075 158.645 94.675 158.815 ;
        RECT 93.565 158.595 93.850 158.645 ;
        RECT 92.150 158.305 93.400 158.475 ;
        RECT 92.150 157.650 92.320 158.305 ;
        RECT 92.495 157.805 92.840 158.135 ;
        RECT 93.070 157.885 93.400 158.305 ;
        RECT 93.570 157.715 93.850 158.595 ;
        RECT 94.030 158.085 94.220 158.465 ;
        RECT 94.400 158.305 94.675 158.645 ;
        RECT 94.845 158.305 95.175 159.445 ;
        RECT 95.435 158.865 95.605 159.275 ;
        RECT 95.775 159.065 96.105 159.445 ;
        RECT 96.750 159.065 97.420 159.445 ;
        RECT 97.655 158.895 97.825 159.275 ;
        RECT 97.995 159.065 98.335 159.445 ;
        RECT 98.505 158.895 98.675 159.275 ;
        RECT 99.015 159.065 99.345 159.445 ;
        RECT 99.515 158.895 99.775 159.275 ;
        RECT 95.435 158.695 97.185 158.865 ;
        RECT 95.410 158.085 95.590 158.445 ;
        RECT 94.030 157.885 95.175 158.085 ;
        RECT 95.405 157.915 95.590 158.085 ;
        RECT 95.410 157.805 95.590 157.915 ;
        RECT 92.150 157.320 92.385 157.650 ;
        RECT 92.555 156.895 92.885 157.635 ;
        RECT 93.120 157.275 93.395 157.715 ;
        RECT 93.570 157.615 93.895 157.715 ;
        RECT 93.565 157.445 93.895 157.615 ;
        RECT 94.065 157.505 95.175 157.715 ;
        RECT 95.760 157.615 95.930 158.695 ;
        RECT 96.250 158.355 96.580 158.525 ;
        RECT 94.065 157.275 94.315 157.505 ;
        RECT 93.120 157.065 94.315 157.275 ;
        RECT 94.485 156.895 94.655 157.335 ;
        RECT 94.825 157.065 95.175 157.505 ;
        RECT 95.435 157.445 95.930 157.615 ;
        RECT 95.435 157.065 95.605 157.445 ;
        RECT 95.775 156.895 96.105 157.275 ;
        RECT 96.275 157.065 96.500 158.355 ;
        RECT 97.015 158.135 97.185 158.695 ;
        RECT 97.495 158.725 98.675 158.895 ;
        RECT 98.845 158.725 99.775 158.895 ;
        RECT 96.675 157.615 96.845 158.135 ;
        RECT 97.015 157.805 97.325 158.135 ;
        RECT 97.495 157.615 97.665 158.725 ;
        RECT 98.845 158.555 99.015 158.725 ;
        RECT 97.835 158.385 99.015 158.555 ;
        RECT 97.835 158.210 98.005 158.385 ;
        RECT 98.165 157.915 98.435 158.085 ;
        RECT 96.675 157.445 97.665 157.615 ;
        RECT 96.670 156.895 97.000 157.275 ;
        RECT 97.270 157.065 97.440 157.445 ;
        RECT 98.170 157.230 98.435 157.915 ;
        RECT 98.610 157.235 98.915 158.215 ;
        RECT 99.085 157.575 99.435 158.115 ;
        RECT 99.605 157.395 99.775 158.725 ;
        RECT 100.410 158.575 100.675 159.275 ;
        RECT 100.845 158.745 101.175 159.445 ;
        RECT 101.345 158.575 102.015 159.275 ;
        RECT 102.520 158.745 102.950 159.445 ;
        RECT 103.130 158.885 103.320 159.275 ;
        RECT 103.490 159.065 103.820 159.445 ;
        RECT 103.130 158.715 103.860 158.885 ;
        RECT 100.410 158.320 102.985 158.575 ;
        RECT 100.405 157.805 100.680 158.135 ;
        RECT 100.850 157.635 101.030 158.320 ;
        RECT 102.815 158.135 102.985 158.320 ;
        RECT 101.200 157.805 101.560 158.135 ;
        RECT 101.850 158.085 102.140 158.135 ;
        RECT 101.845 157.915 102.140 158.085 ;
        RECT 101.850 157.805 102.140 157.915 ;
        RECT 102.310 157.805 102.645 158.135 ;
        RECT 102.815 157.805 103.495 158.135 ;
        RECT 99.095 156.895 99.345 157.395 ;
        RECT 99.515 157.065 99.775 157.395 ;
        RECT 100.415 157.235 101.030 157.635 ;
        RECT 101.200 157.445 102.470 157.635 ;
        RECT 103.665 157.595 103.860 158.715 ;
        RECT 104.175 158.700 104.445 159.445 ;
        RECT 105.075 159.440 111.350 159.445 ;
        RECT 104.615 158.530 104.905 159.270 ;
        RECT 105.075 158.715 105.330 159.440 ;
        RECT 105.515 158.545 105.775 159.270 ;
        RECT 105.945 158.715 106.190 159.440 ;
        RECT 106.375 158.545 106.635 159.270 ;
        RECT 106.805 158.715 107.050 159.440 ;
        RECT 107.235 158.545 107.495 159.270 ;
        RECT 107.665 158.715 107.910 159.440 ;
        RECT 108.080 158.545 108.340 159.270 ;
        RECT 108.510 158.715 108.770 159.440 ;
        RECT 108.940 158.545 109.200 159.270 ;
        RECT 109.370 158.715 109.630 159.440 ;
        RECT 109.800 158.545 110.060 159.270 ;
        RECT 110.230 158.715 110.490 159.440 ;
        RECT 110.660 158.545 110.920 159.270 ;
        RECT 111.090 158.645 111.350 159.440 ;
        RECT 105.515 158.530 110.920 158.545 ;
        RECT 103.040 157.425 103.860 157.595 ;
        RECT 104.175 158.305 110.920 158.530 ;
        RECT 104.175 157.715 105.340 158.305 ;
        RECT 111.520 158.135 111.770 159.270 ;
        RECT 111.950 158.635 112.210 159.445 ;
        RECT 112.385 158.135 112.630 159.275 ;
        RECT 112.810 158.635 113.105 159.445 ;
        RECT 113.745 158.280 114.035 159.445 ;
        RECT 114.215 158.635 114.510 159.445 ;
        RECT 114.690 158.135 114.935 159.275 ;
        RECT 115.110 158.635 115.370 159.445 ;
        RECT 115.970 159.440 122.245 159.445 ;
        RECT 115.550 158.135 115.800 159.270 ;
        RECT 115.970 158.645 116.230 159.440 ;
        RECT 116.400 158.545 116.660 159.270 ;
        RECT 116.830 158.715 117.090 159.440 ;
        RECT 117.260 158.545 117.520 159.270 ;
        RECT 117.690 158.715 117.950 159.440 ;
        RECT 118.120 158.545 118.380 159.270 ;
        RECT 118.550 158.715 118.810 159.440 ;
        RECT 118.980 158.545 119.240 159.270 ;
        RECT 119.410 158.715 119.655 159.440 ;
        RECT 119.825 158.545 120.085 159.270 ;
        RECT 120.270 158.715 120.515 159.440 ;
        RECT 120.685 158.545 120.945 159.270 ;
        RECT 121.130 158.715 121.375 159.440 ;
        RECT 121.545 158.545 121.805 159.270 ;
        RECT 121.990 158.715 122.245 159.440 ;
        RECT 116.400 158.530 121.805 158.545 ;
        RECT 122.415 158.530 122.705 159.270 ;
        RECT 122.875 158.700 123.145 159.445 ;
        RECT 123.415 158.635 123.710 159.445 ;
        RECT 116.400 158.305 123.145 158.530 ;
        RECT 105.510 157.885 112.630 158.135 ;
        RECT 104.175 157.545 110.920 157.715 ;
        RECT 100.415 157.065 100.750 157.235 ;
        RECT 101.710 156.895 102.045 157.275 ;
        RECT 102.635 156.895 102.870 157.335 ;
        RECT 103.040 157.065 103.370 157.425 ;
        RECT 103.540 156.895 103.870 157.255 ;
        RECT 104.175 156.895 104.475 157.375 ;
        RECT 104.645 157.090 104.905 157.545 ;
        RECT 105.075 156.895 105.335 157.375 ;
        RECT 105.515 157.090 105.775 157.545 ;
        RECT 105.945 156.895 106.195 157.375 ;
        RECT 106.375 157.090 106.635 157.545 ;
        RECT 106.805 156.895 107.055 157.375 ;
        RECT 107.235 157.090 107.495 157.545 ;
        RECT 107.665 156.895 107.910 157.375 ;
        RECT 108.080 157.090 108.355 157.545 ;
        RECT 108.525 156.895 108.770 157.375 ;
        RECT 108.940 157.090 109.200 157.545 ;
        RECT 109.370 156.895 109.630 157.375 ;
        RECT 109.800 157.090 110.060 157.545 ;
        RECT 110.230 156.895 110.490 157.375 ;
        RECT 110.660 157.090 110.920 157.545 ;
        RECT 111.090 156.895 111.350 157.455 ;
        RECT 111.520 157.075 111.770 157.885 ;
        RECT 111.950 156.895 112.210 157.420 ;
        RECT 112.380 157.075 112.630 157.885 ;
        RECT 112.800 157.575 113.115 158.135 ;
        RECT 112.810 156.895 113.115 157.405 ;
        RECT 113.745 156.895 114.035 157.620 ;
        RECT 114.205 157.575 114.520 158.135 ;
        RECT 114.690 157.885 121.810 158.135 ;
        RECT 114.205 156.895 114.510 157.405 ;
        RECT 114.690 157.075 114.940 157.885 ;
        RECT 115.110 156.895 115.370 157.420 ;
        RECT 115.550 157.075 115.800 157.885 ;
        RECT 121.980 157.715 123.145 158.305 ;
        RECT 123.890 158.135 124.135 159.275 ;
        RECT 124.310 158.635 124.570 159.445 ;
        RECT 125.170 159.440 131.445 159.445 ;
        RECT 124.750 158.135 125.000 159.270 ;
        RECT 125.170 158.645 125.430 159.440 ;
        RECT 125.600 158.545 125.860 159.270 ;
        RECT 126.030 158.715 126.290 159.440 ;
        RECT 126.460 158.545 126.720 159.270 ;
        RECT 126.890 158.715 127.150 159.440 ;
        RECT 127.320 158.545 127.580 159.270 ;
        RECT 127.750 158.715 128.010 159.440 ;
        RECT 128.180 158.545 128.440 159.270 ;
        RECT 128.610 158.715 128.855 159.440 ;
        RECT 129.025 158.545 129.285 159.270 ;
        RECT 129.470 158.715 129.715 159.440 ;
        RECT 129.885 158.545 130.145 159.270 ;
        RECT 130.330 158.715 130.575 159.440 ;
        RECT 130.745 158.545 131.005 159.270 ;
        RECT 131.190 158.715 131.445 159.440 ;
        RECT 125.600 158.530 131.005 158.545 ;
        RECT 131.615 158.530 131.905 159.270 ;
        RECT 132.075 158.700 132.345 159.445 ;
        RECT 125.600 158.305 132.345 158.530 ;
        RECT 116.400 157.545 123.145 157.715 ;
        RECT 123.405 157.575 123.720 158.135 ;
        RECT 123.890 157.885 131.010 158.135 ;
        RECT 115.970 156.895 116.230 157.455 ;
        RECT 116.400 157.090 116.660 157.545 ;
        RECT 116.830 156.895 117.090 157.375 ;
        RECT 117.260 157.090 117.520 157.545 ;
        RECT 117.690 156.895 117.950 157.375 ;
        RECT 118.120 157.090 118.380 157.545 ;
        RECT 118.550 156.895 118.795 157.375 ;
        RECT 118.965 157.090 119.240 157.545 ;
        RECT 119.410 156.895 119.655 157.375 ;
        RECT 119.825 157.090 120.085 157.545 ;
        RECT 120.265 156.895 120.515 157.375 ;
        RECT 120.685 157.090 120.945 157.545 ;
        RECT 121.125 156.895 121.375 157.375 ;
        RECT 121.545 157.090 121.805 157.545 ;
        RECT 121.985 156.895 122.245 157.375 ;
        RECT 122.415 157.090 122.675 157.545 ;
        RECT 122.845 156.895 123.145 157.375 ;
        RECT 123.405 156.895 123.710 157.405 ;
        RECT 123.890 157.075 124.140 157.885 ;
        RECT 124.310 156.895 124.570 157.420 ;
        RECT 124.750 157.075 125.000 157.885 ;
        RECT 131.180 157.715 132.345 158.305 ;
        RECT 132.610 158.475 132.885 159.275 ;
        RECT 133.055 158.645 133.385 159.445 ;
        RECT 133.555 159.105 134.695 159.275 ;
        RECT 133.555 158.475 133.725 159.105 ;
        RECT 132.610 158.265 133.725 158.475 ;
        RECT 133.895 158.475 134.225 158.935 ;
        RECT 134.395 158.645 134.695 159.105 ;
        RECT 133.895 158.255 134.655 158.475 ;
        RECT 132.610 157.885 133.330 158.085 ;
        RECT 133.500 157.885 134.270 158.085 ;
        RECT 134.440 157.715 134.655 158.255 ;
        RECT 134.905 158.355 136.115 159.445 ;
        RECT 134.905 157.815 135.425 158.355 ;
        RECT 125.600 157.545 132.345 157.715 ;
        RECT 125.170 156.895 125.430 157.455 ;
        RECT 125.600 157.090 125.860 157.545 ;
        RECT 126.030 156.895 126.290 157.375 ;
        RECT 126.460 157.090 126.720 157.545 ;
        RECT 126.890 156.895 127.150 157.375 ;
        RECT 127.320 157.090 127.580 157.545 ;
        RECT 127.750 156.895 127.995 157.375 ;
        RECT 128.165 157.090 128.440 157.545 ;
        RECT 128.610 156.895 128.855 157.375 ;
        RECT 129.025 157.090 129.285 157.545 ;
        RECT 129.465 156.895 129.715 157.375 ;
        RECT 129.885 157.090 130.145 157.545 ;
        RECT 130.325 156.895 130.575 157.375 ;
        RECT 130.745 157.090 131.005 157.545 ;
        RECT 131.185 156.895 131.445 157.375 ;
        RECT 131.615 157.090 131.875 157.545 ;
        RECT 132.045 156.895 132.345 157.375 ;
        RECT 132.610 156.895 132.885 157.715 ;
        RECT 133.055 157.545 134.655 157.715 ;
        RECT 135.595 157.645 136.115 158.185 ;
        RECT 133.055 157.535 134.225 157.545 ;
        RECT 133.055 157.065 133.385 157.535 ;
        RECT 133.555 156.895 133.725 157.365 ;
        RECT 133.895 157.065 134.225 157.535 ;
        RECT 134.395 156.895 134.685 157.365 ;
        RECT 134.905 156.895 136.115 157.645 ;
        RECT 23.500 156.725 136.200 156.895 ;
        RECT 23.585 155.975 24.795 156.725 ;
        RECT 25.145 156.065 25.485 156.725 ;
        RECT 23.585 155.435 24.105 155.975 ;
        RECT 24.275 155.265 24.795 155.805 ;
        RECT 23.585 154.175 24.795 155.265 ;
        RECT 24.965 154.345 25.485 155.895 ;
        RECT 25.655 155.070 26.175 156.555 ;
        RECT 26.345 156.180 31.690 156.725 ;
        RECT 31.865 156.180 37.210 156.725 ;
        RECT 37.385 156.180 42.730 156.725 ;
        RECT 42.905 156.180 48.250 156.725 ;
        RECT 27.930 155.350 28.270 156.180 ;
        RECT 25.655 154.175 25.985 154.900 ;
        RECT 29.750 154.610 30.100 155.860 ;
        RECT 33.450 155.350 33.790 156.180 ;
        RECT 35.270 154.610 35.620 155.860 ;
        RECT 38.970 155.350 39.310 156.180 ;
        RECT 40.790 154.610 41.140 155.860 ;
        RECT 44.490 155.350 44.830 156.180 ;
        RECT 49.345 156.000 49.635 156.725 ;
        RECT 50.730 155.885 50.990 156.725 ;
        RECT 51.165 155.980 51.420 156.555 ;
        RECT 51.590 156.345 51.920 156.725 ;
        RECT 52.135 156.175 52.305 156.555 ;
        RECT 51.590 156.005 52.305 156.175 ;
        RECT 52.570 156.155 52.890 156.555 ;
        RECT 46.310 154.610 46.660 155.860 ;
        RECT 26.345 154.175 31.690 154.610 ;
        RECT 31.865 154.175 37.210 154.610 ;
        RECT 37.385 154.175 42.730 154.610 ;
        RECT 42.905 154.175 48.250 154.610 ;
        RECT 49.345 154.175 49.635 155.340 ;
        RECT 50.730 154.175 50.990 155.325 ;
        RECT 51.165 155.250 51.335 155.980 ;
        RECT 51.590 155.815 51.760 156.005 ;
        RECT 51.505 155.485 51.760 155.815 ;
        RECT 51.590 155.275 51.760 155.485 ;
        RECT 52.040 155.455 52.395 155.825 ;
        RECT 52.570 155.365 52.740 156.155 ;
        RECT 53.060 155.905 53.370 156.725 ;
        RECT 53.540 156.095 53.870 156.555 ;
        RECT 54.040 156.265 54.290 156.725 ;
        RECT 54.480 156.345 56.530 156.555 ;
        RECT 54.480 156.095 55.230 156.175 ;
        RECT 53.540 155.905 55.230 156.095 ;
        RECT 55.400 155.905 55.570 156.345 ;
        RECT 55.740 155.905 56.530 156.175 ;
        RECT 56.305 155.875 56.530 155.905 ;
        RECT 56.710 155.885 56.970 156.725 ;
        RECT 57.145 155.980 57.400 156.555 ;
        RECT 57.570 156.345 57.900 156.725 ;
        RECT 58.115 156.175 58.285 156.555 ;
        RECT 57.570 156.005 58.285 156.175 ;
        RECT 52.910 155.535 53.260 155.735 ;
        RECT 53.540 155.535 54.220 155.735 ;
        RECT 54.430 155.535 55.620 155.735 ;
        RECT 55.800 155.365 56.130 155.735 ;
        RECT 51.165 154.345 51.420 155.250 ;
        RECT 51.590 155.105 52.305 155.275 ;
        RECT 51.590 154.175 51.920 154.935 ;
        RECT 52.135 154.345 52.305 155.105 ;
        RECT 52.570 155.195 56.130 155.365 ;
        RECT 52.570 154.745 52.740 155.195 ;
        RECT 56.330 155.025 56.530 155.875 ;
        RECT 52.570 154.345 52.890 154.745 ;
        RECT 53.060 154.175 53.370 154.975 ;
        RECT 53.540 154.855 56.530 155.025 ;
        RECT 53.540 154.805 54.710 154.855 ;
        RECT 53.540 154.345 53.870 154.805 ;
        RECT 54.040 154.175 54.210 154.635 ;
        RECT 54.380 154.345 54.710 154.805 ;
        RECT 55.740 154.805 56.530 154.855 ;
        RECT 54.880 154.175 55.130 154.635 ;
        RECT 55.320 154.175 55.570 154.635 ;
        RECT 55.740 154.345 55.990 154.805 ;
        RECT 56.240 154.175 56.530 154.635 ;
        RECT 56.710 154.175 56.970 155.325 ;
        RECT 57.145 155.250 57.315 155.980 ;
        RECT 57.570 155.815 57.740 156.005 ;
        RECT 58.550 155.885 58.810 156.725 ;
        RECT 58.985 155.980 59.240 156.555 ;
        RECT 59.410 156.345 59.740 156.725 ;
        RECT 59.955 156.175 60.125 156.555 ;
        RECT 59.410 156.005 60.125 156.175 ;
        RECT 57.485 155.485 57.740 155.815 ;
        RECT 57.570 155.275 57.740 155.485 ;
        RECT 58.020 155.455 58.375 155.825 ;
        RECT 57.145 154.345 57.400 155.250 ;
        RECT 57.570 155.105 58.285 155.275 ;
        RECT 57.570 154.175 57.900 154.935 ;
        RECT 58.115 154.345 58.285 155.105 ;
        RECT 58.550 154.175 58.810 155.325 ;
        RECT 58.985 155.250 59.155 155.980 ;
        RECT 59.410 155.815 59.580 156.005 ;
        RECT 60.385 155.985 60.705 156.360 ;
        RECT 60.960 155.985 61.130 156.725 ;
        RECT 61.380 156.155 61.550 156.360 ;
        RECT 61.795 156.325 62.150 156.725 ;
        RECT 62.325 156.155 62.495 156.505 ;
        RECT 62.695 156.325 63.025 156.725 ;
        RECT 63.195 156.155 63.365 156.505 ;
        RECT 63.535 156.325 63.915 156.725 ;
        RECT 61.380 155.985 61.900 156.155 ;
        RECT 62.325 155.985 63.935 156.155 ;
        RECT 64.105 156.050 64.380 156.395 ;
        RECT 59.325 155.485 59.580 155.815 ;
        RECT 59.410 155.275 59.580 155.485 ;
        RECT 59.860 155.455 60.215 155.825 ;
        RECT 58.985 154.345 59.240 155.250 ;
        RECT 59.410 155.105 60.125 155.275 ;
        RECT 59.410 154.175 59.740 154.935 ;
        RECT 59.955 154.345 60.125 155.105 ;
        RECT 60.385 154.945 60.560 155.985 ;
        RECT 60.730 155.115 61.080 155.815 ;
        RECT 61.250 155.485 61.540 155.815 ;
        RECT 61.710 155.735 61.900 155.985 ;
        RECT 63.765 155.815 63.935 155.985 ;
        RECT 61.710 155.565 62.155 155.735 ;
        RECT 61.710 155.285 61.900 155.565 ;
        RECT 62.550 155.395 62.720 155.815 ;
        RECT 62.940 155.485 63.595 155.815 ;
        RECT 63.765 155.485 64.040 155.815 ;
        RECT 61.295 155.115 61.900 155.285 ;
        RECT 62.070 155.225 62.720 155.395 ;
        RECT 63.765 155.315 63.935 155.485 ;
        RECT 64.210 155.315 64.380 156.050 ;
        RECT 64.550 155.785 64.720 156.725 ;
        RECT 64.990 156.345 67.040 156.555 ;
        RECT 64.990 155.905 65.780 156.175 ;
        RECT 65.950 155.905 66.120 156.345 ;
        RECT 67.230 156.265 67.480 156.725 ;
        RECT 66.290 156.095 67.040 156.175 ;
        RECT 67.650 156.095 67.980 156.555 ;
        RECT 66.290 155.905 67.980 156.095 ;
        RECT 68.150 155.905 68.460 156.725 ;
        RECT 68.630 156.155 68.950 156.555 ;
        RECT 64.990 155.875 65.215 155.905 ;
        RECT 62.070 154.945 62.240 155.225 ;
        RECT 63.275 155.145 63.935 155.315 ;
        RECT 63.275 155.025 63.445 155.145 ;
        RECT 60.385 154.775 62.240 154.945 ;
        RECT 62.410 154.855 63.445 155.025 ;
        RECT 60.385 154.355 60.645 154.775 ;
        RECT 62.410 154.605 62.580 154.855 ;
        RECT 60.815 154.175 61.145 154.605 ;
        RECT 61.835 154.435 62.580 154.605 ;
        RECT 62.805 154.355 63.445 154.685 ;
        RECT 63.615 154.175 63.895 154.975 ;
        RECT 64.105 154.345 64.380 155.315 ;
        RECT 64.550 154.175 64.720 155.370 ;
        RECT 64.990 155.025 65.190 155.875 ;
        RECT 65.390 155.365 65.720 155.735 ;
        RECT 65.900 155.535 67.090 155.735 ;
        RECT 67.300 155.535 67.980 155.735 ;
        RECT 68.260 155.535 68.610 155.735 ;
        RECT 68.780 155.365 68.950 156.155 ;
        RECT 69.675 156.175 69.845 156.555 ;
        RECT 70.025 156.345 70.355 156.725 ;
        RECT 69.675 156.005 70.340 156.175 ;
        RECT 70.535 156.050 70.795 156.555 ;
        RECT 69.605 155.455 69.945 155.825 ;
        RECT 70.170 155.750 70.340 156.005 ;
        RECT 65.390 155.195 68.950 155.365 ;
        RECT 70.170 155.420 70.445 155.750 ;
        RECT 70.170 155.275 70.340 155.420 ;
        RECT 64.990 154.855 67.980 155.025 ;
        RECT 64.990 154.805 65.780 154.855 ;
        RECT 64.990 154.175 65.280 154.635 ;
        RECT 65.530 154.345 65.780 154.805 ;
        RECT 66.810 154.805 67.980 154.855 ;
        RECT 65.950 154.175 66.200 154.635 ;
        RECT 66.390 154.175 66.640 154.635 ;
        RECT 66.810 154.345 67.140 154.805 ;
        RECT 67.310 154.175 67.480 154.635 ;
        RECT 67.650 154.345 67.980 154.805 ;
        RECT 68.150 154.175 68.460 154.975 ;
        RECT 68.780 154.745 68.950 155.195 ;
        RECT 68.630 154.345 68.950 154.745 ;
        RECT 69.665 155.105 70.340 155.275 ;
        RECT 70.615 155.250 70.795 156.050 ;
        RECT 71.025 155.905 71.235 156.725 ;
        RECT 71.405 155.925 71.735 156.555 ;
        RECT 71.405 155.325 71.655 155.925 ;
        RECT 71.905 155.905 72.135 156.725 ;
        RECT 72.435 156.175 72.605 156.555 ;
        RECT 72.785 156.345 73.115 156.725 ;
        RECT 72.435 156.005 73.100 156.175 ;
        RECT 73.295 156.050 73.555 156.555 ;
        RECT 71.825 155.485 72.155 155.735 ;
        RECT 72.365 155.455 72.705 155.825 ;
        RECT 72.930 155.750 73.100 156.005 ;
        RECT 72.930 155.420 73.205 155.750 ;
        RECT 69.665 154.345 69.845 155.105 ;
        RECT 70.025 154.175 70.355 154.935 ;
        RECT 70.525 154.345 70.795 155.250 ;
        RECT 71.025 154.175 71.235 155.315 ;
        RECT 71.405 154.345 71.735 155.325 ;
        RECT 71.905 154.175 72.135 155.315 ;
        RECT 72.930 155.275 73.100 155.420 ;
        RECT 72.425 155.105 73.100 155.275 ;
        RECT 73.375 155.250 73.555 156.050 ;
        RECT 73.735 155.915 74.005 156.725 ;
        RECT 74.175 155.915 74.505 156.555 ;
        RECT 74.675 155.915 74.915 156.725 ;
        RECT 75.105 156.000 75.395 156.725 ;
        RECT 75.720 156.075 76.050 156.540 ;
        RECT 76.220 156.255 76.390 156.725 ;
        RECT 76.560 156.075 76.890 156.555 ;
        RECT 73.725 155.485 74.075 155.735 ;
        RECT 74.245 155.315 74.415 155.915 ;
        RECT 75.720 155.905 76.890 156.075 ;
        RECT 74.585 155.485 74.935 155.735 ;
        RECT 75.565 155.525 76.210 155.735 ;
        RECT 76.380 155.525 76.950 155.735 ;
        RECT 77.120 155.355 77.290 156.555 ;
        RECT 77.830 156.155 78.000 156.360 ;
        RECT 72.425 154.345 72.605 155.105 ;
        RECT 72.785 154.175 73.115 154.935 ;
        RECT 73.285 154.345 73.555 155.250 ;
        RECT 73.735 154.175 74.065 155.315 ;
        RECT 74.245 155.145 74.925 155.315 ;
        RECT 74.595 154.360 74.925 155.145 ;
        RECT 75.105 154.175 75.395 155.340 ;
        RECT 75.780 154.175 76.110 155.275 ;
        RECT 76.585 154.945 77.290 155.355 ;
        RECT 77.460 155.985 78.000 156.155 ;
        RECT 78.280 155.985 78.450 156.725 ;
        RECT 78.845 156.360 79.015 156.385 ;
        RECT 78.715 155.985 79.075 156.360 ;
        RECT 77.460 155.285 77.630 155.985 ;
        RECT 77.800 155.485 78.130 155.815 ;
        RECT 78.300 155.485 78.650 155.815 ;
        RECT 77.460 155.115 78.085 155.285 ;
        RECT 78.300 154.945 78.565 155.485 ;
        RECT 78.820 155.330 79.075 155.985 ;
        RECT 80.225 155.905 80.435 156.725 ;
        RECT 80.605 155.925 80.935 156.555 ;
        RECT 76.585 154.775 78.565 154.945 ;
        RECT 76.585 154.345 76.910 154.775 ;
        RECT 77.080 154.175 77.410 154.595 ;
        RECT 78.155 154.175 78.565 154.605 ;
        RECT 78.735 154.345 79.075 155.330 ;
        RECT 80.605 155.325 80.855 155.925 ;
        RECT 81.105 155.905 81.335 156.725 ;
        RECT 81.550 156.050 81.825 156.395 ;
        RECT 82.015 156.325 82.395 156.725 ;
        RECT 82.565 156.155 82.735 156.505 ;
        RECT 82.905 156.325 83.235 156.725 ;
        RECT 83.405 156.155 83.660 156.505 ;
        RECT 81.025 155.485 81.355 155.735 ;
        RECT 80.225 154.175 80.435 155.315 ;
        RECT 80.605 154.345 80.935 155.325 ;
        RECT 81.550 155.315 81.720 156.050 ;
        RECT 81.995 155.985 83.660 156.155 ;
        RECT 81.995 155.815 82.165 155.985 ;
        RECT 83.845 155.925 84.135 156.725 ;
        RECT 84.305 156.265 84.855 156.555 ;
        RECT 85.025 156.265 85.275 156.725 ;
        RECT 81.890 155.485 82.165 155.815 ;
        RECT 82.335 155.485 83.160 155.815 ;
        RECT 83.330 155.485 83.675 155.815 ;
        RECT 81.995 155.315 82.165 155.485 ;
        RECT 81.105 154.175 81.335 155.315 ;
        RECT 81.550 154.345 81.825 155.315 ;
        RECT 81.995 155.145 82.655 155.315 ;
        RECT 82.965 155.195 83.160 155.485 ;
        RECT 82.485 155.025 82.655 155.145 ;
        RECT 83.330 155.025 83.655 155.315 ;
        RECT 82.035 154.175 82.315 154.975 ;
        RECT 82.485 154.855 83.655 155.025 ;
        RECT 82.485 154.395 83.675 154.685 ;
        RECT 83.845 154.175 84.135 155.315 ;
        RECT 84.305 154.895 84.555 156.265 ;
        RECT 85.905 156.095 86.235 156.455 ;
        RECT 84.845 155.905 86.235 156.095 ;
        RECT 86.625 156.185 86.955 156.555 ;
        RECT 87.125 156.355 87.455 156.725 ;
        RECT 87.645 156.185 87.990 156.555 ;
        RECT 86.625 155.985 87.990 156.185 ;
        RECT 84.845 155.815 85.015 155.905 ;
        RECT 84.725 155.485 85.015 155.815 ;
        RECT 85.185 155.485 85.515 155.735 ;
        RECT 85.745 155.485 86.435 155.735 ;
        RECT 84.845 155.235 85.015 155.485 ;
        RECT 84.845 155.065 85.785 155.235 ;
        RECT 84.305 154.345 84.755 154.895 ;
        RECT 84.945 154.175 85.275 154.895 ;
        RECT 85.485 154.515 85.785 155.065 ;
        RECT 86.120 155.045 86.435 155.485 ;
        RECT 86.625 155.195 86.955 155.805 ;
        RECT 87.125 155.195 87.755 155.815 ;
        RECT 87.925 155.195 88.215 155.815 ;
        RECT 88.385 155.195 88.715 156.555 ;
        RECT 89.050 155.925 89.655 156.555 ;
        RECT 89.915 156.175 90.085 156.555 ;
        RECT 90.300 156.345 90.630 156.725 ;
        RECT 89.915 156.005 90.630 156.175 ;
        RECT 88.925 155.195 89.255 155.735 ;
        RECT 85.955 154.175 86.235 154.845 ;
        RECT 86.625 154.175 86.955 155.015 ;
        RECT 87.125 154.440 87.470 155.195 ;
        RECT 89.425 155.025 89.655 155.925 ;
        RECT 89.825 155.455 90.180 155.825 ;
        RECT 90.460 155.815 90.630 156.005 ;
        RECT 90.800 155.980 91.055 156.555 ;
        RECT 90.460 155.485 90.715 155.815 ;
        RECT 90.460 155.275 90.630 155.485 ;
        RECT 87.645 154.785 89.655 155.025 ;
        RECT 89.915 155.105 90.630 155.275 ;
        RECT 90.885 155.250 91.055 155.980 ;
        RECT 91.230 155.885 91.490 156.725 ;
        RECT 91.755 156.245 92.055 156.725 ;
        RECT 92.225 156.075 92.485 156.530 ;
        RECT 92.655 156.245 92.915 156.725 ;
        RECT 93.095 156.075 93.355 156.530 ;
        RECT 93.525 156.245 93.775 156.725 ;
        RECT 93.955 156.075 94.215 156.530 ;
        RECT 94.385 156.245 94.635 156.725 ;
        RECT 94.815 156.075 95.075 156.530 ;
        RECT 95.245 156.245 95.490 156.725 ;
        RECT 95.660 156.075 95.935 156.530 ;
        RECT 96.105 156.245 96.350 156.725 ;
        RECT 96.520 156.075 96.780 156.530 ;
        RECT 96.950 156.245 97.210 156.725 ;
        RECT 97.380 156.075 97.640 156.530 ;
        RECT 97.810 156.245 98.070 156.725 ;
        RECT 98.240 156.075 98.500 156.530 ;
        RECT 98.670 156.165 98.930 156.725 ;
        RECT 91.755 155.905 98.500 156.075 ;
        RECT 87.645 154.345 87.990 154.785 ;
        RECT 88.200 154.175 88.530 154.555 ;
        RECT 88.715 154.345 88.950 154.785 ;
        RECT 89.120 154.175 89.450 154.615 ;
        RECT 89.915 154.345 90.085 155.105 ;
        RECT 90.300 154.175 90.630 154.935 ;
        RECT 90.800 154.345 91.055 155.250 ;
        RECT 91.230 154.175 91.490 155.325 ;
        RECT 91.755 155.315 92.920 155.905 ;
        RECT 99.100 155.735 99.350 156.545 ;
        RECT 99.530 156.200 99.790 156.725 ;
        RECT 99.960 155.735 100.210 156.545 ;
        RECT 100.390 156.215 100.695 156.725 ;
        RECT 93.090 155.485 100.210 155.735 ;
        RECT 100.380 155.485 100.695 156.045 ;
        RECT 100.865 156.000 101.155 156.725 ;
        RECT 101.330 155.905 101.605 156.725 ;
        RECT 101.775 156.085 102.105 156.555 ;
        RECT 102.275 156.255 102.445 156.725 ;
        RECT 102.615 156.085 102.945 156.555 ;
        RECT 103.115 156.255 103.825 156.725 ;
        RECT 103.995 156.085 104.325 156.555 ;
        RECT 104.495 156.255 104.785 156.725 ;
        RECT 105.555 156.245 105.855 156.725 ;
        RECT 101.775 155.905 104.835 156.085 ;
        RECT 106.025 156.075 106.285 156.530 ;
        RECT 106.455 156.245 106.715 156.725 ;
        RECT 106.895 156.075 107.155 156.530 ;
        RECT 107.325 156.245 107.575 156.725 ;
        RECT 107.755 156.075 108.015 156.530 ;
        RECT 108.185 156.245 108.435 156.725 ;
        RECT 108.615 156.075 108.875 156.530 ;
        RECT 109.045 156.245 109.290 156.725 ;
        RECT 109.460 156.075 109.735 156.530 ;
        RECT 109.905 156.245 110.150 156.725 ;
        RECT 110.320 156.075 110.580 156.530 ;
        RECT 110.750 156.245 111.010 156.725 ;
        RECT 111.180 156.075 111.440 156.530 ;
        RECT 111.610 156.245 111.870 156.725 ;
        RECT 112.040 156.075 112.300 156.530 ;
        RECT 112.470 156.165 112.730 156.725 ;
        RECT 101.375 155.525 102.205 155.735 ;
        RECT 102.375 155.525 103.425 155.735 ;
        RECT 103.615 155.525 104.205 155.735 ;
        RECT 91.755 155.090 98.500 155.315 ;
        RECT 91.755 154.175 92.025 154.920 ;
        RECT 92.195 154.350 92.485 155.090 ;
        RECT 93.095 155.075 98.500 155.090 ;
        RECT 92.655 154.180 92.910 154.905 ;
        RECT 93.095 154.350 93.355 155.075 ;
        RECT 93.525 154.180 93.770 154.905 ;
        RECT 93.955 154.350 94.215 155.075 ;
        RECT 94.385 154.180 94.630 154.905 ;
        RECT 94.815 154.350 95.075 155.075 ;
        RECT 95.245 154.180 95.490 154.905 ;
        RECT 95.660 154.350 95.920 155.075 ;
        RECT 96.090 154.180 96.350 154.905 ;
        RECT 96.520 154.350 96.780 155.075 ;
        RECT 96.950 154.180 97.210 154.905 ;
        RECT 97.380 154.350 97.640 155.075 ;
        RECT 97.810 154.180 98.070 154.905 ;
        RECT 98.240 154.350 98.500 155.075 ;
        RECT 98.670 154.180 98.930 154.975 ;
        RECT 99.100 154.350 99.350 155.485 ;
        RECT 92.655 154.175 98.930 154.180 ;
        RECT 99.530 154.175 99.790 154.985 ;
        RECT 99.965 154.345 100.210 155.485 ;
        RECT 100.390 154.175 100.685 154.985 ;
        RECT 100.865 154.175 101.155 155.340 ;
        RECT 101.390 155.185 103.325 155.355 ;
        RECT 103.615 155.185 103.880 155.525 ;
        RECT 104.375 155.355 104.835 155.905 ;
        RECT 104.075 155.185 104.835 155.355 ;
        RECT 105.555 155.905 112.300 156.075 ;
        RECT 105.555 155.315 106.720 155.905 ;
        RECT 112.900 155.735 113.150 156.545 ;
        RECT 113.330 156.200 113.590 156.725 ;
        RECT 113.760 155.735 114.010 156.545 ;
        RECT 114.190 156.215 114.495 156.725 ;
        RECT 114.685 156.240 115.475 156.505 ;
        RECT 106.890 155.485 114.010 155.735 ;
        RECT 114.180 155.485 114.495 156.045 ;
        RECT 114.665 155.565 115.050 156.045 ;
        RECT 101.390 154.345 101.645 155.185 ;
        RECT 101.815 154.175 102.065 155.015 ;
        RECT 102.235 154.345 102.485 155.185 ;
        RECT 102.655 154.515 102.905 155.015 ;
        RECT 103.075 154.685 103.325 155.185 ;
        RECT 103.655 154.515 103.865 155.015 ;
        RECT 104.075 154.685 104.285 155.185 ;
        RECT 105.555 155.090 112.300 155.315 ;
        RECT 104.455 154.515 104.705 155.015 ;
        RECT 102.655 154.345 104.705 154.515 ;
        RECT 105.555 154.175 105.825 154.920 ;
        RECT 105.995 154.350 106.285 155.090 ;
        RECT 106.895 155.075 112.300 155.090 ;
        RECT 106.455 154.180 106.710 154.905 ;
        RECT 106.895 154.350 107.155 155.075 ;
        RECT 107.325 154.180 107.570 154.905 ;
        RECT 107.755 154.350 108.015 155.075 ;
        RECT 108.185 154.180 108.430 154.905 ;
        RECT 108.615 154.350 108.875 155.075 ;
        RECT 109.045 154.180 109.290 154.905 ;
        RECT 109.460 154.350 109.720 155.075 ;
        RECT 109.890 154.180 110.150 154.905 ;
        RECT 110.320 154.350 110.580 155.075 ;
        RECT 110.750 154.180 111.010 154.905 ;
        RECT 111.180 154.350 111.440 155.075 ;
        RECT 111.610 154.180 111.870 154.905 ;
        RECT 112.040 154.350 112.300 155.075 ;
        RECT 112.470 154.180 112.730 154.975 ;
        RECT 112.900 154.350 113.150 155.485 ;
        RECT 106.455 154.175 112.730 154.180 ;
        RECT 113.330 154.175 113.590 154.985 ;
        RECT 113.765 154.345 114.010 155.485 ;
        RECT 115.220 155.385 115.475 156.240 ;
        RECT 115.645 156.060 115.875 156.505 ;
        RECT 116.055 156.230 116.385 156.725 ;
        RECT 116.560 156.095 116.810 156.555 ;
        RECT 115.645 155.565 116.055 156.060 ;
        RECT 116.640 155.885 116.810 156.095 ;
        RECT 116.980 156.065 117.255 156.725 ;
        RECT 117.425 156.215 117.730 156.725 ;
        RECT 116.240 155.385 116.470 155.815 ;
        RECT 114.680 155.215 116.470 155.385 ;
        RECT 116.640 155.365 117.255 155.885 ;
        RECT 117.425 155.485 117.740 156.045 ;
        RECT 117.910 155.735 118.160 156.545 ;
        RECT 118.330 156.200 118.590 156.725 ;
        RECT 118.770 155.735 119.020 156.545 ;
        RECT 119.190 156.165 119.450 156.725 ;
        RECT 119.620 156.075 119.880 156.530 ;
        RECT 120.050 156.245 120.310 156.725 ;
        RECT 120.480 156.075 120.740 156.530 ;
        RECT 120.910 156.245 121.170 156.725 ;
        RECT 121.340 156.075 121.600 156.530 ;
        RECT 121.770 156.245 122.015 156.725 ;
        RECT 122.185 156.075 122.460 156.530 ;
        RECT 122.630 156.245 122.875 156.725 ;
        RECT 123.045 156.075 123.305 156.530 ;
        RECT 123.485 156.245 123.735 156.725 ;
        RECT 123.905 156.075 124.165 156.530 ;
        RECT 124.345 156.245 124.595 156.725 ;
        RECT 124.765 156.075 125.025 156.530 ;
        RECT 125.205 156.245 125.465 156.725 ;
        RECT 125.635 156.075 125.895 156.530 ;
        RECT 126.065 156.245 126.365 156.725 ;
        RECT 119.620 156.045 126.365 156.075 ;
        RECT 119.620 155.905 126.395 156.045 ;
        RECT 126.625 156.000 126.915 156.725 ;
        RECT 127.100 155.945 127.395 156.725 ;
        RECT 127.955 156.195 128.300 156.555 ;
        RECT 128.760 156.365 129.090 156.725 ;
        RECT 129.295 156.195 129.615 156.555 ;
        RECT 127.955 156.025 129.615 156.195 ;
        RECT 125.200 155.875 126.395 155.905 ;
        RECT 117.910 155.485 125.030 155.735 ;
        RECT 114.190 154.175 114.485 154.985 ;
        RECT 114.680 154.850 114.935 155.215 ;
        RECT 115.105 154.855 115.435 155.045 ;
        RECT 115.660 154.920 115.910 155.215 ;
        RECT 115.105 154.680 115.295 154.855 ;
        RECT 114.665 154.175 115.295 154.680 ;
        RECT 115.475 154.345 115.950 154.685 ;
        RECT 116.135 154.175 116.350 155.020 ;
        RECT 116.655 155.015 116.825 155.365 ;
        RECT 116.550 154.345 116.825 155.015 ;
        RECT 116.995 154.175 117.255 155.185 ;
        RECT 117.435 154.175 117.730 154.985 ;
        RECT 117.910 154.345 118.155 155.485 ;
        RECT 118.330 154.175 118.590 154.985 ;
        RECT 118.770 154.350 119.020 155.485 ;
        RECT 125.200 155.315 126.365 155.875 ;
        RECT 119.620 155.090 126.365 155.315 ;
        RECT 119.620 155.075 125.025 155.090 ;
        RECT 119.190 154.180 119.450 154.975 ;
        RECT 119.620 154.350 119.880 155.075 ;
        RECT 120.050 154.180 120.310 154.905 ;
        RECT 120.480 154.350 120.740 155.075 ;
        RECT 120.910 154.180 121.170 154.905 ;
        RECT 121.340 154.350 121.600 155.075 ;
        RECT 121.770 154.180 122.030 154.905 ;
        RECT 122.200 154.350 122.460 155.075 ;
        RECT 122.630 154.180 122.875 154.905 ;
        RECT 123.045 154.350 123.305 155.075 ;
        RECT 123.490 154.180 123.735 154.905 ;
        RECT 123.905 154.350 124.165 155.075 ;
        RECT 124.350 154.180 124.595 154.905 ;
        RECT 124.765 154.350 125.025 155.075 ;
        RECT 125.210 154.180 125.465 154.905 ;
        RECT 125.635 154.350 125.925 155.090 ;
        RECT 119.190 154.175 125.465 154.180 ;
        RECT 126.095 154.175 126.365 154.920 ;
        RECT 126.625 154.175 126.915 155.340 ;
        RECT 127.145 155.315 127.645 155.775 ;
        RECT 127.815 155.485 128.425 155.815 ;
        RECT 128.605 155.565 128.935 155.735 ;
        RECT 128.605 155.315 128.930 155.565 ;
        RECT 127.145 155.135 128.930 155.315 ;
        RECT 127.110 154.785 129.145 154.955 ;
        RECT 127.110 154.705 128.220 154.785 ;
        RECT 127.110 154.345 127.370 154.705 ;
        RECT 127.540 154.175 127.870 154.535 ;
        RECT 128.050 154.345 128.220 154.705 ;
        RECT 128.475 154.175 128.645 154.615 ;
        RECT 128.815 154.525 129.145 154.785 ;
        RECT 129.315 154.695 129.615 156.025 ;
        RECT 129.795 155.985 130.125 156.725 ;
        RECT 130.920 156.075 131.250 156.540 ;
        RECT 131.420 156.255 131.590 156.725 ;
        RECT 131.760 156.075 132.090 156.555 ;
        RECT 130.920 155.905 132.090 156.075 ;
        RECT 129.800 155.185 130.075 155.815 ;
        RECT 130.765 155.525 131.410 155.735 ;
        RECT 131.580 155.525 132.150 155.735 ;
        RECT 132.320 155.355 132.490 156.555 ;
        RECT 133.030 156.155 133.200 156.360 ;
        RECT 129.785 154.525 130.090 155.015 ;
        RECT 128.815 154.345 130.090 154.525 ;
        RECT 130.980 154.175 131.310 155.275 ;
        RECT 131.785 154.945 132.490 155.355 ;
        RECT 132.660 155.985 133.200 156.155 ;
        RECT 133.480 155.985 133.650 156.725 ;
        RECT 134.045 156.360 134.215 156.385 ;
        RECT 133.915 155.985 134.275 156.360 ;
        RECT 132.660 155.285 132.830 155.985 ;
        RECT 133.000 155.485 133.330 155.815 ;
        RECT 133.500 155.485 133.850 155.815 ;
        RECT 132.660 155.115 133.285 155.285 ;
        RECT 133.500 154.945 133.765 155.485 ;
        RECT 134.020 155.330 134.275 155.985 ;
        RECT 134.905 155.975 136.115 156.725 ;
        RECT 131.785 154.775 133.765 154.945 ;
        RECT 131.785 154.345 132.110 154.775 ;
        RECT 132.280 154.175 132.610 154.595 ;
        RECT 133.355 154.175 133.765 154.605 ;
        RECT 133.935 154.345 134.275 155.330 ;
        RECT 134.905 155.265 135.425 155.805 ;
        RECT 135.595 155.435 136.115 155.975 ;
        RECT 134.905 154.175 136.115 155.265 ;
        RECT 23.500 154.005 136.200 154.175 ;
        RECT 23.585 152.915 24.795 154.005 ;
        RECT 24.965 153.570 30.310 154.005 ;
        RECT 30.485 153.570 35.830 154.005 ;
        RECT 23.585 152.205 24.105 152.745 ;
        RECT 24.275 152.375 24.795 152.915 ;
        RECT 23.585 151.455 24.795 152.205 ;
        RECT 26.550 152.000 26.890 152.830 ;
        RECT 28.370 152.320 28.720 153.570 ;
        RECT 32.070 152.000 32.410 152.830 ;
        RECT 33.890 152.320 34.240 153.570 ;
        RECT 36.465 152.840 36.755 154.005 ;
        RECT 37.925 153.075 38.105 153.835 ;
        RECT 38.285 153.245 38.615 154.005 ;
        RECT 37.925 152.905 38.600 153.075 ;
        RECT 38.785 152.930 39.055 153.835 ;
        RECT 38.430 152.760 38.600 152.905 ;
        RECT 37.865 152.355 38.205 152.725 ;
        RECT 38.430 152.430 38.705 152.760 ;
        RECT 24.965 151.455 30.310 152.000 ;
        RECT 30.485 151.455 35.830 152.000 ;
        RECT 36.465 151.455 36.755 152.180 ;
        RECT 38.430 152.175 38.600 152.430 ;
        RECT 37.935 152.005 38.600 152.175 ;
        RECT 38.875 152.130 39.055 152.930 ;
        RECT 39.225 152.915 40.895 154.005 ;
        RECT 37.935 151.625 38.105 152.005 ;
        RECT 38.285 151.455 38.615 151.835 ;
        RECT 38.795 151.625 39.055 152.130 ;
        RECT 39.225 152.225 39.975 152.745 ;
        RECT 40.145 152.395 40.895 152.915 ;
        RECT 41.155 153.075 41.325 153.835 ;
        RECT 41.505 153.245 41.835 154.005 ;
        RECT 41.155 152.905 41.820 153.075 ;
        RECT 42.005 152.930 42.275 153.835 ;
        RECT 41.650 152.760 41.820 152.905 ;
        RECT 41.085 152.355 41.415 152.725 ;
        RECT 41.650 152.430 41.935 152.760 ;
        RECT 39.225 151.455 40.895 152.225 ;
        RECT 41.650 152.175 41.820 152.430 ;
        RECT 41.155 152.005 41.820 152.175 ;
        RECT 42.105 152.130 42.275 152.930 ;
        RECT 42.445 152.915 44.115 154.005 ;
        RECT 41.155 151.625 41.325 152.005 ;
        RECT 41.505 151.455 41.835 151.835 ;
        RECT 42.015 151.625 42.275 152.130 ;
        RECT 42.445 152.225 43.195 152.745 ;
        RECT 43.365 152.395 44.115 152.915 ;
        RECT 44.375 153.075 44.545 153.835 ;
        RECT 44.760 153.245 45.090 154.005 ;
        RECT 44.375 152.905 45.090 153.075 ;
        RECT 45.260 152.930 45.515 153.835 ;
        RECT 44.285 152.355 44.640 152.725 ;
        RECT 44.920 152.695 45.090 152.905 ;
        RECT 44.920 152.365 45.175 152.695 ;
        RECT 42.445 151.455 44.115 152.225 ;
        RECT 44.920 152.175 45.090 152.365 ;
        RECT 45.345 152.200 45.515 152.930 ;
        RECT 45.690 152.855 45.950 154.005 ;
        RECT 46.125 152.915 47.335 154.005 ;
        RECT 44.375 152.005 45.090 152.175 ;
        RECT 44.375 151.625 44.545 152.005 ;
        RECT 44.760 151.455 45.090 151.835 ;
        RECT 45.260 151.625 45.515 152.200 ;
        RECT 45.690 151.455 45.950 152.295 ;
        RECT 46.125 152.205 46.645 152.745 ;
        RECT 46.815 152.375 47.335 152.915 ;
        RECT 47.585 153.075 47.765 153.835 ;
        RECT 47.945 153.245 48.275 154.005 ;
        RECT 47.585 152.905 48.260 153.075 ;
        RECT 48.445 152.930 48.715 153.835 ;
        RECT 48.090 152.760 48.260 152.905 ;
        RECT 47.525 152.355 47.865 152.725 ;
        RECT 48.090 152.430 48.365 152.760 ;
        RECT 46.125 151.455 47.335 152.205 ;
        RECT 48.090 152.175 48.260 152.430 ;
        RECT 47.595 152.005 48.260 152.175 ;
        RECT 48.535 152.130 48.715 152.930 ;
        RECT 49.345 152.840 49.635 154.005 ;
        RECT 49.805 152.915 51.475 154.005 ;
        RECT 49.805 152.225 50.555 152.745 ;
        RECT 50.725 152.395 51.475 152.915 ;
        RECT 51.645 153.405 51.905 153.825 ;
        RECT 52.075 153.575 52.405 154.005 ;
        RECT 53.070 153.575 53.815 153.745 ;
        RECT 51.645 153.235 53.475 153.405 ;
        RECT 47.595 151.625 47.765 152.005 ;
        RECT 47.945 151.455 48.275 151.835 ;
        RECT 48.455 151.625 48.715 152.130 ;
        RECT 49.345 151.455 49.635 152.180 ;
        RECT 49.805 151.455 51.475 152.225 ;
        RECT 51.645 152.195 51.815 153.235 ;
        RECT 51.985 152.365 52.335 153.065 ;
        RECT 52.550 152.895 53.135 153.065 ;
        RECT 52.505 152.365 52.795 152.695 ;
        RECT 52.965 152.615 53.135 152.895 ;
        RECT 53.305 152.955 53.475 153.235 ;
        RECT 53.645 153.325 53.815 153.575 ;
        RECT 54.040 153.495 54.680 153.825 ;
        RECT 53.645 153.155 54.680 153.325 ;
        RECT 54.850 153.205 55.130 154.005 ;
        RECT 54.510 153.035 54.680 153.155 ;
        RECT 53.305 152.785 53.955 152.955 ;
        RECT 54.510 152.865 55.170 153.035 ;
        RECT 55.340 152.865 55.615 153.835 ;
        RECT 52.965 152.445 53.390 152.615 ;
        RECT 52.965 152.195 53.135 152.445 ;
        RECT 53.785 152.365 53.955 152.785 ;
        RECT 55.000 152.695 55.170 152.865 ;
        RECT 54.175 152.365 54.830 152.695 ;
        RECT 55.000 152.365 55.275 152.695 ;
        RECT 55.000 152.195 55.170 152.365 ;
        RECT 51.645 151.820 51.960 152.195 ;
        RECT 52.215 151.455 52.385 152.195 ;
        RECT 52.635 152.025 53.135 152.195 ;
        RECT 53.575 152.025 55.170 152.195 ;
        RECT 55.445 152.130 55.615 152.865 ;
        RECT 52.635 151.820 52.805 152.025 ;
        RECT 53.030 151.455 53.405 151.855 ;
        RECT 53.575 151.675 53.745 152.025 ;
        RECT 53.930 151.455 54.260 151.855 ;
        RECT 54.430 151.675 54.600 152.025 ;
        RECT 54.770 151.455 55.150 151.855 ;
        RECT 55.340 151.785 55.615 152.130 ;
        RECT 55.785 153.035 56.055 153.805 ;
        RECT 56.225 153.225 56.555 154.005 ;
        RECT 56.760 153.400 56.945 153.805 ;
        RECT 57.115 153.580 57.450 154.005 ;
        RECT 56.760 153.225 57.425 153.400 ;
        RECT 55.785 152.865 56.915 153.035 ;
        RECT 55.785 151.955 55.955 152.865 ;
        RECT 56.125 152.115 56.485 152.695 ;
        RECT 56.665 152.365 56.915 152.865 ;
        RECT 57.085 152.195 57.425 153.225 ;
        RECT 57.705 153.075 57.885 153.835 ;
        RECT 58.065 153.245 58.395 154.005 ;
        RECT 57.705 152.905 58.380 153.075 ;
        RECT 58.565 152.930 58.835 153.835 ;
        RECT 58.210 152.760 58.380 152.905 ;
        RECT 57.645 152.355 57.985 152.725 ;
        RECT 58.210 152.430 58.485 152.760 ;
        RECT 56.740 152.025 57.425 152.195 ;
        RECT 58.210 152.175 58.380 152.430 ;
        RECT 55.785 151.625 56.045 151.955 ;
        RECT 56.255 151.455 56.530 151.935 ;
        RECT 56.740 151.625 56.945 152.025 ;
        RECT 57.715 152.005 58.380 152.175 ;
        RECT 58.655 152.130 58.835 152.930 ;
        RECT 57.115 151.455 57.450 151.855 ;
        RECT 57.715 151.625 57.885 152.005 ;
        RECT 58.065 151.455 58.395 151.835 ;
        RECT 58.575 151.625 58.835 152.130 ;
        RECT 59.925 151.625 60.675 153.835 ;
        RECT 60.925 153.075 61.105 153.835 ;
        RECT 61.285 153.245 61.615 154.005 ;
        RECT 60.925 152.905 61.600 153.075 ;
        RECT 61.785 152.930 62.055 153.835 ;
        RECT 61.430 152.760 61.600 152.905 ;
        RECT 60.865 152.355 61.205 152.725 ;
        RECT 61.430 152.430 61.705 152.760 ;
        RECT 61.430 152.175 61.600 152.430 ;
        RECT 60.935 152.005 61.600 152.175 ;
        RECT 61.875 152.130 62.055 152.930 ;
        RECT 62.225 152.840 62.515 154.005 ;
        RECT 63.695 153.075 63.865 153.835 ;
        RECT 64.080 153.245 64.410 154.005 ;
        RECT 63.695 152.905 64.410 153.075 ;
        RECT 64.580 152.930 64.835 153.835 ;
        RECT 63.605 152.355 63.960 152.725 ;
        RECT 64.240 152.695 64.410 152.905 ;
        RECT 64.240 152.365 64.495 152.695 ;
        RECT 60.935 151.625 61.105 152.005 ;
        RECT 61.285 151.455 61.615 151.835 ;
        RECT 61.795 151.625 62.055 152.130 ;
        RECT 62.225 151.455 62.515 152.180 ;
        RECT 64.240 152.175 64.410 152.365 ;
        RECT 64.665 152.200 64.835 152.930 ;
        RECT 65.010 152.855 65.270 154.005 ;
        RECT 65.525 153.075 65.705 153.835 ;
        RECT 65.885 153.245 66.215 154.005 ;
        RECT 65.525 152.905 66.200 153.075 ;
        RECT 66.385 152.930 66.655 153.835 ;
        RECT 66.030 152.760 66.200 152.905 ;
        RECT 65.465 152.355 65.805 152.725 ;
        RECT 66.030 152.430 66.305 152.760 ;
        RECT 63.695 152.005 64.410 152.175 ;
        RECT 63.695 151.625 63.865 152.005 ;
        RECT 64.080 151.455 64.410 151.835 ;
        RECT 64.580 151.625 64.835 152.200 ;
        RECT 65.010 151.455 65.270 152.295 ;
        RECT 66.030 152.175 66.200 152.430 ;
        RECT 65.535 152.005 66.200 152.175 ;
        RECT 66.475 152.130 66.655 152.930 ;
        RECT 66.825 152.285 67.345 153.835 ;
        RECT 67.515 153.280 67.845 154.005 ;
        RECT 65.535 151.625 65.705 152.005 ;
        RECT 65.885 151.455 66.215 151.835 ;
        RECT 66.395 151.625 66.655 152.130 ;
        RECT 67.005 151.455 67.345 152.115 ;
        RECT 67.515 151.625 68.035 153.110 ;
        RECT 68.285 153.075 68.465 153.835 ;
        RECT 68.645 153.245 68.975 154.005 ;
        RECT 68.285 152.905 68.960 153.075 ;
        RECT 69.145 152.930 69.415 153.835 ;
        RECT 68.790 152.760 68.960 152.905 ;
        RECT 68.225 152.355 68.565 152.725 ;
        RECT 68.790 152.430 69.065 152.760 ;
        RECT 68.790 152.175 68.960 152.430 ;
        RECT 68.295 152.005 68.960 152.175 ;
        RECT 69.235 152.130 69.415 152.930 ;
        RECT 69.735 152.855 70.065 154.005 ;
        RECT 70.235 152.985 70.405 153.835 ;
        RECT 70.575 153.205 70.905 154.005 ;
        RECT 71.075 152.985 71.245 153.835 ;
        RECT 71.425 153.205 71.665 154.005 ;
        RECT 71.835 153.025 72.165 153.835 ;
        RECT 70.235 152.815 71.245 152.985 ;
        RECT 71.450 152.855 72.165 153.025 ;
        RECT 72.425 153.075 72.605 153.835 ;
        RECT 72.785 153.245 73.115 154.005 ;
        RECT 72.425 152.905 73.100 153.075 ;
        RECT 73.285 152.930 73.555 153.835 ;
        RECT 70.235 152.305 70.730 152.815 ;
        RECT 71.450 152.615 71.620 152.855 ;
        RECT 72.930 152.760 73.100 152.905 ;
        RECT 71.120 152.445 71.620 152.615 ;
        RECT 71.790 152.445 72.170 152.685 ;
        RECT 70.235 152.275 70.735 152.305 ;
        RECT 71.450 152.275 71.620 152.445 ;
        RECT 72.365 152.355 72.705 152.725 ;
        RECT 72.930 152.430 73.205 152.760 ;
        RECT 68.295 151.625 68.465 152.005 ;
        RECT 68.645 151.455 68.975 151.835 ;
        RECT 69.155 151.625 69.415 152.130 ;
        RECT 69.735 151.455 70.065 152.255 ;
        RECT 70.235 152.105 71.245 152.275 ;
        RECT 71.450 152.105 72.085 152.275 ;
        RECT 72.930 152.175 73.100 152.430 ;
        RECT 70.235 151.625 70.405 152.105 ;
        RECT 70.575 151.455 70.905 151.935 ;
        RECT 71.075 151.625 71.245 152.105 ;
        RECT 71.495 151.455 71.735 151.935 ;
        RECT 71.915 151.625 72.085 152.105 ;
        RECT 72.435 152.005 73.100 152.175 ;
        RECT 73.375 152.130 73.555 152.930 ;
        RECT 73.805 153.075 73.985 153.835 ;
        RECT 74.165 153.245 74.495 154.005 ;
        RECT 73.805 152.905 74.480 153.075 ;
        RECT 74.665 152.930 74.935 153.835 ;
        RECT 74.310 152.760 74.480 152.905 ;
        RECT 73.745 152.355 74.085 152.725 ;
        RECT 74.310 152.430 74.585 152.760 ;
        RECT 74.310 152.175 74.480 152.430 ;
        RECT 72.435 151.625 72.605 152.005 ;
        RECT 72.785 151.455 73.115 151.835 ;
        RECT 73.295 151.625 73.555 152.130 ;
        RECT 73.815 152.005 74.480 152.175 ;
        RECT 74.755 152.130 74.935 152.930 ;
        RECT 75.105 152.840 75.395 154.005 ;
        RECT 76.565 153.075 76.745 153.835 ;
        RECT 76.925 153.245 77.255 154.005 ;
        RECT 76.565 152.905 77.240 153.075 ;
        RECT 77.425 152.930 77.695 153.835 ;
        RECT 77.070 152.760 77.240 152.905 ;
        RECT 76.505 152.355 76.845 152.725 ;
        RECT 77.070 152.430 77.345 152.760 ;
        RECT 73.815 151.625 73.985 152.005 ;
        RECT 74.165 151.455 74.495 151.835 ;
        RECT 74.675 151.625 74.935 152.130 ;
        RECT 75.105 151.455 75.395 152.180 ;
        RECT 77.070 152.175 77.240 152.430 ;
        RECT 76.575 152.005 77.240 152.175 ;
        RECT 77.515 152.130 77.695 152.930 ;
        RECT 77.945 153.075 78.125 153.835 ;
        RECT 78.305 153.245 78.635 154.005 ;
        RECT 77.945 152.905 78.620 153.075 ;
        RECT 78.805 152.930 79.075 153.835 ;
        RECT 78.450 152.760 78.620 152.905 ;
        RECT 77.885 152.355 78.225 152.725 ;
        RECT 78.450 152.430 78.725 152.760 ;
        RECT 78.450 152.175 78.620 152.430 ;
        RECT 76.575 151.625 76.745 152.005 ;
        RECT 76.925 151.455 77.255 151.835 ;
        RECT 77.435 151.625 77.695 152.130 ;
        RECT 77.955 152.005 78.620 152.175 ;
        RECT 78.895 152.130 79.075 152.930 ;
        RECT 79.255 152.865 79.585 154.005 ;
        RECT 80.115 153.035 80.445 153.820 ;
        RECT 79.765 152.865 80.445 153.035 ;
        RECT 79.245 152.445 79.595 152.695 ;
        RECT 79.765 152.265 79.935 152.865 ;
        RECT 81.090 152.855 81.350 154.005 ;
        RECT 81.525 152.930 81.780 153.835 ;
        RECT 81.950 153.245 82.280 154.005 ;
        RECT 82.495 153.075 82.665 153.835 ;
        RECT 82.965 153.665 84.105 153.835 ;
        RECT 82.965 153.205 83.265 153.665 ;
        RECT 80.105 152.445 80.455 152.695 ;
        RECT 77.955 151.625 78.125 152.005 ;
        RECT 78.305 151.455 78.635 151.835 ;
        RECT 78.815 151.625 79.075 152.130 ;
        RECT 79.255 151.455 79.525 152.265 ;
        RECT 79.695 151.625 80.025 152.265 ;
        RECT 80.195 151.455 80.435 152.265 ;
        RECT 81.090 151.455 81.350 152.295 ;
        RECT 81.525 152.200 81.695 152.930 ;
        RECT 81.950 152.905 82.665 153.075 ;
        RECT 83.435 153.035 83.765 153.495 ;
        RECT 81.950 152.695 82.120 152.905 ;
        RECT 83.005 152.815 83.765 153.035 ;
        RECT 83.935 153.035 84.105 153.665 ;
        RECT 84.275 153.205 84.605 154.005 ;
        RECT 84.775 153.035 85.050 153.835 ;
        RECT 85.280 153.135 85.565 154.005 ;
        RECT 85.735 153.375 85.995 153.835 ;
        RECT 86.170 153.545 86.425 154.005 ;
        RECT 86.595 153.375 86.855 153.835 ;
        RECT 85.735 153.205 86.855 153.375 ;
        RECT 87.025 153.205 87.335 154.005 ;
        RECT 83.935 152.825 85.050 153.035 ;
        RECT 85.735 152.955 85.995 153.205 ;
        RECT 87.505 153.035 87.815 153.835 ;
        RECT 81.865 152.365 82.120 152.695 ;
        RECT 81.525 151.625 81.780 152.200 ;
        RECT 81.950 152.175 82.120 152.365 ;
        RECT 82.400 152.355 82.755 152.725 ;
        RECT 83.005 152.275 83.220 152.815 ;
        RECT 85.240 152.785 85.995 152.955 ;
        RECT 86.785 152.865 87.815 153.035 ;
        RECT 83.390 152.445 84.160 152.645 ;
        RECT 84.330 152.445 85.050 152.645 ;
        RECT 85.240 152.275 85.645 152.785 ;
        RECT 86.785 152.615 86.955 152.865 ;
        RECT 85.815 152.445 86.955 152.615 ;
        RECT 81.950 152.005 82.665 152.175 ;
        RECT 83.005 152.105 84.605 152.275 ;
        RECT 81.950 151.455 82.280 151.835 ;
        RECT 82.495 151.625 82.665 152.005 ;
        RECT 83.435 152.095 84.605 152.105 ;
        RECT 82.975 151.455 83.265 151.925 ;
        RECT 83.435 151.625 83.765 152.095 ;
        RECT 83.935 151.455 84.105 151.925 ;
        RECT 84.275 151.625 84.605 152.095 ;
        RECT 84.775 151.455 85.050 152.275 ;
        RECT 85.240 152.105 86.890 152.275 ;
        RECT 87.125 152.125 87.475 152.695 ;
        RECT 85.285 151.455 85.565 151.935 ;
        RECT 85.735 151.715 85.995 152.105 ;
        RECT 86.170 151.455 86.425 151.935 ;
        RECT 86.595 151.715 86.890 152.105 ;
        RECT 87.645 151.955 87.815 152.865 ;
        RECT 87.985 152.840 88.275 154.005 ;
        RECT 88.445 152.865 88.775 154.005 ;
        RECT 88.945 153.375 89.300 153.835 ;
        RECT 89.470 153.545 90.045 154.005 ;
        RECT 90.215 153.375 90.545 153.835 ;
        RECT 88.945 153.205 90.545 153.375 ;
        RECT 90.745 153.205 91.000 154.005 ;
        RECT 91.755 153.260 92.025 154.005 ;
        RECT 92.655 154.000 98.930 154.005 ;
        RECT 88.945 152.865 89.220 153.205 ;
        RECT 89.400 152.645 89.590 153.025 ;
        RECT 88.445 152.445 89.590 152.645 ;
        RECT 89.770 152.305 90.050 153.205 ;
        RECT 91.170 153.035 91.470 153.230 ;
        RECT 92.195 153.090 92.485 153.830 ;
        RECT 92.655 153.275 92.910 154.000 ;
        RECT 93.095 153.105 93.355 153.830 ;
        RECT 93.525 153.275 93.770 154.000 ;
        RECT 93.955 153.105 94.215 153.830 ;
        RECT 94.385 153.275 94.630 154.000 ;
        RECT 94.815 153.105 95.075 153.830 ;
        RECT 95.245 153.275 95.490 154.000 ;
        RECT 95.660 153.105 95.920 153.830 ;
        RECT 96.090 153.275 96.350 154.000 ;
        RECT 96.520 153.105 96.780 153.830 ;
        RECT 96.950 153.275 97.210 154.000 ;
        RECT 97.380 153.105 97.640 153.830 ;
        RECT 97.810 153.275 98.070 154.000 ;
        RECT 98.240 153.105 98.500 153.830 ;
        RECT 98.670 153.205 98.930 154.000 ;
        RECT 93.095 153.090 98.500 153.105 ;
        RECT 90.220 152.865 91.470 153.035 ;
        RECT 90.220 152.445 90.550 152.865 ;
        RECT 90.780 152.365 91.125 152.695 ;
        RECT 89.770 152.275 90.055 152.305 ;
        RECT 87.070 151.455 87.345 151.935 ;
        RECT 87.515 151.625 87.815 151.955 ;
        RECT 87.985 151.455 88.275 152.180 ;
        RECT 88.445 152.065 89.555 152.275 ;
        RECT 88.445 151.625 88.795 152.065 ;
        RECT 88.965 151.455 89.135 151.895 ;
        RECT 89.305 151.835 89.555 152.065 ;
        RECT 89.725 152.005 90.055 152.275 ;
        RECT 90.225 151.835 90.500 152.275 ;
        RECT 91.300 152.210 91.470 152.865 ;
        RECT 89.305 151.625 90.500 151.835 ;
        RECT 90.735 151.455 91.065 152.195 ;
        RECT 91.235 151.880 91.470 152.210 ;
        RECT 91.755 152.865 98.500 153.090 ;
        RECT 91.755 152.275 92.920 152.865 ;
        RECT 99.100 152.695 99.350 153.830 ;
        RECT 99.530 153.195 99.790 154.005 ;
        RECT 99.965 152.695 100.210 153.835 ;
        RECT 100.390 153.195 100.685 154.005 ;
        RECT 100.865 152.840 101.155 154.005 ;
        RECT 101.415 153.260 101.685 154.005 ;
        RECT 102.315 154.000 108.590 154.005 ;
        RECT 101.855 153.090 102.145 153.830 ;
        RECT 102.315 153.275 102.570 154.000 ;
        RECT 102.755 153.105 103.015 153.830 ;
        RECT 103.185 153.275 103.430 154.000 ;
        RECT 103.615 153.105 103.875 153.830 ;
        RECT 104.045 153.275 104.290 154.000 ;
        RECT 104.475 153.105 104.735 153.830 ;
        RECT 104.905 153.275 105.150 154.000 ;
        RECT 105.320 153.105 105.580 153.830 ;
        RECT 105.750 153.275 106.010 154.000 ;
        RECT 106.180 153.105 106.440 153.830 ;
        RECT 106.610 153.275 106.870 154.000 ;
        RECT 107.040 153.105 107.300 153.830 ;
        RECT 107.470 153.275 107.730 154.000 ;
        RECT 107.900 153.105 108.160 153.830 ;
        RECT 108.330 153.205 108.590 154.000 ;
        RECT 102.755 153.090 108.160 153.105 ;
        RECT 101.415 152.865 108.160 153.090 ;
        RECT 93.090 152.445 100.210 152.695 ;
        RECT 91.755 152.105 98.500 152.275 ;
        RECT 91.755 151.455 92.055 151.935 ;
        RECT 92.225 151.650 92.485 152.105 ;
        RECT 92.655 151.455 92.915 151.935 ;
        RECT 93.095 151.650 93.355 152.105 ;
        RECT 93.525 151.455 93.775 151.935 ;
        RECT 93.955 151.650 94.215 152.105 ;
        RECT 94.385 151.455 94.635 151.935 ;
        RECT 94.815 151.650 95.075 152.105 ;
        RECT 95.245 151.455 95.490 151.935 ;
        RECT 95.660 151.650 95.935 152.105 ;
        RECT 96.105 151.455 96.350 151.935 ;
        RECT 96.520 151.650 96.780 152.105 ;
        RECT 96.950 151.455 97.210 151.935 ;
        RECT 97.380 151.650 97.640 152.105 ;
        RECT 97.810 151.455 98.070 151.935 ;
        RECT 98.240 151.650 98.500 152.105 ;
        RECT 98.670 151.455 98.930 152.015 ;
        RECT 99.100 151.635 99.350 152.445 ;
        RECT 99.530 151.455 99.790 151.980 ;
        RECT 99.960 151.635 100.210 152.445 ;
        RECT 100.380 152.135 100.695 152.695 ;
        RECT 101.415 152.305 102.580 152.865 ;
        RECT 108.760 152.695 109.010 153.830 ;
        RECT 109.190 153.195 109.450 154.005 ;
        RECT 109.625 152.695 109.870 153.835 ;
        RECT 110.050 153.195 110.345 154.005 ;
        RECT 110.525 152.865 110.855 154.005 ;
        RECT 111.025 153.375 111.380 153.835 ;
        RECT 111.550 153.545 112.125 154.005 ;
        RECT 112.295 153.375 112.625 153.835 ;
        RECT 111.025 153.205 112.625 153.375 ;
        RECT 112.825 153.205 113.080 154.005 ;
        RECT 111.025 152.865 111.300 153.205 ;
        RECT 102.750 152.445 109.870 152.695 ;
        RECT 101.385 152.275 102.580 152.305 ;
        RECT 100.390 151.455 100.695 151.965 ;
        RECT 100.865 151.455 101.155 152.180 ;
        RECT 101.385 152.135 108.160 152.275 ;
        RECT 101.415 152.105 108.160 152.135 ;
        RECT 101.415 151.455 101.715 151.935 ;
        RECT 101.885 151.650 102.145 152.105 ;
        RECT 102.315 151.455 102.575 151.935 ;
        RECT 102.755 151.650 103.015 152.105 ;
        RECT 103.185 151.455 103.435 151.935 ;
        RECT 103.615 151.650 103.875 152.105 ;
        RECT 104.045 151.455 104.295 151.935 ;
        RECT 104.475 151.650 104.735 152.105 ;
        RECT 104.905 151.455 105.150 151.935 ;
        RECT 105.320 151.650 105.595 152.105 ;
        RECT 105.765 151.455 106.010 151.935 ;
        RECT 106.180 151.650 106.440 152.105 ;
        RECT 106.610 151.455 106.870 151.935 ;
        RECT 107.040 151.650 107.300 152.105 ;
        RECT 107.470 151.455 107.730 151.935 ;
        RECT 107.900 151.650 108.160 152.105 ;
        RECT 108.330 151.455 108.590 152.015 ;
        RECT 108.760 151.635 109.010 152.445 ;
        RECT 109.190 151.455 109.450 151.980 ;
        RECT 109.620 151.635 109.870 152.445 ;
        RECT 110.040 152.135 110.355 152.695 ;
        RECT 111.480 152.645 111.670 153.025 ;
        RECT 110.525 152.445 111.670 152.645 ;
        RECT 111.850 152.275 112.130 153.205 ;
        RECT 113.250 153.035 113.550 153.230 ;
        RECT 112.300 152.865 113.550 153.035 ;
        RECT 112.300 152.445 112.630 152.865 ;
        RECT 112.860 152.365 113.205 152.695 ;
        RECT 110.525 152.065 111.635 152.275 ;
        RECT 110.050 151.455 110.355 151.965 ;
        RECT 110.525 151.625 110.875 152.065 ;
        RECT 111.045 151.455 111.215 151.895 ;
        RECT 111.385 151.835 111.635 152.065 ;
        RECT 111.805 152.175 112.130 152.275 ;
        RECT 111.805 152.005 112.135 152.175 ;
        RECT 112.305 151.835 112.580 152.275 ;
        RECT 113.380 152.210 113.550 152.865 ;
        RECT 113.745 152.840 114.035 154.005 ;
        RECT 114.265 153.305 114.485 153.835 ;
        RECT 114.655 153.495 114.985 154.005 ;
        RECT 115.155 153.305 115.380 153.835 ;
        RECT 114.265 153.040 115.380 153.305 ;
        RECT 115.550 153.290 115.865 153.835 ;
        RECT 116.055 153.590 116.385 154.005 ;
        RECT 115.550 153.060 116.385 153.290 ;
        RECT 111.385 151.625 112.580 151.835 ;
        RECT 112.815 151.455 113.145 152.195 ;
        RECT 113.315 151.880 113.550 152.210 ;
        RECT 113.745 151.455 114.035 152.180 ;
        RECT 114.215 152.120 114.530 152.695 ;
        RECT 114.205 151.455 114.535 151.935 ;
        RECT 114.720 151.735 115.100 152.695 ;
        RECT 115.550 152.365 115.875 152.780 ;
        RECT 116.045 152.365 116.385 153.060 ;
        RECT 116.045 152.195 116.215 152.365 ;
        RECT 116.555 152.195 116.785 153.835 ;
        RECT 116.955 153.035 117.245 154.005 ;
        RECT 117.515 153.260 117.785 154.005 ;
        RECT 118.415 154.000 124.690 154.005 ;
        RECT 117.955 153.090 118.245 153.830 ;
        RECT 118.415 153.275 118.670 154.000 ;
        RECT 118.855 153.105 119.115 153.830 ;
        RECT 119.285 153.275 119.530 154.000 ;
        RECT 119.715 153.105 119.975 153.830 ;
        RECT 120.145 153.275 120.390 154.000 ;
        RECT 120.575 153.105 120.835 153.830 ;
        RECT 121.005 153.275 121.250 154.000 ;
        RECT 121.420 153.105 121.680 153.830 ;
        RECT 121.850 153.275 122.110 154.000 ;
        RECT 122.280 153.105 122.540 153.830 ;
        RECT 122.710 153.275 122.970 154.000 ;
        RECT 123.140 153.105 123.400 153.830 ;
        RECT 123.570 153.275 123.830 154.000 ;
        RECT 124.000 153.105 124.260 153.830 ;
        RECT 124.430 153.205 124.690 154.000 ;
        RECT 118.855 153.090 124.260 153.105 ;
        RECT 117.515 152.985 124.260 153.090 ;
        RECT 117.485 152.865 124.260 152.985 ;
        RECT 117.485 152.815 118.680 152.865 ;
        RECT 115.475 152.025 116.215 152.195 ;
        RECT 115.475 151.625 115.665 152.025 ;
        RECT 116.385 152.005 116.785 152.195 ;
        RECT 117.515 152.275 118.680 152.815 ;
        RECT 124.860 152.695 125.110 153.830 ;
        RECT 125.290 153.195 125.550 154.005 ;
        RECT 125.725 152.695 125.970 153.835 ;
        RECT 126.150 153.195 126.445 154.005 ;
        RECT 126.625 152.840 126.915 154.005 ;
        RECT 127.085 153.410 127.520 153.835 ;
        RECT 127.690 153.580 128.075 154.005 ;
        RECT 127.085 153.240 128.075 153.410 ;
        RECT 118.850 152.445 125.970 152.695 ;
        RECT 117.515 152.105 124.260 152.275 ;
        RECT 115.885 151.455 116.215 151.815 ;
        RECT 116.385 151.625 116.575 152.005 ;
        RECT 116.745 151.455 117.075 151.835 ;
        RECT 117.515 151.455 117.815 151.935 ;
        RECT 117.985 151.650 118.245 152.105 ;
        RECT 118.415 151.455 118.675 151.935 ;
        RECT 118.855 151.650 119.115 152.105 ;
        RECT 119.285 151.455 119.535 151.935 ;
        RECT 119.715 151.650 119.975 152.105 ;
        RECT 120.145 151.455 120.395 151.935 ;
        RECT 120.575 151.650 120.835 152.105 ;
        RECT 121.005 151.455 121.250 151.935 ;
        RECT 121.420 151.650 121.695 152.105 ;
        RECT 121.865 151.455 122.110 151.935 ;
        RECT 122.280 151.650 122.540 152.105 ;
        RECT 122.710 151.455 122.970 151.935 ;
        RECT 123.140 151.650 123.400 152.105 ;
        RECT 123.570 151.455 123.830 151.935 ;
        RECT 124.000 151.650 124.260 152.105 ;
        RECT 124.430 151.455 124.690 152.015 ;
        RECT 124.860 151.635 125.110 152.445 ;
        RECT 125.290 151.455 125.550 151.980 ;
        RECT 125.720 151.635 125.970 152.445 ;
        RECT 126.140 152.135 126.455 152.695 ;
        RECT 127.085 152.365 127.570 153.070 ;
        RECT 127.740 152.695 128.075 153.240 ;
        RECT 128.245 153.045 128.670 153.835 ;
        RECT 128.840 153.410 129.115 153.835 ;
        RECT 129.285 153.580 129.670 154.005 ;
        RECT 128.840 153.215 129.670 153.410 ;
        RECT 128.245 152.865 129.150 153.045 ;
        RECT 127.740 152.365 128.150 152.695 ;
        RECT 128.320 152.365 129.150 152.865 ;
        RECT 129.320 152.695 129.670 153.215 ;
        RECT 129.840 153.045 130.085 153.835 ;
        RECT 130.275 153.410 130.530 153.835 ;
        RECT 130.700 153.580 131.085 154.005 ;
        RECT 130.275 153.215 131.085 153.410 ;
        RECT 129.840 152.865 130.565 153.045 ;
        RECT 129.320 152.365 129.745 152.695 ;
        RECT 129.915 152.365 130.565 152.865 ;
        RECT 130.735 152.695 131.085 153.215 ;
        RECT 131.255 152.865 131.515 153.835 ;
        RECT 131.695 153.205 132.025 154.005 ;
        RECT 132.205 153.665 133.635 153.835 ;
        RECT 132.205 153.035 132.455 153.665 ;
        RECT 130.735 152.365 131.160 152.695 ;
        RECT 127.740 152.195 128.075 152.365 ;
        RECT 128.320 152.195 128.670 152.365 ;
        RECT 129.320 152.195 129.670 152.365 ;
        RECT 129.915 152.195 130.085 152.365 ;
        RECT 130.735 152.195 131.085 152.365 ;
        RECT 131.330 152.195 131.515 152.865 ;
        RECT 126.150 151.455 126.455 151.965 ;
        RECT 126.625 151.455 126.915 152.180 ;
        RECT 127.085 152.025 128.075 152.195 ;
        RECT 127.085 151.625 127.520 152.025 ;
        RECT 127.690 151.455 128.075 151.855 ;
        RECT 128.245 151.625 128.670 152.195 ;
        RECT 128.860 152.025 129.670 152.195 ;
        RECT 128.860 151.625 129.115 152.025 ;
        RECT 129.285 151.455 129.670 151.855 ;
        RECT 129.840 151.625 130.085 152.195 ;
        RECT 130.275 152.025 131.085 152.195 ;
        RECT 130.275 151.625 130.530 152.025 ;
        RECT 130.700 151.455 131.085 151.855 ;
        RECT 131.255 151.625 131.515 152.195 ;
        RECT 131.685 152.865 132.455 153.035 ;
        RECT 131.685 152.195 131.855 152.865 ;
        RECT 132.025 152.365 132.430 152.695 ;
        RECT 132.645 152.365 132.895 153.495 ;
        RECT 133.095 152.695 133.295 153.495 ;
        RECT 133.465 152.985 133.635 153.665 ;
        RECT 133.805 153.155 134.120 154.005 ;
        RECT 134.295 153.205 134.735 153.835 ;
        RECT 133.465 152.815 134.255 152.985 ;
        RECT 133.095 152.365 133.340 152.695 ;
        RECT 133.525 152.365 133.915 152.645 ;
        RECT 134.085 152.365 134.255 152.815 ;
        RECT 134.425 152.195 134.735 153.205 ;
        RECT 134.905 152.915 136.115 154.005 ;
        RECT 134.905 152.375 135.425 152.915 ;
        RECT 135.595 152.205 136.115 152.745 ;
        RECT 131.685 151.625 132.175 152.195 ;
        RECT 132.345 152.025 133.505 152.195 ;
        RECT 132.345 151.625 132.575 152.025 ;
        RECT 132.745 151.455 133.165 151.855 ;
        RECT 133.335 151.625 133.505 152.025 ;
        RECT 133.675 151.455 134.125 152.195 ;
        RECT 134.295 151.635 134.735 152.195 ;
        RECT 134.905 151.455 136.115 152.205 ;
        RECT 23.500 151.285 136.200 151.455 ;
        RECT 50.705 70.245 110.465 70.695 ;
        RECT 50.705 70.115 110.525 70.245 ;
        RECT 50.485 69.875 110.525 70.115 ;
        RECT 50.485 69.630 52.195 69.875 ;
        RECT 58.775 69.645 60.485 69.875 ;
        RECT 46.190 69.460 50.000 69.630 ;
        RECT 46.190 63.650 46.360 69.460 ;
        RECT 46.840 66.820 47.530 68.980 ;
        RECT 46.840 64.130 47.530 66.290 ;
        RECT 48.010 63.650 48.180 69.460 ;
        RECT 48.660 66.820 49.350 68.980 ;
        RECT 48.660 64.130 49.350 66.290 ;
        RECT 49.830 63.650 50.000 69.460 ;
        RECT 46.190 63.480 50.000 63.650 ;
        RECT 1.470 57.840 13.600 58.010 ;
        RECT 1.470 56.190 1.640 57.840 ;
        RECT 2.120 56.670 4.280 57.360 ;
        RECT 4.810 56.670 6.970 57.360 ;
        RECT 7.450 56.190 7.620 57.840 ;
        RECT 8.100 56.670 10.260 57.360 ;
        RECT 10.790 56.670 12.950 57.360 ;
        RECT 13.430 56.190 13.600 57.840 ;
        RECT 46.190 57.670 46.360 63.480 ;
        RECT 46.840 60.840 47.530 63.000 ;
        RECT 46.840 58.150 47.530 60.310 ;
        RECT 48.010 57.670 48.180 63.480 ;
        RECT 48.660 60.840 49.350 63.000 ;
        RECT 48.660 58.150 49.350 60.310 ;
        RECT 49.830 57.670 50.000 63.480 ;
        RECT 50.480 69.460 52.230 69.630 ;
        RECT 50.480 61.970 50.650 69.460 ;
        RECT 51.190 68.950 51.520 69.120 ;
        RECT 51.050 62.695 51.220 68.735 ;
        RECT 51.490 62.695 51.660 68.735 ;
        RECT 51.190 62.310 51.520 62.480 ;
        RECT 52.060 61.970 52.230 69.460 ;
        RECT 50.480 61.800 52.230 61.970 ;
        RECT 52.655 69.475 58.285 69.645 ;
        RECT 52.655 63.665 52.825 69.475 ;
        RECT 53.305 66.835 53.995 68.995 ;
        RECT 53.305 64.145 53.995 66.305 ;
        RECT 54.475 63.665 54.645 69.475 ;
        RECT 55.125 66.835 55.815 68.995 ;
        RECT 55.125 64.145 55.815 66.305 ;
        RECT 56.295 63.665 56.465 69.475 ;
        RECT 56.945 66.835 57.635 68.995 ;
        RECT 56.945 64.145 57.635 66.305 ;
        RECT 58.115 63.665 58.285 69.475 ;
        RECT 52.655 63.495 58.285 63.665 ;
        RECT 50.460 61.075 52.210 61.245 ;
        RECT 50.460 57.675 50.630 61.075 ;
        RECT 51.170 60.565 51.500 60.735 ;
        RECT 51.030 58.355 51.200 60.395 ;
        RECT 51.470 58.355 51.640 60.395 ;
        RECT 51.170 58.015 51.500 58.185 ;
        RECT 52.040 57.675 52.210 61.075 ;
        RECT 50.460 57.670 52.210 57.675 ;
        RECT 52.655 57.685 52.825 63.495 ;
        RECT 53.305 60.855 53.995 63.015 ;
        RECT 53.305 58.165 53.995 60.325 ;
        RECT 54.475 57.685 54.645 63.495 ;
        RECT 55.125 60.855 55.815 63.015 ;
        RECT 55.125 58.165 55.815 60.325 ;
        RECT 56.295 57.685 56.465 63.495 ;
        RECT 56.945 60.855 57.635 63.015 ;
        RECT 56.945 58.165 57.635 60.325 ;
        RECT 58.115 57.685 58.285 63.495 ;
        RECT 58.775 69.475 60.525 69.645 ;
        RECT 58.775 61.985 58.945 69.475 ;
        RECT 59.485 68.965 59.815 69.135 ;
        RECT 59.345 62.710 59.515 68.750 ;
        RECT 59.785 62.710 59.955 68.750 ;
        RECT 59.485 62.325 59.815 62.495 ;
        RECT 60.355 61.985 60.525 69.475 ;
        RECT 58.775 61.815 60.525 61.985 ;
        RECT 60.985 69.465 66.615 69.635 ;
        RECT 60.985 63.655 61.155 69.465 ;
        RECT 61.635 66.825 62.325 68.985 ;
        RECT 61.635 64.135 62.325 66.295 ;
        RECT 62.805 63.655 62.975 69.465 ;
        RECT 63.455 66.825 64.145 68.985 ;
        RECT 63.455 64.135 64.145 66.295 ;
        RECT 64.625 63.655 64.795 69.465 ;
        RECT 65.275 66.825 65.965 68.985 ;
        RECT 65.275 64.135 65.965 66.295 ;
        RECT 66.445 63.655 66.615 69.465 ;
        RECT 66.915 69.485 69.035 69.875 ;
        RECT 75.425 69.675 77.325 69.875 ;
        RECT 66.915 69.405 69.015 69.485 ;
        RECT 69.280 69.455 74.910 69.625 ;
        RECT 60.985 63.485 66.615 63.655 ;
        RECT 52.655 57.670 58.285 57.685 ;
        RECT 58.765 61.075 60.515 61.245 ;
        RECT 58.765 57.675 58.935 61.075 ;
        RECT 59.475 60.565 59.805 60.735 ;
        RECT 59.335 58.355 59.505 60.395 ;
        RECT 59.775 58.355 59.945 60.395 ;
        RECT 59.475 58.015 59.805 58.185 ;
        RECT 60.345 57.675 60.515 61.075 ;
        RECT 58.765 57.670 60.515 57.675 ;
        RECT 60.985 57.675 61.155 63.485 ;
        RECT 61.635 60.845 62.325 63.005 ;
        RECT 61.635 58.155 62.325 60.315 ;
        RECT 62.805 57.675 62.975 63.485 ;
        RECT 63.455 60.845 64.145 63.005 ;
        RECT 63.455 58.155 64.145 60.315 ;
        RECT 64.625 57.675 64.795 63.485 ;
        RECT 65.275 60.845 65.965 63.005 ;
        RECT 65.275 58.155 65.965 60.315 ;
        RECT 66.445 57.675 66.615 63.485 ;
        RECT 67.090 61.975 67.260 69.405 ;
        RECT 67.800 68.955 68.130 69.125 ;
        RECT 67.660 62.700 67.830 68.740 ;
        RECT 68.100 62.700 68.270 68.740 ;
        RECT 67.800 62.315 68.130 62.485 ;
        RECT 68.670 61.975 68.840 69.405 ;
        RECT 67.090 61.805 68.840 61.975 ;
        RECT 69.280 63.645 69.450 69.455 ;
        RECT 69.930 66.815 70.620 68.975 ;
        RECT 69.930 64.125 70.620 66.285 ;
        RECT 71.100 63.645 71.270 69.455 ;
        RECT 71.750 66.815 72.440 68.975 ;
        RECT 71.750 64.125 72.440 66.285 ;
        RECT 72.920 63.645 73.090 69.455 ;
        RECT 73.570 66.815 74.260 68.975 ;
        RECT 73.570 64.125 74.260 66.285 ;
        RECT 74.740 63.645 74.910 69.455 ;
        RECT 69.280 63.475 74.910 63.645 ;
        RECT 60.985 57.670 66.615 57.675 ;
        RECT 67.025 61.075 68.775 61.245 ;
        RECT 67.025 57.675 67.195 61.075 ;
        RECT 67.735 60.565 68.065 60.735 ;
        RECT 67.595 58.355 67.765 60.395 ;
        RECT 68.035 58.355 68.205 60.395 ;
        RECT 67.735 58.015 68.065 58.185 ;
        RECT 68.605 57.675 68.775 61.075 ;
        RECT 67.025 57.670 68.775 57.675 ;
        RECT 69.280 57.670 69.450 63.475 ;
        RECT 69.930 60.835 70.620 62.995 ;
        RECT 69.930 58.145 70.620 60.305 ;
        RECT 71.100 57.670 71.270 63.475 ;
        RECT 71.750 60.835 72.440 62.995 ;
        RECT 71.750 58.145 72.440 60.305 ;
        RECT 72.920 57.670 73.090 63.475 ;
        RECT 73.570 60.835 74.260 62.995 ;
        RECT 73.570 58.145 74.260 60.305 ;
        RECT 74.740 57.670 74.910 63.475 ;
        RECT 75.470 69.565 77.220 69.675 ;
        RECT 83.865 69.660 85.575 69.875 ;
        RECT 92.195 69.685 93.905 69.875 ;
        RECT 100.485 69.700 102.195 69.875 ;
        RECT 75.470 62.075 75.640 69.565 ;
        RECT 76.180 69.055 76.510 69.225 ;
        RECT 76.040 62.800 76.210 68.840 ;
        RECT 76.480 62.800 76.650 68.840 ;
        RECT 76.180 62.415 76.510 62.585 ;
        RECT 77.050 62.075 77.220 69.565 ;
        RECT 75.470 61.905 77.220 62.075 ;
        RECT 77.725 69.470 83.355 69.640 ;
        RECT 77.725 63.660 77.895 69.470 ;
        RECT 78.375 66.830 79.065 68.990 ;
        RECT 78.375 64.140 79.065 66.300 ;
        RECT 79.545 63.660 79.715 69.470 ;
        RECT 80.195 66.830 80.885 68.990 ;
        RECT 80.195 64.140 80.885 66.300 ;
        RECT 81.365 63.660 81.535 69.470 ;
        RECT 82.015 66.830 82.705 68.990 ;
        RECT 82.015 64.140 82.705 66.300 ;
        RECT 83.185 63.660 83.355 69.470 ;
        RECT 77.725 63.490 83.355 63.660 ;
        RECT 75.445 61.095 77.195 61.265 ;
        RECT 75.445 57.695 75.615 61.095 ;
        RECT 76.155 60.585 76.485 60.755 ;
        RECT 76.015 58.375 76.185 60.415 ;
        RECT 76.455 58.375 76.625 60.415 ;
        RECT 76.155 58.035 76.485 58.205 ;
        RECT 77.025 57.695 77.195 61.095 ;
        RECT 75.445 57.670 77.195 57.695 ;
        RECT 77.725 57.680 77.895 63.490 ;
        RECT 78.375 60.850 79.065 63.010 ;
        RECT 78.375 58.160 79.065 60.320 ;
        RECT 79.545 57.680 79.715 63.490 ;
        RECT 80.195 60.850 80.885 63.010 ;
        RECT 80.195 58.160 80.885 60.320 ;
        RECT 81.365 57.680 81.535 63.490 ;
        RECT 82.015 60.850 82.705 63.010 ;
        RECT 82.015 58.160 82.705 60.320 ;
        RECT 83.185 57.680 83.355 63.490 ;
        RECT 83.860 69.490 85.610 69.660 ;
        RECT 83.860 62.000 84.030 69.490 ;
        RECT 84.570 68.980 84.900 69.150 ;
        RECT 84.430 62.725 84.600 68.765 ;
        RECT 84.870 62.725 85.040 68.765 ;
        RECT 84.570 62.340 84.900 62.510 ;
        RECT 85.440 62.000 85.610 69.490 ;
        RECT 83.860 61.830 85.610 62.000 ;
        RECT 86.055 69.470 91.685 69.640 ;
        RECT 86.055 63.660 86.225 69.470 ;
        RECT 86.705 66.830 87.395 68.990 ;
        RECT 86.705 64.140 87.395 66.300 ;
        RECT 87.875 63.660 88.045 69.470 ;
        RECT 88.525 66.830 89.215 68.990 ;
        RECT 88.525 64.140 89.215 66.300 ;
        RECT 89.695 63.660 89.865 69.470 ;
        RECT 90.345 66.830 91.035 68.990 ;
        RECT 90.345 64.140 91.035 66.300 ;
        RECT 91.515 63.660 91.685 69.470 ;
        RECT 86.055 63.490 91.685 63.660 ;
        RECT 77.725 57.670 83.355 57.680 ;
        RECT 83.795 61.075 85.545 61.245 ;
        RECT 83.795 57.675 83.965 61.075 ;
        RECT 84.505 60.565 84.835 60.735 ;
        RECT 84.365 58.355 84.535 60.395 ;
        RECT 84.805 58.355 84.975 60.395 ;
        RECT 84.505 58.015 84.835 58.185 ;
        RECT 85.375 57.675 85.545 61.075 ;
        RECT 83.795 57.670 85.545 57.675 ;
        RECT 86.055 57.680 86.225 63.490 ;
        RECT 86.705 60.850 87.395 63.010 ;
        RECT 86.705 58.160 87.395 60.320 ;
        RECT 87.875 57.680 88.045 63.490 ;
        RECT 88.525 60.850 89.215 63.010 ;
        RECT 88.525 58.160 89.215 60.320 ;
        RECT 89.695 57.680 89.865 63.490 ;
        RECT 90.345 60.850 91.035 63.010 ;
        RECT 90.345 58.160 91.035 60.320 ;
        RECT 91.515 57.680 91.685 63.490 ;
        RECT 92.190 69.515 93.940 69.685 ;
        RECT 92.190 62.025 92.360 69.515 ;
        RECT 92.900 69.005 93.230 69.175 ;
        RECT 92.760 62.750 92.930 68.790 ;
        RECT 93.200 62.750 93.370 68.790 ;
        RECT 92.900 62.365 93.230 62.535 ;
        RECT 93.770 62.025 93.940 69.515 ;
        RECT 92.190 61.855 93.940 62.025 ;
        RECT 94.385 69.470 100.015 69.640 ;
        RECT 94.385 63.660 94.555 69.470 ;
        RECT 95.035 66.830 95.725 68.990 ;
        RECT 95.035 64.140 95.725 66.300 ;
        RECT 96.205 63.660 96.375 69.470 ;
        RECT 96.855 66.830 97.545 68.990 ;
        RECT 96.855 64.140 97.545 66.300 ;
        RECT 98.025 63.660 98.195 69.470 ;
        RECT 98.675 66.830 99.365 68.990 ;
        RECT 98.675 64.140 99.365 66.300 ;
        RECT 99.845 63.660 100.015 69.470 ;
        RECT 94.385 63.490 100.015 63.660 ;
        RECT 86.055 57.670 91.685 57.680 ;
        RECT 92.180 61.070 93.930 61.240 ;
        RECT 92.180 57.670 92.350 61.070 ;
        RECT 92.890 60.560 93.220 60.730 ;
        RECT 92.750 58.350 92.920 60.390 ;
        RECT 93.190 58.350 93.360 60.390 ;
        RECT 92.890 58.010 93.220 58.180 ;
        RECT 93.760 57.670 93.930 61.070 ;
        RECT 94.385 57.680 94.555 63.490 ;
        RECT 95.035 60.850 95.725 63.010 ;
        RECT 95.035 58.160 95.725 60.320 ;
        RECT 96.205 57.680 96.375 63.490 ;
        RECT 96.855 60.850 97.545 63.010 ;
        RECT 96.855 58.160 97.545 60.320 ;
        RECT 98.025 57.680 98.195 63.490 ;
        RECT 98.675 60.850 99.365 63.010 ;
        RECT 98.675 58.160 99.365 60.320 ;
        RECT 99.845 57.680 100.015 63.490 ;
        RECT 100.485 69.530 102.235 69.700 ;
        RECT 108.815 69.680 110.525 69.875 ;
        RECT 100.485 62.040 100.655 69.530 ;
        RECT 101.195 69.020 101.525 69.190 ;
        RECT 101.055 62.765 101.225 68.805 ;
        RECT 101.495 62.765 101.665 68.805 ;
        RECT 101.195 62.380 101.525 62.550 ;
        RECT 102.065 62.040 102.235 69.530 ;
        RECT 100.485 61.870 102.235 62.040 ;
        RECT 102.690 69.465 108.320 69.635 ;
        RECT 102.690 63.655 102.860 69.465 ;
        RECT 103.340 66.825 104.030 68.985 ;
        RECT 103.340 64.135 104.030 66.295 ;
        RECT 104.510 63.655 104.680 69.465 ;
        RECT 105.160 66.825 105.850 68.985 ;
        RECT 105.160 64.135 105.850 66.295 ;
        RECT 106.330 63.655 106.500 69.465 ;
        RECT 106.980 66.825 107.670 68.985 ;
        RECT 106.980 64.135 107.670 66.295 ;
        RECT 108.150 63.655 108.320 69.465 ;
        RECT 102.690 63.485 108.320 63.655 ;
        RECT 94.385 57.670 100.015 57.680 ;
        RECT 100.420 61.080 102.170 61.250 ;
        RECT 100.420 57.680 100.590 61.080 ;
        RECT 101.130 60.570 101.460 60.740 ;
        RECT 100.990 58.360 101.160 60.400 ;
        RECT 101.430 58.360 101.600 60.400 ;
        RECT 101.130 58.020 101.460 58.190 ;
        RECT 102.000 57.680 102.170 61.080 ;
        RECT 100.420 57.670 102.170 57.680 ;
        RECT 102.690 57.675 102.860 63.485 ;
        RECT 103.340 60.845 104.030 63.005 ;
        RECT 103.340 58.155 104.030 60.315 ;
        RECT 104.510 57.675 104.680 63.485 ;
        RECT 105.160 60.845 105.850 63.005 ;
        RECT 105.160 58.155 105.850 60.315 ;
        RECT 106.330 57.675 106.500 63.485 ;
        RECT 106.980 60.845 107.670 63.005 ;
        RECT 106.980 58.155 107.670 60.315 ;
        RECT 108.150 57.675 108.320 63.485 ;
        RECT 108.785 69.510 110.535 69.680 ;
        RECT 108.785 62.020 108.955 69.510 ;
        RECT 109.495 69.000 109.825 69.170 ;
        RECT 109.355 62.745 109.525 68.785 ;
        RECT 109.795 62.745 109.965 68.785 ;
        RECT 109.495 62.360 109.825 62.530 ;
        RECT 110.365 62.020 110.535 69.510 ;
        RECT 108.785 61.850 110.535 62.020 ;
        RECT 110.990 69.475 114.800 69.645 ;
        RECT 110.990 63.665 111.160 69.475 ;
        RECT 111.640 66.835 112.330 68.995 ;
        RECT 111.640 64.145 112.330 66.305 ;
        RECT 112.810 63.665 112.980 69.475 ;
        RECT 113.460 66.835 114.150 68.995 ;
        RECT 113.460 64.145 114.150 66.305 ;
        RECT 114.630 63.665 114.800 69.475 ;
        RECT 110.990 63.495 114.800 63.665 ;
        RECT 102.690 57.670 108.320 57.675 ;
        RECT 108.785 61.080 110.535 61.250 ;
        RECT 108.785 57.680 108.955 61.080 ;
        RECT 109.495 60.570 109.825 60.740 ;
        RECT 109.355 58.360 109.525 60.400 ;
        RECT 109.795 58.360 109.965 60.400 ;
        RECT 109.495 58.020 109.825 58.190 ;
        RECT 110.365 57.680 110.535 61.080 ;
        RECT 108.785 57.670 110.535 57.680 ;
        RECT 110.990 57.685 111.160 63.495 ;
        RECT 111.640 60.855 112.330 63.015 ;
        RECT 111.640 58.165 112.330 60.325 ;
        RECT 112.810 57.685 112.980 63.495 ;
        RECT 113.460 60.855 114.150 63.015 ;
        RECT 113.460 58.165 114.150 60.325 ;
        RECT 114.630 57.685 114.800 63.495 ;
        RECT 110.990 57.670 114.800 57.685 ;
        RECT 46.190 56.795 114.805 57.670 ;
        RECT 1.470 56.020 13.600 56.190 ;
        RECT 1.470 54.370 1.640 56.020 ;
        RECT 2.120 54.850 4.280 55.540 ;
        RECT 4.810 54.850 6.970 55.540 ;
        RECT 7.450 54.370 7.620 56.020 ;
        RECT 8.100 54.850 10.260 55.540 ;
        RECT 10.790 54.850 12.950 55.540 ;
        RECT 13.430 54.370 13.600 56.020 ;
        RECT 1.470 54.200 13.600 54.370 ;
        RECT 1.470 52.550 1.640 54.200 ;
        RECT 2.120 53.030 4.280 53.720 ;
        RECT 4.810 53.030 6.970 53.720 ;
        RECT 7.450 52.550 7.620 54.200 ;
        RECT 8.100 53.030 10.260 53.720 ;
        RECT 10.790 53.030 12.950 53.720 ;
        RECT 13.430 52.550 13.600 54.200 ;
        RECT 1.470 52.380 31.540 52.550 ;
        RECT 1.470 50.855 1.640 52.380 ;
        RECT 2.120 51.210 4.280 51.900 ;
        RECT 4.810 51.210 6.970 51.900 ;
        RECT 7.450 50.855 7.620 52.380 ;
        RECT 8.100 51.210 10.260 51.900 ;
        RECT 10.790 51.210 12.950 51.900 ;
        RECT 1.470 50.730 9.960 50.855 ;
        RECT 13.430 50.730 13.600 52.380 ;
        RECT 14.080 51.210 16.240 51.900 ;
        RECT 16.770 51.210 18.930 51.900 ;
        RECT 19.410 50.730 19.580 52.380 ;
        RECT 20.060 51.210 22.220 51.900 ;
        RECT 22.750 51.210 24.910 51.900 ;
        RECT 25.390 50.730 25.560 52.380 ;
        RECT 26.040 51.210 28.200 51.900 ;
        RECT 28.730 51.210 30.890 51.900 ;
        RECT 31.370 50.730 31.540 52.380 ;
        RECT 1.470 50.560 31.540 50.730 ;
        RECT 43.490 52.540 61.600 52.550 ;
        RECT 67.490 52.540 85.600 52.550 ;
        RECT 43.490 52.380 85.600 52.540 ;
        RECT 43.490 50.730 43.660 52.380 ;
        RECT 44.140 51.210 46.300 51.900 ;
        RECT 46.830 51.210 48.990 51.900 ;
        RECT 49.470 50.730 49.640 52.380 ;
        RECT 50.120 51.210 52.280 51.900 ;
        RECT 52.810 51.210 54.970 51.900 ;
        RECT 55.450 50.730 55.620 52.380 ;
        RECT 61.430 52.090 67.670 52.380 ;
        RECT 56.100 51.210 58.260 51.900 ;
        RECT 58.790 51.210 60.950 51.900 ;
        RECT 61.430 50.730 61.600 52.090 ;
        RECT 43.490 50.560 61.600 50.730 ;
        RECT 67.490 50.730 67.660 52.090 ;
        RECT 68.140 51.210 70.300 51.900 ;
        RECT 70.830 51.210 72.990 51.900 ;
        RECT 73.470 50.730 73.640 52.380 ;
        RECT 74.120 51.210 76.280 51.900 ;
        RECT 76.810 51.210 78.970 51.900 ;
        RECT 79.450 50.730 79.620 52.380 ;
        RECT 80.100 51.210 82.260 51.900 ;
        RECT 82.790 51.210 84.950 51.900 ;
        RECT 85.430 50.730 85.600 52.380 ;
        RECT 67.490 50.560 85.600 50.730 ;
        RECT 1.585 50.360 9.960 50.560 ;
        RECT 77.790 50.170 80.360 50.560 ;
        RECT 1.450 49.480 27.925 49.960 ;
        RECT 29.450 49.480 55.925 49.960 ;
        RECT 57.450 49.480 83.925 49.960 ;
        RECT 85.450 49.480 111.925 49.960 ;
        RECT 113.450 49.480 139.925 49.960 ;
        RECT 1.435 49.420 27.925 49.480 ;
        RECT 29.435 49.420 55.925 49.480 ;
        RECT 57.435 49.420 83.925 49.480 ;
        RECT 85.435 49.420 111.925 49.480 ;
        RECT 113.435 49.420 139.925 49.480 ;
        RECT 143.470 49.840 149.620 50.010 ;
        RECT 1.435 49.260 27.980 49.420 ;
        RECT 1.435 49.235 14.180 49.260 ;
        RECT 1.435 49.005 5.760 49.235 ;
        RECT 1.470 39.745 1.640 49.005 ;
        RECT 2.365 48.435 4.405 48.605 ;
        RECT 1.980 40.375 2.150 48.375 ;
        RECT 4.620 40.375 4.790 48.375 ;
        RECT 2.365 40.145 4.405 40.315 ;
        RECT 5.130 39.745 5.300 49.005 ;
        RECT 1.470 39.575 5.300 39.745 ;
        RECT 5.590 39.745 5.760 49.005 ;
        RECT 6.390 48.725 8.390 48.895 ;
        RECT 6.160 40.470 6.330 48.510 ;
        RECT 8.450 40.470 8.620 48.510 ;
        RECT 6.390 40.085 8.390 40.255 ;
        RECT 9.020 39.745 9.190 49.235 ;
        RECT 9.820 48.725 11.820 48.895 ;
        RECT 9.590 40.470 9.760 48.510 ;
        RECT 11.880 40.470 12.050 48.510 ;
        RECT 12.450 47.665 14.180 49.235 ;
        RECT 26.230 49.250 27.980 49.260 ;
        RECT 12.450 47.495 20.915 47.665 ;
        RECT 12.450 46.085 14.255 47.495 ;
        RECT 14.595 46.625 14.765 46.955 ;
        RECT 14.980 46.925 20.020 47.095 ;
        RECT 14.980 46.485 20.020 46.655 ;
        RECT 20.235 46.625 20.405 46.955 ;
        RECT 20.745 46.085 20.915 47.495 ;
        RECT 12.450 45.915 20.915 46.085 ;
        RECT 12.450 45.400 14.180 45.915 ;
        RECT 12.450 45.285 23.930 45.400 ;
        RECT 9.820 40.085 11.820 40.255 ;
        RECT 12.450 39.745 12.620 45.285 ;
        RECT 5.590 39.575 12.620 39.745 ;
        RECT 12.900 45.230 23.930 45.285 ;
        RECT 12.900 39.740 13.070 45.230 ;
        RECT 13.700 44.720 17.700 44.890 ;
        RECT 13.470 40.465 13.640 44.505 ;
        RECT 17.760 40.465 17.930 44.505 ;
        RECT 13.700 40.080 17.700 40.250 ;
        RECT 18.330 39.740 18.500 45.230 ;
        RECT 19.130 44.720 23.130 44.890 ;
        RECT 18.900 40.465 19.070 44.505 ;
        RECT 23.190 40.465 23.360 44.505 ;
        RECT 19.130 40.080 23.130 40.250 ;
        RECT 23.760 39.740 23.930 45.230 ;
        RECT 12.900 39.570 23.930 39.740 ;
        RECT 24.205 45.245 25.955 45.415 ;
        RECT 24.205 39.755 24.375 45.245 ;
        RECT 24.915 44.735 25.245 44.905 ;
        RECT 24.775 40.480 24.945 44.520 ;
        RECT 25.215 40.480 25.385 44.520 ;
        RECT 24.915 40.095 25.245 40.265 ;
        RECT 25.785 39.755 25.955 45.245 ;
        RECT 24.205 39.585 25.955 39.755 ;
        RECT 26.230 39.760 26.400 49.250 ;
        RECT 26.940 48.740 27.270 48.910 ;
        RECT 26.800 40.485 26.970 48.525 ;
        RECT 27.240 40.485 27.410 48.525 ;
        RECT 26.940 40.100 27.270 40.270 ;
        RECT 27.810 39.760 27.980 49.250 ;
        RECT 29.435 49.260 55.980 49.420 ;
        RECT 29.435 49.235 42.180 49.260 ;
        RECT 29.435 49.005 33.760 49.235 ;
        RECT 26.230 39.590 27.980 39.760 ;
        RECT 29.470 39.745 29.640 49.005 ;
        RECT 30.365 48.435 32.405 48.605 ;
        RECT 29.980 40.375 30.150 48.375 ;
        RECT 32.620 40.375 32.790 48.375 ;
        RECT 30.365 40.145 32.405 40.315 ;
        RECT 33.130 39.745 33.300 49.005 ;
        RECT 29.470 39.575 33.300 39.745 ;
        RECT 33.590 39.745 33.760 49.005 ;
        RECT 34.390 48.725 36.390 48.895 ;
        RECT 34.160 40.470 34.330 48.510 ;
        RECT 36.450 40.470 36.620 48.510 ;
        RECT 34.390 40.085 36.390 40.255 ;
        RECT 37.020 39.745 37.190 49.235 ;
        RECT 37.820 48.725 39.820 48.895 ;
        RECT 37.590 40.470 37.760 48.510 ;
        RECT 39.880 40.470 40.050 48.510 ;
        RECT 40.450 47.665 42.180 49.235 ;
        RECT 54.230 49.250 55.980 49.260 ;
        RECT 40.450 47.495 48.915 47.665 ;
        RECT 40.450 46.085 42.255 47.495 ;
        RECT 42.595 46.625 42.765 46.955 ;
        RECT 42.980 46.925 48.020 47.095 ;
        RECT 42.980 46.485 48.020 46.655 ;
        RECT 48.235 46.625 48.405 46.955 ;
        RECT 48.745 46.085 48.915 47.495 ;
        RECT 40.450 45.915 48.915 46.085 ;
        RECT 40.450 45.400 42.180 45.915 ;
        RECT 40.450 45.285 51.930 45.400 ;
        RECT 37.820 40.085 39.820 40.255 ;
        RECT 40.450 39.745 40.620 45.285 ;
        RECT 33.590 39.575 40.620 39.745 ;
        RECT 40.900 45.230 51.930 45.285 ;
        RECT 40.900 39.740 41.070 45.230 ;
        RECT 41.700 44.720 45.700 44.890 ;
        RECT 41.470 40.465 41.640 44.505 ;
        RECT 45.760 40.465 45.930 44.505 ;
        RECT 41.700 40.080 45.700 40.250 ;
        RECT 46.330 39.740 46.500 45.230 ;
        RECT 47.130 44.720 51.130 44.890 ;
        RECT 46.900 40.465 47.070 44.505 ;
        RECT 51.190 40.465 51.360 44.505 ;
        RECT 47.130 40.080 51.130 40.250 ;
        RECT 51.760 39.740 51.930 45.230 ;
        RECT 40.900 39.570 51.930 39.740 ;
        RECT 52.205 45.245 53.955 45.415 ;
        RECT 52.205 39.755 52.375 45.245 ;
        RECT 52.915 44.735 53.245 44.905 ;
        RECT 52.775 40.480 52.945 44.520 ;
        RECT 53.215 40.480 53.385 44.520 ;
        RECT 52.915 40.095 53.245 40.265 ;
        RECT 53.785 39.755 53.955 45.245 ;
        RECT 52.205 39.585 53.955 39.755 ;
        RECT 54.230 39.760 54.400 49.250 ;
        RECT 54.940 48.740 55.270 48.910 ;
        RECT 54.800 40.485 54.970 48.525 ;
        RECT 55.240 40.485 55.410 48.525 ;
        RECT 54.940 40.100 55.270 40.270 ;
        RECT 55.810 39.760 55.980 49.250 ;
        RECT 57.435 49.260 83.980 49.420 ;
        RECT 57.435 49.235 70.180 49.260 ;
        RECT 57.435 49.005 61.760 49.235 ;
        RECT 54.230 39.590 55.980 39.760 ;
        RECT 57.470 39.745 57.640 49.005 ;
        RECT 58.365 48.435 60.405 48.605 ;
        RECT 57.980 40.375 58.150 48.375 ;
        RECT 60.620 40.375 60.790 48.375 ;
        RECT 58.365 40.145 60.405 40.315 ;
        RECT 61.130 39.745 61.300 49.005 ;
        RECT 57.470 39.575 61.300 39.745 ;
        RECT 61.590 39.745 61.760 49.005 ;
        RECT 62.390 48.725 64.390 48.895 ;
        RECT 62.160 40.470 62.330 48.510 ;
        RECT 64.450 40.470 64.620 48.510 ;
        RECT 62.390 40.085 64.390 40.255 ;
        RECT 65.020 39.745 65.190 49.235 ;
        RECT 65.820 48.725 67.820 48.895 ;
        RECT 65.590 40.470 65.760 48.510 ;
        RECT 67.880 40.470 68.050 48.510 ;
        RECT 68.450 47.665 70.180 49.235 ;
        RECT 82.230 49.250 83.980 49.260 ;
        RECT 68.450 47.495 76.915 47.665 ;
        RECT 68.450 46.085 70.255 47.495 ;
        RECT 70.595 46.625 70.765 46.955 ;
        RECT 70.980 46.925 76.020 47.095 ;
        RECT 70.980 46.485 76.020 46.655 ;
        RECT 76.235 46.625 76.405 46.955 ;
        RECT 76.745 46.085 76.915 47.495 ;
        RECT 68.450 45.915 76.915 46.085 ;
        RECT 68.450 45.400 70.180 45.915 ;
        RECT 68.450 45.285 79.930 45.400 ;
        RECT 65.820 40.085 67.820 40.255 ;
        RECT 68.450 39.745 68.620 45.285 ;
        RECT 61.590 39.575 68.620 39.745 ;
        RECT 68.900 45.230 79.930 45.285 ;
        RECT 68.900 39.740 69.070 45.230 ;
        RECT 69.700 44.720 73.700 44.890 ;
        RECT 69.470 40.465 69.640 44.505 ;
        RECT 73.760 40.465 73.930 44.505 ;
        RECT 69.700 40.080 73.700 40.250 ;
        RECT 74.330 39.740 74.500 45.230 ;
        RECT 75.130 44.720 79.130 44.890 ;
        RECT 74.900 40.465 75.070 44.505 ;
        RECT 79.190 40.465 79.360 44.505 ;
        RECT 75.130 40.080 79.130 40.250 ;
        RECT 79.760 39.740 79.930 45.230 ;
        RECT 68.900 39.570 79.930 39.740 ;
        RECT 80.205 45.245 81.955 45.415 ;
        RECT 80.205 39.755 80.375 45.245 ;
        RECT 80.915 44.735 81.245 44.905 ;
        RECT 80.775 40.480 80.945 44.520 ;
        RECT 81.215 40.480 81.385 44.520 ;
        RECT 80.915 40.095 81.245 40.265 ;
        RECT 81.785 39.755 81.955 45.245 ;
        RECT 80.205 39.585 81.955 39.755 ;
        RECT 82.230 39.760 82.400 49.250 ;
        RECT 82.940 48.740 83.270 48.910 ;
        RECT 82.800 40.485 82.970 48.525 ;
        RECT 83.240 40.485 83.410 48.525 ;
        RECT 82.940 40.100 83.270 40.270 ;
        RECT 83.810 39.760 83.980 49.250 ;
        RECT 85.435 49.260 111.980 49.420 ;
        RECT 85.435 49.235 98.180 49.260 ;
        RECT 85.435 49.005 89.760 49.235 ;
        RECT 82.230 39.590 83.980 39.760 ;
        RECT 85.470 39.745 85.640 49.005 ;
        RECT 86.365 48.435 88.405 48.605 ;
        RECT 85.980 40.375 86.150 48.375 ;
        RECT 88.620 40.375 88.790 48.375 ;
        RECT 86.365 40.145 88.405 40.315 ;
        RECT 89.130 39.745 89.300 49.005 ;
        RECT 85.470 39.575 89.300 39.745 ;
        RECT 89.590 39.745 89.760 49.005 ;
        RECT 90.390 48.725 92.390 48.895 ;
        RECT 90.160 40.470 90.330 48.510 ;
        RECT 92.450 40.470 92.620 48.510 ;
        RECT 90.390 40.085 92.390 40.255 ;
        RECT 93.020 39.745 93.190 49.235 ;
        RECT 93.820 48.725 95.820 48.895 ;
        RECT 93.590 40.470 93.760 48.510 ;
        RECT 95.880 40.470 96.050 48.510 ;
        RECT 96.450 47.665 98.180 49.235 ;
        RECT 110.230 49.250 111.980 49.260 ;
        RECT 96.450 47.495 104.915 47.665 ;
        RECT 96.450 46.085 98.255 47.495 ;
        RECT 98.595 46.625 98.765 46.955 ;
        RECT 98.980 46.925 104.020 47.095 ;
        RECT 98.980 46.485 104.020 46.655 ;
        RECT 104.235 46.625 104.405 46.955 ;
        RECT 104.745 46.085 104.915 47.495 ;
        RECT 96.450 45.915 104.915 46.085 ;
        RECT 96.450 45.400 98.180 45.915 ;
        RECT 96.450 45.285 107.930 45.400 ;
        RECT 93.820 40.085 95.820 40.255 ;
        RECT 96.450 39.745 96.620 45.285 ;
        RECT 89.590 39.575 96.620 39.745 ;
        RECT 96.900 45.230 107.930 45.285 ;
        RECT 96.900 39.740 97.070 45.230 ;
        RECT 97.700 44.720 101.700 44.890 ;
        RECT 97.470 40.465 97.640 44.505 ;
        RECT 101.760 40.465 101.930 44.505 ;
        RECT 97.700 40.080 101.700 40.250 ;
        RECT 102.330 39.740 102.500 45.230 ;
        RECT 103.130 44.720 107.130 44.890 ;
        RECT 102.900 40.465 103.070 44.505 ;
        RECT 107.190 40.465 107.360 44.505 ;
        RECT 103.130 40.080 107.130 40.250 ;
        RECT 107.760 39.740 107.930 45.230 ;
        RECT 96.900 39.570 107.930 39.740 ;
        RECT 108.205 45.245 109.955 45.415 ;
        RECT 108.205 39.755 108.375 45.245 ;
        RECT 108.915 44.735 109.245 44.905 ;
        RECT 108.775 40.480 108.945 44.520 ;
        RECT 109.215 40.480 109.385 44.520 ;
        RECT 108.915 40.095 109.245 40.265 ;
        RECT 109.785 39.755 109.955 45.245 ;
        RECT 108.205 39.585 109.955 39.755 ;
        RECT 110.230 39.760 110.400 49.250 ;
        RECT 110.940 48.740 111.270 48.910 ;
        RECT 110.800 40.485 110.970 48.525 ;
        RECT 111.240 40.485 111.410 48.525 ;
        RECT 110.940 40.100 111.270 40.270 ;
        RECT 111.810 39.760 111.980 49.250 ;
        RECT 113.435 49.260 139.980 49.420 ;
        RECT 113.435 49.235 126.180 49.260 ;
        RECT 113.435 49.005 117.760 49.235 ;
        RECT 110.230 39.590 111.980 39.760 ;
        RECT 113.470 39.745 113.640 49.005 ;
        RECT 114.365 48.435 116.405 48.605 ;
        RECT 113.980 40.375 114.150 48.375 ;
        RECT 116.620 40.375 116.790 48.375 ;
        RECT 114.365 40.145 116.405 40.315 ;
        RECT 117.130 39.745 117.300 49.005 ;
        RECT 113.470 39.575 117.300 39.745 ;
        RECT 117.590 39.745 117.760 49.005 ;
        RECT 118.390 48.725 120.390 48.895 ;
        RECT 118.160 40.470 118.330 48.510 ;
        RECT 120.450 40.470 120.620 48.510 ;
        RECT 118.390 40.085 120.390 40.255 ;
        RECT 121.020 39.745 121.190 49.235 ;
        RECT 121.820 48.725 123.820 48.895 ;
        RECT 121.590 40.470 121.760 48.510 ;
        RECT 123.880 40.470 124.050 48.510 ;
        RECT 124.450 47.665 126.180 49.235 ;
        RECT 138.230 49.250 139.980 49.260 ;
        RECT 124.450 47.495 132.915 47.665 ;
        RECT 124.450 46.085 126.255 47.495 ;
        RECT 126.595 46.625 126.765 46.955 ;
        RECT 126.980 46.925 132.020 47.095 ;
        RECT 126.980 46.485 132.020 46.655 ;
        RECT 132.235 46.625 132.405 46.955 ;
        RECT 132.745 46.085 132.915 47.495 ;
        RECT 124.450 45.915 132.915 46.085 ;
        RECT 124.450 45.400 126.180 45.915 ;
        RECT 124.450 45.285 135.930 45.400 ;
        RECT 121.820 40.085 123.820 40.255 ;
        RECT 124.450 39.745 124.620 45.285 ;
        RECT 117.590 39.575 124.620 39.745 ;
        RECT 124.900 45.230 135.930 45.285 ;
        RECT 124.900 39.740 125.070 45.230 ;
        RECT 125.700 44.720 129.700 44.890 ;
        RECT 125.470 40.465 125.640 44.505 ;
        RECT 129.760 40.465 129.930 44.505 ;
        RECT 125.700 40.080 129.700 40.250 ;
        RECT 130.330 39.740 130.500 45.230 ;
        RECT 131.130 44.720 135.130 44.890 ;
        RECT 130.900 40.465 131.070 44.505 ;
        RECT 135.190 40.465 135.360 44.505 ;
        RECT 131.130 40.080 135.130 40.250 ;
        RECT 135.760 39.740 135.930 45.230 ;
        RECT 124.900 39.570 135.930 39.740 ;
        RECT 136.205 45.245 137.955 45.415 ;
        RECT 136.205 39.755 136.375 45.245 ;
        RECT 136.915 44.735 137.245 44.905 ;
        RECT 136.775 40.480 136.945 44.520 ;
        RECT 137.215 40.480 137.385 44.520 ;
        RECT 136.915 40.095 137.245 40.265 ;
        RECT 137.785 39.755 137.955 45.245 ;
        RECT 136.205 39.585 137.955 39.755 ;
        RECT 138.230 39.760 138.400 49.250 ;
        RECT 138.940 48.740 139.270 48.910 ;
        RECT 138.800 40.485 138.970 48.525 ;
        RECT 139.240 40.485 139.410 48.525 ;
        RECT 138.940 40.100 139.270 40.270 ;
        RECT 139.810 39.760 139.980 49.250 ;
        RECT 143.470 48.190 143.640 49.840 ;
        RECT 144.120 48.670 146.280 49.360 ;
        RECT 146.810 48.670 148.970 49.360 ;
        RECT 149.450 48.190 149.620 49.840 ;
        RECT 143.470 48.020 149.620 48.190 ;
        RECT 143.470 46.370 143.640 48.020 ;
        RECT 144.120 46.850 146.280 47.540 ;
        RECT 146.810 46.850 148.970 47.540 ;
        RECT 149.450 46.370 149.620 48.020 ;
        RECT 143.470 46.200 149.620 46.370 ;
        RECT 143.470 44.550 143.640 46.200 ;
        RECT 144.120 45.030 146.280 45.720 ;
        RECT 146.810 45.030 148.970 45.720 ;
        RECT 149.450 44.550 149.620 46.200 ;
        RECT 143.470 44.380 155.600 44.550 ;
        RECT 143.470 42.730 143.640 44.380 ;
        RECT 144.120 43.210 146.280 43.900 ;
        RECT 146.810 43.210 148.970 43.900 ;
        RECT 149.450 42.730 149.620 44.380 ;
        RECT 150.100 43.210 152.260 43.900 ;
        RECT 152.790 43.210 154.950 43.900 ;
        RECT 155.430 42.730 155.600 44.380 ;
        RECT 143.470 42.560 155.600 42.730 ;
        RECT 143.470 40.910 143.640 42.560 ;
        RECT 144.120 41.390 146.280 42.080 ;
        RECT 146.810 41.390 148.970 42.080 ;
        RECT 149.450 40.910 149.620 42.560 ;
        RECT 150.100 41.390 152.260 42.080 ;
        RECT 152.790 41.390 154.950 42.080 ;
        RECT 155.430 40.910 155.600 42.560 ;
        RECT 143.470 40.740 155.600 40.910 ;
        RECT 150.780 40.250 154.340 40.740 ;
        RECT 138.230 39.590 139.980 39.760 ;
        RECT 2.130 38.665 24.020 38.835 ;
        RECT 2.130 35.265 2.300 38.665 ;
        RECT 2.930 38.155 6.930 38.325 ;
        RECT 2.700 35.945 2.870 37.985 ;
        RECT 6.990 35.945 7.160 37.985 ;
        RECT 2.930 35.605 6.930 35.775 ;
        RECT 7.560 35.265 7.730 38.665 ;
        RECT 8.360 38.155 12.360 38.325 ;
        RECT 8.130 35.945 8.300 37.985 ;
        RECT 12.420 35.945 12.590 37.985 ;
        RECT 8.360 35.605 12.360 35.775 ;
        RECT 12.990 35.265 13.160 38.665 ;
        RECT 13.790 38.155 17.790 38.325 ;
        RECT 13.560 35.945 13.730 37.985 ;
        RECT 17.850 35.945 18.020 37.985 ;
        RECT 13.790 35.605 17.790 35.775 ;
        RECT 18.420 35.265 18.590 38.665 ;
        RECT 19.220 38.155 23.220 38.325 ;
        RECT 18.990 35.945 19.160 37.985 ;
        RECT 23.280 35.945 23.450 37.985 ;
        RECT 23.850 36.240 24.020 38.665 ;
        RECT 24.290 38.670 26.040 38.840 ;
        RECT 24.290 36.270 24.460 38.670 ;
        RECT 25.000 38.160 25.330 38.330 ;
        RECT 24.860 36.950 25.030 37.990 ;
        RECT 25.300 36.950 25.470 37.990 ;
        RECT 25.000 36.610 25.330 36.780 ;
        RECT 25.870 36.270 26.040 38.670 ;
        RECT 24.290 36.240 26.040 36.270 ;
        RECT 26.315 38.675 28.065 38.845 ;
        RECT 26.315 36.240 26.485 38.675 ;
        RECT 27.025 38.165 27.355 38.335 ;
        RECT 19.220 35.605 23.220 35.775 ;
        RECT 23.850 35.275 26.485 36.240 ;
        RECT 26.885 35.955 27.055 37.995 ;
        RECT 27.325 35.955 27.495 37.995 ;
        RECT 27.025 35.615 27.355 35.785 ;
        RECT 27.895 35.275 28.065 38.675 ;
        RECT 23.850 35.265 28.065 35.275 ;
        RECT 2.130 35.245 28.065 35.265 ;
        RECT 30.130 38.665 52.020 38.835 ;
        RECT 30.130 35.265 30.300 38.665 ;
        RECT 30.930 38.155 34.930 38.325 ;
        RECT 30.700 35.945 30.870 37.985 ;
        RECT 34.990 35.945 35.160 37.985 ;
        RECT 30.930 35.605 34.930 35.775 ;
        RECT 35.560 35.265 35.730 38.665 ;
        RECT 36.360 38.155 40.360 38.325 ;
        RECT 36.130 35.945 36.300 37.985 ;
        RECT 40.420 35.945 40.590 37.985 ;
        RECT 36.360 35.605 40.360 35.775 ;
        RECT 40.990 35.265 41.160 38.665 ;
        RECT 41.790 38.155 45.790 38.325 ;
        RECT 41.560 35.945 41.730 37.985 ;
        RECT 45.850 35.945 46.020 37.985 ;
        RECT 41.790 35.605 45.790 35.775 ;
        RECT 46.420 35.265 46.590 38.665 ;
        RECT 47.220 38.155 51.220 38.325 ;
        RECT 46.990 35.945 47.160 37.985 ;
        RECT 51.280 35.945 51.450 37.985 ;
        RECT 51.850 36.240 52.020 38.665 ;
        RECT 52.290 38.670 54.040 38.840 ;
        RECT 52.290 36.270 52.460 38.670 ;
        RECT 53.000 38.160 53.330 38.330 ;
        RECT 52.860 36.950 53.030 37.990 ;
        RECT 53.300 36.950 53.470 37.990 ;
        RECT 53.000 36.610 53.330 36.780 ;
        RECT 53.870 36.270 54.040 38.670 ;
        RECT 52.290 36.240 54.040 36.270 ;
        RECT 54.315 38.675 56.065 38.845 ;
        RECT 54.315 36.240 54.485 38.675 ;
        RECT 55.025 38.165 55.355 38.335 ;
        RECT 47.220 35.605 51.220 35.775 ;
        RECT 51.850 35.275 54.485 36.240 ;
        RECT 54.885 35.955 55.055 37.995 ;
        RECT 55.325 35.955 55.495 37.995 ;
        RECT 55.025 35.615 55.355 35.785 ;
        RECT 55.895 35.275 56.065 38.675 ;
        RECT 51.850 35.265 56.065 35.275 ;
        RECT 30.130 35.245 56.065 35.265 ;
        RECT 58.130 38.665 80.020 38.835 ;
        RECT 58.130 35.265 58.300 38.665 ;
        RECT 58.930 38.155 62.930 38.325 ;
        RECT 58.700 35.945 58.870 37.985 ;
        RECT 62.990 35.945 63.160 37.985 ;
        RECT 58.930 35.605 62.930 35.775 ;
        RECT 63.560 35.265 63.730 38.665 ;
        RECT 64.360 38.155 68.360 38.325 ;
        RECT 64.130 35.945 64.300 37.985 ;
        RECT 68.420 35.945 68.590 37.985 ;
        RECT 64.360 35.605 68.360 35.775 ;
        RECT 68.990 35.265 69.160 38.665 ;
        RECT 69.790 38.155 73.790 38.325 ;
        RECT 69.560 35.945 69.730 37.985 ;
        RECT 73.850 35.945 74.020 37.985 ;
        RECT 69.790 35.605 73.790 35.775 ;
        RECT 74.420 35.265 74.590 38.665 ;
        RECT 75.220 38.155 79.220 38.325 ;
        RECT 74.990 35.945 75.160 37.985 ;
        RECT 79.280 35.945 79.450 37.985 ;
        RECT 79.850 36.240 80.020 38.665 ;
        RECT 80.290 38.670 82.040 38.840 ;
        RECT 80.290 36.270 80.460 38.670 ;
        RECT 81.000 38.160 81.330 38.330 ;
        RECT 80.860 36.950 81.030 37.990 ;
        RECT 81.300 36.950 81.470 37.990 ;
        RECT 81.000 36.610 81.330 36.780 ;
        RECT 81.870 36.270 82.040 38.670 ;
        RECT 80.290 36.240 82.040 36.270 ;
        RECT 82.315 38.675 84.065 38.845 ;
        RECT 82.315 36.240 82.485 38.675 ;
        RECT 83.025 38.165 83.355 38.335 ;
        RECT 75.220 35.605 79.220 35.775 ;
        RECT 79.850 35.275 82.485 36.240 ;
        RECT 82.885 35.955 83.055 37.995 ;
        RECT 83.325 35.955 83.495 37.995 ;
        RECT 83.025 35.615 83.355 35.785 ;
        RECT 83.895 35.275 84.065 38.675 ;
        RECT 79.850 35.265 84.065 35.275 ;
        RECT 58.130 35.245 84.065 35.265 ;
        RECT 86.130 38.665 108.020 38.835 ;
        RECT 86.130 35.265 86.300 38.665 ;
        RECT 86.930 38.155 90.930 38.325 ;
        RECT 86.700 35.945 86.870 37.985 ;
        RECT 90.990 35.945 91.160 37.985 ;
        RECT 86.930 35.605 90.930 35.775 ;
        RECT 91.560 35.265 91.730 38.665 ;
        RECT 92.360 38.155 96.360 38.325 ;
        RECT 92.130 35.945 92.300 37.985 ;
        RECT 96.420 35.945 96.590 37.985 ;
        RECT 92.360 35.605 96.360 35.775 ;
        RECT 96.990 35.265 97.160 38.665 ;
        RECT 97.790 38.155 101.790 38.325 ;
        RECT 97.560 35.945 97.730 37.985 ;
        RECT 101.850 35.945 102.020 37.985 ;
        RECT 97.790 35.605 101.790 35.775 ;
        RECT 102.420 35.265 102.590 38.665 ;
        RECT 103.220 38.155 107.220 38.325 ;
        RECT 102.990 35.945 103.160 37.985 ;
        RECT 107.280 35.945 107.450 37.985 ;
        RECT 107.850 36.240 108.020 38.665 ;
        RECT 108.290 38.670 110.040 38.840 ;
        RECT 108.290 36.270 108.460 38.670 ;
        RECT 109.000 38.160 109.330 38.330 ;
        RECT 108.860 36.950 109.030 37.990 ;
        RECT 109.300 36.950 109.470 37.990 ;
        RECT 109.000 36.610 109.330 36.780 ;
        RECT 109.870 36.270 110.040 38.670 ;
        RECT 108.290 36.240 110.040 36.270 ;
        RECT 110.315 38.675 112.065 38.845 ;
        RECT 110.315 36.240 110.485 38.675 ;
        RECT 111.025 38.165 111.355 38.335 ;
        RECT 103.220 35.605 107.220 35.775 ;
        RECT 107.850 35.275 110.485 36.240 ;
        RECT 110.885 35.955 111.055 37.995 ;
        RECT 111.325 35.955 111.495 37.995 ;
        RECT 111.025 35.615 111.355 35.785 ;
        RECT 111.895 35.275 112.065 38.675 ;
        RECT 107.850 35.265 112.065 35.275 ;
        RECT 86.130 35.245 112.065 35.265 ;
        RECT 114.130 38.665 136.020 38.835 ;
        RECT 114.130 35.265 114.300 38.665 ;
        RECT 114.930 38.155 118.930 38.325 ;
        RECT 114.700 35.945 114.870 37.985 ;
        RECT 118.990 35.945 119.160 37.985 ;
        RECT 114.930 35.605 118.930 35.775 ;
        RECT 119.560 35.265 119.730 38.665 ;
        RECT 120.360 38.155 124.360 38.325 ;
        RECT 120.130 35.945 120.300 37.985 ;
        RECT 124.420 35.945 124.590 37.985 ;
        RECT 120.360 35.605 124.360 35.775 ;
        RECT 124.990 35.265 125.160 38.665 ;
        RECT 125.790 38.155 129.790 38.325 ;
        RECT 125.560 35.945 125.730 37.985 ;
        RECT 129.850 35.945 130.020 37.985 ;
        RECT 125.790 35.605 129.790 35.775 ;
        RECT 130.420 35.265 130.590 38.665 ;
        RECT 131.220 38.155 135.220 38.325 ;
        RECT 130.990 35.945 131.160 37.985 ;
        RECT 135.280 35.945 135.450 37.985 ;
        RECT 135.850 36.240 136.020 38.665 ;
        RECT 136.290 38.670 138.040 38.840 ;
        RECT 136.290 36.270 136.460 38.670 ;
        RECT 137.000 38.160 137.330 38.330 ;
        RECT 136.860 36.950 137.030 37.990 ;
        RECT 137.300 36.950 137.470 37.990 ;
        RECT 137.000 36.610 137.330 36.780 ;
        RECT 137.870 36.270 138.040 38.670 ;
        RECT 136.290 36.240 138.040 36.270 ;
        RECT 138.315 38.675 140.065 38.845 ;
        RECT 138.315 36.240 138.485 38.675 ;
        RECT 139.025 38.165 139.355 38.335 ;
        RECT 131.220 35.605 135.220 35.775 ;
        RECT 135.850 35.275 138.485 36.240 ;
        RECT 138.885 35.955 139.055 37.995 ;
        RECT 139.325 35.955 139.495 37.995 ;
        RECT 139.025 35.615 139.355 35.785 ;
        RECT 139.895 35.275 140.065 38.675 ;
        RECT 135.850 35.265 140.065 35.275 ;
        RECT 114.130 35.245 140.065 35.265 ;
        RECT 1.475 35.105 28.065 35.245 ;
        RECT 29.475 35.105 56.065 35.245 ;
        RECT 57.475 35.105 84.065 35.245 ;
        RECT 85.475 35.105 112.065 35.245 ;
        RECT 113.475 35.105 140.065 35.245 ;
        RECT 1.475 34.380 28.055 35.105 ;
        RECT 29.475 34.380 56.055 35.105 ;
        RECT 57.475 34.380 84.055 35.105 ;
        RECT 85.475 34.380 112.055 35.105 ;
        RECT 113.475 34.380 140.055 35.105 ;
        RECT 1.450 33.480 27.925 33.960 ;
        RECT 29.450 33.480 55.925 33.960 ;
        RECT 57.450 33.480 83.925 33.960 ;
        RECT 85.450 33.480 111.925 33.960 ;
        RECT 113.450 33.480 139.925 33.960 ;
        RECT 1.435 33.420 27.925 33.480 ;
        RECT 29.435 33.420 55.925 33.480 ;
        RECT 57.435 33.420 83.925 33.480 ;
        RECT 85.435 33.420 111.925 33.480 ;
        RECT 113.435 33.420 139.925 33.480 ;
        RECT 1.435 33.260 27.980 33.420 ;
        RECT 1.435 33.235 14.180 33.260 ;
        RECT 1.435 33.005 5.760 33.235 ;
        RECT 1.470 23.745 1.640 33.005 ;
        RECT 2.365 32.435 4.405 32.605 ;
        RECT 1.980 24.375 2.150 32.375 ;
        RECT 4.620 24.375 4.790 32.375 ;
        RECT 2.365 24.145 4.405 24.315 ;
        RECT 5.130 23.745 5.300 33.005 ;
        RECT 1.470 23.575 5.300 23.745 ;
        RECT 5.590 23.745 5.760 33.005 ;
        RECT 6.390 32.725 8.390 32.895 ;
        RECT 6.160 24.470 6.330 32.510 ;
        RECT 8.450 24.470 8.620 32.510 ;
        RECT 6.390 24.085 8.390 24.255 ;
        RECT 9.020 23.745 9.190 33.235 ;
        RECT 9.820 32.725 11.820 32.895 ;
        RECT 9.590 24.470 9.760 32.510 ;
        RECT 11.880 24.470 12.050 32.510 ;
        RECT 12.450 31.665 14.180 33.235 ;
        RECT 26.230 33.250 27.980 33.260 ;
        RECT 12.450 31.495 20.915 31.665 ;
        RECT 12.450 30.085 14.255 31.495 ;
        RECT 14.595 30.625 14.765 30.955 ;
        RECT 14.980 30.925 20.020 31.095 ;
        RECT 14.980 30.485 20.020 30.655 ;
        RECT 20.235 30.625 20.405 30.955 ;
        RECT 20.745 30.085 20.915 31.495 ;
        RECT 12.450 29.915 20.915 30.085 ;
        RECT 12.450 29.400 14.180 29.915 ;
        RECT 12.450 29.285 23.930 29.400 ;
        RECT 9.820 24.085 11.820 24.255 ;
        RECT 12.450 23.745 12.620 29.285 ;
        RECT 5.590 23.575 12.620 23.745 ;
        RECT 12.900 29.230 23.930 29.285 ;
        RECT 12.900 23.740 13.070 29.230 ;
        RECT 13.700 28.720 17.700 28.890 ;
        RECT 13.470 24.465 13.640 28.505 ;
        RECT 17.760 24.465 17.930 28.505 ;
        RECT 13.700 24.080 17.700 24.250 ;
        RECT 18.330 23.740 18.500 29.230 ;
        RECT 19.130 28.720 23.130 28.890 ;
        RECT 18.900 24.465 19.070 28.505 ;
        RECT 23.190 24.465 23.360 28.505 ;
        RECT 19.130 24.080 23.130 24.250 ;
        RECT 23.760 23.740 23.930 29.230 ;
        RECT 12.900 23.570 23.930 23.740 ;
        RECT 24.205 29.245 25.955 29.415 ;
        RECT 24.205 23.755 24.375 29.245 ;
        RECT 24.915 28.735 25.245 28.905 ;
        RECT 24.775 24.480 24.945 28.520 ;
        RECT 25.215 24.480 25.385 28.520 ;
        RECT 24.915 24.095 25.245 24.265 ;
        RECT 25.785 23.755 25.955 29.245 ;
        RECT 24.205 23.585 25.955 23.755 ;
        RECT 26.230 23.760 26.400 33.250 ;
        RECT 26.940 32.740 27.270 32.910 ;
        RECT 26.800 24.485 26.970 32.525 ;
        RECT 27.240 24.485 27.410 32.525 ;
        RECT 26.940 24.100 27.270 24.270 ;
        RECT 27.810 23.760 27.980 33.250 ;
        RECT 29.435 33.260 55.980 33.420 ;
        RECT 29.435 33.235 42.180 33.260 ;
        RECT 29.435 33.005 33.760 33.235 ;
        RECT 26.230 23.590 27.980 23.760 ;
        RECT 29.470 23.745 29.640 33.005 ;
        RECT 30.365 32.435 32.405 32.605 ;
        RECT 29.980 24.375 30.150 32.375 ;
        RECT 32.620 24.375 32.790 32.375 ;
        RECT 30.365 24.145 32.405 24.315 ;
        RECT 33.130 23.745 33.300 33.005 ;
        RECT 29.470 23.575 33.300 23.745 ;
        RECT 33.590 23.745 33.760 33.005 ;
        RECT 34.390 32.725 36.390 32.895 ;
        RECT 34.160 24.470 34.330 32.510 ;
        RECT 36.450 24.470 36.620 32.510 ;
        RECT 34.390 24.085 36.390 24.255 ;
        RECT 37.020 23.745 37.190 33.235 ;
        RECT 37.820 32.725 39.820 32.895 ;
        RECT 37.590 24.470 37.760 32.510 ;
        RECT 39.880 24.470 40.050 32.510 ;
        RECT 40.450 31.665 42.180 33.235 ;
        RECT 54.230 33.250 55.980 33.260 ;
        RECT 40.450 31.495 48.915 31.665 ;
        RECT 40.450 30.085 42.255 31.495 ;
        RECT 42.595 30.625 42.765 30.955 ;
        RECT 42.980 30.925 48.020 31.095 ;
        RECT 42.980 30.485 48.020 30.655 ;
        RECT 48.235 30.625 48.405 30.955 ;
        RECT 48.745 30.085 48.915 31.495 ;
        RECT 40.450 29.915 48.915 30.085 ;
        RECT 40.450 29.400 42.180 29.915 ;
        RECT 40.450 29.285 51.930 29.400 ;
        RECT 37.820 24.085 39.820 24.255 ;
        RECT 40.450 23.745 40.620 29.285 ;
        RECT 33.590 23.575 40.620 23.745 ;
        RECT 40.900 29.230 51.930 29.285 ;
        RECT 40.900 23.740 41.070 29.230 ;
        RECT 41.700 28.720 45.700 28.890 ;
        RECT 41.470 24.465 41.640 28.505 ;
        RECT 45.760 24.465 45.930 28.505 ;
        RECT 41.700 24.080 45.700 24.250 ;
        RECT 46.330 23.740 46.500 29.230 ;
        RECT 47.130 28.720 51.130 28.890 ;
        RECT 46.900 24.465 47.070 28.505 ;
        RECT 51.190 24.465 51.360 28.505 ;
        RECT 47.130 24.080 51.130 24.250 ;
        RECT 51.760 23.740 51.930 29.230 ;
        RECT 40.900 23.570 51.930 23.740 ;
        RECT 52.205 29.245 53.955 29.415 ;
        RECT 52.205 23.755 52.375 29.245 ;
        RECT 52.915 28.735 53.245 28.905 ;
        RECT 52.775 24.480 52.945 28.520 ;
        RECT 53.215 24.480 53.385 28.520 ;
        RECT 52.915 24.095 53.245 24.265 ;
        RECT 53.785 23.755 53.955 29.245 ;
        RECT 52.205 23.585 53.955 23.755 ;
        RECT 54.230 23.760 54.400 33.250 ;
        RECT 54.940 32.740 55.270 32.910 ;
        RECT 54.800 24.485 54.970 32.525 ;
        RECT 55.240 24.485 55.410 32.525 ;
        RECT 54.940 24.100 55.270 24.270 ;
        RECT 55.810 23.760 55.980 33.250 ;
        RECT 57.435 33.260 83.980 33.420 ;
        RECT 57.435 33.235 70.180 33.260 ;
        RECT 57.435 33.005 61.760 33.235 ;
        RECT 54.230 23.590 55.980 23.760 ;
        RECT 57.470 23.745 57.640 33.005 ;
        RECT 58.365 32.435 60.405 32.605 ;
        RECT 57.980 24.375 58.150 32.375 ;
        RECT 60.620 24.375 60.790 32.375 ;
        RECT 58.365 24.145 60.405 24.315 ;
        RECT 61.130 23.745 61.300 33.005 ;
        RECT 57.470 23.575 61.300 23.745 ;
        RECT 61.590 23.745 61.760 33.005 ;
        RECT 62.390 32.725 64.390 32.895 ;
        RECT 62.160 24.470 62.330 32.510 ;
        RECT 64.450 24.470 64.620 32.510 ;
        RECT 62.390 24.085 64.390 24.255 ;
        RECT 65.020 23.745 65.190 33.235 ;
        RECT 65.820 32.725 67.820 32.895 ;
        RECT 65.590 24.470 65.760 32.510 ;
        RECT 67.880 24.470 68.050 32.510 ;
        RECT 68.450 31.665 70.180 33.235 ;
        RECT 82.230 33.250 83.980 33.260 ;
        RECT 68.450 31.495 76.915 31.665 ;
        RECT 68.450 30.085 70.255 31.495 ;
        RECT 70.595 30.625 70.765 30.955 ;
        RECT 70.980 30.925 76.020 31.095 ;
        RECT 70.980 30.485 76.020 30.655 ;
        RECT 76.235 30.625 76.405 30.955 ;
        RECT 76.745 30.085 76.915 31.495 ;
        RECT 68.450 29.915 76.915 30.085 ;
        RECT 68.450 29.400 70.180 29.915 ;
        RECT 68.450 29.285 79.930 29.400 ;
        RECT 65.820 24.085 67.820 24.255 ;
        RECT 68.450 23.745 68.620 29.285 ;
        RECT 61.590 23.575 68.620 23.745 ;
        RECT 68.900 29.230 79.930 29.285 ;
        RECT 68.900 23.740 69.070 29.230 ;
        RECT 69.700 28.720 73.700 28.890 ;
        RECT 69.470 24.465 69.640 28.505 ;
        RECT 73.760 24.465 73.930 28.505 ;
        RECT 69.700 24.080 73.700 24.250 ;
        RECT 74.330 23.740 74.500 29.230 ;
        RECT 75.130 28.720 79.130 28.890 ;
        RECT 74.900 24.465 75.070 28.505 ;
        RECT 79.190 24.465 79.360 28.505 ;
        RECT 75.130 24.080 79.130 24.250 ;
        RECT 79.760 23.740 79.930 29.230 ;
        RECT 68.900 23.570 79.930 23.740 ;
        RECT 80.205 29.245 81.955 29.415 ;
        RECT 80.205 23.755 80.375 29.245 ;
        RECT 80.915 28.735 81.245 28.905 ;
        RECT 80.775 24.480 80.945 28.520 ;
        RECT 81.215 24.480 81.385 28.520 ;
        RECT 80.915 24.095 81.245 24.265 ;
        RECT 81.785 23.755 81.955 29.245 ;
        RECT 80.205 23.585 81.955 23.755 ;
        RECT 82.230 23.760 82.400 33.250 ;
        RECT 82.940 32.740 83.270 32.910 ;
        RECT 82.800 24.485 82.970 32.525 ;
        RECT 83.240 24.485 83.410 32.525 ;
        RECT 82.940 24.100 83.270 24.270 ;
        RECT 83.810 23.760 83.980 33.250 ;
        RECT 85.435 33.260 111.980 33.420 ;
        RECT 85.435 33.235 98.180 33.260 ;
        RECT 85.435 33.005 89.760 33.235 ;
        RECT 82.230 23.590 83.980 23.760 ;
        RECT 85.470 23.745 85.640 33.005 ;
        RECT 86.365 32.435 88.405 32.605 ;
        RECT 85.980 24.375 86.150 32.375 ;
        RECT 88.620 24.375 88.790 32.375 ;
        RECT 86.365 24.145 88.405 24.315 ;
        RECT 89.130 23.745 89.300 33.005 ;
        RECT 85.470 23.575 89.300 23.745 ;
        RECT 89.590 23.745 89.760 33.005 ;
        RECT 90.390 32.725 92.390 32.895 ;
        RECT 90.160 24.470 90.330 32.510 ;
        RECT 92.450 24.470 92.620 32.510 ;
        RECT 90.390 24.085 92.390 24.255 ;
        RECT 93.020 23.745 93.190 33.235 ;
        RECT 93.820 32.725 95.820 32.895 ;
        RECT 93.590 24.470 93.760 32.510 ;
        RECT 95.880 24.470 96.050 32.510 ;
        RECT 96.450 31.665 98.180 33.235 ;
        RECT 110.230 33.250 111.980 33.260 ;
        RECT 96.450 31.495 104.915 31.665 ;
        RECT 96.450 30.085 98.255 31.495 ;
        RECT 98.595 30.625 98.765 30.955 ;
        RECT 98.980 30.925 104.020 31.095 ;
        RECT 98.980 30.485 104.020 30.655 ;
        RECT 104.235 30.625 104.405 30.955 ;
        RECT 104.745 30.085 104.915 31.495 ;
        RECT 96.450 29.915 104.915 30.085 ;
        RECT 96.450 29.400 98.180 29.915 ;
        RECT 96.450 29.285 107.930 29.400 ;
        RECT 93.820 24.085 95.820 24.255 ;
        RECT 96.450 23.745 96.620 29.285 ;
        RECT 89.590 23.575 96.620 23.745 ;
        RECT 96.900 29.230 107.930 29.285 ;
        RECT 96.900 23.740 97.070 29.230 ;
        RECT 97.700 28.720 101.700 28.890 ;
        RECT 97.470 24.465 97.640 28.505 ;
        RECT 101.760 24.465 101.930 28.505 ;
        RECT 97.700 24.080 101.700 24.250 ;
        RECT 102.330 23.740 102.500 29.230 ;
        RECT 103.130 28.720 107.130 28.890 ;
        RECT 102.900 24.465 103.070 28.505 ;
        RECT 107.190 24.465 107.360 28.505 ;
        RECT 103.130 24.080 107.130 24.250 ;
        RECT 107.760 23.740 107.930 29.230 ;
        RECT 96.900 23.570 107.930 23.740 ;
        RECT 108.205 29.245 109.955 29.415 ;
        RECT 108.205 23.755 108.375 29.245 ;
        RECT 108.915 28.735 109.245 28.905 ;
        RECT 108.775 24.480 108.945 28.520 ;
        RECT 109.215 24.480 109.385 28.520 ;
        RECT 108.915 24.095 109.245 24.265 ;
        RECT 109.785 23.755 109.955 29.245 ;
        RECT 108.205 23.585 109.955 23.755 ;
        RECT 110.230 23.760 110.400 33.250 ;
        RECT 110.940 32.740 111.270 32.910 ;
        RECT 110.800 24.485 110.970 32.525 ;
        RECT 111.240 24.485 111.410 32.525 ;
        RECT 110.940 24.100 111.270 24.270 ;
        RECT 111.810 23.760 111.980 33.250 ;
        RECT 113.435 33.260 139.980 33.420 ;
        RECT 113.435 33.235 126.180 33.260 ;
        RECT 113.435 33.005 117.760 33.235 ;
        RECT 110.230 23.590 111.980 23.760 ;
        RECT 113.470 23.745 113.640 33.005 ;
        RECT 114.365 32.435 116.405 32.605 ;
        RECT 113.980 24.375 114.150 32.375 ;
        RECT 116.620 24.375 116.790 32.375 ;
        RECT 114.365 24.145 116.405 24.315 ;
        RECT 117.130 23.745 117.300 33.005 ;
        RECT 113.470 23.575 117.300 23.745 ;
        RECT 117.590 23.745 117.760 33.005 ;
        RECT 118.390 32.725 120.390 32.895 ;
        RECT 118.160 24.470 118.330 32.510 ;
        RECT 120.450 24.470 120.620 32.510 ;
        RECT 118.390 24.085 120.390 24.255 ;
        RECT 121.020 23.745 121.190 33.235 ;
        RECT 121.820 32.725 123.820 32.895 ;
        RECT 121.590 24.470 121.760 32.510 ;
        RECT 123.880 24.470 124.050 32.510 ;
        RECT 124.450 31.665 126.180 33.235 ;
        RECT 138.230 33.250 139.980 33.260 ;
        RECT 124.450 31.495 132.915 31.665 ;
        RECT 124.450 30.085 126.255 31.495 ;
        RECT 126.595 30.625 126.765 30.955 ;
        RECT 126.980 30.925 132.020 31.095 ;
        RECT 126.980 30.485 132.020 30.655 ;
        RECT 132.235 30.625 132.405 30.955 ;
        RECT 132.745 30.085 132.915 31.495 ;
        RECT 124.450 29.915 132.915 30.085 ;
        RECT 124.450 29.400 126.180 29.915 ;
        RECT 124.450 29.285 135.930 29.400 ;
        RECT 121.820 24.085 123.820 24.255 ;
        RECT 124.450 23.745 124.620 29.285 ;
        RECT 117.590 23.575 124.620 23.745 ;
        RECT 124.900 29.230 135.930 29.285 ;
        RECT 124.900 23.740 125.070 29.230 ;
        RECT 125.700 28.720 129.700 28.890 ;
        RECT 125.470 24.465 125.640 28.505 ;
        RECT 129.760 24.465 129.930 28.505 ;
        RECT 125.700 24.080 129.700 24.250 ;
        RECT 130.330 23.740 130.500 29.230 ;
        RECT 131.130 28.720 135.130 28.890 ;
        RECT 130.900 24.465 131.070 28.505 ;
        RECT 135.190 24.465 135.360 28.505 ;
        RECT 131.130 24.080 135.130 24.250 ;
        RECT 135.760 23.740 135.930 29.230 ;
        RECT 124.900 23.570 135.930 23.740 ;
        RECT 136.205 29.245 137.955 29.415 ;
        RECT 136.205 23.755 136.375 29.245 ;
        RECT 136.915 28.735 137.245 28.905 ;
        RECT 136.775 24.480 136.945 28.520 ;
        RECT 137.215 24.480 137.385 28.520 ;
        RECT 136.915 24.095 137.245 24.265 ;
        RECT 137.785 23.755 137.955 29.245 ;
        RECT 136.205 23.585 137.955 23.755 ;
        RECT 138.230 23.760 138.400 33.250 ;
        RECT 138.940 32.740 139.270 32.910 ;
        RECT 138.800 24.485 138.970 32.525 ;
        RECT 139.240 24.485 139.410 32.525 ;
        RECT 138.940 24.100 139.270 24.270 ;
        RECT 139.810 23.760 139.980 33.250 ;
        RECT 138.230 23.590 139.980 23.760 ;
        RECT 2.130 22.665 24.020 22.835 ;
        RECT 2.130 19.265 2.300 22.665 ;
        RECT 2.930 22.155 6.930 22.325 ;
        RECT 2.700 19.945 2.870 21.985 ;
        RECT 6.990 19.945 7.160 21.985 ;
        RECT 2.930 19.605 6.930 19.775 ;
        RECT 7.560 19.265 7.730 22.665 ;
        RECT 8.360 22.155 12.360 22.325 ;
        RECT 8.130 19.945 8.300 21.985 ;
        RECT 12.420 19.945 12.590 21.985 ;
        RECT 8.360 19.605 12.360 19.775 ;
        RECT 12.990 19.265 13.160 22.665 ;
        RECT 13.790 22.155 17.790 22.325 ;
        RECT 13.560 19.945 13.730 21.985 ;
        RECT 17.850 19.945 18.020 21.985 ;
        RECT 13.790 19.605 17.790 19.775 ;
        RECT 18.420 19.265 18.590 22.665 ;
        RECT 19.220 22.155 23.220 22.325 ;
        RECT 18.990 19.945 19.160 21.985 ;
        RECT 23.280 19.945 23.450 21.985 ;
        RECT 23.850 20.240 24.020 22.665 ;
        RECT 24.290 22.670 26.040 22.840 ;
        RECT 24.290 20.270 24.460 22.670 ;
        RECT 25.000 22.160 25.330 22.330 ;
        RECT 24.860 20.950 25.030 21.990 ;
        RECT 25.300 20.950 25.470 21.990 ;
        RECT 25.000 20.610 25.330 20.780 ;
        RECT 25.870 20.270 26.040 22.670 ;
        RECT 24.290 20.240 26.040 20.270 ;
        RECT 26.315 22.675 28.065 22.845 ;
        RECT 26.315 20.240 26.485 22.675 ;
        RECT 27.025 22.165 27.355 22.335 ;
        RECT 19.220 19.605 23.220 19.775 ;
        RECT 23.850 19.275 26.485 20.240 ;
        RECT 26.885 19.955 27.055 21.995 ;
        RECT 27.325 19.955 27.495 21.995 ;
        RECT 27.025 19.615 27.355 19.785 ;
        RECT 27.895 19.275 28.065 22.675 ;
        RECT 23.850 19.265 28.065 19.275 ;
        RECT 2.130 19.245 28.065 19.265 ;
        RECT 30.130 22.665 52.020 22.835 ;
        RECT 30.130 19.265 30.300 22.665 ;
        RECT 30.930 22.155 34.930 22.325 ;
        RECT 30.700 19.945 30.870 21.985 ;
        RECT 34.990 19.945 35.160 21.985 ;
        RECT 30.930 19.605 34.930 19.775 ;
        RECT 35.560 19.265 35.730 22.665 ;
        RECT 36.360 22.155 40.360 22.325 ;
        RECT 36.130 19.945 36.300 21.985 ;
        RECT 40.420 19.945 40.590 21.985 ;
        RECT 36.360 19.605 40.360 19.775 ;
        RECT 40.990 19.265 41.160 22.665 ;
        RECT 41.790 22.155 45.790 22.325 ;
        RECT 41.560 19.945 41.730 21.985 ;
        RECT 45.850 19.945 46.020 21.985 ;
        RECT 41.790 19.605 45.790 19.775 ;
        RECT 46.420 19.265 46.590 22.665 ;
        RECT 47.220 22.155 51.220 22.325 ;
        RECT 46.990 19.945 47.160 21.985 ;
        RECT 51.280 19.945 51.450 21.985 ;
        RECT 51.850 20.240 52.020 22.665 ;
        RECT 52.290 22.670 54.040 22.840 ;
        RECT 52.290 20.270 52.460 22.670 ;
        RECT 53.000 22.160 53.330 22.330 ;
        RECT 52.860 20.950 53.030 21.990 ;
        RECT 53.300 20.950 53.470 21.990 ;
        RECT 53.000 20.610 53.330 20.780 ;
        RECT 53.870 20.270 54.040 22.670 ;
        RECT 52.290 20.240 54.040 20.270 ;
        RECT 54.315 22.675 56.065 22.845 ;
        RECT 54.315 20.240 54.485 22.675 ;
        RECT 55.025 22.165 55.355 22.335 ;
        RECT 47.220 19.605 51.220 19.775 ;
        RECT 51.850 19.275 54.485 20.240 ;
        RECT 54.885 19.955 55.055 21.995 ;
        RECT 55.325 19.955 55.495 21.995 ;
        RECT 55.025 19.615 55.355 19.785 ;
        RECT 55.895 19.275 56.065 22.675 ;
        RECT 51.850 19.265 56.065 19.275 ;
        RECT 30.130 19.245 56.065 19.265 ;
        RECT 58.130 22.665 80.020 22.835 ;
        RECT 58.130 19.265 58.300 22.665 ;
        RECT 58.930 22.155 62.930 22.325 ;
        RECT 58.700 19.945 58.870 21.985 ;
        RECT 62.990 19.945 63.160 21.985 ;
        RECT 58.930 19.605 62.930 19.775 ;
        RECT 63.560 19.265 63.730 22.665 ;
        RECT 64.360 22.155 68.360 22.325 ;
        RECT 64.130 19.945 64.300 21.985 ;
        RECT 68.420 19.945 68.590 21.985 ;
        RECT 64.360 19.605 68.360 19.775 ;
        RECT 68.990 19.265 69.160 22.665 ;
        RECT 69.790 22.155 73.790 22.325 ;
        RECT 69.560 19.945 69.730 21.985 ;
        RECT 73.850 19.945 74.020 21.985 ;
        RECT 69.790 19.605 73.790 19.775 ;
        RECT 74.420 19.265 74.590 22.665 ;
        RECT 75.220 22.155 79.220 22.325 ;
        RECT 74.990 19.945 75.160 21.985 ;
        RECT 79.280 19.945 79.450 21.985 ;
        RECT 79.850 20.240 80.020 22.665 ;
        RECT 80.290 22.670 82.040 22.840 ;
        RECT 80.290 20.270 80.460 22.670 ;
        RECT 81.000 22.160 81.330 22.330 ;
        RECT 80.860 20.950 81.030 21.990 ;
        RECT 81.300 20.950 81.470 21.990 ;
        RECT 81.000 20.610 81.330 20.780 ;
        RECT 81.870 20.270 82.040 22.670 ;
        RECT 80.290 20.240 82.040 20.270 ;
        RECT 82.315 22.675 84.065 22.845 ;
        RECT 82.315 20.240 82.485 22.675 ;
        RECT 83.025 22.165 83.355 22.335 ;
        RECT 75.220 19.605 79.220 19.775 ;
        RECT 79.850 19.275 82.485 20.240 ;
        RECT 82.885 19.955 83.055 21.995 ;
        RECT 83.325 19.955 83.495 21.995 ;
        RECT 83.025 19.615 83.355 19.785 ;
        RECT 83.895 19.275 84.065 22.675 ;
        RECT 79.850 19.265 84.065 19.275 ;
        RECT 58.130 19.245 84.065 19.265 ;
        RECT 86.130 22.665 108.020 22.835 ;
        RECT 86.130 19.265 86.300 22.665 ;
        RECT 86.930 22.155 90.930 22.325 ;
        RECT 86.700 19.945 86.870 21.985 ;
        RECT 90.990 19.945 91.160 21.985 ;
        RECT 86.930 19.605 90.930 19.775 ;
        RECT 91.560 19.265 91.730 22.665 ;
        RECT 92.360 22.155 96.360 22.325 ;
        RECT 92.130 19.945 92.300 21.985 ;
        RECT 96.420 19.945 96.590 21.985 ;
        RECT 92.360 19.605 96.360 19.775 ;
        RECT 96.990 19.265 97.160 22.665 ;
        RECT 97.790 22.155 101.790 22.325 ;
        RECT 97.560 19.945 97.730 21.985 ;
        RECT 101.850 19.945 102.020 21.985 ;
        RECT 97.790 19.605 101.790 19.775 ;
        RECT 102.420 19.265 102.590 22.665 ;
        RECT 103.220 22.155 107.220 22.325 ;
        RECT 102.990 19.945 103.160 21.985 ;
        RECT 107.280 19.945 107.450 21.985 ;
        RECT 107.850 20.240 108.020 22.665 ;
        RECT 108.290 22.670 110.040 22.840 ;
        RECT 108.290 20.270 108.460 22.670 ;
        RECT 109.000 22.160 109.330 22.330 ;
        RECT 108.860 20.950 109.030 21.990 ;
        RECT 109.300 20.950 109.470 21.990 ;
        RECT 109.000 20.610 109.330 20.780 ;
        RECT 109.870 20.270 110.040 22.670 ;
        RECT 108.290 20.240 110.040 20.270 ;
        RECT 110.315 22.675 112.065 22.845 ;
        RECT 110.315 20.240 110.485 22.675 ;
        RECT 111.025 22.165 111.355 22.335 ;
        RECT 103.220 19.605 107.220 19.775 ;
        RECT 107.850 19.275 110.485 20.240 ;
        RECT 110.885 19.955 111.055 21.995 ;
        RECT 111.325 19.955 111.495 21.995 ;
        RECT 111.025 19.615 111.355 19.785 ;
        RECT 111.895 19.275 112.065 22.675 ;
        RECT 107.850 19.265 112.065 19.275 ;
        RECT 86.130 19.245 112.065 19.265 ;
        RECT 114.130 22.665 136.020 22.835 ;
        RECT 114.130 19.265 114.300 22.665 ;
        RECT 114.930 22.155 118.930 22.325 ;
        RECT 114.700 19.945 114.870 21.985 ;
        RECT 118.990 19.945 119.160 21.985 ;
        RECT 114.930 19.605 118.930 19.775 ;
        RECT 119.560 19.265 119.730 22.665 ;
        RECT 120.360 22.155 124.360 22.325 ;
        RECT 120.130 19.945 120.300 21.985 ;
        RECT 124.420 19.945 124.590 21.985 ;
        RECT 120.360 19.605 124.360 19.775 ;
        RECT 124.990 19.265 125.160 22.665 ;
        RECT 125.790 22.155 129.790 22.325 ;
        RECT 125.560 19.945 125.730 21.985 ;
        RECT 129.850 19.945 130.020 21.985 ;
        RECT 125.790 19.605 129.790 19.775 ;
        RECT 130.420 19.265 130.590 22.665 ;
        RECT 131.220 22.155 135.220 22.325 ;
        RECT 130.990 19.945 131.160 21.985 ;
        RECT 135.280 19.945 135.450 21.985 ;
        RECT 135.850 20.240 136.020 22.665 ;
        RECT 136.290 22.670 138.040 22.840 ;
        RECT 136.290 20.270 136.460 22.670 ;
        RECT 137.000 22.160 137.330 22.330 ;
        RECT 136.860 20.950 137.030 21.990 ;
        RECT 137.300 20.950 137.470 21.990 ;
        RECT 137.000 20.610 137.330 20.780 ;
        RECT 137.870 20.270 138.040 22.670 ;
        RECT 136.290 20.240 138.040 20.270 ;
        RECT 138.315 22.675 140.065 22.845 ;
        RECT 138.315 20.240 138.485 22.675 ;
        RECT 139.025 22.165 139.355 22.335 ;
        RECT 131.220 19.605 135.220 19.775 ;
        RECT 135.850 19.275 138.485 20.240 ;
        RECT 138.885 19.955 139.055 21.995 ;
        RECT 139.325 19.955 139.495 21.995 ;
        RECT 139.025 19.615 139.355 19.785 ;
        RECT 139.895 19.275 140.065 22.675 ;
        RECT 135.850 19.265 140.065 19.275 ;
        RECT 114.130 19.245 140.065 19.265 ;
        RECT 1.475 19.105 28.065 19.245 ;
        RECT 29.475 19.105 56.065 19.245 ;
        RECT 57.475 19.105 84.065 19.245 ;
        RECT 85.475 19.105 112.065 19.245 ;
        RECT 113.475 19.105 140.065 19.245 ;
        RECT 1.475 18.380 28.055 19.105 ;
        RECT 29.475 18.380 56.055 19.105 ;
        RECT 57.475 18.380 84.055 19.105 ;
        RECT 85.475 18.380 112.055 19.105 ;
        RECT 113.475 18.380 140.055 19.105 ;
        RECT 1.450 17.480 27.925 17.960 ;
        RECT 29.450 17.480 55.925 17.960 ;
        RECT 57.450 17.480 83.925 17.960 ;
        RECT 85.450 17.480 111.925 17.960 ;
        RECT 113.450 17.480 139.925 17.960 ;
        RECT 1.435 17.420 27.925 17.480 ;
        RECT 29.435 17.420 55.925 17.480 ;
        RECT 57.435 17.420 83.925 17.480 ;
        RECT 85.435 17.420 111.925 17.480 ;
        RECT 113.435 17.420 139.925 17.480 ;
        RECT 1.435 17.260 27.980 17.420 ;
        RECT 1.435 17.235 14.180 17.260 ;
        RECT 1.435 17.005 5.760 17.235 ;
        RECT 1.470 7.745 1.640 17.005 ;
        RECT 2.365 16.435 4.405 16.605 ;
        RECT 1.980 8.375 2.150 16.375 ;
        RECT 4.620 8.375 4.790 16.375 ;
        RECT 2.365 8.145 4.405 8.315 ;
        RECT 5.130 7.745 5.300 17.005 ;
        RECT 1.470 7.575 5.300 7.745 ;
        RECT 5.590 7.745 5.760 17.005 ;
        RECT 6.390 16.725 8.390 16.895 ;
        RECT 6.160 8.470 6.330 16.510 ;
        RECT 8.450 8.470 8.620 16.510 ;
        RECT 6.390 8.085 8.390 8.255 ;
        RECT 9.020 7.745 9.190 17.235 ;
        RECT 9.820 16.725 11.820 16.895 ;
        RECT 9.590 8.470 9.760 16.510 ;
        RECT 11.880 8.470 12.050 16.510 ;
        RECT 12.450 15.665 14.180 17.235 ;
        RECT 26.230 17.250 27.980 17.260 ;
        RECT 12.450 15.495 20.915 15.665 ;
        RECT 12.450 14.085 14.255 15.495 ;
        RECT 14.595 14.625 14.765 14.955 ;
        RECT 14.980 14.925 20.020 15.095 ;
        RECT 14.980 14.485 20.020 14.655 ;
        RECT 20.235 14.625 20.405 14.955 ;
        RECT 20.745 14.085 20.915 15.495 ;
        RECT 12.450 13.915 20.915 14.085 ;
        RECT 12.450 13.400 14.180 13.915 ;
        RECT 12.450 13.285 23.930 13.400 ;
        RECT 9.820 8.085 11.820 8.255 ;
        RECT 12.450 7.745 12.620 13.285 ;
        RECT 5.590 7.575 12.620 7.745 ;
        RECT 12.900 13.230 23.930 13.285 ;
        RECT 12.900 7.740 13.070 13.230 ;
        RECT 13.700 12.720 17.700 12.890 ;
        RECT 13.470 8.465 13.640 12.505 ;
        RECT 17.760 8.465 17.930 12.505 ;
        RECT 13.700 8.080 17.700 8.250 ;
        RECT 18.330 7.740 18.500 13.230 ;
        RECT 19.130 12.720 23.130 12.890 ;
        RECT 18.900 8.465 19.070 12.505 ;
        RECT 23.190 8.465 23.360 12.505 ;
        RECT 19.130 8.080 23.130 8.250 ;
        RECT 23.760 7.740 23.930 13.230 ;
        RECT 12.900 7.570 23.930 7.740 ;
        RECT 24.205 13.245 25.955 13.415 ;
        RECT 24.205 7.755 24.375 13.245 ;
        RECT 24.915 12.735 25.245 12.905 ;
        RECT 24.775 8.480 24.945 12.520 ;
        RECT 25.215 8.480 25.385 12.520 ;
        RECT 24.915 8.095 25.245 8.265 ;
        RECT 25.785 7.755 25.955 13.245 ;
        RECT 24.205 7.585 25.955 7.755 ;
        RECT 26.230 7.760 26.400 17.250 ;
        RECT 26.940 16.740 27.270 16.910 ;
        RECT 26.800 8.485 26.970 16.525 ;
        RECT 27.240 8.485 27.410 16.525 ;
        RECT 26.940 8.100 27.270 8.270 ;
        RECT 27.810 7.760 27.980 17.250 ;
        RECT 29.435 17.260 55.980 17.420 ;
        RECT 29.435 17.235 42.180 17.260 ;
        RECT 29.435 17.005 33.760 17.235 ;
        RECT 26.230 7.590 27.980 7.760 ;
        RECT 29.470 7.745 29.640 17.005 ;
        RECT 30.365 16.435 32.405 16.605 ;
        RECT 29.980 8.375 30.150 16.375 ;
        RECT 32.620 8.375 32.790 16.375 ;
        RECT 30.365 8.145 32.405 8.315 ;
        RECT 33.130 7.745 33.300 17.005 ;
        RECT 29.470 7.575 33.300 7.745 ;
        RECT 33.590 7.745 33.760 17.005 ;
        RECT 34.390 16.725 36.390 16.895 ;
        RECT 34.160 8.470 34.330 16.510 ;
        RECT 36.450 8.470 36.620 16.510 ;
        RECT 34.390 8.085 36.390 8.255 ;
        RECT 37.020 7.745 37.190 17.235 ;
        RECT 37.820 16.725 39.820 16.895 ;
        RECT 37.590 8.470 37.760 16.510 ;
        RECT 39.880 8.470 40.050 16.510 ;
        RECT 40.450 15.665 42.180 17.235 ;
        RECT 54.230 17.250 55.980 17.260 ;
        RECT 40.450 15.495 48.915 15.665 ;
        RECT 40.450 14.085 42.255 15.495 ;
        RECT 42.595 14.625 42.765 14.955 ;
        RECT 42.980 14.925 48.020 15.095 ;
        RECT 42.980 14.485 48.020 14.655 ;
        RECT 48.235 14.625 48.405 14.955 ;
        RECT 48.745 14.085 48.915 15.495 ;
        RECT 40.450 13.915 48.915 14.085 ;
        RECT 40.450 13.400 42.180 13.915 ;
        RECT 40.450 13.285 51.930 13.400 ;
        RECT 37.820 8.085 39.820 8.255 ;
        RECT 40.450 7.745 40.620 13.285 ;
        RECT 33.590 7.575 40.620 7.745 ;
        RECT 40.900 13.230 51.930 13.285 ;
        RECT 40.900 7.740 41.070 13.230 ;
        RECT 41.700 12.720 45.700 12.890 ;
        RECT 41.470 8.465 41.640 12.505 ;
        RECT 45.760 8.465 45.930 12.505 ;
        RECT 41.700 8.080 45.700 8.250 ;
        RECT 46.330 7.740 46.500 13.230 ;
        RECT 47.130 12.720 51.130 12.890 ;
        RECT 46.900 8.465 47.070 12.505 ;
        RECT 51.190 8.465 51.360 12.505 ;
        RECT 47.130 8.080 51.130 8.250 ;
        RECT 51.760 7.740 51.930 13.230 ;
        RECT 40.900 7.570 51.930 7.740 ;
        RECT 52.205 13.245 53.955 13.415 ;
        RECT 52.205 7.755 52.375 13.245 ;
        RECT 52.915 12.735 53.245 12.905 ;
        RECT 52.775 8.480 52.945 12.520 ;
        RECT 53.215 8.480 53.385 12.520 ;
        RECT 52.915 8.095 53.245 8.265 ;
        RECT 53.785 7.755 53.955 13.245 ;
        RECT 52.205 7.585 53.955 7.755 ;
        RECT 54.230 7.760 54.400 17.250 ;
        RECT 54.940 16.740 55.270 16.910 ;
        RECT 54.800 8.485 54.970 16.525 ;
        RECT 55.240 8.485 55.410 16.525 ;
        RECT 54.940 8.100 55.270 8.270 ;
        RECT 55.810 7.760 55.980 17.250 ;
        RECT 57.435 17.260 83.980 17.420 ;
        RECT 57.435 17.235 70.180 17.260 ;
        RECT 57.435 17.005 61.760 17.235 ;
        RECT 54.230 7.590 55.980 7.760 ;
        RECT 57.470 7.745 57.640 17.005 ;
        RECT 58.365 16.435 60.405 16.605 ;
        RECT 57.980 8.375 58.150 16.375 ;
        RECT 60.620 8.375 60.790 16.375 ;
        RECT 58.365 8.145 60.405 8.315 ;
        RECT 61.130 7.745 61.300 17.005 ;
        RECT 57.470 7.575 61.300 7.745 ;
        RECT 61.590 7.745 61.760 17.005 ;
        RECT 62.390 16.725 64.390 16.895 ;
        RECT 62.160 8.470 62.330 16.510 ;
        RECT 64.450 8.470 64.620 16.510 ;
        RECT 62.390 8.085 64.390 8.255 ;
        RECT 65.020 7.745 65.190 17.235 ;
        RECT 65.820 16.725 67.820 16.895 ;
        RECT 65.590 8.470 65.760 16.510 ;
        RECT 67.880 8.470 68.050 16.510 ;
        RECT 68.450 15.665 70.180 17.235 ;
        RECT 82.230 17.250 83.980 17.260 ;
        RECT 68.450 15.495 76.915 15.665 ;
        RECT 68.450 14.085 70.255 15.495 ;
        RECT 70.595 14.625 70.765 14.955 ;
        RECT 70.980 14.925 76.020 15.095 ;
        RECT 70.980 14.485 76.020 14.655 ;
        RECT 76.235 14.625 76.405 14.955 ;
        RECT 76.745 14.085 76.915 15.495 ;
        RECT 68.450 13.915 76.915 14.085 ;
        RECT 68.450 13.400 70.180 13.915 ;
        RECT 68.450 13.285 79.930 13.400 ;
        RECT 65.820 8.085 67.820 8.255 ;
        RECT 68.450 7.745 68.620 13.285 ;
        RECT 61.590 7.575 68.620 7.745 ;
        RECT 68.900 13.230 79.930 13.285 ;
        RECT 68.900 7.740 69.070 13.230 ;
        RECT 69.700 12.720 73.700 12.890 ;
        RECT 69.470 8.465 69.640 12.505 ;
        RECT 73.760 8.465 73.930 12.505 ;
        RECT 69.700 8.080 73.700 8.250 ;
        RECT 74.330 7.740 74.500 13.230 ;
        RECT 75.130 12.720 79.130 12.890 ;
        RECT 74.900 8.465 75.070 12.505 ;
        RECT 79.190 8.465 79.360 12.505 ;
        RECT 75.130 8.080 79.130 8.250 ;
        RECT 79.760 7.740 79.930 13.230 ;
        RECT 68.900 7.570 79.930 7.740 ;
        RECT 80.205 13.245 81.955 13.415 ;
        RECT 80.205 7.755 80.375 13.245 ;
        RECT 80.915 12.735 81.245 12.905 ;
        RECT 80.775 8.480 80.945 12.520 ;
        RECT 81.215 8.480 81.385 12.520 ;
        RECT 80.915 8.095 81.245 8.265 ;
        RECT 81.785 7.755 81.955 13.245 ;
        RECT 80.205 7.585 81.955 7.755 ;
        RECT 82.230 7.760 82.400 17.250 ;
        RECT 82.940 16.740 83.270 16.910 ;
        RECT 82.800 8.485 82.970 16.525 ;
        RECT 83.240 8.485 83.410 16.525 ;
        RECT 82.940 8.100 83.270 8.270 ;
        RECT 83.810 7.760 83.980 17.250 ;
        RECT 85.435 17.260 111.980 17.420 ;
        RECT 85.435 17.235 98.180 17.260 ;
        RECT 85.435 17.005 89.760 17.235 ;
        RECT 82.230 7.590 83.980 7.760 ;
        RECT 85.470 7.745 85.640 17.005 ;
        RECT 86.365 16.435 88.405 16.605 ;
        RECT 85.980 8.375 86.150 16.375 ;
        RECT 88.620 8.375 88.790 16.375 ;
        RECT 86.365 8.145 88.405 8.315 ;
        RECT 89.130 7.745 89.300 17.005 ;
        RECT 85.470 7.575 89.300 7.745 ;
        RECT 89.590 7.745 89.760 17.005 ;
        RECT 90.390 16.725 92.390 16.895 ;
        RECT 90.160 8.470 90.330 16.510 ;
        RECT 92.450 8.470 92.620 16.510 ;
        RECT 90.390 8.085 92.390 8.255 ;
        RECT 93.020 7.745 93.190 17.235 ;
        RECT 93.820 16.725 95.820 16.895 ;
        RECT 93.590 8.470 93.760 16.510 ;
        RECT 95.880 8.470 96.050 16.510 ;
        RECT 96.450 15.665 98.180 17.235 ;
        RECT 110.230 17.250 111.980 17.260 ;
        RECT 96.450 15.495 104.915 15.665 ;
        RECT 96.450 14.085 98.255 15.495 ;
        RECT 98.595 14.625 98.765 14.955 ;
        RECT 98.980 14.925 104.020 15.095 ;
        RECT 98.980 14.485 104.020 14.655 ;
        RECT 104.235 14.625 104.405 14.955 ;
        RECT 104.745 14.085 104.915 15.495 ;
        RECT 96.450 13.915 104.915 14.085 ;
        RECT 96.450 13.400 98.180 13.915 ;
        RECT 96.450 13.285 107.930 13.400 ;
        RECT 93.820 8.085 95.820 8.255 ;
        RECT 96.450 7.745 96.620 13.285 ;
        RECT 89.590 7.575 96.620 7.745 ;
        RECT 96.900 13.230 107.930 13.285 ;
        RECT 96.900 7.740 97.070 13.230 ;
        RECT 97.700 12.720 101.700 12.890 ;
        RECT 97.470 8.465 97.640 12.505 ;
        RECT 101.760 8.465 101.930 12.505 ;
        RECT 97.700 8.080 101.700 8.250 ;
        RECT 102.330 7.740 102.500 13.230 ;
        RECT 103.130 12.720 107.130 12.890 ;
        RECT 102.900 8.465 103.070 12.505 ;
        RECT 107.190 8.465 107.360 12.505 ;
        RECT 103.130 8.080 107.130 8.250 ;
        RECT 107.760 7.740 107.930 13.230 ;
        RECT 96.900 7.570 107.930 7.740 ;
        RECT 108.205 13.245 109.955 13.415 ;
        RECT 108.205 7.755 108.375 13.245 ;
        RECT 108.915 12.735 109.245 12.905 ;
        RECT 108.775 8.480 108.945 12.520 ;
        RECT 109.215 8.480 109.385 12.520 ;
        RECT 108.915 8.095 109.245 8.265 ;
        RECT 109.785 7.755 109.955 13.245 ;
        RECT 108.205 7.585 109.955 7.755 ;
        RECT 110.230 7.760 110.400 17.250 ;
        RECT 110.940 16.740 111.270 16.910 ;
        RECT 110.800 8.485 110.970 16.525 ;
        RECT 111.240 8.485 111.410 16.525 ;
        RECT 110.940 8.100 111.270 8.270 ;
        RECT 111.810 7.760 111.980 17.250 ;
        RECT 113.435 17.260 139.980 17.420 ;
        RECT 113.435 17.235 126.180 17.260 ;
        RECT 113.435 17.005 117.760 17.235 ;
        RECT 110.230 7.590 111.980 7.760 ;
        RECT 113.470 7.745 113.640 17.005 ;
        RECT 114.365 16.435 116.405 16.605 ;
        RECT 113.980 8.375 114.150 16.375 ;
        RECT 116.620 8.375 116.790 16.375 ;
        RECT 114.365 8.145 116.405 8.315 ;
        RECT 117.130 7.745 117.300 17.005 ;
        RECT 113.470 7.575 117.300 7.745 ;
        RECT 117.590 7.745 117.760 17.005 ;
        RECT 118.390 16.725 120.390 16.895 ;
        RECT 118.160 8.470 118.330 16.510 ;
        RECT 120.450 8.470 120.620 16.510 ;
        RECT 118.390 8.085 120.390 8.255 ;
        RECT 121.020 7.745 121.190 17.235 ;
        RECT 121.820 16.725 123.820 16.895 ;
        RECT 121.590 8.470 121.760 16.510 ;
        RECT 123.880 8.470 124.050 16.510 ;
        RECT 124.450 15.665 126.180 17.235 ;
        RECT 138.230 17.250 139.980 17.260 ;
        RECT 124.450 15.495 132.915 15.665 ;
        RECT 124.450 14.085 126.255 15.495 ;
        RECT 126.595 14.625 126.765 14.955 ;
        RECT 126.980 14.925 132.020 15.095 ;
        RECT 126.980 14.485 132.020 14.655 ;
        RECT 132.235 14.625 132.405 14.955 ;
        RECT 132.745 14.085 132.915 15.495 ;
        RECT 124.450 13.915 132.915 14.085 ;
        RECT 124.450 13.400 126.180 13.915 ;
        RECT 124.450 13.285 135.930 13.400 ;
        RECT 121.820 8.085 123.820 8.255 ;
        RECT 124.450 7.745 124.620 13.285 ;
        RECT 117.590 7.575 124.620 7.745 ;
        RECT 124.900 13.230 135.930 13.285 ;
        RECT 124.900 7.740 125.070 13.230 ;
        RECT 125.700 12.720 129.700 12.890 ;
        RECT 125.470 8.465 125.640 12.505 ;
        RECT 129.760 8.465 129.930 12.505 ;
        RECT 125.700 8.080 129.700 8.250 ;
        RECT 130.330 7.740 130.500 13.230 ;
        RECT 131.130 12.720 135.130 12.890 ;
        RECT 130.900 8.465 131.070 12.505 ;
        RECT 135.190 8.465 135.360 12.505 ;
        RECT 131.130 8.080 135.130 8.250 ;
        RECT 135.760 7.740 135.930 13.230 ;
        RECT 124.900 7.570 135.930 7.740 ;
        RECT 136.205 13.245 137.955 13.415 ;
        RECT 136.205 7.755 136.375 13.245 ;
        RECT 136.915 12.735 137.245 12.905 ;
        RECT 136.775 8.480 136.945 12.520 ;
        RECT 137.215 8.480 137.385 12.520 ;
        RECT 136.915 8.095 137.245 8.265 ;
        RECT 137.785 7.755 137.955 13.245 ;
        RECT 136.205 7.585 137.955 7.755 ;
        RECT 138.230 7.760 138.400 17.250 ;
        RECT 138.940 16.740 139.270 16.910 ;
        RECT 138.800 8.485 138.970 16.525 ;
        RECT 139.240 8.485 139.410 16.525 ;
        RECT 138.940 8.100 139.270 8.270 ;
        RECT 139.810 7.760 139.980 17.250 ;
        RECT 138.230 7.590 139.980 7.760 ;
        RECT 2.130 6.665 24.020 6.835 ;
        RECT 2.130 3.265 2.300 6.665 ;
        RECT 2.930 6.155 6.930 6.325 ;
        RECT 2.700 3.945 2.870 5.985 ;
        RECT 6.990 3.945 7.160 5.985 ;
        RECT 2.930 3.605 6.930 3.775 ;
        RECT 7.560 3.265 7.730 6.665 ;
        RECT 8.360 6.155 12.360 6.325 ;
        RECT 8.130 3.945 8.300 5.985 ;
        RECT 12.420 3.945 12.590 5.985 ;
        RECT 8.360 3.605 12.360 3.775 ;
        RECT 12.990 3.265 13.160 6.665 ;
        RECT 13.790 6.155 17.790 6.325 ;
        RECT 13.560 3.945 13.730 5.985 ;
        RECT 17.850 3.945 18.020 5.985 ;
        RECT 13.790 3.605 17.790 3.775 ;
        RECT 18.420 3.265 18.590 6.665 ;
        RECT 19.220 6.155 23.220 6.325 ;
        RECT 18.990 3.945 19.160 5.985 ;
        RECT 23.280 3.945 23.450 5.985 ;
        RECT 23.850 4.240 24.020 6.665 ;
        RECT 24.290 6.670 26.040 6.840 ;
        RECT 24.290 4.270 24.460 6.670 ;
        RECT 25.000 6.160 25.330 6.330 ;
        RECT 24.860 4.950 25.030 5.990 ;
        RECT 25.300 4.950 25.470 5.990 ;
        RECT 25.000 4.610 25.330 4.780 ;
        RECT 25.870 4.270 26.040 6.670 ;
        RECT 24.290 4.240 26.040 4.270 ;
        RECT 26.315 6.675 28.065 6.845 ;
        RECT 26.315 4.240 26.485 6.675 ;
        RECT 27.025 6.165 27.355 6.335 ;
        RECT 19.220 3.605 23.220 3.775 ;
        RECT 23.850 3.275 26.485 4.240 ;
        RECT 26.885 3.955 27.055 5.995 ;
        RECT 27.325 3.955 27.495 5.995 ;
        RECT 27.025 3.615 27.355 3.785 ;
        RECT 27.895 3.275 28.065 6.675 ;
        RECT 23.850 3.265 28.065 3.275 ;
        RECT 2.130 3.245 28.065 3.265 ;
        RECT 30.130 6.665 52.020 6.835 ;
        RECT 30.130 3.265 30.300 6.665 ;
        RECT 30.930 6.155 34.930 6.325 ;
        RECT 30.700 3.945 30.870 5.985 ;
        RECT 34.990 3.945 35.160 5.985 ;
        RECT 30.930 3.605 34.930 3.775 ;
        RECT 35.560 3.265 35.730 6.665 ;
        RECT 36.360 6.155 40.360 6.325 ;
        RECT 36.130 3.945 36.300 5.985 ;
        RECT 40.420 3.945 40.590 5.985 ;
        RECT 36.360 3.605 40.360 3.775 ;
        RECT 40.990 3.265 41.160 6.665 ;
        RECT 41.790 6.155 45.790 6.325 ;
        RECT 41.560 3.945 41.730 5.985 ;
        RECT 45.850 3.945 46.020 5.985 ;
        RECT 41.790 3.605 45.790 3.775 ;
        RECT 46.420 3.265 46.590 6.665 ;
        RECT 47.220 6.155 51.220 6.325 ;
        RECT 46.990 3.945 47.160 5.985 ;
        RECT 51.280 3.945 51.450 5.985 ;
        RECT 51.850 4.240 52.020 6.665 ;
        RECT 52.290 6.670 54.040 6.840 ;
        RECT 52.290 4.270 52.460 6.670 ;
        RECT 53.000 6.160 53.330 6.330 ;
        RECT 52.860 4.950 53.030 5.990 ;
        RECT 53.300 4.950 53.470 5.990 ;
        RECT 53.000 4.610 53.330 4.780 ;
        RECT 53.870 4.270 54.040 6.670 ;
        RECT 52.290 4.240 54.040 4.270 ;
        RECT 54.315 6.675 56.065 6.845 ;
        RECT 54.315 4.240 54.485 6.675 ;
        RECT 55.025 6.165 55.355 6.335 ;
        RECT 47.220 3.605 51.220 3.775 ;
        RECT 51.850 3.275 54.485 4.240 ;
        RECT 54.885 3.955 55.055 5.995 ;
        RECT 55.325 3.955 55.495 5.995 ;
        RECT 55.025 3.615 55.355 3.785 ;
        RECT 55.895 3.275 56.065 6.675 ;
        RECT 51.850 3.265 56.065 3.275 ;
        RECT 30.130 3.245 56.065 3.265 ;
        RECT 58.130 6.665 80.020 6.835 ;
        RECT 58.130 3.265 58.300 6.665 ;
        RECT 58.930 6.155 62.930 6.325 ;
        RECT 58.700 3.945 58.870 5.985 ;
        RECT 62.990 3.945 63.160 5.985 ;
        RECT 58.930 3.605 62.930 3.775 ;
        RECT 63.560 3.265 63.730 6.665 ;
        RECT 64.360 6.155 68.360 6.325 ;
        RECT 64.130 3.945 64.300 5.985 ;
        RECT 68.420 3.945 68.590 5.985 ;
        RECT 64.360 3.605 68.360 3.775 ;
        RECT 68.990 3.265 69.160 6.665 ;
        RECT 69.790 6.155 73.790 6.325 ;
        RECT 69.560 3.945 69.730 5.985 ;
        RECT 73.850 3.945 74.020 5.985 ;
        RECT 69.790 3.605 73.790 3.775 ;
        RECT 74.420 3.265 74.590 6.665 ;
        RECT 75.220 6.155 79.220 6.325 ;
        RECT 74.990 3.945 75.160 5.985 ;
        RECT 79.280 3.945 79.450 5.985 ;
        RECT 79.850 4.240 80.020 6.665 ;
        RECT 80.290 6.670 82.040 6.840 ;
        RECT 80.290 4.270 80.460 6.670 ;
        RECT 81.000 6.160 81.330 6.330 ;
        RECT 80.860 4.950 81.030 5.990 ;
        RECT 81.300 4.950 81.470 5.990 ;
        RECT 81.000 4.610 81.330 4.780 ;
        RECT 81.870 4.270 82.040 6.670 ;
        RECT 80.290 4.240 82.040 4.270 ;
        RECT 82.315 6.675 84.065 6.845 ;
        RECT 82.315 4.240 82.485 6.675 ;
        RECT 83.025 6.165 83.355 6.335 ;
        RECT 75.220 3.605 79.220 3.775 ;
        RECT 79.850 3.275 82.485 4.240 ;
        RECT 82.885 3.955 83.055 5.995 ;
        RECT 83.325 3.955 83.495 5.995 ;
        RECT 83.025 3.615 83.355 3.785 ;
        RECT 83.895 3.275 84.065 6.675 ;
        RECT 79.850 3.265 84.065 3.275 ;
        RECT 58.130 3.245 84.065 3.265 ;
        RECT 86.130 6.665 108.020 6.835 ;
        RECT 86.130 3.265 86.300 6.665 ;
        RECT 86.930 6.155 90.930 6.325 ;
        RECT 86.700 3.945 86.870 5.985 ;
        RECT 90.990 3.945 91.160 5.985 ;
        RECT 86.930 3.605 90.930 3.775 ;
        RECT 91.560 3.265 91.730 6.665 ;
        RECT 92.360 6.155 96.360 6.325 ;
        RECT 92.130 3.945 92.300 5.985 ;
        RECT 96.420 3.945 96.590 5.985 ;
        RECT 92.360 3.605 96.360 3.775 ;
        RECT 96.990 3.265 97.160 6.665 ;
        RECT 97.790 6.155 101.790 6.325 ;
        RECT 97.560 3.945 97.730 5.985 ;
        RECT 101.850 3.945 102.020 5.985 ;
        RECT 97.790 3.605 101.790 3.775 ;
        RECT 102.420 3.265 102.590 6.665 ;
        RECT 103.220 6.155 107.220 6.325 ;
        RECT 102.990 3.945 103.160 5.985 ;
        RECT 107.280 3.945 107.450 5.985 ;
        RECT 107.850 4.240 108.020 6.665 ;
        RECT 108.290 6.670 110.040 6.840 ;
        RECT 108.290 4.270 108.460 6.670 ;
        RECT 109.000 6.160 109.330 6.330 ;
        RECT 108.860 4.950 109.030 5.990 ;
        RECT 109.300 4.950 109.470 5.990 ;
        RECT 109.000 4.610 109.330 4.780 ;
        RECT 109.870 4.270 110.040 6.670 ;
        RECT 108.290 4.240 110.040 4.270 ;
        RECT 110.315 6.675 112.065 6.845 ;
        RECT 110.315 4.240 110.485 6.675 ;
        RECT 111.025 6.165 111.355 6.335 ;
        RECT 103.220 3.605 107.220 3.775 ;
        RECT 107.850 3.275 110.485 4.240 ;
        RECT 110.885 3.955 111.055 5.995 ;
        RECT 111.325 3.955 111.495 5.995 ;
        RECT 111.025 3.615 111.355 3.785 ;
        RECT 111.895 3.275 112.065 6.675 ;
        RECT 107.850 3.265 112.065 3.275 ;
        RECT 86.130 3.245 112.065 3.265 ;
        RECT 114.130 6.665 136.020 6.835 ;
        RECT 114.130 3.265 114.300 6.665 ;
        RECT 114.930 6.155 118.930 6.325 ;
        RECT 114.700 3.945 114.870 5.985 ;
        RECT 118.990 3.945 119.160 5.985 ;
        RECT 114.930 3.605 118.930 3.775 ;
        RECT 119.560 3.265 119.730 6.665 ;
        RECT 120.360 6.155 124.360 6.325 ;
        RECT 120.130 3.945 120.300 5.985 ;
        RECT 124.420 3.945 124.590 5.985 ;
        RECT 120.360 3.605 124.360 3.775 ;
        RECT 124.990 3.265 125.160 6.665 ;
        RECT 125.790 6.155 129.790 6.325 ;
        RECT 125.560 3.945 125.730 5.985 ;
        RECT 129.850 3.945 130.020 5.985 ;
        RECT 125.790 3.605 129.790 3.775 ;
        RECT 130.420 3.265 130.590 6.665 ;
        RECT 131.220 6.155 135.220 6.325 ;
        RECT 130.990 3.945 131.160 5.985 ;
        RECT 135.280 3.945 135.450 5.985 ;
        RECT 135.850 4.240 136.020 6.665 ;
        RECT 136.290 6.670 138.040 6.840 ;
        RECT 136.290 4.270 136.460 6.670 ;
        RECT 137.000 6.160 137.330 6.330 ;
        RECT 136.860 4.950 137.030 5.990 ;
        RECT 137.300 4.950 137.470 5.990 ;
        RECT 137.000 4.610 137.330 4.780 ;
        RECT 137.870 4.270 138.040 6.670 ;
        RECT 136.290 4.240 138.040 4.270 ;
        RECT 138.315 6.675 140.065 6.845 ;
        RECT 138.315 4.240 138.485 6.675 ;
        RECT 139.025 6.165 139.355 6.335 ;
        RECT 131.220 3.605 135.220 3.775 ;
        RECT 135.850 3.275 138.485 4.240 ;
        RECT 138.885 3.955 139.055 5.995 ;
        RECT 139.325 3.955 139.495 5.995 ;
        RECT 139.025 3.615 139.355 3.785 ;
        RECT 139.895 3.275 140.065 6.675 ;
        RECT 135.850 3.265 140.065 3.275 ;
        RECT 114.130 3.245 140.065 3.265 ;
        RECT 1.475 3.105 28.065 3.245 ;
        RECT 29.475 3.105 56.065 3.245 ;
        RECT 57.475 3.105 84.065 3.245 ;
        RECT 85.475 3.105 112.065 3.245 ;
        RECT 113.475 3.105 140.065 3.245 ;
        RECT 1.475 2.380 28.055 3.105 ;
        RECT 29.475 2.380 56.055 3.105 ;
        RECT 57.475 2.380 84.055 3.105 ;
        RECT 85.475 2.380 112.055 3.105 ;
        RECT 113.475 2.380 140.055 3.105 ;
      LAYER met1 ;
        RECT 99.010 207.030 99.330 207.090 ;
        RECT 133.510 207.030 133.830 207.090 ;
        RECT 99.010 206.890 133.830 207.030 ;
        RECT 99.010 206.830 99.330 206.890 ;
        RECT 133.510 206.830 133.830 206.890 ;
        RECT 102.690 195.810 103.010 195.870 ;
        RECT 121.090 195.810 121.410 195.870 ;
        RECT 102.690 195.670 121.410 195.810 ;
        RECT 102.690 195.610 103.010 195.670 ;
        RECT 121.090 195.610 121.410 195.670 ;
        RECT 88.890 195.470 89.210 195.530 ;
        RECT 93.030 195.470 93.350 195.530 ;
        RECT 88.890 195.330 93.350 195.470 ;
        RECT 88.890 195.270 89.210 195.330 ;
        RECT 93.030 195.270 93.350 195.330 ;
        RECT 99.930 195.470 100.250 195.530 ;
        RECT 125.230 195.470 125.550 195.530 ;
        RECT 99.930 195.330 125.550 195.470 ;
        RECT 99.930 195.270 100.250 195.330 ;
        RECT 125.230 195.270 125.550 195.330 ;
        RECT 125.690 195.470 126.010 195.530 ;
        RECT 131.210 195.470 131.530 195.530 ;
        RECT 125.690 195.330 131.530 195.470 ;
        RECT 125.690 195.270 126.010 195.330 ;
        RECT 131.210 195.270 131.530 195.330 ;
        RECT 23.500 194.650 136.200 195.130 ;
        RECT 66.350 194.450 66.670 194.510 ;
        RECT 67.285 194.450 67.575 194.495 ;
        RECT 66.350 194.310 67.575 194.450 ;
        RECT 66.350 194.250 66.670 194.310 ;
        RECT 67.285 194.265 67.575 194.310 ;
        RECT 76.010 194.450 76.330 194.510 ;
        RECT 76.485 194.450 76.775 194.495 ;
        RECT 76.010 194.310 76.775 194.450 ;
        RECT 76.010 194.250 76.330 194.310 ;
        RECT 76.485 194.265 76.775 194.310 ;
        RECT 85.670 194.450 85.990 194.510 ;
        RECT 89.365 194.450 89.655 194.495 ;
        RECT 85.670 194.310 89.655 194.450 ;
        RECT 85.670 194.250 85.990 194.310 ;
        RECT 89.365 194.265 89.655 194.310 ;
        RECT 92.110 194.450 92.430 194.510 ;
        RECT 93.505 194.450 93.795 194.495 ;
        RECT 92.110 194.310 93.795 194.450 ;
        RECT 92.110 194.250 92.430 194.310 ;
        RECT 93.505 194.265 93.795 194.310 ;
        RECT 95.330 194.450 95.650 194.510 ;
        RECT 95.805 194.450 96.095 194.495 ;
        RECT 95.330 194.310 96.095 194.450 ;
        RECT 95.330 194.250 95.650 194.310 ;
        RECT 95.805 194.265 96.095 194.310 ;
        RECT 98.550 194.250 98.870 194.510 ;
        RECT 101.770 194.450 102.090 194.510 ;
        RECT 102.705 194.450 102.995 194.495 ;
        RECT 101.770 194.310 102.995 194.450 ;
        RECT 101.770 194.250 102.090 194.310 ;
        RECT 102.705 194.265 102.995 194.310 ;
        RECT 104.990 194.450 105.310 194.510 ;
        RECT 105.925 194.450 106.215 194.495 ;
        RECT 104.990 194.310 106.215 194.450 ;
        RECT 104.990 194.250 105.310 194.310 ;
        RECT 105.925 194.265 106.215 194.310 ;
        RECT 114.650 194.450 114.970 194.510 ;
        RECT 115.585 194.450 115.875 194.495 ;
        RECT 122.485 194.450 122.775 194.495 ;
        RECT 114.650 194.310 115.875 194.450 ;
        RECT 114.650 194.250 114.970 194.310 ;
        RECT 115.585 194.265 115.875 194.310 ;
        RECT 120.720 194.310 122.775 194.450 ;
        RECT 93.950 194.110 94.270 194.170 ;
        RECT 107.290 194.110 107.610 194.170 ;
        RECT 77.480 193.970 94.270 194.110 ;
        RECT 26.345 193.770 26.635 193.815 ;
        RECT 27.710 193.770 28.030 193.830 ;
        RECT 26.345 193.630 28.030 193.770 ;
        RECT 26.345 193.585 26.635 193.630 ;
        RECT 27.710 193.570 28.030 193.630 ;
        RECT 34.610 193.770 34.930 193.830 ;
        RECT 37.385 193.770 37.675 193.815 ;
        RECT 34.610 193.630 37.675 193.770 ;
        RECT 34.610 193.570 34.930 193.630 ;
        RECT 37.385 193.585 37.675 193.630 ;
        RECT 38.765 193.585 39.055 193.815 ;
        RECT 39.225 193.770 39.515 193.815 ;
        RECT 41.510 193.770 41.830 193.830 ;
        RECT 39.225 193.630 41.830 193.770 ;
        RECT 39.225 193.585 39.515 193.630 ;
        RECT 24.490 193.430 24.810 193.490 ;
        RECT 26.805 193.430 27.095 193.475 ;
        RECT 24.490 193.290 27.095 193.430 ;
        RECT 38.840 193.430 38.980 193.585 ;
        RECT 41.510 193.570 41.830 193.630 ;
        RECT 63.130 193.770 63.450 193.830 ;
        RECT 63.605 193.770 63.895 193.815 ;
        RECT 63.130 193.630 63.895 193.770 ;
        RECT 63.130 193.570 63.450 193.630 ;
        RECT 63.605 193.585 63.895 193.630 ;
        RECT 67.730 193.770 68.050 193.830 ;
        RECT 68.205 193.770 68.495 193.815 ;
        RECT 67.730 193.630 68.495 193.770 ;
        RECT 67.730 193.570 68.050 193.630 ;
        RECT 68.205 193.585 68.495 193.630 ;
        RECT 72.790 193.770 73.110 193.830 ;
        RECT 77.480 193.815 77.620 193.970 ;
        RECT 93.950 193.910 94.270 193.970 ;
        RECT 97.720 193.970 107.610 194.110 ;
        RECT 73.265 193.770 73.555 193.815 ;
        RECT 72.790 193.630 73.555 193.770 ;
        RECT 72.790 193.570 73.110 193.630 ;
        RECT 73.265 193.585 73.555 193.630 ;
        RECT 77.405 193.585 77.695 193.815 ;
        RECT 79.230 193.570 79.550 193.830 ;
        RECT 81.530 193.570 81.850 193.830 ;
        RECT 82.450 193.770 82.770 193.830 ;
        RECT 82.925 193.770 83.215 193.815 ;
        RECT 82.450 193.630 83.215 193.770 ;
        RECT 82.450 193.570 82.770 193.630 ;
        RECT 82.925 193.585 83.215 193.630 ;
        RECT 87.510 193.770 87.830 193.830 ;
        RECT 88.445 193.770 88.735 193.815 ;
        RECT 87.510 193.630 88.735 193.770 ;
        RECT 87.510 193.570 87.830 193.630 ;
        RECT 88.445 193.585 88.735 193.630 ;
        RECT 91.190 193.570 91.510 193.830 ;
        RECT 92.585 193.770 92.875 193.815 ;
        RECT 92.200 193.630 92.875 193.770 ;
        RECT 41.970 193.430 42.290 193.490 ;
        RECT 38.840 193.290 42.290 193.430 ;
        RECT 24.490 193.230 24.810 193.290 ;
        RECT 26.805 193.245 27.095 193.290 ;
        RECT 41.970 193.230 42.290 193.290 ;
        RECT 83.370 193.430 83.690 193.490 ;
        RECT 84.305 193.430 84.595 193.475 ;
        RECT 83.370 193.290 84.595 193.430 ;
        RECT 83.370 193.230 83.690 193.290 ;
        RECT 84.305 193.245 84.595 193.290 ;
        RECT 45.190 193.090 45.510 193.150 ;
        RECT 78.310 193.090 78.630 193.150 ;
        RECT 92.200 193.135 92.340 193.630 ;
        RECT 92.585 193.585 92.875 193.630 ;
        RECT 93.030 193.770 93.350 193.830 ;
        RECT 97.720 193.815 97.860 193.970 ;
        RECT 107.290 193.910 107.610 193.970 ;
        RECT 110.065 194.110 110.355 194.155 ;
        RECT 120.720 194.110 120.860 194.310 ;
        RECT 122.485 194.265 122.775 194.310 ;
        RECT 110.065 193.970 112.120 194.110 ;
        RECT 110.065 193.925 110.355 193.970 ;
        RECT 111.980 193.830 112.120 193.970 ;
        RECT 117.040 193.970 120.860 194.110 ;
        RECT 94.425 193.770 94.715 193.815 ;
        RECT 93.030 193.630 94.715 193.770 ;
        RECT 93.030 193.570 93.350 193.630 ;
        RECT 94.425 193.585 94.715 193.630 ;
        RECT 96.725 193.585 97.015 193.815 ;
        RECT 97.645 193.585 97.935 193.815 ;
        RECT 96.800 193.430 96.940 193.585 ;
        RECT 100.390 193.570 100.710 193.830 ;
        RECT 103.610 193.570 103.930 193.830 ;
        RECT 105.005 193.770 105.295 193.815 ;
        RECT 106.370 193.770 106.690 193.830 ;
        RECT 105.005 193.630 106.690 193.770 ;
        RECT 105.005 193.585 105.295 193.630 ;
        RECT 106.370 193.570 106.690 193.630 ;
        RECT 106.830 193.570 107.150 193.830 ;
        RECT 108.225 193.770 108.515 193.815 ;
        RECT 110.985 193.770 111.275 193.815 ;
        RECT 108.225 193.630 111.275 193.770 ;
        RECT 108.225 193.585 108.515 193.630 ;
        RECT 110.985 193.585 111.275 193.630 ;
        RECT 110.510 193.430 110.830 193.490 ;
        RECT 96.800 193.290 110.830 193.430 ;
        RECT 110.510 193.230 110.830 193.290 ;
        RECT 111.060 193.150 111.200 193.585 ;
        RECT 111.890 193.570 112.210 193.830 ;
        RECT 112.365 193.585 112.655 193.815 ;
        RECT 112.440 193.430 112.580 193.585 ;
        RECT 116.490 193.570 116.810 193.830 ;
        RECT 117.040 193.475 117.180 193.970 ;
        RECT 120.720 193.815 120.860 193.970 ;
        RECT 130.290 194.110 130.610 194.170 ;
        RECT 131.670 194.110 131.990 194.170 ;
        RECT 132.605 194.110 132.895 194.155 ;
        RECT 130.290 193.970 132.895 194.110 ;
        RECT 130.290 193.910 130.610 193.970 ;
        RECT 117.885 193.585 118.175 193.815 ;
        RECT 120.645 193.585 120.935 193.815 ;
        RECT 116.965 193.430 117.255 193.475 ;
        RECT 112.440 193.290 117.255 193.430 ;
        RECT 116.965 193.245 117.255 193.290 ;
        RECT 45.190 192.950 78.630 193.090 ;
        RECT 45.190 192.890 45.510 192.950 ;
        RECT 78.310 192.890 78.630 192.950 ;
        RECT 92.125 192.905 92.415 193.135 ;
        RECT 98.090 193.090 98.410 193.150 ;
        RECT 99.485 193.090 99.775 193.135 ;
        RECT 94.960 192.950 97.860 193.090 ;
        RECT 19.890 192.750 20.210 192.810 ;
        RECT 25.425 192.750 25.715 192.795 ;
        RECT 19.890 192.610 25.715 192.750 ;
        RECT 19.890 192.550 20.210 192.610 ;
        RECT 25.425 192.565 25.715 192.610 ;
        RECT 37.845 192.750 38.135 192.795 ;
        RECT 38.290 192.750 38.610 192.810 ;
        RECT 37.845 192.610 38.610 192.750 ;
        RECT 37.845 192.565 38.135 192.610 ;
        RECT 38.290 192.550 38.610 192.610 ;
        RECT 40.145 192.750 40.435 192.795 ;
        RECT 47.030 192.750 47.350 192.810 ;
        RECT 40.145 192.610 47.350 192.750 ;
        RECT 40.145 192.565 40.435 192.610 ;
        RECT 47.030 192.550 47.350 192.610 ;
        RECT 64.510 192.550 64.830 192.810 ;
        RECT 74.185 192.750 74.475 192.795 ;
        RECT 76.010 192.750 76.330 192.810 ;
        RECT 74.185 192.610 76.330 192.750 ;
        RECT 74.185 192.565 74.475 192.610 ;
        RECT 76.010 192.550 76.330 192.610 ;
        RECT 80.150 192.550 80.470 192.810 ;
        RECT 81.085 192.750 81.375 192.795 ;
        RECT 81.530 192.750 81.850 192.810 ;
        RECT 81.085 192.610 81.850 192.750 ;
        RECT 81.085 192.565 81.375 192.610 ;
        RECT 81.530 192.550 81.850 192.610 ;
        RECT 82.465 192.750 82.755 192.795 ;
        RECT 94.960 192.750 95.100 192.950 ;
        RECT 82.465 192.610 95.100 192.750 ;
        RECT 82.465 192.565 82.755 192.610 ;
        RECT 95.330 192.550 95.650 192.810 ;
        RECT 97.720 192.750 97.860 192.950 ;
        RECT 98.090 192.950 99.775 193.090 ;
        RECT 98.090 192.890 98.410 192.950 ;
        RECT 99.485 192.905 99.775 192.950 ;
        RECT 100.850 193.090 101.170 193.150 ;
        RECT 103.610 193.090 103.930 193.150 ;
        RECT 107.305 193.090 107.595 193.135 ;
        RECT 110.970 193.090 111.290 193.150 ;
        RECT 115.570 193.090 115.890 193.150 ;
        RECT 117.960 193.090 118.100 193.585 ;
        RECT 122.010 193.570 122.330 193.830 ;
        RECT 123.390 193.570 123.710 193.830 ;
        RECT 125.230 193.570 125.550 193.830 ;
        RECT 127.070 193.570 127.390 193.830 ;
        RECT 129.830 193.570 130.150 193.830 ;
        RECT 130.840 193.815 130.980 193.970 ;
        RECT 131.670 193.910 131.990 193.970 ;
        RECT 132.605 193.925 132.895 193.970 ;
        RECT 133.510 194.110 133.830 194.170 ;
        RECT 134.445 194.110 134.735 194.155 ;
        RECT 133.510 193.970 134.735 194.110 ;
        RECT 133.510 193.910 133.830 193.970 ;
        RECT 134.445 193.925 134.735 193.970 ;
        RECT 130.765 193.585 131.055 193.815 ;
        RECT 131.225 193.585 131.515 193.815 ;
        RECT 123.850 193.230 124.170 193.490 ;
        RECT 126.165 193.430 126.455 193.475 ;
        RECT 130.305 193.430 130.595 193.475 ;
        RECT 131.300 193.430 131.440 193.585 ;
        RECT 133.525 193.430 133.815 193.475 ;
        RECT 126.165 193.290 130.595 193.430 ;
        RECT 126.165 193.245 126.455 193.290 ;
        RECT 130.305 193.245 130.595 193.290 ;
        RECT 130.840 193.290 133.815 193.430 ;
        RECT 100.850 192.950 102.000 193.090 ;
        RECT 100.850 192.890 101.170 192.950 ;
        RECT 101.310 192.750 101.630 192.810 ;
        RECT 97.720 192.610 101.630 192.750 ;
        RECT 101.860 192.750 102.000 192.950 ;
        RECT 103.610 192.950 107.595 193.090 ;
        RECT 103.610 192.890 103.930 192.950 ;
        RECT 107.305 192.905 107.595 192.950 ;
        RECT 108.760 192.950 110.740 193.090 ;
        RECT 104.085 192.750 104.375 192.795 ;
        RECT 108.760 192.750 108.900 192.950 ;
        RECT 101.860 192.610 108.900 192.750 ;
        RECT 101.310 192.550 101.630 192.610 ;
        RECT 104.085 192.565 104.375 192.610 ;
        RECT 109.130 192.550 109.450 192.810 ;
        RECT 110.600 192.750 110.740 192.950 ;
        RECT 110.970 192.950 114.880 193.090 ;
        RECT 110.970 192.890 111.290 192.950 ;
        RECT 112.350 192.750 112.670 192.810 ;
        RECT 110.600 192.610 112.670 192.750 ;
        RECT 112.350 192.550 112.670 192.610 ;
        RECT 113.285 192.750 113.575 192.795 ;
        RECT 114.190 192.750 114.510 192.810 ;
        RECT 113.285 192.610 114.510 192.750 ;
        RECT 114.740 192.750 114.880 192.950 ;
        RECT 115.570 192.950 118.100 193.090 ;
        RECT 118.805 193.090 119.095 193.135 ;
        RECT 129.830 193.090 130.150 193.150 ;
        RECT 118.805 192.950 130.150 193.090 ;
        RECT 115.570 192.890 115.890 192.950 ;
        RECT 118.805 192.905 119.095 192.950 ;
        RECT 129.830 192.890 130.150 192.950 ;
        RECT 120.185 192.750 120.475 192.795 ;
        RECT 114.740 192.610 120.475 192.750 ;
        RECT 113.285 192.565 113.575 192.610 ;
        RECT 114.190 192.550 114.510 192.610 ;
        RECT 120.185 192.565 120.475 192.610 ;
        RECT 121.090 192.550 121.410 192.810 ;
        RECT 124.310 192.550 124.630 192.810 ;
        RECT 125.230 192.750 125.550 192.810 ;
        RECT 128.005 192.750 128.295 192.795 ;
        RECT 125.230 192.610 128.295 192.750 ;
        RECT 125.230 192.550 125.550 192.610 ;
        RECT 128.005 192.565 128.295 192.610 ;
        RECT 128.450 192.750 128.770 192.810 ;
        RECT 130.840 192.750 130.980 193.290 ;
        RECT 133.525 193.245 133.815 193.290 ;
        RECT 131.210 193.090 131.530 193.150 ;
        RECT 133.985 193.090 134.275 193.135 ;
        RECT 131.210 192.950 134.275 193.090 ;
        RECT 131.210 192.890 131.530 192.950 ;
        RECT 133.985 192.905 134.275 192.950 ;
        RECT 128.450 192.610 130.980 192.750 ;
        RECT 128.450 192.550 128.770 192.610 ;
        RECT 132.130 192.550 132.450 192.810 ;
        RECT 132.590 192.550 132.910 192.810 ;
        RECT 23.500 191.930 136.200 192.410 ;
        RECT 27.710 191.530 28.030 191.790 ;
        RECT 38.290 191.530 38.610 191.790 ;
        RECT 48.425 191.730 48.715 191.775 ;
        RECT 50.710 191.730 51.030 191.790 ;
        RECT 48.425 191.590 51.030 191.730 ;
        RECT 48.425 191.545 48.715 191.590 ;
        RECT 50.710 191.530 51.030 191.590 ;
        RECT 67.730 191.530 68.050 191.790 ;
        RECT 78.310 191.730 78.630 191.790 ;
        RECT 81.070 191.730 81.390 191.790 ;
        RECT 78.310 191.590 81.390 191.730 ;
        RECT 78.310 191.530 78.630 191.590 ;
        RECT 81.070 191.530 81.390 191.590 ;
        RECT 87.510 191.530 87.830 191.790 ;
        RECT 91.280 191.590 100.160 191.730 ;
        RECT 91.280 191.450 91.420 191.590 ;
        RECT 48.885 191.390 49.175 191.435 ;
        RECT 67.285 191.390 67.575 191.435 ;
        RECT 69.585 191.390 69.875 191.435 ;
        RECT 48.885 191.250 66.580 191.390 ;
        RECT 48.885 191.205 49.175 191.250 ;
        RECT 41.525 191.050 41.815 191.095 ;
        RECT 44.730 191.050 45.050 191.110 ;
        RECT 41.525 190.910 45.050 191.050 ;
        RECT 41.525 190.865 41.815 190.910 ;
        RECT 44.730 190.850 45.050 190.910 ;
        RECT 53.010 190.850 53.330 191.110 ;
        RECT 56.690 190.850 57.010 191.110 ;
        RECT 26.330 190.510 26.650 190.770 ;
        RECT 28.645 190.710 28.935 190.755 ;
        RECT 34.610 190.710 34.930 190.770 ;
        RECT 28.645 190.570 34.930 190.710 ;
        RECT 28.645 190.525 28.935 190.570 ;
        RECT 34.610 190.510 34.930 190.570 ;
        RECT 44.285 190.710 44.575 190.755 ;
        RECT 45.190 190.710 45.510 190.770 ;
        RECT 44.285 190.570 45.510 190.710 ;
        RECT 44.285 190.525 44.575 190.570 ;
        RECT 45.190 190.510 45.510 190.570 ;
        RECT 47.030 190.510 47.350 190.770 ;
        RECT 50.265 190.710 50.555 190.755 ;
        RECT 50.725 190.710 51.015 190.755 ;
        RECT 50.265 190.570 51.015 190.710 ;
        RECT 50.265 190.525 50.555 190.570 ;
        RECT 50.725 190.525 51.015 190.570 ;
        RECT 51.645 190.525 51.935 190.755 ;
        RECT 40.145 190.370 40.435 190.415 ;
        RECT 41.050 190.370 41.370 190.430 ;
        RECT 40.145 190.230 41.370 190.370 ;
        RECT 40.145 190.185 40.435 190.230 ;
        RECT 41.050 190.170 41.370 190.230 ;
        RECT 43.365 190.370 43.655 190.415 ;
        RECT 43.810 190.370 44.130 190.430 ;
        RECT 43.365 190.230 44.130 190.370 ;
        RECT 43.365 190.185 43.655 190.230 ;
        RECT 43.810 190.170 44.130 190.230 ;
        RECT 48.425 190.370 48.715 190.415 ;
        RECT 48.870 190.370 49.190 190.430 ;
        RECT 48.425 190.230 49.190 190.370 ;
        RECT 51.720 190.370 51.860 190.525 ;
        RECT 52.090 190.510 52.410 190.770 ;
        RECT 53.470 190.510 53.790 190.770 ;
        RECT 59.005 190.710 59.295 190.755 ;
        RECT 64.510 190.710 64.830 190.770 ;
        RECT 59.005 190.570 64.830 190.710 ;
        RECT 59.005 190.525 59.295 190.570 ;
        RECT 64.510 190.510 64.830 190.570 ;
        RECT 65.445 190.525 65.735 190.755 ;
        RECT 52.550 190.370 52.870 190.430 ;
        RECT 58.085 190.370 58.375 190.415 ;
        RECT 51.720 190.230 52.870 190.370 ;
        RECT 48.425 190.185 48.715 190.230 ;
        RECT 48.870 190.170 49.190 190.230 ;
        RECT 52.550 190.170 52.870 190.230 ;
        RECT 55.860 190.230 58.375 190.370 ;
        RECT 65.520 190.370 65.660 190.525 ;
        RECT 65.890 190.510 66.210 190.770 ;
        RECT 66.440 190.710 66.580 191.250 ;
        RECT 67.285 191.250 69.875 191.390 ;
        RECT 67.285 191.205 67.575 191.250 ;
        RECT 69.585 191.205 69.875 191.250 ;
        RECT 76.485 191.390 76.775 191.435 ;
        RECT 82.450 191.390 82.770 191.450 ;
        RECT 76.485 191.250 82.770 191.390 ;
        RECT 76.485 191.205 76.775 191.250 ;
        RECT 82.450 191.190 82.770 191.250 ;
        RECT 85.685 191.390 85.975 191.435 ;
        RECT 91.190 191.390 91.510 191.450 ;
        RECT 85.685 191.250 91.510 191.390 ;
        RECT 85.685 191.205 85.975 191.250 ;
        RECT 91.190 191.190 91.510 191.250 ;
        RECT 92.660 191.250 98.320 191.390 ;
        RECT 76.010 191.050 76.330 191.110 ;
        RECT 80.150 191.050 80.470 191.110 ;
        RECT 92.660 191.050 92.800 191.250 ;
        RECT 94.870 191.050 95.190 191.110 ;
        RECT 73.800 190.910 76.330 191.050 ;
        RECT 67.285 190.710 67.575 190.755 ;
        RECT 66.440 190.570 67.575 190.710 ;
        RECT 67.285 190.525 67.575 190.570 ;
        RECT 68.650 190.510 68.970 190.770 ;
        RECT 69.125 190.710 69.415 190.755 ;
        RECT 70.030 190.710 70.350 190.770 ;
        RECT 69.125 190.570 70.350 190.710 ;
        RECT 69.125 190.525 69.415 190.570 ;
        RECT 70.030 190.510 70.350 190.570 ;
        RECT 70.490 190.510 70.810 190.770 ;
        RECT 73.800 190.710 73.940 190.910 ;
        RECT 76.010 190.850 76.330 190.910 ;
        RECT 76.560 190.910 78.540 191.050 ;
        RECT 71.040 190.570 73.940 190.710 ;
        RECT 74.630 190.710 74.920 190.755 ;
        RECT 75.090 190.710 75.410 190.770 ;
        RECT 74.630 190.570 75.410 190.710 ;
        RECT 71.040 190.370 71.180 190.570 ;
        RECT 74.630 190.525 74.920 190.570 ;
        RECT 75.090 190.510 75.410 190.570 ;
        RECT 65.520 190.230 71.180 190.370 ;
        RECT 19.890 190.030 20.210 190.090 ;
        RECT 25.425 190.030 25.715 190.075 ;
        RECT 19.890 189.890 25.715 190.030 ;
        RECT 19.890 189.830 20.210 189.890 ;
        RECT 25.425 189.845 25.715 189.890 ;
        RECT 40.590 190.030 40.910 190.090 ;
        RECT 42.445 190.030 42.735 190.075 ;
        RECT 40.590 189.890 42.735 190.030 ;
        RECT 40.590 189.830 40.910 189.890 ;
        RECT 42.445 189.845 42.735 189.890 ;
        RECT 46.570 190.030 46.890 190.090 ;
        RECT 47.505 190.030 47.795 190.075 ;
        RECT 49.805 190.030 50.095 190.075 ;
        RECT 46.570 189.890 50.095 190.030 ;
        RECT 46.570 189.830 46.890 189.890 ;
        RECT 47.505 189.845 47.795 189.890 ;
        RECT 49.805 189.845 50.095 189.890 ;
        RECT 51.630 190.030 51.950 190.090 ;
        RECT 53.945 190.030 54.235 190.075 ;
        RECT 51.630 189.890 54.235 190.030 ;
        RECT 51.630 189.830 51.950 189.890 ;
        RECT 53.945 189.845 54.235 189.890 ;
        RECT 55.310 190.030 55.630 190.090 ;
        RECT 55.860 190.075 56.000 190.230 ;
        RECT 58.085 190.185 58.375 190.230 ;
        RECT 71.410 190.170 71.730 190.430 ;
        RECT 76.560 190.370 76.700 190.910 ;
        RECT 78.400 190.770 78.540 190.910 ;
        RECT 80.150 190.910 84.060 191.050 ;
        RECT 80.150 190.850 80.470 190.910 ;
        RECT 76.945 190.525 77.235 190.755 ;
        RECT 74.720 190.230 76.700 190.370 ;
        RECT 74.720 190.090 74.860 190.230 ;
        RECT 55.785 190.030 56.075 190.075 ;
        RECT 55.310 189.890 56.075 190.030 ;
        RECT 55.310 189.830 55.630 189.890 ;
        RECT 55.785 189.845 56.075 189.890 ;
        RECT 56.230 189.830 56.550 190.090 ;
        RECT 64.525 190.030 64.815 190.075 ;
        RECT 66.365 190.030 66.655 190.075 ;
        RECT 66.810 190.030 67.130 190.090 ;
        RECT 64.525 189.890 67.130 190.030 ;
        RECT 64.525 189.845 64.815 189.890 ;
        RECT 66.365 189.845 66.655 189.890 ;
        RECT 66.810 189.830 67.130 189.890 ;
        RECT 70.950 190.030 71.270 190.090 ;
        RECT 73.725 190.030 74.015 190.075 ;
        RECT 70.950 189.890 74.015 190.030 ;
        RECT 70.950 189.830 71.270 189.890 ;
        RECT 73.725 189.845 74.015 189.890 ;
        RECT 74.630 189.830 74.950 190.090 ;
        RECT 76.470 190.030 76.790 190.090 ;
        RECT 77.020 190.030 77.160 190.525 ;
        RECT 78.310 190.510 78.630 190.770 ;
        RECT 78.770 190.710 79.090 190.770 ;
        RECT 82.465 190.710 82.755 190.755 ;
        RECT 78.770 190.570 82.755 190.710 ;
        RECT 78.770 190.510 79.090 190.570 ;
        RECT 82.465 190.525 82.755 190.570 ;
        RECT 83.370 190.510 83.690 190.770 ;
        RECT 83.920 190.755 84.060 190.910 ;
        RECT 89.440 190.910 92.800 191.050 ;
        RECT 83.845 190.710 84.135 190.755 ;
        RECT 85.225 190.710 85.515 190.755 ;
        RECT 83.845 190.570 85.515 190.710 ;
        RECT 83.845 190.525 84.135 190.570 ;
        RECT 85.225 190.525 85.515 190.570 ;
        RECT 86.590 190.510 86.910 190.770 ;
        RECT 88.890 190.710 89.210 190.770 ;
        RECT 89.440 190.755 89.580 190.910 ;
        RECT 89.365 190.710 89.655 190.755 ;
        RECT 88.890 190.570 89.655 190.710 ;
        RECT 88.890 190.510 89.210 190.570 ;
        RECT 89.365 190.525 89.655 190.570 ;
        RECT 90.285 190.710 90.575 190.755 ;
        RECT 92.110 190.710 92.430 190.770 ;
        RECT 92.660 190.755 92.800 190.910 ;
        RECT 93.580 190.910 96.480 191.050 ;
        RECT 90.285 190.570 92.430 190.710 ;
        RECT 90.285 190.525 90.575 190.570 ;
        RECT 92.110 190.510 92.430 190.570 ;
        RECT 92.585 190.525 92.875 190.755 ;
        RECT 93.030 190.710 93.350 190.770 ;
        RECT 93.580 190.755 93.720 190.910 ;
        RECT 94.870 190.850 95.190 190.910 ;
        RECT 96.340 190.760 96.480 190.910 ;
        RECT 96.685 190.760 96.975 190.805 ;
        RECT 93.505 190.710 93.795 190.755 ;
        RECT 93.030 190.570 93.795 190.710 ;
        RECT 79.245 190.370 79.535 190.415 ;
        RECT 81.070 190.370 81.390 190.430 ;
        RECT 79.245 190.230 81.390 190.370 ;
        RECT 79.245 190.185 79.535 190.230 ;
        RECT 81.070 190.170 81.390 190.230 ;
        RECT 81.990 190.370 82.310 190.430 ;
        RECT 86.680 190.370 86.820 190.510 ;
        RECT 91.665 190.370 91.955 190.415 ;
        RECT 81.990 190.230 86.820 190.370 ;
        RECT 89.440 190.230 91.955 190.370 ;
        RECT 92.660 190.370 92.800 190.525 ;
        RECT 93.030 190.510 93.350 190.570 ;
        RECT 93.505 190.525 93.795 190.570 ;
        RECT 94.425 190.525 94.715 190.755 ;
        RECT 95.345 190.525 95.635 190.755 ;
        RECT 96.340 190.620 96.975 190.760 ;
        RECT 98.180 190.755 98.320 191.250 ;
        RECT 100.020 191.050 100.160 191.590 ;
        RECT 100.390 191.530 100.710 191.790 ;
        RECT 106.830 191.730 107.150 191.790 ;
        RECT 111.905 191.730 112.195 191.775 ;
        RECT 106.830 191.590 112.195 191.730 ;
        RECT 106.830 191.530 107.150 191.590 ;
        RECT 111.905 191.545 112.195 191.590 ;
        RECT 112.350 191.730 112.670 191.790 ;
        RECT 125.690 191.730 126.010 191.790 ;
        RECT 112.350 191.590 126.010 191.730 ;
        RECT 112.350 191.530 112.670 191.590 ;
        RECT 125.690 191.530 126.010 191.590 ;
        RECT 127.530 191.730 127.850 191.790 ;
        RECT 128.465 191.730 128.755 191.775 ;
        RECT 127.530 191.590 128.755 191.730 ;
        RECT 127.530 191.530 127.850 191.590 ;
        RECT 128.465 191.545 128.755 191.590 ;
        RECT 104.530 191.390 104.850 191.450 ;
        RECT 104.530 191.250 107.750 191.390 ;
        RECT 104.530 191.190 104.850 191.250 ;
        RECT 107.610 191.050 107.750 191.250 ;
        RECT 133.065 191.205 133.355 191.435 ;
        RECT 100.020 190.910 107.060 191.050 ;
        RECT 107.610 190.910 108.440 191.050 ;
        RECT 106.920 190.770 107.060 190.910 ;
        RECT 108.300 190.770 108.440 190.910 ;
        RECT 108.670 190.850 108.990 191.110 ;
        RECT 109.130 191.050 109.450 191.110 ;
        RECT 113.730 191.050 114.050 191.110 ;
        RECT 114.665 191.050 114.955 191.095 ;
        RECT 116.505 191.050 116.795 191.095 ;
        RECT 121.090 191.050 121.410 191.110 ;
        RECT 133.140 191.050 133.280 191.205 ;
        RECT 109.130 190.910 113.040 191.050 ;
        RECT 109.130 190.850 109.450 190.910 ;
        RECT 96.685 190.575 96.975 190.620 ;
        RECT 98.105 190.525 98.395 190.755 ;
        RECT 99.025 190.710 99.315 190.755 ;
        RECT 99.485 190.710 99.775 190.755 ;
        RECT 99.025 190.570 99.775 190.710 ;
        RECT 99.025 190.525 99.315 190.570 ;
        RECT 99.485 190.525 99.775 190.570 ;
        RECT 94.500 190.370 94.640 190.525 ;
        RECT 92.660 190.230 94.640 190.370 ;
        RECT 95.420 190.370 95.560 190.525 ;
        RECT 97.185 190.370 97.475 190.415 ;
        RECT 99.100 190.370 99.240 190.525 ;
        RECT 102.690 190.510 103.010 190.770 ;
        RECT 106.385 190.525 106.675 190.755 ;
        RECT 106.830 190.710 107.150 190.770 ;
        RECT 107.305 190.710 107.595 190.755 ;
        RECT 106.830 190.570 107.595 190.710 ;
        RECT 95.420 190.230 99.240 190.370 ;
        RECT 81.990 190.170 82.310 190.230 ;
        RECT 89.440 190.090 89.580 190.230 ;
        RECT 91.665 190.185 91.955 190.230 ;
        RECT 97.185 190.185 97.475 190.230 ;
        RECT 77.405 190.030 77.695 190.075 ;
        RECT 76.470 189.890 77.695 190.030 ;
        RECT 76.470 189.830 76.790 189.890 ;
        RECT 77.405 189.845 77.695 189.890 ;
        RECT 89.350 189.830 89.670 190.090 ;
        RECT 90.730 190.030 91.050 190.090 ;
        RECT 91.205 190.030 91.495 190.075 ;
        RECT 90.730 189.890 91.495 190.030 ;
        RECT 90.730 189.830 91.050 189.890 ;
        RECT 91.205 189.845 91.495 189.890 ;
        RECT 95.790 190.030 96.110 190.090 ;
        RECT 96.265 190.030 96.555 190.075 ;
        RECT 95.790 189.890 96.555 190.030 ;
        RECT 95.790 189.830 96.110 189.890 ;
        RECT 96.265 189.845 96.555 189.890 ;
        RECT 96.710 190.030 97.030 190.090 ;
        RECT 98.565 190.030 98.855 190.075 ;
        RECT 96.710 189.890 98.855 190.030 ;
        RECT 106.460 190.030 106.600 190.525 ;
        RECT 106.830 190.510 107.150 190.570 ;
        RECT 107.305 190.525 107.595 190.570 ;
        RECT 108.210 190.510 108.530 190.770 ;
        RECT 108.760 190.710 108.900 190.850 ;
        RECT 110.525 190.710 110.815 190.755 ;
        RECT 110.970 190.710 111.290 190.770 ;
        RECT 108.760 190.570 109.360 190.710 ;
        RECT 109.220 190.415 109.360 190.570 ;
        RECT 110.525 190.570 111.290 190.710 ;
        RECT 110.525 190.525 110.815 190.570 ;
        RECT 110.970 190.510 111.290 190.570 ;
        RECT 111.445 190.710 111.735 190.755 ;
        RECT 111.890 190.710 112.210 190.770 ;
        RECT 112.900 190.755 113.040 190.910 ;
        RECT 113.730 190.910 114.955 191.050 ;
        RECT 113.730 190.850 114.050 190.910 ;
        RECT 114.665 190.865 114.955 190.910 ;
        RECT 115.200 190.910 121.410 191.050 ;
        RECT 111.445 190.570 112.210 190.710 ;
        RECT 111.445 190.525 111.735 190.570 ;
        RECT 111.890 190.510 112.210 190.570 ;
        RECT 112.825 190.525 113.115 190.755 ;
        RECT 113.270 190.710 113.590 190.770 ;
        RECT 115.200 190.710 115.340 190.910 ;
        RECT 116.505 190.865 116.795 190.910 ;
        RECT 121.090 190.850 121.410 190.910 ;
        RECT 131.760 190.910 133.280 191.050 ;
        RECT 113.270 190.570 115.340 190.710 ;
        RECT 113.270 190.510 113.590 190.570 ;
        RECT 115.570 190.510 115.890 190.770 ;
        RECT 123.850 190.710 124.170 190.770 ;
        RECT 127.545 190.710 127.835 190.755 ;
        RECT 123.850 190.570 127.835 190.710 ;
        RECT 123.850 190.510 124.170 190.570 ;
        RECT 127.545 190.525 127.835 190.570 ;
        RECT 130.305 190.710 130.595 190.755 ;
        RECT 131.210 190.710 131.530 190.770 ;
        RECT 131.760 190.755 131.900 190.910 ;
        RECT 130.305 190.570 131.530 190.710 ;
        RECT 130.305 190.525 130.595 190.570 ;
        RECT 131.210 190.510 131.530 190.570 ;
        RECT 131.685 190.525 131.975 190.755 ;
        RECT 132.605 190.710 132.895 190.755 ;
        RECT 133.510 190.710 133.830 190.770 ;
        RECT 132.605 190.570 133.830 190.710 ;
        RECT 132.605 190.525 132.895 190.570 ;
        RECT 133.510 190.510 133.830 190.570 ;
        RECT 134.445 190.710 134.735 190.755 ;
        RECT 134.445 190.570 136.500 190.710 ;
        RECT 134.445 190.525 134.735 190.570 ;
        RECT 109.145 190.185 109.435 190.415 ;
        RECT 109.590 190.170 109.910 190.430 ;
        RECT 117.870 190.170 118.190 190.430 ;
        RECT 123.390 190.370 123.710 190.430 ;
        RECT 118.420 190.230 123.710 190.370 ;
        RECT 118.420 190.030 118.560 190.230 ;
        RECT 123.390 190.170 123.710 190.230 ;
        RECT 124.770 190.370 125.090 190.430 ;
        RECT 133.065 190.370 133.355 190.415 ;
        RECT 124.770 190.230 133.355 190.370 ;
        RECT 124.770 190.170 125.090 190.230 ;
        RECT 133.065 190.185 133.355 190.230 ;
        RECT 106.460 189.890 118.560 190.030 ;
        RECT 118.790 190.030 119.110 190.090 ;
        RECT 124.325 190.030 124.615 190.075 ;
        RECT 118.790 189.890 124.615 190.030 ;
        RECT 96.710 189.830 97.030 189.890 ;
        RECT 98.565 189.845 98.855 189.890 ;
        RECT 118.790 189.830 119.110 189.890 ;
        RECT 124.325 189.845 124.615 189.890 ;
        RECT 129.385 190.030 129.675 190.075 ;
        RECT 130.290 190.030 130.610 190.090 ;
        RECT 129.385 189.890 130.610 190.030 ;
        RECT 129.385 189.845 129.675 189.890 ;
        RECT 130.290 189.830 130.610 189.890 ;
        RECT 133.970 189.830 134.290 190.090 ;
        RECT 23.500 189.210 136.200 189.690 ;
        RECT 26.330 189.010 26.650 189.070 ;
        RECT 27.725 189.010 28.015 189.055 ;
        RECT 26.330 188.870 28.015 189.010 ;
        RECT 26.330 188.810 26.650 188.870 ;
        RECT 27.725 188.825 28.015 188.870 ;
        RECT 39.685 189.010 39.975 189.055 ;
        RECT 40.590 189.010 40.910 189.070 ;
        RECT 39.685 188.870 40.910 189.010 ;
        RECT 39.685 188.825 39.975 188.870 ;
        RECT 40.590 188.810 40.910 188.870 ;
        RECT 46.570 188.810 46.890 189.070 ;
        RECT 47.950 189.010 48.270 189.070 ;
        RECT 52.090 189.010 52.410 189.070 ;
        RECT 47.950 188.870 52.410 189.010 ;
        RECT 47.950 188.810 48.270 188.870 ;
        RECT 52.090 188.810 52.410 188.870 ;
        RECT 53.010 189.010 53.330 189.070 ;
        RECT 58.085 189.010 58.375 189.055 ;
        RECT 53.010 188.870 58.375 189.010 ;
        RECT 53.010 188.810 53.330 188.870 ;
        RECT 58.085 188.825 58.375 188.870 ;
        RECT 60.370 188.810 60.690 189.070 ;
        RECT 75.550 189.010 75.870 189.070 ;
        RECT 78.770 189.010 79.090 189.070 ;
        RECT 80.150 189.010 80.470 189.070 ;
        RECT 81.990 189.010 82.310 189.070 ;
        RECT 75.550 188.870 79.090 189.010 ;
        RECT 75.550 188.810 75.870 188.870 ;
        RECT 78.770 188.810 79.090 188.870 ;
        RECT 79.320 188.870 82.310 189.010 ;
        RECT 43.350 188.670 43.670 188.730 ;
        RECT 56.230 188.670 56.550 188.730 ;
        RECT 63.145 188.670 63.435 188.715 ;
        RECT 67.270 188.670 67.590 188.730 ;
        RECT 43.350 188.530 52.780 188.670 ;
        RECT 43.350 188.470 43.670 188.530 ;
        RECT 28.645 188.145 28.935 188.375 ;
        RECT 40.145 188.330 40.435 188.375 ;
        RECT 41.050 188.330 41.370 188.390 ;
        RECT 40.145 188.190 41.370 188.330 ;
        RECT 40.145 188.145 40.435 188.190 ;
        RECT 28.720 187.310 28.860 188.145 ;
        RECT 41.050 188.130 41.370 188.190 ;
        RECT 44.730 188.130 45.050 188.390 ;
        RECT 45.665 188.145 45.955 188.375 ;
        RECT 40.605 187.990 40.895 188.035 ;
        RECT 44.820 187.990 44.960 188.130 ;
        RECT 40.605 187.850 44.960 187.990 ;
        RECT 45.740 187.990 45.880 188.145 ;
        RECT 47.030 188.130 47.350 188.390 ;
        RECT 47.965 188.145 48.255 188.375 ;
        RECT 46.110 187.990 46.430 188.050 ;
        RECT 48.040 187.990 48.180 188.145 ;
        RECT 51.630 188.130 51.950 188.390 ;
        RECT 52.090 188.130 52.410 188.390 ;
        RECT 52.640 188.330 52.780 188.530 ;
        RECT 56.230 188.530 63.435 188.670 ;
        RECT 56.230 188.470 56.550 188.530 ;
        RECT 63.145 188.485 63.435 188.530 ;
        RECT 65.060 188.530 67.590 188.670 ;
        RECT 53.010 188.375 53.330 188.390 ;
        RECT 53.010 188.330 53.545 188.375 ;
        RECT 52.640 188.190 53.545 188.330 ;
        RECT 53.010 188.145 53.545 188.190 ;
        RECT 55.785 188.330 56.075 188.375 ;
        RECT 59.450 188.330 59.770 188.390 ;
        RECT 55.785 188.190 59.770 188.330 ;
        RECT 55.785 188.145 56.075 188.190 ;
        RECT 53.010 188.130 53.330 188.145 ;
        RECT 59.450 188.130 59.770 188.190 ;
        RECT 59.925 188.330 60.215 188.375 ;
        RECT 61.290 188.330 61.610 188.390 ;
        RECT 59.925 188.190 61.610 188.330 ;
        RECT 59.925 188.145 60.215 188.190 ;
        RECT 61.290 188.130 61.610 188.190 ;
        RECT 62.670 188.130 62.990 188.390 ;
        RECT 63.605 188.330 63.895 188.375 ;
        RECT 64.050 188.330 64.370 188.390 ;
        RECT 65.060 188.375 65.200 188.530 ;
        RECT 67.270 188.470 67.590 188.530 ;
        RECT 69.110 188.670 69.430 188.730 ;
        RECT 69.585 188.670 69.875 188.715 ;
        RECT 69.110 188.530 69.875 188.670 ;
        RECT 69.110 188.470 69.430 188.530 ;
        RECT 69.585 188.485 69.875 188.530 ;
        RECT 63.605 188.190 64.370 188.330 ;
        RECT 63.605 188.145 63.895 188.190 ;
        RECT 64.050 188.130 64.370 188.190 ;
        RECT 64.985 188.145 65.275 188.375 ;
        RECT 65.445 188.145 65.735 188.375 ;
        RECT 66.365 188.330 66.655 188.375 ;
        RECT 70.030 188.330 70.350 188.390 ;
        RECT 66.365 188.190 70.350 188.330 ;
        RECT 66.365 188.145 66.655 188.190 ;
        RECT 56.705 187.990 56.995 188.035 ;
        RECT 60.845 187.990 61.135 188.035 ;
        RECT 45.740 187.850 48.180 187.990 ;
        RECT 51.720 187.850 61.135 187.990 ;
        RECT 40.605 187.805 40.895 187.850 ;
        RECT 46.110 187.790 46.430 187.850 ;
        RECT 37.845 187.650 38.135 187.695 ;
        RECT 41.510 187.650 41.830 187.710 ;
        RECT 37.845 187.510 41.830 187.650 ;
        RECT 37.845 187.465 38.135 187.510 ;
        RECT 41.510 187.450 41.830 187.510 ;
        RECT 47.030 187.650 47.350 187.710 ;
        RECT 51.720 187.650 51.860 187.850 ;
        RECT 56.705 187.805 56.995 187.850 ;
        RECT 60.845 187.805 61.135 187.850 ;
        RECT 47.030 187.510 51.860 187.650 ;
        RECT 52.090 187.650 52.410 187.710 ;
        RECT 65.520 187.650 65.660 188.145 ;
        RECT 70.030 188.130 70.350 188.190 ;
        RECT 70.950 188.130 71.270 188.390 ;
        RECT 71.870 188.330 72.190 188.390 ;
        RECT 79.320 188.330 79.460 188.870 ;
        RECT 80.150 188.810 80.470 188.870 ;
        RECT 81.990 188.810 82.310 188.870 ;
        RECT 82.450 188.810 82.770 189.070 ;
        RECT 83.370 189.010 83.690 189.070 ;
        RECT 101.310 189.010 101.630 189.070 ;
        RECT 136.360 189.010 136.500 190.570 ;
        RECT 83.370 188.870 100.850 189.010 ;
        RECT 83.370 188.810 83.690 188.870 ;
        RECT 79.690 188.670 80.010 188.730 ;
        RECT 84.765 188.670 85.055 188.715 ;
        RECT 92.585 188.670 92.875 188.715 ;
        RECT 79.690 188.530 85.055 188.670 ;
        RECT 79.690 188.470 80.010 188.530 ;
        RECT 84.765 188.485 85.055 188.530 ;
        RECT 90.360 188.530 92.875 188.670 ;
        RECT 90.360 188.390 90.500 188.530 ;
        RECT 92.585 188.485 92.875 188.530 ;
        RECT 71.870 188.190 79.460 188.330 ;
        RECT 71.870 188.130 72.190 188.190 ;
        RECT 80.165 188.145 80.455 188.375 ;
        RECT 81.990 188.330 82.310 188.390 ;
        RECT 84.305 188.330 84.595 188.375 ;
        RECT 81.990 188.190 84.595 188.330 ;
        RECT 67.285 187.990 67.575 188.035 ;
        RECT 69.125 187.990 69.415 188.035 ;
        RECT 67.285 187.850 69.415 187.990 ;
        RECT 67.285 187.805 67.575 187.850 ;
        RECT 69.125 187.805 69.415 187.850 ;
        RECT 70.505 187.990 70.795 188.035 ;
        RECT 71.410 187.990 71.730 188.050 ;
        RECT 70.505 187.850 71.730 187.990 ;
        RECT 70.505 187.805 70.795 187.850 ;
        RECT 71.410 187.790 71.730 187.850 ;
        RECT 79.230 187.990 79.550 188.050 ;
        RECT 80.240 187.990 80.380 188.145 ;
        RECT 81.990 188.130 82.310 188.190 ;
        RECT 84.305 188.145 84.595 188.190 ;
        RECT 88.430 188.330 88.750 188.390 ;
        RECT 89.365 188.330 89.655 188.375 ;
        RECT 88.430 188.190 89.655 188.330 ;
        RECT 88.430 188.130 88.750 188.190 ;
        RECT 89.365 188.145 89.655 188.190 ;
        RECT 90.270 188.130 90.590 188.390 ;
        RECT 90.745 188.330 91.035 188.375 ;
        RECT 92.125 188.330 92.415 188.375 ;
        RECT 90.745 188.190 92.415 188.330 ;
        RECT 92.660 188.330 92.800 188.485 ;
        RECT 93.490 188.470 93.810 188.730 ;
        RECT 96.710 188.470 97.030 188.730 ;
        RECT 100.710 188.670 100.850 188.870 ;
        RECT 101.310 188.870 136.500 189.010 ;
        RECT 101.310 188.810 101.630 188.870 ;
        RECT 104.530 188.670 104.850 188.730 ;
        RECT 97.260 188.530 100.160 188.670 ;
        RECT 100.710 188.530 104.850 188.670 ;
        RECT 95.330 188.330 95.650 188.390 ;
        RECT 95.805 188.330 96.095 188.375 ;
        RECT 92.660 188.190 95.100 188.330 ;
        RECT 90.745 188.145 91.035 188.190 ;
        RECT 92.125 188.145 92.415 188.190 ;
        RECT 79.230 187.850 80.380 187.990 ;
        RECT 79.230 187.790 79.550 187.850 ;
        RECT 80.610 187.790 80.930 188.050 ;
        RECT 81.545 187.990 81.835 188.035 ;
        RECT 85.685 187.990 85.975 188.035 ;
        RECT 92.200 187.990 92.340 188.145 ;
        RECT 94.960 187.990 95.100 188.190 ;
        RECT 95.330 188.190 96.095 188.330 ;
        RECT 95.330 188.130 95.650 188.190 ;
        RECT 95.805 188.145 96.095 188.190 ;
        RECT 96.250 188.330 96.570 188.390 ;
        RECT 97.260 188.330 97.400 188.530 ;
        RECT 96.250 188.190 97.400 188.330 ;
        RECT 96.250 188.130 96.570 188.190 ;
        RECT 97.630 188.130 97.950 188.390 ;
        RECT 98.090 188.130 98.410 188.390 ;
        RECT 99.025 188.145 99.315 188.375 ;
        RECT 99.100 187.990 99.240 188.145 ;
        RECT 99.470 188.130 99.790 188.390 ;
        RECT 100.020 188.330 100.160 188.530 ;
        RECT 104.530 188.470 104.850 188.530 ;
        RECT 105.005 188.670 105.295 188.715 ;
        RECT 108.210 188.670 108.530 188.730 ;
        RECT 140.410 188.670 140.730 188.730 ;
        RECT 105.005 188.530 106.140 188.670 ;
        RECT 105.005 188.485 105.295 188.530 ;
        RECT 101.325 188.330 101.615 188.375 ;
        RECT 100.020 188.190 101.615 188.330 ;
        RECT 101.325 188.145 101.615 188.190 ;
        RECT 101.770 188.130 102.090 188.390 ;
        RECT 102.230 188.330 102.550 188.390 ;
        RECT 103.955 188.330 104.245 188.375 ;
        RECT 102.230 188.320 103.790 188.330 ;
        RECT 103.930 188.320 104.245 188.330 ;
        RECT 102.230 188.190 104.245 188.320 ;
        RECT 102.230 188.130 102.550 188.190 ;
        RECT 103.650 188.180 104.245 188.190 ;
        RECT 103.955 188.145 104.245 188.180 ;
        RECT 105.465 188.145 105.755 188.375 ;
        RECT 106.000 188.330 106.140 188.530 ;
        RECT 107.810 188.530 108.530 188.670 ;
        RECT 106.830 188.330 107.150 188.390 ;
        RECT 107.810 188.375 107.950 188.530 ;
        RECT 108.210 188.470 108.530 188.530 ;
        RECT 128.080 188.530 140.730 188.670 ;
        RECT 106.000 188.190 107.150 188.330 ;
        RECT 81.545 187.850 89.095 187.990 ;
        RECT 92.200 187.850 94.640 187.990 ;
        RECT 94.960 187.850 97.400 187.990 ;
        RECT 81.545 187.805 81.835 187.850 ;
        RECT 85.685 187.805 85.975 187.850 ;
        RECT 52.090 187.510 65.660 187.650 ;
        RECT 75.090 187.650 75.410 187.710 ;
        RECT 82.450 187.650 82.770 187.710 ;
        RECT 75.090 187.510 82.770 187.650 ;
        RECT 47.030 187.450 47.350 187.510 ;
        RECT 52.090 187.450 52.410 187.510 ;
        RECT 75.090 187.450 75.410 187.510 ;
        RECT 82.450 187.450 82.770 187.510 ;
        RECT 87.970 187.650 88.290 187.710 ;
        RECT 88.445 187.650 88.735 187.695 ;
        RECT 87.970 187.510 88.735 187.650 ;
        RECT 88.955 187.650 89.095 187.850 ;
        RECT 94.500 187.650 94.640 187.850 ;
        RECT 94.885 187.650 95.175 187.695 ;
        RECT 88.955 187.510 94.180 187.650 ;
        RECT 94.500 187.510 95.175 187.650 ;
        RECT 97.260 187.650 97.400 187.850 ;
        RECT 98.640 187.850 99.240 187.990 ;
        RECT 98.640 187.650 98.780 187.850 ;
        RECT 103.150 187.790 103.470 188.050 ;
        RECT 105.540 187.990 105.680 188.145 ;
        RECT 106.830 188.130 107.150 188.190 ;
        RECT 107.735 188.145 108.025 188.375 ;
        RECT 111.430 188.330 111.750 188.390 ;
        RECT 108.300 188.190 111.750 188.330 ;
        RECT 108.300 188.050 108.440 188.190 ;
        RECT 111.430 188.130 111.750 188.190 ;
        RECT 114.650 188.330 114.970 188.390 ;
        RECT 116.965 188.330 117.255 188.375 ;
        RECT 114.650 188.190 117.255 188.330 ;
        RECT 114.650 188.130 114.970 188.190 ;
        RECT 116.965 188.145 117.255 188.190 ;
        RECT 117.885 188.330 118.175 188.375 ;
        RECT 118.790 188.330 119.110 188.390 ;
        RECT 117.885 188.190 119.110 188.330 ;
        RECT 117.885 188.145 118.175 188.190 ;
        RECT 118.790 188.130 119.110 188.190 ;
        RECT 121.550 188.330 121.870 188.390 ;
        RECT 128.080 188.375 128.220 188.530 ;
        RECT 140.410 188.470 140.730 188.530 ;
        RECT 125.245 188.330 125.535 188.375 ;
        RECT 121.550 188.190 125.535 188.330 ;
        RECT 121.550 188.130 121.870 188.190 ;
        RECT 125.245 188.145 125.535 188.190 ;
        RECT 128.005 188.145 128.295 188.375 ;
        RECT 129.385 188.145 129.675 188.375 ;
        RECT 130.305 188.145 130.595 188.375 ;
        RECT 130.750 188.330 131.070 188.390 ;
        RECT 131.685 188.330 131.975 188.375 ;
        RECT 130.750 188.190 131.975 188.330 ;
        RECT 103.650 187.850 105.680 187.990 ;
        RECT 97.260 187.510 98.780 187.650 ;
        RECT 101.770 187.650 102.090 187.710 ;
        RECT 103.650 187.650 103.790 187.850 ;
        RECT 108.210 187.790 108.530 188.050 ;
        RECT 108.670 187.990 108.990 188.050 ;
        RECT 124.310 187.990 124.630 188.050 ;
        RECT 129.460 187.990 129.600 188.145 ;
        RECT 108.670 187.850 124.630 187.990 ;
        RECT 108.670 187.790 108.990 187.850 ;
        RECT 124.310 187.790 124.630 187.850 ;
        RECT 128.310 187.850 129.600 187.990 ;
        RECT 101.770 187.510 103.790 187.650 ;
        RECT 105.450 187.650 105.770 187.710 ;
        RECT 106.845 187.650 107.135 187.695 ;
        RECT 105.450 187.510 107.135 187.650 ;
        RECT 87.970 187.450 88.290 187.510 ;
        RECT 88.445 187.465 88.735 187.510 ;
        RECT 38.290 187.310 38.610 187.370 ;
        RECT 42.890 187.310 43.210 187.370 ;
        RECT 28.720 187.170 43.210 187.310 ;
        RECT 38.290 187.110 38.610 187.170 ;
        RECT 42.890 187.110 43.210 187.170 ;
        RECT 48.410 187.310 48.730 187.370 ;
        RECT 48.885 187.310 49.175 187.355 ;
        RECT 48.410 187.170 49.175 187.310 ;
        RECT 48.410 187.110 48.730 187.170 ;
        RECT 48.885 187.125 49.175 187.170 ;
        RECT 49.790 187.310 50.110 187.370 ;
        RECT 50.725 187.310 51.015 187.355 ;
        RECT 49.790 187.170 51.015 187.310 ;
        RECT 49.790 187.110 50.110 187.170 ;
        RECT 50.725 187.125 51.015 187.170 ;
        RECT 53.025 187.310 53.315 187.355 ;
        RECT 53.945 187.310 54.235 187.355 ;
        RECT 53.025 187.170 54.235 187.310 ;
        RECT 53.025 187.125 53.315 187.170 ;
        RECT 53.945 187.125 54.235 187.170 ;
        RECT 54.390 187.310 54.710 187.370 ;
        RECT 67.730 187.310 68.050 187.370 ;
        RECT 54.390 187.170 68.050 187.310 ;
        RECT 54.390 187.110 54.710 187.170 ;
        RECT 67.730 187.110 68.050 187.170 ;
        RECT 68.190 187.110 68.510 187.370 ;
        RECT 76.930 187.310 77.250 187.370 ;
        RECT 78.325 187.310 78.615 187.355 ;
        RECT 76.930 187.170 78.615 187.310 ;
        RECT 76.930 187.110 77.250 187.170 ;
        RECT 78.325 187.125 78.615 187.170 ;
        RECT 87.050 187.310 87.370 187.370 ;
        RECT 93.505 187.310 93.795 187.355 ;
        RECT 87.050 187.170 93.795 187.310 ;
        RECT 94.040 187.310 94.180 187.510 ;
        RECT 94.885 187.465 95.175 187.510 ;
        RECT 101.770 187.450 102.090 187.510 ;
        RECT 105.450 187.450 105.770 187.510 ;
        RECT 106.845 187.465 107.135 187.510 ;
        RECT 98.105 187.310 98.395 187.355 ;
        RECT 94.040 187.170 98.395 187.310 ;
        RECT 87.050 187.110 87.370 187.170 ;
        RECT 93.505 187.125 93.795 187.170 ;
        RECT 98.105 187.125 98.395 187.170 ;
        RECT 100.850 187.310 101.170 187.370 ;
        RECT 104.990 187.310 105.310 187.370 ;
        RECT 100.850 187.170 105.310 187.310 ;
        RECT 100.850 187.110 101.170 187.170 ;
        RECT 104.990 187.110 105.310 187.170 ;
        RECT 106.385 187.310 106.675 187.355 ;
        RECT 107.750 187.310 108.070 187.370 ;
        RECT 106.385 187.170 108.070 187.310 ;
        RECT 106.385 187.125 106.675 187.170 ;
        RECT 107.750 187.110 108.070 187.170 ;
        RECT 110.050 187.310 110.370 187.370 ;
        RECT 110.525 187.310 110.815 187.355 ;
        RECT 126.610 187.310 126.930 187.370 ;
        RECT 110.050 187.170 126.930 187.310 ;
        RECT 110.050 187.110 110.370 187.170 ;
        RECT 110.525 187.125 110.815 187.170 ;
        RECT 126.610 187.110 126.930 187.170 ;
        RECT 127.070 187.310 127.390 187.370 ;
        RECT 128.310 187.310 128.450 187.850 ;
        RECT 129.370 187.650 129.690 187.710 ;
        RECT 130.380 187.650 130.520 188.145 ;
        RECT 130.750 188.130 131.070 188.190 ;
        RECT 131.685 188.145 131.975 188.190 ;
        RECT 133.050 188.130 133.370 188.390 ;
        RECT 129.370 187.510 130.520 187.650 ;
        RECT 132.605 187.650 132.895 187.695 ;
        RECT 134.890 187.650 135.210 187.710 ;
        RECT 132.605 187.510 135.210 187.650 ;
        RECT 129.370 187.450 129.690 187.510 ;
        RECT 132.605 187.465 132.895 187.510 ;
        RECT 134.890 187.450 135.210 187.510 ;
        RECT 127.070 187.170 128.450 187.310 ;
        RECT 131.210 187.310 131.530 187.370 ;
        RECT 133.985 187.310 134.275 187.355 ;
        RECT 131.210 187.170 134.275 187.310 ;
        RECT 127.070 187.110 127.390 187.170 ;
        RECT 131.210 187.110 131.530 187.170 ;
        RECT 133.985 187.125 134.275 187.170 ;
        RECT 23.500 186.490 136.200 186.970 ;
        RECT 33.245 186.290 33.535 186.335 ;
        RECT 47.490 186.290 47.810 186.350 ;
        RECT 33.245 186.150 47.810 186.290 ;
        RECT 33.245 186.105 33.535 186.150 ;
        RECT 47.490 186.090 47.810 186.150 ;
        RECT 52.090 186.090 52.410 186.350 ;
        RECT 52.550 186.290 52.870 186.350 ;
        RECT 53.945 186.290 54.235 186.335 ;
        RECT 52.550 186.150 54.235 186.290 ;
        RECT 52.550 186.090 52.870 186.150 ;
        RECT 53.945 186.105 54.235 186.150 ;
        RECT 60.370 186.090 60.690 186.350 ;
        RECT 65.445 186.290 65.735 186.335 ;
        RECT 65.890 186.290 66.210 186.350 ;
        RECT 65.445 186.150 66.210 186.290 ;
        RECT 65.445 186.105 65.735 186.150 ;
        RECT 65.890 186.090 66.210 186.150 ;
        RECT 70.490 186.290 70.810 186.350 ;
        RECT 72.345 186.290 72.635 186.335 ;
        RECT 70.490 186.150 72.635 186.290 ;
        RECT 70.490 186.090 70.810 186.150 ;
        RECT 72.345 186.105 72.635 186.150 ;
        RECT 76.470 186.090 76.790 186.350 ;
        RECT 85.670 186.290 85.990 186.350 ;
        RECT 80.010 186.150 85.990 186.290 ;
        RECT 35.545 185.950 35.835 185.995 ;
        RECT 36.925 185.950 37.215 185.995 ;
        RECT 44.730 185.950 45.050 186.010 ;
        RECT 35.545 185.810 37.215 185.950 ;
        RECT 35.545 185.765 35.835 185.810 ;
        RECT 36.925 185.765 37.215 185.810 ;
        RECT 40.220 185.810 45.050 185.950 ;
        RECT 40.220 185.655 40.360 185.810 ;
        RECT 44.730 185.750 45.050 185.810 ;
        RECT 49.330 185.750 49.650 186.010 ;
        RECT 60.460 185.950 60.600 186.090 ;
        RECT 56.320 185.810 60.600 185.950 ;
        RECT 62.210 185.950 62.530 186.010 ;
        RECT 64.510 185.950 64.830 186.010 ;
        RECT 73.725 185.950 74.015 185.995 ;
        RECT 80.010 185.950 80.150 186.150 ;
        RECT 85.670 186.090 85.990 186.150 ;
        RECT 93.030 186.090 93.350 186.350 ;
        RECT 93.490 186.290 93.810 186.350 ;
        RECT 95.330 186.290 95.650 186.350 ;
        RECT 93.490 186.150 95.650 186.290 ;
        RECT 93.490 186.090 93.810 186.150 ;
        RECT 95.330 186.090 95.650 186.150 ;
        RECT 97.645 186.290 97.935 186.335 ;
        RECT 99.470 186.290 99.790 186.350 ;
        RECT 97.645 186.150 99.790 186.290 ;
        RECT 97.645 186.105 97.935 186.150 ;
        RECT 99.470 186.090 99.790 186.150 ;
        RECT 99.930 186.290 100.250 186.350 ;
        RECT 100.405 186.290 100.695 186.335 ;
        RECT 99.930 186.150 100.695 186.290 ;
        RECT 99.930 186.090 100.250 186.150 ;
        RECT 100.405 186.105 100.695 186.150 ;
        RECT 101.310 186.090 101.630 186.350 ;
        RECT 104.990 186.090 105.310 186.350 ;
        RECT 106.370 186.090 106.690 186.350 ;
        RECT 110.510 186.090 110.830 186.350 ;
        RECT 116.490 186.290 116.810 186.350 ;
        RECT 117.885 186.290 118.175 186.335 ;
        RECT 111.520 186.150 114.650 186.290 ;
        RECT 81.990 185.950 82.310 186.010 ;
        RECT 62.210 185.810 64.830 185.950 ;
        RECT 40.145 185.425 40.435 185.655 ;
        RECT 43.350 185.610 43.670 185.670 ;
        RECT 44.285 185.610 44.575 185.655 ;
        RECT 54.390 185.610 54.710 185.670 ;
        RECT 56.320 185.655 56.460 185.810 ;
        RECT 62.210 185.750 62.530 185.810 ;
        RECT 64.510 185.750 64.830 185.810 ;
        RECT 71.040 185.810 74.015 185.950 ;
        RECT 41.140 185.470 44.575 185.610 ;
        RECT 34.150 185.070 34.470 185.330 ;
        RECT 34.610 185.070 34.930 185.330 ;
        RECT 36.005 185.270 36.295 185.315 ;
        RECT 39.760 185.270 40.360 185.280 ;
        RECT 41.140 185.270 41.280 185.470 ;
        RECT 43.350 185.410 43.670 185.470 ;
        RECT 44.285 185.425 44.575 185.470 ;
        RECT 45.740 185.470 54.710 185.610 ;
        RECT 45.740 185.330 45.880 185.470 ;
        RECT 54.390 185.410 54.710 185.470 ;
        RECT 56.245 185.425 56.535 185.655 ;
        RECT 56.690 185.410 57.010 185.670 ;
        RECT 62.670 185.610 62.990 185.670 ;
        RECT 64.065 185.610 64.355 185.655 ;
        RECT 65.890 185.610 66.210 185.670 ;
        RECT 71.040 185.655 71.180 185.810 ;
        RECT 73.725 185.765 74.015 185.810 ;
        RECT 76.560 185.810 80.150 185.950 ;
        RECT 80.325 185.810 82.310 185.950 ;
        RECT 60.000 185.470 66.210 185.610 ;
        RECT 36.005 185.140 41.280 185.270 ;
        RECT 36.005 185.130 39.900 185.140 ;
        RECT 40.220 185.130 41.280 185.140 ;
        RECT 36.005 185.085 36.295 185.130 ;
        RECT 41.525 185.085 41.815 185.315 ;
        RECT 41.985 185.270 42.275 185.315 ;
        RECT 42.890 185.270 43.210 185.330 ;
        RECT 43.825 185.270 44.115 185.315 ;
        RECT 41.985 185.130 44.115 185.270 ;
        RECT 41.985 185.085 42.275 185.130 ;
        RECT 36.910 184.930 37.230 184.990 ;
        RECT 39.225 184.930 39.515 184.975 ;
        RECT 36.910 184.790 39.515 184.930 ;
        RECT 41.600 184.930 41.740 185.085 ;
        RECT 42.890 185.070 43.210 185.130 ;
        RECT 43.825 185.085 44.115 185.130 ;
        RECT 44.745 185.270 45.035 185.315 ;
        RECT 45.650 185.270 45.970 185.330 ;
        RECT 44.745 185.130 45.970 185.270 ;
        RECT 44.745 185.085 45.035 185.130 ;
        RECT 44.820 184.930 44.960 185.085 ;
        RECT 45.650 185.070 45.970 185.130 ;
        RECT 46.570 185.070 46.890 185.330 ;
        RECT 47.490 185.270 47.810 185.330 ;
        RECT 47.965 185.270 48.255 185.315 ;
        RECT 47.490 185.130 48.255 185.270 ;
        RECT 47.490 185.070 47.810 185.130 ;
        RECT 47.965 185.085 48.255 185.130 ;
        RECT 48.410 185.070 48.730 185.330 ;
        RECT 49.790 185.070 50.110 185.330 ;
        RECT 51.185 185.270 51.475 185.315 ;
        RECT 59.450 185.270 59.770 185.330 ;
        RECT 60.000 185.315 60.140 185.470 ;
        RECT 62.670 185.410 62.990 185.470 ;
        RECT 64.065 185.425 64.355 185.470 ;
        RECT 65.890 185.410 66.210 185.470 ;
        RECT 70.965 185.425 71.255 185.655 ;
        RECT 75.550 185.610 75.870 185.670 ;
        RECT 71.500 185.470 75.870 185.610 ;
        RECT 51.185 185.130 59.770 185.270 ;
        RECT 51.185 185.085 51.475 185.130 ;
        RECT 41.600 184.790 44.960 184.930 ;
        RECT 36.910 184.730 37.230 184.790 ;
        RECT 39.225 184.745 39.515 184.790 ;
        RECT 38.750 184.390 39.070 184.650 ;
        RECT 41.970 184.590 42.290 184.650 ;
        RECT 42.905 184.590 43.195 184.635 ;
        RECT 41.970 184.450 43.195 184.590 ;
        RECT 41.970 184.390 42.290 184.450 ;
        RECT 42.905 184.405 43.195 184.450 ;
        RECT 46.110 184.390 46.430 184.650 ;
        RECT 48.500 184.590 48.640 185.070 ;
        RECT 48.870 184.930 49.190 184.990 ;
        RECT 49.345 184.930 49.635 184.975 ;
        RECT 51.260 184.930 51.400 185.085 ;
        RECT 59.450 185.070 59.770 185.130 ;
        RECT 59.925 185.085 60.215 185.315 ;
        RECT 60.845 185.085 61.135 185.315 ;
        RECT 48.870 184.790 51.400 184.930 ;
        RECT 58.070 184.930 58.390 184.990 ;
        RECT 60.000 184.930 60.140 185.085 ;
        RECT 58.070 184.790 60.140 184.930 ;
        RECT 60.920 184.930 61.060 185.085 ;
        RECT 63.130 185.070 63.450 185.330 ;
        RECT 63.590 185.070 63.910 185.330 ;
        RECT 64.525 185.270 64.815 185.315 ;
        RECT 64.970 185.270 65.290 185.330 ;
        RECT 64.525 185.130 65.290 185.270 ;
        RECT 64.525 185.085 64.815 185.130 ;
        RECT 64.600 184.930 64.740 185.085 ;
        RECT 64.970 185.070 65.290 185.130 ;
        RECT 69.110 185.070 69.430 185.330 ;
        RECT 70.030 185.070 70.350 185.330 ;
        RECT 70.505 185.270 70.795 185.315 ;
        RECT 71.500 185.270 71.640 185.470 ;
        RECT 75.550 185.410 75.870 185.470 ;
        RECT 70.505 185.130 71.640 185.270 ;
        RECT 70.505 185.085 70.795 185.130 ;
        RECT 71.870 185.070 72.190 185.330 ;
        RECT 72.330 185.270 72.650 185.330 ;
        RECT 74.630 185.270 74.920 185.315 ;
        RECT 76.560 185.270 76.700 185.810 ;
        RECT 76.930 185.410 77.250 185.670 ;
        RECT 77.865 185.610 78.155 185.655 ;
        RECT 80.325 185.610 80.465 185.810 ;
        RECT 81.990 185.750 82.310 185.810 ;
        RECT 93.950 185.950 94.270 186.010 ;
        RECT 98.090 185.950 98.410 186.010 ;
        RECT 93.950 185.810 98.410 185.950 ;
        RECT 93.950 185.750 94.270 185.810 ;
        RECT 98.090 185.750 98.410 185.810 ;
        RECT 99.010 185.750 99.330 186.010 ;
        RECT 103.150 185.950 103.470 186.010 ;
        RECT 100.710 185.810 103.470 185.950 ;
        RECT 77.865 185.470 80.465 185.610 ;
        RECT 80.625 185.610 80.915 185.655 ;
        RECT 87.050 185.610 87.370 185.670 ;
        RECT 100.710 185.610 100.850 185.810 ;
        RECT 103.150 185.750 103.470 185.810 ;
        RECT 104.530 185.750 104.850 186.010 ;
        RECT 106.830 185.950 107.150 186.010 ;
        RECT 109.590 185.950 109.910 186.010 ;
        RECT 106.830 185.810 109.910 185.950 ;
        RECT 106.830 185.750 107.150 185.810 ;
        RECT 109.590 185.750 109.910 185.810 ;
        RECT 80.625 185.470 87.370 185.610 ;
        RECT 77.865 185.425 78.155 185.470 ;
        RECT 80.625 185.425 80.915 185.470 ;
        RECT 87.050 185.410 87.370 185.470 ;
        RECT 99.560 185.470 100.850 185.610 ;
        RECT 101.310 185.610 101.630 185.670 ;
        RECT 102.705 185.610 102.995 185.655 ;
        RECT 105.450 185.610 105.770 185.670 ;
        RECT 101.310 185.470 102.995 185.610 ;
        RECT 72.330 185.130 76.700 185.270 ;
        RECT 72.330 185.070 72.650 185.130 ;
        RECT 74.630 185.085 74.920 185.130 ;
        RECT 77.390 185.070 77.710 185.330 ;
        RECT 78.310 185.070 78.630 185.330 ;
        RECT 79.230 185.270 79.550 185.330 ;
        RECT 85.685 185.270 85.975 185.315 ;
        RECT 79.230 185.130 85.975 185.270 ;
        RECT 79.230 185.070 79.550 185.130 ;
        RECT 85.685 185.085 85.975 185.130 ;
        RECT 90.730 185.270 91.050 185.330 ;
        RECT 92.125 185.270 92.415 185.315 ;
        RECT 90.730 185.130 92.415 185.270 ;
        RECT 90.730 185.070 91.050 185.130 ;
        RECT 92.125 185.085 92.415 185.130 ;
        RECT 92.570 185.270 92.890 185.330 ;
        RECT 93.490 185.270 93.810 185.330 ;
        RECT 92.570 185.130 93.810 185.270 ;
        RECT 92.570 185.070 92.890 185.130 ;
        RECT 93.490 185.070 93.810 185.130 ;
        RECT 93.950 185.270 94.270 185.330 ;
        RECT 94.885 185.270 95.175 185.315 ;
        RECT 93.950 185.130 95.175 185.270 ;
        RECT 93.950 185.070 94.270 185.130 ;
        RECT 94.885 185.085 95.175 185.130 ;
        RECT 95.790 185.070 96.110 185.330 ;
        RECT 96.250 185.070 96.570 185.330 ;
        RECT 96.710 185.315 97.030 185.330 ;
        RECT 96.710 185.085 97.135 185.315 ;
        RECT 98.105 185.270 98.395 185.315 ;
        RECT 98.550 185.270 98.870 185.330 ;
        RECT 99.560 185.315 99.700 185.470 ;
        RECT 101.310 185.410 101.630 185.470 ;
        RECT 102.705 185.425 102.995 185.470 ;
        RECT 103.240 185.470 105.770 185.610 ;
        RECT 103.240 185.330 103.380 185.470 ;
        RECT 105.450 185.410 105.770 185.470 ;
        RECT 98.105 185.130 98.870 185.270 ;
        RECT 98.105 185.085 98.395 185.130 ;
        RECT 96.710 185.070 97.030 185.085 ;
        RECT 98.550 185.070 98.870 185.130 ;
        RECT 99.485 185.085 99.775 185.315 ;
        RECT 100.390 185.070 100.710 185.330 ;
        RECT 100.850 185.270 101.170 185.330 ;
        RECT 100.850 185.250 101.540 185.270 ;
        RECT 101.785 185.250 102.075 185.315 ;
        RECT 100.850 185.130 102.075 185.250 ;
        RECT 100.850 185.070 101.170 185.130 ;
        RECT 101.400 185.110 102.075 185.130 ;
        RECT 101.785 185.085 102.075 185.110 ;
        RECT 103.150 185.070 103.470 185.330 ;
        RECT 103.625 185.270 103.915 185.315 ;
        RECT 103.625 185.130 105.680 185.270 ;
        RECT 103.625 185.085 103.915 185.130 ;
        RECT 60.920 184.790 64.740 184.930 ;
        RECT 69.200 184.930 69.340 185.070 ;
        RECT 82.910 184.930 83.230 184.990 ;
        RECT 69.200 184.790 83.230 184.930 ;
        RECT 48.870 184.730 49.190 184.790 ;
        RECT 49.345 184.745 49.635 184.790 ;
        RECT 58.070 184.730 58.390 184.790 ;
        RECT 82.910 184.730 83.230 184.790 ;
        RECT 84.290 184.930 84.610 184.990 ;
        RECT 105.540 184.930 105.680 185.130 ;
        RECT 105.910 185.070 106.230 185.330 ;
        RECT 107.290 185.070 107.610 185.330 ;
        RECT 107.765 185.270 108.055 185.315 ;
        RECT 108.210 185.270 108.530 185.330 ;
        RECT 107.765 185.130 108.530 185.270 ;
        RECT 107.765 185.085 108.055 185.130 ;
        RECT 108.210 185.070 108.530 185.130 ;
        RECT 108.685 185.270 108.975 185.315 ;
        RECT 109.130 185.270 109.450 185.330 ;
        RECT 111.520 185.315 111.660 186.150 ;
        RECT 111.890 185.750 112.210 186.010 ;
        RECT 114.510 185.950 114.650 186.150 ;
        RECT 116.490 186.150 118.175 186.290 ;
        RECT 116.490 186.090 116.810 186.150 ;
        RECT 117.885 186.105 118.175 186.150 ;
        RECT 121.550 186.090 121.870 186.350 ;
        RECT 133.985 186.290 134.275 186.335 ;
        RECT 137.190 186.290 137.510 186.350 ;
        RECT 133.985 186.150 137.510 186.290 ;
        RECT 133.985 186.105 134.275 186.150 ;
        RECT 137.190 186.090 137.510 186.150 ;
        RECT 122.930 185.950 123.250 186.010 ;
        RECT 114.510 185.810 123.250 185.950 ;
        RECT 122.930 185.750 123.250 185.810 ;
        RECT 111.975 185.315 112.115 185.750 ;
        RECT 129.830 185.610 130.150 185.670 ;
        RECT 115.660 185.470 119.940 185.610 ;
        RECT 108.685 185.130 109.450 185.270 ;
        RECT 108.685 185.085 108.975 185.130 ;
        RECT 109.130 185.070 109.450 185.130 ;
        RECT 111.445 185.085 111.735 185.315 ;
        RECT 111.905 185.085 112.195 185.315 ;
        RECT 112.810 185.070 113.130 185.330 ;
        RECT 113.270 185.070 113.590 185.330 ;
        RECT 113.730 185.270 114.050 185.330 ;
        RECT 114.205 185.270 114.495 185.315 ;
        RECT 113.730 185.130 114.495 185.270 ;
        RECT 113.730 185.070 114.050 185.130 ;
        RECT 114.205 185.085 114.495 185.130 ;
        RECT 115.110 185.070 115.430 185.330 ;
        RECT 115.660 185.315 115.800 185.470 ;
        RECT 115.585 185.085 115.875 185.315 ;
        RECT 116.030 185.270 116.350 185.330 ;
        RECT 118.805 185.270 119.095 185.315 ;
        RECT 116.030 185.130 116.545 185.270 ;
        RECT 118.420 185.130 119.095 185.270 ;
        RECT 119.800 185.270 119.940 185.470 ;
        RECT 129.830 185.470 133.280 185.610 ;
        RECT 129.830 185.410 130.150 185.470 ;
        RECT 127.530 185.270 127.850 185.330 ;
        RECT 119.800 185.130 127.850 185.270 ;
        RECT 116.030 185.070 116.350 185.130 ;
        RECT 116.950 184.930 117.270 184.990 ;
        RECT 84.290 184.790 100.850 184.930 ;
        RECT 105.540 184.790 117.270 184.930 ;
        RECT 84.290 184.730 84.610 184.790 ;
        RECT 50.265 184.590 50.555 184.635 ;
        RECT 48.500 184.450 50.555 184.590 ;
        RECT 50.265 184.405 50.555 184.450 ;
        RECT 55.785 184.590 56.075 184.635 ;
        RECT 61.290 184.590 61.610 184.650 ;
        RECT 55.785 184.450 61.610 184.590 ;
        RECT 55.785 184.405 56.075 184.450 ;
        RECT 61.290 184.390 61.610 184.450 ;
        RECT 63.590 184.590 63.910 184.650 ;
        RECT 73.710 184.590 74.030 184.650 ;
        RECT 63.590 184.450 74.030 184.590 ;
        RECT 63.590 184.390 63.910 184.450 ;
        RECT 73.710 184.390 74.030 184.450 ;
        RECT 74.630 184.390 74.950 184.650 ;
        RECT 75.090 184.590 75.410 184.650 ;
        RECT 77.390 184.590 77.710 184.650 ;
        RECT 75.090 184.450 77.710 184.590 ;
        RECT 75.090 184.390 75.410 184.450 ;
        RECT 77.390 184.390 77.710 184.450 ;
        RECT 78.310 184.590 78.630 184.650 ;
        RECT 79.690 184.590 80.010 184.650 ;
        RECT 81.085 184.590 81.375 184.635 ;
        RECT 78.310 184.450 81.375 184.590 ;
        RECT 78.310 184.390 78.630 184.450 ;
        RECT 79.690 184.390 80.010 184.450 ;
        RECT 81.085 184.405 81.375 184.450 ;
        RECT 81.545 184.590 81.835 184.635 ;
        RECT 81.990 184.590 82.310 184.650 ;
        RECT 81.545 184.450 82.310 184.590 ;
        RECT 81.545 184.405 81.835 184.450 ;
        RECT 81.990 184.390 82.310 184.450 ;
        RECT 83.370 184.390 83.690 184.650 ;
        RECT 83.830 184.390 84.150 184.650 ;
        RECT 86.130 184.390 86.450 184.650 ;
        RECT 91.190 184.390 91.510 184.650 ;
        RECT 100.710 184.590 100.850 184.790 ;
        RECT 116.950 184.730 117.270 184.790 ;
        RECT 117.410 184.730 117.730 184.990 ;
        RECT 102.230 184.590 102.550 184.650 ;
        RECT 100.710 184.450 102.550 184.590 ;
        RECT 102.230 184.390 102.550 184.450 ;
        RECT 104.530 184.590 104.850 184.650 ;
        RECT 107.750 184.590 108.070 184.650 ;
        RECT 104.530 184.450 108.070 184.590 ;
        RECT 104.530 184.390 104.850 184.450 ;
        RECT 107.750 184.390 108.070 184.450 ;
        RECT 109.605 184.590 109.895 184.635 ;
        RECT 112.810 184.590 113.130 184.650 ;
        RECT 109.605 184.450 113.130 184.590 ;
        RECT 109.605 184.405 109.895 184.450 ;
        RECT 112.810 184.390 113.130 184.450 ;
        RECT 114.190 184.590 114.510 184.650 ;
        RECT 118.420 184.590 118.560 185.130 ;
        RECT 118.805 185.085 119.095 185.130 ;
        RECT 127.530 185.070 127.850 185.130 ;
        RECT 128.450 185.270 128.770 185.330 ;
        RECT 129.385 185.270 129.675 185.315 ;
        RECT 128.450 185.130 129.675 185.270 ;
        RECT 128.450 185.070 128.770 185.130 ;
        RECT 129.385 185.085 129.675 185.130 ;
        RECT 130.290 185.070 130.610 185.330 ;
        RECT 131.670 185.070 131.990 185.330 ;
        RECT 133.140 185.315 133.280 185.470 ;
        RECT 133.065 185.085 133.355 185.315 ;
        RECT 128.005 184.930 128.295 184.975 ;
        RECT 128.910 184.930 129.230 184.990 ;
        RECT 128.005 184.790 129.230 184.930 ;
        RECT 128.005 184.745 128.295 184.790 ;
        RECT 128.910 184.730 129.230 184.790 ;
        RECT 114.190 184.450 118.560 184.590 ;
        RECT 119.250 184.590 119.570 184.650 ;
        RECT 124.770 184.590 125.090 184.650 ;
        RECT 119.250 184.450 125.090 184.590 ;
        RECT 114.190 184.390 114.510 184.450 ;
        RECT 119.250 184.390 119.570 184.450 ;
        RECT 124.770 184.390 125.090 184.450 ;
        RECT 132.130 184.590 132.450 184.650 ;
        RECT 132.605 184.590 132.895 184.635 ;
        RECT 132.130 184.450 132.895 184.590 ;
        RECT 132.130 184.390 132.450 184.450 ;
        RECT 132.605 184.405 132.895 184.450 ;
        RECT 23.500 183.770 136.200 184.250 ;
        RECT 34.150 183.570 34.470 183.630 ;
        RECT 35.085 183.570 35.375 183.615 ;
        RECT 34.150 183.430 35.375 183.570 ;
        RECT 34.150 183.370 34.470 183.430 ;
        RECT 35.085 183.385 35.375 183.430 ;
        RECT 36.910 183.370 37.230 183.630 ;
        RECT 37.385 183.570 37.675 183.615 ;
        RECT 38.750 183.570 39.070 183.630 ;
        RECT 39.225 183.570 39.515 183.615 ;
        RECT 41.985 183.570 42.275 183.615 ;
        RECT 37.385 183.430 39.515 183.570 ;
        RECT 37.385 183.385 37.675 183.430 ;
        RECT 38.750 183.370 39.070 183.430 ;
        RECT 39.225 183.385 39.515 183.430 ;
        RECT 39.760 183.430 42.275 183.570 ;
        RECT 38.290 183.230 38.610 183.290 ;
        RECT 39.760 183.230 39.900 183.430 ;
        RECT 41.985 183.385 42.275 183.430 ;
        RECT 44.730 183.570 45.050 183.630 ;
        RECT 56.690 183.570 57.010 183.630 ;
        RECT 44.730 183.430 57.010 183.570 ;
        RECT 44.730 183.370 45.050 183.430 ;
        RECT 56.690 183.370 57.010 183.430 ;
        RECT 57.240 183.430 66.350 183.570 ;
        RECT 45.190 183.230 45.510 183.290 ;
        RECT 53.010 183.230 53.330 183.290 ;
        RECT 57.240 183.230 57.380 183.430 ;
        RECT 66.210 183.290 66.350 183.430 ;
        RECT 67.270 183.370 67.590 183.630 ;
        RECT 76.485 183.385 76.775 183.615 ;
        RECT 78.785 183.570 79.075 183.615 ;
        RECT 80.610 183.570 80.930 183.630 ;
        RECT 86.130 183.570 86.450 183.630 ;
        RECT 78.785 183.430 86.450 183.570 ;
        RECT 78.785 183.385 79.075 183.430 ;
        RECT 38.290 183.090 39.900 183.230 ;
        RECT 41.140 183.090 45.510 183.230 ;
        RECT 38.290 183.030 38.610 183.090 ;
        RECT 37.370 182.890 37.690 182.950 ;
        RECT 41.140 182.935 41.280 183.090 ;
        RECT 45.190 183.030 45.510 183.090 ;
        RECT 45.740 183.090 57.380 183.230 ;
        RECT 62.210 183.230 62.530 183.290 ;
        RECT 63.145 183.230 63.435 183.275 ;
        RECT 62.210 183.090 63.435 183.230 ;
        RECT 66.210 183.230 66.670 183.290 ;
        RECT 70.950 183.230 71.270 183.290 ;
        RECT 66.210 183.090 71.270 183.230 ;
        RECT 76.560 183.230 76.700 183.385 ;
        RECT 80.610 183.370 80.930 183.430 ;
        RECT 86.130 183.370 86.450 183.430 ;
        RECT 88.430 183.370 88.750 183.630 ;
        RECT 90.270 183.570 90.590 183.630 ;
        RECT 93.965 183.570 94.255 183.615 ;
        RECT 90.270 183.430 91.880 183.570 ;
        RECT 90.270 183.370 90.590 183.430 ;
        RECT 79.230 183.230 79.550 183.290 ;
        RECT 91.190 183.275 91.510 183.290 ;
        RECT 76.560 183.090 79.550 183.230 ;
        RECT 40.295 182.890 40.585 182.935 ;
        RECT 37.370 182.750 40.585 182.890 ;
        RECT 37.370 182.690 37.690 182.750 ;
        RECT 40.295 182.705 40.585 182.750 ;
        RECT 41.065 182.890 41.355 182.935 ;
        RECT 41.970 182.890 42.290 182.950 ;
        RECT 41.065 182.750 42.290 182.890 ;
        RECT 41.065 182.705 41.355 182.750 ;
        RECT 41.970 182.690 42.290 182.750 ;
        RECT 42.430 182.690 42.750 182.950 ;
        RECT 42.890 182.890 43.210 182.950 ;
        RECT 45.740 182.890 45.880 183.090 ;
        RECT 53.010 183.030 53.330 183.090 ;
        RECT 62.210 183.030 62.530 183.090 ;
        RECT 63.145 183.045 63.435 183.090 ;
        RECT 66.350 183.030 66.670 183.090 ;
        RECT 70.950 183.030 71.270 183.090 ;
        RECT 79.230 183.030 79.550 183.090 ;
        RECT 90.975 183.045 91.510 183.275 ;
        RECT 91.190 183.030 91.510 183.045 ;
        RECT 42.890 182.750 45.880 182.890 ;
        RECT 46.110 182.890 46.430 182.950 ;
        RECT 47.505 182.890 47.795 182.935 ;
        RECT 46.110 182.750 47.795 182.890 ;
        RECT 42.890 182.690 43.210 182.750 ;
        RECT 46.110 182.690 46.430 182.750 ;
        RECT 47.505 182.705 47.795 182.750 ;
        RECT 50.250 182.690 50.570 182.950 ;
        RECT 51.170 182.690 51.490 182.950 ;
        RECT 63.605 182.705 63.895 182.935 ;
        RECT 64.065 182.705 64.355 182.935 ;
        RECT 64.985 182.890 65.275 182.935 ;
        RECT 65.445 182.890 65.735 182.935 ;
        RECT 64.985 182.750 65.735 182.890 ;
        RECT 64.985 182.705 65.275 182.750 ;
        RECT 65.445 182.705 65.735 182.750 ;
        RECT 65.890 182.890 66.210 182.950 ;
        RECT 67.285 182.890 67.575 182.935 ;
        RECT 75.090 182.890 75.410 182.950 ;
        RECT 75.565 182.890 75.855 182.935 ;
        RECT 65.890 182.750 75.855 182.890 ;
        RECT 38.305 182.550 38.595 182.595 ;
        RECT 44.730 182.550 45.050 182.610 ;
        RECT 62.670 182.550 62.990 182.610 ;
        RECT 63.680 182.550 63.820 182.705 ;
        RECT 38.305 182.410 45.050 182.550 ;
        RECT 38.305 182.365 38.595 182.410 ;
        RECT 44.730 182.350 45.050 182.410 ;
        RECT 48.040 182.410 63.820 182.550 ;
        RECT 64.140 182.550 64.280 182.705 ;
        RECT 65.890 182.690 66.210 182.750 ;
        RECT 67.285 182.705 67.575 182.750 ;
        RECT 75.090 182.690 75.410 182.750 ;
        RECT 75.565 182.705 75.855 182.750 ;
        RECT 76.485 182.705 76.775 182.935 ;
        RECT 77.405 182.705 77.695 182.935 ;
        RECT 80.610 182.890 80.930 182.950 ;
        RECT 81.085 182.890 81.375 182.935 ;
        RECT 80.610 182.750 81.375 182.890 ;
        RECT 64.140 182.410 65.200 182.550 ;
        RECT 47.490 182.210 47.810 182.270 ;
        RECT 48.040 182.255 48.180 182.410 ;
        RECT 62.670 182.350 62.990 182.410 ;
        RECT 65.060 182.270 65.200 182.410 ;
        RECT 66.810 182.350 67.130 182.610 ;
        RECT 73.710 182.550 74.030 182.610 ;
        RECT 76.560 182.550 76.700 182.705 ;
        RECT 73.710 182.410 76.700 182.550 ;
        RECT 73.710 182.350 74.030 182.410 ;
        RECT 47.965 182.210 48.255 182.255 ;
        RECT 47.490 182.070 48.255 182.210 ;
        RECT 47.490 182.010 47.810 182.070 ;
        RECT 47.965 182.025 48.255 182.070 ;
        RECT 48.410 182.210 48.730 182.270 ;
        RECT 50.725 182.210 51.015 182.255 ;
        RECT 48.410 182.070 51.015 182.210 ;
        RECT 48.410 182.010 48.730 182.070 ;
        RECT 50.725 182.025 51.015 182.070 ;
        RECT 58.990 182.210 59.310 182.270 ;
        RECT 62.225 182.210 62.515 182.255 ;
        RECT 58.990 182.070 62.515 182.210 ;
        RECT 58.990 182.010 59.310 182.070 ;
        RECT 62.225 182.025 62.515 182.070 ;
        RECT 64.970 182.010 65.290 182.270 ;
        RECT 67.730 182.210 68.050 182.270 ;
        RECT 77.480 182.210 77.620 182.705 ;
        RECT 80.610 182.690 80.930 182.750 ;
        RECT 81.085 182.705 81.375 182.750 ;
        RECT 82.005 182.890 82.295 182.935 ;
        RECT 84.290 182.890 84.610 182.950 ;
        RECT 82.005 182.750 84.610 182.890 ;
        RECT 82.005 182.705 82.295 182.750 ;
        RECT 84.290 182.690 84.610 182.750 ;
        RECT 89.365 182.705 89.655 182.935 ;
        RECT 78.770 182.350 79.090 182.610 ;
        RECT 65.520 182.070 67.500 182.210 ;
        RECT 42.430 181.870 42.750 181.930 ;
        RECT 45.190 181.870 45.510 181.930 ;
        RECT 46.110 181.870 46.430 181.930 ;
        RECT 56.690 181.870 57.010 181.930 ;
        RECT 42.430 181.730 57.010 181.870 ;
        RECT 42.430 181.670 42.750 181.730 ;
        RECT 45.190 181.670 45.510 181.730 ;
        RECT 46.110 181.670 46.430 181.730 ;
        RECT 56.690 181.670 57.010 181.730 ;
        RECT 60.830 181.870 61.150 181.930 ;
        RECT 65.520 181.870 65.660 182.070 ;
        RECT 60.830 181.730 65.660 181.870 ;
        RECT 60.830 181.670 61.150 181.730 ;
        RECT 65.890 181.670 66.210 181.930 ;
        RECT 67.360 181.870 67.500 182.070 ;
        RECT 67.730 182.070 77.620 182.210 ;
        RECT 89.440 182.210 89.580 182.705 ;
        RECT 89.810 182.690 90.130 182.950 ;
        RECT 91.740 182.935 91.880 183.430 ;
        RECT 93.965 183.430 96.940 183.570 ;
        RECT 93.965 183.385 94.255 183.430 ;
        RECT 96.250 183.230 96.570 183.290 ;
        RECT 95.420 183.090 96.570 183.230 ;
        RECT 90.285 182.705 90.575 182.935 ;
        RECT 91.665 182.705 91.955 182.935 ;
        RECT 93.045 182.705 93.335 182.935 ;
        RECT 90.360 182.550 90.500 182.705 ;
        RECT 90.730 182.550 91.050 182.610 ;
        RECT 90.360 182.410 91.050 182.550 ;
        RECT 90.730 182.350 91.050 182.410 ;
        RECT 92.570 182.550 92.890 182.610 ;
        RECT 93.120 182.550 93.260 182.705 ;
        RECT 94.410 182.690 94.730 182.950 ;
        RECT 95.420 182.935 95.560 183.090 ;
        RECT 96.250 183.030 96.570 183.090 ;
        RECT 95.345 182.705 95.635 182.935 ;
        RECT 95.790 182.690 96.110 182.950 ;
        RECT 92.570 182.410 93.260 182.550 ;
        RECT 92.570 182.350 92.890 182.410 ;
        RECT 96.265 182.365 96.555 182.595 ;
        RECT 96.800 182.550 96.940 183.430 ;
        RECT 97.170 183.370 97.490 183.630 ;
        RECT 98.090 183.370 98.410 183.630 ;
        RECT 104.070 183.570 104.390 183.630 ;
        RECT 101.400 183.430 104.390 183.570 ;
        RECT 97.260 183.230 97.400 183.370 ;
        RECT 99.945 183.230 100.235 183.275 ;
        RECT 97.260 183.090 100.235 183.230 ;
        RECT 99.945 183.045 100.235 183.090 ;
        RECT 97.170 182.690 97.490 182.950 ;
        RECT 99.485 182.705 99.775 182.935 ;
        RECT 99.560 182.550 99.700 182.705 ;
        RECT 100.390 182.690 100.710 182.950 ;
        RECT 101.400 182.935 101.540 183.430 ;
        RECT 104.070 183.370 104.390 183.430 ;
        RECT 104.545 183.570 104.835 183.615 ;
        RECT 110.065 183.570 110.355 183.615 ;
        RECT 111.430 183.570 111.750 183.630 ;
        RECT 104.545 183.430 111.750 183.570 ;
        RECT 104.545 183.385 104.835 183.430 ;
        RECT 110.065 183.385 110.355 183.430 ;
        RECT 111.430 183.370 111.750 183.430 ;
        RECT 113.745 183.570 114.035 183.615 ;
        RECT 123.390 183.570 123.710 183.630 ;
        RECT 123.865 183.570 124.155 183.615 ;
        RECT 113.745 183.430 119.480 183.570 ;
        RECT 113.745 183.385 114.035 183.430 ;
        RECT 102.230 183.230 102.550 183.290 ;
        RECT 105.910 183.230 106.230 183.290 ;
        RECT 106.845 183.230 107.135 183.275 ;
        RECT 107.750 183.230 108.070 183.290 ;
        RECT 109.590 183.275 109.910 183.290 ;
        RECT 102.230 183.090 105.680 183.230 ;
        RECT 102.230 183.030 102.550 183.090 ;
        RECT 101.325 182.705 101.615 182.935 ;
        RECT 102.690 182.690 103.010 182.950 ;
        RECT 103.610 182.690 103.930 182.950 ;
        RECT 104.085 182.705 104.375 182.935 ;
        RECT 104.530 182.890 104.850 182.950 ;
        RECT 105.540 182.935 105.680 183.090 ;
        RECT 105.910 183.090 107.135 183.230 ;
        RECT 105.910 183.030 106.230 183.090 ;
        RECT 106.845 183.045 107.135 183.090 ;
        RECT 107.380 183.090 108.070 183.230 ;
        RECT 105.005 182.890 105.295 182.935 ;
        RECT 104.530 182.750 105.295 182.890 ;
        RECT 100.850 182.550 101.170 182.610 ;
        RECT 96.800 182.410 101.170 182.550 ;
        RECT 104.160 182.550 104.300 182.705 ;
        RECT 104.530 182.690 104.850 182.750 ;
        RECT 105.005 182.705 105.295 182.750 ;
        RECT 105.465 182.705 105.755 182.935 ;
        RECT 106.370 182.690 106.690 182.950 ;
        RECT 107.380 182.935 107.520 183.090 ;
        RECT 107.750 183.030 108.070 183.090 ;
        RECT 109.515 183.045 109.910 183.275 ;
        RECT 109.590 183.030 109.910 183.045 ;
        RECT 107.305 182.705 107.595 182.935 ;
        RECT 108.685 182.705 108.975 182.935 ;
        RECT 110.525 182.890 110.815 182.935 ;
        RECT 110.970 182.890 111.290 182.950 ;
        RECT 110.525 182.750 111.290 182.890 ;
        RECT 111.520 182.890 111.660 183.370 ;
        RECT 112.810 183.230 113.130 183.290 ;
        RECT 112.810 183.090 116.260 183.230 ;
        RECT 112.810 183.030 113.130 183.090 ;
        RECT 116.120 182.935 116.260 183.090 ;
        RECT 113.745 182.890 114.035 182.935 ;
        RECT 115.585 182.890 115.875 182.935 ;
        RECT 111.520 182.750 114.035 182.890 ;
        RECT 110.525 182.705 110.815 182.750 ;
        RECT 108.760 182.550 108.900 182.705 ;
        RECT 110.970 182.690 111.290 182.750 ;
        RECT 113.745 182.705 114.035 182.750 ;
        RECT 114.280 182.750 115.875 182.890 ;
        RECT 111.445 182.550 111.735 182.595 ;
        RECT 111.905 182.550 112.195 182.595 ;
        RECT 114.280 182.550 114.420 182.750 ;
        RECT 115.585 182.705 115.875 182.750 ;
        RECT 116.045 182.890 116.335 182.935 ;
        RECT 116.490 182.890 116.810 182.950 ;
        RECT 116.045 182.750 116.810 182.890 ;
        RECT 116.045 182.705 116.335 182.750 ;
        RECT 116.490 182.690 116.810 182.750 ;
        RECT 117.655 182.890 117.945 182.935 ;
        RECT 118.790 182.890 119.110 182.950 ;
        RECT 117.655 182.750 119.110 182.890 ;
        RECT 117.655 182.705 117.945 182.750 ;
        RECT 118.790 182.690 119.110 182.750 ;
        RECT 104.160 182.410 105.215 182.550 ;
        RECT 108.760 182.410 110.740 182.550 ;
        RECT 94.410 182.210 94.730 182.270 ;
        RECT 89.440 182.070 94.730 182.210 ;
        RECT 67.730 182.010 68.050 182.070 ;
        RECT 94.410 182.010 94.730 182.070 ;
        RECT 77.390 181.870 77.710 181.930 ;
        RECT 67.360 181.730 77.710 181.870 ;
        RECT 77.390 181.670 77.710 181.730 ;
        RECT 77.850 181.670 78.170 181.930 ;
        RECT 81.545 181.870 81.835 181.915 ;
        RECT 84.750 181.870 85.070 181.930 ;
        RECT 81.545 181.730 85.070 181.870 ;
        RECT 81.545 181.685 81.835 181.730 ;
        RECT 84.750 181.670 85.070 181.730 ;
        RECT 87.050 181.870 87.370 181.930 ;
        RECT 96.340 181.870 96.480 182.365 ;
        RECT 100.850 182.350 101.170 182.410 ;
        RECT 105.075 182.270 105.215 182.410 ;
        RECT 110.600 182.270 110.740 182.410 ;
        RECT 111.445 182.410 112.195 182.550 ;
        RECT 111.445 182.365 111.735 182.410 ;
        RECT 111.905 182.365 112.195 182.410 ;
        RECT 112.440 182.410 114.420 182.550 ;
        RECT 102.230 182.010 102.550 182.270 ;
        RECT 104.990 182.010 105.310 182.270 ;
        RECT 105.910 182.210 106.230 182.270 ;
        RECT 108.670 182.210 108.990 182.270 ;
        RECT 105.910 182.070 108.990 182.210 ;
        RECT 105.910 182.010 106.230 182.070 ;
        RECT 108.670 182.010 108.990 182.070 ;
        RECT 110.510 182.010 110.830 182.270 ;
        RECT 110.970 182.210 111.290 182.270 ;
        RECT 112.440 182.210 112.580 182.410 ;
        RECT 114.665 182.365 114.955 182.595 ;
        RECT 116.950 182.550 117.270 182.610 ;
        RECT 118.345 182.550 118.635 182.595 ;
        RECT 116.950 182.410 118.635 182.550 ;
        RECT 119.340 182.550 119.480 183.430 ;
        RECT 123.390 183.430 124.155 183.570 ;
        RECT 123.390 183.370 123.710 183.430 ;
        RECT 123.865 183.385 124.155 183.430 ;
        RECT 124.770 183.370 125.090 183.630 ;
        RECT 133.065 183.570 133.355 183.615 ;
        RECT 133.970 183.570 134.290 183.630 ;
        RECT 125.320 183.430 132.360 183.570 ;
        RECT 120.185 183.230 120.475 183.275 ;
        RECT 122.025 183.230 122.315 183.275 ;
        RECT 120.185 183.090 122.315 183.230 ;
        RECT 120.185 183.045 120.475 183.090 ;
        RECT 122.025 183.045 122.315 183.090 ;
        RECT 122.470 183.030 122.790 183.290 ;
        RECT 124.310 183.230 124.630 183.290 ;
        RECT 125.320 183.230 125.460 183.430 ;
        RECT 124.310 183.090 125.460 183.230 ;
        RECT 126.150 183.230 126.470 183.290 ;
        RECT 132.220 183.230 132.360 183.430 ;
        RECT 133.065 183.430 134.290 183.570 ;
        RECT 133.065 183.385 133.355 183.430 ;
        RECT 133.970 183.370 134.290 183.430 ;
        RECT 126.150 183.090 130.520 183.230 ;
        RECT 132.220 183.090 132.820 183.230 ;
        RECT 124.310 183.030 124.630 183.090 ;
        RECT 126.150 183.030 126.470 183.090 ;
        RECT 119.710 182.890 120.030 182.950 ;
        RECT 122.930 182.935 123.250 182.950 ;
        RECT 120.645 182.890 120.935 182.935 ;
        RECT 119.710 182.750 120.935 182.890 ;
        RECT 119.710 182.690 120.030 182.750 ;
        RECT 120.645 182.705 120.935 182.750 ;
        RECT 121.110 182.705 121.400 182.935 ;
        RECT 122.930 182.890 123.260 182.935 ;
        RECT 122.930 182.750 123.445 182.890 ;
        RECT 122.930 182.705 123.260 182.750 ;
        RECT 121.185 182.550 121.325 182.705 ;
        RECT 122.930 182.690 123.250 182.705 ;
        RECT 125.690 182.690 126.010 182.950 ;
        RECT 126.610 182.890 126.930 182.950 ;
        RECT 127.085 182.890 127.375 182.935 ;
        RECT 126.610 182.750 127.375 182.890 ;
        RECT 126.610 182.690 126.930 182.750 ;
        RECT 127.085 182.705 127.375 182.750 ;
        RECT 127.530 182.890 127.850 182.950 ;
        RECT 128.005 182.890 128.295 182.935 ;
        RECT 127.530 182.750 128.295 182.890 ;
        RECT 127.530 182.690 127.850 182.750 ;
        RECT 128.005 182.705 128.295 182.750 ;
        RECT 129.370 182.690 129.690 182.950 ;
        RECT 130.380 182.935 130.520 183.090 ;
        RECT 130.305 182.705 130.595 182.935 ;
        RECT 131.685 182.890 131.975 182.935 ;
        RECT 132.130 182.890 132.450 182.950 ;
        RECT 132.680 182.935 132.820 183.090 ;
        RECT 131.685 182.750 132.450 182.890 ;
        RECT 131.685 182.705 131.975 182.750 ;
        RECT 132.130 182.690 132.450 182.750 ;
        RECT 132.605 182.705 132.895 182.935 ;
        RECT 133.985 182.890 134.275 182.935 ;
        RECT 139.030 182.890 139.350 182.950 ;
        RECT 133.985 182.750 139.350 182.890 ;
        RECT 133.985 182.705 134.275 182.750 ;
        RECT 139.030 182.690 139.350 182.750 ;
        RECT 119.340 182.410 121.325 182.550 ;
        RECT 110.970 182.070 112.580 182.210 ;
        RECT 114.740 182.210 114.880 182.365 ;
        RECT 116.950 182.350 117.270 182.410 ;
        RECT 118.345 182.365 118.635 182.410 ;
        RECT 128.465 182.210 128.755 182.255 ;
        RECT 114.740 182.070 128.755 182.210 ;
        RECT 110.970 182.010 111.290 182.070 ;
        RECT 128.465 182.025 128.755 182.070 ;
        RECT 87.050 181.730 96.480 181.870 ;
        RECT 101.310 181.870 101.630 181.930 ;
        RECT 102.690 181.870 103.010 181.930 ;
        RECT 101.310 181.730 103.010 181.870 ;
        RECT 87.050 181.670 87.370 181.730 ;
        RECT 101.310 181.670 101.630 181.730 ;
        RECT 102.690 181.670 103.010 181.730 ;
        RECT 103.165 181.870 103.455 181.915 ;
        RECT 107.750 181.870 108.070 181.930 ;
        RECT 103.165 181.730 108.070 181.870 ;
        RECT 103.165 181.685 103.455 181.730 ;
        RECT 107.750 181.670 108.070 181.730 ;
        RECT 108.225 181.870 108.515 181.915 ;
        RECT 109.130 181.870 109.450 181.930 ;
        RECT 108.225 181.730 109.450 181.870 ;
        RECT 108.225 181.685 108.515 181.730 ;
        RECT 109.130 181.670 109.450 181.730 ;
        RECT 23.500 181.050 136.200 181.530 ;
        RECT 35.545 180.850 35.835 180.895 ;
        RECT 36.910 180.850 37.230 180.910 ;
        RECT 35.545 180.710 37.230 180.850 ;
        RECT 35.545 180.665 35.835 180.710 ;
        RECT 36.910 180.650 37.230 180.710 ;
        RECT 39.685 180.850 39.975 180.895 ;
        RECT 41.050 180.850 41.370 180.910 ;
        RECT 39.685 180.710 41.370 180.850 ;
        RECT 39.685 180.665 39.975 180.710 ;
        RECT 41.050 180.650 41.370 180.710 ;
        RECT 44.730 180.850 45.050 180.910 ;
        RECT 45.205 180.850 45.495 180.895 ;
        RECT 44.730 180.710 45.495 180.850 ;
        RECT 44.730 180.650 45.050 180.710 ;
        RECT 45.205 180.665 45.495 180.710 ;
        RECT 47.030 180.850 47.350 180.910 ;
        RECT 48.425 180.850 48.715 180.895 ;
        RECT 47.030 180.710 48.715 180.850 ;
        RECT 47.030 180.650 47.350 180.710 ;
        RECT 48.425 180.665 48.715 180.710 ;
        RECT 52.090 180.850 52.410 180.910 ;
        RECT 53.930 180.850 54.250 180.910 ;
        RECT 56.705 180.850 56.995 180.895 ;
        RECT 62.685 180.850 62.975 180.895 ;
        RECT 63.130 180.850 63.450 180.910 ;
        RECT 52.090 180.710 60.600 180.850 ;
        RECT 52.090 180.650 52.410 180.710 ;
        RECT 53.930 180.650 54.250 180.710 ;
        RECT 56.705 180.665 56.995 180.710 ;
        RECT 34.610 180.510 34.930 180.570 ;
        RECT 35.085 180.510 35.375 180.555 ;
        RECT 39.225 180.510 39.515 180.555 ;
        RECT 46.110 180.510 46.430 180.570 ;
        RECT 34.610 180.370 39.515 180.510 ;
        RECT 34.610 180.310 34.930 180.370 ;
        RECT 35.085 180.325 35.375 180.370 ;
        RECT 39.225 180.325 39.515 180.370 ;
        RECT 39.760 180.370 46.430 180.510 ;
        RECT 36.005 180.170 36.295 180.215 ;
        RECT 39.760 180.170 39.900 180.370 ;
        RECT 46.110 180.310 46.430 180.370 ;
        RECT 49.805 180.510 50.095 180.555 ;
        RECT 50.250 180.510 50.570 180.570 ;
        RECT 52.565 180.510 52.855 180.555 ;
        RECT 49.805 180.370 52.855 180.510 ;
        RECT 49.805 180.325 50.095 180.370 ;
        RECT 50.250 180.310 50.570 180.370 ;
        RECT 52.565 180.325 52.855 180.370 ;
        RECT 57.165 180.325 57.455 180.555 ;
        RECT 36.005 180.030 39.900 180.170 ;
        RECT 36.005 179.985 36.295 180.030 ;
        RECT 40.130 179.970 40.450 180.230 ;
        RECT 44.730 180.170 45.050 180.230 ;
        RECT 47.505 180.170 47.795 180.215 ;
        RECT 44.730 180.030 47.795 180.170 ;
        RECT 44.730 179.970 45.050 180.030 ;
        RECT 47.505 179.985 47.795 180.030 ;
        RECT 47.965 180.170 48.255 180.215 ;
        RECT 50.725 180.170 51.015 180.215 ;
        RECT 57.240 180.170 57.380 180.325 ;
        RECT 47.965 180.030 57.380 180.170 ;
        RECT 47.965 179.985 48.255 180.030 ;
        RECT 50.725 179.985 51.015 180.030 ;
        RECT 57.625 179.985 57.915 180.215 ;
        RECT 19.890 179.830 20.210 179.890 ;
        RECT 24.965 179.830 25.255 179.875 ;
        RECT 19.890 179.690 25.255 179.830 ;
        RECT 19.890 179.630 20.210 179.690 ;
        RECT 24.965 179.645 25.255 179.690 ;
        RECT 26.345 179.830 26.635 179.875 ;
        RECT 27.710 179.830 28.030 179.890 ;
        RECT 26.345 179.690 28.030 179.830 ;
        RECT 26.345 179.645 26.635 179.690 ;
        RECT 27.710 179.630 28.030 179.690 ;
        RECT 34.625 179.645 34.915 179.875 ;
        RECT 34.700 179.490 34.840 179.645 ;
        RECT 36.910 179.630 37.230 179.890 ;
        RECT 38.750 179.630 39.070 179.890 ;
        RECT 40.605 179.645 40.895 179.875 ;
        RECT 38.840 179.490 38.980 179.630 ;
        RECT 34.700 179.350 38.980 179.490 ;
        RECT 40.680 179.490 40.820 179.645 ;
        RECT 41.050 179.630 41.370 179.890 ;
        RECT 46.125 179.645 46.415 179.875 ;
        RECT 46.585 179.830 46.875 179.875 ;
        RECT 48.410 179.830 48.730 179.890 ;
        RECT 46.585 179.690 48.730 179.830 ;
        RECT 46.585 179.645 46.875 179.690 ;
        RECT 41.510 179.490 41.830 179.550 ;
        RECT 40.680 179.350 41.830 179.490 ;
        RECT 46.200 179.490 46.340 179.645 ;
        RECT 48.410 179.630 48.730 179.690 ;
        RECT 49.345 179.645 49.635 179.875 ;
        RECT 50.265 179.645 50.555 179.875 ;
        RECT 48.870 179.490 49.190 179.550 ;
        RECT 49.420 179.490 49.560 179.645 ;
        RECT 46.200 179.350 49.560 179.490 ;
        RECT 50.340 179.490 50.480 179.645 ;
        RECT 51.630 179.630 51.950 179.890 ;
        RECT 52.090 179.630 52.410 179.890 ;
        RECT 53.025 179.830 53.315 179.875 ;
        RECT 53.025 179.690 54.620 179.830 ;
        RECT 53.025 179.645 53.315 179.690 ;
        RECT 51.170 179.490 51.490 179.550 ;
        RECT 53.945 179.490 54.235 179.535 ;
        RECT 50.340 179.350 54.235 179.490 ;
        RECT 41.510 179.290 41.830 179.350 ;
        RECT 48.870 179.290 49.190 179.350 ;
        RECT 51.170 179.290 51.490 179.350 ;
        RECT 53.945 179.305 54.235 179.350 ;
        RECT 37.370 179.150 37.690 179.210 ;
        RECT 37.845 179.150 38.135 179.195 ;
        RECT 37.370 179.010 38.135 179.150 ;
        RECT 54.480 179.150 54.620 179.690 ;
        RECT 54.865 179.645 55.155 179.875 ;
        RECT 55.770 179.830 56.090 179.890 ;
        RECT 56.245 179.830 56.535 179.875 ;
        RECT 55.770 179.690 56.535 179.830 ;
        RECT 57.700 179.830 57.840 179.985 ;
        RECT 58.070 179.830 58.390 179.890 ;
        RECT 60.460 179.875 60.600 180.710 ;
        RECT 62.685 180.710 63.450 180.850 ;
        RECT 62.685 180.665 62.975 180.710 ;
        RECT 63.130 180.650 63.450 180.710 ;
        RECT 65.430 180.850 65.750 180.910 ;
        RECT 68.190 180.850 68.510 180.910 ;
        RECT 65.430 180.710 68.510 180.850 ;
        RECT 65.430 180.650 65.750 180.710 ;
        RECT 68.190 180.650 68.510 180.710 ;
        RECT 78.310 180.650 78.630 180.910 ;
        RECT 83.830 180.850 84.150 180.910 ;
        RECT 81.160 180.710 84.150 180.850 ;
        RECT 61.765 180.510 62.055 180.555 ;
        RECT 62.210 180.510 62.530 180.570 ;
        RECT 69.570 180.510 69.890 180.570 ;
        RECT 61.765 180.370 62.530 180.510 ;
        RECT 61.765 180.325 62.055 180.370 ;
        RECT 62.210 180.310 62.530 180.370 ;
        RECT 63.680 180.370 69.890 180.510 ;
        RECT 63.680 180.170 63.820 180.370 ;
        RECT 69.570 180.310 69.890 180.370 ;
        RECT 80.610 180.310 80.930 180.570 ;
        RECT 81.160 180.555 81.300 180.710 ;
        RECT 83.830 180.650 84.150 180.710 ;
        RECT 93.950 180.650 94.270 180.910 ;
        RECT 94.870 180.650 95.190 180.910 ;
        RECT 95.805 180.665 96.095 180.895 ;
        RECT 103.150 180.850 103.470 180.910 ;
        RECT 105.910 180.850 106.230 180.910 ;
        RECT 107.750 180.850 108.070 180.910 ;
        RECT 110.970 180.850 111.290 180.910 ;
        RECT 111.890 180.850 112.210 180.910 ;
        RECT 103.150 180.710 106.230 180.850 ;
        RECT 81.085 180.325 81.375 180.555 ;
        RECT 83.370 180.510 83.690 180.570 ;
        RECT 84.305 180.510 84.595 180.555 ;
        RECT 83.370 180.370 84.595 180.510 ;
        RECT 83.370 180.310 83.690 180.370 ;
        RECT 84.305 180.325 84.595 180.370 ;
        RECT 89.810 180.510 90.130 180.570 ;
        RECT 95.880 180.510 96.020 180.665 ;
        RECT 103.150 180.650 103.470 180.710 ;
        RECT 105.910 180.650 106.230 180.710 ;
        RECT 106.460 180.710 107.520 180.850 ;
        RECT 98.105 180.510 98.395 180.555 ;
        RECT 89.810 180.370 98.395 180.510 ;
        RECT 89.810 180.310 90.130 180.370 ;
        RECT 98.105 180.325 98.395 180.370 ;
        RECT 61.840 180.030 63.820 180.170 ;
        RECT 64.050 180.170 64.370 180.230 ;
        RECT 65.905 180.170 66.195 180.215 ;
        RECT 70.950 180.170 71.270 180.230 ;
        RECT 64.050 180.030 66.195 180.170 ;
        RECT 57.700 179.690 58.390 179.830 ;
        RECT 54.940 179.490 55.080 179.645 ;
        RECT 55.770 179.630 56.090 179.690 ;
        RECT 56.245 179.645 56.535 179.690 ;
        RECT 58.070 179.630 58.390 179.690 ;
        RECT 58.620 179.690 60.140 179.830 ;
        RECT 55.310 179.490 55.630 179.550 ;
        RECT 58.620 179.490 58.760 179.690 ;
        RECT 60.000 179.550 60.140 179.690 ;
        RECT 60.385 179.645 60.675 179.875 ;
        RECT 60.830 179.630 61.150 179.890 ;
        RECT 61.840 179.875 61.980 180.030 ;
        RECT 64.050 179.970 64.370 180.030 ;
        RECT 65.905 179.985 66.195 180.030 ;
        RECT 69.200 180.030 71.270 180.170 ;
        RECT 61.765 179.645 62.055 179.875 ;
        RECT 63.590 179.630 63.910 179.890 ;
        RECT 67.270 179.875 67.590 179.890 ;
        RECT 69.200 179.875 69.340 180.030 ;
        RECT 70.950 179.970 71.270 180.030 ;
        RECT 76.470 180.170 76.790 180.230 ;
        RECT 78.785 180.170 79.075 180.215 ;
        RECT 86.145 180.170 86.435 180.215 ;
        RECT 76.470 180.030 79.075 180.170 ;
        RECT 76.470 179.970 76.790 180.030 ;
        RECT 78.785 179.985 79.075 180.030 ;
        RECT 81.620 180.030 86.435 180.170 ;
        RECT 69.570 179.875 69.890 179.890 ;
        RECT 65.215 179.830 65.505 179.875 ;
        RECT 67.260 179.830 67.590 179.875 ;
        RECT 65.215 179.690 66.580 179.830 ;
        RECT 67.075 179.690 67.590 179.830 ;
        RECT 65.215 179.645 65.505 179.690 ;
        RECT 54.940 179.350 58.760 179.490 ;
        RECT 55.310 179.290 55.630 179.350 ;
        RECT 58.990 179.290 59.310 179.550 ;
        RECT 59.910 179.290 60.230 179.550 ;
        RECT 62.670 179.490 62.990 179.550 ;
        RECT 64.065 179.490 64.355 179.535 ;
        RECT 62.670 179.350 64.355 179.490 ;
        RECT 62.670 179.290 62.990 179.350 ;
        RECT 64.065 179.305 64.355 179.350 ;
        RECT 64.530 179.305 64.820 179.535 ;
        RECT 59.080 179.150 59.220 179.290 ;
        RECT 54.480 179.010 59.220 179.150 ;
        RECT 64.600 179.150 64.740 179.305 ;
        RECT 65.890 179.150 66.210 179.210 ;
        RECT 66.440 179.195 66.580 179.690 ;
        RECT 67.260 179.645 67.590 179.690 ;
        RECT 69.120 179.645 69.410 179.875 ;
        RECT 69.550 179.830 69.890 179.875 ;
        RECT 69.550 179.690 70.050 179.830 ;
        RECT 69.550 179.645 69.890 179.690 ;
        RECT 67.270 179.630 67.590 179.645 ;
        RECT 69.570 179.630 69.890 179.645 ;
        RECT 77.390 179.630 77.710 179.890 ;
        RECT 77.850 179.630 78.170 179.890 ;
        RECT 80.165 179.830 80.455 179.875 ;
        RECT 81.070 179.830 81.390 179.890 ;
        RECT 81.620 179.875 81.760 180.030 ;
        RECT 86.145 179.985 86.435 180.030 ;
        RECT 91.665 180.170 91.955 180.215 ;
        RECT 94.410 180.170 94.730 180.230 ;
        RECT 95.790 180.170 96.110 180.230 ;
        RECT 91.665 180.030 96.110 180.170 ;
        RECT 91.665 179.985 91.955 180.030 ;
        RECT 94.410 179.970 94.730 180.030 ;
        RECT 95.790 179.970 96.110 180.030 ;
        RECT 96.250 180.170 96.570 180.230 ;
        RECT 104.990 180.170 105.310 180.230 ;
        RECT 106.460 180.170 106.600 180.710 ;
        RECT 107.380 180.510 107.520 180.710 ;
        RECT 107.750 180.710 112.210 180.850 ;
        RECT 107.750 180.650 108.070 180.710 ;
        RECT 110.970 180.650 111.290 180.710 ;
        RECT 111.890 180.650 112.210 180.710 ;
        RECT 112.825 180.850 113.115 180.895 ;
        RECT 113.270 180.850 113.590 180.910 ;
        RECT 112.825 180.710 113.590 180.850 ;
        RECT 112.825 180.665 113.115 180.710 ;
        RECT 113.270 180.650 113.590 180.710 ;
        RECT 113.730 180.850 114.050 180.910 ;
        RECT 129.370 180.850 129.690 180.910 ;
        RECT 113.730 180.710 129.690 180.850 ;
        RECT 113.730 180.650 114.050 180.710 ;
        RECT 129.370 180.650 129.690 180.710 ;
        RECT 133.050 180.650 133.370 180.910 ;
        RECT 114.190 180.510 114.510 180.570 ;
        RECT 115.570 180.510 115.890 180.570 ;
        RECT 107.380 180.370 115.890 180.510 ;
        RECT 114.190 180.310 114.510 180.370 ;
        RECT 115.570 180.310 115.890 180.370 ;
        RECT 121.090 180.510 121.410 180.570 ;
        RECT 121.090 180.370 134.200 180.510 ;
        RECT 121.090 180.310 121.410 180.370 ;
        RECT 110.065 180.170 110.355 180.215 ;
        RECT 113.270 180.170 113.590 180.230 ;
        RECT 121.550 180.170 121.870 180.230 ;
        RECT 96.250 180.030 105.310 180.170 ;
        RECT 96.250 179.970 96.570 180.030 ;
        RECT 104.990 179.970 105.310 180.030 ;
        RECT 106.000 180.030 106.600 180.170 ;
        RECT 107.380 180.030 108.900 180.170 ;
        RECT 80.165 179.690 81.390 179.830 ;
        RECT 80.165 179.645 80.455 179.690 ;
        RECT 81.070 179.630 81.390 179.690 ;
        RECT 81.545 179.645 81.835 179.875 ;
        RECT 81.990 179.830 82.310 179.890 ;
        RECT 83.385 179.830 83.675 179.875 ;
        RECT 81.990 179.690 83.675 179.830 ;
        RECT 81.990 179.630 82.310 179.690 ;
        RECT 83.385 179.645 83.675 179.690 ;
        RECT 83.845 179.645 84.135 179.875 ;
        RECT 67.730 179.290 68.050 179.550 ;
        RECT 68.190 179.290 68.510 179.550 ;
        RECT 77.940 179.490 78.080 179.630 ;
        RECT 77.480 179.350 78.080 179.490 ;
        RECT 80.610 179.490 80.930 179.550 ;
        RECT 83.920 179.490 84.060 179.645 ;
        RECT 84.750 179.630 85.070 179.890 ;
        RECT 85.670 179.630 85.990 179.890 ;
        RECT 86.605 179.830 86.895 179.875 ;
        RECT 88.445 179.830 88.735 179.875 ;
        RECT 86.605 179.690 88.735 179.830 ;
        RECT 86.605 179.645 86.895 179.690 ;
        RECT 88.445 179.645 88.735 179.690 ;
        RECT 86.680 179.490 86.820 179.645 ;
        RECT 89.350 179.630 89.670 179.890 ;
        RECT 90.270 179.630 90.590 179.890 ;
        RECT 91.190 179.875 91.510 179.890 ;
        RECT 90.975 179.645 91.510 179.875 ;
        RECT 93.045 179.830 93.335 179.875 ;
        RECT 95.330 179.830 95.650 179.890 ;
        RECT 99.025 179.830 99.315 179.875 ;
        RECT 93.045 179.690 93.445 179.830 ;
        RECT 95.330 179.690 99.315 179.830 ;
        RECT 93.045 179.645 93.335 179.690 ;
        RECT 91.190 179.630 91.510 179.645 ;
        RECT 80.610 179.350 86.820 179.490 ;
        RECT 64.600 179.010 66.210 179.150 ;
        RECT 37.370 178.950 37.690 179.010 ;
        RECT 37.845 178.965 38.135 179.010 ;
        RECT 65.890 178.950 66.210 179.010 ;
        RECT 66.365 178.965 66.655 179.195 ;
        RECT 67.820 179.150 67.960 179.290 ;
        RECT 77.480 179.150 77.620 179.350 ;
        RECT 80.610 179.290 80.930 179.350 ;
        RECT 89.810 179.290 90.130 179.550 ;
        RECT 92.585 179.490 92.875 179.535 ;
        RECT 93.120 179.490 93.260 179.645 ;
        RECT 95.330 179.630 95.650 179.690 ;
        RECT 99.025 179.645 99.315 179.690 ;
        RECT 99.485 179.645 99.775 179.875 ;
        RECT 100.850 179.830 101.170 179.890 ;
        RECT 101.325 179.830 101.615 179.875 ;
        RECT 102.230 179.830 102.550 179.890 ;
        RECT 100.850 179.690 102.550 179.830 ;
        RECT 92.585 179.350 97.400 179.490 ;
        RECT 92.585 179.305 92.875 179.350 ;
        RECT 67.820 179.010 77.620 179.150 ;
        RECT 78.310 179.150 78.630 179.210 ;
        RECT 79.245 179.150 79.535 179.195 ;
        RECT 78.310 179.010 79.535 179.150 ;
        RECT 78.310 178.950 78.630 179.010 ;
        RECT 79.245 178.965 79.535 179.010 ;
        RECT 81.990 179.150 82.310 179.210 ;
        RECT 82.465 179.150 82.755 179.195 ;
        RECT 81.990 179.010 82.755 179.150 ;
        RECT 81.990 178.950 82.310 179.010 ;
        RECT 82.465 178.965 82.755 179.010 ;
        RECT 95.760 179.150 96.050 179.195 ;
        RECT 96.710 179.150 97.030 179.210 ;
        RECT 95.760 179.010 97.030 179.150 ;
        RECT 97.260 179.150 97.400 179.350 ;
        RECT 97.630 179.290 97.950 179.550 ;
        RECT 98.550 179.490 98.870 179.550 ;
        RECT 99.560 179.490 99.700 179.645 ;
        RECT 100.850 179.630 101.170 179.690 ;
        RECT 101.325 179.645 101.615 179.690 ;
        RECT 102.230 179.630 102.550 179.690 ;
        RECT 102.690 179.630 103.010 179.890 ;
        RECT 103.610 179.630 103.930 179.890 ;
        RECT 104.070 179.830 104.390 179.890 ;
        RECT 105.450 179.830 105.770 179.890 ;
        RECT 106.000 179.875 106.140 180.030 ;
        RECT 106.770 179.875 107.090 179.890 ;
        RECT 104.070 179.690 105.770 179.830 ;
        RECT 104.070 179.630 104.390 179.690 ;
        RECT 105.450 179.630 105.770 179.690 ;
        RECT 105.925 179.645 106.215 179.875 ;
        RECT 106.770 179.645 107.135 179.875 ;
        RECT 106.770 179.630 107.090 179.645 ;
        RECT 98.550 179.350 99.700 179.490 ;
        RECT 104.530 179.490 104.850 179.550 ;
        RECT 107.380 179.490 107.520 180.030 ;
        RECT 107.750 179.630 108.070 179.890 ;
        RECT 108.760 179.875 108.900 180.030 ;
        RECT 110.065 180.030 113.590 180.170 ;
        RECT 110.065 179.985 110.355 180.030 ;
        RECT 113.270 179.970 113.590 180.030 ;
        RECT 114.510 180.030 121.870 180.170 ;
        RECT 108.685 179.830 108.975 179.875 ;
        RECT 110.510 179.830 110.830 179.890 ;
        RECT 108.685 179.690 110.830 179.830 ;
        RECT 108.685 179.645 108.975 179.690 ;
        RECT 110.510 179.630 110.830 179.690 ;
        RECT 111.430 179.630 111.750 179.890 ;
        RECT 111.890 179.630 112.210 179.890 ;
        RECT 114.510 179.830 114.650 180.030 ;
        RECT 121.550 179.970 121.870 180.030 ;
        RECT 112.860 179.690 114.650 179.830 ;
        RECT 120.630 179.830 120.950 179.890 ;
        RECT 134.060 179.875 134.200 180.370 ;
        RECT 123.405 179.830 123.695 179.875 ;
        RECT 120.630 179.690 123.695 179.830 ;
        RECT 104.530 179.350 107.520 179.490 ;
        RECT 98.550 179.290 98.870 179.350 ;
        RECT 104.530 179.290 104.850 179.350 ;
        RECT 108.225 179.305 108.515 179.535 ;
        RECT 110.985 179.490 111.275 179.535 ;
        RECT 112.860 179.490 113.000 179.690 ;
        RECT 120.630 179.630 120.950 179.690 ;
        RECT 123.405 179.645 123.695 179.690 ;
        RECT 133.985 179.645 134.275 179.875 ;
        RECT 110.985 179.350 113.000 179.490 ;
        RECT 110.985 179.305 111.275 179.350 ;
        RECT 99.470 179.150 99.790 179.210 ;
        RECT 97.260 179.010 99.790 179.150 ;
        RECT 95.760 178.965 96.050 179.010 ;
        RECT 96.710 178.950 97.030 179.010 ;
        RECT 99.470 178.950 99.790 179.010 ;
        RECT 102.245 179.150 102.535 179.195 ;
        RECT 103.610 179.150 103.930 179.210 ;
        RECT 102.245 179.010 103.930 179.150 ;
        RECT 108.300 179.150 108.440 179.305 ;
        RECT 114.650 179.290 114.970 179.550 ;
        RECT 122.930 179.290 123.250 179.550 ;
        RECT 108.670 179.150 108.990 179.210 ;
        RECT 108.300 179.010 108.990 179.150 ;
        RECT 102.245 178.965 102.535 179.010 ;
        RECT 103.610 178.950 103.930 179.010 ;
        RECT 108.670 178.950 108.990 179.010 ;
        RECT 109.605 179.150 109.895 179.195 ;
        RECT 110.510 179.150 110.830 179.210 ;
        RECT 109.605 179.010 110.830 179.150 ;
        RECT 109.605 178.965 109.895 179.010 ;
        RECT 110.510 178.950 110.830 179.010 ;
        RECT 123.390 179.150 123.710 179.210 ;
        RECT 129.845 179.150 130.135 179.195 ;
        RECT 131.210 179.150 131.530 179.210 ;
        RECT 123.390 179.010 131.530 179.150 ;
        RECT 123.390 178.950 123.710 179.010 ;
        RECT 129.845 178.965 130.135 179.010 ;
        RECT 131.210 178.950 131.530 179.010 ;
        RECT 23.500 178.330 136.200 178.810 ;
        RECT 39.685 178.130 39.975 178.175 ;
        RECT 41.970 178.130 42.290 178.190 ;
        RECT 45.665 178.130 45.955 178.175 ;
        RECT 39.685 177.990 42.290 178.130 ;
        RECT 39.685 177.945 39.975 177.990 ;
        RECT 41.970 177.930 42.290 177.990 ;
        RECT 43.900 177.990 45.955 178.130 ;
        RECT 37.845 177.790 38.135 177.835 ;
        RECT 38.290 177.790 38.610 177.850 ;
        RECT 41.050 177.790 41.370 177.850 ;
        RECT 43.900 177.835 44.040 177.990 ;
        RECT 45.665 177.945 45.955 177.990 ;
        RECT 48.870 177.930 49.190 178.190 ;
        RECT 51.630 178.130 51.950 178.190 ;
        RECT 52.105 178.130 52.395 178.175 ;
        RECT 51.630 177.990 52.395 178.130 ;
        RECT 51.630 177.930 51.950 177.990 ;
        RECT 52.105 177.945 52.395 177.990 ;
        RECT 63.145 178.130 63.435 178.175 ;
        RECT 64.050 178.130 64.370 178.190 ;
        RECT 63.145 177.990 64.370 178.130 ;
        RECT 63.145 177.945 63.435 177.990 ;
        RECT 64.050 177.930 64.370 177.990 ;
        RECT 67.270 178.130 67.590 178.190 ;
        RECT 89.810 178.130 90.130 178.190 ;
        RECT 67.270 177.990 90.130 178.130 ;
        RECT 67.270 177.930 67.590 177.990 ;
        RECT 89.810 177.930 90.130 177.990 ;
        RECT 92.585 178.130 92.875 178.175 ;
        RECT 93.950 178.130 94.270 178.190 ;
        RECT 92.585 177.990 94.270 178.130 ;
        RECT 92.585 177.945 92.875 177.990 ;
        RECT 93.950 177.930 94.270 177.990 ;
        RECT 95.790 177.930 96.110 178.190 ;
        RECT 104.990 177.930 105.310 178.190 ;
        RECT 105.925 178.130 106.215 178.175 ;
        RECT 108.210 178.130 108.530 178.190 ;
        RECT 116.490 178.130 116.810 178.190 ;
        RECT 105.925 177.990 116.810 178.130 ;
        RECT 105.925 177.945 106.215 177.990 ;
        RECT 108.210 177.930 108.530 177.990 ;
        RECT 116.490 177.930 116.810 177.990 ;
        RECT 121.550 178.130 121.870 178.190 ;
        RECT 125.690 178.130 126.010 178.190 ;
        RECT 127.545 178.130 127.835 178.175 ;
        RECT 121.550 177.990 125.000 178.130 ;
        RECT 121.550 177.930 121.870 177.990 ;
        RECT 43.825 177.790 44.115 177.835 ;
        RECT 37.845 177.650 38.610 177.790 ;
        RECT 37.845 177.605 38.135 177.650 ;
        RECT 38.290 177.590 38.610 177.650 ;
        RECT 39.300 177.650 44.115 177.790 ;
        RECT 26.330 177.250 26.650 177.510 ;
        RECT 39.300 177.495 39.440 177.650 ;
        RECT 41.050 177.590 41.370 177.650 ;
        RECT 43.825 177.605 44.115 177.650 ;
        RECT 44.270 177.790 44.590 177.850 ;
        RECT 44.745 177.790 45.035 177.835 ;
        RECT 49.330 177.790 49.650 177.850 ;
        RECT 49.805 177.790 50.095 177.835 ;
        RECT 44.270 177.650 46.800 177.790 ;
        RECT 44.270 177.590 44.590 177.650 ;
        RECT 44.745 177.605 45.035 177.650 ;
        RECT 36.005 177.450 36.295 177.495 ;
        RECT 39.225 177.450 39.515 177.495 ;
        RECT 36.005 177.310 39.515 177.450 ;
        RECT 36.005 177.265 36.295 177.310 ;
        RECT 39.225 177.265 39.515 177.310 ;
        RECT 39.670 177.450 39.990 177.510 ;
        RECT 46.660 177.495 46.800 177.650 ;
        RECT 49.330 177.650 50.095 177.790 ;
        RECT 64.140 177.790 64.280 177.930 ;
        RECT 78.770 177.790 79.090 177.850 ;
        RECT 82.910 177.790 83.230 177.850 ;
        RECT 83.385 177.790 83.675 177.835 ;
        RECT 64.140 177.650 82.680 177.790 ;
        RECT 49.330 177.590 49.650 177.650 ;
        RECT 49.805 177.605 50.095 177.650 ;
        RECT 78.770 177.590 79.090 177.650 ;
        RECT 40.145 177.450 40.435 177.495 ;
        RECT 39.670 177.310 40.435 177.450 ;
        RECT 39.670 177.250 39.990 177.310 ;
        RECT 40.145 177.265 40.435 177.310 ;
        RECT 43.365 177.265 43.655 177.495 ;
        RECT 45.205 177.265 45.495 177.495 ;
        RECT 46.585 177.265 46.875 177.495 ;
        RECT 50.250 177.450 50.570 177.510 ;
        RECT 50.725 177.450 51.015 177.495 ;
        RECT 50.250 177.310 51.015 177.450 ;
        RECT 37.370 177.110 37.690 177.170 ;
        RECT 43.440 177.110 43.580 177.265 ;
        RECT 45.280 177.110 45.420 177.265 ;
        RECT 50.250 177.250 50.570 177.310 ;
        RECT 50.725 177.265 51.015 177.310 ;
        RECT 51.170 177.250 51.490 177.510 ;
        RECT 51.630 177.250 51.950 177.510 ;
        RECT 52.565 177.265 52.855 177.495 ;
        RECT 37.370 176.970 45.420 177.110 ;
        RECT 48.410 177.110 48.730 177.170 ;
        RECT 52.640 177.110 52.780 177.265 ;
        RECT 64.510 177.250 64.830 177.510 ;
        RECT 64.970 177.250 65.290 177.510 ;
        RECT 66.825 177.450 67.115 177.495 ;
        RECT 65.980 177.310 67.115 177.450 ;
        RECT 48.410 176.970 52.780 177.110 ;
        RECT 57.610 177.110 57.930 177.170 ;
        RECT 58.990 177.110 59.310 177.170 ;
        RECT 60.845 177.110 61.135 177.155 ;
        RECT 57.610 176.970 61.135 177.110 ;
        RECT 37.370 176.910 37.690 176.970 ;
        RECT 48.410 176.910 48.730 176.970 ;
        RECT 57.610 176.910 57.930 176.970 ;
        RECT 58.990 176.910 59.310 176.970 ;
        RECT 60.845 176.925 61.135 176.970 ;
        RECT 63.590 177.110 63.910 177.170 ;
        RECT 65.980 177.110 66.120 177.310 ;
        RECT 66.825 177.265 67.115 177.310 ;
        RECT 69.570 177.450 69.890 177.510 ;
        RECT 76.470 177.450 76.790 177.510 ;
        RECT 80.165 177.450 80.455 177.495 ;
        RECT 80.610 177.450 80.930 177.510 ;
        RECT 69.570 177.310 76.790 177.450 ;
        RECT 69.570 177.250 69.890 177.310 ;
        RECT 76.470 177.250 76.790 177.310 ;
        RECT 78.400 177.310 80.930 177.450 ;
        RECT 82.540 177.450 82.680 177.650 ;
        RECT 82.910 177.650 83.675 177.790 ;
        RECT 82.910 177.590 83.230 177.650 ;
        RECT 83.385 177.605 83.675 177.650 ;
        RECT 92.125 177.790 92.415 177.835 ;
        RECT 96.250 177.790 96.570 177.850 ;
        RECT 92.125 177.650 96.570 177.790 ;
        RECT 92.125 177.605 92.415 177.650 ;
        RECT 96.250 177.590 96.570 177.650 ;
        RECT 97.645 177.790 97.935 177.835 ;
        RECT 104.070 177.790 104.390 177.850 ;
        RECT 97.645 177.650 104.390 177.790 ;
        RECT 105.080 177.790 105.220 177.930 ;
        RECT 106.385 177.790 106.675 177.835 ;
        RECT 105.080 177.650 106.675 177.790 ;
        RECT 97.645 177.605 97.935 177.650 ;
        RECT 91.650 177.450 91.970 177.510 ;
        RECT 82.540 177.310 91.970 177.450 ;
        RECT 63.590 176.970 66.120 177.110 ;
        RECT 63.590 176.910 63.910 176.970 ;
        RECT 66.350 176.910 66.670 177.170 ;
        RECT 70.490 177.110 70.810 177.170 ;
        RECT 78.400 177.110 78.540 177.310 ;
        RECT 80.165 177.265 80.455 177.310 ;
        RECT 80.610 177.250 80.930 177.310 ;
        RECT 91.650 177.250 91.970 177.310 ;
        RECT 93.490 177.250 93.810 177.510 ;
        RECT 93.965 177.265 94.255 177.495 ;
        RECT 70.490 176.970 78.540 177.110 ;
        RECT 78.770 177.110 79.090 177.170 ;
        RECT 81.545 177.110 81.835 177.155 ;
        RECT 78.770 176.970 81.835 177.110 ;
        RECT 70.490 176.910 70.810 176.970 ;
        RECT 78.770 176.910 79.090 176.970 ;
        RECT 81.545 176.925 81.835 176.970 ;
        RECT 82.450 176.910 82.770 177.170 ;
        RECT 91.740 177.110 91.880 177.250 ;
        RECT 94.040 177.110 94.180 177.265 ;
        RECT 94.410 177.250 94.730 177.510 ;
        RECT 95.345 177.450 95.635 177.495 ;
        RECT 95.790 177.450 96.110 177.510 ;
        RECT 96.725 177.450 97.015 177.495 ;
        RECT 95.345 177.310 97.015 177.450 ;
        RECT 95.345 177.265 95.635 177.310 ;
        RECT 95.790 177.250 96.110 177.310 ;
        RECT 96.725 177.265 97.015 177.310 ;
        RECT 94.870 177.110 95.190 177.170 ;
        RECT 91.740 176.970 95.190 177.110 ;
        RECT 94.870 176.910 95.190 176.970 ;
        RECT 38.765 176.770 39.055 176.815 ;
        RECT 44.270 176.770 44.590 176.830 ;
        RECT 38.765 176.630 44.590 176.770 ;
        RECT 38.765 176.585 39.055 176.630 ;
        RECT 44.270 176.570 44.590 176.630 ;
        RECT 44.730 176.570 45.050 176.830 ;
        RECT 47.030 176.770 47.350 176.830 ;
        RECT 51.630 176.770 51.950 176.830 ;
        RECT 47.030 176.630 51.950 176.770 ;
        RECT 47.030 176.570 47.350 176.630 ;
        RECT 51.630 176.570 51.950 176.630 ;
        RECT 59.910 176.770 60.230 176.830 ;
        RECT 62.210 176.770 62.530 176.830 ;
        RECT 80.625 176.770 80.915 176.815 ;
        RECT 59.910 176.630 62.530 176.770 ;
        RECT 59.910 176.570 60.230 176.630 ;
        RECT 62.210 176.570 62.530 176.630 ;
        RECT 62.760 176.630 80.915 176.770 ;
        RECT 18.970 176.430 19.290 176.490 ;
        RECT 25.425 176.430 25.715 176.475 ;
        RECT 18.970 176.290 25.715 176.430 ;
        RECT 18.970 176.230 19.290 176.290 ;
        RECT 25.425 176.245 25.715 176.290 ;
        RECT 37.830 176.430 38.150 176.490 ;
        RECT 39.670 176.430 39.990 176.490 ;
        RECT 37.830 176.290 39.990 176.430 ;
        RECT 37.830 176.230 38.150 176.290 ;
        RECT 39.670 176.230 39.990 176.290 ;
        RECT 40.130 176.430 40.450 176.490 ;
        RECT 41.970 176.430 42.290 176.490 ;
        RECT 40.130 176.290 42.290 176.430 ;
        RECT 40.130 176.230 40.450 176.290 ;
        RECT 41.970 176.230 42.290 176.290 ;
        RECT 47.505 176.430 47.795 176.475 ;
        RECT 48.410 176.430 48.730 176.490 ;
        RECT 47.505 176.290 48.730 176.430 ;
        RECT 47.505 176.245 47.795 176.290 ;
        RECT 48.410 176.230 48.730 176.290 ;
        RECT 49.805 176.430 50.095 176.475 ;
        RECT 62.760 176.430 62.900 176.630 ;
        RECT 80.625 176.585 80.915 176.630 ;
        RECT 88.430 176.770 88.750 176.830 ;
        RECT 93.490 176.770 93.810 176.830 ;
        RECT 97.720 176.770 97.860 177.605 ;
        RECT 104.070 177.590 104.390 177.650 ;
        RECT 106.385 177.605 106.675 177.650 ;
        RECT 109.130 177.790 109.450 177.850 ;
        RECT 123.390 177.790 123.710 177.850 ;
        RECT 124.325 177.790 124.615 177.835 ;
        RECT 109.130 177.650 121.320 177.790 ;
        RECT 109.130 177.590 109.450 177.650 ;
        RECT 99.025 177.265 99.315 177.495 ;
        RECT 100.405 177.450 100.695 177.495 ;
        RECT 100.850 177.450 101.170 177.510 ;
        RECT 100.405 177.310 101.170 177.450 ;
        RECT 100.405 177.265 100.695 177.310 ;
        RECT 99.100 177.110 99.240 177.265 ;
        RECT 100.850 177.250 101.170 177.310 ;
        RECT 102.245 177.265 102.535 177.495 ;
        RECT 101.770 177.110 102.090 177.170 ;
        RECT 99.100 176.970 102.090 177.110 ;
        RECT 102.320 177.110 102.460 177.265 ;
        RECT 103.150 177.250 103.470 177.510 ;
        RECT 104.530 177.250 104.850 177.510 ;
        RECT 104.990 177.250 105.310 177.510 ;
        RECT 105.450 177.450 105.770 177.510 ;
        RECT 116.490 177.495 116.810 177.510 ;
        RECT 121.180 177.495 121.320 177.650 ;
        RECT 123.390 177.650 124.615 177.790 ;
        RECT 124.860 177.790 125.000 177.990 ;
        RECT 125.690 177.990 127.835 178.130 ;
        RECT 125.690 177.930 126.010 177.990 ;
        RECT 127.545 177.945 127.835 177.990 ;
        RECT 128.925 177.790 129.215 177.835 ;
        RECT 124.860 177.650 129.215 177.790 ;
        RECT 123.390 177.590 123.710 177.650 ;
        RECT 124.325 177.605 124.615 177.650 ;
        RECT 128.925 177.605 129.215 177.650 ;
        RECT 129.370 177.590 129.690 177.850 ;
        RECT 132.130 177.790 132.450 177.850 ;
        RECT 132.130 177.650 133.280 177.790 ;
        RECT 132.130 177.590 132.450 177.650 ;
        RECT 115.585 177.450 115.875 177.495 ;
        RECT 105.450 177.310 115.875 177.450 ;
        RECT 105.450 177.250 105.770 177.310 ;
        RECT 115.585 177.265 115.875 177.310 ;
        RECT 116.475 177.265 116.810 177.495 ;
        RECT 121.105 177.265 121.395 177.495 ;
        RECT 121.550 177.450 121.870 177.510 ;
        RECT 122.025 177.450 122.315 177.495 ;
        RECT 121.550 177.310 122.315 177.450 ;
        RECT 116.490 177.250 116.810 177.265 ;
        RECT 121.550 177.250 121.870 177.310 ;
        RECT 122.025 177.265 122.315 177.310 ;
        RECT 122.470 177.450 122.790 177.510 ;
        RECT 125.230 177.450 125.550 177.510 ;
        RECT 122.470 177.310 125.550 177.450 ;
        RECT 122.470 177.250 122.790 177.310 ;
        RECT 125.230 177.250 125.550 177.310 ;
        RECT 128.450 177.250 128.770 177.510 ;
        RECT 129.830 177.250 130.150 177.510 ;
        RECT 130.765 177.265 131.055 177.495 ;
        RECT 131.210 177.450 131.530 177.510 ;
        RECT 131.685 177.450 131.975 177.495 ;
        RECT 131.210 177.310 131.975 177.450 ;
        RECT 116.045 177.110 116.335 177.155 ;
        RECT 130.840 177.110 130.980 177.265 ;
        RECT 131.210 177.250 131.530 177.310 ;
        RECT 131.685 177.265 131.975 177.310 ;
        RECT 132.590 177.250 132.910 177.510 ;
        RECT 133.140 177.495 133.280 177.650 ;
        RECT 133.065 177.265 133.355 177.495 ;
        RECT 133.985 177.110 134.275 177.155 ;
        RECT 102.320 176.970 105.680 177.110 ;
        RECT 101.770 176.910 102.090 176.970 ;
        RECT 88.430 176.630 93.260 176.770 ;
        RECT 88.430 176.570 88.750 176.630 ;
        RECT 49.805 176.290 62.900 176.430 ;
        RECT 63.130 176.430 63.450 176.490 ;
        RECT 63.605 176.430 63.895 176.475 ;
        RECT 63.130 176.290 63.895 176.430 ;
        RECT 93.120 176.430 93.260 176.630 ;
        RECT 93.490 176.630 97.860 176.770 ;
        RECT 100.390 176.770 100.710 176.830 ;
        RECT 104.530 176.770 104.850 176.830 ;
        RECT 100.390 176.630 104.850 176.770 ;
        RECT 93.490 176.570 93.810 176.630 ;
        RECT 100.390 176.570 100.710 176.630 ;
        RECT 104.530 176.570 104.850 176.630 ;
        RECT 98.105 176.430 98.395 176.475 ;
        RECT 99.010 176.430 99.330 176.490 ;
        RECT 93.120 176.290 99.330 176.430 ;
        RECT 49.805 176.245 50.095 176.290 ;
        RECT 63.130 176.230 63.450 176.290 ;
        RECT 63.605 176.245 63.895 176.290 ;
        RECT 98.105 176.245 98.395 176.290 ;
        RECT 99.010 176.230 99.330 176.290 ;
        RECT 99.930 176.230 100.250 176.490 ;
        RECT 103.150 176.430 103.470 176.490 ;
        RECT 103.625 176.430 103.915 176.475 ;
        RECT 103.150 176.290 103.915 176.430 ;
        RECT 105.540 176.430 105.680 176.970 ;
        RECT 116.045 176.970 129.600 177.110 ;
        RECT 130.840 176.970 134.275 177.110 ;
        RECT 116.045 176.925 116.335 176.970 ;
        RECT 110.970 176.770 111.290 176.830 ;
        RECT 125.230 176.770 125.550 176.830 ;
        RECT 110.970 176.630 125.550 176.770 ;
        RECT 110.970 176.570 111.290 176.630 ;
        RECT 125.230 176.570 125.550 176.630 ;
        RECT 109.130 176.430 109.450 176.490 ;
        RECT 105.540 176.290 109.450 176.430 ;
        RECT 103.150 176.230 103.470 176.290 ;
        RECT 103.625 176.245 103.915 176.290 ;
        RECT 109.130 176.230 109.450 176.290 ;
        RECT 113.745 176.430 114.035 176.475 ;
        RECT 114.190 176.430 114.510 176.490 ;
        RECT 120.170 176.430 120.490 176.490 ;
        RECT 113.745 176.290 120.490 176.430 ;
        RECT 113.745 176.245 114.035 176.290 ;
        RECT 114.190 176.230 114.510 176.290 ;
        RECT 120.170 176.230 120.490 176.290 ;
        RECT 121.550 176.230 121.870 176.490 ;
        RECT 123.405 176.430 123.695 176.475 ;
        RECT 123.850 176.430 124.170 176.490 ;
        RECT 123.405 176.290 124.170 176.430 ;
        RECT 129.460 176.430 129.600 176.970 ;
        RECT 133.985 176.925 134.275 176.970 ;
        RECT 132.145 176.770 132.435 176.815 ;
        RECT 134.430 176.770 134.750 176.830 ;
        RECT 132.145 176.630 134.750 176.770 ;
        RECT 132.145 176.585 132.435 176.630 ;
        RECT 134.430 176.570 134.750 176.630 ;
        RECT 129.830 176.430 130.150 176.490 ;
        RECT 129.460 176.290 130.150 176.430 ;
        RECT 123.405 176.245 123.695 176.290 ;
        RECT 123.850 176.230 124.170 176.290 ;
        RECT 129.830 176.230 130.150 176.290 ;
        RECT 23.500 175.610 136.200 176.090 ;
        RECT 27.710 175.410 28.030 175.470 ;
        RECT 39.210 175.410 39.530 175.470 ;
        RECT 46.570 175.410 46.890 175.470 ;
        RECT 54.850 175.410 55.170 175.470 ;
        RECT 27.710 175.270 32.540 175.410 ;
        RECT 27.710 175.210 28.030 175.270 ;
        RECT 32.400 175.115 32.540 175.270 ;
        RECT 39.210 175.270 55.170 175.410 ;
        RECT 39.210 175.210 39.530 175.270 ;
        RECT 46.570 175.210 46.890 175.270 ;
        RECT 54.850 175.210 55.170 175.270 ;
        RECT 56.690 175.410 57.010 175.470 ;
        RECT 67.270 175.410 67.590 175.470 ;
        RECT 56.690 175.270 67.590 175.410 ;
        RECT 56.690 175.210 57.010 175.270 ;
        RECT 67.270 175.210 67.590 175.270 ;
        RECT 67.730 175.410 68.050 175.470 ;
        RECT 68.205 175.410 68.495 175.455 ;
        RECT 72.805 175.410 73.095 175.455 ;
        RECT 67.730 175.270 73.095 175.410 ;
        RECT 67.730 175.210 68.050 175.270 ;
        RECT 68.205 175.225 68.495 175.270 ;
        RECT 72.805 175.225 73.095 175.270 ;
        RECT 82.925 175.410 83.215 175.455 ;
        RECT 84.750 175.410 85.070 175.470 ;
        RECT 99.470 175.410 99.790 175.470 ;
        RECT 115.570 175.410 115.890 175.470 ;
        RECT 128.450 175.410 128.770 175.470 ;
        RECT 82.925 175.270 85.070 175.410 ;
        RECT 82.925 175.225 83.215 175.270 ;
        RECT 84.750 175.210 85.070 175.270 ;
        RECT 85.300 175.270 99.240 175.410 ;
        RECT 29.105 174.885 29.395 175.115 ;
        RECT 32.325 175.070 32.615 175.115 ;
        RECT 34.610 175.070 34.930 175.130 ;
        RECT 32.325 174.930 34.930 175.070 ;
        RECT 32.325 174.885 32.615 174.930 ;
        RECT 27.710 174.530 28.030 174.790 ;
        RECT 25.870 174.390 26.190 174.450 ;
        RECT 26.345 174.390 26.635 174.435 ;
        RECT 29.180 174.390 29.320 174.885 ;
        RECT 34.610 174.870 34.930 174.930 ;
        RECT 44.270 175.070 44.590 175.130 ;
        RECT 48.410 175.070 48.730 175.130 ;
        RECT 44.270 174.930 48.730 175.070 ;
        RECT 44.270 174.870 44.590 174.930 ;
        RECT 48.410 174.870 48.730 174.930 ;
        RECT 50.250 174.870 50.570 175.130 ;
        RECT 57.610 175.070 57.930 175.130 ;
        RECT 64.065 175.070 64.355 175.115 ;
        RECT 57.610 174.930 64.355 175.070 ;
        RECT 57.610 174.870 57.930 174.930 ;
        RECT 64.065 174.885 64.355 174.930 ;
        RECT 64.985 175.070 65.275 175.115 ;
        RECT 69.570 175.070 69.890 175.130 ;
        RECT 85.300 175.070 85.440 175.270 ;
        RECT 93.490 175.070 93.810 175.130 ;
        RECT 64.985 174.930 69.890 175.070 ;
        RECT 64.985 174.885 65.275 174.930 ;
        RECT 69.570 174.870 69.890 174.930 ;
        RECT 71.040 174.930 85.440 175.070 ;
        RECT 92.660 174.930 93.810 175.070 ;
        RECT 38.750 174.730 39.070 174.790 ;
        RECT 39.350 174.730 39.640 174.775 ;
        RECT 33.780 174.590 39.640 174.730 ;
        RECT 33.780 174.435 33.920 174.590 ;
        RECT 38.750 174.530 39.070 174.590 ;
        RECT 39.350 174.545 39.640 174.590 ;
        RECT 47.505 174.730 47.795 174.775 ;
        RECT 67.745 174.730 68.035 174.775 ;
        RECT 68.190 174.730 68.510 174.790 ;
        RECT 71.040 174.730 71.180 174.930 ;
        RECT 47.505 174.590 66.580 174.730 ;
        RECT 47.505 174.545 47.795 174.590 ;
        RECT 30.945 174.390 31.235 174.435 ;
        RECT 33.705 174.390 33.995 174.435 ;
        RECT 25.870 174.250 33.995 174.390 ;
        RECT 25.870 174.190 26.190 174.250 ;
        RECT 26.345 174.205 26.635 174.250 ;
        RECT 30.945 174.205 31.235 174.250 ;
        RECT 33.705 174.205 33.995 174.250 ;
        RECT 34.610 174.390 34.930 174.450 ;
        RECT 36.925 174.390 37.215 174.435 ;
        RECT 41.510 174.390 41.830 174.450 ;
        RECT 34.610 174.250 37.215 174.390 ;
        RECT 34.610 174.190 34.930 174.250 ;
        RECT 36.925 174.205 37.215 174.250 ;
        RECT 37.460 174.250 41.830 174.390 ;
        RECT 37.460 174.050 37.600 174.250 ;
        RECT 41.510 174.190 41.830 174.250 ;
        RECT 44.270 174.190 44.590 174.450 ;
        RECT 45.205 174.205 45.495 174.435 ;
        RECT 31.710 173.910 37.600 174.050 ;
        RECT 38.305 174.050 38.595 174.095 ;
        RECT 40.590 174.050 40.910 174.110 ;
        RECT 38.305 173.910 40.910 174.050 ;
        RECT 26.805 173.710 27.095 173.755 ;
        RECT 28.630 173.710 28.950 173.770 ;
        RECT 26.805 173.570 28.950 173.710 ;
        RECT 26.805 173.525 27.095 173.570 ;
        RECT 28.630 173.510 28.950 173.570 ;
        RECT 30.025 173.710 30.315 173.755 ;
        RECT 31.710 173.710 31.850 173.910 ;
        RECT 38.305 173.865 38.595 173.910 ;
        RECT 40.590 173.850 40.910 173.910 ;
        RECT 41.050 174.050 41.370 174.110 ;
        RECT 43.810 174.050 44.130 174.110 ;
        RECT 45.280 174.050 45.420 174.205 ;
        RECT 46.570 174.190 46.890 174.450 ;
        RECT 48.870 174.190 49.190 174.450 ;
        RECT 50.265 174.390 50.555 174.435 ;
        RECT 50.710 174.390 51.030 174.450 ;
        RECT 50.265 174.250 51.030 174.390 ;
        RECT 50.265 174.205 50.555 174.250 ;
        RECT 50.710 174.190 51.030 174.250 ;
        RECT 56.705 174.390 56.995 174.435 ;
        RECT 58.070 174.390 58.390 174.450 ;
        RECT 56.705 174.250 58.390 174.390 ;
        RECT 56.705 174.205 56.995 174.250 ;
        RECT 58.070 174.190 58.390 174.250 ;
        RECT 62.210 174.390 62.530 174.450 ;
        RECT 62.685 174.390 62.975 174.435 ;
        RECT 65.890 174.390 66.210 174.450 ;
        RECT 66.440 174.435 66.580 174.590 ;
        RECT 67.745 174.590 71.180 174.730 ;
        RECT 71.410 174.730 71.730 174.790 ;
        RECT 71.885 174.730 72.175 174.775 ;
        RECT 71.410 174.590 72.175 174.730 ;
        RECT 67.745 174.545 68.035 174.590 ;
        RECT 68.190 174.530 68.510 174.590 ;
        RECT 71.410 174.530 71.730 174.590 ;
        RECT 71.885 174.545 72.175 174.590 ;
        RECT 76.010 174.530 76.330 174.790 ;
        RECT 76.560 174.590 78.540 174.730 ;
        RECT 62.210 174.250 66.210 174.390 ;
        RECT 62.210 174.190 62.530 174.250 ;
        RECT 62.685 174.205 62.975 174.250 ;
        RECT 65.890 174.190 66.210 174.250 ;
        RECT 66.365 174.390 66.655 174.435 ;
        RECT 67.270 174.390 67.590 174.450 ;
        RECT 66.365 174.250 67.590 174.390 ;
        RECT 66.365 174.205 66.655 174.250 ;
        RECT 67.270 174.190 67.590 174.250 ;
        RECT 69.585 174.205 69.875 174.435 ;
        RECT 70.965 174.205 71.255 174.435 ;
        RECT 72.345 174.205 72.635 174.435 ;
        RECT 73.265 174.390 73.555 174.435 ;
        RECT 74.170 174.390 74.490 174.450 ;
        RECT 73.265 174.250 74.490 174.390 ;
        RECT 73.265 174.205 73.555 174.250 ;
        RECT 41.050 173.910 45.420 174.050 ;
        RECT 49.345 174.050 49.635 174.095 ;
        RECT 49.790 174.050 50.110 174.110 ;
        RECT 63.130 174.050 63.450 174.110 ;
        RECT 69.660 174.050 69.800 174.205 ;
        RECT 49.345 173.910 57.840 174.050 ;
        RECT 41.050 173.850 41.370 173.910 ;
        RECT 43.810 173.850 44.130 173.910 ;
        RECT 49.345 173.865 49.635 173.910 ;
        RECT 49.790 173.850 50.110 173.910 ;
        RECT 30.025 173.570 31.850 173.710 ;
        RECT 30.025 173.525 30.315 173.570 ;
        RECT 33.230 173.510 33.550 173.770 ;
        RECT 35.530 173.510 35.850 173.770 ;
        RECT 37.830 173.710 38.150 173.770 ;
        RECT 38.765 173.710 39.055 173.755 ;
        RECT 39.670 173.710 39.990 173.770 ;
        RECT 37.830 173.570 39.990 173.710 ;
        RECT 37.830 173.510 38.150 173.570 ;
        RECT 38.765 173.525 39.055 173.570 ;
        RECT 39.670 173.510 39.990 173.570 ;
        RECT 40.145 173.710 40.435 173.755 ;
        RECT 47.030 173.710 47.350 173.770 ;
        RECT 40.145 173.570 47.350 173.710 ;
        RECT 40.145 173.525 40.435 173.570 ;
        RECT 47.030 173.510 47.350 173.570 ;
        RECT 47.950 173.710 48.270 173.770 ;
        RECT 57.150 173.710 57.470 173.770 ;
        RECT 47.950 173.570 57.470 173.710 ;
        RECT 57.700 173.710 57.840 173.910 ;
        RECT 63.130 173.910 69.800 174.050 ;
        RECT 63.130 173.850 63.450 173.910 ;
        RECT 66.810 173.710 67.130 173.770 ;
        RECT 57.700 173.570 67.130 173.710 ;
        RECT 47.950 173.510 48.270 173.570 ;
        RECT 57.150 173.510 57.470 173.570 ;
        RECT 66.810 173.510 67.130 173.570 ;
        RECT 69.125 173.710 69.415 173.755 ;
        RECT 69.570 173.710 69.890 173.770 ;
        RECT 69.125 173.570 69.890 173.710 ;
        RECT 69.125 173.525 69.415 173.570 ;
        RECT 69.570 173.510 69.890 173.570 ;
        RECT 70.045 173.710 70.335 173.755 ;
        RECT 70.490 173.710 70.810 173.770 ;
        RECT 70.045 173.570 70.810 173.710 ;
        RECT 71.040 173.710 71.180 174.205 ;
        RECT 71.410 174.050 71.730 174.110 ;
        RECT 72.420 174.050 72.560 174.205 ;
        RECT 74.170 174.190 74.490 174.250 ;
        RECT 75.550 174.390 75.870 174.450 ;
        RECT 76.560 174.390 76.700 174.590 ;
        RECT 75.550 174.250 76.700 174.390 ;
        RECT 75.550 174.190 75.870 174.250 ;
        RECT 76.945 174.205 77.235 174.435 ;
        RECT 77.405 174.390 77.695 174.435 ;
        RECT 77.850 174.390 78.170 174.450 ;
        RECT 77.405 174.250 78.170 174.390 ;
        RECT 78.400 174.390 78.540 174.590 ;
        RECT 78.770 174.530 79.090 174.790 ;
        RECT 79.230 174.730 79.550 174.790 ;
        RECT 89.810 174.730 90.130 174.790 ;
        RECT 92.660 174.730 92.800 174.930 ;
        RECT 93.490 174.870 93.810 174.930 ;
        RECT 94.870 175.070 95.190 175.130 ;
        RECT 97.170 175.070 97.490 175.130 ;
        RECT 94.870 174.930 97.490 175.070 ;
        RECT 99.100 175.070 99.240 175.270 ;
        RECT 99.470 175.270 114.650 175.410 ;
        RECT 99.470 175.210 99.790 175.270 ;
        RECT 106.370 175.070 106.690 175.130 ;
        RECT 107.750 175.070 108.070 175.130 ;
        RECT 99.100 174.930 108.070 175.070 ;
        RECT 94.870 174.870 95.190 174.930 ;
        RECT 97.170 174.870 97.490 174.930 ;
        RECT 106.370 174.870 106.690 174.930 ;
        RECT 107.750 174.870 108.070 174.930 ;
        RECT 108.210 175.070 108.530 175.130 ;
        RECT 108.210 174.930 109.820 175.070 ;
        RECT 108.210 174.870 108.530 174.930 ;
        RECT 79.230 174.590 84.060 174.730 ;
        RECT 79.230 174.530 79.550 174.590 ;
        RECT 79.690 174.390 80.010 174.450 ;
        RECT 78.400 174.250 80.010 174.390 ;
        RECT 77.405 174.205 77.695 174.250 ;
        RECT 74.630 174.050 74.950 174.110 ;
        RECT 71.410 173.910 74.950 174.050 ;
        RECT 71.410 173.850 71.730 173.910 ;
        RECT 74.630 173.850 74.950 173.910 ;
        RECT 75.640 173.710 75.780 174.190 ;
        RECT 77.020 174.050 77.160 174.205 ;
        RECT 77.850 174.190 78.170 174.250 ;
        RECT 79.690 174.190 80.010 174.250 ;
        RECT 80.150 174.390 80.470 174.450 ;
        RECT 80.625 174.390 80.915 174.435 ;
        RECT 80.150 174.250 80.915 174.390 ;
        RECT 80.150 174.190 80.470 174.250 ;
        RECT 80.625 174.205 80.915 174.250 ;
        RECT 81.070 174.190 81.390 174.450 ;
        RECT 81.550 174.390 81.840 174.435 ;
        RECT 81.990 174.390 82.310 174.450 ;
        RECT 81.550 174.250 82.310 174.390 ;
        RECT 81.550 174.205 81.840 174.250 ;
        RECT 81.990 174.190 82.310 174.250 ;
        RECT 82.450 174.190 82.770 174.450 ;
        RECT 83.920 174.435 84.060 174.590 ;
        RECT 89.810 174.590 92.800 174.730 ;
        RECT 89.810 174.530 90.130 174.590 ;
        RECT 83.845 174.205 84.135 174.435 ;
        RECT 84.305 174.390 84.595 174.435 ;
        RECT 86.130 174.390 86.450 174.450 ;
        RECT 84.305 174.250 86.450 174.390 ;
        RECT 84.305 174.205 84.595 174.250 ;
        RECT 86.130 174.190 86.450 174.250 ;
        RECT 86.590 174.190 86.910 174.450 ;
        RECT 88.430 174.390 88.750 174.450 ;
        RECT 89.365 174.390 89.655 174.435 ;
        RECT 88.430 174.250 89.655 174.390 ;
        RECT 88.430 174.190 88.750 174.250 ;
        RECT 89.365 174.205 89.655 174.250 ;
        RECT 90.285 174.205 90.575 174.435 ;
        RECT 81.160 174.050 81.300 174.190 ;
        RECT 77.020 173.910 81.300 174.050 ;
        RECT 82.925 173.865 83.215 174.095 ;
        RECT 85.210 174.050 85.530 174.110 ;
        RECT 90.360 174.050 90.500 174.205 ;
        RECT 91.650 174.190 91.970 174.450 ;
        RECT 92.660 174.435 92.800 174.590 ;
        RECT 97.630 174.730 97.950 174.790 ;
        RECT 104.990 174.730 105.310 174.790 ;
        RECT 108.670 174.730 108.990 174.790 ;
        RECT 97.630 174.590 104.300 174.730 ;
        RECT 97.630 174.530 97.950 174.590 ;
        RECT 92.585 174.205 92.875 174.435 ;
        RECT 93.505 174.390 93.795 174.435 ;
        RECT 94.410 174.390 94.730 174.450 ;
        RECT 93.505 174.250 94.730 174.390 ;
        RECT 93.505 174.205 93.795 174.250 ;
        RECT 94.410 174.190 94.730 174.250 ;
        RECT 100.850 174.390 101.170 174.450 ;
        RECT 104.160 174.435 104.300 174.590 ;
        RECT 104.990 174.590 108.990 174.730 ;
        RECT 104.990 174.530 105.310 174.590 ;
        RECT 108.670 174.530 108.990 174.590 ;
        RECT 109.130 174.530 109.450 174.790 ;
        RECT 109.680 174.775 109.820 174.930 ;
        RECT 112.810 174.870 113.130 175.130 ;
        RECT 114.510 175.070 114.650 175.270 ;
        RECT 115.570 175.270 128.770 175.410 ;
        RECT 115.570 175.210 115.890 175.270 ;
        RECT 128.450 175.210 128.770 175.270 ;
        RECT 139.950 175.070 140.270 175.130 ;
        RECT 114.510 174.930 140.270 175.070 ;
        RECT 139.950 174.870 140.270 174.930 ;
        RECT 109.605 174.545 109.895 174.775 ;
        RECT 110.050 174.530 110.370 174.790 ;
        RECT 111.445 174.730 111.735 174.775 ;
        RECT 115.110 174.730 115.430 174.790 ;
        RECT 111.445 174.590 115.430 174.730 ;
        RECT 111.445 174.545 111.735 174.590 ;
        RECT 115.110 174.530 115.430 174.590 ;
        RECT 123.045 174.590 133.280 174.730 ;
        RECT 103.165 174.390 103.455 174.435 ;
        RECT 100.850 174.250 103.455 174.390 ;
        RECT 100.850 174.190 101.170 174.250 ;
        RECT 103.165 174.205 103.455 174.250 ;
        RECT 104.085 174.205 104.375 174.435 ;
        RECT 104.530 174.390 104.850 174.450 ;
        RECT 106.830 174.390 107.150 174.450 ;
        RECT 104.530 174.250 107.150 174.390 ;
        RECT 104.530 174.190 104.850 174.250 ;
        RECT 106.830 174.190 107.150 174.250 ;
        RECT 108.210 174.190 108.530 174.450 ;
        RECT 108.760 174.390 108.900 174.530 ;
        RECT 110.525 174.390 110.815 174.435 ;
        RECT 108.760 174.250 110.815 174.390 ;
        RECT 110.525 174.205 110.815 174.250 ;
        RECT 111.890 174.390 112.210 174.450 ;
        RECT 112.365 174.390 112.655 174.435 ;
        RECT 111.890 174.250 112.655 174.390 ;
        RECT 111.890 174.190 112.210 174.250 ;
        RECT 112.365 174.205 112.655 174.250 ;
        RECT 113.270 174.190 113.590 174.450 ;
        RECT 113.730 174.390 114.050 174.450 ;
        RECT 123.045 174.390 123.185 174.590 ;
        RECT 113.730 174.250 123.185 174.390 ;
        RECT 113.730 174.190 114.050 174.250 ;
        RECT 123.390 174.190 123.710 174.450 ;
        RECT 133.140 174.435 133.280 174.590 ;
        RECT 133.065 174.205 133.355 174.435 ;
        RECT 85.210 173.910 90.500 174.050 ;
        RECT 91.190 174.050 91.510 174.110 ;
        RECT 92.125 174.050 92.415 174.095 ;
        RECT 91.190 173.910 92.415 174.050 ;
        RECT 71.040 173.570 75.780 173.710 ;
        RECT 78.325 173.710 78.615 173.755 ;
        RECT 79.230 173.710 79.550 173.770 ;
        RECT 78.325 173.570 79.550 173.710 ;
        RECT 83.000 173.710 83.140 173.865 ;
        RECT 85.210 173.850 85.530 173.910 ;
        RECT 91.190 173.850 91.510 173.910 ;
        RECT 92.125 173.865 92.415 173.910 ;
        RECT 93.030 174.050 93.350 174.110 ;
        RECT 100.390 174.050 100.710 174.110 ;
        RECT 93.030 173.910 100.710 174.050 ;
        RECT 84.750 173.710 85.070 173.770 ;
        RECT 83.000 173.570 85.070 173.710 ;
        RECT 70.045 173.525 70.335 173.570 ;
        RECT 70.490 173.510 70.810 173.570 ;
        RECT 78.325 173.525 78.615 173.570 ;
        RECT 79.230 173.510 79.550 173.570 ;
        RECT 84.750 173.510 85.070 173.570 ;
        RECT 86.145 173.710 86.435 173.755 ;
        RECT 86.590 173.710 86.910 173.770 ;
        RECT 86.145 173.570 86.910 173.710 ;
        RECT 86.145 173.525 86.435 173.570 ;
        RECT 86.590 173.510 86.910 173.570 ;
        RECT 87.510 173.510 87.830 173.770 ;
        RECT 89.810 173.510 90.130 173.770 ;
        RECT 90.730 173.510 91.050 173.770 ;
        RECT 92.200 173.710 92.340 173.865 ;
        RECT 93.030 173.850 93.350 173.910 ;
        RECT 100.390 173.850 100.710 173.910 ;
        RECT 102.690 173.850 103.010 174.110 ;
        RECT 103.240 173.910 113.960 174.050 ;
        RECT 94.410 173.710 94.730 173.770 ;
        RECT 95.790 173.710 96.110 173.770 ;
        RECT 92.200 173.570 96.110 173.710 ;
        RECT 94.410 173.510 94.730 173.570 ;
        RECT 95.790 173.510 96.110 173.570 ;
        RECT 96.250 173.510 96.570 173.770 ;
        RECT 99.010 173.710 99.330 173.770 ;
        RECT 101.310 173.710 101.630 173.770 ;
        RECT 99.010 173.570 101.630 173.710 ;
        RECT 99.010 173.510 99.330 173.570 ;
        RECT 101.310 173.510 101.630 173.570 ;
        RECT 102.230 173.710 102.550 173.770 ;
        RECT 103.240 173.710 103.380 173.910 ;
        RECT 102.230 173.570 103.380 173.710 ;
        RECT 103.625 173.710 103.915 173.755 ;
        RECT 105.450 173.710 105.770 173.770 ;
        RECT 103.625 173.570 105.770 173.710 ;
        RECT 102.230 173.510 102.550 173.570 ;
        RECT 103.625 173.525 103.915 173.570 ;
        RECT 105.450 173.510 105.770 173.570 ;
        RECT 107.290 173.710 107.610 173.770 ;
        RECT 113.270 173.710 113.590 173.770 ;
        RECT 107.290 173.570 113.590 173.710 ;
        RECT 113.820 173.710 113.960 173.910 ;
        RECT 114.190 173.850 114.510 174.110 ;
        RECT 123.850 174.050 124.170 174.110 ;
        RECT 128.910 174.050 129.230 174.110 ;
        RECT 130.750 174.050 131.070 174.110 ;
        RECT 131.225 174.050 131.515 174.095 ;
        RECT 123.850 173.910 127.760 174.050 ;
        RECT 123.850 173.850 124.170 173.910 ;
        RECT 120.645 173.710 120.935 173.755 ;
        RECT 113.820 173.570 120.935 173.710 ;
        RECT 107.290 173.510 107.610 173.570 ;
        RECT 113.270 173.510 113.590 173.570 ;
        RECT 120.645 173.525 120.935 173.570 ;
        RECT 121.550 173.710 121.870 173.770 ;
        RECT 127.070 173.710 127.390 173.770 ;
        RECT 121.550 173.570 127.390 173.710 ;
        RECT 127.620 173.710 127.760 173.910 ;
        RECT 128.910 173.910 131.515 174.050 ;
        RECT 128.910 173.850 129.230 173.910 ;
        RECT 130.750 173.850 131.070 173.910 ;
        RECT 131.225 173.865 131.515 173.910 ;
        RECT 133.985 173.710 134.275 173.755 ;
        RECT 127.620 173.570 134.275 173.710 ;
        RECT 121.550 173.510 121.870 173.570 ;
        RECT 127.070 173.510 127.390 173.570 ;
        RECT 133.985 173.525 134.275 173.570 ;
        RECT 23.500 172.890 136.200 173.370 ;
        RECT 25.870 172.490 26.190 172.750 ;
        RECT 26.330 172.690 26.650 172.750 ;
        RECT 27.725 172.690 28.015 172.735 ;
        RECT 26.330 172.550 28.015 172.690 ;
        RECT 26.330 172.490 26.650 172.550 ;
        RECT 27.725 172.505 28.015 172.550 ;
        RECT 38.290 172.490 38.610 172.750 ;
        RECT 41.510 172.690 41.830 172.750 ;
        RECT 54.390 172.690 54.710 172.750 ;
        RECT 41.510 172.550 54.710 172.690 ;
        RECT 41.510 172.490 41.830 172.550 ;
        RECT 54.390 172.490 54.710 172.550 ;
        RECT 61.290 172.690 61.610 172.750 ;
        RECT 65.905 172.690 66.195 172.735 ;
        RECT 61.290 172.550 66.195 172.690 ;
        RECT 61.290 172.490 61.610 172.550 ;
        RECT 65.905 172.505 66.195 172.550 ;
        RECT 66.825 172.690 67.115 172.735 ;
        RECT 70.030 172.690 70.350 172.750 ;
        RECT 66.825 172.550 70.350 172.690 ;
        RECT 66.825 172.505 67.115 172.550 ;
        RECT 70.030 172.490 70.350 172.550 ;
        RECT 70.950 172.490 71.270 172.750 ;
        RECT 82.450 172.690 82.770 172.750 ;
        RECT 78.400 172.550 82.770 172.690 ;
        RECT 40.605 172.350 40.895 172.395 ;
        RECT 35.160 172.210 40.895 172.350 ;
        RECT 21.730 172.010 22.050 172.070 ;
        RECT 25.425 172.010 25.715 172.055 ;
        RECT 21.730 171.870 25.715 172.010 ;
        RECT 21.730 171.810 22.050 171.870 ;
        RECT 25.425 171.825 25.715 171.870 ;
        RECT 28.630 171.810 28.950 172.070 ;
        RECT 34.610 172.010 34.930 172.070 ;
        RECT 35.160 172.055 35.300 172.210 ;
        RECT 40.605 172.165 40.895 172.210 ;
        RECT 50.250 172.350 50.570 172.410 ;
        RECT 50.250 172.210 77.620 172.350 ;
        RECT 50.250 172.150 50.570 172.210 ;
        RECT 35.085 172.010 35.375 172.055 ;
        RECT 34.610 171.870 35.375 172.010 ;
        RECT 34.610 171.810 34.930 171.870 ;
        RECT 35.085 171.825 35.375 171.870 ;
        RECT 37.830 171.810 38.150 172.070 ;
        RECT 38.765 172.010 39.055 172.055 ;
        RECT 39.210 172.010 39.530 172.070 ;
        RECT 38.765 171.870 39.530 172.010 ;
        RECT 38.765 171.825 39.055 171.870 ;
        RECT 39.210 171.810 39.530 171.870 ;
        RECT 39.670 172.010 39.990 172.070 ;
        RECT 42.430 172.010 42.750 172.070 ;
        RECT 39.670 171.870 42.750 172.010 ;
        RECT 39.670 171.810 39.990 171.870 ;
        RECT 42.430 171.810 42.750 171.870 ;
        RECT 43.365 171.825 43.655 172.055 ;
        RECT 43.825 172.010 44.115 172.055 ;
        RECT 46.110 172.010 46.430 172.070 ;
        RECT 43.825 171.870 46.430 172.010 ;
        RECT 43.825 171.825 44.115 171.870 ;
        RECT 36.005 171.670 36.295 171.715 ;
        RECT 38.290 171.670 38.610 171.730 ;
        RECT 43.440 171.670 43.580 171.825 ;
        RECT 46.110 171.810 46.430 171.870 ;
        RECT 59.450 172.010 59.770 172.070 ;
        RECT 63.605 172.010 63.895 172.055 ;
        RECT 65.430 172.010 65.750 172.070 ;
        RECT 59.450 171.870 65.750 172.010 ;
        RECT 59.450 171.810 59.770 171.870 ;
        RECT 63.605 171.825 63.895 171.870 ;
        RECT 65.430 171.810 65.750 171.870 ;
        RECT 66.135 172.010 66.425 172.055 ;
        RECT 66.810 172.010 67.130 172.070 ;
        RECT 66.135 171.870 67.130 172.010 ;
        RECT 66.135 171.825 66.425 171.870 ;
        RECT 66.810 171.810 67.130 171.870 ;
        RECT 67.270 172.010 67.590 172.070 ;
        RECT 67.745 172.010 68.035 172.055 ;
        RECT 67.270 171.870 68.035 172.010 ;
        RECT 67.270 171.810 67.590 171.870 ;
        RECT 67.745 171.825 68.035 171.870 ;
        RECT 68.190 172.010 68.510 172.070 ;
        RECT 69.125 172.010 69.415 172.055 ;
        RECT 68.190 171.870 69.415 172.010 ;
        RECT 68.190 171.810 68.510 171.870 ;
        RECT 69.125 171.825 69.415 171.870 ;
        RECT 69.570 172.010 69.890 172.070 ;
        RECT 72.805 172.010 73.095 172.055 ;
        RECT 69.570 171.870 73.095 172.010 ;
        RECT 69.570 171.810 69.890 171.870 ;
        RECT 72.805 171.825 73.095 171.870 ;
        RECT 76.470 171.810 76.790 172.070 ;
        RECT 76.930 171.810 77.250 172.070 ;
        RECT 46.570 171.670 46.890 171.730 ;
        RECT 68.650 171.670 68.970 171.730 ;
        RECT 36.005 171.530 38.610 171.670 ;
        RECT 36.005 171.485 36.295 171.530 ;
        RECT 38.290 171.470 38.610 171.530 ;
        RECT 38.840 171.530 68.970 171.670 ;
        RECT 35.530 171.330 35.850 171.390 ;
        RECT 38.840 171.330 38.980 171.530 ;
        RECT 46.570 171.470 46.890 171.530 ;
        RECT 68.650 171.470 68.970 171.530 ;
        RECT 71.870 171.470 72.190 171.730 ;
        RECT 72.345 171.485 72.635 171.715 ;
        RECT 73.250 171.670 73.570 171.730 ;
        RECT 74.630 171.670 74.950 171.730 ;
        RECT 73.250 171.530 74.950 171.670 ;
        RECT 77.480 171.670 77.620 172.210 ;
        RECT 77.850 171.810 78.170 172.070 ;
        RECT 78.400 172.055 78.540 172.550 ;
        RECT 82.450 172.490 82.770 172.550 ;
        RECT 86.130 172.490 86.450 172.750 ;
        RECT 90.745 172.505 91.035 172.735 ;
        RECT 91.280 172.550 94.180 172.690 ;
        RECT 81.530 172.150 81.850 172.410 ;
        RECT 90.820 172.350 90.960 172.505 ;
        RECT 87.140 172.210 90.960 172.350 ;
        RECT 78.325 171.825 78.615 172.055 ;
        RECT 79.230 171.810 79.550 172.070 ;
        RECT 79.705 171.825 79.995 172.055 ;
        RECT 80.170 172.010 80.460 172.055 ;
        RECT 80.610 172.010 80.930 172.070 ;
        RECT 80.170 171.870 80.930 172.010 ;
        RECT 80.170 171.825 80.460 171.870 ;
        RECT 79.780 171.670 79.920 171.825 ;
        RECT 80.610 171.810 80.930 171.870 ;
        RECT 82.925 172.010 83.215 172.055 ;
        RECT 86.605 172.010 86.895 172.055 ;
        RECT 82.925 171.870 86.895 172.010 ;
        RECT 82.925 171.825 83.215 171.870 ;
        RECT 86.605 171.825 86.895 171.870 ;
        RECT 83.000 171.670 83.140 171.825 ;
        RECT 77.480 171.530 79.920 171.670 ;
        RECT 80.700 171.530 83.140 171.670 ;
        RECT 35.530 171.190 38.980 171.330 ;
        RECT 39.685 171.330 39.975 171.375 ;
        RECT 41.050 171.330 41.370 171.390 ;
        RECT 39.685 171.190 41.370 171.330 ;
        RECT 35.530 171.130 35.850 171.190 ;
        RECT 39.685 171.145 39.975 171.190 ;
        RECT 41.050 171.130 41.370 171.190 ;
        RECT 42.430 171.130 42.750 171.390 ;
        RECT 42.890 171.330 43.210 171.390 ;
        RECT 45.190 171.330 45.510 171.390 ;
        RECT 42.890 171.190 45.510 171.330 ;
        RECT 42.890 171.130 43.210 171.190 ;
        RECT 45.190 171.130 45.510 171.190 ;
        RECT 57.150 171.330 57.470 171.390 ;
        RECT 68.190 171.330 68.510 171.390 ;
        RECT 71.410 171.330 71.730 171.390 ;
        RECT 57.150 171.190 68.510 171.330 ;
        RECT 57.150 171.130 57.470 171.190 ;
        RECT 68.190 171.130 68.510 171.190 ;
        RECT 69.660 171.190 71.730 171.330 ;
        RECT 40.590 170.990 40.910 171.050 ;
        RECT 41.510 170.990 41.830 171.050 ;
        RECT 40.590 170.850 41.830 170.990 ;
        RECT 40.590 170.790 40.910 170.850 ;
        RECT 41.510 170.790 41.830 170.850 ;
        RECT 44.745 170.990 45.035 171.035 ;
        RECT 45.650 170.990 45.970 171.050 ;
        RECT 44.745 170.850 45.970 170.990 ;
        RECT 44.745 170.805 45.035 170.850 ;
        RECT 45.650 170.790 45.970 170.850 ;
        RECT 64.065 170.990 64.355 171.035 ;
        RECT 65.890 170.990 66.210 171.050 ;
        RECT 69.660 171.035 69.800 171.190 ;
        RECT 71.410 171.130 71.730 171.190 ;
        RECT 64.065 170.850 66.210 170.990 ;
        RECT 64.065 170.805 64.355 170.850 ;
        RECT 65.890 170.790 66.210 170.850 ;
        RECT 69.585 170.805 69.875 171.035 ;
        RECT 70.490 170.790 70.810 171.050 ;
        RECT 70.950 170.990 71.270 171.050 ;
        RECT 72.420 170.990 72.560 171.485 ;
        RECT 73.250 171.470 73.570 171.530 ;
        RECT 74.630 171.470 74.950 171.530 ;
        RECT 77.865 171.330 78.155 171.375 ;
        RECT 80.150 171.330 80.470 171.390 ;
        RECT 77.865 171.190 80.470 171.330 ;
        RECT 77.865 171.145 78.155 171.190 ;
        RECT 80.150 171.130 80.470 171.190 ;
        RECT 70.950 170.850 72.560 170.990 ;
        RECT 77.390 170.990 77.710 171.050 ;
        RECT 80.700 170.990 80.840 171.530 ;
        RECT 84.765 171.485 85.055 171.715 ;
        RECT 85.225 171.670 85.515 171.715 ;
        RECT 86.130 171.670 86.450 171.730 ;
        RECT 85.225 171.530 86.450 171.670 ;
        RECT 85.225 171.485 85.515 171.530 ;
        RECT 81.990 171.330 82.310 171.390 ;
        RECT 84.840 171.330 84.980 171.485 ;
        RECT 86.130 171.470 86.450 171.530 ;
        RECT 87.140 171.330 87.280 172.210 ;
        RECT 90.745 172.010 91.035 172.055 ;
        RECT 91.280 172.010 91.420 172.550 ;
        RECT 94.040 172.410 94.180 172.550 ;
        RECT 94.870 172.490 95.190 172.750 ;
        RECT 99.470 172.690 99.790 172.750 ;
        RECT 99.470 172.550 131.440 172.690 ;
        RECT 99.470 172.490 99.790 172.550 ;
        RECT 93.045 172.350 93.335 172.395 ;
        RECT 92.200 172.210 93.335 172.350 ;
        RECT 90.745 171.870 91.420 172.010 ;
        RECT 91.630 172.010 91.920 172.055 ;
        RECT 92.200 172.010 92.340 172.210 ;
        RECT 93.045 172.165 93.335 172.210 ;
        RECT 93.950 172.350 94.270 172.410 ;
        RECT 94.425 172.350 94.715 172.395 ;
        RECT 93.950 172.210 94.715 172.350 ;
        RECT 94.960 172.350 95.100 172.490 ;
        RECT 99.930 172.350 100.250 172.410 ;
        RECT 117.870 172.350 118.190 172.410 ;
        RECT 118.345 172.350 118.635 172.395 ;
        RECT 94.960 172.210 98.320 172.350 ;
        RECT 93.950 172.150 94.270 172.210 ;
        RECT 94.425 172.165 94.715 172.210 ;
        RECT 91.630 171.870 92.340 172.010 ;
        RECT 90.745 171.825 91.035 171.870 ;
        RECT 91.630 171.825 91.970 171.870 ;
        RECT 92.560 171.825 92.850 172.055 ;
        RECT 88.430 171.470 88.750 171.730 ;
        RECT 88.905 171.670 89.195 171.715 ;
        RECT 88.905 171.530 90.960 171.670 ;
        RECT 91.650 171.640 91.970 171.825 ;
        RECT 92.635 171.670 92.775 171.825 ;
        RECT 93.490 171.810 93.810 172.070 ;
        RECT 95.345 172.010 95.635 172.055 ;
        RECT 94.500 171.870 95.635 172.010 ;
        RECT 94.500 171.730 94.640 171.870 ;
        RECT 95.345 171.825 95.635 171.870 ;
        RECT 96.250 172.010 96.570 172.070 ;
        RECT 98.180 172.055 98.320 172.210 ;
        RECT 99.930 172.210 116.720 172.350 ;
        RECT 99.930 172.150 100.250 172.210 ;
        RECT 96.250 171.870 97.860 172.010 ;
        RECT 96.250 171.810 96.570 171.870 ;
        RECT 93.950 171.670 94.270 171.730 ;
        RECT 92.635 171.530 94.270 171.670 ;
        RECT 88.905 171.485 89.195 171.530 ;
        RECT 81.990 171.190 87.280 171.330 ;
        RECT 90.820 171.330 90.960 171.530 ;
        RECT 93.950 171.470 94.270 171.530 ;
        RECT 94.410 171.470 94.730 171.730 ;
        RECT 96.725 171.485 97.015 171.715 ;
        RECT 97.185 171.485 97.475 171.715 ;
        RECT 97.720 171.670 97.860 171.870 ;
        RECT 98.105 171.825 98.395 172.055 ;
        RECT 99.010 172.010 99.330 172.070 ;
        RECT 99.485 172.010 99.775 172.055 ;
        RECT 100.405 172.010 100.695 172.055 ;
        RECT 99.010 171.870 99.775 172.010 ;
        RECT 99.010 171.810 99.330 171.870 ;
        RECT 99.485 171.825 99.775 171.870 ;
        RECT 100.020 171.870 100.695 172.010 ;
        RECT 100.020 171.670 100.160 171.870 ;
        RECT 100.405 171.825 100.695 171.870 ;
        RECT 102.230 171.810 102.550 172.070 ;
        RECT 102.705 171.825 102.995 172.055 ;
        RECT 103.150 172.010 103.470 172.070 ;
        RECT 106.370 172.010 106.690 172.070 ;
        RECT 103.150 171.870 106.690 172.010 ;
        RECT 97.720 171.530 100.160 171.670 ;
        RECT 101.770 171.670 102.090 171.730 ;
        RECT 102.780 171.670 102.920 171.825 ;
        RECT 103.150 171.810 103.470 171.870 ;
        RECT 106.370 171.810 106.690 171.870 ;
        RECT 109.130 172.010 109.450 172.070 ;
        RECT 114.665 172.010 114.955 172.055 ;
        RECT 116.030 172.010 116.350 172.070 ;
        RECT 109.130 171.870 114.420 172.010 ;
        RECT 109.130 171.810 109.450 171.870 ;
        RECT 101.770 171.530 102.920 171.670 ;
        RECT 93.490 171.330 93.810 171.390 ;
        RECT 95.790 171.330 96.110 171.390 ;
        RECT 90.820 171.190 91.190 171.330 ;
        RECT 81.990 171.130 82.310 171.190 ;
        RECT 77.390 170.850 80.840 170.990 ;
        RECT 84.290 170.990 84.610 171.050 ;
        RECT 89.825 170.990 90.115 171.035 ;
        RECT 84.290 170.850 90.115 170.990 ;
        RECT 91.050 170.990 91.190 171.190 ;
        RECT 93.490 171.190 96.110 171.330 ;
        RECT 93.490 171.130 93.810 171.190 ;
        RECT 95.790 171.130 96.110 171.190 ;
        RECT 94.425 170.990 94.715 171.035 ;
        RECT 91.050 170.850 94.715 170.990 ;
        RECT 96.800 170.990 96.940 171.485 ;
        RECT 97.260 171.330 97.400 171.485 ;
        RECT 101.770 171.470 102.090 171.530 ;
        RECT 104.085 171.485 104.375 171.715 ;
        RECT 105.005 171.670 105.295 171.715 ;
        RECT 113.730 171.670 114.050 171.730 ;
        RECT 105.005 171.530 114.050 171.670 ;
        RECT 114.280 171.670 114.420 171.870 ;
        RECT 114.665 171.870 116.350 172.010 ;
        RECT 116.580 172.010 116.720 172.210 ;
        RECT 117.870 172.210 118.635 172.350 ;
        RECT 117.870 172.150 118.190 172.210 ;
        RECT 118.345 172.165 118.635 172.210 ;
        RECT 118.790 172.350 119.110 172.410 ;
        RECT 121.105 172.350 121.395 172.395 ;
        RECT 118.790 172.210 125.460 172.350 ;
        RECT 118.790 172.150 119.110 172.210 ;
        RECT 121.105 172.165 121.395 172.210 ;
        RECT 120.185 172.010 120.475 172.055 ;
        RECT 116.580 171.870 120.475 172.010 ;
        RECT 114.665 171.825 114.955 171.870 ;
        RECT 116.030 171.810 116.350 171.870 ;
        RECT 120.185 171.825 120.475 171.870 ;
        RECT 121.565 171.825 121.855 172.055 ;
        RECT 122.930 172.010 123.250 172.070 ;
        RECT 123.405 172.010 123.695 172.055 ;
        RECT 122.930 171.870 123.695 172.010 ;
        RECT 121.640 171.670 121.780 171.825 ;
        RECT 122.930 171.810 123.250 171.870 ;
        RECT 123.405 171.825 123.695 171.870 ;
        RECT 124.770 171.810 125.090 172.070 ;
        RECT 125.320 172.010 125.460 172.210 ;
        RECT 127.070 172.150 127.390 172.410 ;
        RECT 127.530 172.150 127.850 172.410 ;
        RECT 125.320 171.870 128.450 172.010 ;
        RECT 125.690 171.670 126.010 171.730 ;
        RECT 114.280 171.530 126.010 171.670 ;
        RECT 105.005 171.485 105.295 171.530 ;
        RECT 98.090 171.330 98.410 171.390 ;
        RECT 97.260 171.190 98.410 171.330 ;
        RECT 104.160 171.330 104.300 171.485 ;
        RECT 113.730 171.470 114.050 171.530 ;
        RECT 125.690 171.470 126.010 171.530 ;
        RECT 126.150 171.670 126.470 171.730 ;
        RECT 127.530 171.670 127.850 171.730 ;
        RECT 126.150 171.530 127.850 171.670 ;
        RECT 128.310 171.670 128.450 171.870 ;
        RECT 128.910 171.810 129.230 172.070 ;
        RECT 131.300 172.055 131.440 172.550 ;
        RECT 131.225 171.825 131.515 172.055 ;
        RECT 131.670 171.810 131.990 172.070 ;
        RECT 132.605 171.825 132.895 172.055 ;
        RECT 129.485 171.670 129.775 171.715 ;
        RECT 128.310 171.530 129.775 171.670 ;
        RECT 126.150 171.470 126.470 171.530 ;
        RECT 127.530 171.470 127.850 171.530 ;
        RECT 129.485 171.485 129.775 171.530 ;
        RECT 131.210 171.330 131.530 171.390 ;
        RECT 132.680 171.330 132.820 171.825 ;
        RECT 133.050 171.810 133.370 172.070 ;
        RECT 104.160 171.190 132.820 171.330 ;
        RECT 98.090 171.130 98.410 171.190 ;
        RECT 131.210 171.130 131.530 171.190 ;
        RECT 97.170 170.990 97.490 171.050 ;
        RECT 96.800 170.850 97.490 170.990 ;
        RECT 70.950 170.790 71.270 170.850 ;
        RECT 77.390 170.790 77.710 170.850 ;
        RECT 84.290 170.790 84.610 170.850 ;
        RECT 89.825 170.805 90.115 170.850 ;
        RECT 94.425 170.805 94.715 170.850 ;
        RECT 97.170 170.790 97.490 170.850 ;
        RECT 98.550 170.990 98.870 171.050 ;
        RECT 99.025 170.990 99.315 171.035 ;
        RECT 98.550 170.850 99.315 170.990 ;
        RECT 98.550 170.790 98.870 170.850 ;
        RECT 99.025 170.805 99.315 170.850 ;
        RECT 100.405 170.990 100.695 171.035 ;
        RECT 105.910 170.990 106.230 171.050 ;
        RECT 100.405 170.850 106.230 170.990 ;
        RECT 100.405 170.805 100.695 170.850 ;
        RECT 105.910 170.790 106.230 170.850 ;
        RECT 108.210 170.790 108.530 171.050 ;
        RECT 111.890 170.990 112.210 171.050 ;
        RECT 126.150 170.990 126.470 171.050 ;
        RECT 111.890 170.850 126.470 170.990 ;
        RECT 111.890 170.790 112.210 170.850 ;
        RECT 126.150 170.790 126.470 170.850 ;
        RECT 128.450 170.990 128.770 171.050 ;
        RECT 130.305 170.990 130.595 171.035 ;
        RECT 128.450 170.850 130.595 170.990 ;
        RECT 128.450 170.790 128.770 170.850 ;
        RECT 130.305 170.805 130.595 170.850 ;
        RECT 133.970 170.790 134.290 171.050 ;
        RECT 23.500 170.170 136.200 170.650 ;
        RECT 44.745 169.970 45.035 170.015 ;
        RECT 46.110 169.970 46.430 170.030 ;
        RECT 44.745 169.830 46.430 169.970 ;
        RECT 44.745 169.785 45.035 169.830 ;
        RECT 46.110 169.770 46.430 169.830 ;
        RECT 58.085 169.970 58.375 170.015 ;
        RECT 59.450 169.970 59.770 170.030 ;
        RECT 58.085 169.830 59.770 169.970 ;
        RECT 58.085 169.785 58.375 169.830 ;
        RECT 59.450 169.770 59.770 169.830 ;
        RECT 59.925 169.970 60.215 170.015 ;
        RECT 63.130 169.970 63.450 170.030 ;
        RECT 59.925 169.830 63.450 169.970 ;
        RECT 59.925 169.785 60.215 169.830 ;
        RECT 63.130 169.770 63.450 169.830 ;
        RECT 65.890 169.770 66.210 170.030 ;
        RECT 69.570 169.970 69.890 170.030 ;
        RECT 67.335 169.830 69.890 169.970 ;
        RECT 27.725 169.445 28.015 169.675 ;
        RECT 37.830 169.630 38.150 169.690 ;
        RECT 41.970 169.630 42.290 169.690 ;
        RECT 42.905 169.630 43.195 169.675 ;
        RECT 45.190 169.630 45.510 169.690 ;
        RECT 67.335 169.630 67.475 169.830 ;
        RECT 69.570 169.770 69.890 169.830 ;
        RECT 71.870 169.970 72.190 170.030 ;
        RECT 77.850 169.970 78.170 170.030 ;
        RECT 79.705 169.970 79.995 170.015 ;
        RECT 71.870 169.830 74.860 169.970 ;
        RECT 71.870 169.770 72.190 169.830 ;
        RECT 37.830 169.490 38.980 169.630 ;
        RECT 26.345 168.950 26.635 168.995 ;
        RECT 27.800 168.950 27.940 169.445 ;
        RECT 37.830 169.430 38.150 169.490 ;
        RECT 38.840 169.335 38.980 169.490 ;
        RECT 41.970 169.490 67.475 169.630 ;
        RECT 68.650 169.630 68.970 169.690 ;
        RECT 70.045 169.630 70.335 169.675 ;
        RECT 68.650 169.490 73.020 169.630 ;
        RECT 41.970 169.430 42.290 169.490 ;
        RECT 42.905 169.445 43.195 169.490 ;
        RECT 45.190 169.430 45.510 169.490 ;
        RECT 68.650 169.430 68.970 169.490 ;
        RECT 70.045 169.445 70.335 169.490 ;
        RECT 38.765 169.290 39.055 169.335 ;
        RECT 43.365 169.290 43.655 169.335 ;
        RECT 46.110 169.290 46.430 169.350 ;
        RECT 62.210 169.290 62.530 169.350 ;
        RECT 38.765 169.150 43.120 169.290 ;
        RECT 38.765 169.105 39.055 169.150 ;
        RECT 42.980 169.010 43.120 169.150 ;
        RECT 43.365 169.150 46.430 169.290 ;
        RECT 43.365 169.105 43.655 169.150 ;
        RECT 46.110 169.090 46.430 169.150 ;
        RECT 56.320 169.150 62.530 169.290 ;
        RECT 56.320 169.010 56.460 169.150 ;
        RECT 62.210 169.090 62.530 169.150 ;
        RECT 66.350 169.290 66.670 169.350 ;
        RECT 70.505 169.290 70.795 169.335 ;
        RECT 72.330 169.290 72.650 169.350 ;
        RECT 66.350 169.150 70.795 169.290 ;
        RECT 66.350 169.090 66.670 169.150 ;
        RECT 70.505 169.105 70.795 169.150 ;
        RECT 71.500 169.150 72.650 169.290 ;
        RECT 26.345 168.810 27.940 168.950 ;
        RECT 28.645 168.950 28.935 168.995 ;
        RECT 37.830 168.950 38.150 169.010 ;
        RECT 28.645 168.810 38.150 168.950 ;
        RECT 26.345 168.765 26.635 168.810 ;
        RECT 28.645 168.765 28.935 168.810 ;
        RECT 37.830 168.750 38.150 168.810 ;
        RECT 39.685 168.950 39.975 168.995 ;
        RECT 41.050 168.950 41.370 169.010 ;
        RECT 39.685 168.810 41.370 168.950 ;
        RECT 39.685 168.765 39.975 168.810 ;
        RECT 41.050 168.750 41.370 168.810 ;
        RECT 41.985 168.765 42.275 168.995 ;
        RECT 38.750 168.610 39.070 168.670 ;
        RECT 42.060 168.610 42.200 168.765 ;
        RECT 42.890 168.750 43.210 169.010 ;
        RECT 43.825 168.950 44.115 168.995 ;
        RECT 44.270 168.950 44.590 169.010 ;
        RECT 43.825 168.810 44.590 168.950 ;
        RECT 43.825 168.765 44.115 168.810 ;
        RECT 44.270 168.750 44.590 168.810 ;
        RECT 45.650 168.750 45.970 169.010 ;
        RECT 46.585 168.950 46.875 168.995 ;
        RECT 47.030 168.950 47.350 169.010 ;
        RECT 46.585 168.810 47.350 168.950 ;
        RECT 46.585 168.765 46.875 168.810 ;
        RECT 47.030 168.750 47.350 168.810 ;
        RECT 56.230 168.750 56.550 169.010 ;
        RECT 57.610 168.750 57.930 169.010 ;
        RECT 59.450 168.750 59.770 169.010 ;
        RECT 60.385 168.950 60.675 168.995 ;
        RECT 66.810 168.950 67.130 169.010 ;
        RECT 60.385 168.810 67.130 168.950 ;
        RECT 60.385 168.765 60.675 168.810 ;
        RECT 66.810 168.750 67.130 168.810 ;
        RECT 67.270 168.750 67.590 169.010 ;
        RECT 67.745 168.765 68.035 168.995 ;
        RECT 58.070 168.610 58.390 168.670 ;
        RECT 67.820 168.610 67.960 168.765 ;
        RECT 68.190 168.750 68.510 169.010 ;
        RECT 69.125 168.765 69.415 168.995 ;
        RECT 69.585 168.950 69.875 168.995 ;
        RECT 70.030 168.950 70.350 169.010 ;
        RECT 71.500 168.995 71.640 169.150 ;
        RECT 72.330 169.090 72.650 169.150 ;
        RECT 69.585 168.810 70.350 168.950 ;
        RECT 69.585 168.765 69.875 168.810 ;
        RECT 68.650 168.610 68.970 168.670 ;
        RECT 38.750 168.470 57.840 168.610 ;
        RECT 38.750 168.410 39.070 168.470 ;
        RECT 21.730 168.270 22.050 168.330 ;
        RECT 25.425 168.270 25.715 168.315 ;
        RECT 21.730 168.130 25.715 168.270 ;
        RECT 21.730 168.070 22.050 168.130 ;
        RECT 25.425 168.085 25.715 168.130 ;
        RECT 40.130 168.270 40.450 168.330 ;
        RECT 40.605 168.270 40.895 168.315 ;
        RECT 40.130 168.130 40.895 168.270 ;
        RECT 40.130 168.070 40.450 168.130 ;
        RECT 40.605 168.085 40.895 168.130 ;
        RECT 41.050 168.070 41.370 168.330 ;
        RECT 47.505 168.270 47.795 168.315 ;
        RECT 51.630 168.270 51.950 168.330 ;
        RECT 47.505 168.130 51.950 168.270 ;
        RECT 57.700 168.270 57.840 168.470 ;
        RECT 58.070 168.470 67.500 168.610 ;
        RECT 67.820 168.470 68.970 168.610 ;
        RECT 69.200 168.610 69.340 168.765 ;
        RECT 70.030 168.750 70.350 168.810 ;
        RECT 71.425 168.765 71.715 168.995 ;
        RECT 71.870 168.750 72.190 169.010 ;
        RECT 72.880 168.995 73.020 169.490 ;
        RECT 74.720 169.335 74.860 169.830 ;
        RECT 77.850 169.830 79.995 169.970 ;
        RECT 77.850 169.770 78.170 169.830 ;
        RECT 79.705 169.785 79.995 169.830 ;
        RECT 85.210 169.970 85.530 170.030 ;
        RECT 85.685 169.970 85.975 170.015 ;
        RECT 85.210 169.830 85.975 169.970 ;
        RECT 85.210 169.770 85.530 169.830 ;
        RECT 85.685 169.785 85.975 169.830 ;
        RECT 86.590 169.970 86.910 170.030 ;
        RECT 87.525 169.970 87.815 170.015 ;
        RECT 90.745 169.970 91.035 170.015 ;
        RECT 93.950 169.970 94.270 170.030 ;
        RECT 94.425 169.970 94.715 170.015 ;
        RECT 86.590 169.830 87.815 169.970 ;
        RECT 76.010 169.630 76.330 169.690 ;
        RECT 83.385 169.630 83.675 169.675 ;
        RECT 76.010 169.490 83.675 169.630 ;
        RECT 76.010 169.430 76.330 169.490 ;
        RECT 83.385 169.445 83.675 169.490 ;
        RECT 74.645 169.290 74.935 169.335 ;
        RECT 78.770 169.290 79.090 169.350 ;
        RECT 84.290 169.290 84.610 169.350 ;
        RECT 74.645 169.150 79.090 169.290 ;
        RECT 74.645 169.105 74.935 169.150 ;
        RECT 78.770 169.090 79.090 169.150 ;
        RECT 81.160 169.150 84.610 169.290 ;
        RECT 81.160 168.995 81.300 169.150 ;
        RECT 84.290 169.090 84.610 169.150 ;
        RECT 72.805 168.765 73.095 168.995 ;
        RECT 80.625 168.950 80.915 168.995 ;
        RECT 73.340 168.810 80.915 168.950 ;
        RECT 70.490 168.610 70.810 168.670 ;
        RECT 73.340 168.610 73.480 168.810 ;
        RECT 80.625 168.765 80.915 168.810 ;
        RECT 81.085 168.765 81.375 168.995 ;
        RECT 81.990 168.750 82.310 169.010 ;
        RECT 83.385 168.950 83.675 168.995 ;
        RECT 83.830 168.950 84.150 169.010 ;
        RECT 83.385 168.810 84.150 168.950 ;
        RECT 83.385 168.765 83.675 168.810 ;
        RECT 83.830 168.750 84.150 168.810 ;
        RECT 85.760 168.670 85.900 169.785 ;
        RECT 86.590 169.770 86.910 169.830 ;
        RECT 87.525 169.785 87.815 169.830 ;
        RECT 89.470 169.830 91.035 169.970 ;
        RECT 86.130 169.630 86.450 169.690 ;
        RECT 89.470 169.630 89.610 169.830 ;
        RECT 90.745 169.785 91.035 169.830 ;
        RECT 92.200 169.830 94.715 169.970 ;
        RECT 86.130 169.490 89.610 169.630 ;
        RECT 86.130 169.430 86.450 169.490 ;
        RECT 91.190 169.430 91.510 169.690 ;
        RECT 92.200 169.290 92.340 169.830 ;
        RECT 93.950 169.770 94.270 169.830 ;
        RECT 94.425 169.785 94.715 169.830 ;
        RECT 99.930 169.770 100.250 170.030 ;
        RECT 102.230 169.970 102.550 170.030 ;
        RECT 104.990 169.970 105.310 170.030 ;
        RECT 102.230 169.830 105.310 169.970 ;
        RECT 102.230 169.770 102.550 169.830 ;
        RECT 104.990 169.770 105.310 169.830 ;
        RECT 109.590 169.970 109.910 170.030 ;
        RECT 112.825 169.970 113.115 170.015 ;
        RECT 115.570 169.970 115.890 170.030 ;
        RECT 109.590 169.830 111.200 169.970 ;
        RECT 109.590 169.770 109.910 169.830 ;
        RECT 94.870 169.630 95.190 169.690 ;
        RECT 100.390 169.630 100.710 169.690 ;
        RECT 101.770 169.630 102.090 169.690 ;
        RECT 109.130 169.630 109.450 169.690 ;
        RECT 110.525 169.630 110.815 169.675 ;
        RECT 94.870 169.490 95.560 169.630 ;
        RECT 94.870 169.430 95.190 169.490 ;
        RECT 95.420 169.335 95.560 169.490 ;
        RECT 100.390 169.490 106.600 169.630 ;
        RECT 100.390 169.430 100.710 169.490 ;
        RECT 101.770 169.430 102.090 169.490 ;
        RECT 89.435 169.150 92.340 169.290 ;
        RECT 89.435 169.050 89.575 169.150 ;
        RECT 95.345 169.105 95.635 169.335 ;
        RECT 97.170 169.290 97.490 169.350 ;
        RECT 105.005 169.290 105.295 169.335 ;
        RECT 97.170 169.150 105.295 169.290 ;
        RECT 97.170 169.090 97.490 169.150 ;
        RECT 105.005 169.105 105.295 169.150 ;
        RECT 88.980 169.045 89.575 169.050 ;
        RECT 86.145 168.765 86.435 168.995 ;
        RECT 86.605 168.950 86.895 168.995 ;
        RECT 87.970 168.950 88.290 169.010 ;
        RECT 86.605 168.810 88.290 168.950 ;
        RECT 88.880 168.910 89.575 169.045 ;
        RECT 88.880 168.815 89.170 168.910 ;
        RECT 86.605 168.765 86.895 168.810 ;
        RECT 69.200 168.470 73.480 168.610 ;
        RECT 73.725 168.610 74.015 168.655 ;
        RECT 74.170 168.610 74.490 168.670 ;
        RECT 73.725 168.470 74.490 168.610 ;
        RECT 58.070 168.410 58.390 168.470 ;
        RECT 66.350 168.270 66.670 168.330 ;
        RECT 57.700 168.130 66.670 168.270 ;
        RECT 67.360 168.270 67.500 168.470 ;
        RECT 68.650 168.410 68.970 168.470 ;
        RECT 70.490 168.410 70.810 168.470 ;
        RECT 73.725 168.425 74.015 168.470 ;
        RECT 74.170 168.410 74.490 168.470 ;
        RECT 74.630 168.610 74.950 168.670 ;
        RECT 79.705 168.610 79.995 168.655 ;
        RECT 80.150 168.610 80.470 168.670 ;
        RECT 82.465 168.610 82.755 168.655 ;
        RECT 74.630 168.470 80.470 168.610 ;
        RECT 74.630 168.410 74.950 168.470 ;
        RECT 79.705 168.425 79.995 168.470 ;
        RECT 80.150 168.410 80.470 168.470 ;
        RECT 80.700 168.470 82.755 168.610 ;
        RECT 70.965 168.270 71.255 168.315 ;
        RECT 73.250 168.270 73.570 168.330 ;
        RECT 67.360 168.130 73.570 168.270 ;
        RECT 47.505 168.085 47.795 168.130 ;
        RECT 51.630 168.070 51.950 168.130 ;
        RECT 66.350 168.070 66.670 168.130 ;
        RECT 70.965 168.085 71.255 168.130 ;
        RECT 73.250 168.070 73.570 168.130 ;
        RECT 76.930 168.270 77.250 168.330 ;
        RECT 80.700 168.270 80.840 168.470 ;
        RECT 82.465 168.425 82.755 168.470 ;
        RECT 82.910 168.610 83.230 168.670 ;
        RECT 85.225 168.610 85.515 168.655 ;
        RECT 82.910 168.470 85.515 168.610 ;
        RECT 82.910 168.410 83.230 168.470 ;
        RECT 85.225 168.425 85.515 168.470 ;
        RECT 85.670 168.410 85.990 168.670 ;
        RECT 86.220 168.610 86.360 168.765 ;
        RECT 87.970 168.750 88.290 168.810 ;
        RECT 89.825 168.765 90.115 168.995 ;
        RECT 87.510 168.610 87.830 168.670 ;
        RECT 86.220 168.470 87.830 168.610 ;
        RECT 87.510 168.410 87.830 168.470 ;
        RECT 89.365 168.425 89.655 168.655 ;
        RECT 89.900 168.610 90.040 168.765 ;
        RECT 90.730 168.750 91.050 169.010 ;
        RECT 92.110 168.750 92.430 169.010 ;
        RECT 92.570 168.750 92.890 169.010 ;
        RECT 93.030 168.750 93.350 169.010 ;
        RECT 93.965 168.950 94.255 168.995 ;
        RECT 94.410 168.950 94.730 169.010 ;
        RECT 95.805 168.950 96.095 168.995 ;
        RECT 93.965 168.810 94.730 168.950 ;
        RECT 93.965 168.765 94.255 168.810 ;
        RECT 94.410 168.750 94.730 168.810 ;
        RECT 94.960 168.810 96.095 168.950 ;
        RECT 94.960 168.670 95.100 168.810 ;
        RECT 95.805 168.765 96.095 168.810 ;
        RECT 97.630 168.750 97.950 169.010 ;
        RECT 98.550 168.750 98.870 169.010 ;
        RECT 99.010 168.750 99.330 169.010 ;
        RECT 99.560 168.810 101.540 168.950 ;
        RECT 93.490 168.610 93.810 168.670 ;
        RECT 89.900 168.470 93.810 168.610 ;
        RECT 76.930 168.130 80.840 168.270 ;
        RECT 84.305 168.270 84.595 168.315 ;
        RECT 84.750 168.270 85.070 168.330 ;
        RECT 84.305 168.130 85.070 168.270 ;
        RECT 89.435 168.270 89.575 168.425 ;
        RECT 93.490 168.410 93.810 168.470 ;
        RECT 94.870 168.410 95.190 168.670 ;
        RECT 97.185 168.425 97.475 168.655 ;
        RECT 97.720 168.610 97.860 168.750 ;
        RECT 99.560 168.610 99.700 168.810 ;
        RECT 97.720 168.470 99.700 168.610 ;
        RECT 99.945 168.425 100.235 168.655 ;
        RECT 101.400 168.610 101.540 168.810 ;
        RECT 101.770 168.750 102.090 169.010 ;
        RECT 102.230 168.750 102.550 169.010 ;
        RECT 102.705 168.765 102.995 168.995 ;
        RECT 102.780 168.610 102.920 168.765 ;
        RECT 103.610 168.750 103.930 169.010 ;
        RECT 105.910 168.750 106.230 169.010 ;
        RECT 106.460 168.950 106.600 169.490 ;
        RECT 109.130 169.490 110.815 169.630 ;
        RECT 111.060 169.630 111.200 169.830 ;
        RECT 112.825 169.830 115.890 169.970 ;
        RECT 112.825 169.785 113.115 169.830 ;
        RECT 115.570 169.770 115.890 169.830 ;
        RECT 120.630 169.770 120.950 170.030 ;
        RECT 124.785 169.630 125.075 169.675 ;
        RECT 111.060 169.490 125.075 169.630 ;
        RECT 109.130 169.430 109.450 169.490 ;
        RECT 110.525 169.445 110.815 169.490 ;
        RECT 124.785 169.445 125.075 169.490 ;
        RECT 126.150 169.630 126.470 169.690 ;
        RECT 133.970 169.630 134.290 169.690 ;
        RECT 126.150 169.490 134.290 169.630 ;
        RECT 126.150 169.430 126.470 169.490 ;
        RECT 133.970 169.430 134.290 169.490 ;
        RECT 107.305 169.290 107.595 169.335 ;
        RECT 110.085 169.290 110.375 169.335 ;
        RECT 107.305 169.150 110.375 169.290 ;
        RECT 107.305 169.105 107.595 169.150 ;
        RECT 110.085 169.105 110.375 169.150 ;
        RECT 112.810 169.290 113.130 169.350 ;
        RECT 121.090 169.290 121.410 169.350 ;
        RECT 112.810 169.150 121.410 169.290 ;
        RECT 112.810 169.090 113.130 169.150 ;
        RECT 121.090 169.090 121.410 169.150 ;
        RECT 125.320 169.150 128.450 169.290 ;
        RECT 125.320 169.010 125.460 169.150 ;
        RECT 107.750 168.950 108.070 169.010 ;
        RECT 108.225 168.950 108.515 168.995 ;
        RECT 106.460 168.810 108.515 168.950 ;
        RECT 107.750 168.750 108.070 168.810 ;
        RECT 108.225 168.765 108.515 168.810 ;
        RECT 108.685 168.765 108.975 168.995 ;
        RECT 101.400 168.470 102.920 168.610 ;
        RECT 104.070 168.610 104.390 168.670 ;
        RECT 108.760 168.610 108.900 168.765 ;
        RECT 112.350 168.750 112.670 169.010 ;
        RECT 125.230 168.750 125.550 169.010 ;
        RECT 125.690 168.750 126.010 169.010 ;
        RECT 128.310 168.950 128.450 169.150 ;
        RECT 133.525 168.950 133.815 168.995 ;
        RECT 128.310 168.810 133.815 168.950 ;
        RECT 133.525 168.765 133.815 168.810 ;
        RECT 104.070 168.470 108.900 168.610 ;
        RECT 109.130 168.610 109.450 168.670 ;
        RECT 114.205 168.610 114.495 168.655 ;
        RECT 109.130 168.470 114.495 168.610 ;
        RECT 89.810 168.270 90.130 168.330 ;
        RECT 89.435 168.130 90.130 168.270 ;
        RECT 97.260 168.270 97.400 168.425 ;
        RECT 98.550 168.270 98.870 168.330 ;
        RECT 97.260 168.130 98.870 168.270 ;
        RECT 100.020 168.270 100.160 168.425 ;
        RECT 104.070 168.410 104.390 168.470 ;
        RECT 109.130 168.410 109.450 168.470 ;
        RECT 114.205 168.425 114.495 168.470 ;
        RECT 100.405 168.270 100.695 168.315 ;
        RECT 100.020 168.130 100.695 168.270 ;
        RECT 76.930 168.070 77.250 168.130 ;
        RECT 84.305 168.085 84.595 168.130 ;
        RECT 84.750 168.070 85.070 168.130 ;
        RECT 89.810 168.070 90.130 168.130 ;
        RECT 98.550 168.070 98.870 168.130 ;
        RECT 100.405 168.085 100.695 168.130 ;
        RECT 23.500 167.450 136.200 167.930 ;
        RECT 37.830 167.050 38.150 167.310 ;
        RECT 42.905 167.250 43.195 167.295 ;
        RECT 48.870 167.250 49.190 167.310 ;
        RECT 38.380 167.110 42.660 167.250 ;
        RECT 20.810 166.570 21.130 166.630 ;
        RECT 25.425 166.570 25.715 166.615 ;
        RECT 20.810 166.430 25.715 166.570 ;
        RECT 20.810 166.370 21.130 166.430 ;
        RECT 25.425 166.385 25.715 166.430 ;
        RECT 37.370 166.570 37.690 166.630 ;
        RECT 38.380 166.570 38.520 167.110 ;
        RECT 39.685 166.910 39.975 166.955 ;
        RECT 42.520 166.910 42.660 167.110 ;
        RECT 42.905 167.110 49.190 167.250 ;
        RECT 42.905 167.065 43.195 167.110 ;
        RECT 48.870 167.050 49.190 167.110 ;
        RECT 50.710 167.250 51.030 167.310 ;
        RECT 53.010 167.250 53.330 167.310 ;
        RECT 50.710 167.110 51.400 167.250 ;
        RECT 50.710 167.050 51.030 167.110 ;
        RECT 51.260 166.955 51.400 167.110 ;
        RECT 51.720 167.110 53.330 167.250 ;
        RECT 51.720 166.955 51.860 167.110 ;
        RECT 53.010 167.050 53.330 167.110 ;
        RECT 53.470 167.250 53.790 167.310 ;
        RECT 55.310 167.250 55.630 167.310 ;
        RECT 57.165 167.250 57.455 167.295 ;
        RECT 58.070 167.250 58.390 167.310 ;
        RECT 53.470 167.110 55.080 167.250 ;
        RECT 53.470 167.050 53.790 167.110 ;
        RECT 52.090 166.955 52.410 166.970 ;
        RECT 39.685 166.770 42.200 166.910 ;
        RECT 42.520 166.770 50.480 166.910 ;
        RECT 39.685 166.725 39.975 166.770 ;
        RECT 37.370 166.430 38.520 166.570 ;
        RECT 37.370 166.370 37.690 166.430 ;
        RECT 38.750 166.370 39.070 166.630 ;
        RECT 40.130 166.370 40.450 166.630 ;
        RECT 40.605 166.570 40.895 166.615 ;
        RECT 41.050 166.570 41.370 166.630 ;
        RECT 42.060 166.615 42.200 166.770 ;
        RECT 40.605 166.430 41.370 166.570 ;
        RECT 40.605 166.385 40.895 166.430 ;
        RECT 41.050 166.370 41.370 166.430 ;
        RECT 41.525 166.385 41.815 166.615 ;
        RECT 41.985 166.385 42.275 166.615 ;
        RECT 44.285 166.570 44.575 166.615 ;
        RECT 44.730 166.570 45.050 166.630 ;
        RECT 45.280 166.615 45.420 166.770 ;
        RECT 50.340 166.630 50.480 166.770 ;
        RECT 51.185 166.725 51.475 166.955 ;
        RECT 51.645 166.725 51.935 166.955 ;
        RECT 52.090 166.725 52.525 166.955 ;
        RECT 54.940 166.910 55.080 167.110 ;
        RECT 55.310 167.110 58.390 167.250 ;
        RECT 55.310 167.050 55.630 167.110 ;
        RECT 57.165 167.065 57.455 167.110 ;
        RECT 58.070 167.050 58.390 167.110 ;
        RECT 60.385 167.250 60.675 167.295 ;
        RECT 60.830 167.250 61.150 167.310 ;
        RECT 60.385 167.110 61.150 167.250 ;
        RECT 60.385 167.065 60.675 167.110 ;
        RECT 60.830 167.050 61.150 167.110 ;
        RECT 73.710 167.250 74.030 167.310 ;
        RECT 74.185 167.250 74.475 167.295 ;
        RECT 73.710 167.110 74.475 167.250 ;
        RECT 73.710 167.050 74.030 167.110 ;
        RECT 74.185 167.065 74.475 167.110 ;
        RECT 85.210 167.250 85.530 167.310 ;
        RECT 94.410 167.250 94.730 167.310 ;
        RECT 85.210 167.110 94.730 167.250 ;
        RECT 85.210 167.050 85.530 167.110 ;
        RECT 74.630 166.910 74.950 166.970 ;
        RECT 54.940 166.770 74.950 166.910 ;
        RECT 52.090 166.710 52.410 166.725 ;
        RECT 74.630 166.710 74.950 166.770 ;
        RECT 76.010 166.910 76.330 166.970 ;
        RECT 80.150 166.910 80.470 166.970 ;
        RECT 81.545 166.910 81.835 166.955 ;
        RECT 88.430 166.910 88.750 166.970 ;
        RECT 93.120 166.955 93.260 167.110 ;
        RECT 94.410 167.050 94.730 167.110 ;
        RECT 95.790 167.250 96.110 167.310 ;
        RECT 96.265 167.250 96.555 167.295 ;
        RECT 95.790 167.110 96.555 167.250 ;
        RECT 95.790 167.050 96.110 167.110 ;
        RECT 96.265 167.065 96.555 167.110 ;
        RECT 96.710 167.250 97.030 167.310 ;
        RECT 99.930 167.250 100.250 167.310 ;
        RECT 102.705 167.250 102.995 167.295 ;
        RECT 107.305 167.250 107.595 167.295 ;
        RECT 123.390 167.250 123.710 167.310 ;
        RECT 96.710 167.110 102.995 167.250 ;
        RECT 96.710 167.050 97.030 167.110 ;
        RECT 99.930 167.050 100.250 167.110 ;
        RECT 102.705 167.065 102.995 167.110 ;
        RECT 103.240 167.110 107.060 167.250 ;
        RECT 76.010 166.770 77.160 166.910 ;
        RECT 76.010 166.710 76.330 166.770 ;
        RECT 44.285 166.430 45.050 166.570 ;
        RECT 44.285 166.385 44.575 166.430 ;
        RECT 26.345 165.890 26.635 165.935 ;
        RECT 41.600 165.890 41.740 166.385 ;
        RECT 44.730 166.370 45.050 166.430 ;
        RECT 45.205 166.385 45.495 166.615 ;
        RECT 45.650 166.370 45.970 166.630 ;
        RECT 46.110 166.370 46.430 166.630 ;
        RECT 46.570 166.570 46.890 166.630 ;
        RECT 47.045 166.570 47.335 166.615 ;
        RECT 46.570 166.430 47.335 166.570 ;
        RECT 46.570 166.370 46.890 166.430 ;
        RECT 47.045 166.385 47.335 166.430 ;
        RECT 50.250 166.560 50.570 166.630 ;
        RECT 50.725 166.560 51.015 166.615 ;
        RECT 50.250 166.420 51.015 166.560 ;
        RECT 47.120 166.230 47.260 166.385 ;
        RECT 50.250 166.370 50.570 166.420 ;
        RECT 50.725 166.385 51.015 166.420 ;
        RECT 53.010 166.370 53.330 166.630 ;
        RECT 54.390 166.370 54.710 166.630 ;
        RECT 54.850 166.370 55.170 166.630 ;
        RECT 55.310 166.370 55.630 166.630 ;
        RECT 56.245 166.570 56.535 166.615 ;
        RECT 57.150 166.570 57.470 166.630 ;
        RECT 58.990 166.570 59.310 166.630 ;
        RECT 59.465 166.570 59.755 166.615 ;
        RECT 56.245 166.430 58.760 166.570 ;
        RECT 56.245 166.385 56.535 166.430 ;
        RECT 57.150 166.370 57.470 166.430 ;
        RECT 48.870 166.230 49.190 166.290 ;
        RECT 58.620 166.230 58.760 166.430 ;
        RECT 58.990 166.430 59.755 166.570 ;
        RECT 58.990 166.370 59.310 166.430 ;
        RECT 59.465 166.385 59.755 166.430 ;
        RECT 59.910 166.370 60.230 166.630 ;
        RECT 60.370 166.570 60.690 166.630 ;
        RECT 60.845 166.570 61.135 166.615 ;
        RECT 62.670 166.570 62.990 166.630 ;
        RECT 60.370 166.430 62.990 166.570 ;
        RECT 60.370 166.370 60.690 166.430 ;
        RECT 60.845 166.385 61.135 166.430 ;
        RECT 62.670 166.370 62.990 166.430 ;
        RECT 73.725 166.570 74.015 166.615 ;
        RECT 75.090 166.570 75.410 166.630 ;
        RECT 73.725 166.430 75.410 166.570 ;
        RECT 73.725 166.385 74.015 166.430 ;
        RECT 75.090 166.370 75.410 166.430 ;
        RECT 75.550 166.370 75.870 166.630 ;
        RECT 76.485 166.385 76.775 166.615 ;
        RECT 77.020 166.570 77.160 166.770 ;
        RECT 80.150 166.770 81.835 166.910 ;
        RECT 80.150 166.710 80.470 166.770 ;
        RECT 81.545 166.725 81.835 166.770 ;
        RECT 83.000 166.770 88.750 166.910 ;
        RECT 77.405 166.570 77.695 166.615 ;
        RECT 77.020 166.430 77.695 166.570 ;
        RECT 77.405 166.385 77.695 166.430 ;
        RECT 71.870 166.230 72.190 166.290 ;
        RECT 47.120 166.090 49.190 166.230 ;
        RECT 48.870 166.030 49.190 166.090 ;
        RECT 56.170 166.090 58.300 166.230 ;
        RECT 58.620 166.090 72.190 166.230 ;
        RECT 41.970 165.890 42.290 165.950 ;
        RECT 50.710 165.890 51.030 165.950 ;
        RECT 56.170 165.890 56.310 166.090 ;
        RECT 26.345 165.750 31.850 165.890 ;
        RECT 41.600 165.750 56.310 165.890 ;
        RECT 56.690 165.890 57.010 165.950 ;
        RECT 57.625 165.890 57.915 165.935 ;
        RECT 56.690 165.750 57.915 165.890 ;
        RECT 58.160 165.890 58.300 166.090 ;
        RECT 71.870 166.030 72.190 166.090 ;
        RECT 73.250 166.230 73.570 166.290 ;
        RECT 76.560 166.230 76.700 166.385 ;
        RECT 77.850 166.370 78.170 166.630 ;
        RECT 78.770 166.370 79.090 166.630 ;
        RECT 83.000 166.615 83.140 166.770 ;
        RECT 88.430 166.710 88.750 166.770 ;
        RECT 93.045 166.725 93.335 166.955 ;
        RECT 93.490 166.710 93.810 166.970 ;
        RECT 101.310 166.910 101.630 166.970 ;
        RECT 103.240 166.910 103.380 167.110 ;
        RECT 94.960 166.770 100.620 166.910 ;
        RECT 82.925 166.385 83.215 166.615 ;
        RECT 84.750 166.370 85.070 166.630 ;
        RECT 86.145 166.385 86.435 166.615 ;
        RECT 87.525 166.570 87.815 166.615 ;
        RECT 87.970 166.570 88.290 166.630 ;
        RECT 87.525 166.430 88.290 166.570 ;
        RECT 87.525 166.385 87.815 166.430 ;
        RECT 73.250 166.090 76.700 166.230 ;
        RECT 76.930 166.230 77.250 166.290 ;
        RECT 86.220 166.230 86.360 166.385 ;
        RECT 87.970 166.370 88.290 166.430 ;
        RECT 90.285 166.570 90.575 166.615 ;
        RECT 91.190 166.570 91.510 166.630 ;
        RECT 90.285 166.430 91.510 166.570 ;
        RECT 90.285 166.385 90.575 166.430 ;
        RECT 91.190 166.370 91.510 166.430 ;
        RECT 92.110 166.570 92.430 166.630 ;
        RECT 92.585 166.570 92.875 166.615 ;
        RECT 94.425 166.570 94.715 166.615 ;
        RECT 92.110 166.430 92.875 166.570 ;
        RECT 92.110 166.370 92.430 166.430 ;
        RECT 92.585 166.385 92.875 166.430 ;
        RECT 93.120 166.430 94.715 166.570 ;
        RECT 92.200 166.230 92.340 166.370 ;
        RECT 93.120 166.290 93.260 166.430 ;
        RECT 94.425 166.385 94.715 166.430 ;
        RECT 76.930 166.090 86.360 166.230 ;
        RECT 89.440 166.090 92.340 166.230 ;
        RECT 73.250 166.030 73.570 166.090 ;
        RECT 76.930 166.030 77.250 166.090 ;
        RECT 79.230 165.890 79.550 165.950 ;
        RECT 87.510 165.890 87.830 165.950 ;
        RECT 58.160 165.750 79.550 165.890 ;
        RECT 26.345 165.705 26.635 165.750 ;
        RECT 31.710 165.550 31.850 165.750 ;
        RECT 41.970 165.690 42.290 165.750 ;
        RECT 50.710 165.690 51.030 165.750 ;
        RECT 56.690 165.690 57.010 165.750 ;
        RECT 57.625 165.705 57.915 165.750 ;
        RECT 79.230 165.690 79.550 165.750 ;
        RECT 79.780 165.750 87.830 165.890 ;
        RECT 47.490 165.550 47.810 165.610 ;
        RECT 31.710 165.410 47.810 165.550 ;
        RECT 47.490 165.350 47.810 165.410 ;
        RECT 47.950 165.350 48.270 165.610 ;
        RECT 49.790 165.350 50.110 165.610 ;
        RECT 50.250 165.550 50.570 165.610 ;
        RECT 79.780 165.550 79.920 165.750 ;
        RECT 87.510 165.690 87.830 165.750 ;
        RECT 88.445 165.890 88.735 165.935 ;
        RECT 88.890 165.890 89.210 165.950 ;
        RECT 89.440 165.935 89.580 166.090 ;
        RECT 93.030 166.030 93.350 166.290 ;
        RECT 93.950 166.230 94.270 166.290 ;
        RECT 94.960 166.230 95.100 166.770 ;
        RECT 95.790 166.370 96.110 166.630 ;
        RECT 97.185 166.570 97.475 166.615 ;
        RECT 96.340 166.430 97.475 166.570 ;
        RECT 96.340 166.290 96.480 166.430 ;
        RECT 97.185 166.385 97.475 166.430 ;
        RECT 97.630 166.370 97.950 166.630 ;
        RECT 98.090 166.370 98.410 166.630 ;
        RECT 100.480 166.615 100.620 166.770 ;
        RECT 101.310 166.770 103.380 166.910 ;
        RECT 103.625 166.910 103.915 166.955 ;
        RECT 105.910 166.910 106.230 166.970 ;
        RECT 103.625 166.770 106.230 166.910 ;
        RECT 101.310 166.710 101.630 166.770 ;
        RECT 103.625 166.725 103.915 166.770 ;
        RECT 105.910 166.710 106.230 166.770 ;
        RECT 99.025 166.385 99.315 166.615 ;
        RECT 100.405 166.385 100.695 166.615 ;
        RECT 93.950 166.090 95.100 166.230 ;
        RECT 93.950 166.030 94.270 166.090 ;
        RECT 96.250 166.030 96.570 166.290 ;
        RECT 96.710 166.230 97.030 166.290 ;
        RECT 99.100 166.230 99.240 166.385 ;
        RECT 104.070 166.370 104.390 166.630 ;
        RECT 104.990 166.570 105.310 166.630 ;
        RECT 104.795 166.430 105.310 166.570 ;
        RECT 104.990 166.370 105.310 166.430 ;
        RECT 105.450 166.370 105.770 166.630 ;
        RECT 106.920 166.615 107.060 167.110 ;
        RECT 107.305 167.110 123.710 167.250 ;
        RECT 107.305 167.065 107.595 167.110 ;
        RECT 123.390 167.050 123.710 167.110 ;
        RECT 126.150 167.250 126.470 167.310 ;
        RECT 130.290 167.250 130.610 167.310 ;
        RECT 126.150 167.110 130.610 167.250 ;
        RECT 126.150 167.050 126.470 167.110 ;
        RECT 130.290 167.050 130.610 167.110 ;
        RECT 133.050 167.250 133.370 167.310 ;
        RECT 133.525 167.250 133.815 167.295 ;
        RECT 133.050 167.110 133.815 167.250 ;
        RECT 133.050 167.050 133.370 167.110 ;
        RECT 133.525 167.065 133.815 167.110 ;
        RECT 107.750 166.910 108.070 166.970 ;
        RECT 107.750 166.770 109.360 166.910 ;
        RECT 107.750 166.710 108.070 166.770 ;
        RECT 109.220 166.615 109.360 166.770 ;
        RECT 118.790 166.710 119.110 166.970 ;
        RECT 122.010 166.910 122.330 166.970 ;
        RECT 122.010 166.770 127.300 166.910 ;
        RECT 122.010 166.710 122.330 166.770 ;
        RECT 127.160 166.630 127.300 166.770 ;
        RECT 106.845 166.385 107.135 166.615 ;
        RECT 108.225 166.385 108.515 166.615 ;
        RECT 109.145 166.385 109.435 166.615 ;
        RECT 109.605 166.570 109.895 166.615 ;
        RECT 110.050 166.570 110.370 166.630 ;
        RECT 109.605 166.430 110.370 166.570 ;
        RECT 109.605 166.385 109.895 166.430 ;
        RECT 105.925 166.230 106.215 166.275 ;
        RECT 108.300 166.230 108.440 166.385 ;
        RECT 110.050 166.370 110.370 166.430 ;
        RECT 112.350 166.570 112.670 166.630 ;
        RECT 123.850 166.570 124.170 166.630 ;
        RECT 112.350 166.430 124.170 166.570 ;
        RECT 112.350 166.370 112.670 166.430 ;
        RECT 123.850 166.370 124.170 166.430 ;
        RECT 124.310 166.570 124.630 166.630 ;
        RECT 124.785 166.570 125.075 166.615 ;
        RECT 124.310 166.430 125.075 166.570 ;
        RECT 124.310 166.370 124.630 166.430 ;
        RECT 124.785 166.385 125.075 166.430 ;
        RECT 126.150 166.370 126.470 166.630 ;
        RECT 127.070 166.370 127.390 166.630 ;
        RECT 132.145 166.570 132.435 166.615 ;
        RECT 132.590 166.570 132.910 166.630 ;
        RECT 132.145 166.430 132.910 166.570 ;
        RECT 132.145 166.385 132.435 166.430 ;
        RECT 132.590 166.370 132.910 166.430 ;
        RECT 133.050 166.370 133.370 166.630 ;
        RECT 133.510 166.570 133.830 166.630 ;
        RECT 134.445 166.570 134.735 166.615 ;
        RECT 133.510 166.430 134.735 166.570 ;
        RECT 133.510 166.370 133.830 166.430 ;
        RECT 134.445 166.385 134.735 166.430 ;
        RECT 96.710 166.090 106.215 166.230 ;
        RECT 96.710 166.030 97.030 166.090 ;
        RECT 105.925 166.045 106.215 166.090 ;
        RECT 106.460 166.090 108.440 166.230 ;
        RECT 88.445 165.750 89.210 165.890 ;
        RECT 88.445 165.705 88.735 165.750 ;
        RECT 88.890 165.690 89.210 165.750 ;
        RECT 89.365 165.705 89.655 165.935 ;
        RECT 89.810 165.890 90.130 165.950 ;
        RECT 91.665 165.890 91.955 165.935 ;
        RECT 106.460 165.890 106.600 166.090 ;
        RECT 108.670 166.030 108.990 166.290 ;
        RECT 121.550 166.230 121.870 166.290 ;
        RECT 125.705 166.230 125.995 166.275 ;
        RECT 126.610 166.230 126.930 166.290 ;
        RECT 129.845 166.230 130.135 166.275 ;
        RECT 121.550 166.090 125.460 166.230 ;
        RECT 121.550 166.030 121.870 166.090 ;
        RECT 123.865 165.890 124.155 165.935 ;
        RECT 89.810 165.750 106.600 165.890 ;
        RECT 106.920 165.750 124.155 165.890 ;
        RECT 125.320 165.890 125.460 166.090 ;
        RECT 125.705 166.090 126.930 166.230 ;
        RECT 125.705 166.045 125.995 166.090 ;
        RECT 126.610 166.030 126.930 166.090 ;
        RECT 127.160 166.090 130.135 166.230 ;
        RECT 127.160 165.890 127.300 166.090 ;
        RECT 129.845 166.045 130.135 166.090 ;
        RECT 125.320 165.750 127.300 165.890 ;
        RECT 127.990 165.890 128.310 165.950 ;
        RECT 129.385 165.890 129.675 165.935 ;
        RECT 127.990 165.750 129.675 165.890 ;
        RECT 89.810 165.690 90.130 165.750 ;
        RECT 91.665 165.705 91.955 165.750 ;
        RECT 50.250 165.410 79.920 165.550 ;
        RECT 82.005 165.550 82.295 165.595 ;
        RECT 83.370 165.550 83.690 165.610 ;
        RECT 82.005 165.410 83.690 165.550 ;
        RECT 50.250 165.350 50.570 165.410 ;
        RECT 82.005 165.365 82.295 165.410 ;
        RECT 83.370 165.350 83.690 165.410 ;
        RECT 83.830 165.350 84.150 165.610 ;
        RECT 85.670 165.350 85.990 165.610 ;
        RECT 87.050 165.350 87.370 165.610 ;
        RECT 87.970 165.550 88.290 165.610 ;
        RECT 90.745 165.550 91.035 165.595 ;
        RECT 87.970 165.410 91.035 165.550 ;
        RECT 87.970 165.350 88.290 165.410 ;
        RECT 90.745 165.365 91.035 165.410 ;
        RECT 91.190 165.550 91.510 165.610 ;
        RECT 93.950 165.550 94.270 165.610 ;
        RECT 91.190 165.410 94.270 165.550 ;
        RECT 91.190 165.350 91.510 165.410 ;
        RECT 93.950 165.350 94.270 165.410 ;
        RECT 94.870 165.550 95.190 165.610 ;
        RECT 99.485 165.550 99.775 165.595 ;
        RECT 94.870 165.410 99.775 165.550 ;
        RECT 94.870 165.350 95.190 165.410 ;
        RECT 99.485 165.365 99.775 165.410 ;
        RECT 101.310 165.550 101.630 165.610 ;
        RECT 101.785 165.550 102.075 165.595 ;
        RECT 101.310 165.410 102.075 165.550 ;
        RECT 101.310 165.350 101.630 165.410 ;
        RECT 101.785 165.365 102.075 165.410 ;
        RECT 102.705 165.550 102.995 165.595 ;
        RECT 103.150 165.550 103.470 165.610 ;
        RECT 102.705 165.410 103.470 165.550 ;
        RECT 102.705 165.365 102.995 165.410 ;
        RECT 103.150 165.350 103.470 165.410 ;
        RECT 106.370 165.550 106.690 165.610 ;
        RECT 106.920 165.550 107.060 165.750 ;
        RECT 123.865 165.705 124.155 165.750 ;
        RECT 127.990 165.690 128.310 165.750 ;
        RECT 129.385 165.705 129.675 165.750 ;
        RECT 106.370 165.410 107.060 165.550 ;
        RECT 112.810 165.550 113.130 165.610 ;
        RECT 114.190 165.550 114.510 165.610 ;
        RECT 116.045 165.550 116.335 165.595 ;
        RECT 112.810 165.410 116.335 165.550 ;
        RECT 106.370 165.350 106.690 165.410 ;
        RECT 112.810 165.350 113.130 165.410 ;
        RECT 114.190 165.350 114.510 165.410 ;
        RECT 116.045 165.365 116.335 165.410 ;
        RECT 126.165 165.550 126.455 165.595 ;
        RECT 127.530 165.550 127.850 165.610 ;
        RECT 126.165 165.410 127.850 165.550 ;
        RECT 126.165 165.365 126.455 165.410 ;
        RECT 127.530 165.350 127.850 165.410 ;
        RECT 128.925 165.550 129.215 165.595 ;
        RECT 129.830 165.550 130.150 165.610 ;
        RECT 128.925 165.410 130.150 165.550 ;
        RECT 128.925 165.365 129.215 165.410 ;
        RECT 129.830 165.350 130.150 165.410 ;
        RECT 131.210 165.350 131.530 165.610 ;
        RECT 23.500 164.730 136.200 165.210 ;
        RECT 40.605 164.530 40.895 164.575 ;
        RECT 45.190 164.530 45.510 164.590 ;
        RECT 40.605 164.390 45.510 164.530 ;
        RECT 40.605 164.345 40.895 164.390 ;
        RECT 45.190 164.330 45.510 164.390 ;
        RECT 50.265 164.530 50.555 164.575 ;
        RECT 51.170 164.530 51.490 164.590 ;
        RECT 50.265 164.390 51.490 164.530 ;
        RECT 50.265 164.345 50.555 164.390 ;
        RECT 51.170 164.330 51.490 164.390 ;
        RECT 56.690 164.530 57.010 164.590 ;
        RECT 58.530 164.530 58.850 164.590 ;
        RECT 56.690 164.390 58.850 164.530 ;
        RECT 56.690 164.330 57.010 164.390 ;
        RECT 58.530 164.330 58.850 164.390 ;
        RECT 61.290 164.330 61.610 164.590 ;
        RECT 61.750 164.530 62.070 164.590 ;
        RECT 63.145 164.530 63.435 164.575 ;
        RECT 61.750 164.390 63.435 164.530 ;
        RECT 61.750 164.330 62.070 164.390 ;
        RECT 63.145 164.345 63.435 164.390 ;
        RECT 71.870 164.530 72.190 164.590 ;
        RECT 75.550 164.530 75.870 164.590 ;
        RECT 81.530 164.530 81.850 164.590 ;
        RECT 71.870 164.390 75.870 164.530 ;
        RECT 71.870 164.330 72.190 164.390 ;
        RECT 75.550 164.330 75.870 164.390 ;
        RECT 77.020 164.390 81.850 164.530 ;
        RECT 40.145 164.190 40.435 164.235 ;
        RECT 41.510 164.190 41.830 164.250 ;
        RECT 40.145 164.050 41.830 164.190 ;
        RECT 40.145 164.005 40.435 164.050 ;
        RECT 41.510 163.990 41.830 164.050 ;
        RECT 42.430 164.190 42.750 164.250 ;
        RECT 43.365 164.190 43.655 164.235 ;
        RECT 44.270 164.190 44.590 164.250 ;
        RECT 42.430 164.050 44.590 164.190 ;
        RECT 42.430 163.990 42.750 164.050 ;
        RECT 43.365 164.005 43.655 164.050 ;
        RECT 44.270 163.990 44.590 164.050 ;
        RECT 47.490 164.190 47.810 164.250 ;
        RECT 55.310 164.190 55.630 164.250 ;
        RECT 57.610 164.190 57.930 164.250 ;
        RECT 47.490 164.050 59.680 164.190 ;
        RECT 47.490 163.990 47.810 164.050 ;
        RECT 55.310 163.990 55.630 164.050 ;
        RECT 57.610 163.990 57.930 164.050 ;
        RECT 43.810 163.650 44.130 163.910 ;
        RECT 49.790 163.850 50.110 163.910 ;
        RECT 47.580 163.710 50.110 163.850 ;
        RECT 47.580 163.555 47.720 163.710 ;
        RECT 49.790 163.650 50.110 163.710 ;
        RECT 54.405 163.850 54.695 163.895 ;
        RECT 59.540 163.850 59.680 164.050 ;
        RECT 74.170 163.990 74.490 164.250 ;
        RECT 60.830 163.850 61.150 163.910 ;
        RECT 54.405 163.710 58.760 163.850 ;
        RECT 54.405 163.665 54.695 163.710 ;
        RECT 47.505 163.325 47.795 163.555 ;
        RECT 47.950 163.310 48.270 163.570 ;
        RECT 48.870 163.310 49.190 163.570 ;
        RECT 49.345 163.510 49.635 163.555 ;
        RECT 53.470 163.510 53.790 163.570 ;
        RECT 49.345 163.370 53.790 163.510 ;
        RECT 49.345 163.325 49.635 163.370 ;
        RECT 53.470 163.310 53.790 163.370 ;
        RECT 53.930 163.310 54.250 163.570 ;
        RECT 54.865 163.325 55.155 163.555 ;
        RECT 38.290 162.970 38.610 163.230 ;
        RECT 41.510 162.970 41.830 163.230 ;
        RECT 54.940 163.170 55.080 163.325 ;
        RECT 55.310 163.310 55.630 163.570 ;
        RECT 56.230 163.555 56.550 163.570 ;
        RECT 56.095 163.510 56.550 163.555 ;
        RECT 56.095 163.370 57.840 163.510 ;
        RECT 56.095 163.325 56.550 163.370 ;
        RECT 56.230 163.310 56.550 163.325 ;
        RECT 56.690 163.170 57.010 163.230 ;
        RECT 54.940 163.030 57.010 163.170 ;
        RECT 57.700 163.170 57.840 163.370 ;
        RECT 58.070 163.310 58.390 163.570 ;
        RECT 58.620 163.555 58.760 163.710 ;
        RECT 59.540 163.710 61.150 163.850 ;
        RECT 59.540 163.555 59.680 163.710 ;
        RECT 60.830 163.650 61.150 163.710 ;
        RECT 73.250 163.850 73.570 163.910 ;
        RECT 75.090 163.850 75.410 163.910 ;
        RECT 73.250 163.710 75.410 163.850 ;
        RECT 73.250 163.650 73.570 163.710 ;
        RECT 75.090 163.650 75.410 163.710 ;
        RECT 58.545 163.325 58.835 163.555 ;
        RECT 59.465 163.325 59.755 163.555 ;
        RECT 60.385 163.510 60.675 163.555 ;
        RECT 63.130 163.510 63.450 163.570 ;
        RECT 60.385 163.370 63.450 163.510 ;
        RECT 60.385 163.325 60.675 163.370 ;
        RECT 63.130 163.310 63.450 163.370 ;
        RECT 64.050 163.310 64.370 163.570 ;
        RECT 66.350 163.510 66.670 163.570 ;
        RECT 72.345 163.510 72.635 163.555 ;
        RECT 66.350 163.370 72.635 163.510 ;
        RECT 66.350 163.310 66.670 163.370 ;
        RECT 72.345 163.325 72.635 163.370 ;
        RECT 58.990 163.170 59.310 163.230 ;
        RECT 59.925 163.170 60.215 163.215 ;
        RECT 57.700 163.030 60.215 163.170 ;
        RECT 72.420 163.170 72.560 163.325 ;
        RECT 73.710 163.310 74.030 163.570 ;
        RECT 75.550 163.310 75.870 163.570 ;
        RECT 77.020 163.555 77.160 164.390 ;
        RECT 81.530 164.330 81.850 164.390 ;
        RECT 81.990 164.530 82.310 164.590 ;
        RECT 82.925 164.530 83.215 164.575 ;
        RECT 89.810 164.530 90.130 164.590 ;
        RECT 97.630 164.530 97.950 164.590 ;
        RECT 81.990 164.390 83.215 164.530 ;
        RECT 81.990 164.330 82.310 164.390 ;
        RECT 82.925 164.345 83.215 164.390 ;
        RECT 84.840 164.390 90.130 164.530 ;
        RECT 77.865 164.190 78.155 164.235 ;
        RECT 84.840 164.190 84.980 164.390 ;
        RECT 89.810 164.330 90.130 164.390 ;
        RECT 91.280 164.390 97.950 164.530 ;
        RECT 77.865 164.050 84.980 164.190 ;
        RECT 85.225 164.190 85.515 164.235 ;
        RECT 86.130 164.190 86.450 164.250 ;
        RECT 85.225 164.050 86.450 164.190 ;
        RECT 77.865 164.005 78.155 164.050 ;
        RECT 85.225 164.005 85.515 164.050 ;
        RECT 86.130 163.990 86.450 164.050 ;
        RECT 88.890 163.850 89.210 163.910 ;
        RECT 79.320 163.710 89.210 163.850 ;
        RECT 79.320 163.555 79.460 163.710 ;
        RECT 88.890 163.650 89.210 163.710 ;
        RECT 76.945 163.325 77.235 163.555 ;
        RECT 79.245 163.325 79.535 163.555 ;
        RECT 79.705 163.325 79.995 163.555 ;
        RECT 80.150 163.510 80.470 163.570 ;
        RECT 81.990 163.555 82.310 163.570 ;
        RECT 80.150 163.370 80.665 163.510 ;
        RECT 74.185 163.170 74.475 163.215 ;
        RECT 72.420 163.030 74.475 163.170 ;
        RECT 56.690 162.970 57.010 163.030 ;
        RECT 58.990 162.970 59.310 163.030 ;
        RECT 59.925 162.985 60.215 163.030 ;
        RECT 74.185 162.985 74.475 163.030 ;
        RECT 74.630 163.170 74.950 163.230 ;
        RECT 78.310 163.170 78.630 163.230 ;
        RECT 74.630 163.030 78.630 163.170 ;
        RECT 74.630 162.970 74.950 163.030 ;
        RECT 78.310 162.970 78.630 163.030 ;
        RECT 57.150 162.630 57.470 162.890 ;
        RECT 71.425 162.830 71.715 162.875 ;
        RECT 72.330 162.830 72.650 162.890 ;
        RECT 71.425 162.690 72.650 162.830 ;
        RECT 71.425 162.645 71.715 162.690 ;
        RECT 72.330 162.630 72.650 162.690 ;
        RECT 73.265 162.830 73.555 162.875 ;
        RECT 73.710 162.830 74.030 162.890 ;
        RECT 75.105 162.830 75.395 162.875 ;
        RECT 77.390 162.830 77.710 162.890 ;
        RECT 73.265 162.690 77.710 162.830 ;
        RECT 73.265 162.645 73.555 162.690 ;
        RECT 73.710 162.630 74.030 162.690 ;
        RECT 75.105 162.645 75.395 162.690 ;
        RECT 77.390 162.630 77.710 162.690 ;
        RECT 78.770 162.630 79.090 162.890 ;
        RECT 79.780 162.830 79.920 163.325 ;
        RECT 80.150 163.310 80.470 163.370 ;
        RECT 81.990 163.325 82.320 163.555 ;
        RECT 81.990 163.310 82.310 163.325 ;
        RECT 83.830 163.310 84.150 163.570 ;
        RECT 84.290 163.310 84.610 163.570 ;
        RECT 86.145 163.510 86.435 163.555 ;
        RECT 86.590 163.510 86.910 163.570 ;
        RECT 86.145 163.370 86.910 163.510 ;
        RECT 86.145 163.325 86.435 163.370 ;
        RECT 86.590 163.310 86.910 163.370 ;
        RECT 87.510 163.510 87.830 163.570 ;
        RECT 90.270 163.555 90.590 163.570 ;
        RECT 89.365 163.510 89.655 163.555 ;
        RECT 87.510 163.370 89.655 163.510 ;
        RECT 87.510 163.310 87.830 163.370 ;
        RECT 89.365 163.325 89.655 163.370 ;
        RECT 90.135 163.325 90.590 163.555 ;
        RECT 90.270 163.310 90.590 163.325 ;
        RECT 81.070 162.970 81.390 163.230 ;
        RECT 81.545 163.170 81.835 163.215 ;
        RECT 84.380 163.170 84.520 163.310 ;
        RECT 91.280 163.215 91.420 164.390 ;
        RECT 97.630 164.330 97.950 164.390 ;
        RECT 98.105 164.530 98.395 164.575 ;
        RECT 100.390 164.530 100.710 164.590 ;
        RECT 98.105 164.390 100.710 164.530 ;
        RECT 98.105 164.345 98.395 164.390 ;
        RECT 100.390 164.330 100.710 164.390 ;
        RECT 102.690 164.530 103.010 164.590 ;
        RECT 121.550 164.530 121.870 164.590 ;
        RECT 102.690 164.390 121.870 164.530 ;
        RECT 102.690 164.330 103.010 164.390 ;
        RECT 121.550 164.330 121.870 164.390 ;
        RECT 124.770 164.330 125.090 164.590 ;
        RECT 92.110 164.190 92.430 164.250 ;
        RECT 99.010 164.190 99.330 164.250 ;
        RECT 92.110 164.050 99.330 164.190 ;
        RECT 92.110 163.990 92.430 164.050 ;
        RECT 99.010 163.990 99.330 164.050 ;
        RECT 99.930 164.190 100.250 164.250 ;
        RECT 105.925 164.190 106.215 164.235 ;
        RECT 110.510 164.190 110.830 164.250 ;
        RECT 99.930 164.050 110.830 164.190 ;
        RECT 99.930 163.990 100.250 164.050 ;
        RECT 105.925 164.005 106.215 164.050 ;
        RECT 110.510 163.990 110.830 164.050 ;
        RECT 120.645 164.005 120.935 164.235 ;
        RECT 95.790 163.850 96.110 163.910 ;
        RECT 120.720 163.850 120.860 164.005 ;
        RECT 93.120 163.710 120.860 163.850 ;
        RECT 129.370 163.850 129.690 163.910 ;
        RECT 129.370 163.710 133.280 163.850 ;
        RECT 93.120 163.555 93.260 163.710 ;
        RECT 95.790 163.650 96.110 163.710 ;
        RECT 129.370 163.650 129.690 163.710 ;
        RECT 93.045 163.325 93.335 163.555 ;
        RECT 94.425 163.510 94.715 163.555 ;
        RECT 98.090 163.510 98.410 163.570 ;
        RECT 94.425 163.370 98.410 163.510 ;
        RECT 94.425 163.325 94.715 163.370 ;
        RECT 81.545 163.030 84.520 163.170 ;
        RECT 85.225 163.170 85.515 163.215 ;
        RECT 91.205 163.170 91.495 163.215 ;
        RECT 85.225 163.030 91.495 163.170 ;
        RECT 81.545 162.985 81.835 163.030 ;
        RECT 85.225 162.985 85.515 163.030 ;
        RECT 91.205 162.985 91.495 163.030 ;
        RECT 92.570 162.970 92.890 163.230 ;
        RECT 82.910 162.830 83.230 162.890 ;
        RECT 79.780 162.690 83.230 162.830 ;
        RECT 82.910 162.630 83.230 162.690 ;
        RECT 84.290 162.630 84.610 162.890 ;
        RECT 87.525 162.830 87.815 162.875 ;
        RECT 88.430 162.830 88.750 162.890 ;
        RECT 87.525 162.690 88.750 162.830 ;
        RECT 87.525 162.645 87.815 162.690 ;
        RECT 88.430 162.630 88.750 162.690 ;
        RECT 92.110 162.830 92.430 162.890 ;
        RECT 94.500 162.830 94.640 163.325 ;
        RECT 98.090 163.310 98.410 163.370 ;
        RECT 99.010 163.310 99.330 163.570 ;
        RECT 99.470 163.510 99.790 163.570 ;
        RECT 99.945 163.510 100.235 163.555 ;
        RECT 99.470 163.370 100.235 163.510 ;
        RECT 99.470 163.310 99.790 163.370 ;
        RECT 99.945 163.325 100.235 163.370 ;
        RECT 100.390 163.310 100.710 163.570 ;
        RECT 100.850 163.510 101.170 163.570 ;
        RECT 102.705 163.510 102.995 163.555 ;
        RECT 100.850 163.370 102.995 163.510 ;
        RECT 100.850 163.310 101.170 163.370 ;
        RECT 102.705 163.325 102.995 163.370 ;
        RECT 103.150 163.310 103.470 163.570 ;
        RECT 104.070 163.310 104.390 163.570 ;
        RECT 113.285 163.510 113.575 163.555 ;
        RECT 120.630 163.510 120.950 163.570 ;
        RECT 113.285 163.370 120.950 163.510 ;
        RECT 113.285 163.325 113.575 163.370 ;
        RECT 120.630 163.310 120.950 163.370 ;
        RECT 130.750 163.510 131.070 163.570 ;
        RECT 133.140 163.555 133.280 163.710 ;
        RECT 132.145 163.510 132.435 163.555 ;
        RECT 130.750 163.370 132.435 163.510 ;
        RECT 130.750 163.310 131.070 163.370 ;
        RECT 132.145 163.325 132.435 163.370 ;
        RECT 133.065 163.510 133.355 163.555 ;
        RECT 133.510 163.510 133.830 163.570 ;
        RECT 133.065 163.370 133.830 163.510 ;
        RECT 133.065 163.325 133.355 163.370 ;
        RECT 133.510 163.310 133.830 163.370 ;
        RECT 96.725 163.170 97.015 163.215 ;
        RECT 101.770 163.170 102.090 163.230 ;
        RECT 96.725 163.030 102.090 163.170 ;
        RECT 96.725 162.985 97.015 163.030 ;
        RECT 101.770 162.970 102.090 163.030 ;
        RECT 114.190 162.970 114.510 163.230 ;
        RECT 92.110 162.690 94.640 162.830 ;
        RECT 99.470 162.830 99.790 162.890 ;
        RECT 100.865 162.830 101.155 162.875 ;
        RECT 103.610 162.830 103.930 162.890 ;
        RECT 105.450 162.830 105.770 162.890 ;
        RECT 99.470 162.690 105.770 162.830 ;
        RECT 92.110 162.630 92.430 162.690 ;
        RECT 99.470 162.630 99.790 162.690 ;
        RECT 100.865 162.645 101.155 162.690 ;
        RECT 103.610 162.630 103.930 162.690 ;
        RECT 105.450 162.630 105.770 162.690 ;
        RECT 133.970 162.630 134.290 162.890 ;
        RECT 23.500 162.010 136.200 162.490 ;
        RECT 41.970 161.810 42.290 161.870 ;
        RECT 42.905 161.810 43.195 161.855 ;
        RECT 41.970 161.670 43.195 161.810 ;
        RECT 41.970 161.610 42.290 161.670 ;
        RECT 42.905 161.625 43.195 161.670 ;
        RECT 45.665 161.810 45.955 161.855 ;
        RECT 50.250 161.810 50.570 161.870 ;
        RECT 45.665 161.670 50.570 161.810 ;
        RECT 45.665 161.625 45.955 161.670 ;
        RECT 39.225 161.470 39.515 161.515 ;
        RECT 41.050 161.470 41.370 161.530 ;
        RECT 39.225 161.330 41.370 161.470 ;
        RECT 39.225 161.285 39.515 161.330 ;
        RECT 41.050 161.270 41.370 161.330 ;
        RECT 41.510 161.470 41.830 161.530 ;
        RECT 45.740 161.470 45.880 161.625 ;
        RECT 50.250 161.610 50.570 161.670 ;
        RECT 56.690 161.810 57.010 161.870 ;
        RECT 59.910 161.810 60.230 161.870 ;
        RECT 61.305 161.810 61.595 161.855 ;
        RECT 76.565 161.810 76.855 161.855 ;
        RECT 56.690 161.670 61.595 161.810 ;
        RECT 56.690 161.610 57.010 161.670 ;
        RECT 59.910 161.610 60.230 161.670 ;
        RECT 61.305 161.625 61.595 161.670 ;
        RECT 72.420 161.670 76.855 161.810 ;
        RECT 72.420 161.530 72.560 161.670 ;
        RECT 76.565 161.625 76.855 161.670 ;
        RECT 78.310 161.810 78.630 161.870 ;
        RECT 78.865 161.810 79.155 161.855 ;
        RECT 82.005 161.810 82.295 161.855 ;
        RECT 84.290 161.810 84.610 161.870 ;
        RECT 78.310 161.670 79.155 161.810 ;
        RECT 78.310 161.610 78.630 161.670 ;
        RECT 78.865 161.625 79.155 161.670 ;
        RECT 80.325 161.670 84.610 161.810 ;
        RECT 41.510 161.330 45.880 161.470 ;
        RECT 41.510 161.270 41.830 161.330 ;
        RECT 38.290 161.130 38.610 161.190 ;
        RECT 43.825 161.130 44.115 161.175 ;
        RECT 44.270 161.130 44.590 161.190 ;
        RECT 44.820 161.175 44.960 161.330 ;
        RECT 46.110 161.270 46.430 161.530 ;
        RECT 62.225 161.470 62.515 161.515 ;
        RECT 58.620 161.330 62.515 161.470 ;
        RECT 38.290 160.990 44.590 161.130 ;
        RECT 38.290 160.930 38.610 160.990 ;
        RECT 43.825 160.945 44.115 160.990 ;
        RECT 44.270 160.930 44.590 160.990 ;
        RECT 44.745 160.945 45.035 161.175 ;
        RECT 55.310 161.130 55.630 161.190 ;
        RECT 55.785 161.130 56.075 161.175 ;
        RECT 55.310 160.990 56.075 161.130 ;
        RECT 55.310 160.930 55.630 160.990 ;
        RECT 55.785 160.945 56.075 160.990 ;
        RECT 56.690 160.930 57.010 161.190 ;
        RECT 58.620 161.175 58.760 161.330 ;
        RECT 62.225 161.285 62.515 161.330 ;
        RECT 63.130 161.470 63.450 161.530 ;
        RECT 65.905 161.470 66.195 161.515 ;
        RECT 63.130 161.330 66.195 161.470 ;
        RECT 63.130 161.270 63.450 161.330 ;
        RECT 65.905 161.285 66.195 161.330 ;
        RECT 72.330 161.270 72.650 161.530 ;
        RECT 74.630 161.470 74.950 161.530 ;
        RECT 73.340 161.330 74.950 161.470 ;
        RECT 58.545 160.945 58.835 161.175 ;
        RECT 44.360 160.110 44.500 160.930 ;
        RECT 56.245 160.790 56.535 160.835 ;
        RECT 58.620 160.790 58.760 160.945 ;
        RECT 58.990 160.930 59.310 161.190 ;
        RECT 59.465 161.130 59.755 161.175 ;
        RECT 59.465 160.990 60.140 161.130 ;
        RECT 59.465 160.945 59.755 160.990 ;
        RECT 56.245 160.650 58.760 160.790 ;
        RECT 56.245 160.605 56.535 160.650 ;
        RECT 57.625 160.450 57.915 160.495 ;
        RECT 59.450 160.450 59.770 160.510 ;
        RECT 57.625 160.310 59.770 160.450 ;
        RECT 60.000 160.450 60.140 160.990 ;
        RECT 60.370 160.930 60.690 161.190 ;
        RECT 60.845 160.945 61.135 161.175 ;
        RECT 61.750 161.130 62.070 161.190 ;
        RECT 63.605 161.130 63.895 161.175 ;
        RECT 64.050 161.130 64.370 161.190 ;
        RECT 61.750 160.990 64.370 161.130 ;
        RECT 60.920 160.790 61.060 160.945 ;
        RECT 61.750 160.930 62.070 160.990 ;
        RECT 63.605 160.945 63.895 160.990 ;
        RECT 64.050 160.930 64.370 160.990 ;
        RECT 64.525 160.945 64.815 161.175 ;
        RECT 64.970 161.130 65.290 161.190 ;
        RECT 65.445 161.130 65.735 161.175 ;
        RECT 64.970 160.990 65.735 161.130 ;
        RECT 64.600 160.790 64.740 160.945 ;
        RECT 64.970 160.930 65.290 160.990 ;
        RECT 65.445 160.945 65.735 160.990 ;
        RECT 66.350 160.930 66.670 161.190 ;
        RECT 73.340 161.175 73.480 161.330 ;
        RECT 74.630 161.270 74.950 161.330 ;
        RECT 75.550 161.470 75.870 161.530 ;
        RECT 77.865 161.470 78.155 161.515 ;
        RECT 75.550 161.330 78.155 161.470 ;
        RECT 75.550 161.270 75.870 161.330 ;
        RECT 77.865 161.285 78.155 161.330 ;
        RECT 73.265 160.945 73.555 161.175 ;
        RECT 73.725 160.945 74.015 161.175 ;
        RECT 80.325 161.130 80.465 161.670 ;
        RECT 82.005 161.625 82.295 161.670 ;
        RECT 84.290 161.610 84.610 161.670 ;
        RECT 88.890 161.810 89.210 161.870 ;
        RECT 93.030 161.810 93.350 161.870 ;
        RECT 88.890 161.670 93.350 161.810 ;
        RECT 88.890 161.610 89.210 161.670 ;
        RECT 93.030 161.610 93.350 161.670 ;
        RECT 93.965 161.810 94.255 161.855 ;
        RECT 94.410 161.810 94.730 161.870 ;
        RECT 103.150 161.810 103.470 161.870 ;
        RECT 124.770 161.810 125.090 161.870 ;
        RECT 93.965 161.670 103.470 161.810 ;
        RECT 93.965 161.625 94.255 161.670 ;
        RECT 94.410 161.610 94.730 161.670 ;
        RECT 103.150 161.610 103.470 161.670 ;
        RECT 122.100 161.670 125.090 161.810 ;
        RECT 82.925 161.470 83.215 161.515 ;
        RECT 92.125 161.470 92.415 161.515 ;
        RECT 96.250 161.470 96.570 161.530 ;
        RECT 99.010 161.470 99.330 161.530 ;
        RECT 116.490 161.470 116.810 161.530 ;
        RECT 122.100 161.515 122.240 161.670 ;
        RECT 124.770 161.610 125.090 161.670 ;
        RECT 82.925 161.330 98.780 161.470 ;
        RECT 82.925 161.285 83.215 161.330 ;
        RECT 92.125 161.285 92.415 161.330 ;
        RECT 96.250 161.270 96.570 161.330 ;
        RECT 76.640 160.990 80.465 161.130 ;
        RECT 66.440 160.790 66.580 160.930 ;
        RECT 60.920 160.650 63.820 160.790 ;
        RECT 64.600 160.650 66.580 160.790 ;
        RECT 60.830 160.450 61.150 160.510 ;
        RECT 63.680 160.495 63.820 160.650 ;
        RECT 60.000 160.310 61.150 160.450 ;
        RECT 57.625 160.265 57.915 160.310 ;
        RECT 59.450 160.250 59.770 160.310 ;
        RECT 60.830 160.250 61.150 160.310 ;
        RECT 63.605 160.265 63.895 160.495 ;
        RECT 64.510 160.450 64.830 160.510 ;
        RECT 73.800 160.450 73.940 160.945 ;
        RECT 74.630 160.790 74.950 160.850 ;
        RECT 76.640 160.790 76.780 160.990 ;
        RECT 81.545 160.945 81.835 161.175 ;
        RECT 84.305 160.945 84.595 161.175 ;
        RECT 84.765 161.130 85.055 161.175 ;
        RECT 85.210 161.130 85.530 161.190 ;
        RECT 84.765 160.990 85.530 161.130 ;
        RECT 84.765 160.945 85.055 160.990 ;
        RECT 79.230 160.790 79.550 160.850 ;
        RECT 81.620 160.790 81.760 160.945 ;
        RECT 84.380 160.790 84.520 160.945 ;
        RECT 85.210 160.930 85.530 160.990 ;
        RECT 85.670 160.930 85.990 161.190 ;
        RECT 86.130 160.930 86.450 161.190 ;
        RECT 87.050 161.130 87.370 161.190 ;
        RECT 87.985 161.130 88.275 161.175 ;
        RECT 87.050 160.990 88.275 161.130 ;
        RECT 87.050 160.930 87.370 160.990 ;
        RECT 87.985 160.945 88.275 160.990 ;
        RECT 88.890 161.130 89.210 161.190 ;
        RECT 90.270 161.130 90.590 161.190 ;
        RECT 91.205 161.130 91.495 161.175 ;
        RECT 88.890 160.990 91.495 161.130 ;
        RECT 88.890 160.930 89.210 160.990 ;
        RECT 90.270 160.930 90.590 160.990 ;
        RECT 91.205 160.945 91.495 160.990 ;
        RECT 92.200 160.990 96.020 161.130 ;
        RECT 74.630 160.650 76.780 160.790 ;
        RECT 77.020 160.650 81.760 160.790 ;
        RECT 82.540 160.650 84.520 160.790 ;
        RECT 74.630 160.590 74.950 160.650 ;
        RECT 75.550 160.450 75.870 160.510 ;
        RECT 77.020 160.450 77.160 160.650 ;
        RECT 79.230 160.590 79.550 160.650 ;
        RECT 64.510 160.310 75.870 160.450 ;
        RECT 63.130 160.110 63.450 160.170 ;
        RECT 44.360 159.970 63.450 160.110 ;
        RECT 63.680 160.110 63.820 160.265 ;
        RECT 64.510 160.250 64.830 160.310 ;
        RECT 75.550 160.250 75.870 160.310 ;
        RECT 76.100 160.310 77.160 160.450 ;
        RECT 70.030 160.110 70.350 160.170 ;
        RECT 72.345 160.110 72.635 160.155 ;
        RECT 63.680 159.970 72.635 160.110 ;
        RECT 63.130 159.910 63.450 159.970 ;
        RECT 70.030 159.910 70.350 159.970 ;
        RECT 72.345 159.925 72.635 159.970 ;
        RECT 74.630 159.910 74.950 160.170 ;
        RECT 75.090 160.110 75.410 160.170 ;
        RECT 76.100 160.110 76.240 160.310 ;
        RECT 77.390 160.250 77.710 160.510 ;
        RECT 81.070 160.450 81.390 160.510 ;
        RECT 82.540 160.450 82.680 160.650 ;
        RECT 81.070 160.310 82.680 160.450 ;
        RECT 81.070 160.250 81.390 160.310 ;
        RECT 82.910 160.250 83.230 160.510 ;
        RECT 83.830 160.450 84.150 160.510 ;
        RECT 89.825 160.450 90.115 160.495 ;
        RECT 92.200 160.450 92.340 160.990 ;
        RECT 95.880 160.850 96.020 160.990 ;
        RECT 97.170 160.930 97.490 161.190 ;
        RECT 98.640 161.175 98.780 161.330 ;
        RECT 99.010 161.330 116.810 161.470 ;
        RECT 99.010 161.270 99.330 161.330 ;
        RECT 116.490 161.270 116.810 161.330 ;
        RECT 122.025 161.285 122.315 161.515 ;
        RECT 129.370 161.470 129.690 161.530 ;
        RECT 122.560 161.330 129.690 161.470 ;
        RECT 98.565 160.945 98.855 161.175 ;
        RECT 100.405 160.945 100.695 161.175 ;
        RECT 101.325 161.130 101.615 161.175 ;
        RECT 101.770 161.130 102.090 161.190 ;
        RECT 104.070 161.130 104.390 161.190 ;
        RECT 101.325 160.990 104.390 161.130 ;
        RECT 101.325 160.945 101.615 160.990 ;
        RECT 92.585 160.605 92.875 160.835 ;
        RECT 95.330 160.790 95.650 160.850 ;
        RECT 94.500 160.650 95.650 160.790 ;
        RECT 83.830 160.310 92.340 160.450 ;
        RECT 83.830 160.250 84.150 160.310 ;
        RECT 89.825 160.265 90.115 160.310 ;
        RECT 75.090 159.970 76.240 160.110 ;
        RECT 76.485 160.110 76.775 160.155 ;
        RECT 77.850 160.110 78.170 160.170 ;
        RECT 78.785 160.110 79.075 160.155 ;
        RECT 76.485 159.970 79.075 160.110 ;
        RECT 75.090 159.910 75.410 159.970 ;
        RECT 76.485 159.925 76.775 159.970 ;
        RECT 77.850 159.910 78.170 159.970 ;
        RECT 78.785 159.925 79.075 159.970 ;
        RECT 79.230 160.110 79.550 160.170 ;
        RECT 79.705 160.110 79.995 160.155 ;
        RECT 79.230 159.970 79.995 160.110 ;
        RECT 79.230 159.910 79.550 159.970 ;
        RECT 79.705 159.925 79.995 159.970 ;
        RECT 80.610 160.110 80.930 160.170 ;
        RECT 83.385 160.110 83.675 160.155 ;
        RECT 80.610 159.970 83.675 160.110 ;
        RECT 80.610 159.910 80.930 159.970 ;
        RECT 83.385 159.925 83.675 159.970 ;
        RECT 90.270 159.910 90.590 160.170 ;
        RECT 91.190 160.110 91.510 160.170 ;
        RECT 92.660 160.110 92.800 160.605 ;
        RECT 94.500 160.510 94.640 160.650 ;
        RECT 95.330 160.590 95.650 160.650 ;
        RECT 95.790 160.790 96.110 160.850 ;
        RECT 96.265 160.790 96.555 160.835 ;
        RECT 95.790 160.650 96.555 160.790 ;
        RECT 95.790 160.590 96.110 160.650 ;
        RECT 96.265 160.605 96.555 160.650 ;
        RECT 98.090 160.590 98.410 160.850 ;
        RECT 99.010 160.590 99.330 160.850 ;
        RECT 99.485 160.790 99.775 160.835 ;
        RECT 99.930 160.790 100.250 160.850 ;
        RECT 99.485 160.650 100.250 160.790 ;
        RECT 100.480 160.790 100.620 160.945 ;
        RECT 101.770 160.930 102.090 160.990 ;
        RECT 104.070 160.930 104.390 160.990 ;
        RECT 104.530 161.130 104.850 161.190 ;
        RECT 106.845 161.130 107.135 161.175 ;
        RECT 109.605 161.130 109.895 161.175 ;
        RECT 104.530 160.990 107.135 161.130 ;
        RECT 104.530 160.930 104.850 160.990 ;
        RECT 106.845 160.945 107.135 160.990 ;
        RECT 107.380 160.990 109.895 161.130 ;
        RECT 103.610 160.790 103.930 160.850 ;
        RECT 100.480 160.650 103.930 160.790 ;
        RECT 99.485 160.605 99.775 160.650 ;
        RECT 99.930 160.590 100.250 160.650 ;
        RECT 103.610 160.590 103.930 160.650 ;
        RECT 105.005 160.790 105.295 160.835 ;
        RECT 107.380 160.790 107.520 160.990 ;
        RECT 109.605 160.945 109.895 160.990 ;
        RECT 113.730 161.130 114.050 161.190 ;
        RECT 122.560 161.175 122.700 161.330 ;
        RECT 129.370 161.270 129.690 161.330 ;
        RECT 129.830 161.470 130.150 161.530 ;
        RECT 129.830 161.330 133.740 161.470 ;
        RECT 129.830 161.270 130.150 161.330 ;
        RECT 120.185 161.130 120.475 161.175 ;
        RECT 113.730 160.990 120.475 161.130 ;
        RECT 113.730 160.930 114.050 160.990 ;
        RECT 120.185 160.945 120.475 160.990 ;
        RECT 120.645 161.130 120.935 161.175 ;
        RECT 120.645 160.990 122.240 161.130 ;
        RECT 120.645 160.945 120.935 160.990 ;
        RECT 122.100 160.850 122.240 160.990 ;
        RECT 122.485 160.945 122.775 161.175 ;
        RECT 122.945 160.945 123.235 161.175 ;
        RECT 105.005 160.650 107.520 160.790 ;
        RECT 105.005 160.605 105.295 160.650 ;
        RECT 108.225 160.605 108.515 160.835 ;
        RECT 108.685 160.790 108.975 160.835 ;
        RECT 110.050 160.790 110.370 160.850 ;
        RECT 108.685 160.650 110.370 160.790 ;
        RECT 108.685 160.605 108.975 160.650 ;
        RECT 94.410 160.250 94.730 160.510 ;
        RECT 94.870 160.450 95.190 160.510 ;
        RECT 108.300 160.450 108.440 160.605 ;
        RECT 110.050 160.590 110.370 160.650 ;
        RECT 110.510 160.790 110.830 160.850 ;
        RECT 121.090 160.790 121.410 160.850 ;
        RECT 121.565 160.790 121.855 160.835 ;
        RECT 110.510 160.650 120.400 160.790 ;
        RECT 110.510 160.590 110.830 160.650 ;
        RECT 94.870 160.310 108.440 160.450 ;
        RECT 94.870 160.250 95.190 160.310 ;
        RECT 116.030 160.250 116.350 160.510 ;
        RECT 97.630 160.110 97.950 160.170 ;
        RECT 98.550 160.110 98.870 160.170 ;
        RECT 91.190 159.970 98.870 160.110 ;
        RECT 91.190 159.910 91.510 159.970 ;
        RECT 97.630 159.910 97.950 159.970 ;
        RECT 98.550 159.910 98.870 159.970 ;
        RECT 119.250 159.910 119.570 160.170 ;
        RECT 120.260 160.110 120.400 160.650 ;
        RECT 121.090 160.650 121.855 160.790 ;
        RECT 121.090 160.590 121.410 160.650 ;
        RECT 121.565 160.605 121.855 160.650 ;
        RECT 122.010 160.590 122.330 160.850 ;
        RECT 123.020 160.790 123.160 160.945 ;
        RECT 123.850 160.930 124.170 161.190 ;
        RECT 124.770 161.175 125.090 161.190 ;
        RECT 124.325 160.945 124.615 161.175 ;
        RECT 124.770 161.130 125.100 161.175 ;
        RECT 130.305 161.130 130.595 161.175 ;
        RECT 124.770 160.990 125.285 161.130 ;
        RECT 128.310 160.990 130.595 161.130 ;
        RECT 124.770 160.945 125.100 160.990 ;
        RECT 122.560 160.650 123.160 160.790 ;
        RECT 120.630 160.450 120.950 160.510 ;
        RECT 122.560 160.450 122.700 160.650 ;
        RECT 120.630 160.310 122.700 160.450 ;
        RECT 120.630 160.250 120.950 160.310 ;
        RECT 124.400 160.110 124.540 160.945 ;
        RECT 124.770 160.930 125.090 160.945 ;
        RECT 125.705 160.450 125.995 160.495 ;
        RECT 128.310 160.450 128.450 160.990 ;
        RECT 130.305 160.945 130.595 160.990 ;
        RECT 131.210 160.930 131.530 161.190 ;
        RECT 132.130 160.930 132.450 161.190 ;
        RECT 133.600 161.175 133.740 161.330 ;
        RECT 133.525 160.945 133.815 161.175 ;
        RECT 128.910 160.790 129.230 160.850 ;
        RECT 133.985 160.790 134.275 160.835 ;
        RECT 128.910 160.650 134.275 160.790 ;
        RECT 128.910 160.590 129.230 160.650 ;
        RECT 133.985 160.605 134.275 160.650 ;
        RECT 125.705 160.310 128.450 160.450 ;
        RECT 125.705 160.265 125.995 160.310 ;
        RECT 129.370 160.250 129.690 160.510 ;
        RECT 120.260 159.970 124.540 160.110 ;
        RECT 23.500 159.290 136.200 159.770 ;
        RECT 54.865 159.090 55.155 159.135 ;
        RECT 58.070 159.090 58.390 159.150 ;
        RECT 54.865 158.950 58.390 159.090 ;
        RECT 54.865 158.905 55.155 158.950 ;
        RECT 58.070 158.890 58.390 158.950 ;
        RECT 61.765 159.090 62.055 159.135 ;
        RECT 68.190 159.090 68.510 159.150 ;
        RECT 61.765 158.950 68.510 159.090 ;
        RECT 61.765 158.905 62.055 158.950 ;
        RECT 68.190 158.890 68.510 158.950 ;
        RECT 69.110 158.890 69.430 159.150 ;
        RECT 70.965 158.905 71.255 159.135 ;
        RECT 72.330 159.090 72.650 159.150 ;
        RECT 73.710 159.090 74.030 159.150 ;
        RECT 72.330 158.950 74.030 159.090 ;
        RECT 53.930 158.750 54.250 158.810 ;
        RECT 57.625 158.750 57.915 158.795 ;
        RECT 53.930 158.610 57.380 158.750 ;
        RECT 53.930 158.550 54.250 158.610 ;
        RECT 54.850 158.410 55.170 158.470 ;
        RECT 57.240 158.410 57.380 158.610 ;
        RECT 57.625 158.610 70.720 158.750 ;
        RECT 57.625 158.565 57.915 158.610 ;
        RECT 59.465 158.410 59.755 158.455 ;
        RECT 63.145 158.410 63.435 158.455 ;
        RECT 65.445 158.410 65.735 158.455 ;
        RECT 69.570 158.410 69.890 158.470 ;
        RECT 54.850 158.270 56.920 158.410 ;
        RECT 57.240 158.270 59.220 158.410 ;
        RECT 54.850 158.210 55.170 158.270 ;
        RECT 56.780 158.115 56.920 158.270 ;
        RECT 53.485 158.070 53.775 158.115 ;
        RECT 55.325 158.070 55.615 158.115 ;
        RECT 56.705 158.070 56.995 158.115 ;
        RECT 58.530 158.070 58.850 158.130 ;
        RECT 59.080 158.115 59.220 158.270 ;
        RECT 59.465 158.270 65.200 158.410 ;
        RECT 59.465 158.225 59.755 158.270 ;
        RECT 63.145 158.225 63.435 158.270 ;
        RECT 65.060 158.130 65.200 158.270 ;
        RECT 65.445 158.270 69.890 158.410 ;
        RECT 65.445 158.225 65.735 158.270 ;
        RECT 69.570 158.210 69.890 158.270 ;
        RECT 53.485 157.930 56.460 158.070 ;
        RECT 53.485 157.885 53.775 157.930 ;
        RECT 55.325 157.885 55.615 157.930 ;
        RECT 54.850 157.530 55.170 157.790 ;
        RECT 56.320 157.450 56.460 157.930 ;
        RECT 56.705 157.930 58.850 158.070 ;
        RECT 56.705 157.885 56.995 157.930 ;
        RECT 58.530 157.870 58.850 157.930 ;
        RECT 59.005 157.885 59.295 158.115 ;
        RECT 60.370 157.870 60.690 158.130 ;
        RECT 60.845 157.885 61.135 158.115 ;
        RECT 61.290 158.070 61.610 158.130 ;
        RECT 62.670 158.070 62.990 158.130 ;
        RECT 61.290 157.930 62.990 158.070 ;
        RECT 60.920 157.730 61.060 157.885 ;
        RECT 61.290 157.870 61.610 157.930 ;
        RECT 62.670 157.870 62.990 157.930 ;
        RECT 64.050 157.870 64.370 158.130 ;
        RECT 64.525 157.885 64.815 158.115 ;
        RECT 64.970 158.070 65.290 158.130 ;
        RECT 65.905 158.070 66.195 158.115 ;
        RECT 64.970 157.930 66.195 158.070 ;
        RECT 64.600 157.730 64.740 157.885 ;
        RECT 64.970 157.870 65.290 157.930 ;
        RECT 65.905 157.885 66.195 157.930 ;
        RECT 67.270 157.870 67.590 158.130 ;
        RECT 68.665 158.070 68.955 158.115 ;
        RECT 68.280 157.930 68.955 158.070 ;
        RECT 70.580 158.070 70.720 158.610 ;
        RECT 71.040 158.410 71.180 158.905 ;
        RECT 72.330 158.890 72.650 158.950 ;
        RECT 73.710 158.890 74.030 158.950 ;
        RECT 75.090 158.890 75.410 159.150 ;
        RECT 76.010 159.090 76.330 159.150 ;
        RECT 76.485 159.090 76.775 159.135 ;
        RECT 77.865 159.090 78.155 159.135 ;
        RECT 76.010 158.950 76.775 159.090 ;
        RECT 76.010 158.890 76.330 158.950 ;
        RECT 76.485 158.905 76.775 158.950 ;
        RECT 77.020 158.950 78.155 159.090 ;
        RECT 71.885 158.750 72.175 158.795 ;
        RECT 77.020 158.750 77.160 158.950 ;
        RECT 77.865 158.905 78.155 158.950 ;
        RECT 79.705 159.090 79.995 159.135 ;
        RECT 81.070 159.090 81.390 159.150 ;
        RECT 82.910 159.090 83.230 159.150 ;
        RECT 79.705 158.950 81.390 159.090 ;
        RECT 79.705 158.905 79.995 158.950 ;
        RECT 81.070 158.890 81.390 158.950 ;
        RECT 82.080 158.950 83.230 159.090 ;
        RECT 71.885 158.610 77.160 158.750 ;
        RECT 71.885 158.565 72.175 158.610 ;
        RECT 76.560 158.470 76.700 158.610 ;
        RECT 77.405 158.565 77.695 158.795 ;
        RECT 82.080 158.750 82.220 158.950 ;
        RECT 82.910 158.890 83.230 158.950 ;
        RECT 83.370 158.890 83.690 159.150 ;
        RECT 85.670 159.090 85.990 159.150 ;
        RECT 86.605 159.090 86.895 159.135 ;
        RECT 85.670 158.950 86.895 159.090 ;
        RECT 85.670 158.890 85.990 158.950 ;
        RECT 86.605 158.905 86.895 158.950 ;
        RECT 87.050 159.090 87.370 159.150 ;
        RECT 118.330 159.090 118.650 159.150 ;
        RECT 87.050 158.950 90.960 159.090 ;
        RECT 87.050 158.890 87.370 158.950 ;
        RECT 83.460 158.750 83.600 158.890 ;
        RECT 81.160 158.610 82.220 158.750 ;
        RECT 82.540 158.610 90.040 158.750 ;
        RECT 72.805 158.410 73.095 158.455 ;
        RECT 76.010 158.410 76.330 158.470 ;
        RECT 71.040 158.270 76.330 158.410 ;
        RECT 72.805 158.225 73.095 158.270 ;
        RECT 76.010 158.210 76.330 158.270 ;
        RECT 76.470 158.210 76.790 158.470 ;
        RECT 77.480 158.410 77.620 158.565 ;
        RECT 81.160 158.410 81.300 158.610 ;
        RECT 77.480 158.270 81.300 158.410 ;
        RECT 72.345 158.070 72.635 158.115 ;
        RECT 73.250 158.070 73.570 158.130 ;
        RECT 70.580 157.930 73.570 158.070 ;
        RECT 68.280 157.730 68.420 157.930 ;
        RECT 68.665 157.885 68.955 157.930 ;
        RECT 72.345 157.885 72.635 157.930 ;
        RECT 73.250 157.870 73.570 157.930 ;
        RECT 73.710 157.870 74.030 158.130 ;
        RECT 74.170 158.070 74.490 158.130 ;
        RECT 77.390 158.070 77.710 158.130 ;
        RECT 77.865 158.070 78.155 158.115 ;
        RECT 74.170 157.930 76.240 158.070 ;
        RECT 74.170 157.870 74.490 157.930 ;
        RECT 60.460 157.590 64.740 157.730 ;
        RECT 66.440 157.590 68.420 157.730 ;
        RECT 53.945 157.390 54.235 157.435 ;
        RECT 55.310 157.390 55.630 157.450 ;
        RECT 55.785 157.390 56.075 157.435 ;
        RECT 53.945 157.250 56.075 157.390 ;
        RECT 53.945 157.205 54.235 157.250 ;
        RECT 55.310 157.190 55.630 157.250 ;
        RECT 55.785 157.205 56.075 157.250 ;
        RECT 56.230 157.390 56.550 157.450 ;
        RECT 60.460 157.390 60.600 157.590 ;
        RECT 66.440 157.450 66.580 157.590 ;
        RECT 70.030 157.530 70.350 157.790 ;
        RECT 71.125 157.730 71.415 157.775 ;
        RECT 74.260 157.730 74.400 157.870 ;
        RECT 71.125 157.590 74.400 157.730 ;
        RECT 71.125 157.545 71.415 157.590 ;
        RECT 75.550 157.530 75.870 157.790 ;
        RECT 76.100 157.730 76.240 157.930 ;
        RECT 77.390 157.930 78.155 158.070 ;
        RECT 77.390 157.870 77.710 157.930 ;
        RECT 77.865 157.885 78.155 157.930 ;
        RECT 78.325 158.070 78.615 158.115 ;
        RECT 79.230 158.070 79.550 158.130 ;
        RECT 78.325 157.930 79.550 158.070 ;
        RECT 78.325 157.885 78.615 157.930 ;
        RECT 79.230 157.870 79.550 157.930 ;
        RECT 79.690 158.070 80.010 158.130 ;
        RECT 80.165 158.070 80.455 158.115 ;
        RECT 80.610 158.070 80.930 158.130 ;
        RECT 81.160 158.115 81.300 158.270 ;
        RECT 82.540 158.115 82.680 158.610 ;
        RECT 83.370 158.410 83.690 158.470 ;
        RECT 84.765 158.410 85.055 158.455 ;
        RECT 83.370 158.270 85.055 158.410 ;
        RECT 83.370 158.210 83.690 158.270 ;
        RECT 84.765 158.225 85.055 158.270 ;
        RECT 85.210 158.210 85.530 158.470 ;
        RECT 79.690 157.930 80.930 158.070 ;
        RECT 79.690 157.870 80.010 157.930 ;
        RECT 80.165 157.885 80.455 157.930 ;
        RECT 80.610 157.870 80.930 157.930 ;
        RECT 81.085 157.885 81.375 158.115 ;
        RECT 82.465 157.885 82.755 158.115 ;
        RECT 82.910 158.070 83.230 158.130 ;
        RECT 84.305 158.070 84.595 158.115 ;
        RECT 82.910 157.930 84.595 158.070 ;
        RECT 82.910 157.870 83.230 157.930 ;
        RECT 84.305 157.885 84.595 157.930 ;
        RECT 85.670 158.070 85.990 158.130 ;
        RECT 89.900 158.115 90.040 158.610 ;
        RECT 90.820 158.455 90.960 158.950 ;
        RECT 91.280 158.950 118.650 159.090 ;
        RECT 91.280 158.795 91.420 158.950 ;
        RECT 118.330 158.890 118.650 158.950 ;
        RECT 118.790 159.090 119.110 159.150 ;
        RECT 120.645 159.090 120.935 159.135 ;
        RECT 118.790 158.950 120.935 159.090 ;
        RECT 118.790 158.890 119.110 158.950 ;
        RECT 120.645 158.905 120.935 158.950 ;
        RECT 122.470 159.090 122.790 159.150 ;
        RECT 127.070 159.090 127.390 159.150 ;
        RECT 122.470 158.950 127.390 159.090 ;
        RECT 122.470 158.890 122.790 158.950 ;
        RECT 127.070 158.890 127.390 158.950 ;
        RECT 91.205 158.565 91.495 158.795 ;
        RECT 92.110 158.750 92.430 158.810 ;
        RECT 93.505 158.750 93.795 158.795 ;
        RECT 92.110 158.610 93.795 158.750 ;
        RECT 92.110 158.550 92.430 158.610 ;
        RECT 93.505 158.565 93.795 158.610 ;
        RECT 93.950 158.750 94.270 158.810 ;
        RECT 95.790 158.750 96.110 158.810 ;
        RECT 93.950 158.610 96.110 158.750 ;
        RECT 93.950 158.550 94.270 158.610 ;
        RECT 95.790 158.550 96.110 158.610 ;
        RECT 100.390 158.750 100.710 158.810 ;
        RECT 103.625 158.750 103.915 158.795 ;
        RECT 100.390 158.610 103.915 158.750 ;
        RECT 100.390 158.550 100.710 158.610 ;
        RECT 103.625 158.565 103.915 158.610 ;
        RECT 104.070 158.750 104.390 158.810 ;
        RECT 129.845 158.750 130.135 158.795 ;
        RECT 104.070 158.610 130.135 158.750 ;
        RECT 104.070 158.550 104.390 158.610 ;
        RECT 129.845 158.565 130.135 158.610 ;
        RECT 90.745 158.225 91.035 158.455 ;
        RECT 93.030 158.410 93.350 158.470 ;
        RECT 104.545 158.410 104.835 158.455 ;
        RECT 93.030 158.270 104.835 158.410 ;
        RECT 93.030 158.210 93.350 158.270 ;
        RECT 88.445 158.070 88.735 158.115 ;
        RECT 85.670 157.930 88.735 158.070 ;
        RECT 85.670 157.870 85.990 157.930 ;
        RECT 88.445 157.885 88.735 157.930 ;
        RECT 88.905 157.885 89.195 158.115 ;
        RECT 89.825 158.070 90.115 158.115 ;
        RECT 91.190 158.070 91.510 158.130 ;
        RECT 89.825 157.930 91.510 158.070 ;
        RECT 89.825 157.885 90.115 157.930 ;
        RECT 76.565 157.730 76.855 157.775 ;
        RECT 76.100 157.590 76.855 157.730 ;
        RECT 76.565 157.545 76.855 157.590 ;
        RECT 78.770 157.730 79.090 157.790 ;
        RECT 88.980 157.730 89.120 157.885 ;
        RECT 91.190 157.870 91.510 157.930 ;
        RECT 92.585 158.070 92.875 158.115 ;
        RECT 93.950 158.070 94.270 158.130 ;
        RECT 92.585 157.930 94.270 158.070 ;
        RECT 92.585 157.885 92.875 157.930 ;
        RECT 93.950 157.870 94.270 157.930 ;
        RECT 94.410 157.870 94.730 158.130 ;
        RECT 95.330 157.870 95.650 158.130 ;
        RECT 98.105 158.070 98.395 158.115 ;
        RECT 99.470 158.070 99.790 158.130 ;
        RECT 98.105 157.930 99.790 158.070 ;
        RECT 98.105 157.885 98.395 157.930 ;
        RECT 99.470 157.870 99.790 157.930 ;
        RECT 100.390 157.870 100.710 158.130 ;
        RECT 101.400 158.115 101.540 158.270 ;
        RECT 104.545 158.225 104.835 158.270 ;
        RECT 106.830 158.410 107.150 158.470 ;
        RECT 118.330 158.410 118.650 158.470 ;
        RECT 123.850 158.410 124.170 158.470 ;
        RECT 106.830 158.270 118.100 158.410 ;
        RECT 106.830 158.210 107.150 158.270 ;
        RECT 101.325 157.885 101.615 158.115 ;
        RECT 101.770 157.870 102.090 158.130 ;
        RECT 102.250 158.070 102.540 158.115 ;
        RECT 102.690 158.070 103.010 158.130 ;
        RECT 102.250 157.930 103.010 158.070 ;
        RECT 102.250 157.885 102.540 157.930 ;
        RECT 102.690 157.870 103.010 157.930 ;
        RECT 112.810 157.870 113.130 158.130 ;
        RECT 114.205 158.070 114.495 158.115 ;
        RECT 114.650 158.070 114.970 158.130 ;
        RECT 114.205 157.930 114.970 158.070 ;
        RECT 117.960 158.070 118.100 158.270 ;
        RECT 118.330 158.270 124.170 158.410 ;
        RECT 118.330 158.210 118.650 158.270 ;
        RECT 123.850 158.210 124.170 158.270 ;
        RECT 124.770 158.070 125.090 158.130 ;
        RECT 117.960 157.930 125.090 158.070 ;
        RECT 129.920 158.070 130.060 158.565 ;
        RECT 132.605 158.070 132.895 158.115 ;
        RECT 129.920 157.930 132.895 158.070 ;
        RECT 114.205 157.885 114.495 157.930 ;
        RECT 114.650 157.870 114.970 157.930 ;
        RECT 124.770 157.870 125.090 157.930 ;
        RECT 132.605 157.885 132.895 157.930 ;
        RECT 133.510 157.870 133.830 158.130 ;
        RECT 99.025 157.730 99.315 157.775 ;
        RECT 103.150 157.730 103.470 157.790 ;
        RECT 78.770 157.590 89.120 157.730 ;
        RECT 89.900 157.590 103.470 157.730 ;
        RECT 78.770 157.530 79.090 157.590 ;
        RECT 56.230 157.250 60.600 157.390 ;
        RECT 56.230 157.190 56.550 157.250 ;
        RECT 66.350 157.190 66.670 157.450 ;
        RECT 68.205 157.390 68.495 157.435 ;
        RECT 73.710 157.390 74.030 157.450 ;
        RECT 68.205 157.250 74.030 157.390 ;
        RECT 68.205 157.205 68.495 157.250 ;
        RECT 73.710 157.190 74.030 157.250 ;
        RECT 76.010 157.390 76.330 157.450 ;
        RECT 79.690 157.390 80.010 157.450 ;
        RECT 76.010 157.250 80.010 157.390 ;
        RECT 76.010 157.190 76.330 157.250 ;
        RECT 79.690 157.190 80.010 157.250 ;
        RECT 81.530 157.390 81.850 157.450 ;
        RECT 82.910 157.390 83.230 157.450 ;
        RECT 81.530 157.250 83.230 157.390 ;
        RECT 81.530 157.190 81.850 157.250 ;
        RECT 82.910 157.190 83.230 157.250 ;
        RECT 83.385 157.390 83.675 157.435 ;
        RECT 87.050 157.390 87.370 157.450 ;
        RECT 83.385 157.250 87.370 157.390 ;
        RECT 83.385 157.205 83.675 157.250 ;
        RECT 87.050 157.190 87.370 157.250 ;
        RECT 87.510 157.390 87.830 157.450 ;
        RECT 89.350 157.390 89.670 157.450 ;
        RECT 89.900 157.390 90.040 157.590 ;
        RECT 99.025 157.545 99.315 157.590 ;
        RECT 103.150 157.530 103.470 157.590 ;
        RECT 117.410 157.730 117.730 157.790 ;
        RECT 123.405 157.730 123.695 157.775 ;
        RECT 117.410 157.590 123.695 157.730 ;
        RECT 117.410 157.530 117.730 157.590 ;
        RECT 123.405 157.545 123.695 157.590 ;
        RECT 87.510 157.250 90.040 157.390 ;
        RECT 87.510 157.190 87.830 157.250 ;
        RECT 89.350 157.190 89.670 157.250 ;
        RECT 90.270 157.190 90.590 157.450 ;
        RECT 91.650 157.390 91.970 157.450 ;
        RECT 96.265 157.390 96.555 157.435 ;
        RECT 91.650 157.250 96.555 157.390 ;
        RECT 91.650 157.190 91.970 157.250 ;
        RECT 96.265 157.205 96.555 157.250 ;
        RECT 98.550 157.390 98.870 157.450 ;
        RECT 105.910 157.390 106.230 157.450 ;
        RECT 112.810 157.390 113.130 157.450 ;
        RECT 98.550 157.250 113.130 157.390 ;
        RECT 98.550 157.190 98.870 157.250 ;
        RECT 105.910 157.190 106.230 157.250 ;
        RECT 112.810 157.190 113.130 157.250 ;
        RECT 115.570 157.390 115.890 157.450 ;
        RECT 120.630 157.390 120.950 157.450 ;
        RECT 115.570 157.250 120.950 157.390 ;
        RECT 115.570 157.190 115.890 157.250 ;
        RECT 120.630 157.190 120.950 157.250 ;
        RECT 121.550 157.390 121.870 157.450 ;
        RECT 133.065 157.390 133.355 157.435 ;
        RECT 121.550 157.250 133.355 157.390 ;
        RECT 121.550 157.190 121.870 157.250 ;
        RECT 133.065 157.205 133.355 157.250 ;
        RECT 23.500 156.570 136.200 157.050 ;
        RECT 51.185 156.370 51.475 156.415 ;
        RECT 52.090 156.370 52.410 156.430 ;
        RECT 53.010 156.370 53.330 156.430 ;
        RECT 51.185 156.230 53.330 156.370 ;
        RECT 51.185 156.185 51.475 156.230 ;
        RECT 52.090 156.170 52.410 156.230 ;
        RECT 53.010 156.170 53.330 156.230 ;
        RECT 54.850 156.370 55.170 156.430 ;
        RECT 55.770 156.370 56.090 156.430 ;
        RECT 57.165 156.370 57.455 156.415 ;
        RECT 54.850 156.230 57.455 156.370 ;
        RECT 54.850 156.170 55.170 156.230 ;
        RECT 55.770 156.170 56.090 156.230 ;
        RECT 57.165 156.185 57.455 156.230 ;
        RECT 64.065 156.370 64.355 156.415 ;
        RECT 66.350 156.370 66.670 156.430 ;
        RECT 68.190 156.370 68.510 156.430 ;
        RECT 64.065 156.230 66.670 156.370 ;
        RECT 64.065 156.185 64.355 156.230 ;
        RECT 66.350 156.170 66.670 156.230 ;
        RECT 66.900 156.230 68.510 156.370 ;
        RECT 56.230 155.830 56.550 156.090 ;
        RECT 64.970 155.830 65.290 156.090 ;
        RECT 66.900 156.030 67.040 156.230 ;
        RECT 68.190 156.170 68.510 156.230 ;
        RECT 70.505 156.370 70.795 156.415 ;
        RECT 71.410 156.370 71.730 156.430 ;
        RECT 70.505 156.230 71.730 156.370 ;
        RECT 70.505 156.185 70.795 156.230 ;
        RECT 71.410 156.170 71.730 156.230 ;
        RECT 72.330 156.170 72.650 156.430 ;
        RECT 78.770 156.170 79.090 156.430 ;
        RECT 79.230 156.170 79.550 156.430 ;
        RECT 80.625 156.370 80.915 156.415 ;
        RECT 81.070 156.370 81.390 156.430 ;
        RECT 80.625 156.230 81.390 156.370 ;
        RECT 80.625 156.185 80.915 156.230 ;
        RECT 81.070 156.170 81.390 156.230 ;
        RECT 81.545 156.370 81.835 156.415 ;
        RECT 81.990 156.370 82.310 156.430 ;
        RECT 81.545 156.230 82.310 156.370 ;
        RECT 81.545 156.185 81.835 156.230 ;
        RECT 81.990 156.170 82.310 156.230 ;
        RECT 84.290 156.170 84.610 156.430 ;
        RECT 88.445 156.370 88.735 156.415 ;
        RECT 90.270 156.370 90.590 156.430 ;
        RECT 88.445 156.230 90.590 156.370 ;
        RECT 88.445 156.185 88.735 156.230 ;
        RECT 90.270 156.170 90.590 156.230 ;
        RECT 93.965 156.370 94.255 156.415 ;
        RECT 94.870 156.370 95.190 156.430 ;
        RECT 93.965 156.230 95.190 156.370 ;
        RECT 93.965 156.185 94.255 156.230 ;
        RECT 72.420 156.030 72.560 156.170 ;
        RECT 66.210 155.890 67.040 156.030 ;
        RECT 67.820 155.890 72.560 156.030 ;
        RECT 74.170 156.030 74.490 156.090 ;
        RECT 79.320 156.030 79.460 156.170 ;
        RECT 85.670 156.030 85.990 156.090 ;
        RECT 94.040 156.030 94.180 156.185 ;
        RECT 94.870 156.170 95.190 156.230 ;
        RECT 101.770 156.170 102.090 156.430 ;
        RECT 107.765 156.370 108.055 156.415 ;
        RECT 110.050 156.370 110.370 156.430 ;
        RECT 114.190 156.370 114.510 156.430 ;
        RECT 127.990 156.370 128.310 156.430 ;
        RECT 107.765 156.230 114.510 156.370 ;
        RECT 107.765 156.185 108.055 156.230 ;
        RECT 110.050 156.170 110.370 156.230 ;
        RECT 114.190 156.170 114.510 156.230 ;
        RECT 126.240 156.230 128.310 156.370 ;
        RECT 74.170 155.890 74.860 156.030 ;
        RECT 52.105 155.505 52.395 155.735 ;
        RECT 52.180 155.350 52.320 155.505 ;
        RECT 53.010 155.490 53.330 155.750 ;
        RECT 53.945 155.690 54.235 155.735 ;
        RECT 54.390 155.690 54.710 155.750 ;
        RECT 53.945 155.550 54.710 155.690 ;
        RECT 53.945 155.505 54.235 155.550 ;
        RECT 54.390 155.490 54.710 155.550 ;
        RECT 54.850 155.490 55.170 155.750 ;
        RECT 58.070 155.490 58.390 155.750 ;
        RECT 59.910 155.490 60.230 155.750 ;
        RECT 61.305 155.690 61.595 155.735 ;
        RECT 60.460 155.550 61.595 155.690 ;
        RECT 58.530 155.350 58.850 155.410 ;
        RECT 52.180 155.210 58.850 155.350 ;
        RECT 58.530 155.150 58.850 155.210 ;
        RECT 58.990 155.350 59.310 155.410 ;
        RECT 60.460 155.350 60.600 155.550 ;
        RECT 61.305 155.505 61.595 155.550 ;
        RECT 62.210 155.690 62.530 155.750 ;
        RECT 63.145 155.690 63.435 155.735 ;
        RECT 62.210 155.550 63.435 155.690 ;
        RECT 62.210 155.490 62.530 155.550 ;
        RECT 63.145 155.505 63.435 155.550 ;
        RECT 58.990 155.210 60.600 155.350 ;
        RECT 60.830 155.350 61.150 155.410 ;
        RECT 66.210 155.350 66.350 155.890 ;
        RECT 67.820 155.750 67.960 155.890 ;
        RECT 74.170 155.830 74.490 155.890 ;
        RECT 66.825 155.505 67.115 155.735 ;
        RECT 60.830 155.210 66.350 155.350 ;
        RECT 66.900 155.350 67.040 155.505 ;
        RECT 67.730 155.490 68.050 155.750 ;
        RECT 68.190 155.490 68.510 155.750 ;
        RECT 69.570 155.490 69.890 155.750 ;
        RECT 71.870 155.490 72.190 155.750 ;
        RECT 72.330 155.490 72.650 155.750 ;
        RECT 73.250 155.690 73.570 155.750 ;
        RECT 74.720 155.735 74.860 155.890 ;
        RECT 75.640 155.890 79.460 156.030 ;
        RECT 82.540 155.890 85.990 156.030 ;
        RECT 75.640 155.735 75.780 155.890 ;
        RECT 73.725 155.690 74.015 155.735 ;
        RECT 73.250 155.550 74.015 155.690 ;
        RECT 73.250 155.490 73.570 155.550 ;
        RECT 73.725 155.505 74.015 155.550 ;
        RECT 74.645 155.505 74.935 155.735 ;
        RECT 75.565 155.505 75.855 155.735 ;
        RECT 76.470 155.490 76.790 155.750 ;
        RECT 77.865 155.690 78.155 155.735 ;
        RECT 79.230 155.690 79.550 155.750 ;
        RECT 77.865 155.550 79.550 155.690 ;
        RECT 77.865 155.505 78.155 155.550 ;
        RECT 70.950 155.350 71.270 155.410 ;
        RECT 66.900 155.210 71.270 155.350 ;
        RECT 58.990 155.150 59.310 155.210 ;
        RECT 60.830 155.150 61.150 155.210 ;
        RECT 53.010 155.010 53.330 155.070 ;
        RECT 66.900 155.010 67.040 155.210 ;
        RECT 70.950 155.150 71.270 155.210 ;
        RECT 71.425 155.350 71.715 155.395 ;
        RECT 72.790 155.350 73.110 155.410 ;
        RECT 71.425 155.210 73.110 155.350 ;
        RECT 71.425 155.165 71.715 155.210 ;
        RECT 72.790 155.150 73.110 155.210 ;
        RECT 74.185 155.350 74.475 155.395 ;
        RECT 77.390 155.350 77.710 155.410 ;
        RECT 74.185 155.210 77.710 155.350 ;
        RECT 74.185 155.165 74.475 155.210 ;
        RECT 77.390 155.150 77.710 155.210 ;
        RECT 77.940 155.010 78.080 155.505 ;
        RECT 79.230 155.490 79.550 155.550 ;
        RECT 80.150 155.690 80.470 155.750 ;
        RECT 81.085 155.690 81.375 155.735 ;
        RECT 80.150 155.550 81.375 155.690 ;
        RECT 80.150 155.490 80.470 155.550 ;
        RECT 81.085 155.505 81.375 155.550 ;
        RECT 81.530 155.690 81.850 155.750 ;
        RECT 82.540 155.735 82.680 155.890 ;
        RECT 85.670 155.830 85.990 155.890 ;
        RECT 86.220 155.890 94.180 156.030 ;
        RECT 95.330 156.030 95.650 156.090 ;
        RECT 112.810 156.030 113.130 156.090 ;
        RECT 114.665 156.030 114.955 156.075 ;
        RECT 95.330 155.890 101.080 156.030 ;
        RECT 82.465 155.690 82.755 155.735 ;
        RECT 81.530 155.550 82.755 155.690 ;
        RECT 81.530 155.490 81.850 155.550 ;
        RECT 82.465 155.505 82.755 155.550 ;
        RECT 83.370 155.490 83.690 155.750 ;
        RECT 85.210 155.490 85.530 155.750 ;
        RECT 86.220 155.735 86.360 155.890 ;
        RECT 95.330 155.830 95.650 155.890 ;
        RECT 86.145 155.505 86.435 155.735 ;
        RECT 87.050 155.490 87.370 155.750 ;
        RECT 87.970 155.490 88.290 155.750 ;
        RECT 89.810 155.490 90.130 155.750 ;
        RECT 100.405 155.505 100.695 155.735 ;
        RECT 100.940 155.690 101.080 155.890 ;
        RECT 112.810 155.890 114.955 156.030 ;
        RECT 112.810 155.830 113.130 155.890 ;
        RECT 114.665 155.845 114.955 155.890 ;
        RECT 115.585 155.845 115.875 156.075 ;
        RECT 117.425 156.030 117.715 156.075 ;
        RECT 117.870 156.030 118.190 156.090 ;
        RECT 126.240 156.075 126.380 156.230 ;
        RECT 127.990 156.170 128.310 156.230 ;
        RECT 129.385 156.370 129.675 156.415 ;
        RECT 132.130 156.370 132.450 156.430 ;
        RECT 129.385 156.230 132.450 156.370 ;
        RECT 129.385 156.185 129.675 156.230 ;
        RECT 132.130 156.170 132.450 156.230 ;
        RECT 133.050 156.370 133.370 156.430 ;
        RECT 133.985 156.370 134.275 156.415 ;
        RECT 133.050 156.230 134.275 156.370 ;
        RECT 133.050 156.170 133.370 156.230 ;
        RECT 133.985 156.185 134.275 156.230 ;
        RECT 117.425 155.890 118.190 156.030 ;
        RECT 117.425 155.845 117.715 155.890 ;
        RECT 101.325 155.690 101.615 155.735 ;
        RECT 100.940 155.550 101.615 155.690 ;
        RECT 101.325 155.505 101.615 155.550 ;
        RECT 78.310 155.350 78.630 155.410 ;
        RECT 86.605 155.350 86.895 155.395 ;
        RECT 88.905 155.350 89.195 155.395 ;
        RECT 78.310 155.210 86.895 155.350 ;
        RECT 78.310 155.150 78.630 155.210 ;
        RECT 86.605 155.165 86.895 155.210 ;
        RECT 87.140 155.210 89.195 155.350 ;
        RECT 53.010 154.870 67.040 155.010 ;
        RECT 71.500 154.870 78.080 155.010 ;
        RECT 53.010 154.810 53.330 154.870 ;
        RECT 21.730 154.670 22.050 154.730 ;
        RECT 24.965 154.670 25.255 154.715 ;
        RECT 21.730 154.530 25.255 154.670 ;
        RECT 21.730 154.470 22.050 154.530 ;
        RECT 24.965 154.485 25.255 154.530 ;
        RECT 54.390 154.670 54.710 154.730 ;
        RECT 59.005 154.670 59.295 154.715 ;
        RECT 62.210 154.670 62.530 154.730 ;
        RECT 63.220 154.715 63.360 154.870 ;
        RECT 54.390 154.530 62.530 154.670 ;
        RECT 54.390 154.470 54.710 154.530 ;
        RECT 59.005 154.485 59.295 154.530 ;
        RECT 62.210 154.470 62.530 154.530 ;
        RECT 63.145 154.485 63.435 154.715 ;
        RECT 63.590 154.670 63.910 154.730 ;
        RECT 71.500 154.670 71.640 154.870 ;
        RECT 63.590 154.530 71.640 154.670 ;
        RECT 71.870 154.670 72.190 154.730 ;
        RECT 72.790 154.670 73.110 154.730 ;
        RECT 71.870 154.530 73.110 154.670 ;
        RECT 63.590 154.470 63.910 154.530 ;
        RECT 71.870 154.470 72.190 154.530 ;
        RECT 72.790 154.470 73.110 154.530 ;
        RECT 73.265 154.670 73.555 154.715 ;
        RECT 74.170 154.670 74.490 154.730 ;
        RECT 73.265 154.530 74.490 154.670 ;
        RECT 73.265 154.485 73.555 154.530 ;
        RECT 74.170 154.470 74.490 154.530 ;
        RECT 74.630 154.670 74.950 154.730 ;
        RECT 78.770 154.670 79.090 154.730 ;
        RECT 74.630 154.530 79.090 154.670 ;
        RECT 74.630 154.470 74.950 154.530 ;
        RECT 78.770 154.470 79.090 154.530 ;
        RECT 80.610 154.670 80.930 154.730 ;
        RECT 82.465 154.670 82.755 154.715 ;
        RECT 80.610 154.530 82.755 154.670 ;
        RECT 80.610 154.470 80.930 154.530 ;
        RECT 82.465 154.485 82.755 154.530 ;
        RECT 82.910 154.670 83.230 154.730 ;
        RECT 86.590 154.670 86.910 154.730 ;
        RECT 87.140 154.670 87.280 155.210 ;
        RECT 88.905 155.165 89.195 155.210 ;
        RECT 89.365 155.010 89.655 155.055 ;
        RECT 100.480 155.010 100.620 155.505 ;
        RECT 103.150 155.490 103.470 155.750 ;
        RECT 114.190 155.490 114.510 155.750 ;
        RECT 103.610 155.150 103.930 155.410 ;
        RECT 110.510 155.350 110.830 155.410 ;
        RECT 115.660 155.350 115.800 155.845 ;
        RECT 117.870 155.830 118.190 155.890 ;
        RECT 126.165 155.845 126.455 156.075 ;
        RECT 127.070 156.030 127.390 156.090 ;
        RECT 134.890 156.030 135.210 156.090 ;
        RECT 127.070 155.890 130.980 156.030 ;
        RECT 127.070 155.830 127.390 155.890 ;
        RECT 121.090 155.690 121.410 155.750 ;
        RECT 128.005 155.690 128.295 155.735 ;
        RECT 121.090 155.550 128.295 155.690 ;
        RECT 121.090 155.490 121.410 155.550 ;
        RECT 128.005 155.505 128.295 155.550 ;
        RECT 129.830 155.490 130.150 155.750 ;
        RECT 130.840 155.735 130.980 155.890 ;
        RECT 131.760 155.890 135.210 156.030 ;
        RECT 131.760 155.735 131.900 155.890 ;
        RECT 134.890 155.830 135.210 155.890 ;
        RECT 130.765 155.505 131.055 155.735 ;
        RECT 131.685 155.505 131.975 155.735 ;
        RECT 133.065 155.505 133.355 155.735 ;
        RECT 110.510 155.210 115.800 155.350 ;
        RECT 127.085 155.350 127.375 155.395 ;
        RECT 128.450 155.350 128.770 155.410 ;
        RECT 127.085 155.210 128.770 155.350 ;
        RECT 110.510 155.150 110.830 155.210 ;
        RECT 127.085 155.165 127.375 155.210 ;
        RECT 128.450 155.150 128.770 155.210 ;
        RECT 114.650 155.010 114.970 155.070 ;
        RECT 133.140 155.010 133.280 155.505 ;
        RECT 89.365 154.870 93.720 155.010 ;
        RECT 100.480 154.870 114.970 155.010 ;
        RECT 89.365 154.825 89.655 154.870 ;
        RECT 82.910 154.530 87.280 154.670 ;
        RECT 88.890 154.670 89.210 154.730 ;
        RECT 90.745 154.670 91.035 154.715 ;
        RECT 88.890 154.530 91.035 154.670 ;
        RECT 93.580 154.670 93.720 154.870 ;
        RECT 114.650 154.810 114.970 154.870 ;
        RECT 115.200 154.870 133.280 155.010 ;
        RECT 100.850 154.670 101.170 154.730 ;
        RECT 93.580 154.530 101.170 154.670 ;
        RECT 82.910 154.470 83.230 154.530 ;
        RECT 86.590 154.470 86.910 154.530 ;
        RECT 88.890 154.470 89.210 154.530 ;
        RECT 90.745 154.485 91.035 154.530 ;
        RECT 100.850 154.470 101.170 154.530 ;
        RECT 104.990 154.670 105.310 154.730 ;
        RECT 115.200 154.670 115.340 154.870 ;
        RECT 104.990 154.530 115.340 154.670 ;
        RECT 115.585 154.670 115.875 154.715 ;
        RECT 116.030 154.670 116.350 154.730 ;
        RECT 115.585 154.530 116.350 154.670 ;
        RECT 104.990 154.470 105.310 154.530 ;
        RECT 115.585 154.485 115.875 154.530 ;
        RECT 116.030 154.470 116.350 154.530 ;
        RECT 116.490 154.470 116.810 154.730 ;
        RECT 23.500 153.850 136.200 154.330 ;
        RECT 38.765 153.650 39.055 153.695 ;
        RECT 41.050 153.650 41.370 153.710 ;
        RECT 38.765 153.510 41.370 153.650 ;
        RECT 38.765 153.465 39.055 153.510 ;
        RECT 41.050 153.450 41.370 153.510 ;
        RECT 46.110 153.650 46.430 153.710 ;
        RECT 48.425 153.650 48.715 153.695 ;
        RECT 46.110 153.510 48.715 153.650 ;
        RECT 46.110 153.450 46.430 153.510 ;
        RECT 48.425 153.465 48.715 153.510 ;
        RECT 54.405 153.650 54.695 153.695 ;
        RECT 54.850 153.650 55.170 153.710 ;
        RECT 54.405 153.510 55.170 153.650 ;
        RECT 54.405 153.465 54.695 153.510 ;
        RECT 54.850 153.450 55.170 153.510 ;
        RECT 55.310 153.450 55.630 153.710 ;
        RECT 58.530 153.650 58.850 153.710 ;
        RECT 72.790 153.650 73.110 153.710 ;
        RECT 87.050 153.650 87.370 153.710 ;
        RECT 93.965 153.650 94.255 153.695 ;
        RECT 100.390 153.650 100.710 153.710 ;
        RECT 58.530 153.510 65.660 153.650 ;
        RECT 58.530 153.450 58.850 153.510 ;
        RECT 41.985 153.310 42.275 153.355 ;
        RECT 59.910 153.310 60.230 153.370 ;
        RECT 41.985 153.170 60.230 153.310 ;
        RECT 41.985 153.125 42.275 153.170 ;
        RECT 59.910 153.110 60.230 153.170 ;
        RECT 61.750 153.110 62.070 153.370 ;
        RECT 64.525 153.125 64.815 153.355 ;
        RECT 65.520 153.310 65.660 153.510 ;
        RECT 72.790 153.510 83.600 153.650 ;
        RECT 72.790 153.450 73.110 153.510 ;
        RECT 76.930 153.310 77.250 153.370 ;
        RECT 65.520 153.170 77.250 153.310 ;
        RECT 52.090 152.770 52.410 153.030 ;
        RECT 57.150 152.970 57.470 153.030 ;
        RECT 52.640 152.830 57.470 152.970 ;
        RECT 60.000 152.970 60.140 153.110 ;
        RECT 64.600 152.970 64.740 153.125 ;
        RECT 76.930 153.110 77.250 153.170 ;
        RECT 77.405 153.310 77.695 153.355 ;
        RECT 82.910 153.310 83.230 153.370 ;
        RECT 83.460 153.355 83.600 153.510 ;
        RECT 87.050 153.510 100.710 153.650 ;
        RECT 87.050 153.450 87.370 153.510 ;
        RECT 93.965 153.465 94.255 153.510 ;
        RECT 100.390 153.450 100.710 153.510 ;
        RECT 100.850 153.650 101.170 153.710 ;
        RECT 104.070 153.650 104.390 153.710 ;
        RECT 100.850 153.510 104.390 153.650 ;
        RECT 100.850 153.450 101.170 153.510 ;
        RECT 104.070 153.450 104.390 153.510 ;
        RECT 112.365 153.650 112.655 153.695 ;
        RECT 114.190 153.650 114.510 153.710 ;
        RECT 112.365 153.510 114.510 153.650 ;
        RECT 112.365 153.465 112.655 153.510 ;
        RECT 114.190 153.450 114.510 153.510 ;
        RECT 134.430 153.450 134.750 153.710 ;
        RECT 77.405 153.170 83.230 153.310 ;
        RECT 77.405 153.125 77.695 153.170 ;
        RECT 82.910 153.110 83.230 153.170 ;
        RECT 83.385 153.125 83.675 153.355 ;
        RECT 107.290 153.310 107.610 153.370 ;
        RECT 115.110 153.310 115.430 153.370 ;
        RECT 107.290 153.170 115.430 153.310 ;
        RECT 107.290 153.110 107.610 153.170 ;
        RECT 115.110 153.110 115.430 153.170 ;
        RECT 132.590 153.110 132.910 153.370 ;
        RECT 67.730 152.970 68.050 153.030 ;
        RECT 114.650 152.970 114.970 153.030 ;
        RECT 117.410 152.970 117.730 153.030 ;
        RECT 60.000 152.830 63.820 152.970 ;
        RECT 64.600 152.830 68.050 152.970 ;
        RECT 37.370 152.630 37.690 152.690 ;
        RECT 37.845 152.630 38.135 152.675 ;
        RECT 37.370 152.490 38.135 152.630 ;
        RECT 37.370 152.430 37.690 152.490 ;
        RECT 37.845 152.445 38.135 152.490 ;
        RECT 40.590 152.630 40.910 152.690 ;
        RECT 41.065 152.630 41.355 152.675 ;
        RECT 40.590 152.490 41.355 152.630 ;
        RECT 40.590 152.430 40.910 152.490 ;
        RECT 41.065 152.445 41.355 152.490 ;
        RECT 44.270 152.430 44.590 152.690 ;
        RECT 47.030 152.630 47.350 152.690 ;
        RECT 52.640 152.675 52.780 152.830 ;
        RECT 57.150 152.770 57.470 152.830 ;
        RECT 47.505 152.630 47.795 152.675 ;
        RECT 47.030 152.490 47.795 152.630 ;
        RECT 47.030 152.430 47.350 152.490 ;
        RECT 47.505 152.445 47.795 152.490 ;
        RECT 52.565 152.445 52.855 152.675 ;
        RECT 45.280 152.150 49.100 152.290 ;
        RECT 45.280 151.995 45.420 152.150 ;
        RECT 45.205 151.765 45.495 151.995 ;
        RECT 48.960 151.950 49.100 152.150 ;
        RECT 52.640 151.950 52.780 152.445 ;
        RECT 54.390 152.430 54.710 152.690 ;
        RECT 56.690 152.630 57.010 152.690 ;
        RECT 63.680 152.675 63.820 152.830 ;
        RECT 67.730 152.770 68.050 152.830 ;
        RECT 71.960 152.830 113.500 152.970 ;
        RECT 57.625 152.630 57.915 152.675 ;
        RECT 60.845 152.630 61.135 152.675 ;
        RECT 56.690 152.490 57.915 152.630 ;
        RECT 56.690 152.430 57.010 152.490 ;
        RECT 57.625 152.445 57.915 152.490 ;
        RECT 60.460 152.490 61.135 152.630 ;
        RECT 53.470 152.290 53.790 152.350 ;
        RECT 56.245 152.290 56.535 152.335 ;
        RECT 53.470 152.150 56.535 152.290 ;
        RECT 53.470 152.090 53.790 152.150 ;
        RECT 56.245 152.105 56.535 152.150 ;
        RECT 57.165 152.290 57.455 152.335 ;
        RECT 58.070 152.290 58.390 152.350 ;
        RECT 57.165 152.150 58.390 152.290 ;
        RECT 57.165 152.105 57.455 152.150 ;
        RECT 58.070 152.090 58.390 152.150 ;
        RECT 60.460 152.010 60.600 152.490 ;
        RECT 60.845 152.445 61.135 152.490 ;
        RECT 63.605 152.445 63.895 152.675 ;
        RECT 65.430 152.430 65.750 152.690 ;
        RECT 68.190 152.430 68.510 152.690 ;
        RECT 71.960 152.675 72.100 152.830 ;
        RECT 71.885 152.445 72.175 152.675 ;
        RECT 72.345 152.630 72.635 152.675 ;
        RECT 72.790 152.630 73.110 152.690 ;
        RECT 72.345 152.490 73.110 152.630 ;
        RECT 72.345 152.445 72.635 152.490 ;
        RECT 72.790 152.430 73.110 152.490 ;
        RECT 73.710 152.430 74.030 152.690 ;
        RECT 76.470 152.430 76.790 152.690 ;
        RECT 77.865 152.445 78.155 152.675 ;
        RECT 78.770 152.630 79.090 152.690 ;
        RECT 79.245 152.630 79.535 152.675 ;
        RECT 78.770 152.490 79.535 152.630 ;
        RECT 70.490 152.090 70.810 152.350 ;
        RECT 77.940 152.290 78.080 152.445 ;
        RECT 78.770 152.430 79.090 152.490 ;
        RECT 79.245 152.445 79.535 152.490 ;
        RECT 79.690 152.630 80.010 152.690 ;
        RECT 80.165 152.630 80.455 152.675 ;
        RECT 79.690 152.490 80.455 152.630 ;
        RECT 79.690 152.430 80.010 152.490 ;
        RECT 80.165 152.445 80.455 152.490 ;
        RECT 82.450 152.430 82.770 152.690 ;
        RECT 83.845 152.445 84.135 152.675 ;
        RECT 84.765 152.445 85.055 152.675 ;
        RECT 83.370 152.290 83.690 152.350 ;
        RECT 77.940 152.150 83.690 152.290 ;
        RECT 83.370 152.090 83.690 152.150 ;
        RECT 48.960 151.810 52.780 151.950 ;
        RECT 60.370 151.750 60.690 152.010 ;
        RECT 66.350 151.750 66.670 152.010 ;
        RECT 67.730 151.750 68.050 152.010 ;
        RECT 69.110 151.750 69.430 152.010 ;
        RECT 73.250 151.750 73.570 152.010 ;
        RECT 74.630 151.750 74.950 152.010 ;
        RECT 78.770 151.750 79.090 152.010 ;
        RECT 79.705 151.950 79.995 151.995 ;
        RECT 81.070 151.950 81.390 152.010 ;
        RECT 79.705 151.810 81.390 151.950 ;
        RECT 79.705 151.765 79.995 151.810 ;
        RECT 81.070 151.750 81.390 151.810 ;
        RECT 81.530 151.750 81.850 152.010 ;
        RECT 83.920 151.950 84.060 152.445 ;
        RECT 84.840 152.290 84.980 152.445 ;
        RECT 87.050 152.430 87.370 152.690 ;
        RECT 88.430 152.430 88.750 152.690 ;
        RECT 89.350 152.630 89.670 152.690 ;
        RECT 90.745 152.630 91.035 152.675 ;
        RECT 89.350 152.490 91.035 152.630 ;
        RECT 89.350 152.430 89.670 152.490 ;
        RECT 90.745 152.445 91.035 152.490 ;
        RECT 100.405 152.630 100.695 152.675 ;
        RECT 107.290 152.630 107.610 152.690 ;
        RECT 100.405 152.490 107.610 152.630 ;
        RECT 100.405 152.445 100.695 152.490 ;
        RECT 107.290 152.430 107.610 152.490 ;
        RECT 110.050 152.430 110.370 152.690 ;
        RECT 110.510 152.430 110.830 152.690 ;
        RECT 112.810 152.430 113.130 152.690 ;
        RECT 113.360 152.630 113.500 152.830 ;
        RECT 114.650 152.830 117.730 152.970 ;
        RECT 114.650 152.770 114.970 152.830 ;
        RECT 117.410 152.770 117.730 152.830 ;
        RECT 117.870 152.970 118.190 153.030 ;
        RECT 127.085 152.970 127.375 153.015 ;
        RECT 117.870 152.830 127.375 152.970 ;
        RECT 117.870 152.770 118.190 152.830 ;
        RECT 127.085 152.785 127.375 152.830 ;
        RECT 128.465 152.970 128.755 153.015 ;
        RECT 129.830 152.970 130.150 153.030 ;
        RECT 128.465 152.830 130.150 152.970 ;
        RECT 128.465 152.785 128.755 152.830 ;
        RECT 129.830 152.770 130.150 152.830 ;
        RECT 130.290 152.970 130.610 153.030 ;
        RECT 133.065 152.970 133.355 153.015 ;
        RECT 130.290 152.830 133.355 152.970 ;
        RECT 130.290 152.770 130.610 152.830 ;
        RECT 133.065 152.785 133.355 152.830 ;
        RECT 115.585 152.630 115.875 152.675 ;
        RECT 119.250 152.630 119.570 152.690 ;
        RECT 113.360 152.490 114.880 152.630 ;
        RECT 89.825 152.290 90.115 152.335 ;
        RECT 96.710 152.290 97.030 152.350 ;
        RECT 84.840 152.150 97.030 152.290 ;
        RECT 89.825 152.105 90.115 152.150 ;
        RECT 96.710 152.090 97.030 152.150 ;
        RECT 101.325 152.290 101.615 152.335 ;
        RECT 103.610 152.290 103.930 152.350 ;
        RECT 101.325 152.150 103.930 152.290 ;
        RECT 101.325 152.105 101.615 152.150 ;
        RECT 101.400 151.950 101.540 152.105 ;
        RECT 103.610 152.090 103.930 152.150 ;
        RECT 104.070 152.290 104.390 152.350 ;
        RECT 114.205 152.290 114.495 152.335 ;
        RECT 104.070 152.150 114.495 152.290 ;
        RECT 114.740 152.290 114.880 152.490 ;
        RECT 115.585 152.490 119.570 152.630 ;
        RECT 115.585 152.445 115.875 152.490 ;
        RECT 119.250 152.430 119.570 152.490 ;
        RECT 132.130 152.430 132.450 152.690 ;
        RECT 133.525 152.445 133.815 152.675 ;
        RECT 114.740 152.150 116.260 152.290 ;
        RECT 104.070 152.090 104.390 152.150 ;
        RECT 114.205 152.105 114.495 152.150 ;
        RECT 83.920 151.810 101.540 151.950 ;
        RECT 114.665 151.950 114.955 151.995 ;
        RECT 115.570 151.950 115.890 152.010 ;
        RECT 114.665 151.810 115.890 151.950 ;
        RECT 116.120 151.950 116.260 152.150 ;
        RECT 116.490 152.090 116.810 152.350 ;
        RECT 126.150 152.090 126.470 152.350 ;
        RECT 126.610 152.290 126.930 152.350 ;
        RECT 133.600 152.290 133.740 152.445 ;
        RECT 126.610 152.150 133.740 152.290 ;
        RECT 126.610 152.090 126.930 152.150 ;
        RECT 129.370 151.950 129.690 152.010 ;
        RECT 116.120 151.810 129.690 151.950 ;
        RECT 114.665 151.765 114.955 151.810 ;
        RECT 115.570 151.750 115.890 151.810 ;
        RECT 129.370 151.750 129.690 151.810 ;
        RECT 23.500 151.130 136.200 151.610 ;
        RECT 73.710 150.930 74.030 150.990 ;
        RECT 101.770 150.930 102.090 150.990 ;
        RECT 73.710 150.790 102.090 150.930 ;
        RECT 73.710 150.730 74.030 150.790 ;
        RECT 101.770 150.730 102.090 150.790 ;
        RECT 76.470 150.590 76.790 150.650 ;
        RECT 91.650 150.590 91.970 150.650 ;
        RECT 76.470 150.450 91.970 150.590 ;
        RECT 76.470 150.390 76.790 150.450 ;
        RECT 91.650 150.390 91.970 150.450 ;
        RECT 72.330 150.250 72.650 150.310 ;
        RECT 116.490 150.250 116.810 150.310 ;
        RECT 72.330 150.110 116.810 150.250 ;
        RECT 72.330 150.050 72.650 150.110 ;
        RECT 116.490 150.050 116.810 150.110 ;
        RECT 68.190 149.910 68.510 149.970 ;
        RECT 92.570 149.910 92.890 149.970 ;
        RECT 68.190 149.770 92.890 149.910 ;
        RECT 68.190 149.710 68.510 149.770 ;
        RECT 92.570 149.710 92.890 149.770 ;
        RECT 65.430 149.570 65.750 149.630 ;
        RECT 101.310 149.570 101.630 149.630 ;
        RECT 65.430 149.430 101.630 149.570 ;
        RECT 65.430 149.370 65.750 149.430 ;
        RECT 101.310 149.370 101.630 149.430 ;
        RECT 83.370 149.230 83.690 149.290 ;
        RECT 116.030 149.230 116.350 149.290 ;
        RECT 83.370 149.090 116.350 149.230 ;
        RECT 83.370 149.030 83.690 149.090 ;
        RECT 116.030 149.030 116.350 149.090 ;
        RECT 58.070 148.890 58.390 148.950 ;
        RECT 81.530 148.890 81.850 148.950 ;
        RECT 92.110 148.890 92.430 148.950 ;
        RECT 58.070 148.750 80.150 148.890 ;
        RECT 58.070 148.690 58.390 148.750 ;
        RECT 80.010 148.550 80.150 148.750 ;
        RECT 81.530 148.750 92.430 148.890 ;
        RECT 81.530 148.690 81.850 148.750 ;
        RECT 92.110 148.690 92.430 148.750 ;
        RECT 88.430 148.550 88.750 148.610 ;
        RECT 95.330 148.550 95.650 148.610 ;
        RECT 80.010 148.410 95.650 148.550 ;
        RECT 88.430 148.350 88.750 148.410 ;
        RECT 95.330 148.350 95.650 148.410 ;
        RECT 74.170 147.190 74.490 147.250 ;
        RECT 111.430 147.190 111.750 147.250 ;
        RECT 74.170 147.050 111.750 147.190 ;
        RECT 74.170 146.990 74.490 147.050 ;
        RECT 111.430 146.990 111.750 147.050 ;
        RECT 73.250 146.850 73.570 146.910 ;
        RECT 104.990 146.850 105.310 146.910 ;
        RECT 73.250 146.710 105.310 146.850 ;
        RECT 73.250 146.650 73.570 146.710 ;
        RECT 104.990 146.650 105.310 146.710 ;
        RECT 78.770 146.510 79.090 146.570 ;
        RECT 98.550 146.510 98.870 146.570 ;
        RECT 78.770 146.370 98.870 146.510 ;
        RECT 78.770 146.310 79.090 146.370 ;
        RECT 98.550 146.310 98.870 146.370 ;
        RECT 69.110 146.170 69.430 146.230 ;
        RECT 108.210 146.170 108.530 146.230 ;
        RECT 69.110 146.030 108.530 146.170 ;
        RECT 69.110 145.970 69.430 146.030 ;
        RECT 108.210 145.970 108.530 146.030 ;
        RECT 74.630 145.830 74.950 145.890 ;
        RECT 101.770 145.830 102.090 145.890 ;
        RECT 74.630 145.690 102.090 145.830 ;
        RECT 74.630 145.630 74.950 145.690 ;
        RECT 101.770 145.630 102.090 145.690 ;
        RECT 82.910 145.490 83.230 145.550 ;
        RECT 95.330 145.490 95.650 145.550 ;
        RECT 82.910 145.350 95.650 145.490 ;
        RECT 82.910 145.290 83.230 145.350 ;
        RECT 95.330 145.290 95.650 145.350 ;
        RECT 67.730 143.790 68.050 143.850 ;
        RECT 127.530 143.790 127.850 143.850 ;
        RECT 67.730 143.650 127.850 143.790 ;
        RECT 67.730 143.590 68.050 143.650 ;
        RECT 127.530 143.590 127.850 143.650 ;
        RECT 70.490 141.070 70.810 141.130 ;
        RECT 114.650 141.070 114.970 141.130 ;
        RECT 70.490 140.930 114.970 141.070 ;
        RECT 70.490 140.870 70.810 140.930 ;
        RECT 114.650 140.870 114.970 140.930 ;
        RECT 77.445 70.840 78.085 70.845 ;
        RECT 50.550 70.835 78.085 70.840 ;
        RECT 81.075 70.840 81.805 70.845 ;
        RECT 81.075 70.835 110.655 70.840 ;
        RECT 50.550 70.300 110.655 70.835 ;
        RECT 50.245 69.600 110.655 70.300 ;
        RECT 50.245 69.435 75.895 69.600 ;
        RECT 76.885 69.435 110.655 69.600 ;
        RECT 46.890 68.900 47.480 68.950 ;
        RECT 48.710 68.900 49.300 68.950 ;
        RECT 46.890 66.945 49.300 68.900 ;
        RECT 50.245 68.670 50.705 69.435 ;
        RECT 51.205 68.920 51.520 69.210 ;
        RECT 51.020 68.670 51.250 68.715 ;
        RECT 50.245 68.000 51.250 68.670 ;
        RECT 46.890 66.845 47.480 66.945 ;
        RECT 48.710 66.845 49.300 66.945 ;
        RECT 46.890 65.940 47.480 66.265 ;
        RECT 48.710 65.960 49.300 66.265 ;
        RECT 46.870 60.920 47.495 65.940 ;
        RECT 48.685 60.940 49.310 65.960 ;
        RECT 50.655 62.795 51.250 68.000 ;
        RECT 51.020 62.715 51.250 62.795 ;
        RECT 51.460 68.655 51.690 68.715 ;
        RECT 53.355 68.670 53.945 68.965 ;
        RECT 51.950 68.655 53.945 68.670 ;
        RECT 51.460 66.885 53.945 68.655 ;
        RECT 51.460 65.275 52.365 66.885 ;
        RECT 53.355 66.860 53.945 66.885 ;
        RECT 55.175 68.870 55.765 68.965 ;
        RECT 56.995 68.870 57.585 68.965 ;
        RECT 55.175 67.085 57.585 68.870 ;
        RECT 58.540 68.670 59.000 69.435 ;
        RECT 59.505 68.945 59.820 69.235 ;
        RECT 59.505 68.935 59.795 68.945 ;
        RECT 61.685 68.755 62.275 68.955 ;
        RECT 59.315 68.670 59.545 68.730 ;
        RECT 58.540 67.840 59.545 68.670 ;
        RECT 55.175 66.860 55.765 67.085 ;
        RECT 56.995 66.860 57.585 67.085 ;
        RECT 53.355 66.100 53.945 66.280 ;
        RECT 55.175 66.100 55.765 66.280 ;
        RECT 51.460 62.820 52.490 65.275 ;
        RECT 53.355 64.315 55.765 66.100 ;
        RECT 56.995 65.950 57.585 66.280 ;
        RECT 53.355 64.175 53.945 64.315 ;
        RECT 55.175 64.175 55.765 64.315 ;
        RECT 56.970 64.175 57.585 65.950 ;
        RECT 56.970 62.985 57.500 64.175 ;
        RECT 51.460 62.715 51.690 62.820 ;
        RECT 51.215 62.510 51.545 62.515 ;
        RECT 51.210 62.280 51.545 62.510 ;
        RECT 51.215 62.255 51.545 62.280 ;
        RECT 51.215 62.085 51.475 62.255 ;
        RECT 50.880 61.085 51.880 62.085 ;
        RECT 46.890 60.865 47.480 60.920 ;
        RECT 48.710 60.865 49.300 60.940 ;
        RECT 51.215 60.765 51.545 61.085 ;
        RECT 51.190 60.550 51.545 60.765 ;
        RECT 51.190 60.535 51.480 60.550 ;
        RECT 51.000 60.315 51.230 60.375 ;
        RECT 46.890 60.195 47.480 60.285 ;
        RECT 46.770 57.670 47.495 60.195 ;
        RECT 48.710 60.185 49.300 60.285 ;
        RECT 48.705 58.090 49.300 60.185 ;
        RECT 50.565 59.530 51.230 60.315 ;
        RECT 50.205 58.445 51.230 59.530 ;
        RECT 48.705 57.670 49.300 57.680 ;
        RECT 50.205 57.670 50.665 58.445 ;
        RECT 51.000 58.375 51.230 58.445 ;
        RECT 51.440 60.305 51.670 60.375 ;
        RECT 52.115 60.305 52.490 62.820 ;
        RECT 53.355 62.805 53.945 62.985 ;
        RECT 55.175 62.805 55.765 62.985 ;
        RECT 53.355 61.020 55.765 62.805 ;
        RECT 53.355 60.880 53.945 61.020 ;
        RECT 55.175 60.880 55.765 61.020 ;
        RECT 56.970 61.005 57.585 62.985 ;
        RECT 58.870 62.795 59.545 67.840 ;
        RECT 59.315 62.730 59.545 62.795 ;
        RECT 59.755 68.675 59.985 68.730 ;
        RECT 60.180 68.675 62.275 68.755 ;
        RECT 59.755 66.970 62.275 68.675 ;
        RECT 59.755 65.390 60.700 66.970 ;
        RECT 61.685 66.850 62.275 66.970 ;
        RECT 63.505 68.705 64.095 68.955 ;
        RECT 65.325 68.705 65.915 68.955 ;
        RECT 63.505 66.920 65.915 68.705 ;
        RECT 66.875 68.650 67.335 69.435 ;
        RECT 67.820 68.920 68.135 69.210 ;
        RECT 67.630 68.650 67.860 68.720 ;
        RECT 66.875 67.850 67.860 68.650 ;
        RECT 63.505 66.850 64.095 66.920 ;
        RECT 65.325 66.850 65.915 66.920 ;
        RECT 61.685 66.015 62.275 66.270 ;
        RECT 63.505 66.015 64.095 66.270 ;
        RECT 59.755 62.840 60.880 65.390 ;
        RECT 61.685 64.230 64.095 66.015 ;
        RECT 65.325 65.940 65.915 66.270 ;
        RECT 61.685 64.165 62.275 64.230 ;
        RECT 63.505 64.165 64.095 64.230 ;
        RECT 59.755 62.730 59.985 62.840 ;
        RECT 59.505 62.495 59.795 62.525 ;
        RECT 59.495 62.080 59.825 62.495 ;
        RECT 59.165 61.080 60.165 62.080 ;
        RECT 56.995 60.880 57.585 61.005 ;
        RECT 59.495 60.530 59.825 61.080 ;
        RECT 51.440 58.485 52.515 60.305 ;
        RECT 51.440 58.375 51.670 58.485 ;
        RECT 51.190 57.930 51.505 58.220 ;
        RECT 53.355 58.195 53.945 60.300 ;
        RECT 55.175 60.085 55.765 60.300 ;
        RECT 55.995 60.085 56.590 60.160 ;
        RECT 56.995 60.085 57.585 60.300 ;
        RECT 59.305 60.285 59.535 60.375 ;
        RECT 59.745 60.295 59.975 60.375 ;
        RECT 60.505 60.295 60.880 62.840 ;
        RECT 61.685 62.845 62.275 62.975 ;
        RECT 63.505 62.845 64.095 62.975 ;
        RECT 61.685 61.060 64.095 62.845 ;
        RECT 61.685 60.870 62.275 61.060 ;
        RECT 63.505 60.870 64.095 61.060 ;
        RECT 65.315 60.920 65.940 65.940 ;
        RECT 67.225 62.775 67.860 67.850 ;
        RECT 67.630 62.720 67.860 62.775 ;
        RECT 68.070 68.700 68.300 68.720 ;
        RECT 68.070 68.680 68.995 68.700 ;
        RECT 69.980 68.680 70.570 68.945 ;
        RECT 68.070 66.865 70.570 68.680 ;
        RECT 68.070 65.265 68.995 66.865 ;
        RECT 69.980 66.840 70.570 66.865 ;
        RECT 71.800 68.760 72.390 68.945 ;
        RECT 73.620 68.760 74.210 68.945 ;
        RECT 71.800 66.945 74.210 68.760 ;
        RECT 75.250 68.790 75.710 69.435 ;
        RECT 76.185 69.045 76.500 69.335 ;
        RECT 76.200 69.025 76.490 69.045 ;
        RECT 76.010 68.790 76.240 68.820 ;
        RECT 75.250 68.230 76.240 68.790 ;
        RECT 71.800 66.840 72.390 66.945 ;
        RECT 73.620 66.840 74.210 66.945 ;
        RECT 69.980 66.120 70.570 66.260 ;
        RECT 71.800 66.120 72.390 66.260 ;
        RECT 68.070 62.865 69.070 65.265 ;
        RECT 69.980 64.305 72.390 66.120 ;
        RECT 69.980 64.155 70.570 64.305 ;
        RECT 71.800 64.155 72.390 64.305 ;
        RECT 73.620 65.980 74.210 66.260 ;
        RECT 68.070 62.720 68.300 62.865 ;
        RECT 67.785 62.285 68.110 62.515 ;
        RECT 67.785 61.965 68.045 62.285 ;
        RECT 67.525 60.965 68.525 61.965 ;
        RECT 65.325 60.870 65.915 60.920 ;
        RECT 67.785 60.765 68.045 60.965 ;
        RECT 67.755 60.535 68.045 60.765 ;
        RECT 55.175 58.300 57.585 60.085 ;
        RECT 58.950 59.680 59.550 60.285 ;
        RECT 55.175 58.195 55.765 58.300 ;
        RECT 56.995 58.195 57.585 58.300 ;
        RECT 58.630 58.415 59.550 59.680 ;
        RECT 59.745 58.605 60.880 60.295 ;
        RECT 59.745 58.475 60.795 58.605 ;
        RECT 58.630 57.670 59.090 58.415 ;
        RECT 59.305 58.375 59.535 58.415 ;
        RECT 59.745 58.375 59.975 58.475 ;
        RECT 59.495 57.940 59.810 58.230 ;
        RECT 61.685 58.185 62.275 60.290 ;
        RECT 63.505 60.025 64.095 60.290 ;
        RECT 64.250 60.025 64.840 60.090 ;
        RECT 65.325 60.025 65.915 60.290 ;
        RECT 67.565 60.275 67.795 60.375 ;
        RECT 63.505 58.240 65.915 60.025 ;
        RECT 67.175 59.690 67.795 60.275 ;
        RECT 63.505 58.185 64.095 58.240 ;
        RECT 65.325 58.185 65.915 58.240 ;
        RECT 66.825 58.405 67.795 59.690 ;
        RECT 61.700 58.160 62.245 58.185 ;
        RECT 66.825 57.670 67.285 58.405 ;
        RECT 67.565 58.375 67.795 58.405 ;
        RECT 68.005 60.280 68.235 60.375 ;
        RECT 68.695 60.280 69.070 62.865 ;
        RECT 69.980 62.815 70.570 62.965 ;
        RECT 71.800 62.815 72.390 62.965 ;
        RECT 69.980 61.000 72.390 62.815 ;
        RECT 69.980 60.860 70.570 61.000 ;
        RECT 71.800 60.860 72.390 61.000 ;
        RECT 73.620 60.960 74.245 65.980 ;
        RECT 75.570 62.915 76.240 68.230 ;
        RECT 76.010 62.820 76.240 62.915 ;
        RECT 76.450 68.750 76.680 68.820 ;
        RECT 76.450 68.700 77.350 68.750 ;
        RECT 78.425 68.700 79.015 68.960 ;
        RECT 76.450 66.885 79.015 68.700 ;
        RECT 76.450 65.315 77.350 66.885 ;
        RECT 78.425 66.855 79.015 66.885 ;
        RECT 80.245 68.820 80.835 68.960 ;
        RECT 82.065 68.820 82.655 68.960 ;
        RECT 80.245 67.005 82.655 68.820 ;
        RECT 83.675 68.700 84.135 69.435 ;
        RECT 84.590 68.960 84.905 69.250 ;
        RECT 84.590 68.950 84.880 68.960 ;
        RECT 86.755 68.760 87.345 68.960 ;
        RECT 84.905 68.745 87.345 68.760 ;
        RECT 84.400 68.700 84.630 68.745 ;
        RECT 83.675 68.210 84.630 68.700 ;
        RECT 80.245 66.855 80.835 67.005 ;
        RECT 82.065 66.855 82.655 67.005 ;
        RECT 78.425 66.020 79.015 66.275 ;
        RECT 80.245 66.020 80.835 66.275 ;
        RECT 82.065 66.205 82.655 66.275 ;
        RECT 76.450 62.915 77.475 65.315 ;
        RECT 78.425 64.205 80.835 66.020 ;
        RECT 78.425 64.170 79.015 64.205 ;
        RECT 80.245 64.170 80.835 64.205 ;
        RECT 76.450 62.820 76.680 62.915 ;
        RECT 76.200 62.385 76.490 62.615 ;
        RECT 76.210 62.125 76.460 62.385 ;
        RECT 75.925 61.125 76.925 62.125 ;
        RECT 73.620 60.860 74.210 60.960 ;
        RECT 76.210 60.785 76.460 61.125 ;
        RECT 76.175 60.555 76.465 60.785 ;
        RECT 75.985 60.315 76.215 60.395 ;
        RECT 68.005 58.460 69.090 60.280 ;
        RECT 69.980 60.130 70.570 60.280 ;
        RECT 68.005 58.375 68.235 58.460 ;
        RECT 67.755 58.195 68.045 58.215 ;
        RECT 67.755 57.985 68.110 58.195 ;
        RECT 69.970 58.175 70.570 60.130 ;
        RECT 71.800 60.035 72.390 60.280 ;
        RECT 73.620 60.035 74.210 60.280 ;
        RECT 71.800 58.220 74.210 60.035 ;
        RECT 75.550 59.830 76.215 60.315 ;
        RECT 75.230 59.780 76.215 59.830 ;
        RECT 71.800 58.175 72.390 58.220 ;
        RECT 73.620 58.175 74.210 58.220 ;
        RECT 75.080 58.445 76.215 59.780 ;
        RECT 69.970 58.140 70.515 58.175 ;
        RECT 67.795 57.905 68.110 57.985 ;
        RECT 75.080 57.710 75.690 58.445 ;
        RECT 75.985 58.395 76.215 58.445 ;
        RECT 76.425 60.305 76.655 60.395 ;
        RECT 77.100 60.305 77.475 62.915 ;
        RECT 78.425 62.715 79.015 62.980 ;
        RECT 80.245 62.715 80.835 62.980 ;
        RECT 78.425 60.900 80.835 62.715 ;
        RECT 78.425 60.875 79.015 60.900 ;
        RECT 80.245 60.875 80.835 60.900 ;
        RECT 82.045 60.885 82.665 66.205 ;
        RECT 84.045 62.825 84.630 68.210 ;
        RECT 84.400 62.745 84.630 62.825 ;
        RECT 84.840 66.945 87.345 68.745 ;
        RECT 84.840 65.250 85.730 66.945 ;
        RECT 86.755 66.855 87.345 66.945 ;
        RECT 88.575 68.800 89.165 68.960 ;
        RECT 90.395 68.800 90.985 68.960 ;
        RECT 88.575 66.985 90.985 68.800 ;
        RECT 92.130 68.750 92.590 69.435 ;
        RECT 92.905 68.995 93.220 69.285 ;
        RECT 92.920 68.975 93.210 68.995 ;
        RECT 92.730 68.750 92.960 68.770 ;
        RECT 92.130 67.930 92.960 68.750 ;
        RECT 88.575 66.855 89.165 66.985 ;
        RECT 90.395 66.855 90.985 66.985 ;
        RECT 86.755 66.060 87.345 66.275 ;
        RECT 88.575 66.060 89.165 66.275 ;
        RECT 84.840 62.815 85.955 65.250 ;
        RECT 86.755 64.245 89.165 66.060 ;
        RECT 90.395 65.980 90.985 66.275 ;
        RECT 86.755 64.170 87.345 64.245 ;
        RECT 88.575 64.170 89.165 64.245 ;
        RECT 84.840 62.745 85.070 62.815 ;
        RECT 84.585 62.540 84.835 62.550 ;
        RECT 84.585 62.310 84.880 62.540 ;
        RECT 84.585 62.085 84.835 62.310 ;
        RECT 84.370 61.085 85.370 62.085 ;
        RECT 82.065 60.875 82.655 60.885 ;
        RECT 84.585 60.765 84.835 61.085 ;
        RECT 84.525 60.565 84.835 60.765 ;
        RECT 84.525 60.535 84.815 60.565 ;
        RECT 76.425 58.485 77.475 60.305 ;
        RECT 84.335 60.295 84.565 60.375 ;
        RECT 76.425 58.395 76.655 58.485 ;
        RECT 76.175 58.220 76.465 58.235 ;
        RECT 76.160 57.930 76.475 58.220 ;
        RECT 78.425 58.175 79.015 60.295 ;
        RECT 80.245 60.055 80.835 60.295 ;
        RECT 82.065 60.055 82.655 60.295 ;
        RECT 80.245 58.240 82.655 60.055 ;
        RECT 83.915 59.840 84.565 60.295 ;
        RECT 80.245 58.190 80.835 58.240 ;
        RECT 82.065 58.190 82.655 58.240 ;
        RECT 83.475 58.395 84.565 59.840 ;
        RECT 74.235 57.670 75.690 57.710 ;
        RECT 83.475 57.670 83.935 58.395 ;
        RECT 84.335 58.375 84.565 58.395 ;
        RECT 84.775 60.255 85.005 60.375 ;
        RECT 85.580 60.255 85.955 62.815 ;
        RECT 86.755 62.795 87.345 62.980 ;
        RECT 88.575 62.795 89.165 62.980 ;
        RECT 86.755 60.980 89.165 62.795 ;
        RECT 86.755 60.875 87.345 60.980 ;
        RECT 88.575 60.875 89.165 60.980 ;
        RECT 90.370 60.960 90.995 65.980 ;
        RECT 92.300 62.875 92.960 67.930 ;
        RECT 92.730 62.770 92.960 62.875 ;
        RECT 93.170 68.685 93.400 68.770 ;
        RECT 93.170 68.680 94.090 68.685 ;
        RECT 95.085 68.680 95.675 68.960 ;
        RECT 93.170 66.865 95.675 68.680 ;
        RECT 93.170 65.275 94.090 66.865 ;
        RECT 95.085 66.855 95.675 66.865 ;
        RECT 96.905 68.780 97.495 68.960 ;
        RECT 98.725 68.780 99.315 68.960 ;
        RECT 96.905 66.965 99.315 68.780 ;
        RECT 100.370 68.710 100.830 69.435 ;
        RECT 101.210 68.970 101.525 69.260 ;
        RECT 101.025 68.710 101.255 68.785 ;
        RECT 100.370 67.980 101.255 68.710 ;
        RECT 96.905 66.855 97.495 66.965 ;
        RECT 98.725 66.855 99.315 66.965 ;
        RECT 95.085 66.020 95.675 66.275 ;
        RECT 96.905 66.020 97.495 66.275 ;
        RECT 98.725 66.020 99.315 66.275 ;
        RECT 93.170 62.850 94.285 65.275 ;
        RECT 95.085 64.205 97.505 66.020 ;
        RECT 95.085 64.170 95.675 64.205 ;
        RECT 96.905 64.170 97.495 64.205 ;
        RECT 93.170 62.770 93.400 62.850 ;
        RECT 92.920 62.335 93.210 62.565 ;
        RECT 92.920 62.070 93.170 62.335 ;
        RECT 92.640 61.070 93.640 62.070 ;
        RECT 90.395 60.875 90.985 60.960 ;
        RECT 92.920 60.760 93.170 61.070 ;
        RECT 92.910 60.530 93.200 60.760 ;
        RECT 92.720 60.315 92.950 60.370 ;
        RECT 84.775 58.465 85.955 60.255 ;
        RECT 86.755 60.280 87.345 60.295 ;
        RECT 84.775 58.435 85.840 58.465 ;
        RECT 84.775 58.375 85.005 58.435 ;
        RECT 86.755 58.260 87.350 60.280 ;
        RECT 88.575 60.075 89.165 60.295 ;
        RECT 90.395 60.075 90.985 60.295 ;
        RECT 88.575 58.260 90.985 60.075 ;
        RECT 92.320 59.850 92.950 60.315 ;
        RECT 84.515 57.940 84.830 58.230 ;
        RECT 86.755 58.190 87.345 58.260 ;
        RECT 88.575 58.190 89.165 58.260 ;
        RECT 89.385 58.175 89.975 58.260 ;
        RECT 90.395 58.190 90.985 58.260 ;
        RECT 91.910 58.415 92.950 59.850 ;
        RECT 91.910 57.670 92.370 58.415 ;
        RECT 92.720 58.370 92.950 58.415 ;
        RECT 93.160 60.245 93.390 60.370 ;
        RECT 93.910 60.245 94.285 62.850 ;
        RECT 95.085 62.775 95.675 62.980 ;
        RECT 96.905 62.775 97.495 62.980 ;
        RECT 95.085 60.960 97.495 62.775 ;
        RECT 98.690 61.000 99.315 66.020 ;
        RECT 100.580 62.835 101.255 67.980 ;
        RECT 101.025 62.785 101.255 62.835 ;
        RECT 101.465 68.680 101.695 68.785 ;
        RECT 103.390 68.680 103.980 68.955 ;
        RECT 101.465 66.865 103.980 68.680 ;
        RECT 101.465 65.375 102.370 66.865 ;
        RECT 103.390 66.850 103.980 66.865 ;
        RECT 105.210 68.780 105.800 68.955 ;
        RECT 107.030 68.780 107.620 68.955 ;
        RECT 105.210 66.965 107.620 68.780 ;
        RECT 108.645 68.710 109.105 69.435 ;
        RECT 109.525 69.200 109.840 69.275 ;
        RECT 109.515 68.985 109.840 69.200 ;
        RECT 109.515 68.970 109.805 68.985 ;
        RECT 111.690 68.780 112.280 68.965 ;
        RECT 113.510 68.780 114.100 68.965 ;
        RECT 109.325 68.710 109.555 68.765 ;
        RECT 108.645 67.750 109.555 68.710 ;
        RECT 105.210 66.850 105.800 66.965 ;
        RECT 107.030 66.850 107.620 66.965 ;
        RECT 103.390 66.020 103.980 66.270 ;
        RECT 105.210 66.020 105.800 66.270 ;
        RECT 101.465 62.825 102.505 65.375 ;
        RECT 103.390 64.205 105.800 66.020 ;
        RECT 103.390 64.165 103.980 64.205 ;
        RECT 105.210 64.165 105.800 64.205 ;
        RECT 107.030 66.000 107.620 66.270 ;
        RECT 107.030 64.165 107.680 66.000 ;
        RECT 107.055 62.975 107.680 64.165 ;
        RECT 101.465 62.785 101.695 62.825 ;
        RECT 101.170 62.100 101.515 62.590 ;
        RECT 100.945 61.100 101.945 62.100 ;
        RECT 95.085 60.875 95.675 60.960 ;
        RECT 96.905 60.875 97.495 60.960 ;
        RECT 98.725 60.875 99.315 61.000 ;
        RECT 101.170 60.770 101.515 61.100 ;
        RECT 101.150 60.555 101.515 60.770 ;
        RECT 101.150 60.540 101.440 60.555 ;
        RECT 100.960 60.305 101.190 60.380 ;
        RECT 93.160 58.490 94.285 60.245 ;
        RECT 95.085 60.200 95.675 60.295 ;
        RECT 93.160 58.425 94.200 58.490 ;
        RECT 93.160 58.370 93.390 58.425 ;
        RECT 92.910 58.195 93.200 58.210 ;
        RECT 92.910 57.980 93.250 58.195 ;
        RECT 95.070 58.190 95.675 60.200 ;
        RECT 96.905 60.075 97.495 60.295 ;
        RECT 98.725 60.075 99.315 60.295 ;
        RECT 96.880 58.260 99.315 60.075 ;
        RECT 100.630 59.810 101.190 60.305 ;
        RECT 96.905 58.190 97.495 58.260 ;
        RECT 98.725 58.190 99.315 58.260 ;
        RECT 100.200 58.405 101.190 59.810 ;
        RECT 95.070 58.170 95.615 58.190 ;
        RECT 92.935 57.905 93.250 57.980 ;
        RECT 100.200 57.670 100.660 58.405 ;
        RECT 100.960 58.380 101.190 58.405 ;
        RECT 101.400 60.280 101.630 60.380 ;
        RECT 102.130 60.280 102.505 62.825 ;
        RECT 103.390 62.775 103.980 62.975 ;
        RECT 105.210 62.775 105.800 62.975 ;
        RECT 103.390 60.960 105.800 62.775 ;
        RECT 103.390 60.870 103.980 60.960 ;
        RECT 105.210 60.870 105.800 60.960 ;
        RECT 107.030 60.980 107.680 62.975 ;
        RECT 108.895 62.835 109.555 67.750 ;
        RECT 109.325 62.765 109.555 62.835 ;
        RECT 109.765 68.745 109.995 68.765 ;
        RECT 109.765 66.160 110.550 68.745 ;
        RECT 111.690 66.965 114.100 68.780 ;
        RECT 111.690 66.860 112.280 66.965 ;
        RECT 113.510 66.860 114.100 66.965 ;
        RECT 111.690 66.160 112.280 66.280 ;
        RECT 109.765 64.345 112.280 66.160 ;
        RECT 113.510 66.040 114.100 66.280 ;
        RECT 109.765 63.580 110.550 64.345 ;
        RECT 111.690 64.175 112.280 64.345 ;
        RECT 113.445 64.175 114.100 66.040 ;
        RECT 109.765 62.845 110.590 63.580 ;
        RECT 109.765 62.765 109.995 62.845 ;
        RECT 109.515 62.505 109.805 62.560 ;
        RECT 109.515 62.495 110.030 62.505 ;
        RECT 109.485 62.060 110.030 62.495 ;
        RECT 110.260 62.265 110.590 62.845 ;
        RECT 111.510 62.695 112.510 63.695 ;
        RECT 113.445 62.985 114.070 64.175 ;
        RECT 109.035 61.060 110.035 62.060 ;
        RECT 110.330 61.265 110.590 62.265 ;
        RECT 107.030 60.870 107.620 60.980 ;
        RECT 109.485 60.595 110.030 61.060 ;
        RECT 110.305 60.970 110.590 61.265 ;
        RECT 111.620 61.010 112.335 62.695 ;
        RECT 113.445 61.020 114.100 62.985 ;
        RECT 109.485 60.585 109.960 60.595 ;
        RECT 109.515 60.570 109.960 60.585 ;
        RECT 109.515 60.540 109.805 60.570 ;
        RECT 109.325 60.335 109.555 60.380 ;
        RECT 101.400 58.590 102.505 60.280 ;
        RECT 103.390 60.180 103.980 60.290 ;
        RECT 101.400 58.460 102.465 58.590 ;
        RECT 101.400 58.380 101.630 58.460 ;
        RECT 101.210 58.220 101.525 58.230 ;
        RECT 101.150 57.990 101.525 58.220 ;
        RECT 103.375 58.185 103.980 60.180 ;
        RECT 105.210 60.135 105.800 60.290 ;
        RECT 107.030 60.135 107.620 60.290 ;
        RECT 105.210 58.320 107.620 60.135 ;
        RECT 108.975 59.900 109.555 60.335 ;
        RECT 105.210 58.185 105.800 58.320 ;
        RECT 103.375 58.160 103.920 58.185 ;
        RECT 106.145 58.170 106.690 58.320 ;
        RECT 107.030 58.185 107.620 58.320 ;
        RECT 108.555 58.435 109.555 59.900 ;
        RECT 101.210 57.940 101.525 57.990 ;
        RECT 108.555 57.670 109.015 58.435 ;
        RECT 109.325 58.380 109.555 58.435 ;
        RECT 109.765 60.320 109.995 60.380 ;
        RECT 110.260 60.320 110.590 60.970 ;
        RECT 111.690 60.975 112.295 61.010 ;
        RECT 111.690 60.880 112.280 60.975 ;
        RECT 113.510 60.880 114.100 61.020 ;
        RECT 109.765 58.825 110.590 60.320 ;
        RECT 111.690 60.115 112.280 60.300 ;
        RECT 113.510 60.115 114.100 60.300 ;
        RECT 109.765 58.440 110.365 58.825 ;
        RECT 109.765 58.380 109.995 58.440 ;
        RECT 111.690 58.300 114.100 60.115 ;
        RECT 109.490 57.930 109.805 58.220 ;
        RECT 111.690 58.195 112.280 58.300 ;
        RECT 113.510 58.195 114.100 58.300 ;
        RECT 10.970 57.310 13.930 57.410 ;
        RECT 2.150 57.280 4.255 57.310 ;
        RECT 2.090 56.720 4.255 57.280 ;
        RECT 4.835 57.280 6.940 57.310 ;
        RECT 8.130 57.280 10.235 57.310 ;
        RECT 4.835 56.720 10.235 57.280 ;
        RECT 10.815 56.720 13.930 57.310 ;
        RECT 46.190 57.190 114.805 57.670 ;
        RECT 2.090 55.490 3.990 56.720 ;
        RECT 4.890 56.680 10.190 56.720 ;
        RECT 10.970 56.630 13.930 56.720 ;
        RECT 46.180 56.610 114.810 57.190 ;
        RECT 2.090 54.900 4.255 55.490 ;
        RECT 4.835 55.480 6.940 55.490 ;
        RECT 8.130 55.480 10.235 55.490 ;
        RECT 4.835 54.900 10.235 55.480 ;
        RECT 10.815 54.900 12.920 55.490 ;
        RECT 2.090 54.880 3.990 54.900 ;
        RECT 4.890 54.880 10.190 54.900 ;
        RECT 2.290 53.670 4.190 53.680 ;
        RECT 4.890 53.670 10.190 53.680 ;
        RECT 10.890 53.670 12.790 54.900 ;
        RECT 2.150 53.080 4.255 53.670 ;
        RECT 4.835 53.080 10.235 53.670 ;
        RECT 10.815 53.080 12.920 53.670 ;
        RECT 2.290 51.850 4.190 53.080 ;
        RECT 61.420 52.540 61.630 52.570 ;
        RECT 61.420 52.090 67.670 52.540 ;
        RECT 61.420 52.060 61.630 52.090 ;
        RECT 10.890 51.875 13.215 51.880 ;
        RECT 10.890 51.850 16.180 51.875 ;
        RECT 25.745 51.850 26.120 51.945 ;
        RECT 41.065 51.875 46.190 51.880 ;
        RECT 28.820 51.850 46.190 51.875 ;
        RECT 46.890 51.850 52.190 51.980 ;
        RECT 52.890 51.850 58.190 51.880 ;
        RECT 58.890 51.850 70.290 51.880 ;
        RECT 70.890 51.850 76.190 51.880 ;
        RECT 76.890 51.850 82.190 51.880 ;
        RECT 2.150 51.260 4.255 51.850 ;
        RECT 4.835 51.780 6.940 51.850 ;
        RECT 8.130 51.780 10.235 51.850 ;
        RECT 4.835 51.260 10.235 51.780 ;
        RECT 10.815 51.260 16.215 51.850 ;
        RECT 16.795 51.260 22.195 51.850 ;
        RECT 22.775 51.810 24.880 51.850 ;
        RECT 25.745 51.810 28.175 51.850 ;
        RECT 22.775 51.260 28.175 51.810 ;
        RECT 28.755 51.270 46.275 51.850 ;
        RECT 28.755 51.260 30.860 51.270 ;
        RECT 41.065 51.260 46.275 51.270 ;
        RECT 46.855 51.280 52.255 51.850 ;
        RECT 46.855 51.260 48.960 51.280 ;
        RECT 50.150 51.260 52.255 51.280 ;
        RECT 52.835 51.260 58.235 51.850 ;
        RECT 58.815 51.260 70.290 51.850 ;
        RECT 70.855 51.260 76.255 51.850 ;
        RECT 76.835 51.280 82.235 51.850 ;
        RECT 76.835 51.260 78.940 51.280 ;
        RECT 80.130 51.260 82.235 51.280 ;
        RECT 82.815 51.260 84.920 51.850 ;
        RECT 4.890 51.180 10.190 51.260 ;
        RECT 10.890 51.180 16.180 51.260 ;
        RECT 16.840 51.255 22.160 51.260 ;
        RECT 12.720 51.170 16.180 51.180 ;
        RECT 1.560 50.360 9.985 50.855 ;
        RECT 10.520 50.500 11.025 50.595 ;
        RECT 17.030 50.500 17.285 51.255 ;
        RECT 22.810 51.215 28.130 51.260 ;
        RECT 28.855 50.575 29.260 51.260 ;
        RECT 41.065 51.180 46.190 51.260 ;
        RECT 47.135 50.630 47.510 51.260 ;
        RECT 52.890 51.180 58.190 51.260 ;
        RECT 58.890 51.180 70.290 51.260 ;
        RECT 70.890 51.180 76.190 51.260 ;
        RECT 59.065 50.680 59.470 51.180 ;
        RECT 10.520 50.245 17.285 50.500 ;
        RECT 10.520 50.150 11.025 50.245 ;
        RECT 26.565 50.170 29.260 50.575 ;
        RECT 38.555 50.255 47.510 50.630 ;
        RECT 54.665 50.275 59.470 50.680 ;
        RECT 71.015 50.655 71.365 51.180 ;
        RECT 81.780 50.735 82.120 51.260 ;
        RECT 82.970 51.160 84.910 51.260 ;
        RECT 83.130 50.755 83.525 51.160 ;
        RECT 66.565 50.305 71.365 50.655 ;
        RECT 77.790 50.170 80.360 50.690 ;
        RECT 81.750 50.395 82.150 50.735 ;
        RECT 82.710 50.360 83.525 50.755 ;
        RECT 84.470 51.100 84.910 51.160 ;
        RECT 144.190 51.100 146.190 51.180 ;
        RECT 84.470 50.660 146.190 51.100 ;
        RECT 27.490 49.960 30.190 49.980 ;
        RECT 55.390 49.960 58.090 49.980 ;
        RECT 83.490 49.960 85.790 49.980 ;
        RECT 111.590 49.960 113.890 49.980 ;
        RECT 1.450 49.280 139.925 49.960 ;
        RECT 144.190 49.310 146.190 50.660 ;
        RECT 1.450 49.260 27.925 49.280 ;
        RECT 29.450 49.260 55.925 49.280 ;
        RECT 57.450 49.260 83.925 49.280 ;
        RECT 85.450 49.260 111.925 49.280 ;
        RECT 113.450 49.260 139.925 49.280 ;
        RECT 2.420 48.635 4.330 49.260 ;
        RECT 6.420 48.925 8.305 48.930 ;
        RECT 9.865 48.925 11.750 48.930 ;
        RECT 6.410 48.695 8.370 48.925 ;
        RECT 9.840 48.695 11.800 48.925 ;
        RECT 2.385 48.405 4.385 48.635 ;
        RECT 6.130 48.410 6.360 48.490 ;
        RECT 1.590 48.355 2.085 48.375 ;
        RECT 1.590 45.060 2.180 48.355 ;
        RECT 4.590 48.275 4.820 48.355 ;
        RECT 4.560 45.060 4.820 48.275 ;
        RECT 1.590 43.245 4.820 45.060 ;
        RECT 1.590 40.395 2.180 43.245 ;
        RECT 3.075 40.640 3.335 40.960 ;
        RECT 4.560 40.645 4.820 43.245 ;
        RECT 5.890 40.990 6.360 48.410 ;
        RECT 6.850 41.775 7.740 48.695 ;
        RECT 8.420 48.390 8.650 48.490 ;
        RECT 8.420 48.380 8.775 48.390 ;
        RECT 9.560 48.380 9.790 48.490 ;
        RECT 3.130 40.480 3.280 40.640 ;
        RECT 1.590 35.255 2.085 40.395 ;
        RECT 3.105 40.345 3.310 40.480 ;
        RECT 4.590 40.395 4.820 40.645 ;
        RECT 5.610 40.550 6.360 40.990 ;
        RECT 6.780 40.775 7.795 41.775 ;
        RECT 2.385 40.115 4.385 40.345 ;
        RECT 5.610 38.355 5.980 40.550 ;
        RECT 6.130 40.490 6.360 40.550 ;
        RECT 6.850 40.285 7.740 40.775 ;
        RECT 8.420 40.580 9.790 48.380 ;
        RECT 10.325 43.635 11.215 48.695 ;
        RECT 11.850 48.410 12.080 48.490 ;
        RECT 10.320 42.015 11.220 43.635 ;
        RECT 10.325 41.605 11.215 42.015 ;
        RECT 10.250 40.605 11.280 41.605 ;
        RECT 11.850 40.625 12.225 48.410 ;
        RECT 12.500 48.025 14.180 49.260 ;
        RECT 15.015 48.025 19.940 48.035 ;
        RECT 12.500 47.545 19.940 48.025 ;
        RECT 12.500 45.285 14.180 47.545 ;
        RECT 15.015 47.125 19.940 47.545 ;
        RECT 14.520 46.935 14.775 46.960 ;
        RECT 14.520 46.920 14.795 46.935 ;
        RECT 14.490 46.645 14.825 46.920 ;
        RECT 15.000 46.895 20.000 47.125 ;
        RECT 20.210 46.935 20.465 46.960 ;
        RECT 14.520 46.630 14.775 46.645 ;
        RECT 15.000 46.455 20.000 46.685 ;
        RECT 20.205 46.645 20.465 46.935 ;
        RECT 20.210 46.630 20.465 46.645 ;
        RECT 15.045 46.445 19.900 46.455 ;
        RECT 15.045 44.920 17.690 44.925 ;
        RECT 13.720 44.720 17.690 44.920 ;
        RECT 13.720 44.690 17.680 44.720 ;
        RECT 12.560 44.335 12.895 44.610 ;
        RECT 13.440 44.440 13.670 44.485 ;
        RECT 8.420 40.560 8.775 40.580 ;
        RECT 8.420 40.490 8.650 40.560 ;
        RECT 9.560 40.490 9.790 40.580 ;
        RECT 10.320 40.465 11.230 40.605 ;
        RECT 11.850 40.490 12.240 40.625 ;
        RECT 10.310 40.285 11.320 40.465 ;
        RECT 6.410 40.055 8.370 40.285 ;
        RECT 9.840 40.055 11.800 40.285 ;
        RECT 7.135 39.065 7.465 40.055 ;
        RECT 9.865 40.050 11.750 40.055 ;
        RECT 12.045 38.355 12.240 40.490 ;
        RECT 12.630 38.830 12.820 44.335 ;
        RECT 13.250 43.105 13.670 44.440 ;
        RECT 14.975 43.105 16.320 44.690 ;
        RECT 13.250 41.720 16.320 43.105 ;
        RECT 13.250 40.990 13.670 41.720 ;
        RECT 13.245 40.485 13.670 40.990 ;
        RECT 12.630 38.640 12.945 38.830 ;
        RECT 2.950 38.125 6.910 38.355 ;
        RECT 8.380 38.125 12.340 38.355 ;
        RECT 12.755 38.130 12.945 38.640 ;
        RECT 2.670 37.515 2.900 37.965 ;
        RECT 4.150 37.515 4.940 38.125 ;
        RECT 2.670 37.210 4.940 37.515 ;
        RECT 2.615 37.195 4.940 37.210 ;
        RECT 2.530 36.350 4.940 37.195 ;
        RECT 2.530 35.975 2.900 36.350 ;
        RECT 2.670 35.965 2.900 35.975 ;
        RECT 4.150 35.805 4.940 36.350 ;
        RECT 6.960 37.880 7.190 37.965 ;
        RECT 8.100 37.880 8.330 37.965 ;
        RECT 6.960 36.055 8.330 37.880 ;
        RECT 6.960 35.965 7.190 36.055 ;
        RECT 2.950 35.575 6.910 35.805 ;
        RECT 2.530 35.255 2.755 35.265 ;
        RECT 7.430 35.255 7.920 36.055 ;
        RECT 8.100 35.965 8.330 36.055 ;
        RECT 9.815 37.745 11.155 38.125 ;
        RECT 12.390 37.745 12.620 37.965 ;
        RECT 9.815 36.150 12.620 37.745 ;
        RECT 9.815 35.805 11.155 36.150 ;
        RECT 12.390 35.965 12.620 36.150 ;
        RECT 8.380 35.575 12.340 35.805 ;
        RECT 12.770 35.785 12.945 38.130 ;
        RECT 13.245 37.965 13.540 40.485 ;
        RECT 14.975 40.280 16.320 41.720 ;
        RECT 17.730 44.390 17.960 44.485 ;
        RECT 18.205 44.390 18.695 46.445 ;
        RECT 19.265 44.920 19.900 44.925 ;
        RECT 19.150 44.690 23.110 44.920 ;
        RECT 18.870 44.390 19.100 44.485 ;
        RECT 17.730 40.565 19.100 44.390 ;
        RECT 17.730 40.485 17.960 40.565 ;
        RECT 18.870 40.485 19.100 40.565 ;
        RECT 20.525 40.280 21.870 44.690 ;
        RECT 23.160 44.420 23.390 44.485 ;
        RECT 24.045 44.425 24.520 49.260 ;
        RECT 25.845 48.455 26.525 49.260 ;
        RECT 26.945 48.735 27.280 48.985 ;
        RECT 26.960 48.710 27.250 48.735 ;
        RECT 30.420 48.635 32.330 49.260 ;
        RECT 34.420 48.925 36.305 48.930 ;
        RECT 37.865 48.925 39.750 48.930 ;
        RECT 34.410 48.695 36.370 48.925 ;
        RECT 37.840 48.695 39.800 48.925 ;
        RECT 26.770 48.455 27.000 48.505 ;
        RECT 25.845 47.955 27.000 48.455 ;
        RECT 24.915 44.735 25.250 44.985 ;
        RECT 24.935 44.705 25.225 44.735 ;
        RECT 24.745 44.425 24.975 44.500 ;
        RECT 23.160 40.485 23.615 44.420 ;
        RECT 24.045 43.680 24.975 44.425 ;
        RECT 24.380 40.565 24.975 43.680 ;
        RECT 24.745 40.500 24.975 40.565 ;
        RECT 25.185 44.475 25.415 44.500 ;
        RECT 25.185 40.920 25.695 44.475 ;
        RECT 25.185 40.550 25.880 40.920 ;
        RECT 26.380 40.600 27.000 47.955 ;
        RECT 25.185 40.500 25.415 40.550 ;
        RECT 13.720 40.250 17.680 40.280 ;
        RECT 19.150 40.250 23.110 40.280 ;
        RECT 13.720 40.090 23.110 40.250 ;
        RECT 13.720 40.050 17.680 40.090 ;
        RECT 19.150 40.050 23.110 40.090 ;
        RECT 23.275 38.660 23.615 40.485 ;
        RECT 24.925 38.660 25.345 40.305 ;
        RECT 23.275 38.505 25.345 38.660 ;
        RECT 23.350 38.390 25.345 38.505 ;
        RECT 13.810 38.125 17.770 38.355 ;
        RECT 19.240 38.125 23.200 38.355 ;
        RECT 13.245 37.205 13.760 37.965 ;
        RECT 13.315 36.025 13.760 37.205 ;
        RECT 13.530 35.965 13.760 36.025 ;
        RECT 15.190 35.805 16.145 38.125 ;
        RECT 17.820 37.900 18.050 37.965 ;
        RECT 18.960 37.900 19.190 37.965 ;
        RECT 17.820 36.030 19.190 37.900 ;
        RECT 17.820 35.965 18.050 36.030 ;
        RECT 12.755 35.255 12.945 35.785 ;
        RECT 13.810 35.575 17.770 35.805 ;
        RECT 18.225 35.255 18.780 36.030 ;
        RECT 18.960 35.965 19.190 36.030 ;
        RECT 20.635 35.805 21.590 38.125 ;
        RECT 23.350 37.970 23.615 38.390 ;
        RECT 24.925 38.115 25.345 38.390 ;
        RECT 25.580 39.355 25.880 40.550 ;
        RECT 26.770 40.505 27.000 40.600 ;
        RECT 27.210 48.430 27.440 48.505 ;
        RECT 27.210 41.110 27.985 48.430 ;
        RECT 30.385 48.405 32.385 48.635 ;
        RECT 34.130 48.410 34.360 48.490 ;
        RECT 29.950 45.060 30.180 48.355 ;
        RECT 32.590 48.275 32.820 48.355 ;
        RECT 32.560 45.060 32.820 48.275 ;
        RECT 29.950 43.245 32.820 45.060 ;
        RECT 27.210 40.580 28.060 41.110 ;
        RECT 29.950 40.825 30.180 43.245 ;
        RECT 27.210 40.505 27.440 40.580 ;
        RECT 26.875 39.825 27.390 40.315 ;
        RECT 27.690 39.825 28.060 40.580 ;
        RECT 29.590 40.395 30.180 40.825 ;
        RECT 31.075 40.640 31.335 40.960 ;
        RECT 32.560 40.645 32.820 43.245 ;
        RECT 33.890 40.990 34.360 48.410 ;
        RECT 34.850 41.775 35.740 48.695 ;
        RECT 36.420 48.390 36.650 48.490 ;
        RECT 36.420 48.380 36.775 48.390 ;
        RECT 37.560 48.380 37.790 48.490 ;
        RECT 31.130 40.480 31.280 40.640 ;
        RECT 26.875 39.360 27.385 39.825 ;
        RECT 26.510 39.355 27.385 39.360 ;
        RECT 25.580 38.950 27.385 39.355 ;
        RECT 25.580 38.110 25.880 38.950 ;
        RECT 26.510 38.935 27.385 38.950 ;
        RECT 26.875 38.825 27.385 38.935 ;
        RECT 26.875 38.125 27.390 38.825 ;
        RECT 27.615 38.795 28.615 39.825 ;
        RECT 23.275 37.965 23.615 37.970 ;
        RECT 23.250 36.020 23.615 37.965 ;
        RECT 24.830 37.900 25.060 37.970 ;
        RECT 24.335 37.230 25.060 37.900 ;
        RECT 24.325 37.040 25.060 37.230 ;
        RECT 24.325 36.240 24.680 37.040 ;
        RECT 24.830 36.970 25.060 37.040 ;
        RECT 25.270 37.925 25.500 37.970 ;
        RECT 25.640 37.925 25.880 38.110 ;
        RECT 25.270 37.595 25.880 37.925 ;
        RECT 26.855 37.870 27.085 37.975 ;
        RECT 25.270 37.040 25.765 37.595 ;
        RECT 25.270 36.970 25.500 37.040 ;
        RECT 25.020 36.785 25.310 36.810 ;
        RECT 25.005 36.535 25.340 36.785 ;
        RECT 26.625 36.765 27.085 37.870 ;
        RECT 26.305 36.240 27.085 36.765 ;
        RECT 23.885 36.060 27.085 36.240 ;
        RECT 23.250 35.965 23.480 36.020 ;
        RECT 19.240 35.575 23.200 35.805 ;
        RECT 23.885 35.620 26.690 36.060 ;
        RECT 26.855 35.975 27.085 36.060 ;
        RECT 27.295 37.910 27.525 37.975 ;
        RECT 27.690 37.910 28.060 38.795 ;
        RECT 27.295 37.585 28.060 37.910 ;
        RECT 27.295 36.045 28.055 37.585 ;
        RECT 27.295 35.975 27.525 36.045 ;
        RECT 27.045 35.795 27.335 35.815 ;
        RECT 23.885 35.255 26.350 35.620 ;
        RECT 27.020 35.545 27.355 35.795 ;
        RECT 29.590 35.280 30.085 40.395 ;
        RECT 31.105 40.345 31.310 40.480 ;
        RECT 32.590 40.395 32.820 40.645 ;
        RECT 33.610 40.550 34.360 40.990 ;
        RECT 34.780 40.775 35.795 41.775 ;
        RECT 30.385 40.115 32.385 40.345 ;
        RECT 33.610 38.355 33.980 40.550 ;
        RECT 34.130 40.490 34.360 40.550 ;
        RECT 34.850 40.285 35.740 40.775 ;
        RECT 36.420 40.580 37.790 48.380 ;
        RECT 38.325 43.635 39.215 48.695 ;
        RECT 39.850 48.410 40.080 48.490 ;
        RECT 38.320 42.015 39.220 43.635 ;
        RECT 38.325 41.605 39.215 42.015 ;
        RECT 38.250 40.605 39.280 41.605 ;
        RECT 39.850 40.625 40.225 48.410 ;
        RECT 40.500 48.025 42.180 49.260 ;
        RECT 43.015 48.025 47.940 48.035 ;
        RECT 40.500 47.545 47.940 48.025 ;
        RECT 40.500 45.285 42.180 47.545 ;
        RECT 43.015 47.125 47.940 47.545 ;
        RECT 42.520 46.935 42.775 46.960 ;
        RECT 42.520 46.920 42.795 46.935 ;
        RECT 42.490 46.645 42.825 46.920 ;
        RECT 43.000 46.895 48.000 47.125 ;
        RECT 48.210 46.935 48.465 46.960 ;
        RECT 42.520 46.630 42.775 46.645 ;
        RECT 43.000 46.455 48.000 46.685 ;
        RECT 48.205 46.645 48.465 46.935 ;
        RECT 48.210 46.630 48.465 46.645 ;
        RECT 43.045 46.445 47.900 46.455 ;
        RECT 43.045 44.920 45.690 44.925 ;
        RECT 41.720 44.720 45.690 44.920 ;
        RECT 41.720 44.690 45.680 44.720 ;
        RECT 40.560 44.335 40.895 44.610 ;
        RECT 41.440 44.440 41.670 44.485 ;
        RECT 36.420 40.560 36.775 40.580 ;
        RECT 36.420 40.490 36.650 40.560 ;
        RECT 37.560 40.490 37.790 40.580 ;
        RECT 38.320 40.465 39.230 40.605 ;
        RECT 39.850 40.490 40.240 40.625 ;
        RECT 38.310 40.285 39.320 40.465 ;
        RECT 34.410 40.055 36.370 40.285 ;
        RECT 37.840 40.055 39.800 40.285 ;
        RECT 35.120 39.340 35.470 40.055 ;
        RECT 37.865 40.050 39.750 40.055 ;
        RECT 40.045 38.355 40.240 40.490 ;
        RECT 40.630 38.830 40.820 44.335 ;
        RECT 41.250 43.105 41.670 44.440 ;
        RECT 42.975 43.105 44.320 44.690 ;
        RECT 41.250 41.720 44.320 43.105 ;
        RECT 41.250 40.990 41.670 41.720 ;
        RECT 41.245 40.485 41.670 40.990 ;
        RECT 40.630 38.640 40.945 38.830 ;
        RECT 30.950 38.125 34.910 38.355 ;
        RECT 36.380 38.125 40.340 38.355 ;
        RECT 40.755 38.130 40.945 38.640 ;
        RECT 30.670 37.515 30.900 37.965 ;
        RECT 32.150 37.515 32.940 38.125 ;
        RECT 30.670 37.210 32.940 37.515 ;
        RECT 30.615 37.195 32.940 37.210 ;
        RECT 30.530 36.350 32.940 37.195 ;
        RECT 30.530 35.975 30.900 36.350 ;
        RECT 30.670 35.965 30.900 35.975 ;
        RECT 32.150 35.805 32.940 36.350 ;
        RECT 34.960 37.880 35.190 37.965 ;
        RECT 36.100 37.880 36.330 37.965 ;
        RECT 34.960 36.055 36.330 37.880 ;
        RECT 34.960 35.965 35.190 36.055 ;
        RECT 30.950 35.575 34.910 35.805 ;
        RECT 27.990 35.255 30.085 35.280 ;
        RECT 30.530 35.255 30.755 35.265 ;
        RECT 35.430 35.255 35.920 36.055 ;
        RECT 36.100 35.965 36.330 36.055 ;
        RECT 37.815 37.745 39.155 38.125 ;
        RECT 40.390 37.745 40.620 37.965 ;
        RECT 37.815 36.150 40.620 37.745 ;
        RECT 37.815 35.805 39.155 36.150 ;
        RECT 40.390 35.965 40.620 36.150 ;
        RECT 36.380 35.575 40.340 35.805 ;
        RECT 40.770 35.785 40.945 38.130 ;
        RECT 41.245 37.965 41.540 40.485 ;
        RECT 42.975 40.280 44.320 41.720 ;
        RECT 45.730 44.390 45.960 44.485 ;
        RECT 46.205 44.390 46.695 46.445 ;
        RECT 47.265 44.920 47.900 44.925 ;
        RECT 47.150 44.690 51.110 44.920 ;
        RECT 46.870 44.390 47.100 44.485 ;
        RECT 45.730 40.565 47.100 44.390 ;
        RECT 45.730 40.485 45.960 40.565 ;
        RECT 46.870 40.485 47.100 40.565 ;
        RECT 48.525 40.280 49.870 44.690 ;
        RECT 51.160 44.420 51.390 44.485 ;
        RECT 52.045 44.425 52.520 49.260 ;
        RECT 53.845 48.455 54.525 49.260 ;
        RECT 54.945 48.735 55.280 48.985 ;
        RECT 54.960 48.710 55.250 48.735 ;
        RECT 58.420 48.635 60.330 49.260 ;
        RECT 62.420 48.925 64.305 48.930 ;
        RECT 65.865 48.925 67.750 48.930 ;
        RECT 62.410 48.695 64.370 48.925 ;
        RECT 65.840 48.695 67.800 48.925 ;
        RECT 54.770 48.455 55.000 48.505 ;
        RECT 53.845 47.955 55.000 48.455 ;
        RECT 52.915 44.735 53.250 44.985 ;
        RECT 52.935 44.705 53.225 44.735 ;
        RECT 52.745 44.425 52.975 44.500 ;
        RECT 51.160 40.485 51.615 44.420 ;
        RECT 52.045 43.680 52.975 44.425 ;
        RECT 52.380 40.565 52.975 43.680 ;
        RECT 52.745 40.500 52.975 40.565 ;
        RECT 53.185 44.475 53.415 44.500 ;
        RECT 53.185 40.920 53.695 44.475 ;
        RECT 53.185 40.550 53.880 40.920 ;
        RECT 54.380 40.600 55.000 47.955 ;
        RECT 53.185 40.500 53.415 40.550 ;
        RECT 41.720 40.250 45.680 40.280 ;
        RECT 47.150 40.250 51.110 40.280 ;
        RECT 41.720 40.090 51.110 40.250 ;
        RECT 41.720 40.050 45.680 40.090 ;
        RECT 47.150 40.050 51.110 40.090 ;
        RECT 51.275 38.660 51.615 40.485 ;
        RECT 52.925 38.660 53.345 40.305 ;
        RECT 51.275 38.505 53.345 38.660 ;
        RECT 51.350 38.390 53.345 38.505 ;
        RECT 41.810 38.125 45.770 38.355 ;
        RECT 47.240 38.125 51.200 38.355 ;
        RECT 41.245 37.205 41.760 37.965 ;
        RECT 41.315 36.025 41.760 37.205 ;
        RECT 41.530 35.965 41.760 36.025 ;
        RECT 43.190 35.805 44.145 38.125 ;
        RECT 45.820 37.900 46.050 37.965 ;
        RECT 46.960 37.900 47.190 37.965 ;
        RECT 45.820 36.030 47.190 37.900 ;
        RECT 45.820 35.965 46.050 36.030 ;
        RECT 40.755 35.255 40.945 35.785 ;
        RECT 41.810 35.575 45.770 35.805 ;
        RECT 46.225 35.255 46.780 36.030 ;
        RECT 46.960 35.965 47.190 36.030 ;
        RECT 48.635 35.805 49.590 38.125 ;
        RECT 51.350 37.970 51.615 38.390 ;
        RECT 52.925 38.115 53.345 38.390 ;
        RECT 53.580 39.355 53.880 40.550 ;
        RECT 54.770 40.505 55.000 40.600 ;
        RECT 55.210 48.430 55.440 48.505 ;
        RECT 55.210 41.110 55.985 48.430 ;
        RECT 58.385 48.405 60.385 48.635 ;
        RECT 62.130 48.410 62.360 48.490 ;
        RECT 57.950 45.060 58.180 48.355 ;
        RECT 60.590 48.275 60.820 48.355 ;
        RECT 60.560 45.060 60.820 48.275 ;
        RECT 57.950 43.245 60.820 45.060 ;
        RECT 55.210 40.580 56.060 41.110 ;
        RECT 57.950 40.825 58.180 43.245 ;
        RECT 55.210 40.505 55.440 40.580 ;
        RECT 54.875 39.825 55.390 40.315 ;
        RECT 54.875 39.360 55.385 39.825 ;
        RECT 55.690 39.795 56.060 40.580 ;
        RECT 57.590 40.395 58.180 40.825 ;
        RECT 59.075 40.640 59.335 40.960 ;
        RECT 60.560 40.645 60.820 43.245 ;
        RECT 61.890 40.990 62.360 48.410 ;
        RECT 62.850 41.775 63.740 48.695 ;
        RECT 64.420 48.390 64.650 48.490 ;
        RECT 64.420 48.380 64.775 48.390 ;
        RECT 65.560 48.380 65.790 48.490 ;
        RECT 59.130 40.480 59.280 40.640 ;
        RECT 54.510 39.355 55.385 39.360 ;
        RECT 53.580 38.950 55.385 39.355 ;
        RECT 53.580 38.110 53.880 38.950 ;
        RECT 54.510 38.935 55.385 38.950 ;
        RECT 54.875 38.825 55.385 38.935 ;
        RECT 54.875 38.125 55.390 38.825 ;
        RECT 55.585 38.795 56.615 39.795 ;
        RECT 51.275 37.965 51.615 37.970 ;
        RECT 51.250 36.020 51.615 37.965 ;
        RECT 52.830 37.900 53.060 37.970 ;
        RECT 52.335 37.230 53.060 37.900 ;
        RECT 52.325 37.040 53.060 37.230 ;
        RECT 52.325 36.240 52.680 37.040 ;
        RECT 52.830 36.970 53.060 37.040 ;
        RECT 53.270 37.925 53.500 37.970 ;
        RECT 53.640 37.925 53.880 38.110 ;
        RECT 53.270 37.595 53.880 37.925 ;
        RECT 54.855 37.870 55.085 37.975 ;
        RECT 53.270 37.040 53.765 37.595 ;
        RECT 53.270 36.970 53.500 37.040 ;
        RECT 53.020 36.785 53.310 36.810 ;
        RECT 53.005 36.535 53.340 36.785 ;
        RECT 54.625 36.765 55.085 37.870 ;
        RECT 54.305 36.240 55.085 36.765 ;
        RECT 51.885 36.060 55.085 36.240 ;
        RECT 51.250 35.965 51.480 36.020 ;
        RECT 47.240 35.575 51.200 35.805 ;
        RECT 51.885 35.620 54.690 36.060 ;
        RECT 54.855 35.975 55.085 36.060 ;
        RECT 55.295 37.910 55.525 37.975 ;
        RECT 55.690 37.910 56.060 38.795 ;
        RECT 55.295 37.585 56.060 37.910 ;
        RECT 55.295 36.045 56.055 37.585 ;
        RECT 55.295 35.975 55.525 36.045 ;
        RECT 55.045 35.795 55.335 35.815 ;
        RECT 51.885 35.255 54.350 35.620 ;
        RECT 55.020 35.545 55.355 35.795 ;
        RECT 57.590 35.280 58.085 40.395 ;
        RECT 59.105 40.345 59.310 40.480 ;
        RECT 60.590 40.395 60.820 40.645 ;
        RECT 61.610 40.550 62.360 40.990 ;
        RECT 62.780 40.775 63.795 41.775 ;
        RECT 58.385 40.115 60.385 40.345 ;
        RECT 61.610 38.355 61.980 40.550 ;
        RECT 62.130 40.490 62.360 40.550 ;
        RECT 62.850 40.285 63.740 40.775 ;
        RECT 64.420 40.580 65.790 48.380 ;
        RECT 66.325 43.635 67.215 48.695 ;
        RECT 67.850 48.410 68.080 48.490 ;
        RECT 66.320 42.015 67.220 43.635 ;
        RECT 66.325 41.605 67.215 42.015 ;
        RECT 66.250 40.605 67.280 41.605 ;
        RECT 67.850 40.625 68.225 48.410 ;
        RECT 68.500 48.025 70.180 49.260 ;
        RECT 71.015 48.025 75.940 48.035 ;
        RECT 68.500 47.545 75.940 48.025 ;
        RECT 68.500 45.285 70.180 47.545 ;
        RECT 71.015 47.125 75.940 47.545 ;
        RECT 70.520 46.935 70.775 46.960 ;
        RECT 70.520 46.920 70.795 46.935 ;
        RECT 70.490 46.645 70.825 46.920 ;
        RECT 71.000 46.895 76.000 47.125 ;
        RECT 76.210 46.935 76.465 46.960 ;
        RECT 70.520 46.630 70.775 46.645 ;
        RECT 71.000 46.455 76.000 46.685 ;
        RECT 76.205 46.645 76.465 46.935 ;
        RECT 76.210 46.630 76.465 46.645 ;
        RECT 71.045 46.445 75.900 46.455 ;
        RECT 71.045 44.920 73.690 44.925 ;
        RECT 69.720 44.720 73.690 44.920 ;
        RECT 69.720 44.690 73.680 44.720 ;
        RECT 68.560 44.335 68.895 44.610 ;
        RECT 69.440 44.440 69.670 44.485 ;
        RECT 64.420 40.560 64.775 40.580 ;
        RECT 64.420 40.490 64.650 40.560 ;
        RECT 65.560 40.490 65.790 40.580 ;
        RECT 66.320 40.465 67.230 40.605 ;
        RECT 67.850 40.490 68.240 40.625 ;
        RECT 66.310 40.285 67.320 40.465 ;
        RECT 62.410 40.055 64.370 40.285 ;
        RECT 65.840 40.055 67.800 40.285 ;
        RECT 63.115 39.230 63.460 40.055 ;
        RECT 65.865 40.050 67.750 40.055 ;
        RECT 68.045 38.355 68.240 40.490 ;
        RECT 68.630 38.830 68.820 44.335 ;
        RECT 69.250 43.105 69.670 44.440 ;
        RECT 70.975 43.105 72.320 44.690 ;
        RECT 69.250 41.720 72.320 43.105 ;
        RECT 69.250 40.990 69.670 41.720 ;
        RECT 69.245 40.485 69.670 40.990 ;
        RECT 68.630 38.640 68.945 38.830 ;
        RECT 58.950 38.125 62.910 38.355 ;
        RECT 64.380 38.125 68.340 38.355 ;
        RECT 68.755 38.130 68.945 38.640 ;
        RECT 58.670 37.515 58.900 37.965 ;
        RECT 60.150 37.515 60.940 38.125 ;
        RECT 58.670 37.210 60.940 37.515 ;
        RECT 58.615 37.195 60.940 37.210 ;
        RECT 58.530 36.350 60.940 37.195 ;
        RECT 58.530 35.975 58.900 36.350 ;
        RECT 58.670 35.965 58.900 35.975 ;
        RECT 60.150 35.805 60.940 36.350 ;
        RECT 62.960 37.880 63.190 37.965 ;
        RECT 64.100 37.880 64.330 37.965 ;
        RECT 62.960 36.055 64.330 37.880 ;
        RECT 62.960 35.965 63.190 36.055 ;
        RECT 58.950 35.575 62.910 35.805 ;
        RECT 55.590 35.255 58.085 35.280 ;
        RECT 58.530 35.255 58.755 35.265 ;
        RECT 63.430 35.255 63.920 36.055 ;
        RECT 64.100 35.965 64.330 36.055 ;
        RECT 65.815 37.745 67.155 38.125 ;
        RECT 68.390 37.745 68.620 37.965 ;
        RECT 65.815 36.150 68.620 37.745 ;
        RECT 65.815 35.805 67.155 36.150 ;
        RECT 68.390 35.965 68.620 36.150 ;
        RECT 64.380 35.575 68.340 35.805 ;
        RECT 68.770 35.785 68.945 38.130 ;
        RECT 69.245 37.965 69.540 40.485 ;
        RECT 70.975 40.280 72.320 41.720 ;
        RECT 73.730 44.390 73.960 44.485 ;
        RECT 74.205 44.390 74.695 46.445 ;
        RECT 75.265 44.920 75.900 44.925 ;
        RECT 75.150 44.690 79.110 44.920 ;
        RECT 74.870 44.390 75.100 44.485 ;
        RECT 73.730 40.565 75.100 44.390 ;
        RECT 73.730 40.485 73.960 40.565 ;
        RECT 74.870 40.485 75.100 40.565 ;
        RECT 76.525 40.280 77.870 44.690 ;
        RECT 79.160 44.420 79.390 44.485 ;
        RECT 80.045 44.425 80.520 49.260 ;
        RECT 81.845 48.455 82.525 49.260 ;
        RECT 82.945 48.735 83.280 48.985 ;
        RECT 82.960 48.710 83.250 48.735 ;
        RECT 86.420 48.635 88.330 49.260 ;
        RECT 90.420 48.925 92.305 48.930 ;
        RECT 93.865 48.925 95.750 48.930 ;
        RECT 90.410 48.695 92.370 48.925 ;
        RECT 93.840 48.695 95.800 48.925 ;
        RECT 82.770 48.455 83.000 48.505 ;
        RECT 81.845 47.955 83.000 48.455 ;
        RECT 80.915 44.735 81.250 44.985 ;
        RECT 80.935 44.705 81.225 44.735 ;
        RECT 80.745 44.425 80.975 44.500 ;
        RECT 79.160 40.485 79.615 44.420 ;
        RECT 80.045 43.680 80.975 44.425 ;
        RECT 80.380 40.565 80.975 43.680 ;
        RECT 80.745 40.500 80.975 40.565 ;
        RECT 81.185 44.475 81.415 44.500 ;
        RECT 81.185 40.920 81.695 44.475 ;
        RECT 81.185 40.550 81.880 40.920 ;
        RECT 82.380 40.600 83.000 47.955 ;
        RECT 81.185 40.500 81.415 40.550 ;
        RECT 69.720 40.250 73.680 40.280 ;
        RECT 75.150 40.250 79.110 40.280 ;
        RECT 69.720 40.090 79.110 40.250 ;
        RECT 69.720 40.050 73.680 40.090 ;
        RECT 75.150 40.050 79.110 40.090 ;
        RECT 79.275 38.660 79.615 40.485 ;
        RECT 80.925 38.660 81.345 40.305 ;
        RECT 79.275 38.505 81.345 38.660 ;
        RECT 79.350 38.390 81.345 38.505 ;
        RECT 69.810 38.125 73.770 38.355 ;
        RECT 75.240 38.125 79.200 38.355 ;
        RECT 69.245 37.205 69.760 37.965 ;
        RECT 69.315 36.025 69.760 37.205 ;
        RECT 69.530 35.965 69.760 36.025 ;
        RECT 71.190 35.805 72.145 38.125 ;
        RECT 73.820 37.900 74.050 37.965 ;
        RECT 74.960 37.900 75.190 37.965 ;
        RECT 73.820 36.030 75.190 37.900 ;
        RECT 73.820 35.965 74.050 36.030 ;
        RECT 68.755 35.255 68.945 35.785 ;
        RECT 69.810 35.575 73.770 35.805 ;
        RECT 74.225 35.255 74.780 36.030 ;
        RECT 74.960 35.965 75.190 36.030 ;
        RECT 76.635 35.805 77.590 38.125 ;
        RECT 79.350 37.970 79.615 38.390 ;
        RECT 80.925 38.115 81.345 38.390 ;
        RECT 81.580 39.355 81.880 40.550 ;
        RECT 82.770 40.505 83.000 40.600 ;
        RECT 83.210 48.430 83.440 48.505 ;
        RECT 83.210 41.110 83.985 48.430 ;
        RECT 86.385 48.405 88.385 48.635 ;
        RECT 90.130 48.410 90.360 48.490 ;
        RECT 85.950 45.060 86.180 48.355 ;
        RECT 88.590 48.275 88.820 48.355 ;
        RECT 88.560 45.060 88.820 48.275 ;
        RECT 85.950 43.245 88.820 45.060 ;
        RECT 83.210 40.580 84.060 41.110 ;
        RECT 85.950 40.825 86.180 43.245 ;
        RECT 83.210 40.505 83.440 40.580 ;
        RECT 82.875 39.825 83.390 40.315 ;
        RECT 82.875 39.360 83.385 39.825 ;
        RECT 83.690 39.795 84.060 40.580 ;
        RECT 85.590 40.395 86.180 40.825 ;
        RECT 87.075 40.640 87.335 40.960 ;
        RECT 88.560 40.645 88.820 43.245 ;
        RECT 89.890 40.990 90.360 48.410 ;
        RECT 90.850 41.775 91.740 48.695 ;
        RECT 92.420 48.390 92.650 48.490 ;
        RECT 92.420 48.380 92.775 48.390 ;
        RECT 93.560 48.380 93.790 48.490 ;
        RECT 87.130 40.480 87.280 40.640 ;
        RECT 82.510 39.355 83.385 39.360 ;
        RECT 81.580 38.950 83.385 39.355 ;
        RECT 81.580 38.110 81.880 38.950 ;
        RECT 82.510 38.935 83.385 38.950 ;
        RECT 82.875 38.825 83.385 38.935 ;
        RECT 82.875 38.125 83.390 38.825 ;
        RECT 83.585 38.795 84.615 39.795 ;
        RECT 79.275 37.965 79.615 37.970 ;
        RECT 79.250 36.020 79.615 37.965 ;
        RECT 80.830 37.900 81.060 37.970 ;
        RECT 80.335 37.230 81.060 37.900 ;
        RECT 80.325 37.040 81.060 37.230 ;
        RECT 80.325 36.240 80.680 37.040 ;
        RECT 80.830 36.970 81.060 37.040 ;
        RECT 81.270 37.925 81.500 37.970 ;
        RECT 81.640 37.925 81.880 38.110 ;
        RECT 81.270 37.595 81.880 37.925 ;
        RECT 82.855 37.870 83.085 37.975 ;
        RECT 81.270 37.040 81.765 37.595 ;
        RECT 81.270 36.970 81.500 37.040 ;
        RECT 81.020 36.785 81.310 36.810 ;
        RECT 81.005 36.535 81.340 36.785 ;
        RECT 82.625 36.765 83.085 37.870 ;
        RECT 82.305 36.240 83.085 36.765 ;
        RECT 79.885 36.060 83.085 36.240 ;
        RECT 79.250 35.965 79.480 36.020 ;
        RECT 79.885 35.960 82.690 36.060 ;
        RECT 82.855 35.975 83.085 36.060 ;
        RECT 83.295 37.910 83.525 37.975 ;
        RECT 83.690 37.910 84.060 38.795 ;
        RECT 83.295 37.585 84.060 37.910 ;
        RECT 83.295 36.045 84.055 37.585 ;
        RECT 83.295 35.975 83.525 36.045 ;
        RECT 75.240 35.575 79.200 35.805 ;
        RECT 79.830 35.785 82.690 35.960 ;
        RECT 83.045 35.795 83.335 35.815 ;
        RECT 79.870 35.620 82.690 35.785 ;
        RECT 79.870 35.255 82.350 35.620 ;
        RECT 83.020 35.545 83.355 35.795 ;
        RECT 85.590 35.280 86.085 40.395 ;
        RECT 87.105 40.345 87.310 40.480 ;
        RECT 88.590 40.395 88.820 40.645 ;
        RECT 89.610 40.550 90.360 40.990 ;
        RECT 90.780 40.775 91.795 41.775 ;
        RECT 86.385 40.115 88.385 40.345 ;
        RECT 89.610 38.355 89.980 40.550 ;
        RECT 90.130 40.490 90.360 40.550 ;
        RECT 90.850 40.285 91.740 40.775 ;
        RECT 92.420 40.580 93.790 48.380 ;
        RECT 94.325 43.635 95.215 48.695 ;
        RECT 95.850 48.410 96.080 48.490 ;
        RECT 94.320 42.015 95.220 43.635 ;
        RECT 94.325 41.605 95.215 42.015 ;
        RECT 94.250 40.605 95.280 41.605 ;
        RECT 95.850 40.625 96.225 48.410 ;
        RECT 96.500 48.025 98.180 49.260 ;
        RECT 99.015 48.025 103.940 48.035 ;
        RECT 96.500 47.545 103.940 48.025 ;
        RECT 96.500 45.285 98.180 47.545 ;
        RECT 99.015 47.125 103.940 47.545 ;
        RECT 98.520 46.935 98.775 46.960 ;
        RECT 98.520 46.920 98.795 46.935 ;
        RECT 98.490 46.645 98.825 46.920 ;
        RECT 99.000 46.895 104.000 47.125 ;
        RECT 104.210 46.935 104.465 46.960 ;
        RECT 98.520 46.630 98.775 46.645 ;
        RECT 99.000 46.455 104.000 46.685 ;
        RECT 104.205 46.645 104.465 46.935 ;
        RECT 104.210 46.630 104.465 46.645 ;
        RECT 99.045 46.445 103.900 46.455 ;
        RECT 99.045 44.920 101.690 44.925 ;
        RECT 97.720 44.720 101.690 44.920 ;
        RECT 97.720 44.690 101.680 44.720 ;
        RECT 96.560 44.335 96.895 44.610 ;
        RECT 97.440 44.440 97.670 44.485 ;
        RECT 92.420 40.560 92.775 40.580 ;
        RECT 92.420 40.490 92.650 40.560 ;
        RECT 93.560 40.490 93.790 40.580 ;
        RECT 94.320 40.465 95.230 40.605 ;
        RECT 95.850 40.490 96.240 40.625 ;
        RECT 94.310 40.285 95.320 40.465 ;
        RECT 90.410 40.055 92.370 40.285 ;
        RECT 93.840 40.055 95.800 40.285 ;
        RECT 91.095 39.170 91.495 40.055 ;
        RECT 93.865 40.050 95.750 40.055 ;
        RECT 96.045 38.355 96.240 40.490 ;
        RECT 96.630 38.830 96.820 44.335 ;
        RECT 97.250 43.105 97.670 44.440 ;
        RECT 98.975 43.105 100.320 44.690 ;
        RECT 97.250 41.720 100.320 43.105 ;
        RECT 97.250 40.990 97.670 41.720 ;
        RECT 97.245 40.485 97.670 40.990 ;
        RECT 96.630 38.640 96.945 38.830 ;
        RECT 86.950 38.125 90.910 38.355 ;
        RECT 92.380 38.125 96.340 38.355 ;
        RECT 96.755 38.130 96.945 38.640 ;
        RECT 86.670 37.515 86.900 37.965 ;
        RECT 88.150 37.515 88.940 38.125 ;
        RECT 86.670 37.210 88.940 37.515 ;
        RECT 86.615 37.195 88.940 37.210 ;
        RECT 86.530 36.350 88.940 37.195 ;
        RECT 86.530 35.975 86.900 36.350 ;
        RECT 86.670 35.965 86.900 35.975 ;
        RECT 88.150 35.805 88.940 36.350 ;
        RECT 90.960 37.880 91.190 37.965 ;
        RECT 92.100 37.880 92.330 37.965 ;
        RECT 90.960 36.055 92.330 37.880 ;
        RECT 90.960 35.965 91.190 36.055 ;
        RECT 86.950 35.575 90.910 35.805 ;
        RECT 83.590 35.255 86.085 35.280 ;
        RECT 86.530 35.255 86.755 35.265 ;
        RECT 91.430 35.255 91.920 36.055 ;
        RECT 92.100 35.965 92.330 36.055 ;
        RECT 93.815 37.745 95.155 38.125 ;
        RECT 96.390 37.745 96.620 37.965 ;
        RECT 93.815 36.150 96.620 37.745 ;
        RECT 93.815 35.805 95.155 36.150 ;
        RECT 96.390 35.965 96.620 36.150 ;
        RECT 92.380 35.575 96.340 35.805 ;
        RECT 96.770 35.785 96.945 38.130 ;
        RECT 97.245 37.965 97.540 40.485 ;
        RECT 98.975 40.280 100.320 41.720 ;
        RECT 101.730 44.390 101.960 44.485 ;
        RECT 102.205 44.390 102.695 46.445 ;
        RECT 103.265 44.920 103.900 44.925 ;
        RECT 103.150 44.690 107.110 44.920 ;
        RECT 102.870 44.390 103.100 44.485 ;
        RECT 101.730 40.565 103.100 44.390 ;
        RECT 101.730 40.485 101.960 40.565 ;
        RECT 102.870 40.485 103.100 40.565 ;
        RECT 104.525 40.280 105.870 44.690 ;
        RECT 107.160 44.420 107.390 44.485 ;
        RECT 108.045 44.425 108.520 49.260 ;
        RECT 109.845 48.455 110.525 49.260 ;
        RECT 110.945 48.735 111.280 48.985 ;
        RECT 110.960 48.710 111.250 48.735 ;
        RECT 114.420 48.635 116.330 49.260 ;
        RECT 118.420 48.925 120.305 48.930 ;
        RECT 121.865 48.925 123.750 48.930 ;
        RECT 118.410 48.695 120.370 48.925 ;
        RECT 121.840 48.695 123.800 48.925 ;
        RECT 110.770 48.455 111.000 48.505 ;
        RECT 109.845 47.955 111.000 48.455 ;
        RECT 108.915 44.735 109.250 44.985 ;
        RECT 108.935 44.705 109.225 44.735 ;
        RECT 108.745 44.425 108.975 44.500 ;
        RECT 107.160 40.485 107.615 44.420 ;
        RECT 108.045 43.680 108.975 44.425 ;
        RECT 108.380 40.565 108.975 43.680 ;
        RECT 108.745 40.500 108.975 40.565 ;
        RECT 109.185 44.475 109.415 44.500 ;
        RECT 109.185 40.920 109.695 44.475 ;
        RECT 109.185 40.550 109.880 40.920 ;
        RECT 110.380 40.600 111.000 47.955 ;
        RECT 109.185 40.500 109.415 40.550 ;
        RECT 97.720 40.250 101.680 40.280 ;
        RECT 103.150 40.250 107.110 40.280 ;
        RECT 97.720 40.090 107.110 40.250 ;
        RECT 97.720 40.050 101.680 40.090 ;
        RECT 103.150 40.050 107.110 40.090 ;
        RECT 107.275 38.660 107.615 40.485 ;
        RECT 108.925 38.660 109.345 40.305 ;
        RECT 107.275 38.505 109.345 38.660 ;
        RECT 107.350 38.390 109.345 38.505 ;
        RECT 97.810 38.125 101.770 38.355 ;
        RECT 103.240 38.125 107.200 38.355 ;
        RECT 97.245 37.205 97.760 37.965 ;
        RECT 97.315 36.025 97.760 37.205 ;
        RECT 97.530 35.965 97.760 36.025 ;
        RECT 99.190 35.805 100.145 38.125 ;
        RECT 101.820 37.900 102.050 37.965 ;
        RECT 102.960 37.900 103.190 37.965 ;
        RECT 101.820 36.030 103.190 37.900 ;
        RECT 101.820 35.965 102.050 36.030 ;
        RECT 96.755 35.255 96.945 35.785 ;
        RECT 97.810 35.575 101.770 35.805 ;
        RECT 102.225 35.255 102.780 36.030 ;
        RECT 102.960 35.965 103.190 36.030 ;
        RECT 104.635 35.805 105.590 38.125 ;
        RECT 107.350 37.970 107.615 38.390 ;
        RECT 108.925 38.115 109.345 38.390 ;
        RECT 109.580 39.355 109.880 40.550 ;
        RECT 110.770 40.505 111.000 40.600 ;
        RECT 111.210 48.430 111.440 48.505 ;
        RECT 111.210 41.110 111.985 48.430 ;
        RECT 114.385 48.405 116.385 48.635 ;
        RECT 118.130 48.410 118.360 48.490 ;
        RECT 113.950 45.060 114.180 48.355 ;
        RECT 116.590 48.275 116.820 48.355 ;
        RECT 116.560 45.060 116.820 48.275 ;
        RECT 113.950 43.245 116.820 45.060 ;
        RECT 111.210 40.580 112.060 41.110 ;
        RECT 113.950 40.825 114.180 43.245 ;
        RECT 111.210 40.505 111.440 40.580 ;
        RECT 110.875 39.825 111.390 40.315 ;
        RECT 110.875 39.360 111.385 39.825 ;
        RECT 111.690 39.795 112.060 40.580 ;
        RECT 113.590 40.395 114.180 40.825 ;
        RECT 115.075 40.640 115.335 40.960 ;
        RECT 116.560 40.645 116.820 43.245 ;
        RECT 117.890 40.990 118.360 48.410 ;
        RECT 118.850 41.775 119.740 48.695 ;
        RECT 120.420 48.390 120.650 48.490 ;
        RECT 120.420 48.380 120.775 48.390 ;
        RECT 121.560 48.380 121.790 48.490 ;
        RECT 115.130 40.480 115.280 40.640 ;
        RECT 110.510 39.355 111.385 39.360 ;
        RECT 109.580 38.950 111.385 39.355 ;
        RECT 109.580 38.110 109.880 38.950 ;
        RECT 110.510 38.935 111.385 38.950 ;
        RECT 110.875 38.825 111.385 38.935 ;
        RECT 110.875 38.125 111.390 38.825 ;
        RECT 111.585 38.795 112.615 39.795 ;
        RECT 107.275 37.965 107.615 37.970 ;
        RECT 107.250 36.020 107.615 37.965 ;
        RECT 108.830 37.900 109.060 37.970 ;
        RECT 108.335 37.230 109.060 37.900 ;
        RECT 108.325 37.040 109.060 37.230 ;
        RECT 108.325 36.240 108.680 37.040 ;
        RECT 108.830 36.970 109.060 37.040 ;
        RECT 109.270 37.925 109.500 37.970 ;
        RECT 109.640 37.925 109.880 38.110 ;
        RECT 109.270 37.595 109.880 37.925 ;
        RECT 110.855 37.870 111.085 37.975 ;
        RECT 109.270 37.040 109.765 37.595 ;
        RECT 109.270 36.970 109.500 37.040 ;
        RECT 109.020 36.785 109.310 36.810 ;
        RECT 109.005 36.535 109.340 36.785 ;
        RECT 110.625 36.765 111.085 37.870 ;
        RECT 110.305 36.240 111.085 36.765 ;
        RECT 107.885 36.060 111.085 36.240 ;
        RECT 107.250 35.965 107.480 36.020 ;
        RECT 103.240 35.575 107.200 35.805 ;
        RECT 107.885 35.620 110.690 36.060 ;
        RECT 110.855 35.975 111.085 36.060 ;
        RECT 111.295 37.910 111.525 37.975 ;
        RECT 111.690 37.910 112.060 38.795 ;
        RECT 111.295 37.585 112.060 37.910 ;
        RECT 111.295 36.045 112.055 37.585 ;
        RECT 111.295 35.975 111.525 36.045 ;
        RECT 111.045 35.795 111.335 35.815 ;
        RECT 107.885 35.255 110.350 35.620 ;
        RECT 111.020 35.545 111.355 35.795 ;
        RECT 113.590 35.280 114.085 40.395 ;
        RECT 115.105 40.345 115.310 40.480 ;
        RECT 116.590 40.395 116.820 40.645 ;
        RECT 117.610 40.550 118.360 40.990 ;
        RECT 118.780 40.775 119.795 41.775 ;
        RECT 114.385 40.115 116.385 40.345 ;
        RECT 117.610 38.355 117.980 40.550 ;
        RECT 118.130 40.490 118.360 40.550 ;
        RECT 118.850 40.285 119.740 40.775 ;
        RECT 120.420 40.580 121.790 48.380 ;
        RECT 122.325 43.635 123.215 48.695 ;
        RECT 123.850 48.410 124.080 48.490 ;
        RECT 122.320 42.015 123.220 43.635 ;
        RECT 122.325 41.605 123.215 42.015 ;
        RECT 122.250 40.605 123.280 41.605 ;
        RECT 123.850 40.625 124.225 48.410 ;
        RECT 124.500 48.025 126.180 49.260 ;
        RECT 127.015 48.025 131.940 48.035 ;
        RECT 124.500 47.545 131.940 48.025 ;
        RECT 124.500 45.285 126.180 47.545 ;
        RECT 127.015 47.125 131.940 47.545 ;
        RECT 126.520 46.935 126.775 46.960 ;
        RECT 126.520 46.920 126.795 46.935 ;
        RECT 126.490 46.645 126.825 46.920 ;
        RECT 127.000 46.895 132.000 47.125 ;
        RECT 132.210 46.935 132.465 46.960 ;
        RECT 126.520 46.630 126.775 46.645 ;
        RECT 127.000 46.455 132.000 46.685 ;
        RECT 132.205 46.645 132.465 46.935 ;
        RECT 132.210 46.630 132.465 46.645 ;
        RECT 127.045 46.445 131.900 46.455 ;
        RECT 127.045 44.920 129.690 44.925 ;
        RECT 125.720 44.720 129.690 44.920 ;
        RECT 125.720 44.690 129.680 44.720 ;
        RECT 124.560 44.335 124.895 44.610 ;
        RECT 125.440 44.440 125.670 44.485 ;
        RECT 120.420 40.560 120.775 40.580 ;
        RECT 120.420 40.490 120.650 40.560 ;
        RECT 121.560 40.490 121.790 40.580 ;
        RECT 122.320 40.465 123.230 40.605 ;
        RECT 123.850 40.490 124.240 40.625 ;
        RECT 122.310 40.285 123.320 40.465 ;
        RECT 118.410 40.055 120.370 40.285 ;
        RECT 121.840 40.055 123.800 40.285 ;
        RECT 119.145 39.135 119.430 40.055 ;
        RECT 121.865 40.050 123.750 40.055 ;
        RECT 124.045 38.355 124.240 40.490 ;
        RECT 124.630 38.830 124.820 44.335 ;
        RECT 125.250 43.105 125.670 44.440 ;
        RECT 126.975 43.105 128.320 44.690 ;
        RECT 125.250 41.720 128.320 43.105 ;
        RECT 125.250 40.990 125.670 41.720 ;
        RECT 125.245 40.485 125.670 40.990 ;
        RECT 124.630 38.640 124.945 38.830 ;
        RECT 114.950 38.125 118.910 38.355 ;
        RECT 120.380 38.125 124.340 38.355 ;
        RECT 124.755 38.130 124.945 38.640 ;
        RECT 114.670 37.515 114.900 37.965 ;
        RECT 116.150 37.515 116.940 38.125 ;
        RECT 114.670 37.210 116.940 37.515 ;
        RECT 114.615 37.195 116.940 37.210 ;
        RECT 114.530 36.350 116.940 37.195 ;
        RECT 114.530 35.975 114.900 36.350 ;
        RECT 114.670 35.965 114.900 35.975 ;
        RECT 116.150 35.805 116.940 36.350 ;
        RECT 118.960 37.880 119.190 37.965 ;
        RECT 120.100 37.880 120.330 37.965 ;
        RECT 118.960 36.055 120.330 37.880 ;
        RECT 118.960 35.965 119.190 36.055 ;
        RECT 114.950 35.575 118.910 35.805 ;
        RECT 111.490 35.255 114.190 35.280 ;
        RECT 114.530 35.255 114.755 35.265 ;
        RECT 119.430 35.255 119.920 36.055 ;
        RECT 120.100 35.965 120.330 36.055 ;
        RECT 121.815 37.745 123.155 38.125 ;
        RECT 124.390 37.745 124.620 37.965 ;
        RECT 121.815 36.150 124.620 37.745 ;
        RECT 121.815 35.805 123.155 36.150 ;
        RECT 124.390 35.965 124.620 36.150 ;
        RECT 120.380 35.575 124.340 35.805 ;
        RECT 124.770 35.785 124.945 38.130 ;
        RECT 125.245 37.965 125.540 40.485 ;
        RECT 126.975 40.280 128.320 41.720 ;
        RECT 129.730 44.390 129.960 44.485 ;
        RECT 130.205 44.390 130.695 46.445 ;
        RECT 131.265 44.920 131.900 44.925 ;
        RECT 131.150 44.690 135.110 44.920 ;
        RECT 130.870 44.390 131.100 44.485 ;
        RECT 129.730 40.565 131.100 44.390 ;
        RECT 129.730 40.485 129.960 40.565 ;
        RECT 130.870 40.485 131.100 40.565 ;
        RECT 132.525 40.280 133.870 44.690 ;
        RECT 135.160 44.420 135.390 44.485 ;
        RECT 136.045 44.425 136.520 49.260 ;
        RECT 137.845 48.455 138.525 49.260 ;
        RECT 138.945 48.735 139.280 48.985 ;
        RECT 138.960 48.710 139.250 48.735 ;
        RECT 144.150 48.720 146.255 49.310 ;
        RECT 146.835 48.720 148.940 49.310 ;
        RECT 138.770 48.455 139.000 48.505 ;
        RECT 137.845 47.955 139.000 48.455 ;
        RECT 136.915 44.735 137.250 44.985 ;
        RECT 136.935 44.705 137.225 44.735 ;
        RECT 136.745 44.425 136.975 44.500 ;
        RECT 135.160 40.485 135.615 44.420 ;
        RECT 136.045 43.680 136.975 44.425 ;
        RECT 136.380 40.565 136.975 43.680 ;
        RECT 136.745 40.500 136.975 40.565 ;
        RECT 137.185 44.475 137.415 44.500 ;
        RECT 137.185 40.920 137.695 44.475 ;
        RECT 137.185 40.550 137.880 40.920 ;
        RECT 138.380 40.600 139.000 47.955 ;
        RECT 137.185 40.500 137.415 40.550 ;
        RECT 125.720 40.250 129.680 40.280 ;
        RECT 131.150 40.250 135.110 40.280 ;
        RECT 125.720 40.090 135.110 40.250 ;
        RECT 125.720 40.050 129.680 40.090 ;
        RECT 131.150 40.050 135.110 40.090 ;
        RECT 135.275 38.660 135.615 40.485 ;
        RECT 136.925 38.660 137.345 40.305 ;
        RECT 135.275 38.505 137.345 38.660 ;
        RECT 135.350 38.390 137.345 38.505 ;
        RECT 125.810 38.125 129.770 38.355 ;
        RECT 131.240 38.125 135.200 38.355 ;
        RECT 125.245 37.205 125.760 37.965 ;
        RECT 125.315 36.025 125.760 37.205 ;
        RECT 125.530 35.965 125.760 36.025 ;
        RECT 127.190 35.805 128.145 38.125 ;
        RECT 129.820 37.900 130.050 37.965 ;
        RECT 130.960 37.900 131.190 37.965 ;
        RECT 129.820 36.030 131.190 37.900 ;
        RECT 129.820 35.965 130.050 36.030 ;
        RECT 124.755 35.255 124.945 35.785 ;
        RECT 125.810 35.575 129.770 35.805 ;
        RECT 130.225 35.255 130.780 36.030 ;
        RECT 130.960 35.965 131.190 36.030 ;
        RECT 132.635 35.805 133.590 38.125 ;
        RECT 135.350 37.970 135.615 38.390 ;
        RECT 136.925 38.115 137.345 38.390 ;
        RECT 137.580 39.355 137.880 40.550 ;
        RECT 138.770 40.505 139.000 40.600 ;
        RECT 139.210 48.430 139.440 48.505 ;
        RECT 139.210 41.110 139.985 48.430 ;
        RECT 146.860 47.490 148.890 48.720 ;
        RECT 144.150 46.900 146.255 47.490 ;
        RECT 146.835 46.900 148.940 47.490 ;
        RECT 144.160 45.670 146.190 46.900 ;
        RECT 146.890 46.880 148.890 46.900 ;
        RECT 146.890 45.670 154.890 45.680 ;
        RECT 144.150 45.080 146.255 45.670 ;
        RECT 146.835 45.180 154.890 45.670 ;
        RECT 146.835 45.080 148.940 45.180 ;
        RECT 144.190 43.850 146.190 43.880 ;
        RECT 144.150 43.260 146.255 43.850 ;
        RECT 146.835 43.780 148.940 43.850 ;
        RECT 149.425 43.780 149.925 44.125 ;
        RECT 152.890 43.850 154.890 45.180 ;
        RECT 150.130 43.780 152.235 43.850 ;
        RECT 146.835 43.280 152.235 43.780 ;
        RECT 146.835 43.260 148.940 43.280 ;
        RECT 150.130 43.260 152.235 43.280 ;
        RECT 152.815 43.260 154.920 43.850 ;
        RECT 144.190 42.945 146.190 43.260 ;
        RECT 141.790 42.505 146.190 42.945 ;
        RECT 144.190 42.030 146.190 42.505 ;
        RECT 144.150 41.440 146.255 42.030 ;
        RECT 146.835 41.980 148.940 42.030 ;
        RECT 150.130 41.980 152.235 42.030 ;
        RECT 146.835 41.480 152.235 41.980 ;
        RECT 146.835 41.440 148.940 41.480 ;
        RECT 149.530 41.440 152.235 41.480 ;
        RECT 152.815 41.440 154.920 42.030 ;
        RECT 149.530 41.240 150.310 41.440 ;
        RECT 139.210 40.580 140.060 41.110 ;
        RECT 149.530 41.035 150.030 41.240 ;
        RECT 139.210 40.505 139.440 40.580 ;
        RECT 138.875 39.825 139.390 40.315 ;
        RECT 138.875 39.360 139.385 39.825 ;
        RECT 139.690 39.795 140.060 40.580 ;
        RECT 142.350 40.535 150.030 41.035 ;
        RECT 153.565 40.995 154.355 41.440 ;
        RECT 150.785 40.205 154.355 40.995 ;
        RECT 150.785 40.055 151.575 40.205 ;
        RECT 138.510 39.355 139.385 39.360 ;
        RECT 137.580 38.950 139.385 39.355 ;
        RECT 137.580 38.110 137.880 38.950 ;
        RECT 138.510 38.935 139.385 38.950 ;
        RECT 138.875 38.825 139.385 38.935 ;
        RECT 138.875 38.125 139.390 38.825 ;
        RECT 139.585 38.795 140.615 39.795 ;
        RECT 141.105 39.265 151.575 40.055 ;
        RECT 135.275 37.965 135.615 37.970 ;
        RECT 135.250 36.020 135.615 37.965 ;
        RECT 136.830 37.900 137.060 37.970 ;
        RECT 136.335 37.230 137.060 37.900 ;
        RECT 136.325 37.040 137.060 37.230 ;
        RECT 136.325 36.240 136.680 37.040 ;
        RECT 136.830 36.970 137.060 37.040 ;
        RECT 137.270 37.925 137.500 37.970 ;
        RECT 137.640 37.925 137.880 38.110 ;
        RECT 137.270 37.595 137.880 37.925 ;
        RECT 138.855 37.870 139.085 37.975 ;
        RECT 137.270 37.040 137.765 37.595 ;
        RECT 137.270 36.970 137.500 37.040 ;
        RECT 137.020 36.785 137.310 36.810 ;
        RECT 137.005 36.535 137.340 36.785 ;
        RECT 138.625 36.765 139.085 37.870 ;
        RECT 138.305 36.240 139.085 36.765 ;
        RECT 135.885 36.060 139.085 36.240 ;
        RECT 135.250 35.965 135.480 36.020 ;
        RECT 131.240 35.575 135.200 35.805 ;
        RECT 135.885 35.620 138.690 36.060 ;
        RECT 138.855 35.975 139.085 36.060 ;
        RECT 139.295 37.910 139.525 37.975 ;
        RECT 139.690 37.910 140.060 38.795 ;
        RECT 139.295 37.585 140.060 37.910 ;
        RECT 139.295 36.045 140.055 37.585 ;
        RECT 139.295 35.975 139.525 36.045 ;
        RECT 139.045 35.795 139.335 35.815 ;
        RECT 135.885 35.335 138.350 35.620 ;
        RECT 139.020 35.545 139.355 35.795 ;
        RECT 141.105 35.335 141.895 39.265 ;
        RECT 135.885 35.255 141.895 35.335 ;
        RECT 1.475 34.545 141.895 35.255 ;
        RECT 1.475 34.380 140.080 34.545 ;
        RECT 27.790 33.960 30.490 33.980 ;
        RECT 55.390 33.960 57.990 33.980 ;
        RECT 83.390 33.960 86.290 33.980 ;
        RECT 111.190 33.960 114.190 33.980 ;
        RECT 1.450 33.280 139.925 33.960 ;
        RECT 1.450 33.260 27.925 33.280 ;
        RECT 29.450 33.260 83.925 33.280 ;
        RECT 85.450 33.260 111.925 33.280 ;
        RECT 113.450 33.260 139.925 33.280 ;
        RECT 2.420 32.635 4.330 33.260 ;
        RECT 6.420 32.925 8.305 32.930 ;
        RECT 9.865 32.925 11.750 32.930 ;
        RECT 6.410 32.695 8.370 32.925 ;
        RECT 9.840 32.695 11.800 32.925 ;
        RECT 2.385 32.405 4.385 32.635 ;
        RECT 6.130 32.410 6.360 32.490 ;
        RECT 1.950 29.060 2.180 32.355 ;
        RECT 4.590 32.275 4.820 32.355 ;
        RECT 4.560 29.060 4.820 32.275 ;
        RECT 1.950 27.245 4.820 29.060 ;
        RECT 1.950 24.825 2.180 27.245 ;
        RECT 1.590 24.395 2.180 24.825 ;
        RECT 3.075 24.640 3.335 24.960 ;
        RECT 4.560 24.645 4.820 27.245 ;
        RECT 5.890 24.990 6.360 32.410 ;
        RECT 6.850 25.775 7.740 32.695 ;
        RECT 8.420 32.390 8.650 32.490 ;
        RECT 8.420 32.380 8.775 32.390 ;
        RECT 9.560 32.380 9.790 32.490 ;
        RECT 3.130 24.480 3.280 24.640 ;
        RECT 1.590 19.255 2.085 24.395 ;
        RECT 3.105 24.345 3.310 24.480 ;
        RECT 4.590 24.395 4.820 24.645 ;
        RECT 5.610 24.550 6.360 24.990 ;
        RECT 6.780 24.775 7.795 25.775 ;
        RECT 2.385 24.115 4.385 24.345 ;
        RECT 5.610 22.355 5.980 24.550 ;
        RECT 6.130 24.490 6.360 24.550 ;
        RECT 6.850 24.285 7.740 24.775 ;
        RECT 8.420 24.580 9.790 32.380 ;
        RECT 10.325 27.635 11.215 32.695 ;
        RECT 11.850 32.410 12.080 32.490 ;
        RECT 10.320 26.015 11.220 27.635 ;
        RECT 10.325 25.605 11.215 26.015 ;
        RECT 10.250 24.605 11.280 25.605 ;
        RECT 11.850 24.625 12.225 32.410 ;
        RECT 12.500 32.025 14.180 33.260 ;
        RECT 15.015 32.025 19.940 32.035 ;
        RECT 12.500 31.545 19.940 32.025 ;
        RECT 12.500 29.285 14.180 31.545 ;
        RECT 15.015 31.125 19.940 31.545 ;
        RECT 14.520 30.935 14.775 30.960 ;
        RECT 14.520 30.920 14.795 30.935 ;
        RECT 14.490 30.645 14.825 30.920 ;
        RECT 15.000 30.895 20.000 31.125 ;
        RECT 20.210 30.935 20.465 30.960 ;
        RECT 14.520 30.630 14.775 30.645 ;
        RECT 15.000 30.455 20.000 30.685 ;
        RECT 20.205 30.645 20.465 30.935 ;
        RECT 20.210 30.630 20.465 30.645 ;
        RECT 15.045 30.445 19.900 30.455 ;
        RECT 15.045 28.920 17.690 28.925 ;
        RECT 13.720 28.720 17.690 28.920 ;
        RECT 13.720 28.690 17.680 28.720 ;
        RECT 12.560 28.335 12.895 28.610 ;
        RECT 13.440 28.440 13.670 28.485 ;
        RECT 8.420 24.560 8.775 24.580 ;
        RECT 8.420 24.490 8.650 24.560 ;
        RECT 9.560 24.490 9.790 24.580 ;
        RECT 10.320 24.465 11.230 24.605 ;
        RECT 11.850 24.490 12.240 24.625 ;
        RECT 10.310 24.285 11.320 24.465 ;
        RECT 6.410 24.055 8.370 24.285 ;
        RECT 9.840 24.055 11.800 24.285 ;
        RECT 7.165 23.035 7.495 24.055 ;
        RECT 9.865 24.050 11.750 24.055 ;
        RECT 12.045 22.355 12.240 24.490 ;
        RECT 12.630 22.830 12.820 28.335 ;
        RECT 13.250 27.105 13.670 28.440 ;
        RECT 14.975 27.105 16.320 28.690 ;
        RECT 13.250 25.720 16.320 27.105 ;
        RECT 13.250 24.990 13.670 25.720 ;
        RECT 13.245 24.485 13.670 24.990 ;
        RECT 12.630 22.640 12.945 22.830 ;
        RECT 2.950 22.125 6.910 22.355 ;
        RECT 8.380 22.125 12.340 22.355 ;
        RECT 12.755 22.130 12.945 22.640 ;
        RECT 2.670 21.515 2.900 21.965 ;
        RECT 4.150 21.515 4.940 22.125 ;
        RECT 2.670 21.210 4.940 21.515 ;
        RECT 2.615 21.195 4.940 21.210 ;
        RECT 2.530 20.350 4.940 21.195 ;
        RECT 2.530 19.975 2.900 20.350 ;
        RECT 2.670 19.965 2.900 19.975 ;
        RECT 4.150 19.805 4.940 20.350 ;
        RECT 6.960 21.880 7.190 21.965 ;
        RECT 8.100 21.880 8.330 21.965 ;
        RECT 6.960 20.055 8.330 21.880 ;
        RECT 6.960 19.965 7.190 20.055 ;
        RECT 2.950 19.575 6.910 19.805 ;
        RECT 2.530 19.255 2.755 19.265 ;
        RECT 7.430 19.255 7.920 20.055 ;
        RECT 8.100 19.965 8.330 20.055 ;
        RECT 9.815 21.745 11.155 22.125 ;
        RECT 12.390 21.745 12.620 21.965 ;
        RECT 9.815 20.150 12.620 21.745 ;
        RECT 9.815 19.805 11.155 20.150 ;
        RECT 12.390 19.965 12.620 20.150 ;
        RECT 8.380 19.575 12.340 19.805 ;
        RECT 12.770 19.785 12.945 22.130 ;
        RECT 13.245 21.965 13.540 24.485 ;
        RECT 14.975 24.280 16.320 25.720 ;
        RECT 17.730 28.390 17.960 28.485 ;
        RECT 18.205 28.390 18.695 30.445 ;
        RECT 19.265 28.920 19.900 28.925 ;
        RECT 19.150 28.690 23.110 28.920 ;
        RECT 18.870 28.390 19.100 28.485 ;
        RECT 17.730 24.565 19.100 28.390 ;
        RECT 17.730 24.485 17.960 24.565 ;
        RECT 18.870 24.485 19.100 24.565 ;
        RECT 20.525 24.280 21.870 28.690 ;
        RECT 23.160 28.420 23.390 28.485 ;
        RECT 24.045 28.425 24.520 33.260 ;
        RECT 25.845 32.455 26.525 33.260 ;
        RECT 26.945 32.735 27.280 32.985 ;
        RECT 26.960 32.710 27.250 32.735 ;
        RECT 30.420 32.635 32.330 33.260 ;
        RECT 34.420 32.925 36.305 32.930 ;
        RECT 37.865 32.925 39.750 32.930 ;
        RECT 34.410 32.695 36.370 32.925 ;
        RECT 37.840 32.695 39.800 32.925 ;
        RECT 26.770 32.455 27.000 32.505 ;
        RECT 25.845 31.955 27.000 32.455 ;
        RECT 24.915 28.735 25.250 28.985 ;
        RECT 24.935 28.705 25.225 28.735 ;
        RECT 24.745 28.425 24.975 28.500 ;
        RECT 23.160 24.485 23.615 28.420 ;
        RECT 24.045 27.680 24.975 28.425 ;
        RECT 24.380 24.565 24.975 27.680 ;
        RECT 24.745 24.500 24.975 24.565 ;
        RECT 25.185 28.475 25.415 28.500 ;
        RECT 25.185 24.920 25.695 28.475 ;
        RECT 25.185 24.550 25.880 24.920 ;
        RECT 26.380 24.600 27.000 31.955 ;
        RECT 25.185 24.500 25.415 24.550 ;
        RECT 13.720 24.250 17.680 24.280 ;
        RECT 19.150 24.250 23.110 24.280 ;
        RECT 13.720 24.090 23.110 24.250 ;
        RECT 13.720 24.050 17.680 24.090 ;
        RECT 19.150 24.050 23.110 24.090 ;
        RECT 23.275 22.660 23.615 24.485 ;
        RECT 24.925 22.660 25.345 24.305 ;
        RECT 23.275 22.505 25.345 22.660 ;
        RECT 23.350 22.390 25.345 22.505 ;
        RECT 13.810 22.125 17.770 22.355 ;
        RECT 19.240 22.125 23.200 22.355 ;
        RECT 13.245 21.205 13.760 21.965 ;
        RECT 13.315 20.025 13.760 21.205 ;
        RECT 13.530 19.965 13.760 20.025 ;
        RECT 15.190 19.805 16.145 22.125 ;
        RECT 17.820 21.900 18.050 21.965 ;
        RECT 18.960 21.900 19.190 21.965 ;
        RECT 17.820 20.030 19.190 21.900 ;
        RECT 17.820 19.965 18.050 20.030 ;
        RECT 12.755 19.255 12.945 19.785 ;
        RECT 13.810 19.575 17.770 19.805 ;
        RECT 18.225 19.255 18.780 20.030 ;
        RECT 18.960 19.965 19.190 20.030 ;
        RECT 20.635 19.805 21.590 22.125 ;
        RECT 23.350 21.970 23.615 22.390 ;
        RECT 24.925 22.115 25.345 22.390 ;
        RECT 25.580 23.355 25.880 24.550 ;
        RECT 26.770 24.505 27.000 24.600 ;
        RECT 27.210 32.430 27.440 32.505 ;
        RECT 27.210 25.110 27.985 32.430 ;
        RECT 30.385 32.405 32.385 32.635 ;
        RECT 34.130 32.410 34.360 32.490 ;
        RECT 29.950 29.060 30.180 32.355 ;
        RECT 32.590 32.275 32.820 32.355 ;
        RECT 32.560 29.060 32.820 32.275 ;
        RECT 29.950 27.245 32.820 29.060 ;
        RECT 27.210 24.580 28.060 25.110 ;
        RECT 29.950 24.825 30.180 27.245 ;
        RECT 27.210 24.505 27.440 24.580 ;
        RECT 26.875 23.825 27.390 24.315 ;
        RECT 27.690 23.825 28.060 24.580 ;
        RECT 29.590 24.395 30.180 24.825 ;
        RECT 31.075 24.640 31.335 24.960 ;
        RECT 32.560 24.645 32.820 27.245 ;
        RECT 33.890 24.990 34.360 32.410 ;
        RECT 34.850 25.775 35.740 32.695 ;
        RECT 36.420 32.390 36.650 32.490 ;
        RECT 36.420 32.380 36.775 32.390 ;
        RECT 37.560 32.380 37.790 32.490 ;
        RECT 31.130 24.480 31.280 24.640 ;
        RECT 26.875 23.360 27.385 23.825 ;
        RECT 26.510 23.355 27.385 23.360 ;
        RECT 25.580 22.950 27.385 23.355 ;
        RECT 25.580 22.110 25.880 22.950 ;
        RECT 26.510 22.935 27.385 22.950 ;
        RECT 26.875 22.825 27.385 22.935 ;
        RECT 26.875 22.125 27.390 22.825 ;
        RECT 27.615 22.795 28.615 23.825 ;
        RECT 23.275 21.965 23.615 21.970 ;
        RECT 23.250 20.020 23.615 21.965 ;
        RECT 24.830 21.900 25.060 21.970 ;
        RECT 24.335 21.230 25.060 21.900 ;
        RECT 24.325 21.040 25.060 21.230 ;
        RECT 24.325 20.240 24.680 21.040 ;
        RECT 24.830 20.970 25.060 21.040 ;
        RECT 25.270 21.925 25.500 21.970 ;
        RECT 25.640 21.925 25.880 22.110 ;
        RECT 25.270 21.595 25.880 21.925 ;
        RECT 26.855 21.870 27.085 21.975 ;
        RECT 25.270 21.040 25.765 21.595 ;
        RECT 25.270 20.970 25.500 21.040 ;
        RECT 25.020 20.785 25.310 20.810 ;
        RECT 25.005 20.535 25.340 20.785 ;
        RECT 26.625 20.765 27.085 21.870 ;
        RECT 26.305 20.240 27.085 20.765 ;
        RECT 23.885 20.060 27.085 20.240 ;
        RECT 23.250 19.965 23.480 20.020 ;
        RECT 19.240 19.575 23.200 19.805 ;
        RECT 23.885 19.620 26.690 20.060 ;
        RECT 26.855 19.975 27.085 20.060 ;
        RECT 27.295 21.910 27.525 21.975 ;
        RECT 27.690 21.910 28.060 22.795 ;
        RECT 27.295 21.585 28.060 21.910 ;
        RECT 27.295 20.045 28.055 21.585 ;
        RECT 27.295 19.975 27.525 20.045 ;
        RECT 27.045 19.795 27.335 19.815 ;
        RECT 23.885 19.255 26.350 19.620 ;
        RECT 27.020 19.545 27.355 19.795 ;
        RECT 29.590 19.280 30.085 24.395 ;
        RECT 31.105 24.345 31.310 24.480 ;
        RECT 32.590 24.395 32.820 24.645 ;
        RECT 33.610 24.550 34.360 24.990 ;
        RECT 34.780 24.775 35.795 25.775 ;
        RECT 30.385 24.115 32.385 24.345 ;
        RECT 33.610 22.355 33.980 24.550 ;
        RECT 34.130 24.490 34.360 24.550 ;
        RECT 34.850 24.285 35.740 24.775 ;
        RECT 36.420 24.580 37.790 32.380 ;
        RECT 38.325 27.635 39.215 32.695 ;
        RECT 39.850 32.410 40.080 32.490 ;
        RECT 38.320 26.015 39.220 27.635 ;
        RECT 38.325 25.605 39.215 26.015 ;
        RECT 38.250 24.605 39.280 25.605 ;
        RECT 39.850 24.625 40.225 32.410 ;
        RECT 40.500 32.025 42.180 33.260 ;
        RECT 43.015 32.025 47.940 32.035 ;
        RECT 40.500 31.545 47.940 32.025 ;
        RECT 40.500 29.285 42.180 31.545 ;
        RECT 43.015 31.125 47.940 31.545 ;
        RECT 42.520 30.935 42.775 30.960 ;
        RECT 42.520 30.920 42.795 30.935 ;
        RECT 42.490 30.645 42.825 30.920 ;
        RECT 43.000 30.895 48.000 31.125 ;
        RECT 48.210 30.935 48.465 30.960 ;
        RECT 42.520 30.630 42.775 30.645 ;
        RECT 43.000 30.455 48.000 30.685 ;
        RECT 48.205 30.645 48.465 30.935 ;
        RECT 48.210 30.630 48.465 30.645 ;
        RECT 43.045 30.445 47.900 30.455 ;
        RECT 43.045 28.920 45.690 28.925 ;
        RECT 41.720 28.720 45.690 28.920 ;
        RECT 41.720 28.690 45.680 28.720 ;
        RECT 40.560 28.335 40.895 28.610 ;
        RECT 41.440 28.440 41.670 28.485 ;
        RECT 36.420 24.560 36.775 24.580 ;
        RECT 36.420 24.490 36.650 24.560 ;
        RECT 37.560 24.490 37.790 24.580 ;
        RECT 38.320 24.465 39.230 24.605 ;
        RECT 39.850 24.490 40.240 24.625 ;
        RECT 38.310 24.285 39.320 24.465 ;
        RECT 34.410 24.055 36.370 24.285 ;
        RECT 37.840 24.055 39.800 24.285 ;
        RECT 35.115 23.005 35.465 24.055 ;
        RECT 37.865 24.050 39.750 24.055 ;
        RECT 40.045 22.355 40.240 24.490 ;
        RECT 40.630 22.830 40.820 28.335 ;
        RECT 41.250 27.105 41.670 28.440 ;
        RECT 42.975 27.105 44.320 28.690 ;
        RECT 41.250 25.720 44.320 27.105 ;
        RECT 41.250 24.990 41.670 25.720 ;
        RECT 41.245 24.485 41.670 24.990 ;
        RECT 40.630 22.640 40.945 22.830 ;
        RECT 30.950 22.125 34.910 22.355 ;
        RECT 36.380 22.125 40.340 22.355 ;
        RECT 40.755 22.130 40.945 22.640 ;
        RECT 30.670 21.515 30.900 21.965 ;
        RECT 32.150 21.515 32.940 22.125 ;
        RECT 30.670 21.210 32.940 21.515 ;
        RECT 30.615 21.195 32.940 21.210 ;
        RECT 30.530 20.350 32.940 21.195 ;
        RECT 30.530 19.975 30.900 20.350 ;
        RECT 30.670 19.965 30.900 19.975 ;
        RECT 32.150 19.805 32.940 20.350 ;
        RECT 34.960 21.880 35.190 21.965 ;
        RECT 36.100 21.880 36.330 21.965 ;
        RECT 34.960 20.055 36.330 21.880 ;
        RECT 34.960 19.965 35.190 20.055 ;
        RECT 30.950 19.575 34.910 19.805 ;
        RECT 27.890 19.255 30.085 19.280 ;
        RECT 30.530 19.255 30.755 19.265 ;
        RECT 35.430 19.255 35.920 20.055 ;
        RECT 36.100 19.965 36.330 20.055 ;
        RECT 37.815 21.745 39.155 22.125 ;
        RECT 40.390 21.745 40.620 21.965 ;
        RECT 37.815 20.150 40.620 21.745 ;
        RECT 37.815 19.805 39.155 20.150 ;
        RECT 40.390 19.965 40.620 20.150 ;
        RECT 36.380 19.575 40.340 19.805 ;
        RECT 40.770 19.785 40.945 22.130 ;
        RECT 41.245 21.965 41.540 24.485 ;
        RECT 42.975 24.280 44.320 25.720 ;
        RECT 45.730 28.390 45.960 28.485 ;
        RECT 46.205 28.390 46.695 30.445 ;
        RECT 47.265 28.920 47.900 28.925 ;
        RECT 47.150 28.690 51.110 28.920 ;
        RECT 46.870 28.390 47.100 28.485 ;
        RECT 45.730 24.565 47.100 28.390 ;
        RECT 45.730 24.485 45.960 24.565 ;
        RECT 46.870 24.485 47.100 24.565 ;
        RECT 48.525 24.280 49.870 28.690 ;
        RECT 51.160 28.420 51.390 28.485 ;
        RECT 52.045 28.425 52.520 33.260 ;
        RECT 53.845 32.455 54.525 33.260 ;
        RECT 55.390 33.180 57.990 33.260 ;
        RECT 54.945 32.735 55.280 32.985 ;
        RECT 54.960 32.710 55.250 32.735 ;
        RECT 58.420 32.635 60.330 33.260 ;
        RECT 62.420 32.925 64.305 32.930 ;
        RECT 65.865 32.925 67.750 32.930 ;
        RECT 62.410 32.695 64.370 32.925 ;
        RECT 65.840 32.695 67.800 32.925 ;
        RECT 54.770 32.455 55.000 32.505 ;
        RECT 53.845 31.955 55.000 32.455 ;
        RECT 52.915 28.735 53.250 28.985 ;
        RECT 52.935 28.705 53.225 28.735 ;
        RECT 52.745 28.425 52.975 28.500 ;
        RECT 51.160 24.485 51.615 28.420 ;
        RECT 52.045 27.680 52.975 28.425 ;
        RECT 52.380 24.565 52.975 27.680 ;
        RECT 52.745 24.500 52.975 24.565 ;
        RECT 53.185 28.475 53.415 28.500 ;
        RECT 53.185 24.920 53.695 28.475 ;
        RECT 53.185 24.550 53.880 24.920 ;
        RECT 54.380 24.600 55.000 31.955 ;
        RECT 53.185 24.500 53.415 24.550 ;
        RECT 41.720 24.250 45.680 24.280 ;
        RECT 47.150 24.250 51.110 24.280 ;
        RECT 41.720 24.090 51.110 24.250 ;
        RECT 41.720 24.050 45.680 24.090 ;
        RECT 47.150 24.050 51.110 24.090 ;
        RECT 51.275 22.660 51.615 24.485 ;
        RECT 52.925 22.660 53.345 24.305 ;
        RECT 51.275 22.505 53.345 22.660 ;
        RECT 51.350 22.390 53.345 22.505 ;
        RECT 41.810 22.125 45.770 22.355 ;
        RECT 47.240 22.125 51.200 22.355 ;
        RECT 41.245 21.205 41.760 21.965 ;
        RECT 41.315 20.025 41.760 21.205 ;
        RECT 41.530 19.965 41.760 20.025 ;
        RECT 43.190 19.805 44.145 22.125 ;
        RECT 45.820 21.900 46.050 21.965 ;
        RECT 46.960 21.900 47.190 21.965 ;
        RECT 45.820 20.030 47.190 21.900 ;
        RECT 45.820 19.965 46.050 20.030 ;
        RECT 40.755 19.255 40.945 19.785 ;
        RECT 41.810 19.575 45.770 19.805 ;
        RECT 46.225 19.255 46.780 20.030 ;
        RECT 46.960 19.965 47.190 20.030 ;
        RECT 48.635 19.805 49.590 22.125 ;
        RECT 51.350 21.970 51.615 22.390 ;
        RECT 52.925 22.115 53.345 22.390 ;
        RECT 53.580 23.355 53.880 24.550 ;
        RECT 54.770 24.505 55.000 24.600 ;
        RECT 55.210 32.430 55.440 32.505 ;
        RECT 55.210 25.110 55.985 32.430 ;
        RECT 58.385 32.405 60.385 32.635 ;
        RECT 62.130 32.410 62.360 32.490 ;
        RECT 57.950 29.060 58.180 32.355 ;
        RECT 60.590 32.275 60.820 32.355 ;
        RECT 60.560 29.060 60.820 32.275 ;
        RECT 57.950 27.245 60.820 29.060 ;
        RECT 55.210 24.580 56.060 25.110 ;
        RECT 57.950 24.825 58.180 27.245 ;
        RECT 55.210 24.505 55.440 24.580 ;
        RECT 54.875 23.825 55.390 24.315 ;
        RECT 54.875 23.360 55.385 23.825 ;
        RECT 55.690 23.795 56.060 24.580 ;
        RECT 57.590 24.395 58.180 24.825 ;
        RECT 59.075 24.640 59.335 24.960 ;
        RECT 60.560 24.645 60.820 27.245 ;
        RECT 61.890 24.990 62.360 32.410 ;
        RECT 62.850 25.775 63.740 32.695 ;
        RECT 64.420 32.390 64.650 32.490 ;
        RECT 64.420 32.380 64.775 32.390 ;
        RECT 65.560 32.380 65.790 32.490 ;
        RECT 59.130 24.480 59.280 24.640 ;
        RECT 54.510 23.355 55.385 23.360 ;
        RECT 53.580 22.950 55.385 23.355 ;
        RECT 53.580 22.110 53.880 22.950 ;
        RECT 54.510 22.935 55.385 22.950 ;
        RECT 54.875 22.825 55.385 22.935 ;
        RECT 54.875 22.125 55.390 22.825 ;
        RECT 55.585 22.795 56.615 23.795 ;
        RECT 51.275 21.965 51.615 21.970 ;
        RECT 51.250 20.020 51.615 21.965 ;
        RECT 52.830 21.900 53.060 21.970 ;
        RECT 52.335 21.230 53.060 21.900 ;
        RECT 52.325 21.040 53.060 21.230 ;
        RECT 52.325 20.240 52.680 21.040 ;
        RECT 52.830 20.970 53.060 21.040 ;
        RECT 53.270 21.925 53.500 21.970 ;
        RECT 53.640 21.925 53.880 22.110 ;
        RECT 53.270 21.595 53.880 21.925 ;
        RECT 54.855 21.870 55.085 21.975 ;
        RECT 53.270 21.040 53.765 21.595 ;
        RECT 53.270 20.970 53.500 21.040 ;
        RECT 53.020 20.785 53.310 20.810 ;
        RECT 53.005 20.535 53.340 20.785 ;
        RECT 54.625 20.765 55.085 21.870 ;
        RECT 54.305 20.240 55.085 20.765 ;
        RECT 51.885 20.060 55.085 20.240 ;
        RECT 51.250 19.965 51.480 20.020 ;
        RECT 47.240 19.575 51.200 19.805 ;
        RECT 51.885 19.620 54.690 20.060 ;
        RECT 54.855 19.975 55.085 20.060 ;
        RECT 55.295 21.910 55.525 21.975 ;
        RECT 55.690 21.910 56.060 22.795 ;
        RECT 55.295 21.585 56.060 21.910 ;
        RECT 55.295 20.045 56.055 21.585 ;
        RECT 55.295 19.975 55.525 20.045 ;
        RECT 55.045 19.795 55.335 19.815 ;
        RECT 51.885 19.255 54.350 19.620 ;
        RECT 55.020 19.545 55.355 19.795 ;
        RECT 57.590 19.280 58.085 24.395 ;
        RECT 59.105 24.345 59.310 24.480 ;
        RECT 60.590 24.395 60.820 24.645 ;
        RECT 61.610 24.550 62.360 24.990 ;
        RECT 62.780 24.775 63.795 25.775 ;
        RECT 58.385 24.115 60.385 24.345 ;
        RECT 61.610 22.355 61.980 24.550 ;
        RECT 62.130 24.490 62.360 24.550 ;
        RECT 62.850 24.285 63.740 24.775 ;
        RECT 64.420 24.580 65.790 32.380 ;
        RECT 66.325 27.635 67.215 32.695 ;
        RECT 67.850 32.410 68.080 32.490 ;
        RECT 66.320 26.015 67.220 27.635 ;
        RECT 66.325 25.605 67.215 26.015 ;
        RECT 66.250 24.605 67.280 25.605 ;
        RECT 67.850 24.625 68.225 32.410 ;
        RECT 68.500 32.025 70.180 33.260 ;
        RECT 71.015 32.025 75.940 32.035 ;
        RECT 68.500 31.545 75.940 32.025 ;
        RECT 68.500 29.285 70.180 31.545 ;
        RECT 71.015 31.125 75.940 31.545 ;
        RECT 70.520 30.935 70.775 30.960 ;
        RECT 70.520 30.920 70.795 30.935 ;
        RECT 70.490 30.645 70.825 30.920 ;
        RECT 71.000 30.895 76.000 31.125 ;
        RECT 76.210 30.935 76.465 30.960 ;
        RECT 70.520 30.630 70.775 30.645 ;
        RECT 71.000 30.455 76.000 30.685 ;
        RECT 76.205 30.645 76.465 30.935 ;
        RECT 76.210 30.630 76.465 30.645 ;
        RECT 71.045 30.445 75.900 30.455 ;
        RECT 71.045 28.920 73.690 28.925 ;
        RECT 69.720 28.720 73.690 28.920 ;
        RECT 69.720 28.690 73.680 28.720 ;
        RECT 68.560 28.335 68.895 28.610 ;
        RECT 69.440 28.440 69.670 28.485 ;
        RECT 64.420 24.560 64.775 24.580 ;
        RECT 64.420 24.490 64.650 24.560 ;
        RECT 65.560 24.490 65.790 24.580 ;
        RECT 66.320 24.465 67.230 24.605 ;
        RECT 67.850 24.490 68.240 24.625 ;
        RECT 66.310 24.285 67.320 24.465 ;
        RECT 62.410 24.055 64.370 24.285 ;
        RECT 65.840 24.055 67.800 24.285 ;
        RECT 63.165 23.050 63.510 24.055 ;
        RECT 65.865 24.050 67.750 24.055 ;
        RECT 68.045 22.355 68.240 24.490 ;
        RECT 68.630 22.830 68.820 28.335 ;
        RECT 69.250 27.105 69.670 28.440 ;
        RECT 70.975 27.105 72.320 28.690 ;
        RECT 69.250 25.720 72.320 27.105 ;
        RECT 69.250 24.990 69.670 25.720 ;
        RECT 69.245 24.485 69.670 24.990 ;
        RECT 68.630 22.640 68.945 22.830 ;
        RECT 58.950 22.125 62.910 22.355 ;
        RECT 64.380 22.125 68.340 22.355 ;
        RECT 68.755 22.130 68.945 22.640 ;
        RECT 58.670 21.515 58.900 21.965 ;
        RECT 60.150 21.515 60.940 22.125 ;
        RECT 58.670 21.210 60.940 21.515 ;
        RECT 58.615 21.195 60.940 21.210 ;
        RECT 58.530 20.350 60.940 21.195 ;
        RECT 58.530 19.975 58.900 20.350 ;
        RECT 58.670 19.965 58.900 19.975 ;
        RECT 60.150 19.805 60.940 20.350 ;
        RECT 62.960 21.880 63.190 21.965 ;
        RECT 64.100 21.880 64.330 21.965 ;
        RECT 62.960 20.055 64.330 21.880 ;
        RECT 62.960 19.965 63.190 20.055 ;
        RECT 58.950 19.575 62.910 19.805 ;
        RECT 55.490 19.255 58.085 19.280 ;
        RECT 58.530 19.255 58.755 19.265 ;
        RECT 63.430 19.255 63.920 20.055 ;
        RECT 64.100 19.965 64.330 20.055 ;
        RECT 65.815 21.745 67.155 22.125 ;
        RECT 68.390 21.745 68.620 21.965 ;
        RECT 65.815 20.150 68.620 21.745 ;
        RECT 65.815 19.805 67.155 20.150 ;
        RECT 68.390 19.965 68.620 20.150 ;
        RECT 64.380 19.575 68.340 19.805 ;
        RECT 68.770 19.785 68.945 22.130 ;
        RECT 69.245 21.965 69.540 24.485 ;
        RECT 70.975 24.280 72.320 25.720 ;
        RECT 73.730 28.390 73.960 28.485 ;
        RECT 74.205 28.390 74.695 30.445 ;
        RECT 75.265 28.920 75.900 28.925 ;
        RECT 75.150 28.690 79.110 28.920 ;
        RECT 74.870 28.390 75.100 28.485 ;
        RECT 73.730 24.565 75.100 28.390 ;
        RECT 73.730 24.485 73.960 24.565 ;
        RECT 74.870 24.485 75.100 24.565 ;
        RECT 76.525 24.280 77.870 28.690 ;
        RECT 79.160 28.420 79.390 28.485 ;
        RECT 80.045 28.425 80.520 33.260 ;
        RECT 81.845 32.455 82.525 33.260 ;
        RECT 82.945 32.735 83.280 32.985 ;
        RECT 82.960 32.710 83.250 32.735 ;
        RECT 86.420 32.635 88.330 33.260 ;
        RECT 90.420 32.925 92.305 32.930 ;
        RECT 93.865 32.925 95.750 32.930 ;
        RECT 90.410 32.695 92.370 32.925 ;
        RECT 93.840 32.695 95.800 32.925 ;
        RECT 82.770 32.455 83.000 32.505 ;
        RECT 81.845 31.955 83.000 32.455 ;
        RECT 80.915 28.735 81.250 28.985 ;
        RECT 80.935 28.705 81.225 28.735 ;
        RECT 80.745 28.425 80.975 28.500 ;
        RECT 79.160 24.485 79.615 28.420 ;
        RECT 80.045 27.680 80.975 28.425 ;
        RECT 80.380 24.565 80.975 27.680 ;
        RECT 80.745 24.500 80.975 24.565 ;
        RECT 81.185 28.475 81.415 28.500 ;
        RECT 81.185 24.920 81.695 28.475 ;
        RECT 81.185 24.550 81.880 24.920 ;
        RECT 82.380 24.600 83.000 31.955 ;
        RECT 81.185 24.500 81.415 24.550 ;
        RECT 69.720 24.250 73.680 24.280 ;
        RECT 75.150 24.250 79.110 24.280 ;
        RECT 69.720 24.090 79.110 24.250 ;
        RECT 69.720 24.050 73.680 24.090 ;
        RECT 75.150 24.050 79.110 24.090 ;
        RECT 79.275 22.660 79.615 24.485 ;
        RECT 80.925 22.660 81.345 24.305 ;
        RECT 79.275 22.505 81.345 22.660 ;
        RECT 79.350 22.390 81.345 22.505 ;
        RECT 69.810 22.125 73.770 22.355 ;
        RECT 75.240 22.125 79.200 22.355 ;
        RECT 69.245 21.205 69.760 21.965 ;
        RECT 69.315 20.025 69.760 21.205 ;
        RECT 69.530 19.965 69.760 20.025 ;
        RECT 71.190 19.805 72.145 22.125 ;
        RECT 73.820 21.900 74.050 21.965 ;
        RECT 74.960 21.900 75.190 21.965 ;
        RECT 73.820 20.030 75.190 21.900 ;
        RECT 73.820 19.965 74.050 20.030 ;
        RECT 68.755 19.255 68.945 19.785 ;
        RECT 69.810 19.575 73.770 19.805 ;
        RECT 74.225 19.255 74.780 20.030 ;
        RECT 74.960 19.965 75.190 20.030 ;
        RECT 76.635 19.805 77.590 22.125 ;
        RECT 79.350 21.970 79.615 22.390 ;
        RECT 80.925 22.115 81.345 22.390 ;
        RECT 81.580 23.355 81.880 24.550 ;
        RECT 82.770 24.505 83.000 24.600 ;
        RECT 83.210 32.430 83.440 32.505 ;
        RECT 83.210 25.110 83.985 32.430 ;
        RECT 86.385 32.405 88.385 32.635 ;
        RECT 90.130 32.410 90.360 32.490 ;
        RECT 85.950 29.060 86.180 32.355 ;
        RECT 88.590 32.275 88.820 32.355 ;
        RECT 88.560 29.060 88.820 32.275 ;
        RECT 85.950 27.245 88.820 29.060 ;
        RECT 83.210 24.580 84.060 25.110 ;
        RECT 85.950 24.825 86.180 27.245 ;
        RECT 83.210 24.505 83.440 24.580 ;
        RECT 82.875 23.825 83.390 24.315 ;
        RECT 82.875 23.360 83.385 23.825 ;
        RECT 83.690 23.795 84.060 24.580 ;
        RECT 85.590 24.395 86.180 24.825 ;
        RECT 87.075 24.640 87.335 24.960 ;
        RECT 88.560 24.645 88.820 27.245 ;
        RECT 89.890 24.990 90.360 32.410 ;
        RECT 90.850 25.775 91.740 32.695 ;
        RECT 92.420 32.390 92.650 32.490 ;
        RECT 92.420 32.380 92.775 32.390 ;
        RECT 93.560 32.380 93.790 32.490 ;
        RECT 87.130 24.480 87.280 24.640 ;
        RECT 82.510 23.355 83.385 23.360 ;
        RECT 81.580 22.950 83.385 23.355 ;
        RECT 81.580 22.110 81.880 22.950 ;
        RECT 82.510 22.935 83.385 22.950 ;
        RECT 82.875 22.825 83.385 22.935 ;
        RECT 82.875 22.125 83.390 22.825 ;
        RECT 83.615 22.795 84.645 23.795 ;
        RECT 79.275 21.965 79.615 21.970 ;
        RECT 79.250 20.020 79.615 21.965 ;
        RECT 80.830 21.900 81.060 21.970 ;
        RECT 80.335 21.230 81.060 21.900 ;
        RECT 80.325 21.040 81.060 21.230 ;
        RECT 80.325 20.240 80.680 21.040 ;
        RECT 80.830 20.970 81.060 21.040 ;
        RECT 81.270 21.925 81.500 21.970 ;
        RECT 81.640 21.925 81.880 22.110 ;
        RECT 81.270 21.595 81.880 21.925 ;
        RECT 82.855 21.870 83.085 21.975 ;
        RECT 81.270 21.040 81.765 21.595 ;
        RECT 81.270 20.970 81.500 21.040 ;
        RECT 81.020 20.785 81.310 20.810 ;
        RECT 81.005 20.535 81.340 20.785 ;
        RECT 82.625 20.765 83.085 21.870 ;
        RECT 82.305 20.240 83.085 20.765 ;
        RECT 79.885 20.060 83.085 20.240 ;
        RECT 79.250 19.965 79.480 20.020 ;
        RECT 75.240 19.575 79.200 19.805 ;
        RECT 79.885 19.620 82.690 20.060 ;
        RECT 82.855 19.975 83.085 20.060 ;
        RECT 83.295 21.910 83.525 21.975 ;
        RECT 83.690 21.910 84.060 22.795 ;
        RECT 83.295 21.585 84.060 21.910 ;
        RECT 83.295 20.045 84.055 21.585 ;
        RECT 83.295 19.975 83.525 20.045 ;
        RECT 83.045 19.795 83.335 19.815 ;
        RECT 79.885 19.255 82.350 19.620 ;
        RECT 83.020 19.545 83.355 19.795 ;
        RECT 85.590 19.280 86.085 24.395 ;
        RECT 87.105 24.345 87.310 24.480 ;
        RECT 88.590 24.395 88.820 24.645 ;
        RECT 89.610 24.550 90.360 24.990 ;
        RECT 90.780 24.775 91.795 25.775 ;
        RECT 86.385 24.115 88.385 24.345 ;
        RECT 89.610 22.355 89.980 24.550 ;
        RECT 90.130 24.490 90.360 24.550 ;
        RECT 90.850 24.285 91.740 24.775 ;
        RECT 92.420 24.580 93.790 32.380 ;
        RECT 94.325 27.635 95.215 32.695 ;
        RECT 95.850 32.410 96.080 32.490 ;
        RECT 94.320 26.015 95.220 27.635 ;
        RECT 94.325 25.605 95.215 26.015 ;
        RECT 94.250 24.605 95.280 25.605 ;
        RECT 95.850 24.625 96.225 32.410 ;
        RECT 96.500 32.025 98.180 33.260 ;
        RECT 99.015 32.025 103.940 32.035 ;
        RECT 96.500 31.545 103.940 32.025 ;
        RECT 96.500 29.285 98.180 31.545 ;
        RECT 99.015 31.125 103.940 31.545 ;
        RECT 98.520 30.935 98.775 30.960 ;
        RECT 98.520 30.920 98.795 30.935 ;
        RECT 98.490 30.645 98.825 30.920 ;
        RECT 99.000 30.895 104.000 31.125 ;
        RECT 104.210 30.935 104.465 30.960 ;
        RECT 98.520 30.630 98.775 30.645 ;
        RECT 99.000 30.455 104.000 30.685 ;
        RECT 104.205 30.645 104.465 30.935 ;
        RECT 104.210 30.630 104.465 30.645 ;
        RECT 99.045 30.445 103.900 30.455 ;
        RECT 99.045 28.920 101.690 28.925 ;
        RECT 97.720 28.720 101.690 28.920 ;
        RECT 97.720 28.690 101.680 28.720 ;
        RECT 96.560 28.335 96.895 28.610 ;
        RECT 97.440 28.440 97.670 28.485 ;
        RECT 92.420 24.560 92.775 24.580 ;
        RECT 92.420 24.490 92.650 24.560 ;
        RECT 93.560 24.490 93.790 24.580 ;
        RECT 94.320 24.465 95.230 24.605 ;
        RECT 95.850 24.490 96.240 24.625 ;
        RECT 94.310 24.285 95.320 24.465 ;
        RECT 90.410 24.055 92.370 24.285 ;
        RECT 93.840 24.055 95.800 24.285 ;
        RECT 91.125 22.980 91.525 24.055 ;
        RECT 93.865 24.050 95.750 24.055 ;
        RECT 96.045 22.355 96.240 24.490 ;
        RECT 96.630 22.830 96.820 28.335 ;
        RECT 97.250 27.105 97.670 28.440 ;
        RECT 98.975 27.105 100.320 28.690 ;
        RECT 97.250 25.720 100.320 27.105 ;
        RECT 97.250 24.990 97.670 25.720 ;
        RECT 97.245 24.485 97.670 24.990 ;
        RECT 96.630 22.640 96.945 22.830 ;
        RECT 86.950 22.125 90.910 22.355 ;
        RECT 92.380 22.125 96.340 22.355 ;
        RECT 96.755 22.130 96.945 22.640 ;
        RECT 86.670 21.515 86.900 21.965 ;
        RECT 88.150 21.515 88.940 22.125 ;
        RECT 86.670 21.210 88.940 21.515 ;
        RECT 86.615 21.195 88.940 21.210 ;
        RECT 86.530 20.350 88.940 21.195 ;
        RECT 86.530 19.975 86.900 20.350 ;
        RECT 86.670 19.965 86.900 19.975 ;
        RECT 88.150 19.805 88.940 20.350 ;
        RECT 90.960 21.880 91.190 21.965 ;
        RECT 92.100 21.880 92.330 21.965 ;
        RECT 90.960 20.055 92.330 21.880 ;
        RECT 90.960 19.965 91.190 20.055 ;
        RECT 86.950 19.575 90.910 19.805 ;
        RECT 83.790 19.255 86.085 19.280 ;
        RECT 86.530 19.255 86.755 19.265 ;
        RECT 91.430 19.255 91.920 20.055 ;
        RECT 92.100 19.965 92.330 20.055 ;
        RECT 93.815 21.745 95.155 22.125 ;
        RECT 96.390 21.745 96.620 21.965 ;
        RECT 93.815 20.150 96.620 21.745 ;
        RECT 93.815 19.805 95.155 20.150 ;
        RECT 96.390 19.965 96.620 20.150 ;
        RECT 92.380 19.575 96.340 19.805 ;
        RECT 96.770 19.785 96.945 22.130 ;
        RECT 97.245 21.965 97.540 24.485 ;
        RECT 98.975 24.280 100.320 25.720 ;
        RECT 101.730 28.390 101.960 28.485 ;
        RECT 102.205 28.390 102.695 30.445 ;
        RECT 103.265 28.920 103.900 28.925 ;
        RECT 103.150 28.690 107.110 28.920 ;
        RECT 102.870 28.390 103.100 28.485 ;
        RECT 101.730 24.565 103.100 28.390 ;
        RECT 101.730 24.485 101.960 24.565 ;
        RECT 102.870 24.485 103.100 24.565 ;
        RECT 104.525 24.280 105.870 28.690 ;
        RECT 107.160 28.420 107.390 28.485 ;
        RECT 108.045 28.425 108.520 33.260 ;
        RECT 109.845 32.455 110.525 33.260 ;
        RECT 110.945 32.735 111.280 32.985 ;
        RECT 110.960 32.710 111.250 32.735 ;
        RECT 114.420 32.635 116.330 33.260 ;
        RECT 118.420 32.925 120.305 32.930 ;
        RECT 121.865 32.925 123.750 32.930 ;
        RECT 118.410 32.695 120.370 32.925 ;
        RECT 121.840 32.695 123.800 32.925 ;
        RECT 110.770 32.455 111.000 32.505 ;
        RECT 109.845 31.955 111.000 32.455 ;
        RECT 108.915 28.735 109.250 28.985 ;
        RECT 108.935 28.705 109.225 28.735 ;
        RECT 108.745 28.425 108.975 28.500 ;
        RECT 107.160 24.485 107.615 28.420 ;
        RECT 108.045 27.680 108.975 28.425 ;
        RECT 108.380 24.565 108.975 27.680 ;
        RECT 108.745 24.500 108.975 24.565 ;
        RECT 109.185 28.475 109.415 28.500 ;
        RECT 109.185 24.920 109.695 28.475 ;
        RECT 109.185 24.550 109.880 24.920 ;
        RECT 110.380 24.600 111.000 31.955 ;
        RECT 109.185 24.500 109.415 24.550 ;
        RECT 97.720 24.250 101.680 24.280 ;
        RECT 103.150 24.250 107.110 24.280 ;
        RECT 97.720 24.090 107.110 24.250 ;
        RECT 97.720 24.050 101.680 24.090 ;
        RECT 103.150 24.050 107.110 24.090 ;
        RECT 107.275 22.660 107.615 24.485 ;
        RECT 108.925 22.660 109.345 24.305 ;
        RECT 107.275 22.505 109.345 22.660 ;
        RECT 107.350 22.390 109.345 22.505 ;
        RECT 97.810 22.125 101.770 22.355 ;
        RECT 103.240 22.125 107.200 22.355 ;
        RECT 97.245 21.205 97.760 21.965 ;
        RECT 97.315 20.025 97.760 21.205 ;
        RECT 97.530 19.965 97.760 20.025 ;
        RECT 99.190 19.805 100.145 22.125 ;
        RECT 101.820 21.900 102.050 21.965 ;
        RECT 102.960 21.900 103.190 21.965 ;
        RECT 101.820 20.030 103.190 21.900 ;
        RECT 101.820 19.965 102.050 20.030 ;
        RECT 96.755 19.255 96.945 19.785 ;
        RECT 97.810 19.575 101.770 19.805 ;
        RECT 102.225 19.255 102.780 20.030 ;
        RECT 102.960 19.965 103.190 20.030 ;
        RECT 104.635 19.805 105.590 22.125 ;
        RECT 107.350 21.970 107.615 22.390 ;
        RECT 108.925 22.115 109.345 22.390 ;
        RECT 109.580 23.355 109.880 24.550 ;
        RECT 110.770 24.505 111.000 24.600 ;
        RECT 111.210 32.430 111.440 32.505 ;
        RECT 111.210 25.110 111.985 32.430 ;
        RECT 114.385 32.405 116.385 32.635 ;
        RECT 118.130 32.410 118.360 32.490 ;
        RECT 113.950 29.060 114.180 32.355 ;
        RECT 116.590 32.275 116.820 32.355 ;
        RECT 116.560 29.060 116.820 32.275 ;
        RECT 113.950 27.245 116.820 29.060 ;
        RECT 111.210 24.580 112.060 25.110 ;
        RECT 113.950 24.825 114.180 27.245 ;
        RECT 111.210 24.505 111.440 24.580 ;
        RECT 110.875 23.825 111.390 24.315 ;
        RECT 110.875 23.360 111.385 23.825 ;
        RECT 111.690 23.795 112.060 24.580 ;
        RECT 113.590 24.395 114.180 24.825 ;
        RECT 115.075 24.640 115.335 24.960 ;
        RECT 116.560 24.645 116.820 27.245 ;
        RECT 117.890 24.990 118.360 32.410 ;
        RECT 118.850 25.775 119.740 32.695 ;
        RECT 120.420 32.390 120.650 32.490 ;
        RECT 120.420 32.380 120.775 32.390 ;
        RECT 121.560 32.380 121.790 32.490 ;
        RECT 115.130 24.480 115.280 24.640 ;
        RECT 110.510 23.355 111.385 23.360 ;
        RECT 109.580 22.950 111.385 23.355 ;
        RECT 109.580 22.110 109.880 22.950 ;
        RECT 110.510 22.935 111.385 22.950 ;
        RECT 110.875 22.825 111.385 22.935 ;
        RECT 110.875 22.125 111.390 22.825 ;
        RECT 111.585 22.795 112.615 23.795 ;
        RECT 107.275 21.965 107.615 21.970 ;
        RECT 107.250 20.020 107.615 21.965 ;
        RECT 108.830 21.900 109.060 21.970 ;
        RECT 108.335 21.230 109.060 21.900 ;
        RECT 108.325 21.040 109.060 21.230 ;
        RECT 108.325 20.240 108.680 21.040 ;
        RECT 108.830 20.970 109.060 21.040 ;
        RECT 109.270 21.925 109.500 21.970 ;
        RECT 109.640 21.925 109.880 22.110 ;
        RECT 109.270 21.595 109.880 21.925 ;
        RECT 110.855 21.870 111.085 21.975 ;
        RECT 109.270 21.040 109.765 21.595 ;
        RECT 109.270 20.970 109.500 21.040 ;
        RECT 109.020 20.785 109.310 20.810 ;
        RECT 109.005 20.535 109.340 20.785 ;
        RECT 110.625 20.765 111.085 21.870 ;
        RECT 110.305 20.240 111.085 20.765 ;
        RECT 107.885 20.060 111.085 20.240 ;
        RECT 107.250 19.965 107.480 20.020 ;
        RECT 103.240 19.575 107.200 19.805 ;
        RECT 107.885 19.620 110.690 20.060 ;
        RECT 110.855 19.975 111.085 20.060 ;
        RECT 111.295 21.910 111.525 21.975 ;
        RECT 111.690 21.910 112.060 22.795 ;
        RECT 111.295 21.585 112.060 21.910 ;
        RECT 111.295 20.045 112.055 21.585 ;
        RECT 111.295 19.975 111.525 20.045 ;
        RECT 111.045 19.795 111.335 19.815 ;
        RECT 107.885 19.255 110.350 19.620 ;
        RECT 111.020 19.545 111.355 19.795 ;
        RECT 113.590 19.255 114.085 24.395 ;
        RECT 115.105 24.345 115.310 24.480 ;
        RECT 116.590 24.395 116.820 24.645 ;
        RECT 117.610 24.550 118.360 24.990 ;
        RECT 118.780 24.775 119.795 25.775 ;
        RECT 114.385 24.115 116.385 24.345 ;
        RECT 117.610 22.355 117.980 24.550 ;
        RECT 118.130 24.490 118.360 24.550 ;
        RECT 118.850 24.285 119.740 24.775 ;
        RECT 120.420 24.580 121.790 32.380 ;
        RECT 122.325 27.635 123.215 32.695 ;
        RECT 123.850 32.410 124.080 32.490 ;
        RECT 122.320 26.015 123.220 27.635 ;
        RECT 122.325 25.605 123.215 26.015 ;
        RECT 122.250 24.605 123.280 25.605 ;
        RECT 123.850 24.625 124.225 32.410 ;
        RECT 124.500 32.025 126.180 33.260 ;
        RECT 127.015 32.025 131.940 32.035 ;
        RECT 124.500 31.545 131.940 32.025 ;
        RECT 124.500 29.285 126.180 31.545 ;
        RECT 127.015 31.125 131.940 31.545 ;
        RECT 126.520 30.935 126.775 30.960 ;
        RECT 126.520 30.920 126.795 30.935 ;
        RECT 126.490 30.645 126.825 30.920 ;
        RECT 127.000 30.895 132.000 31.125 ;
        RECT 132.210 30.935 132.465 30.960 ;
        RECT 126.520 30.630 126.775 30.645 ;
        RECT 127.000 30.455 132.000 30.685 ;
        RECT 132.205 30.645 132.465 30.935 ;
        RECT 132.210 30.630 132.465 30.645 ;
        RECT 127.045 30.445 131.900 30.455 ;
        RECT 127.045 28.920 129.690 28.925 ;
        RECT 125.720 28.720 129.690 28.920 ;
        RECT 125.720 28.690 129.680 28.720 ;
        RECT 124.560 28.335 124.895 28.610 ;
        RECT 125.440 28.440 125.670 28.485 ;
        RECT 120.420 24.560 120.775 24.580 ;
        RECT 120.420 24.490 120.650 24.560 ;
        RECT 121.560 24.490 121.790 24.580 ;
        RECT 122.320 24.465 123.230 24.605 ;
        RECT 123.850 24.490 124.240 24.625 ;
        RECT 122.310 24.285 123.320 24.465 ;
        RECT 118.410 24.055 120.370 24.285 ;
        RECT 121.840 24.055 123.800 24.285 ;
        RECT 119.160 23.115 119.445 24.055 ;
        RECT 121.865 24.050 123.750 24.055 ;
        RECT 124.045 22.355 124.240 24.490 ;
        RECT 124.630 22.830 124.820 28.335 ;
        RECT 125.250 27.105 125.670 28.440 ;
        RECT 126.975 27.105 128.320 28.690 ;
        RECT 125.250 25.720 128.320 27.105 ;
        RECT 125.250 24.990 125.670 25.720 ;
        RECT 125.245 24.485 125.670 24.990 ;
        RECT 124.630 22.640 124.945 22.830 ;
        RECT 114.950 22.125 118.910 22.355 ;
        RECT 120.380 22.125 124.340 22.355 ;
        RECT 124.755 22.130 124.945 22.640 ;
        RECT 114.670 21.515 114.900 21.965 ;
        RECT 116.150 21.515 116.940 22.125 ;
        RECT 114.670 21.210 116.940 21.515 ;
        RECT 114.615 21.195 116.940 21.210 ;
        RECT 114.530 20.350 116.940 21.195 ;
        RECT 114.530 19.975 114.900 20.350 ;
        RECT 114.670 19.965 114.900 19.975 ;
        RECT 116.150 19.805 116.940 20.350 ;
        RECT 118.960 21.880 119.190 21.965 ;
        RECT 120.100 21.880 120.330 21.965 ;
        RECT 118.960 20.055 120.330 21.880 ;
        RECT 118.960 19.965 119.190 20.055 ;
        RECT 114.950 19.575 118.910 19.805 ;
        RECT 114.530 19.255 114.755 19.265 ;
        RECT 119.430 19.255 119.920 20.055 ;
        RECT 120.100 19.965 120.330 20.055 ;
        RECT 121.815 21.745 123.155 22.125 ;
        RECT 124.390 21.745 124.620 21.965 ;
        RECT 121.815 20.150 124.620 21.745 ;
        RECT 121.815 19.805 123.155 20.150 ;
        RECT 124.390 19.965 124.620 20.150 ;
        RECT 120.380 19.575 124.340 19.805 ;
        RECT 124.770 19.785 124.945 22.130 ;
        RECT 125.245 21.965 125.540 24.485 ;
        RECT 126.975 24.280 128.320 25.720 ;
        RECT 129.730 28.390 129.960 28.485 ;
        RECT 130.205 28.390 130.695 30.445 ;
        RECT 131.265 28.920 131.900 28.925 ;
        RECT 131.150 28.690 135.110 28.920 ;
        RECT 130.870 28.390 131.100 28.485 ;
        RECT 129.730 24.565 131.100 28.390 ;
        RECT 129.730 24.485 129.960 24.565 ;
        RECT 130.870 24.485 131.100 24.565 ;
        RECT 132.525 24.280 133.870 28.690 ;
        RECT 135.160 28.420 135.390 28.485 ;
        RECT 136.045 28.425 136.520 33.260 ;
        RECT 137.845 32.455 138.525 33.260 ;
        RECT 138.945 32.735 139.280 32.985 ;
        RECT 138.960 32.710 139.250 32.735 ;
        RECT 138.770 32.455 139.000 32.505 ;
        RECT 137.845 31.955 139.000 32.455 ;
        RECT 136.915 28.735 137.250 28.985 ;
        RECT 136.935 28.705 137.225 28.735 ;
        RECT 136.745 28.425 136.975 28.500 ;
        RECT 135.160 24.485 135.615 28.420 ;
        RECT 136.045 27.680 136.975 28.425 ;
        RECT 136.380 24.565 136.975 27.680 ;
        RECT 136.745 24.500 136.975 24.565 ;
        RECT 137.185 28.475 137.415 28.500 ;
        RECT 137.185 24.920 137.695 28.475 ;
        RECT 137.185 24.550 137.880 24.920 ;
        RECT 138.380 24.600 139.000 31.955 ;
        RECT 137.185 24.500 137.415 24.550 ;
        RECT 125.720 24.250 129.680 24.280 ;
        RECT 131.150 24.250 135.110 24.280 ;
        RECT 125.720 24.090 135.110 24.250 ;
        RECT 125.720 24.050 129.680 24.090 ;
        RECT 131.150 24.050 135.110 24.090 ;
        RECT 135.275 22.660 135.615 24.485 ;
        RECT 136.925 22.660 137.345 24.305 ;
        RECT 135.275 22.505 137.345 22.660 ;
        RECT 135.350 22.390 137.345 22.505 ;
        RECT 125.810 22.125 129.770 22.355 ;
        RECT 131.240 22.125 135.200 22.355 ;
        RECT 125.245 21.205 125.760 21.965 ;
        RECT 125.315 20.025 125.760 21.205 ;
        RECT 125.530 19.965 125.760 20.025 ;
        RECT 127.190 19.805 128.145 22.125 ;
        RECT 129.820 21.900 130.050 21.965 ;
        RECT 130.960 21.900 131.190 21.965 ;
        RECT 129.820 20.030 131.190 21.900 ;
        RECT 129.820 19.965 130.050 20.030 ;
        RECT 124.755 19.255 124.945 19.785 ;
        RECT 125.810 19.575 129.770 19.805 ;
        RECT 130.225 19.255 130.780 20.030 ;
        RECT 130.960 19.965 131.190 20.030 ;
        RECT 132.635 19.805 133.590 22.125 ;
        RECT 135.350 21.970 135.615 22.390 ;
        RECT 136.925 22.115 137.345 22.390 ;
        RECT 137.580 23.355 137.880 24.550 ;
        RECT 138.770 24.505 139.000 24.600 ;
        RECT 139.210 32.430 139.440 32.505 ;
        RECT 139.210 25.110 139.985 32.430 ;
        RECT 139.210 24.580 140.060 25.110 ;
        RECT 139.210 24.505 139.440 24.580 ;
        RECT 138.875 23.825 139.390 24.315 ;
        RECT 138.875 23.360 139.385 23.825 ;
        RECT 139.690 23.795 140.060 24.580 ;
        RECT 138.510 23.355 139.385 23.360 ;
        RECT 137.580 22.950 139.385 23.355 ;
        RECT 137.580 22.110 137.880 22.950 ;
        RECT 138.510 22.935 139.385 22.950 ;
        RECT 138.875 22.825 139.385 22.935 ;
        RECT 138.875 22.125 139.390 22.825 ;
        RECT 139.615 22.795 140.645 23.795 ;
        RECT 135.275 21.965 135.615 21.970 ;
        RECT 135.250 20.020 135.615 21.965 ;
        RECT 136.830 21.900 137.060 21.970 ;
        RECT 136.335 21.230 137.060 21.900 ;
        RECT 136.325 21.040 137.060 21.230 ;
        RECT 136.325 20.240 136.680 21.040 ;
        RECT 136.830 20.970 137.060 21.040 ;
        RECT 137.270 21.925 137.500 21.970 ;
        RECT 137.640 21.925 137.880 22.110 ;
        RECT 137.270 21.595 137.880 21.925 ;
        RECT 138.855 21.870 139.085 21.975 ;
        RECT 137.270 21.040 137.765 21.595 ;
        RECT 137.270 20.970 137.500 21.040 ;
        RECT 137.020 20.785 137.310 20.810 ;
        RECT 137.005 20.535 137.340 20.785 ;
        RECT 138.625 20.765 139.085 21.870 ;
        RECT 138.305 20.240 139.085 20.765 ;
        RECT 135.885 20.060 139.085 20.240 ;
        RECT 135.250 19.965 135.480 20.020 ;
        RECT 131.240 19.575 135.200 19.805 ;
        RECT 135.885 19.620 138.690 20.060 ;
        RECT 138.855 19.975 139.085 20.060 ;
        RECT 139.295 21.910 139.525 21.975 ;
        RECT 139.690 21.910 140.060 22.795 ;
        RECT 139.295 21.585 140.060 21.910 ;
        RECT 139.295 20.045 140.055 21.585 ;
        RECT 139.295 19.975 139.525 20.045 ;
        RECT 139.045 19.795 139.335 19.815 ;
        RECT 135.885 19.255 138.350 19.620 ;
        RECT 139.020 19.545 139.355 19.795 ;
        RECT 1.475 18.380 112.080 19.255 ;
        RECT 113.475 18.380 140.080 19.255 ;
        RECT 27.790 17.960 30.690 17.980 ;
        RECT 55.390 17.960 57.890 17.980 ;
        RECT 68.845 17.960 69.785 17.985 ;
        RECT 83.690 17.960 86.190 17.980 ;
        RECT 1.450 17.280 111.925 17.960 ;
        RECT 1.450 17.260 27.925 17.280 ;
        RECT 29.450 17.260 55.925 17.280 ;
        RECT 57.450 17.260 83.925 17.280 ;
        RECT 85.450 17.260 111.925 17.280 ;
        RECT 113.450 17.260 139.925 17.960 ;
        RECT 2.420 16.635 4.330 17.260 ;
        RECT 6.420 16.925 8.305 16.930 ;
        RECT 9.865 16.925 11.750 16.930 ;
        RECT 6.410 16.695 8.370 16.925 ;
        RECT 9.840 16.695 11.800 16.925 ;
        RECT 2.385 16.405 4.385 16.635 ;
        RECT 6.130 16.410 6.360 16.490 ;
        RECT 1.950 13.060 2.180 16.355 ;
        RECT 4.590 16.275 4.820 16.355 ;
        RECT 4.560 13.060 4.820 16.275 ;
        RECT 1.950 11.245 4.820 13.060 ;
        RECT 1.950 8.825 2.180 11.245 ;
        RECT 1.590 8.395 2.180 8.825 ;
        RECT 3.075 8.640 3.335 8.960 ;
        RECT 4.560 8.645 4.820 11.245 ;
        RECT 5.890 8.990 6.360 16.410 ;
        RECT 6.850 9.775 7.740 16.695 ;
        RECT 8.420 16.390 8.650 16.490 ;
        RECT 8.420 16.380 8.775 16.390 ;
        RECT 9.560 16.380 9.790 16.490 ;
        RECT 3.130 8.480 3.280 8.640 ;
        RECT 1.590 3.255 2.085 8.395 ;
        RECT 3.105 8.345 3.310 8.480 ;
        RECT 4.590 8.395 4.820 8.645 ;
        RECT 5.610 8.550 6.360 8.990 ;
        RECT 6.780 8.775 7.795 9.775 ;
        RECT 2.385 8.115 4.385 8.345 ;
        RECT 5.610 6.355 5.980 8.550 ;
        RECT 6.130 8.490 6.360 8.550 ;
        RECT 6.850 8.285 7.740 8.775 ;
        RECT 8.420 8.580 9.790 16.380 ;
        RECT 10.325 11.635 11.215 16.695 ;
        RECT 11.850 16.410 12.080 16.490 ;
        RECT 10.320 10.015 11.220 11.635 ;
        RECT 10.325 9.605 11.215 10.015 ;
        RECT 10.250 8.605 11.280 9.605 ;
        RECT 11.850 8.625 12.225 16.410 ;
        RECT 12.500 16.025 14.180 17.260 ;
        RECT 15.015 16.025 19.940 16.035 ;
        RECT 12.500 15.545 19.940 16.025 ;
        RECT 12.500 13.285 14.180 15.545 ;
        RECT 15.015 15.125 19.940 15.545 ;
        RECT 14.520 14.935 14.775 14.960 ;
        RECT 14.520 14.920 14.795 14.935 ;
        RECT 14.490 14.645 14.825 14.920 ;
        RECT 15.000 14.895 20.000 15.125 ;
        RECT 20.210 14.935 20.465 14.960 ;
        RECT 14.520 14.630 14.775 14.645 ;
        RECT 15.000 14.455 20.000 14.685 ;
        RECT 20.205 14.645 20.465 14.935 ;
        RECT 20.210 14.630 20.465 14.645 ;
        RECT 15.045 14.445 19.900 14.455 ;
        RECT 15.045 12.920 17.690 12.925 ;
        RECT 13.720 12.720 17.690 12.920 ;
        RECT 13.720 12.690 17.680 12.720 ;
        RECT 12.560 12.335 12.895 12.610 ;
        RECT 13.440 12.440 13.670 12.485 ;
        RECT 8.420 8.560 8.775 8.580 ;
        RECT 8.420 8.490 8.650 8.560 ;
        RECT 9.560 8.490 9.790 8.580 ;
        RECT 10.320 8.465 11.230 8.605 ;
        RECT 11.850 8.490 12.240 8.625 ;
        RECT 10.310 8.285 11.320 8.465 ;
        RECT 6.410 8.055 8.370 8.285 ;
        RECT 9.840 8.055 11.800 8.285 ;
        RECT 7.130 7.085 7.460 8.055 ;
        RECT 9.865 8.050 11.750 8.055 ;
        RECT 12.045 6.355 12.240 8.490 ;
        RECT 12.630 6.830 12.820 12.335 ;
        RECT 13.250 11.105 13.670 12.440 ;
        RECT 14.975 11.105 16.320 12.690 ;
        RECT 13.250 9.720 16.320 11.105 ;
        RECT 13.250 8.990 13.670 9.720 ;
        RECT 13.245 8.485 13.670 8.990 ;
        RECT 12.630 6.640 12.945 6.830 ;
        RECT 2.950 6.125 6.910 6.355 ;
        RECT 8.380 6.125 12.340 6.355 ;
        RECT 12.755 6.130 12.945 6.640 ;
        RECT 2.670 5.515 2.900 5.965 ;
        RECT 4.150 5.515 4.940 6.125 ;
        RECT 2.670 5.210 4.940 5.515 ;
        RECT 2.615 5.195 4.940 5.210 ;
        RECT 2.530 4.350 4.940 5.195 ;
        RECT 2.530 3.975 2.900 4.350 ;
        RECT 2.670 3.965 2.900 3.975 ;
        RECT 4.150 3.805 4.940 4.350 ;
        RECT 6.960 5.880 7.190 5.965 ;
        RECT 8.100 5.880 8.330 5.965 ;
        RECT 6.960 4.055 8.330 5.880 ;
        RECT 6.960 3.965 7.190 4.055 ;
        RECT 2.950 3.575 6.910 3.805 ;
        RECT 2.530 3.255 2.755 3.265 ;
        RECT 7.430 3.255 7.920 4.055 ;
        RECT 8.100 3.965 8.330 4.055 ;
        RECT 9.815 5.745 11.155 6.125 ;
        RECT 12.390 5.745 12.620 5.965 ;
        RECT 9.815 4.150 12.620 5.745 ;
        RECT 9.815 3.805 11.155 4.150 ;
        RECT 12.390 3.965 12.620 4.150 ;
        RECT 8.380 3.575 12.340 3.805 ;
        RECT 12.770 3.785 12.945 6.130 ;
        RECT 13.245 5.965 13.540 8.485 ;
        RECT 14.975 8.280 16.320 9.720 ;
        RECT 17.730 12.390 17.960 12.485 ;
        RECT 18.205 12.390 18.695 14.445 ;
        RECT 19.265 12.920 19.900 12.925 ;
        RECT 19.150 12.690 23.110 12.920 ;
        RECT 18.870 12.390 19.100 12.485 ;
        RECT 17.730 8.565 19.100 12.390 ;
        RECT 17.730 8.485 17.960 8.565 ;
        RECT 18.870 8.485 19.100 8.565 ;
        RECT 20.525 8.280 21.870 12.690 ;
        RECT 23.160 12.420 23.390 12.485 ;
        RECT 24.045 12.425 24.520 17.260 ;
        RECT 25.845 16.455 26.525 17.260 ;
        RECT 26.945 16.735 27.280 16.985 ;
        RECT 26.960 16.710 27.250 16.735 ;
        RECT 30.420 16.635 32.330 17.260 ;
        RECT 34.420 16.925 36.305 16.930 ;
        RECT 37.865 16.925 39.750 16.930 ;
        RECT 34.410 16.695 36.370 16.925 ;
        RECT 37.840 16.695 39.800 16.925 ;
        RECT 26.770 16.455 27.000 16.505 ;
        RECT 25.845 15.955 27.000 16.455 ;
        RECT 24.915 12.735 25.250 12.985 ;
        RECT 24.935 12.705 25.225 12.735 ;
        RECT 24.745 12.425 24.975 12.500 ;
        RECT 23.160 8.485 23.615 12.420 ;
        RECT 24.045 11.680 24.975 12.425 ;
        RECT 24.380 8.565 24.975 11.680 ;
        RECT 24.745 8.500 24.975 8.565 ;
        RECT 25.185 12.475 25.415 12.500 ;
        RECT 25.185 8.920 25.695 12.475 ;
        RECT 25.185 8.550 25.880 8.920 ;
        RECT 26.380 8.600 27.000 15.955 ;
        RECT 25.185 8.500 25.415 8.550 ;
        RECT 13.720 8.250 17.680 8.280 ;
        RECT 19.150 8.250 23.110 8.280 ;
        RECT 13.720 8.090 23.110 8.250 ;
        RECT 13.720 8.050 17.680 8.090 ;
        RECT 19.150 8.050 23.110 8.090 ;
        RECT 23.275 6.660 23.615 8.485 ;
        RECT 24.925 6.660 25.345 8.305 ;
        RECT 23.275 6.505 25.345 6.660 ;
        RECT 23.350 6.390 25.345 6.505 ;
        RECT 13.810 6.125 17.770 6.355 ;
        RECT 19.240 6.125 23.200 6.355 ;
        RECT 13.245 5.205 13.760 5.965 ;
        RECT 13.315 4.025 13.760 5.205 ;
        RECT 13.530 3.965 13.760 4.025 ;
        RECT 15.190 3.805 16.145 6.125 ;
        RECT 17.820 5.900 18.050 5.965 ;
        RECT 18.960 5.900 19.190 5.965 ;
        RECT 17.820 4.030 19.190 5.900 ;
        RECT 17.820 3.965 18.050 4.030 ;
        RECT 12.755 3.255 12.945 3.785 ;
        RECT 13.810 3.575 17.770 3.805 ;
        RECT 18.225 3.255 18.780 4.030 ;
        RECT 18.960 3.965 19.190 4.030 ;
        RECT 20.635 3.805 21.590 6.125 ;
        RECT 23.350 5.970 23.615 6.390 ;
        RECT 24.925 6.115 25.345 6.390 ;
        RECT 25.580 7.355 25.880 8.550 ;
        RECT 26.770 8.505 27.000 8.600 ;
        RECT 27.210 16.430 27.440 16.505 ;
        RECT 27.210 9.110 27.985 16.430 ;
        RECT 30.385 16.405 32.385 16.635 ;
        RECT 34.130 16.410 34.360 16.490 ;
        RECT 29.950 13.060 30.180 16.355 ;
        RECT 32.590 16.275 32.820 16.355 ;
        RECT 32.560 13.060 32.820 16.275 ;
        RECT 29.950 11.245 32.820 13.060 ;
        RECT 27.210 8.580 28.060 9.110 ;
        RECT 29.950 8.825 30.180 11.245 ;
        RECT 27.210 8.505 27.440 8.580 ;
        RECT 26.875 7.825 27.390 8.315 ;
        RECT 27.690 7.825 28.060 8.580 ;
        RECT 29.590 8.395 30.180 8.825 ;
        RECT 31.075 8.640 31.335 8.960 ;
        RECT 32.560 8.645 32.820 11.245 ;
        RECT 33.890 8.990 34.360 16.410 ;
        RECT 34.850 9.775 35.740 16.695 ;
        RECT 36.420 16.390 36.650 16.490 ;
        RECT 36.420 16.380 36.775 16.390 ;
        RECT 37.560 16.380 37.790 16.490 ;
        RECT 31.130 8.480 31.280 8.640 ;
        RECT 26.875 7.360 27.385 7.825 ;
        RECT 26.510 7.355 27.385 7.360 ;
        RECT 25.580 6.950 27.385 7.355 ;
        RECT 25.580 6.110 25.880 6.950 ;
        RECT 26.510 6.935 27.385 6.950 ;
        RECT 26.875 6.825 27.385 6.935 ;
        RECT 26.875 6.125 27.390 6.825 ;
        RECT 27.615 6.795 28.615 7.825 ;
        RECT 23.275 5.965 23.615 5.970 ;
        RECT 23.250 4.020 23.615 5.965 ;
        RECT 24.830 5.900 25.060 5.970 ;
        RECT 24.335 5.230 25.060 5.900 ;
        RECT 24.325 5.040 25.060 5.230 ;
        RECT 24.325 4.240 24.680 5.040 ;
        RECT 24.830 4.970 25.060 5.040 ;
        RECT 25.270 5.925 25.500 5.970 ;
        RECT 25.640 5.925 25.880 6.110 ;
        RECT 25.270 5.595 25.880 5.925 ;
        RECT 26.855 5.870 27.085 5.975 ;
        RECT 25.270 5.040 25.765 5.595 ;
        RECT 25.270 4.970 25.500 5.040 ;
        RECT 25.020 4.785 25.310 4.810 ;
        RECT 25.005 4.535 25.340 4.785 ;
        RECT 26.625 4.765 27.085 5.870 ;
        RECT 26.305 4.240 27.085 4.765 ;
        RECT 23.885 4.060 27.085 4.240 ;
        RECT 23.250 3.965 23.480 4.020 ;
        RECT 19.240 3.575 23.200 3.805 ;
        RECT 23.885 3.620 26.690 4.060 ;
        RECT 26.855 3.975 27.085 4.060 ;
        RECT 27.295 5.910 27.525 5.975 ;
        RECT 27.690 5.910 28.060 6.795 ;
        RECT 27.295 5.585 28.060 5.910 ;
        RECT 27.295 4.045 28.055 5.585 ;
        RECT 27.295 3.975 27.525 4.045 ;
        RECT 27.045 3.795 27.335 3.815 ;
        RECT 23.885 3.255 26.350 3.620 ;
        RECT 27.020 3.545 27.355 3.795 ;
        RECT 29.590 3.280 30.085 8.395 ;
        RECT 31.105 8.345 31.310 8.480 ;
        RECT 32.590 8.395 32.820 8.645 ;
        RECT 33.610 8.550 34.360 8.990 ;
        RECT 34.780 8.775 35.795 9.775 ;
        RECT 30.385 8.115 32.385 8.345 ;
        RECT 33.610 6.355 33.980 8.550 ;
        RECT 34.130 8.490 34.360 8.550 ;
        RECT 34.850 8.285 35.740 8.775 ;
        RECT 36.420 8.580 37.790 16.380 ;
        RECT 38.325 11.635 39.215 16.695 ;
        RECT 39.850 16.410 40.080 16.490 ;
        RECT 38.320 10.015 39.220 11.635 ;
        RECT 38.325 9.605 39.215 10.015 ;
        RECT 38.250 8.605 39.280 9.605 ;
        RECT 39.850 8.625 40.225 16.410 ;
        RECT 40.500 16.025 42.180 17.260 ;
        RECT 43.015 16.025 47.940 16.035 ;
        RECT 40.500 15.545 47.940 16.025 ;
        RECT 40.500 13.285 42.180 15.545 ;
        RECT 43.015 15.125 47.940 15.545 ;
        RECT 42.520 14.935 42.775 14.960 ;
        RECT 42.520 14.920 42.795 14.935 ;
        RECT 42.490 14.645 42.825 14.920 ;
        RECT 43.000 14.895 48.000 15.125 ;
        RECT 48.210 14.935 48.465 14.960 ;
        RECT 42.520 14.630 42.775 14.645 ;
        RECT 43.000 14.455 48.000 14.685 ;
        RECT 48.205 14.645 48.465 14.935 ;
        RECT 48.210 14.630 48.465 14.645 ;
        RECT 43.045 14.445 47.900 14.455 ;
        RECT 43.045 12.920 45.690 12.925 ;
        RECT 41.720 12.720 45.690 12.920 ;
        RECT 41.720 12.690 45.680 12.720 ;
        RECT 40.560 12.335 40.895 12.610 ;
        RECT 41.440 12.440 41.670 12.485 ;
        RECT 36.420 8.560 36.775 8.580 ;
        RECT 36.420 8.490 36.650 8.560 ;
        RECT 37.560 8.490 37.790 8.580 ;
        RECT 38.320 8.465 39.230 8.605 ;
        RECT 39.850 8.490 40.240 8.625 ;
        RECT 38.310 8.285 39.320 8.465 ;
        RECT 34.410 8.055 36.370 8.285 ;
        RECT 37.840 8.055 39.800 8.285 ;
        RECT 35.210 7.040 35.560 8.055 ;
        RECT 37.865 8.050 39.750 8.055 ;
        RECT 40.045 6.355 40.240 8.490 ;
        RECT 40.630 6.830 40.820 12.335 ;
        RECT 41.250 11.105 41.670 12.440 ;
        RECT 42.975 11.105 44.320 12.690 ;
        RECT 41.250 9.720 44.320 11.105 ;
        RECT 41.250 8.990 41.670 9.720 ;
        RECT 41.245 8.485 41.670 8.990 ;
        RECT 40.630 6.640 40.945 6.830 ;
        RECT 30.950 6.125 34.910 6.355 ;
        RECT 36.380 6.125 40.340 6.355 ;
        RECT 40.755 6.130 40.945 6.640 ;
        RECT 30.670 5.515 30.900 5.965 ;
        RECT 32.150 5.515 32.940 6.125 ;
        RECT 30.670 5.210 32.940 5.515 ;
        RECT 30.615 5.195 32.940 5.210 ;
        RECT 30.530 4.350 32.940 5.195 ;
        RECT 30.530 3.975 30.900 4.350 ;
        RECT 30.670 3.965 30.900 3.975 ;
        RECT 32.150 3.805 32.940 4.350 ;
        RECT 34.960 5.880 35.190 5.965 ;
        RECT 36.100 5.880 36.330 5.965 ;
        RECT 34.960 4.055 36.330 5.880 ;
        RECT 34.960 3.965 35.190 4.055 ;
        RECT 30.950 3.575 34.910 3.805 ;
        RECT 27.990 3.255 30.090 3.280 ;
        RECT 30.530 3.255 30.755 3.265 ;
        RECT 35.430 3.255 35.920 4.055 ;
        RECT 36.100 3.965 36.330 4.055 ;
        RECT 37.815 5.745 39.155 6.125 ;
        RECT 40.390 5.745 40.620 5.965 ;
        RECT 37.815 4.150 40.620 5.745 ;
        RECT 37.815 3.805 39.155 4.150 ;
        RECT 40.390 3.965 40.620 4.150 ;
        RECT 36.380 3.575 40.340 3.805 ;
        RECT 40.770 3.785 40.945 6.130 ;
        RECT 41.245 5.965 41.540 8.485 ;
        RECT 42.975 8.280 44.320 9.720 ;
        RECT 45.730 12.390 45.960 12.485 ;
        RECT 46.205 12.390 46.695 14.445 ;
        RECT 47.265 12.920 47.900 12.925 ;
        RECT 47.150 12.690 51.110 12.920 ;
        RECT 46.870 12.390 47.100 12.485 ;
        RECT 45.730 8.565 47.100 12.390 ;
        RECT 45.730 8.485 45.960 8.565 ;
        RECT 46.870 8.485 47.100 8.565 ;
        RECT 48.525 8.280 49.870 12.690 ;
        RECT 51.160 12.420 51.390 12.485 ;
        RECT 52.045 12.425 52.520 17.260 ;
        RECT 53.845 16.455 54.525 17.260 ;
        RECT 54.945 16.735 55.280 16.985 ;
        RECT 54.960 16.710 55.250 16.735 ;
        RECT 58.420 16.635 60.330 17.260 ;
        RECT 62.420 16.925 64.305 16.930 ;
        RECT 65.865 16.925 67.750 16.930 ;
        RECT 62.410 16.695 64.370 16.925 ;
        RECT 65.840 16.695 67.800 16.925 ;
        RECT 54.770 16.455 55.000 16.505 ;
        RECT 53.845 15.955 55.000 16.455 ;
        RECT 52.915 12.735 53.250 12.985 ;
        RECT 52.935 12.705 53.225 12.735 ;
        RECT 52.745 12.425 52.975 12.500 ;
        RECT 51.160 8.485 51.615 12.420 ;
        RECT 52.045 11.680 52.975 12.425 ;
        RECT 52.380 8.565 52.975 11.680 ;
        RECT 52.745 8.500 52.975 8.565 ;
        RECT 53.185 12.475 53.415 12.500 ;
        RECT 53.185 8.920 53.695 12.475 ;
        RECT 53.185 8.550 53.880 8.920 ;
        RECT 54.380 8.600 55.000 15.955 ;
        RECT 53.185 8.500 53.415 8.550 ;
        RECT 41.720 8.250 45.680 8.280 ;
        RECT 47.150 8.250 51.110 8.280 ;
        RECT 41.720 8.090 51.110 8.250 ;
        RECT 41.720 8.050 45.680 8.090 ;
        RECT 47.150 8.050 51.110 8.090 ;
        RECT 51.275 6.660 51.615 8.485 ;
        RECT 52.925 6.660 53.345 8.305 ;
        RECT 51.275 6.505 53.345 6.660 ;
        RECT 51.350 6.390 53.345 6.505 ;
        RECT 41.810 6.125 45.770 6.355 ;
        RECT 47.240 6.125 51.200 6.355 ;
        RECT 41.245 5.205 41.760 5.965 ;
        RECT 41.315 4.025 41.760 5.205 ;
        RECT 41.530 3.965 41.760 4.025 ;
        RECT 43.190 3.805 44.145 6.125 ;
        RECT 45.820 5.900 46.050 5.965 ;
        RECT 46.960 5.900 47.190 5.965 ;
        RECT 45.820 4.030 47.190 5.900 ;
        RECT 45.820 3.965 46.050 4.030 ;
        RECT 40.755 3.255 40.945 3.785 ;
        RECT 41.810 3.575 45.770 3.805 ;
        RECT 46.225 3.255 46.780 4.030 ;
        RECT 46.960 3.965 47.190 4.030 ;
        RECT 48.635 3.805 49.590 6.125 ;
        RECT 51.350 5.970 51.615 6.390 ;
        RECT 52.925 6.115 53.345 6.390 ;
        RECT 53.580 7.355 53.880 8.550 ;
        RECT 54.770 8.505 55.000 8.600 ;
        RECT 55.210 16.430 55.440 16.505 ;
        RECT 55.210 9.110 55.985 16.430 ;
        RECT 58.385 16.405 60.385 16.635 ;
        RECT 62.130 16.410 62.360 16.490 ;
        RECT 57.950 13.060 58.180 16.355 ;
        RECT 60.590 16.275 60.820 16.355 ;
        RECT 60.560 13.060 60.820 16.275 ;
        RECT 57.950 11.245 60.820 13.060 ;
        RECT 55.210 8.580 56.060 9.110 ;
        RECT 57.950 8.825 58.180 11.245 ;
        RECT 55.210 8.505 55.440 8.580 ;
        RECT 54.875 7.825 55.390 8.315 ;
        RECT 54.875 7.360 55.385 7.825 ;
        RECT 55.690 7.795 56.060 8.580 ;
        RECT 57.590 8.395 58.180 8.825 ;
        RECT 59.075 8.640 59.335 8.960 ;
        RECT 60.560 8.645 60.820 11.245 ;
        RECT 61.890 8.990 62.360 16.410 ;
        RECT 62.850 9.775 63.740 16.695 ;
        RECT 64.420 16.390 64.650 16.490 ;
        RECT 64.420 16.380 64.775 16.390 ;
        RECT 65.560 16.380 65.790 16.490 ;
        RECT 59.130 8.480 59.280 8.640 ;
        RECT 54.510 7.355 55.385 7.360 ;
        RECT 53.580 6.950 55.385 7.355 ;
        RECT 53.580 6.110 53.880 6.950 ;
        RECT 54.510 6.935 55.385 6.950 ;
        RECT 54.875 6.825 55.385 6.935 ;
        RECT 54.875 6.125 55.390 6.825 ;
        RECT 55.615 6.795 56.645 7.795 ;
        RECT 51.275 5.965 51.615 5.970 ;
        RECT 51.250 4.020 51.615 5.965 ;
        RECT 52.830 5.900 53.060 5.970 ;
        RECT 52.335 5.230 53.060 5.900 ;
        RECT 52.325 5.040 53.060 5.230 ;
        RECT 52.325 4.240 52.680 5.040 ;
        RECT 52.830 4.970 53.060 5.040 ;
        RECT 53.270 5.925 53.500 5.970 ;
        RECT 53.640 5.925 53.880 6.110 ;
        RECT 53.270 5.595 53.880 5.925 ;
        RECT 54.855 5.870 55.085 5.975 ;
        RECT 53.270 5.040 53.765 5.595 ;
        RECT 53.270 4.970 53.500 5.040 ;
        RECT 53.020 4.785 53.310 4.810 ;
        RECT 53.005 4.535 53.340 4.785 ;
        RECT 54.625 4.765 55.085 5.870 ;
        RECT 54.305 4.240 55.085 4.765 ;
        RECT 51.885 4.060 55.085 4.240 ;
        RECT 51.250 3.965 51.480 4.020 ;
        RECT 47.240 3.575 51.200 3.805 ;
        RECT 51.885 3.620 54.690 4.060 ;
        RECT 54.855 3.975 55.085 4.060 ;
        RECT 55.295 5.910 55.525 5.975 ;
        RECT 55.690 5.910 56.060 6.795 ;
        RECT 55.295 5.585 56.060 5.910 ;
        RECT 55.295 4.045 56.055 5.585 ;
        RECT 55.295 3.975 55.525 4.045 ;
        RECT 55.045 3.795 55.335 3.815 ;
        RECT 51.885 3.255 54.350 3.620 ;
        RECT 55.020 3.545 55.355 3.795 ;
        RECT 57.590 3.280 58.085 8.395 ;
        RECT 59.105 8.345 59.310 8.480 ;
        RECT 60.590 8.395 60.820 8.645 ;
        RECT 61.610 8.550 62.360 8.990 ;
        RECT 62.780 8.775 63.795 9.775 ;
        RECT 58.385 8.115 60.385 8.345 ;
        RECT 61.610 6.355 61.980 8.550 ;
        RECT 62.130 8.490 62.360 8.550 ;
        RECT 62.850 8.285 63.740 8.775 ;
        RECT 64.420 8.580 65.790 16.380 ;
        RECT 66.325 11.635 67.215 16.695 ;
        RECT 67.850 16.410 68.080 16.490 ;
        RECT 66.320 10.015 67.220 11.635 ;
        RECT 66.325 9.605 67.215 10.015 ;
        RECT 66.250 8.605 67.280 9.605 ;
        RECT 67.850 8.625 68.225 16.410 ;
        RECT 68.500 16.025 70.180 17.260 ;
        RECT 71.015 16.025 75.940 16.035 ;
        RECT 68.500 15.545 75.940 16.025 ;
        RECT 68.500 13.285 70.180 15.545 ;
        RECT 71.015 15.125 75.940 15.545 ;
        RECT 70.520 14.935 70.775 14.960 ;
        RECT 70.520 14.920 70.795 14.935 ;
        RECT 70.490 14.645 70.825 14.920 ;
        RECT 71.000 14.895 76.000 15.125 ;
        RECT 76.210 14.935 76.465 14.960 ;
        RECT 70.520 14.630 70.775 14.645 ;
        RECT 71.000 14.455 76.000 14.685 ;
        RECT 76.205 14.645 76.465 14.935 ;
        RECT 76.210 14.630 76.465 14.645 ;
        RECT 71.045 14.445 75.900 14.455 ;
        RECT 71.045 12.920 73.690 12.925 ;
        RECT 69.720 12.720 73.690 12.920 ;
        RECT 69.720 12.690 73.680 12.720 ;
        RECT 68.560 12.335 68.895 12.610 ;
        RECT 69.440 12.440 69.670 12.485 ;
        RECT 64.420 8.560 64.775 8.580 ;
        RECT 64.420 8.490 64.650 8.560 ;
        RECT 65.560 8.490 65.790 8.580 ;
        RECT 66.320 8.465 67.230 8.605 ;
        RECT 67.850 8.490 68.240 8.625 ;
        RECT 66.310 8.285 67.320 8.465 ;
        RECT 62.410 8.055 64.370 8.285 ;
        RECT 65.840 8.055 67.800 8.285 ;
        RECT 63.125 7.090 63.470 8.055 ;
        RECT 65.865 8.050 67.750 8.055 ;
        RECT 68.045 6.355 68.240 8.490 ;
        RECT 68.630 6.830 68.820 12.335 ;
        RECT 69.250 11.105 69.670 12.440 ;
        RECT 70.975 11.105 72.320 12.690 ;
        RECT 69.250 9.720 72.320 11.105 ;
        RECT 69.250 8.990 69.670 9.720 ;
        RECT 69.245 8.485 69.670 8.990 ;
        RECT 68.630 6.640 68.945 6.830 ;
        RECT 58.950 6.125 62.910 6.355 ;
        RECT 64.380 6.125 68.340 6.355 ;
        RECT 68.755 6.130 68.945 6.640 ;
        RECT 58.670 5.515 58.900 5.965 ;
        RECT 60.150 5.515 60.940 6.125 ;
        RECT 58.670 5.210 60.940 5.515 ;
        RECT 58.615 5.195 60.940 5.210 ;
        RECT 58.530 4.350 60.940 5.195 ;
        RECT 58.530 3.975 58.900 4.350 ;
        RECT 58.670 3.965 58.900 3.975 ;
        RECT 60.150 3.805 60.940 4.350 ;
        RECT 62.960 5.880 63.190 5.965 ;
        RECT 64.100 5.880 64.330 5.965 ;
        RECT 62.960 4.055 64.330 5.880 ;
        RECT 62.960 3.965 63.190 4.055 ;
        RECT 58.950 3.575 62.910 3.805 ;
        RECT 55.790 3.255 58.085 3.280 ;
        RECT 58.530 3.255 58.755 3.265 ;
        RECT 63.430 3.255 63.920 4.055 ;
        RECT 64.100 3.965 64.330 4.055 ;
        RECT 65.815 5.745 67.155 6.125 ;
        RECT 68.390 5.745 68.620 5.965 ;
        RECT 65.815 4.150 68.620 5.745 ;
        RECT 65.815 3.805 67.155 4.150 ;
        RECT 68.390 3.965 68.620 4.150 ;
        RECT 64.380 3.575 68.340 3.805 ;
        RECT 68.770 3.785 68.945 6.130 ;
        RECT 69.245 5.965 69.540 8.485 ;
        RECT 70.975 8.280 72.320 9.720 ;
        RECT 73.730 12.390 73.960 12.485 ;
        RECT 74.205 12.390 74.695 14.445 ;
        RECT 75.265 12.920 75.900 12.925 ;
        RECT 75.150 12.690 79.110 12.920 ;
        RECT 74.870 12.390 75.100 12.485 ;
        RECT 73.730 8.565 75.100 12.390 ;
        RECT 73.730 8.485 73.960 8.565 ;
        RECT 74.870 8.485 75.100 8.565 ;
        RECT 76.525 8.280 77.870 12.690 ;
        RECT 79.160 12.420 79.390 12.485 ;
        RECT 80.045 12.425 80.520 17.260 ;
        RECT 81.845 16.455 82.525 17.260 ;
        RECT 82.945 16.735 83.280 16.985 ;
        RECT 82.960 16.710 83.250 16.735 ;
        RECT 86.420 16.635 88.330 17.260 ;
        RECT 90.420 16.925 92.305 16.930 ;
        RECT 93.865 16.925 95.750 16.930 ;
        RECT 90.410 16.695 92.370 16.925 ;
        RECT 93.840 16.695 95.800 16.925 ;
        RECT 82.770 16.455 83.000 16.505 ;
        RECT 81.845 15.955 83.000 16.455 ;
        RECT 80.915 12.735 81.250 12.985 ;
        RECT 80.935 12.705 81.225 12.735 ;
        RECT 80.745 12.425 80.975 12.500 ;
        RECT 79.160 8.485 79.615 12.420 ;
        RECT 80.045 11.680 80.975 12.425 ;
        RECT 80.380 8.565 80.975 11.680 ;
        RECT 80.745 8.500 80.975 8.565 ;
        RECT 81.185 12.475 81.415 12.500 ;
        RECT 81.185 8.920 81.695 12.475 ;
        RECT 81.185 8.550 81.880 8.920 ;
        RECT 82.380 8.600 83.000 15.955 ;
        RECT 81.185 8.500 81.415 8.550 ;
        RECT 69.720 8.250 73.680 8.280 ;
        RECT 75.150 8.250 79.110 8.280 ;
        RECT 69.720 8.090 79.110 8.250 ;
        RECT 69.720 8.050 73.680 8.090 ;
        RECT 75.150 8.050 79.110 8.090 ;
        RECT 79.275 6.660 79.615 8.485 ;
        RECT 80.925 6.660 81.345 8.305 ;
        RECT 79.275 6.505 81.345 6.660 ;
        RECT 79.350 6.390 81.345 6.505 ;
        RECT 69.810 6.125 73.770 6.355 ;
        RECT 75.240 6.125 79.200 6.355 ;
        RECT 69.245 5.205 69.760 5.965 ;
        RECT 69.315 4.025 69.760 5.205 ;
        RECT 69.530 3.965 69.760 4.025 ;
        RECT 71.190 3.805 72.145 6.125 ;
        RECT 73.820 5.900 74.050 5.965 ;
        RECT 74.960 5.900 75.190 5.965 ;
        RECT 73.820 4.030 75.190 5.900 ;
        RECT 73.820 3.965 74.050 4.030 ;
        RECT 68.755 3.255 68.945 3.785 ;
        RECT 69.810 3.575 73.770 3.805 ;
        RECT 74.225 3.255 74.780 4.030 ;
        RECT 74.960 3.965 75.190 4.030 ;
        RECT 76.635 3.805 77.590 6.125 ;
        RECT 79.350 5.970 79.615 6.390 ;
        RECT 80.925 6.115 81.345 6.390 ;
        RECT 81.580 7.355 81.880 8.550 ;
        RECT 82.770 8.505 83.000 8.600 ;
        RECT 83.210 16.430 83.440 16.505 ;
        RECT 83.210 9.110 83.985 16.430 ;
        RECT 86.385 16.405 88.385 16.635 ;
        RECT 90.130 16.410 90.360 16.490 ;
        RECT 85.950 13.060 86.180 16.355 ;
        RECT 88.590 16.275 88.820 16.355 ;
        RECT 88.560 13.060 88.820 16.275 ;
        RECT 85.950 11.245 88.820 13.060 ;
        RECT 83.210 8.580 84.060 9.110 ;
        RECT 85.950 8.825 86.180 11.245 ;
        RECT 83.210 8.505 83.440 8.580 ;
        RECT 82.875 7.825 83.390 8.315 ;
        RECT 82.875 7.360 83.385 7.825 ;
        RECT 83.690 7.795 84.060 8.580 ;
        RECT 85.590 8.395 86.180 8.825 ;
        RECT 87.075 8.640 87.335 8.960 ;
        RECT 88.560 8.645 88.820 11.245 ;
        RECT 89.890 8.990 90.360 16.410 ;
        RECT 90.850 9.775 91.740 16.695 ;
        RECT 92.420 16.390 92.650 16.490 ;
        RECT 92.420 16.380 92.775 16.390 ;
        RECT 93.560 16.380 93.790 16.490 ;
        RECT 87.130 8.480 87.280 8.640 ;
        RECT 82.510 7.355 83.385 7.360 ;
        RECT 81.580 6.950 83.385 7.355 ;
        RECT 81.580 6.110 81.880 6.950 ;
        RECT 82.510 6.935 83.385 6.950 ;
        RECT 82.875 6.825 83.385 6.935 ;
        RECT 82.875 6.125 83.390 6.825 ;
        RECT 83.615 6.795 84.645 7.795 ;
        RECT 79.275 5.965 79.615 5.970 ;
        RECT 79.250 4.020 79.615 5.965 ;
        RECT 80.830 5.900 81.060 5.970 ;
        RECT 80.335 5.230 81.060 5.900 ;
        RECT 80.325 5.040 81.060 5.230 ;
        RECT 80.325 4.240 80.680 5.040 ;
        RECT 80.830 4.970 81.060 5.040 ;
        RECT 81.270 5.925 81.500 5.970 ;
        RECT 81.640 5.925 81.880 6.110 ;
        RECT 81.270 5.595 81.880 5.925 ;
        RECT 82.855 5.870 83.085 5.975 ;
        RECT 81.270 5.040 81.765 5.595 ;
        RECT 81.270 4.970 81.500 5.040 ;
        RECT 81.020 4.785 81.310 4.810 ;
        RECT 81.005 4.535 81.340 4.785 ;
        RECT 82.625 4.765 83.085 5.870 ;
        RECT 82.305 4.240 83.085 4.765 ;
        RECT 79.885 4.060 83.085 4.240 ;
        RECT 79.250 3.965 79.480 4.020 ;
        RECT 75.240 3.575 79.200 3.805 ;
        RECT 79.885 3.620 82.690 4.060 ;
        RECT 82.855 3.975 83.085 4.060 ;
        RECT 83.295 5.910 83.525 5.975 ;
        RECT 83.690 5.910 84.060 6.795 ;
        RECT 83.295 5.585 84.060 5.910 ;
        RECT 83.295 4.045 84.055 5.585 ;
        RECT 83.295 3.975 83.525 4.045 ;
        RECT 83.045 3.795 83.335 3.815 ;
        RECT 79.885 3.255 82.350 3.620 ;
        RECT 83.020 3.545 83.355 3.795 ;
        RECT 85.590 3.280 86.085 8.395 ;
        RECT 87.105 8.345 87.310 8.480 ;
        RECT 88.590 8.395 88.820 8.645 ;
        RECT 89.610 8.550 90.360 8.990 ;
        RECT 90.780 8.775 91.795 9.775 ;
        RECT 86.385 8.115 88.385 8.345 ;
        RECT 89.610 6.355 89.980 8.550 ;
        RECT 90.130 8.490 90.360 8.550 ;
        RECT 90.850 8.285 91.740 8.775 ;
        RECT 92.420 8.580 93.790 16.380 ;
        RECT 94.325 11.635 95.215 16.695 ;
        RECT 95.850 16.410 96.080 16.490 ;
        RECT 94.320 10.015 95.220 11.635 ;
        RECT 94.325 9.605 95.215 10.015 ;
        RECT 94.250 8.605 95.280 9.605 ;
        RECT 95.850 8.625 96.225 16.410 ;
        RECT 96.500 16.025 98.180 17.260 ;
        RECT 99.015 16.025 103.940 16.035 ;
        RECT 96.500 15.545 103.940 16.025 ;
        RECT 96.500 13.285 98.180 15.545 ;
        RECT 99.015 15.125 103.940 15.545 ;
        RECT 98.520 14.935 98.775 14.960 ;
        RECT 98.520 14.920 98.795 14.935 ;
        RECT 98.490 14.645 98.825 14.920 ;
        RECT 99.000 14.895 104.000 15.125 ;
        RECT 104.210 14.935 104.465 14.960 ;
        RECT 98.520 14.630 98.775 14.645 ;
        RECT 99.000 14.455 104.000 14.685 ;
        RECT 104.205 14.645 104.465 14.935 ;
        RECT 104.210 14.630 104.465 14.645 ;
        RECT 99.045 14.445 103.900 14.455 ;
        RECT 99.045 12.920 101.690 12.925 ;
        RECT 97.720 12.720 101.690 12.920 ;
        RECT 97.720 12.690 101.680 12.720 ;
        RECT 96.560 12.335 96.895 12.610 ;
        RECT 97.440 12.440 97.670 12.485 ;
        RECT 92.420 8.560 92.775 8.580 ;
        RECT 92.420 8.490 92.650 8.560 ;
        RECT 93.560 8.490 93.790 8.580 ;
        RECT 94.320 8.465 95.230 8.605 ;
        RECT 95.850 8.490 96.240 8.625 ;
        RECT 94.310 8.285 95.320 8.465 ;
        RECT 90.410 8.055 92.370 8.285 ;
        RECT 93.840 8.055 95.800 8.285 ;
        RECT 91.095 6.975 91.495 8.055 ;
        RECT 93.865 8.050 95.750 8.055 ;
        RECT 96.045 6.355 96.240 8.490 ;
        RECT 96.630 6.830 96.820 12.335 ;
        RECT 97.250 11.105 97.670 12.440 ;
        RECT 98.975 11.105 100.320 12.690 ;
        RECT 97.250 9.720 100.320 11.105 ;
        RECT 97.250 8.990 97.670 9.720 ;
        RECT 97.245 8.485 97.670 8.990 ;
        RECT 96.630 6.640 96.945 6.830 ;
        RECT 86.950 6.125 90.910 6.355 ;
        RECT 92.380 6.125 96.340 6.355 ;
        RECT 96.755 6.130 96.945 6.640 ;
        RECT 86.670 5.515 86.900 5.965 ;
        RECT 88.150 5.515 88.940 6.125 ;
        RECT 86.670 5.210 88.940 5.515 ;
        RECT 86.615 5.195 88.940 5.210 ;
        RECT 86.530 4.350 88.940 5.195 ;
        RECT 86.530 3.975 86.900 4.350 ;
        RECT 86.670 3.965 86.900 3.975 ;
        RECT 88.150 3.805 88.940 4.350 ;
        RECT 90.960 5.880 91.190 5.965 ;
        RECT 92.100 5.880 92.330 5.965 ;
        RECT 90.960 4.055 92.330 5.880 ;
        RECT 90.960 3.965 91.190 4.055 ;
        RECT 86.950 3.575 90.910 3.805 ;
        RECT 83.890 3.255 86.085 3.280 ;
        RECT 86.530 3.255 86.755 3.265 ;
        RECT 91.430 3.255 91.920 4.055 ;
        RECT 92.100 3.965 92.330 4.055 ;
        RECT 93.815 5.745 95.155 6.125 ;
        RECT 96.390 5.745 96.620 5.965 ;
        RECT 93.815 4.150 96.620 5.745 ;
        RECT 93.815 3.805 95.155 4.150 ;
        RECT 96.390 3.965 96.620 4.150 ;
        RECT 92.380 3.575 96.340 3.805 ;
        RECT 96.770 3.785 96.945 6.130 ;
        RECT 97.245 5.965 97.540 8.485 ;
        RECT 98.975 8.280 100.320 9.720 ;
        RECT 101.730 12.390 101.960 12.485 ;
        RECT 102.205 12.390 102.695 14.445 ;
        RECT 103.265 12.920 103.900 12.925 ;
        RECT 103.150 12.690 107.110 12.920 ;
        RECT 102.870 12.390 103.100 12.485 ;
        RECT 101.730 8.565 103.100 12.390 ;
        RECT 101.730 8.485 101.960 8.565 ;
        RECT 102.870 8.485 103.100 8.565 ;
        RECT 104.525 8.280 105.870 12.690 ;
        RECT 107.160 12.420 107.390 12.485 ;
        RECT 108.045 12.425 108.520 17.260 ;
        RECT 109.845 16.455 110.525 17.260 ;
        RECT 110.945 16.735 111.280 16.985 ;
        RECT 110.960 16.710 111.250 16.735 ;
        RECT 114.420 16.635 116.330 17.260 ;
        RECT 118.420 16.925 120.305 16.930 ;
        RECT 121.865 16.925 123.750 16.930 ;
        RECT 118.410 16.695 120.370 16.925 ;
        RECT 121.840 16.695 123.800 16.925 ;
        RECT 110.770 16.455 111.000 16.505 ;
        RECT 109.845 15.955 111.000 16.455 ;
        RECT 108.915 12.735 109.250 12.985 ;
        RECT 108.935 12.705 109.225 12.735 ;
        RECT 108.745 12.425 108.975 12.500 ;
        RECT 107.160 8.485 107.615 12.420 ;
        RECT 108.045 11.680 108.975 12.425 ;
        RECT 108.380 8.565 108.975 11.680 ;
        RECT 108.745 8.500 108.975 8.565 ;
        RECT 109.185 12.475 109.415 12.500 ;
        RECT 109.185 8.920 109.695 12.475 ;
        RECT 109.185 8.550 109.880 8.920 ;
        RECT 110.380 8.600 111.000 15.955 ;
        RECT 109.185 8.500 109.415 8.550 ;
        RECT 97.720 8.250 101.680 8.280 ;
        RECT 103.150 8.250 107.110 8.280 ;
        RECT 97.720 8.090 107.110 8.250 ;
        RECT 97.720 8.050 101.680 8.090 ;
        RECT 103.150 8.050 107.110 8.090 ;
        RECT 107.275 6.660 107.615 8.485 ;
        RECT 108.925 6.660 109.345 8.305 ;
        RECT 107.275 6.505 109.345 6.660 ;
        RECT 107.350 6.390 109.345 6.505 ;
        RECT 97.810 6.125 101.770 6.355 ;
        RECT 103.240 6.125 107.200 6.355 ;
        RECT 97.245 5.205 97.760 5.965 ;
        RECT 97.315 4.025 97.760 5.205 ;
        RECT 97.530 3.965 97.760 4.025 ;
        RECT 99.190 3.805 100.145 6.125 ;
        RECT 101.820 5.900 102.050 5.965 ;
        RECT 102.960 5.900 103.190 5.965 ;
        RECT 101.820 4.030 103.190 5.900 ;
        RECT 101.820 3.965 102.050 4.030 ;
        RECT 96.755 3.255 96.945 3.785 ;
        RECT 97.810 3.575 101.770 3.805 ;
        RECT 102.225 3.255 102.780 4.030 ;
        RECT 102.960 3.965 103.190 4.030 ;
        RECT 104.635 3.805 105.590 6.125 ;
        RECT 107.350 5.970 107.615 6.390 ;
        RECT 108.925 6.115 109.345 6.390 ;
        RECT 109.580 7.355 109.880 8.550 ;
        RECT 110.770 8.505 111.000 8.600 ;
        RECT 111.210 16.430 111.440 16.505 ;
        RECT 111.210 9.110 111.985 16.430 ;
        RECT 114.385 16.405 116.385 16.635 ;
        RECT 118.130 16.410 118.360 16.490 ;
        RECT 113.950 13.060 114.180 16.355 ;
        RECT 116.590 16.275 116.820 16.355 ;
        RECT 116.560 13.060 116.820 16.275 ;
        RECT 113.950 11.245 116.820 13.060 ;
        RECT 111.210 8.580 112.060 9.110 ;
        RECT 113.950 8.825 114.180 11.245 ;
        RECT 111.210 8.505 111.440 8.580 ;
        RECT 110.875 7.825 111.390 8.315 ;
        RECT 110.875 7.360 111.385 7.825 ;
        RECT 111.690 7.795 112.060 8.580 ;
        RECT 113.590 8.395 114.180 8.825 ;
        RECT 115.075 8.640 115.335 8.960 ;
        RECT 116.560 8.645 116.820 11.245 ;
        RECT 117.890 8.990 118.360 16.410 ;
        RECT 118.850 9.775 119.740 16.695 ;
        RECT 120.420 16.390 120.650 16.490 ;
        RECT 120.420 16.380 120.775 16.390 ;
        RECT 121.560 16.380 121.790 16.490 ;
        RECT 115.130 8.480 115.280 8.640 ;
        RECT 110.510 7.355 111.385 7.360 ;
        RECT 109.580 6.950 111.385 7.355 ;
        RECT 109.580 6.110 109.880 6.950 ;
        RECT 110.510 6.935 111.385 6.950 ;
        RECT 110.875 6.825 111.385 6.935 ;
        RECT 110.875 6.125 111.390 6.825 ;
        RECT 111.615 6.795 112.645 7.795 ;
        RECT 107.275 5.965 107.615 5.970 ;
        RECT 107.250 4.020 107.615 5.965 ;
        RECT 108.830 5.900 109.060 5.970 ;
        RECT 108.335 5.230 109.060 5.900 ;
        RECT 108.325 5.040 109.060 5.230 ;
        RECT 108.325 4.240 108.680 5.040 ;
        RECT 108.830 4.970 109.060 5.040 ;
        RECT 109.270 5.925 109.500 5.970 ;
        RECT 109.640 5.925 109.880 6.110 ;
        RECT 109.270 5.595 109.880 5.925 ;
        RECT 110.855 5.870 111.085 5.975 ;
        RECT 109.270 5.040 109.765 5.595 ;
        RECT 109.270 4.970 109.500 5.040 ;
        RECT 109.020 4.785 109.310 4.810 ;
        RECT 109.005 4.535 109.340 4.785 ;
        RECT 110.625 4.765 111.085 5.870 ;
        RECT 110.305 4.240 111.085 4.765 ;
        RECT 107.885 4.060 111.085 4.240 ;
        RECT 107.250 3.965 107.480 4.020 ;
        RECT 103.240 3.575 107.200 3.805 ;
        RECT 107.885 3.620 110.690 4.060 ;
        RECT 110.855 3.975 111.085 4.060 ;
        RECT 111.295 5.910 111.525 5.975 ;
        RECT 111.690 5.910 112.060 6.795 ;
        RECT 111.295 5.585 112.060 5.910 ;
        RECT 111.295 4.045 112.055 5.585 ;
        RECT 111.295 3.975 111.525 4.045 ;
        RECT 111.045 3.795 111.335 3.815 ;
        RECT 107.885 3.255 110.350 3.620 ;
        RECT 111.020 3.545 111.355 3.795 ;
        RECT 113.590 3.280 114.085 8.395 ;
        RECT 115.105 8.345 115.310 8.480 ;
        RECT 116.590 8.395 116.820 8.645 ;
        RECT 117.610 8.550 118.360 8.990 ;
        RECT 118.780 8.775 119.795 9.775 ;
        RECT 114.385 8.115 116.385 8.345 ;
        RECT 117.610 6.355 117.980 8.550 ;
        RECT 118.130 8.490 118.360 8.550 ;
        RECT 118.850 8.285 119.740 8.775 ;
        RECT 120.420 8.580 121.790 16.380 ;
        RECT 122.325 11.635 123.215 16.695 ;
        RECT 123.850 16.410 124.080 16.490 ;
        RECT 122.320 10.015 123.220 11.635 ;
        RECT 122.325 9.605 123.215 10.015 ;
        RECT 122.250 8.605 123.280 9.605 ;
        RECT 123.850 8.625 124.225 16.410 ;
        RECT 124.500 16.025 126.180 17.260 ;
        RECT 127.015 16.025 131.940 16.035 ;
        RECT 124.500 15.545 131.940 16.025 ;
        RECT 124.500 13.285 126.180 15.545 ;
        RECT 127.015 15.125 131.940 15.545 ;
        RECT 126.520 14.935 126.775 14.960 ;
        RECT 126.520 14.920 126.795 14.935 ;
        RECT 126.490 14.645 126.825 14.920 ;
        RECT 127.000 14.895 132.000 15.125 ;
        RECT 132.210 14.935 132.465 14.960 ;
        RECT 126.520 14.630 126.775 14.645 ;
        RECT 127.000 14.455 132.000 14.685 ;
        RECT 132.205 14.645 132.465 14.935 ;
        RECT 132.210 14.630 132.465 14.645 ;
        RECT 127.045 14.445 131.900 14.455 ;
        RECT 127.045 12.920 129.690 12.925 ;
        RECT 125.720 12.720 129.690 12.920 ;
        RECT 125.720 12.690 129.680 12.720 ;
        RECT 124.560 12.335 124.895 12.610 ;
        RECT 125.440 12.440 125.670 12.485 ;
        RECT 120.420 8.560 120.775 8.580 ;
        RECT 120.420 8.490 120.650 8.560 ;
        RECT 121.560 8.490 121.790 8.580 ;
        RECT 122.320 8.465 123.230 8.605 ;
        RECT 123.850 8.490 124.240 8.625 ;
        RECT 122.310 8.285 123.320 8.465 ;
        RECT 118.410 8.055 120.370 8.285 ;
        RECT 121.840 8.055 123.800 8.285 ;
        RECT 119.150 7.155 119.435 8.055 ;
        RECT 121.865 8.050 123.750 8.055 ;
        RECT 124.045 6.355 124.240 8.490 ;
        RECT 124.630 6.830 124.820 12.335 ;
        RECT 125.250 11.105 125.670 12.440 ;
        RECT 126.975 11.105 128.320 12.690 ;
        RECT 125.250 9.720 128.320 11.105 ;
        RECT 125.250 8.990 125.670 9.720 ;
        RECT 125.245 8.485 125.670 8.990 ;
        RECT 124.630 6.640 124.945 6.830 ;
        RECT 114.950 6.125 118.910 6.355 ;
        RECT 120.380 6.125 124.340 6.355 ;
        RECT 124.755 6.130 124.945 6.640 ;
        RECT 114.670 5.515 114.900 5.965 ;
        RECT 116.150 5.515 116.940 6.125 ;
        RECT 114.670 5.210 116.940 5.515 ;
        RECT 114.615 5.195 116.940 5.210 ;
        RECT 114.530 4.350 116.940 5.195 ;
        RECT 114.530 3.975 114.900 4.350 ;
        RECT 114.670 3.965 114.900 3.975 ;
        RECT 116.150 3.805 116.940 4.350 ;
        RECT 118.960 5.880 119.190 5.965 ;
        RECT 120.100 5.880 120.330 5.965 ;
        RECT 118.960 4.055 120.330 5.880 ;
        RECT 118.960 3.965 119.190 4.055 ;
        RECT 114.950 3.575 118.910 3.805 ;
        RECT 111.590 3.255 114.085 3.280 ;
        RECT 114.530 3.255 114.755 3.265 ;
        RECT 119.430 3.255 119.920 4.055 ;
        RECT 120.100 3.965 120.330 4.055 ;
        RECT 121.815 5.745 123.155 6.125 ;
        RECT 124.390 5.745 124.620 5.965 ;
        RECT 121.815 4.150 124.620 5.745 ;
        RECT 121.815 3.805 123.155 4.150 ;
        RECT 124.390 3.965 124.620 4.150 ;
        RECT 120.380 3.575 124.340 3.805 ;
        RECT 124.770 3.785 124.945 6.130 ;
        RECT 125.245 5.965 125.540 8.485 ;
        RECT 126.975 8.280 128.320 9.720 ;
        RECT 129.730 12.390 129.960 12.485 ;
        RECT 130.205 12.390 130.695 14.445 ;
        RECT 131.265 12.920 131.900 12.925 ;
        RECT 131.150 12.690 135.110 12.920 ;
        RECT 130.870 12.390 131.100 12.485 ;
        RECT 129.730 8.565 131.100 12.390 ;
        RECT 129.730 8.485 129.960 8.565 ;
        RECT 130.870 8.485 131.100 8.565 ;
        RECT 132.525 8.280 133.870 12.690 ;
        RECT 135.160 12.420 135.390 12.485 ;
        RECT 136.045 12.425 136.520 17.260 ;
        RECT 137.845 16.455 138.525 17.260 ;
        RECT 138.945 16.735 139.280 16.985 ;
        RECT 138.960 16.710 139.250 16.735 ;
        RECT 138.770 16.455 139.000 16.505 ;
        RECT 137.845 15.955 139.000 16.455 ;
        RECT 136.915 12.735 137.250 12.985 ;
        RECT 136.935 12.705 137.225 12.735 ;
        RECT 136.745 12.425 136.975 12.500 ;
        RECT 135.160 8.485 135.615 12.420 ;
        RECT 136.045 11.680 136.975 12.425 ;
        RECT 136.380 8.565 136.975 11.680 ;
        RECT 136.745 8.500 136.975 8.565 ;
        RECT 137.185 12.475 137.415 12.500 ;
        RECT 137.185 8.920 137.695 12.475 ;
        RECT 137.185 8.550 137.880 8.920 ;
        RECT 138.380 8.600 139.000 15.955 ;
        RECT 137.185 8.500 137.415 8.550 ;
        RECT 125.720 8.250 129.680 8.280 ;
        RECT 131.150 8.250 135.110 8.280 ;
        RECT 125.720 8.090 135.110 8.250 ;
        RECT 125.720 8.050 129.680 8.090 ;
        RECT 131.150 8.050 135.110 8.090 ;
        RECT 135.275 6.660 135.615 8.485 ;
        RECT 136.925 6.660 137.345 8.305 ;
        RECT 135.275 6.505 137.345 6.660 ;
        RECT 135.350 6.390 137.345 6.505 ;
        RECT 125.810 6.125 129.770 6.355 ;
        RECT 131.240 6.125 135.200 6.355 ;
        RECT 125.245 5.205 125.760 5.965 ;
        RECT 125.315 4.025 125.760 5.205 ;
        RECT 125.530 3.965 125.760 4.025 ;
        RECT 127.190 3.805 128.145 6.125 ;
        RECT 129.820 5.900 130.050 5.965 ;
        RECT 130.960 5.900 131.190 5.965 ;
        RECT 129.820 4.030 131.190 5.900 ;
        RECT 129.820 3.965 130.050 4.030 ;
        RECT 124.755 3.255 124.945 3.785 ;
        RECT 125.810 3.575 129.770 3.805 ;
        RECT 130.225 3.255 130.780 4.030 ;
        RECT 130.960 3.965 131.190 4.030 ;
        RECT 132.635 3.805 133.590 6.125 ;
        RECT 135.350 5.970 135.615 6.390 ;
        RECT 136.925 6.115 137.345 6.390 ;
        RECT 137.580 7.355 137.880 8.550 ;
        RECT 138.770 8.505 139.000 8.600 ;
        RECT 139.210 16.430 139.440 16.505 ;
        RECT 139.210 9.110 139.985 16.430 ;
        RECT 139.210 8.580 140.060 9.110 ;
        RECT 139.210 8.505 139.440 8.580 ;
        RECT 138.875 7.825 139.390 8.315 ;
        RECT 138.875 7.360 139.385 7.825 ;
        RECT 139.690 7.795 140.060 8.580 ;
        RECT 138.510 7.355 139.385 7.360 ;
        RECT 137.580 6.950 139.385 7.355 ;
        RECT 137.580 6.110 137.880 6.950 ;
        RECT 138.510 6.935 139.385 6.950 ;
        RECT 138.875 6.825 139.385 6.935 ;
        RECT 138.875 6.125 139.390 6.825 ;
        RECT 139.615 6.795 140.645 7.795 ;
        RECT 135.275 5.965 135.615 5.970 ;
        RECT 135.250 4.020 135.615 5.965 ;
        RECT 136.830 5.900 137.060 5.970 ;
        RECT 136.335 5.230 137.060 5.900 ;
        RECT 136.325 5.040 137.060 5.230 ;
        RECT 136.325 4.240 136.680 5.040 ;
        RECT 136.830 4.970 137.060 5.040 ;
        RECT 137.270 5.925 137.500 5.970 ;
        RECT 137.640 5.925 137.880 6.110 ;
        RECT 137.270 5.595 137.880 5.925 ;
        RECT 138.855 5.870 139.085 5.975 ;
        RECT 137.270 5.040 137.765 5.595 ;
        RECT 137.270 4.970 137.500 5.040 ;
        RECT 137.020 4.785 137.310 4.810 ;
        RECT 137.005 4.535 137.340 4.785 ;
        RECT 138.625 4.765 139.085 5.870 ;
        RECT 138.305 4.240 139.085 4.765 ;
        RECT 135.885 4.060 139.085 4.240 ;
        RECT 135.250 3.965 135.480 4.020 ;
        RECT 131.240 3.575 135.200 3.805 ;
        RECT 135.885 3.620 138.690 4.060 ;
        RECT 138.855 3.975 139.085 4.060 ;
        RECT 139.295 5.910 139.525 5.975 ;
        RECT 139.690 5.910 140.060 6.795 ;
        RECT 139.295 5.585 140.060 5.910 ;
        RECT 139.295 4.045 140.055 5.585 ;
        RECT 139.295 3.975 139.525 4.045 ;
        RECT 139.045 3.795 139.335 3.815 ;
        RECT 135.885 3.255 138.350 3.620 ;
        RECT 139.020 3.545 139.355 3.795 ;
        RECT 1.475 2.380 140.080 3.255 ;
      LAYER met2 ;
        RECT 63.150 206.840 63.430 207.340 ;
        RECT 66.370 206.840 66.650 207.340 ;
        RECT 72.810 206.840 73.090 207.340 ;
        RECT 76.030 206.840 76.310 207.340 ;
        RECT 79.250 206.840 79.530 207.340 ;
        RECT 82.470 206.840 82.750 207.340 ;
        RECT 85.690 206.840 85.970 207.340 ;
        RECT 88.910 206.840 89.190 207.340 ;
        RECT 92.130 206.840 92.410 207.340 ;
        RECT 95.350 206.840 95.630 207.340 ;
        RECT 98.570 206.840 98.850 207.340 ;
        RECT 24.510 195.045 24.790 195.415 ;
        RECT 24.580 193.520 24.720 195.045 ;
        RECT 42.350 194.705 43.890 195.075 ;
        RECT 63.220 193.860 63.360 206.840 ;
        RECT 66.440 194.540 66.580 206.840 ;
        RECT 66.380 194.220 66.640 194.540 ;
        RECT 72.880 193.860 73.020 206.840 ;
        RECT 76.100 194.540 76.240 206.840 ;
        RECT 76.040 194.220 76.300 194.540 ;
        RECT 79.320 193.860 79.460 206.840 ;
        RECT 82.540 193.860 82.680 206.840 ;
        RECT 85.760 194.540 85.900 206.840 ;
        RECT 88.980 195.560 89.120 206.840 ;
        RECT 88.920 195.240 89.180 195.560 ;
        RECT 92.200 194.540 92.340 206.840 ;
        RECT 93.060 195.240 93.320 195.560 ;
        RECT 85.700 194.220 85.960 194.540 ;
        RECT 92.140 194.220 92.400 194.540 ;
        RECT 93.120 193.860 93.260 195.240 ;
        RECT 95.420 194.540 95.560 206.840 ;
        RECT 98.640 196.660 98.780 206.840 ;
        RECT 99.040 206.800 99.300 207.120 ;
        RECT 101.790 206.840 102.070 207.340 ;
        RECT 105.010 206.840 105.290 207.340 ;
        RECT 108.230 206.840 108.510 207.340 ;
        RECT 111.450 206.840 111.730 207.340 ;
        RECT 114.670 206.840 114.950 207.340 ;
        RECT 117.890 206.860 118.170 207.340 ;
        RECT 118.420 207.020 119.480 207.160 ;
        RECT 118.420 206.860 118.560 207.020 ;
        RECT 117.890 206.840 118.560 206.860 ;
        RECT 98.180 196.520 98.780 196.660 ;
        RECT 95.360 194.220 95.620 194.540 ;
        RECT 93.980 193.880 94.240 194.200 ;
        RECT 27.740 193.540 28.000 193.860 ;
        RECT 34.640 193.540 34.900 193.860 ;
        RECT 41.540 193.540 41.800 193.860 ;
        RECT 63.160 193.540 63.420 193.860 ;
        RECT 67.760 193.540 68.020 193.860 ;
        RECT 72.820 193.540 73.080 193.860 ;
        RECT 79.260 193.540 79.520 193.860 ;
        RECT 81.560 193.540 81.820 193.860 ;
        RECT 82.480 193.540 82.740 193.860 ;
        RECT 87.540 193.540 87.800 193.860 ;
        RECT 91.220 193.540 91.480 193.860 ;
        RECT 93.060 193.540 93.320 193.860 ;
        RECT 24.520 193.200 24.780 193.520 ;
        RECT 19.920 192.520 20.180 192.840 ;
        RECT 19.980 192.015 20.120 192.520 ;
        RECT 19.910 191.645 20.190 192.015 ;
        RECT 27.800 191.820 27.940 193.540 ;
        RECT 27.740 191.500 28.000 191.820 ;
        RECT 34.700 190.800 34.840 193.540 ;
        RECT 38.320 192.520 38.580 192.840 ;
        RECT 38.380 191.820 38.520 192.520 ;
        RECT 39.050 191.985 40.590 192.355 ;
        RECT 38.320 191.500 38.580 191.820 ;
        RECT 26.360 190.480 26.620 190.800 ;
        RECT 34.640 190.480 34.900 190.800 ;
        RECT 19.920 189.800 20.180 190.120 ;
        RECT 19.980 188.615 20.120 189.800 ;
        RECT 26.420 189.100 26.560 190.480 ;
        RECT 26.360 188.780 26.620 189.100 ;
        RECT 19.910 188.245 20.190 188.615 ;
        RECT 34.700 185.360 34.840 190.480 ;
        RECT 41.080 190.140 41.340 190.460 ;
        RECT 40.620 189.800 40.880 190.120 ;
        RECT 40.680 189.100 40.820 189.800 ;
        RECT 40.620 188.780 40.880 189.100 ;
        RECT 41.140 188.420 41.280 190.140 ;
        RECT 41.080 188.100 41.340 188.420 ;
        RECT 38.320 187.080 38.580 187.400 ;
        RECT 34.180 185.040 34.440 185.360 ;
        RECT 34.640 185.215 34.900 185.360 ;
        RECT 34.240 183.660 34.380 185.040 ;
        RECT 34.630 184.845 34.910 185.215 ;
        RECT 36.940 184.700 37.200 185.020 ;
        RECT 37.000 183.660 37.140 184.700 ;
        RECT 34.180 183.340 34.440 183.660 ;
        RECT 36.940 183.340 37.200 183.660 ;
        RECT 37.000 180.940 37.140 183.340 ;
        RECT 38.380 183.320 38.520 187.080 ;
        RECT 39.050 186.545 40.590 186.915 ;
        RECT 38.780 184.360 39.040 184.680 ;
        RECT 38.840 183.660 38.980 184.360 ;
        RECT 38.780 183.340 39.040 183.660 ;
        RECT 38.320 183.000 38.580 183.320 ;
        RECT 37.400 182.660 37.660 182.980 ;
        RECT 36.940 180.620 37.200 180.940 ;
        RECT 34.640 180.280 34.900 180.600 ;
        RECT 19.920 179.600 20.180 179.920 ;
        RECT 27.740 179.600 28.000 179.920 ;
        RECT 19.980 178.415 20.120 179.600 ;
        RECT 19.910 178.045 20.190 178.415 ;
        RECT 26.360 177.220 26.620 177.540 ;
        RECT 19.000 176.200 19.260 176.520 ;
        RECT 19.060 175.015 19.200 176.200 ;
        RECT 18.990 174.645 19.270 175.015 ;
        RECT 25.900 174.160 26.160 174.480 ;
        RECT 25.960 172.780 26.100 174.160 ;
        RECT 26.420 172.780 26.560 177.220 ;
        RECT 27.800 175.500 27.940 179.600 ;
        RECT 27.740 175.180 28.000 175.500 ;
        RECT 27.800 174.820 27.940 175.180 ;
        RECT 34.700 175.160 34.840 180.280 ;
        RECT 36.940 179.600 37.200 179.920 ;
        RECT 34.640 174.840 34.900 175.160 ;
        RECT 27.740 174.500 28.000 174.820 ;
        RECT 34.700 174.480 34.840 174.840 ;
        RECT 34.640 174.160 34.900 174.480 ;
        RECT 28.660 173.480 28.920 173.800 ;
        RECT 33.260 173.480 33.520 173.800 ;
        RECT 25.900 172.460 26.160 172.780 ;
        RECT 26.360 172.460 26.620 172.780 ;
        RECT 28.720 172.100 28.860 173.480 ;
        RECT 33.320 172.295 33.460 173.480 ;
        RECT 21.760 171.780 22.020 172.100 ;
        RECT 28.660 171.780 28.920 172.100 ;
        RECT 33.250 171.925 33.530 172.295 ;
        RECT 34.700 172.100 34.840 174.160 ;
        RECT 35.560 173.480 35.820 173.800 ;
        RECT 34.640 171.780 34.900 172.100 ;
        RECT 21.820 171.615 21.960 171.780 ;
        RECT 21.750 171.245 22.030 171.615 ;
        RECT 35.620 171.420 35.760 173.480 ;
        RECT 37.000 172.295 37.140 179.600 ;
        RECT 37.460 179.240 37.600 182.660 ;
        RECT 39.050 181.105 40.590 181.475 ;
        RECT 41.140 180.940 41.280 188.100 ;
        RECT 41.600 187.740 41.740 193.540 ;
        RECT 42.000 193.200 42.260 193.520 ;
        RECT 42.060 189.010 42.200 193.200 ;
        RECT 45.220 192.860 45.480 193.180 ;
        RECT 44.760 190.820 45.020 191.140 ;
        RECT 43.840 190.370 44.100 190.460 ;
        RECT 43.840 190.230 44.500 190.370 ;
        RECT 43.840 190.140 44.100 190.230 ;
        RECT 42.350 189.265 43.890 189.635 ;
        RECT 42.060 188.870 42.660 189.010 ;
        RECT 42.520 188.860 42.660 188.870 ;
        RECT 42.520 188.760 43.580 188.860 ;
        RECT 42.520 188.720 43.640 188.760 ;
        RECT 43.380 188.440 43.640 188.720 ;
        RECT 41.540 187.420 41.800 187.740 ;
        RECT 42.920 187.080 43.180 187.400 ;
        RECT 42.980 185.360 43.120 187.080 ;
        RECT 43.440 185.700 43.580 188.440 ;
        RECT 43.380 185.380 43.640 185.700 ;
        RECT 42.920 185.040 43.180 185.360 ;
        RECT 42.000 184.360 42.260 184.680 ;
        RECT 42.060 183.570 42.200 184.360 ;
        RECT 42.350 183.825 43.890 184.195 ;
        RECT 42.060 183.430 43.120 183.570 ;
        RECT 42.980 182.980 43.120 183.430 ;
        RECT 42.000 182.660 42.260 182.980 ;
        RECT 42.460 182.660 42.720 182.980 ;
        RECT 42.920 182.660 43.180 182.980 ;
        RECT 41.080 180.620 41.340 180.940 ;
        RECT 40.160 179.940 40.420 180.260 ;
        RECT 38.780 179.600 39.040 179.920 ;
        RECT 37.400 178.920 37.660 179.240 ;
        RECT 37.460 177.200 37.600 178.920 ;
        RECT 38.320 177.620 38.580 177.880 ;
        RECT 38.840 177.620 38.980 179.600 ;
        RECT 38.320 177.560 38.980 177.620 ;
        RECT 38.380 177.480 38.980 177.560 ;
        RECT 37.400 176.880 37.660 177.200 ;
        RECT 36.930 171.925 37.210 172.295 ;
        RECT 35.560 171.100 35.820 171.420 ;
        RECT 21.760 168.215 22.020 168.360 ;
        RECT 21.750 167.845 22.030 168.215 ;
        RECT 37.460 166.660 37.600 176.880 ;
        RECT 37.860 176.200 38.120 176.520 ;
        RECT 37.920 173.800 38.060 176.200 ;
        RECT 38.380 175.410 38.520 177.480 ;
        RECT 39.700 177.220 39.960 177.540 ;
        RECT 39.760 176.520 39.900 177.220 ;
        RECT 40.220 176.520 40.360 179.940 ;
        RECT 41.080 179.775 41.340 179.920 ;
        RECT 41.070 179.405 41.350 179.775 ;
        RECT 41.540 179.260 41.800 179.580 ;
        RECT 41.080 177.560 41.340 177.880 ;
        RECT 39.700 176.200 39.960 176.520 ;
        RECT 40.160 176.200 40.420 176.520 ;
        RECT 39.050 175.665 40.590 176.035 ;
        RECT 38.380 175.270 38.980 175.410 ;
        RECT 38.840 174.820 38.980 175.270 ;
        RECT 39.240 175.180 39.500 175.500 ;
        RECT 38.780 174.500 39.040 174.820 ;
        RECT 37.860 173.480 38.120 173.800 ;
        RECT 38.840 172.860 38.980 174.500 ;
        RECT 38.380 172.780 38.980 172.860 ;
        RECT 38.320 172.720 38.980 172.780 ;
        RECT 38.320 172.460 38.580 172.720 ;
        RECT 39.300 172.100 39.440 175.180 ;
        RECT 41.140 175.070 41.280 177.560 ;
        RECT 40.680 174.930 41.280 175.070 ;
        RECT 40.680 174.140 40.820 174.930 ;
        RECT 41.600 174.480 41.740 179.260 ;
        RECT 42.060 178.220 42.200 182.660 ;
        RECT 42.520 181.960 42.660 182.660 ;
        RECT 42.460 181.640 42.720 181.960 ;
        RECT 44.360 179.775 44.500 190.230 ;
        RECT 44.820 188.420 44.960 190.820 ;
        RECT 45.280 190.800 45.420 192.860 ;
        RECT 47.060 192.520 47.320 192.840 ;
        RECT 64.540 192.520 64.800 192.840 ;
        RECT 47.120 190.800 47.260 192.520 ;
        RECT 50.740 191.500 51.000 191.820 ;
        RECT 45.220 190.480 45.480 190.800 ;
        RECT 47.060 190.480 47.320 190.800 ;
        RECT 44.760 188.100 45.020 188.420 ;
        RECT 44.820 186.040 44.960 188.100 ;
        RECT 44.760 185.720 45.020 186.040 ;
        RECT 44.820 183.660 44.960 185.720 ;
        RECT 44.760 183.340 45.020 183.660 ;
        RECT 44.820 182.640 44.960 183.340 ;
        RECT 45.280 183.320 45.420 190.480 ;
        RECT 48.900 190.140 49.160 190.460 ;
        RECT 46.600 189.800 46.860 190.120 ;
        RECT 46.660 189.100 46.800 189.800 ;
        RECT 46.600 188.780 46.860 189.100 ;
        RECT 47.980 188.780 48.240 189.100 ;
        RECT 47.060 188.100 47.320 188.420 ;
        RECT 46.140 187.760 46.400 188.080 ;
        RECT 45.680 185.040 45.940 185.360 ;
        RECT 45.220 183.000 45.480 183.320 ;
        RECT 44.760 182.320 45.020 182.640 ;
        RECT 44.820 180.940 44.960 182.320 ;
        RECT 45.220 181.640 45.480 181.960 ;
        RECT 44.760 180.620 45.020 180.940 ;
        RECT 44.760 179.940 45.020 180.260 ;
        RECT 44.290 179.405 44.570 179.775 ;
        RECT 42.350 178.385 43.890 178.755 ;
        RECT 42.000 177.900 42.260 178.220 ;
        RECT 44.300 177.790 44.560 177.880 ;
        RECT 43.900 177.650 44.560 177.790 ;
        RECT 42.000 176.200 42.260 176.520 ;
        RECT 41.540 174.160 41.800 174.480 ;
        RECT 40.620 173.820 40.880 174.140 ;
        RECT 41.080 173.820 41.340 174.140 ;
        RECT 39.700 173.480 39.960 173.800 ;
        RECT 39.760 172.100 39.900 173.480 ;
        RECT 37.860 171.780 38.120 172.100 ;
        RECT 39.240 171.780 39.500 172.100 ;
        RECT 39.700 171.780 39.960 172.100 ;
        RECT 37.920 169.720 38.060 171.780 ;
        RECT 38.320 171.440 38.580 171.760 ;
        RECT 37.860 169.400 38.120 169.720 ;
        RECT 38.380 169.460 38.520 171.440 ;
        RECT 40.680 171.080 40.820 173.820 ;
        RECT 41.140 171.420 41.280 173.820 ;
        RECT 41.600 172.780 41.740 174.160 ;
        RECT 41.540 172.460 41.800 172.780 ;
        RECT 41.080 171.100 41.340 171.420 ;
        RECT 40.620 170.760 40.880 171.080 ;
        RECT 39.050 170.225 40.590 170.595 ;
        RECT 38.380 169.320 38.980 169.460 ;
        RECT 37.860 168.720 38.120 169.040 ;
        RECT 37.920 167.340 38.060 168.720 ;
        RECT 38.840 168.700 38.980 169.320 ;
        RECT 41.140 169.040 41.280 171.100 ;
        RECT 41.540 170.760 41.800 171.080 ;
        RECT 41.080 168.720 41.340 169.040 ;
        RECT 38.780 168.380 39.040 168.700 ;
        RECT 37.860 167.020 38.120 167.340 ;
        RECT 37.920 166.855 38.060 167.020 ;
        RECT 20.840 166.340 21.100 166.660 ;
        RECT 37.400 166.340 37.660 166.660 ;
        RECT 37.850 166.485 38.130 166.855 ;
        RECT 38.840 166.660 38.980 168.380 ;
        RECT 40.160 168.040 40.420 168.360 ;
        RECT 41.080 168.040 41.340 168.360 ;
        RECT 40.220 166.660 40.360 168.040 ;
        RECT 41.140 166.660 41.280 168.040 ;
        RECT 38.780 166.340 39.040 166.660 ;
        RECT 40.160 166.340 40.420 166.660 ;
        RECT 41.080 166.340 41.340 166.660 ;
        RECT 20.900 164.815 21.040 166.340 ;
        RECT 20.830 164.445 21.110 164.815 ;
        RECT 39.050 164.785 40.590 165.155 ;
        RECT 41.600 164.280 41.740 170.760 ;
        RECT 42.060 169.720 42.200 176.200 ;
        RECT 43.900 174.140 44.040 177.650 ;
        RECT 44.300 177.560 44.560 177.650 ;
        RECT 44.820 176.860 44.960 179.940 ;
        RECT 45.280 176.940 45.420 181.640 ;
        RECT 45.740 181.020 45.880 185.040 ;
        RECT 46.200 184.680 46.340 187.760 ;
        RECT 47.120 187.740 47.260 188.100 ;
        RECT 47.060 187.420 47.320 187.740 ;
        RECT 46.600 185.040 46.860 185.360 ;
        RECT 46.140 184.360 46.400 184.680 ;
        RECT 46.200 182.980 46.340 184.360 ;
        RECT 46.140 182.660 46.400 182.980 ;
        RECT 46.660 182.380 46.800 185.040 ;
        RECT 46.200 182.240 46.800 182.380 ;
        RECT 46.200 181.960 46.340 182.240 ;
        RECT 46.140 181.640 46.400 181.960 ;
        RECT 45.740 180.880 46.800 181.020 ;
        RECT 47.120 180.940 47.260 187.420 ;
        RECT 47.520 186.060 47.780 186.380 ;
        RECT 47.580 185.360 47.720 186.060 ;
        RECT 47.520 185.040 47.780 185.360 ;
        RECT 48.040 185.215 48.180 188.780 ;
        RECT 48.440 187.080 48.700 187.400 ;
        RECT 48.500 185.360 48.640 187.080 ;
        RECT 47.970 184.845 48.250 185.215 ;
        RECT 48.440 185.040 48.700 185.360 ;
        RECT 48.960 185.020 49.100 190.140 ;
        RECT 49.820 187.080 50.080 187.400 ;
        RECT 49.360 185.720 49.620 186.040 ;
        RECT 47.520 181.980 47.780 182.300 ;
        RECT 46.140 180.280 46.400 180.600 ;
        RECT 44.300 176.540 44.560 176.860 ;
        RECT 44.760 176.540 45.020 176.860 ;
        RECT 45.280 176.800 45.880 176.940 ;
        RECT 44.360 175.160 44.500 176.540 ;
        RECT 44.300 174.840 44.560 175.160 ;
        RECT 44.360 174.480 44.500 174.840 ;
        RECT 44.300 174.160 44.560 174.480 ;
        RECT 43.840 173.820 44.100 174.140 ;
        RECT 45.740 173.710 45.880 176.800 ;
        RECT 45.280 173.570 45.880 173.710 ;
        RECT 42.350 172.945 43.890 173.315 ;
        RECT 42.460 171.780 42.720 172.100 ;
        RECT 42.520 171.420 42.660 171.780 ;
        RECT 45.280 171.420 45.420 173.570 ;
        RECT 46.200 172.100 46.340 180.280 ;
        RECT 46.660 175.500 46.800 180.880 ;
        RECT 47.060 180.620 47.320 180.940 ;
        RECT 47.060 176.540 47.320 176.860 ;
        RECT 46.600 175.180 46.860 175.500 ;
        RECT 46.600 174.160 46.860 174.480 ;
        RECT 46.140 171.780 46.400 172.100 ;
        RECT 42.460 171.100 42.720 171.420 ;
        RECT 42.920 171.100 43.180 171.420 ;
        RECT 45.220 171.100 45.480 171.420 ;
        RECT 42.000 169.400 42.260 169.720 ;
        RECT 42.520 168.950 42.660 171.100 ;
        RECT 42.980 169.040 43.120 171.100 ;
        RECT 45.680 170.760 45.940 171.080 ;
        RECT 45.220 169.400 45.480 169.720 ;
        RECT 42.060 168.810 42.660 168.950 ;
        RECT 42.060 167.250 42.200 168.810 ;
        RECT 42.920 168.720 43.180 169.040 ;
        RECT 44.300 168.720 44.560 169.040 ;
        RECT 42.350 167.505 43.890 167.875 ;
        RECT 42.060 167.110 42.660 167.250 ;
        RECT 42.000 165.660 42.260 165.980 ;
        RECT 41.540 163.960 41.800 164.280 ;
        RECT 41.600 163.260 41.740 163.960 ;
        RECT 38.320 162.940 38.580 163.260 ;
        RECT 41.540 162.940 41.800 163.260 ;
        RECT 38.380 161.220 38.520 162.940 ;
        RECT 41.600 161.560 41.740 162.940 ;
        RECT 42.060 161.900 42.200 165.660 ;
        RECT 42.520 164.280 42.660 167.110 ;
        RECT 44.360 166.740 44.500 168.720 ;
        RECT 44.750 167.845 45.030 168.215 ;
        RECT 43.900 166.600 44.500 166.740 ;
        RECT 44.820 166.660 44.960 167.845 ;
        RECT 42.460 163.960 42.720 164.280 ;
        RECT 43.900 163.940 44.040 166.600 ;
        RECT 44.760 166.340 45.020 166.660 ;
        RECT 45.280 166.060 45.420 169.400 ;
        RECT 45.740 169.040 45.880 170.760 ;
        RECT 46.200 170.255 46.340 171.780 ;
        RECT 46.660 171.760 46.800 174.160 ;
        RECT 47.120 173.800 47.260 176.540 ;
        RECT 47.060 173.480 47.320 173.800 ;
        RECT 46.600 171.440 46.860 171.760 ;
        RECT 46.130 169.885 46.410 170.255 ;
        RECT 46.140 169.740 46.400 169.885 ;
        RECT 46.200 169.380 46.340 169.740 ;
        RECT 46.140 169.290 46.400 169.380 ;
        RECT 46.140 169.150 46.800 169.290 ;
        RECT 46.140 169.060 46.400 169.150 ;
        RECT 45.680 168.720 45.940 169.040 ;
        RECT 45.740 166.660 45.880 168.720 ;
        RECT 46.660 166.660 46.800 169.150 ;
        RECT 47.120 169.040 47.260 173.480 ;
        RECT 47.060 168.720 47.320 169.040 ;
        RECT 47.580 166.855 47.720 181.980 ;
        RECT 48.040 173.800 48.180 184.845 ;
        RECT 48.900 184.700 49.160 185.020 ;
        RECT 48.440 181.980 48.700 182.300 ;
        RECT 48.500 179.920 48.640 181.980 ;
        RECT 48.440 179.600 48.700 179.920 ;
        RECT 48.900 179.260 49.160 179.580 ;
        RECT 48.960 178.220 49.100 179.260 ;
        RECT 48.900 177.900 49.160 178.220 ;
        RECT 49.420 177.880 49.560 185.720 ;
        RECT 49.880 185.360 50.020 187.080 ;
        RECT 49.820 185.040 50.080 185.360 ;
        RECT 50.280 182.660 50.540 182.980 ;
        RECT 50.340 180.600 50.480 182.660 ;
        RECT 50.280 180.280 50.540 180.600 ;
        RECT 49.360 177.560 49.620 177.880 ;
        RECT 50.280 177.450 50.540 177.540 ;
        RECT 49.880 177.310 50.540 177.450 ;
        RECT 48.440 176.880 48.700 177.200 ;
        RECT 48.500 176.520 48.640 176.880 ;
        RECT 48.440 176.200 48.700 176.520 ;
        RECT 48.500 175.160 48.640 176.200 ;
        RECT 48.440 174.840 48.700 175.160 ;
        RECT 48.900 174.160 49.160 174.480 ;
        RECT 47.980 173.480 48.240 173.800 ;
        RECT 48.960 167.340 49.100 174.160 ;
        RECT 49.880 174.140 50.020 177.310 ;
        RECT 50.280 177.220 50.540 177.310 ;
        RECT 50.280 174.840 50.540 175.160 ;
        RECT 49.820 173.820 50.080 174.140 ;
        RECT 50.340 172.440 50.480 174.840 ;
        RECT 50.800 174.480 50.940 191.500 ;
        RECT 53.040 190.820 53.300 191.140 ;
        RECT 56.720 190.820 56.980 191.140 ;
        RECT 52.120 190.480 52.380 190.800 ;
        RECT 51.660 189.800 51.920 190.120 ;
        RECT 51.720 188.420 51.860 189.800 ;
        RECT 52.180 189.100 52.320 190.480 ;
        RECT 52.580 190.140 52.840 190.460 ;
        RECT 52.120 188.780 52.380 189.100 ;
        RECT 52.180 188.420 52.320 188.780 ;
        RECT 51.660 188.100 51.920 188.420 ;
        RECT 52.120 188.100 52.380 188.420 ;
        RECT 52.120 187.420 52.380 187.740 ;
        RECT 52.180 186.380 52.320 187.420 ;
        RECT 52.640 186.380 52.780 190.140 ;
        RECT 53.100 189.100 53.240 190.820 ;
        RECT 53.500 190.480 53.760 190.800 ;
        RECT 53.040 188.780 53.300 189.100 ;
        RECT 53.040 188.330 53.300 188.420 ;
        RECT 53.560 188.330 53.700 190.480 ;
        RECT 55.340 189.800 55.600 190.120 ;
        RECT 56.260 189.800 56.520 190.120 ;
        RECT 53.040 188.190 53.700 188.330 ;
        RECT 53.040 188.100 53.300 188.190 ;
        RECT 54.420 187.080 54.680 187.400 ;
        RECT 52.120 186.060 52.380 186.380 ;
        RECT 52.580 186.060 52.840 186.380 ;
        RECT 54.480 185.700 54.620 187.080 ;
        RECT 54.420 185.380 54.680 185.700 ;
        RECT 53.040 183.000 53.300 183.320 ;
        RECT 51.200 182.660 51.460 182.980 ;
        RECT 51.260 179.580 51.400 182.660 ;
        RECT 52.120 180.620 52.380 180.940 ;
        RECT 52.180 179.920 52.320 180.620 ;
        RECT 51.660 179.600 51.920 179.920 ;
        RECT 52.120 179.600 52.380 179.920 ;
        RECT 51.200 179.260 51.460 179.580 ;
        RECT 51.720 178.220 51.860 179.600 ;
        RECT 51.660 177.900 51.920 178.220 ;
        RECT 51.200 177.220 51.460 177.540 ;
        RECT 51.660 177.220 51.920 177.540 ;
        RECT 50.740 174.160 51.000 174.480 ;
        RECT 50.280 172.120 50.540 172.440 ;
        RECT 48.900 167.020 49.160 167.340 ;
        RECT 50.270 167.165 50.550 167.535 ;
        RECT 45.680 166.340 45.940 166.660 ;
        RECT 46.140 166.340 46.400 166.660 ;
        RECT 46.600 166.340 46.860 166.660 ;
        RECT 47.510 166.485 47.790 166.855 ;
        RECT 50.340 166.660 50.480 167.165 ;
        RECT 50.740 167.020 51.000 167.340 ;
        RECT 50.280 166.340 50.540 166.660 ;
        RECT 46.200 166.060 46.340 166.340 ;
        RECT 45.280 165.920 46.340 166.060 ;
        RECT 48.900 166.000 49.160 166.320 ;
        RECT 45.280 164.620 45.420 165.920 ;
        RECT 47.520 165.320 47.780 165.640 ;
        RECT 47.980 165.320 48.240 165.640 ;
        RECT 45.220 164.300 45.480 164.620 ;
        RECT 46.130 164.445 46.410 164.815 ;
        RECT 44.300 163.960 44.560 164.280 ;
        RECT 43.840 163.620 44.100 163.940 ;
        RECT 43.900 163.455 44.040 163.620 ;
        RECT 43.830 163.085 44.110 163.455 ;
        RECT 42.350 162.065 43.890 162.435 ;
        RECT 42.000 161.580 42.260 161.900 ;
        RECT 41.080 161.240 41.340 161.560 ;
        RECT 41.540 161.240 41.800 161.560 ;
        RECT 38.320 160.900 38.580 161.220 ;
        RECT 39.050 159.345 40.590 159.715 ;
        RECT 41.140 158.015 41.280 161.240 ;
        RECT 44.360 161.220 44.500 163.960 ;
        RECT 46.200 161.560 46.340 164.445 ;
        RECT 47.580 164.280 47.720 165.320 ;
        RECT 47.520 163.960 47.780 164.280 ;
        RECT 48.040 163.600 48.180 165.320 ;
        RECT 48.960 163.600 49.100 166.000 ;
        RECT 50.800 165.980 50.940 167.020 ;
        RECT 50.740 165.660 51.000 165.980 ;
        RECT 49.820 165.320 50.080 165.640 ;
        RECT 50.280 165.320 50.540 165.640 ;
        RECT 49.880 163.940 50.020 165.320 ;
        RECT 49.820 163.620 50.080 163.940 ;
        RECT 47.980 163.280 48.240 163.600 ;
        RECT 48.900 163.280 49.160 163.600 ;
        RECT 50.340 161.900 50.480 165.320 ;
        RECT 51.260 164.620 51.400 177.220 ;
        RECT 51.720 176.860 51.860 177.220 ;
        RECT 51.660 176.540 51.920 176.860 ;
        RECT 51.660 168.040 51.920 168.360 ;
        RECT 53.100 168.215 53.240 183.000 ;
        RECT 53.960 180.620 54.220 180.940 ;
        RECT 51.720 166.910 51.860 168.040 ;
        RECT 53.030 167.845 53.310 168.215 ;
        RECT 53.100 167.340 53.240 167.845 ;
        RECT 53.040 167.020 53.300 167.340 ;
        RECT 53.500 167.020 53.760 167.340 ;
        RECT 52.120 166.910 52.380 167.000 ;
        RECT 51.720 166.770 52.380 166.910 ;
        RECT 52.120 166.680 52.380 166.770 ;
        RECT 53.030 166.485 53.310 166.855 ;
        RECT 53.040 166.340 53.300 166.485 ;
        RECT 53.030 165.805 53.310 166.175 ;
        RECT 51.200 164.300 51.460 164.620 ;
        RECT 50.280 161.580 50.540 161.900 ;
        RECT 46.140 161.240 46.400 161.560 ;
        RECT 44.300 160.900 44.560 161.220 ;
        RECT 41.070 157.645 41.350 158.015 ;
        RECT 21.760 154.615 22.020 154.760 ;
        RECT 21.750 154.245 22.030 154.615 ;
        RECT 39.050 153.905 40.590 154.275 ;
        RECT 41.140 153.740 41.280 157.645 ;
        RECT 42.350 156.625 43.890 156.995 ;
        RECT 46.200 153.740 46.340 161.240 ;
        RECT 53.100 156.460 53.240 165.805 ;
        RECT 53.560 163.600 53.700 167.020 ;
        RECT 54.020 166.175 54.160 180.620 ;
        RECT 55.400 179.580 55.540 189.800 ;
        RECT 56.320 188.760 56.460 189.800 ;
        RECT 56.260 188.440 56.520 188.760 ;
        RECT 56.780 185.700 56.920 190.820 ;
        RECT 64.600 190.800 64.740 192.520 ;
        RECT 67.820 191.820 67.960 193.540 ;
        RECT 78.340 192.860 78.600 193.180 ;
        RECT 76.040 192.520 76.300 192.840 ;
        RECT 67.760 191.500 68.020 191.820 ;
        RECT 76.100 191.140 76.240 192.520 ;
        RECT 78.400 191.820 78.540 192.860 ;
        RECT 81.620 192.840 81.760 193.540 ;
        RECT 83.400 193.200 83.660 193.520 ;
        RECT 80.180 192.520 80.440 192.840 ;
        RECT 81.560 192.520 81.820 192.840 ;
        RECT 78.340 191.500 78.600 191.820 ;
        RECT 80.240 191.140 80.380 192.520 ;
        RECT 81.100 191.500 81.360 191.820 ;
        RECT 76.040 190.820 76.300 191.140 ;
        RECT 80.180 190.820 80.440 191.140 ;
        RECT 64.540 190.480 64.800 190.800 ;
        RECT 65.920 190.480 66.180 190.800 ;
        RECT 68.680 190.480 68.940 190.800 ;
        RECT 70.060 190.480 70.320 190.800 ;
        RECT 70.520 190.480 70.780 190.800 ;
        RECT 60.400 188.780 60.660 189.100 ;
        RECT 59.480 188.100 59.740 188.420 ;
        RECT 59.540 185.780 59.680 188.100 ;
        RECT 60.460 186.380 60.600 188.780 ;
        RECT 61.320 188.100 61.580 188.420 ;
        RECT 62.700 188.100 62.960 188.420 ;
        RECT 64.080 188.100 64.340 188.420 ;
        RECT 60.400 186.060 60.660 186.380 ;
        RECT 56.720 185.380 56.980 185.700 ;
        RECT 59.540 185.640 60.600 185.780 ;
        RECT 56.780 183.660 56.920 185.380 ;
        RECT 59.480 185.040 59.740 185.360 ;
        RECT 58.100 184.700 58.360 185.020 ;
        RECT 56.720 183.340 56.980 183.660 ;
        RECT 56.720 181.640 56.980 181.960 ;
        RECT 55.800 179.600 56.060 179.920 ;
        RECT 55.340 179.260 55.600 179.580 ;
        RECT 54.880 175.180 55.140 175.500 ;
        RECT 54.420 172.460 54.680 172.780 ;
        RECT 54.480 168.895 54.620 172.460 ;
        RECT 54.410 168.525 54.690 168.895 ;
        RECT 54.480 166.660 54.620 168.525 ;
        RECT 54.940 166.855 55.080 175.180 ;
        RECT 55.340 167.020 55.600 167.340 ;
        RECT 54.420 166.340 54.680 166.660 ;
        RECT 54.870 166.485 55.150 166.855 ;
        RECT 55.400 166.660 55.540 167.020 ;
        RECT 54.880 166.340 55.140 166.485 ;
        RECT 55.340 166.340 55.600 166.660 ;
        RECT 53.950 165.805 54.230 166.175 ;
        RECT 53.950 165.125 54.230 165.495 ;
        RECT 54.020 163.600 54.160 165.125 ;
        RECT 53.500 163.280 53.760 163.600 ;
        RECT 53.960 163.280 54.220 163.600 ;
        RECT 54.020 158.840 54.160 163.280 ;
        RECT 54.940 159.090 55.080 166.340 ;
        RECT 55.340 163.960 55.600 164.280 ;
        RECT 55.400 163.600 55.540 163.960 ;
        RECT 55.340 163.280 55.600 163.600 ;
        RECT 55.340 160.900 55.600 161.220 ;
        RECT 54.480 158.950 55.080 159.090 ;
        RECT 53.960 158.520 54.220 158.840 ;
        RECT 52.120 156.140 52.380 156.460 ;
        RECT 53.040 156.140 53.300 156.460 ;
        RECT 41.080 153.420 41.340 153.740 ;
        RECT 46.140 153.420 46.400 153.740 ;
        RECT 52.180 153.060 52.320 156.140 ;
        RECT 53.100 155.780 53.240 156.140 ;
        RECT 54.480 155.780 54.620 158.950 ;
        RECT 54.880 158.180 55.140 158.500 ;
        RECT 54.940 157.820 55.080 158.180 ;
        RECT 54.880 157.500 55.140 157.820 ;
        RECT 55.400 157.480 55.540 160.900 ;
        RECT 55.340 157.160 55.600 157.480 ;
        RECT 54.880 156.140 55.140 156.460 ;
        RECT 54.940 155.780 55.080 156.140 ;
        RECT 53.040 155.460 53.300 155.780 ;
        RECT 54.420 155.460 54.680 155.780 ;
        RECT 54.880 155.460 55.140 155.780 ;
        RECT 53.100 155.100 53.240 155.460 ;
        RECT 53.040 154.780 53.300 155.100 ;
        RECT 54.480 154.760 54.620 155.460 ;
        RECT 54.420 154.440 54.680 154.760 ;
        RECT 52.120 152.740 52.380 153.060 ;
        RECT 54.480 152.720 54.620 154.440 ;
        RECT 54.940 153.740 55.080 155.460 ;
        RECT 55.400 153.740 55.540 157.160 ;
        RECT 55.860 156.460 56.000 179.600 ;
        RECT 56.780 175.500 56.920 181.640 ;
        RECT 58.160 179.920 58.300 184.700 ;
        RECT 59.020 181.980 59.280 182.300 ;
        RECT 58.100 179.600 58.360 179.920 ;
        RECT 59.080 179.580 59.220 181.980 ;
        RECT 59.020 179.260 59.280 179.580 ;
        RECT 59.080 177.200 59.220 179.260 ;
        RECT 57.640 176.880 57.900 177.200 ;
        RECT 59.020 176.880 59.280 177.200 ;
        RECT 56.720 175.180 56.980 175.500 ;
        RECT 56.260 168.720 56.520 169.040 ;
        RECT 56.320 163.600 56.460 168.720 ;
        RECT 56.780 165.980 56.920 175.180 ;
        RECT 57.700 175.160 57.840 176.880 ;
        RECT 57.640 174.840 57.900 175.160 ;
        RECT 57.180 173.480 57.440 173.800 ;
        RECT 57.240 171.420 57.380 173.480 ;
        RECT 57.180 171.100 57.440 171.420 ;
        RECT 57.700 169.040 57.840 174.840 ;
        RECT 58.100 174.160 58.360 174.480 ;
        RECT 57.640 168.720 57.900 169.040 ;
        RECT 57.170 167.165 57.450 167.535 ;
        RECT 57.240 166.660 57.380 167.165 ;
        RECT 57.180 166.340 57.440 166.660 ;
        RECT 56.720 165.660 56.980 165.980 ;
        RECT 56.780 164.620 56.920 165.660 ;
        RECT 56.720 164.300 56.980 164.620 ;
        RECT 57.700 164.280 57.840 168.720 ;
        RECT 58.160 168.700 58.300 174.160 ;
        RECT 59.540 172.100 59.680 185.040 ;
        RECT 59.940 179.260 60.200 179.580 ;
        RECT 60.000 176.860 60.140 179.260 ;
        RECT 59.940 176.540 60.200 176.860 ;
        RECT 59.480 171.780 59.740 172.100 ;
        RECT 60.460 170.935 60.600 185.640 ;
        RECT 61.380 184.680 61.520 188.100 ;
        RECT 62.240 185.720 62.500 186.040 ;
        RECT 61.320 184.590 61.580 184.680 ;
        RECT 61.320 184.450 61.980 184.590 ;
        RECT 61.320 184.360 61.580 184.450 ;
        RECT 60.860 181.640 61.120 181.960 ;
        RECT 60.920 179.920 61.060 181.640 ;
        RECT 60.860 179.600 61.120 179.920 ;
        RECT 61.320 172.460 61.580 172.780 ;
        RECT 60.390 170.565 60.670 170.935 ;
        RECT 60.460 170.140 60.600 170.565 ;
        RECT 59.540 170.060 60.600 170.140 ;
        RECT 59.480 170.000 60.600 170.060 ;
        RECT 59.480 169.740 59.740 170.000 ;
        RECT 59.480 168.720 59.740 169.040 ;
        RECT 58.100 168.380 58.360 168.700 ;
        RECT 58.160 167.340 58.300 168.380 ;
        RECT 58.100 167.020 58.360 167.340 ;
        RECT 59.010 166.485 59.290 166.855 ;
        RECT 59.020 166.340 59.280 166.485 ;
        RECT 58.560 164.300 58.820 164.620 ;
        RECT 57.170 163.765 57.450 164.135 ;
        RECT 57.640 163.960 57.900 164.280 ;
        RECT 56.260 163.280 56.520 163.600 ;
        RECT 56.720 162.940 56.980 163.260 ;
        RECT 56.780 161.900 56.920 162.940 ;
        RECT 57.240 162.920 57.380 163.765 ;
        RECT 58.100 163.280 58.360 163.600 ;
        RECT 57.180 162.600 57.440 162.920 ;
        RECT 56.720 161.580 56.980 161.900 ;
        RECT 56.720 160.900 56.980 161.220 ;
        RECT 56.260 157.390 56.520 157.480 ;
        RECT 56.780 157.390 56.920 160.900 ;
        RECT 58.160 160.735 58.300 163.280 ;
        RECT 58.090 160.365 58.370 160.735 ;
        RECT 58.160 159.180 58.300 160.365 ;
        RECT 58.100 158.860 58.360 159.180 ;
        RECT 58.620 158.580 58.760 164.300 ;
        RECT 59.020 162.940 59.280 163.260 ;
        RECT 59.080 161.220 59.220 162.940 ;
        RECT 59.020 160.900 59.280 161.220 ;
        RECT 59.540 160.540 59.680 168.720 ;
        RECT 60.460 166.660 60.600 170.000 ;
        RECT 60.860 167.020 61.120 167.340 ;
        RECT 59.940 166.340 60.200 166.660 ;
        RECT 60.400 166.340 60.660 166.660 ;
        RECT 60.000 161.900 60.140 166.340 ;
        RECT 60.920 164.700 61.060 167.020 ;
        RECT 60.460 164.560 61.060 164.700 ;
        RECT 61.380 164.620 61.520 172.460 ;
        RECT 61.840 165.495 61.980 184.450 ;
        RECT 62.300 183.320 62.440 185.720 ;
        RECT 62.760 185.700 62.900 188.100 ;
        RECT 64.140 186.575 64.280 188.100 ;
        RECT 64.070 186.205 64.350 186.575 ;
        RECT 62.700 185.380 62.960 185.700 ;
        RECT 63.160 185.040 63.420 185.360 ;
        RECT 63.620 185.040 63.880 185.360 ;
        RECT 62.240 183.000 62.500 183.320 ;
        RECT 62.700 182.320 62.960 182.640 ;
        RECT 62.240 180.280 62.500 180.600 ;
        RECT 62.300 177.735 62.440 180.280 ;
        RECT 62.760 179.580 62.900 182.320 ;
        RECT 63.220 180.940 63.360 185.040 ;
        RECT 63.680 184.680 63.820 185.040 ;
        RECT 63.620 184.360 63.880 184.680 ;
        RECT 64.140 183.230 64.280 186.205 ;
        RECT 64.600 186.040 64.740 190.480 ;
        RECT 65.980 186.380 66.120 190.480 ;
        RECT 66.840 189.975 67.100 190.120 ;
        RECT 66.830 189.605 67.110 189.975 ;
        RECT 65.920 186.060 66.180 186.380 ;
        RECT 64.540 185.720 64.800 186.040 ;
        RECT 63.680 183.090 64.280 183.230 ;
        RECT 63.160 180.620 63.420 180.940 ;
        RECT 63.150 180.085 63.430 180.455 ;
        RECT 62.700 179.260 62.960 179.580 ;
        RECT 62.230 177.365 62.510 177.735 ;
        RECT 62.240 176.540 62.500 176.860 ;
        RECT 62.300 174.480 62.440 176.540 ;
        RECT 63.220 176.520 63.360 180.085 ;
        RECT 63.680 179.920 63.820 183.090 ;
        RECT 64.080 179.940 64.340 180.260 ;
        RECT 63.620 179.600 63.880 179.920 ;
        RECT 63.680 177.200 63.820 179.600 ;
        RECT 64.140 178.220 64.280 179.940 ;
        RECT 64.080 177.900 64.340 178.220 ;
        RECT 64.600 177.540 64.740 185.720 ;
        RECT 65.920 185.380 66.180 185.700 ;
        RECT 65.000 185.040 65.260 185.360 ;
        RECT 65.060 182.300 65.200 185.040 ;
        RECT 65.980 182.980 66.120 185.380 ;
        RECT 66.380 183.000 66.640 183.320 ;
        RECT 65.920 182.660 66.180 182.980 ;
        RECT 65.000 181.980 65.260 182.300 ;
        RECT 65.060 180.850 65.200 181.980 ;
        RECT 65.920 181.640 66.180 181.960 ;
        RECT 65.460 180.850 65.720 180.940 ;
        RECT 65.060 180.710 65.720 180.850 ;
        RECT 65.460 180.620 65.720 180.710 ;
        RECT 65.980 180.455 66.120 181.640 ;
        RECT 65.910 180.085 66.190 180.455 ;
        RECT 65.920 178.920 66.180 179.240 ;
        RECT 64.540 177.220 64.800 177.540 ;
        RECT 64.990 177.365 65.270 177.735 ;
        RECT 65.000 177.220 65.260 177.365 ;
        RECT 63.620 176.880 63.880 177.200 ;
        RECT 63.160 176.200 63.420 176.520 ;
        RECT 65.980 174.480 66.120 178.920 ;
        RECT 66.440 177.200 66.580 183.000 ;
        RECT 66.900 182.640 67.040 189.605 ;
        RECT 67.300 188.440 67.560 188.760 ;
        RECT 67.360 183.660 67.500 188.440 ;
        RECT 67.760 187.080 68.020 187.400 ;
        RECT 68.220 187.080 68.480 187.400 ;
        RECT 67.300 183.340 67.560 183.660 ;
        RECT 66.840 182.320 67.100 182.640 ;
        RECT 66.380 176.880 66.640 177.200 ;
        RECT 62.240 174.160 62.500 174.480 ;
        RECT 65.920 174.160 66.180 174.480 ;
        RECT 62.300 169.380 62.440 174.160 ;
        RECT 63.160 173.820 63.420 174.140 ;
        RECT 63.220 170.060 63.360 173.820 ;
        RECT 66.900 173.800 67.040 182.320 ;
        RECT 67.820 182.300 67.960 187.080 ;
        RECT 68.280 185.895 68.420 187.080 ;
        RECT 68.210 185.525 68.490 185.895 ;
        RECT 67.760 181.980 68.020 182.300 ;
        RECT 68.220 180.620 68.480 180.940 ;
        RECT 67.300 179.600 67.560 179.920 ;
        RECT 67.360 178.220 67.500 179.600 ;
        RECT 68.280 179.580 68.420 180.620 ;
        RECT 68.740 180.455 68.880 190.480 ;
        RECT 69.140 188.440 69.400 188.760 ;
        RECT 69.200 185.360 69.340 188.440 ;
        RECT 70.120 188.420 70.260 190.480 ;
        RECT 70.060 188.100 70.320 188.420 ;
        RECT 70.120 185.780 70.260 188.100 ;
        RECT 70.580 186.380 70.720 190.480 ;
        RECT 71.430 190.285 71.710 190.655 ;
        RECT 75.120 190.480 75.380 190.800 ;
        RECT 71.440 190.140 71.700 190.285 ;
        RECT 70.980 189.800 71.240 190.120 ;
        RECT 74.660 189.800 74.920 190.120 ;
        RECT 71.040 188.420 71.180 189.800 ;
        RECT 70.980 188.100 71.240 188.420 ;
        RECT 71.900 188.100 72.160 188.420 ;
        RECT 71.440 187.760 71.700 188.080 ;
        RECT 70.520 186.060 70.780 186.380 ;
        RECT 70.120 185.640 70.720 185.780 ;
        RECT 69.140 185.040 69.400 185.360 ;
        RECT 70.060 185.040 70.320 185.360 ;
        RECT 68.670 180.085 68.950 180.455 ;
        RECT 69.600 180.280 69.860 180.600 ;
        RECT 67.760 179.260 68.020 179.580 ;
        RECT 68.220 179.260 68.480 179.580 ;
        RECT 67.300 177.900 67.560 178.220 ;
        RECT 67.820 177.620 67.960 179.260 ;
        RECT 68.280 179.095 68.420 179.260 ;
        RECT 68.210 178.725 68.490 179.095 ;
        RECT 67.360 177.480 67.960 177.620 ;
        RECT 67.360 175.500 67.500 177.480 ;
        RECT 67.300 175.180 67.560 175.500 ;
        RECT 67.760 175.180 68.020 175.500 ;
        RECT 67.300 174.160 67.560 174.480 ;
        RECT 65.450 173.285 65.730 173.655 ;
        RECT 66.840 173.480 67.100 173.800 ;
        RECT 65.520 172.100 65.660 173.285 ;
        RECT 66.900 172.100 67.040 173.480 ;
        RECT 67.360 172.100 67.500 174.160 ;
        RECT 65.460 171.780 65.720 172.100 ;
        RECT 66.840 171.780 67.100 172.100 ;
        RECT 67.300 171.780 67.560 172.100 ;
        RECT 65.920 170.760 66.180 171.080 ;
        RECT 65.980 170.060 66.120 170.760 ;
        RECT 63.160 169.740 63.420 170.060 ;
        RECT 65.920 169.740 66.180 170.060 ;
        RECT 62.240 169.060 62.500 169.380 ;
        RECT 66.380 169.060 66.640 169.380 ;
        RECT 66.440 168.360 66.580 169.060 ;
        RECT 66.900 169.040 67.040 171.780 ;
        RECT 66.840 168.720 67.100 169.040 ;
        RECT 67.300 168.950 67.560 169.040 ;
        RECT 67.820 168.950 67.960 175.180 ;
        RECT 68.220 174.500 68.480 174.820 ;
        RECT 68.280 172.100 68.420 174.500 ;
        RECT 68.220 171.780 68.480 172.100 ;
        RECT 68.280 171.420 68.420 171.780 ;
        RECT 68.740 171.760 68.880 180.085 ;
        RECT 69.660 179.920 69.800 180.280 ;
        RECT 69.600 179.830 69.860 179.920 ;
        RECT 69.200 179.690 69.860 179.830 ;
        RECT 68.680 171.440 68.940 171.760 ;
        RECT 68.220 171.100 68.480 171.420 ;
        RECT 68.680 169.400 68.940 169.720 ;
        RECT 67.300 168.810 67.960 168.950 ;
        RECT 67.300 168.720 67.560 168.810 ;
        RECT 68.220 168.720 68.480 169.040 ;
        RECT 66.380 168.040 66.640 168.360 ;
        RECT 62.700 166.340 62.960 166.660 ;
        RECT 61.770 165.125 62.050 165.495 ;
        RECT 61.840 164.620 61.980 165.125 ;
        RECT 59.940 161.580 60.200 161.900 ;
        RECT 60.460 161.220 60.600 164.560 ;
        RECT 61.320 164.300 61.580 164.620 ;
        RECT 61.780 164.300 62.040 164.620 ;
        RECT 60.860 163.620 61.120 163.940 ;
        RECT 60.400 160.900 60.660 161.220 ;
        RECT 60.920 160.540 61.060 163.620 ;
        RECT 61.840 161.220 61.980 164.300 ;
        RECT 61.780 160.900 62.040 161.220 ;
        RECT 59.480 160.220 59.740 160.540 ;
        RECT 60.860 160.220 61.120 160.540 ;
        RECT 56.260 157.250 56.920 157.390 ;
        RECT 58.160 158.440 58.760 158.580 ;
        RECT 56.260 157.160 56.520 157.250 ;
        RECT 55.800 156.140 56.060 156.460 ;
        RECT 55.860 155.975 56.000 156.140 ;
        RECT 56.320 156.120 56.460 157.160 ;
        RECT 58.160 156.370 58.300 158.440 ;
        RECT 62.760 158.160 62.900 166.340 ;
        RECT 64.070 163.765 64.350 164.135 ;
        RECT 64.140 163.600 64.280 163.765 ;
        RECT 66.440 163.600 66.580 168.040 ;
        RECT 63.160 163.280 63.420 163.600 ;
        RECT 64.080 163.280 64.340 163.600 ;
        RECT 66.380 163.280 66.640 163.600 ;
        RECT 63.220 161.560 63.360 163.280 ;
        RECT 63.160 161.240 63.420 161.560 ;
        RECT 64.080 160.900 64.340 161.220 ;
        RECT 65.000 160.900 65.260 161.220 ;
        RECT 66.380 160.900 66.640 161.220 ;
        RECT 63.160 159.880 63.420 160.200 ;
        RECT 58.560 158.070 58.820 158.160 ;
        RECT 60.400 158.070 60.660 158.160 ;
        RECT 61.320 158.070 61.580 158.160 ;
        RECT 58.560 157.930 61.580 158.070 ;
        RECT 58.560 157.840 58.820 157.930 ;
        RECT 60.400 157.840 60.660 157.930 ;
        RECT 61.320 157.840 61.580 157.930 ;
        RECT 62.700 157.840 62.960 158.160 ;
        RECT 57.240 156.230 59.220 156.370 ;
        RECT 55.790 155.605 56.070 155.975 ;
        RECT 56.260 155.800 56.520 156.120 ;
        RECT 54.880 153.420 55.140 153.740 ;
        RECT 55.340 153.420 55.600 153.740 ;
        RECT 57.240 153.060 57.380 156.230 ;
        RECT 58.100 155.460 58.360 155.780 ;
        RECT 57.180 152.740 57.440 153.060 ;
        RECT 37.400 152.400 37.660 152.720 ;
        RECT 40.620 152.400 40.880 152.720 ;
        RECT 44.300 152.400 44.560 152.720 ;
        RECT 47.060 152.400 47.320 152.720 ;
        RECT 54.420 152.400 54.680 152.720 ;
        RECT 56.720 152.400 56.980 152.720 ;
        RECT 37.460 140.990 37.600 152.400 ;
        RECT 40.680 140.990 40.820 152.400 ;
        RECT 42.350 151.185 43.890 151.555 ;
        RECT 44.360 147.020 44.500 152.400 ;
        RECT 43.900 146.880 44.500 147.020 ;
        RECT 43.900 140.990 44.040 146.880 ;
        RECT 47.120 140.990 47.260 152.400 ;
        RECT 53.500 152.060 53.760 152.380 ;
        RECT 53.560 140.990 53.700 152.060 ;
        RECT 56.780 140.990 56.920 152.400 ;
        RECT 58.160 152.380 58.300 155.460 ;
        RECT 59.080 155.440 59.220 156.230 ;
        RECT 59.940 155.460 60.200 155.780 ;
        RECT 60.850 155.605 61.130 155.975 ;
        RECT 58.560 155.120 58.820 155.440 ;
        RECT 59.020 155.120 59.280 155.440 ;
        RECT 58.620 153.740 58.760 155.120 ;
        RECT 58.560 153.420 58.820 153.740 ;
        RECT 60.000 153.400 60.140 155.460 ;
        RECT 60.920 155.440 61.060 155.605 ;
        RECT 62.240 155.460 62.500 155.780 ;
        RECT 60.860 155.120 61.120 155.440 ;
        RECT 62.300 154.760 62.440 155.460 ;
        RECT 62.240 154.440 62.500 154.760 ;
        RECT 63.220 154.670 63.360 159.880 ;
        RECT 64.140 159.375 64.280 160.900 ;
        RECT 64.530 160.365 64.810 160.735 ;
        RECT 64.540 160.220 64.800 160.365 ;
        RECT 64.070 159.005 64.350 159.375 ;
        RECT 64.140 158.160 64.280 159.005 ;
        RECT 65.060 158.160 65.200 160.900 ;
        RECT 64.080 157.840 64.340 158.160 ;
        RECT 65.000 157.840 65.260 158.160 ;
        RECT 65.060 156.120 65.200 157.840 ;
        RECT 66.440 157.480 66.580 160.900 ;
        RECT 67.290 159.005 67.570 159.375 ;
        RECT 68.280 159.180 68.420 168.720 ;
        RECT 68.740 168.700 68.880 169.400 ;
        RECT 68.680 168.380 68.940 168.700 ;
        RECT 68.670 167.845 68.950 168.215 ;
        RECT 67.360 158.160 67.500 159.005 ;
        RECT 68.220 158.860 68.480 159.180 ;
        RECT 68.210 158.325 68.490 158.695 ;
        RECT 67.300 157.840 67.560 158.160 ;
        RECT 66.380 157.160 66.640 157.480 ;
        RECT 66.440 156.460 66.580 157.160 ;
        RECT 68.280 156.460 68.420 158.325 ;
        RECT 66.380 156.140 66.640 156.460 ;
        RECT 68.220 156.140 68.480 156.460 ;
        RECT 65.000 155.800 65.260 156.120 ;
        RECT 68.280 155.780 68.420 156.140 ;
        RECT 67.760 155.460 68.020 155.780 ;
        RECT 68.220 155.460 68.480 155.780 ;
        RECT 63.620 154.670 63.880 154.760 ;
        RECT 63.220 154.530 63.880 154.670 ;
        RECT 63.620 154.440 63.880 154.530 ;
        RECT 61.770 153.565 62.050 153.935 ;
        RECT 61.840 153.400 61.980 153.565 ;
        RECT 59.940 153.080 60.200 153.400 ;
        RECT 61.780 153.080 62.040 153.400 ;
        RECT 67.820 153.060 67.960 155.460 ;
        RECT 68.740 153.935 68.880 167.845 ;
        RECT 69.200 159.180 69.340 179.690 ;
        RECT 69.600 179.600 69.860 179.690 ;
        RECT 69.600 177.220 69.860 177.540 ;
        RECT 69.660 175.160 69.800 177.220 ;
        RECT 69.600 174.840 69.860 175.160 ;
        RECT 69.600 173.480 69.860 173.800 ;
        RECT 69.660 172.100 69.800 173.480 ;
        RECT 70.120 172.780 70.260 185.040 ;
        RECT 70.580 177.200 70.720 185.640 ;
        RECT 70.970 184.845 71.250 185.215 ;
        RECT 71.040 183.320 71.180 184.845 ;
        RECT 70.980 183.000 71.240 183.320 ;
        RECT 71.040 180.260 71.180 183.000 ;
        RECT 70.980 179.940 71.240 180.260 ;
        RECT 70.520 176.880 70.780 177.200 ;
        RECT 71.500 174.820 71.640 187.760 ;
        RECT 71.960 185.360 72.100 188.100 ;
        RECT 71.900 185.040 72.160 185.360 ;
        RECT 72.360 185.040 72.620 185.360 ;
        RECT 71.890 180.765 72.170 181.135 ;
        RECT 71.440 174.500 71.700 174.820 ;
        RECT 71.440 173.820 71.700 174.140 ;
        RECT 70.520 173.710 70.780 173.800 ;
        RECT 70.520 173.570 71.180 173.710 ;
        RECT 70.520 173.480 70.780 173.570 ;
        RECT 70.060 172.460 70.320 172.780 ;
        RECT 70.510 172.605 70.790 172.975 ;
        RECT 71.040 172.780 71.180 173.570 ;
        RECT 69.600 171.780 69.860 172.100 ;
        RECT 70.580 171.500 70.720 172.605 ;
        RECT 70.980 172.460 71.240 172.780 ;
        RECT 70.120 171.360 70.720 171.500 ;
        RECT 71.500 171.420 71.640 173.820 ;
        RECT 71.960 172.180 72.100 180.765 ;
        RECT 72.420 172.975 72.560 185.040 ;
        RECT 74.720 184.680 74.860 189.800 ;
        RECT 75.180 187.740 75.320 190.480 ;
        RECT 75.580 188.780 75.840 189.100 ;
        RECT 75.120 187.420 75.380 187.740 ;
        RECT 75.640 185.700 75.780 188.780 ;
        RECT 75.580 185.380 75.840 185.700 ;
        RECT 73.740 184.360 74.000 184.680 ;
        RECT 74.660 184.360 74.920 184.680 ;
        RECT 75.120 184.360 75.380 184.680 ;
        RECT 73.800 182.640 73.940 184.360 ;
        RECT 75.180 182.980 75.320 184.360 ;
        RECT 75.120 182.660 75.380 182.980 ;
        RECT 73.740 182.320 74.000 182.640 ;
        RECT 72.810 177.365 73.090 177.735 ;
        RECT 72.350 172.605 72.630 172.975 ;
        RECT 71.960 172.040 72.560 172.180 ;
        RECT 71.900 171.440 72.160 171.760 ;
        RECT 69.600 169.970 69.860 170.060 ;
        RECT 70.120 169.970 70.260 171.360 ;
        RECT 71.440 171.100 71.700 171.420 ;
        RECT 70.520 170.760 70.780 171.080 ;
        RECT 70.980 170.760 71.240 171.080 ;
        RECT 69.600 169.830 70.260 169.970 ;
        RECT 69.600 169.740 69.860 169.830 ;
        RECT 70.120 169.040 70.260 169.830 ;
        RECT 70.060 168.720 70.320 169.040 ;
        RECT 70.580 168.700 70.720 170.760 ;
        RECT 70.520 168.380 70.780 168.700 ;
        RECT 71.040 160.620 71.180 170.760 ;
        RECT 71.960 170.060 72.100 171.440 ;
        RECT 72.420 170.255 72.560 172.040 ;
        RECT 71.900 169.740 72.160 170.060 ;
        RECT 72.350 169.885 72.630 170.255 ;
        RECT 71.430 169.205 71.710 169.575 ;
        RECT 72.420 169.380 72.560 169.885 ;
        RECT 69.660 160.480 71.180 160.620 ;
        RECT 69.140 158.860 69.400 159.180 ;
        RECT 69.660 158.500 69.800 160.480 ;
        RECT 70.060 159.880 70.320 160.200 ;
        RECT 69.600 158.180 69.860 158.500 ;
        RECT 70.120 157.820 70.260 159.880 ;
        RECT 70.060 157.500 70.320 157.820 ;
        RECT 71.500 156.460 71.640 169.205 ;
        RECT 72.360 169.060 72.620 169.380 ;
        RECT 71.900 168.720 72.160 169.040 ;
        RECT 71.960 166.320 72.100 168.720 ;
        RECT 71.900 166.000 72.160 166.320 ;
        RECT 71.960 164.620 72.100 166.000 ;
        RECT 71.900 164.300 72.160 164.620 ;
        RECT 72.360 162.600 72.620 162.920 ;
        RECT 72.420 161.560 72.560 162.600 ;
        RECT 72.360 161.240 72.620 161.560 ;
        RECT 72.360 158.860 72.620 159.180 ;
        RECT 72.420 156.460 72.560 158.860 ;
        RECT 71.440 156.140 71.700 156.460 ;
        RECT 72.360 156.140 72.620 156.460 ;
        RECT 69.600 155.460 69.860 155.780 ;
        RECT 71.900 155.460 72.160 155.780 ;
        RECT 72.360 155.460 72.620 155.780 ;
        RECT 69.660 154.615 69.800 155.460 ;
        RECT 70.980 155.120 71.240 155.440 ;
        RECT 71.960 155.295 72.100 155.460 ;
        RECT 71.040 154.670 71.180 155.120 ;
        RECT 71.890 154.925 72.170 155.295 ;
        RECT 71.900 154.670 72.160 154.760 ;
        RECT 69.590 154.245 69.870 154.615 ;
        RECT 71.040 154.530 72.160 154.670 ;
        RECT 71.900 154.440 72.160 154.530 ;
        RECT 68.670 153.565 68.950 153.935 ;
        RECT 67.760 152.740 68.020 153.060 ;
        RECT 65.460 152.400 65.720 152.720 ;
        RECT 68.220 152.400 68.480 152.720 ;
        RECT 58.100 152.060 58.360 152.380 ;
        RECT 58.160 148.980 58.300 152.060 ;
        RECT 60.400 151.720 60.660 152.040 ;
        RECT 60.460 149.855 60.600 151.720 ;
        RECT 60.390 149.485 60.670 149.855 ;
        RECT 65.520 149.660 65.660 152.400 ;
        RECT 66.380 151.720 66.640 152.040 ;
        RECT 67.760 151.720 68.020 152.040 ;
        RECT 65.460 149.340 65.720 149.660 ;
        RECT 58.100 148.660 58.360 148.980 ;
        RECT 66.440 141.015 66.580 151.720 ;
        RECT 67.820 143.880 67.960 151.720 ;
        RECT 68.280 150.000 68.420 152.400 ;
        RECT 70.520 152.060 70.780 152.380 ;
        RECT 69.140 151.720 69.400 152.040 ;
        RECT 68.220 149.680 68.480 150.000 ;
        RECT 69.200 146.260 69.340 151.720 ;
        RECT 69.140 145.940 69.400 146.260 ;
        RECT 67.760 143.560 68.020 143.880 ;
        RECT 70.580 141.160 70.720 152.060 ;
        RECT 72.420 150.340 72.560 155.460 ;
        RECT 72.880 155.440 73.020 177.365 ;
        RECT 73.270 173.285 73.550 173.655 ;
        RECT 73.340 171.760 73.480 173.285 ;
        RECT 73.280 171.440 73.540 171.760 ;
        RECT 73.280 168.270 73.540 168.360 ;
        RECT 73.800 168.270 73.940 182.320 ;
        RECT 75.640 174.480 75.780 185.380 ;
        RECT 76.100 185.100 76.240 190.820 ;
        RECT 78.340 190.480 78.600 190.800 ;
        RECT 78.800 190.480 79.060 190.800 ;
        RECT 76.500 189.800 76.760 190.120 ;
        RECT 76.560 186.380 76.700 189.800 ;
        RECT 78.400 187.935 78.540 190.480 ;
        RECT 78.860 189.100 79.000 190.480 ;
        RECT 81.160 190.460 81.300 191.500 ;
        RECT 81.100 190.140 81.360 190.460 ;
        RECT 78.800 188.780 79.060 189.100 ;
        RECT 80.180 188.780 80.440 189.100 ;
        RECT 79.720 188.440 79.980 188.760 ;
        RECT 78.330 187.565 78.610 187.935 ;
        RECT 79.260 187.760 79.520 188.080 ;
        RECT 76.960 187.080 77.220 187.400 ;
        RECT 76.500 186.060 76.760 186.380 ;
        RECT 77.020 185.700 77.160 187.080 ;
        RECT 76.960 185.380 77.220 185.700 ;
        RECT 79.320 185.360 79.460 187.760 ;
        RECT 76.100 184.960 77.160 185.100 ;
        RECT 77.420 185.040 77.680 185.360 ;
        RECT 78.340 185.215 78.600 185.360 ;
        RECT 76.500 179.940 76.760 180.260 ;
        RECT 76.560 177.540 76.700 179.940 ;
        RECT 76.500 177.220 76.760 177.540 ;
        RECT 76.560 175.695 76.700 177.220 ;
        RECT 76.490 175.325 76.770 175.695 ;
        RECT 76.040 174.500 76.300 174.820 ;
        RECT 74.200 174.160 74.460 174.480 ;
        RECT 75.580 174.160 75.840 174.480 ;
        RECT 74.260 168.700 74.400 174.160 ;
        RECT 74.660 173.820 74.920 174.140 ;
        RECT 74.720 172.975 74.860 173.820 ;
        RECT 74.650 172.605 74.930 172.975 ;
        RECT 75.110 171.925 75.390 172.295 ;
        RECT 74.660 171.440 74.920 171.760 ;
        RECT 74.720 168.700 74.860 171.440 ;
        RECT 74.200 168.380 74.460 168.700 ;
        RECT 74.660 168.380 74.920 168.700 ;
        RECT 73.280 168.130 73.940 168.270 ;
        RECT 73.280 168.040 73.540 168.130 ;
        RECT 73.340 166.320 73.480 168.040 ;
        RECT 74.260 167.535 74.400 168.380 ;
        RECT 73.740 167.020 74.000 167.340 ;
        RECT 74.190 167.165 74.470 167.535 ;
        RECT 73.800 166.855 73.940 167.020 ;
        RECT 73.730 166.485 74.010 166.855 ;
        RECT 74.660 166.680 74.920 167.000 ;
        RECT 73.280 166.000 73.540 166.320 ;
        RECT 73.280 163.620 73.540 163.940 ;
        RECT 73.340 158.160 73.480 163.620 ;
        RECT 73.800 163.600 73.940 166.485 ;
        RECT 74.200 163.960 74.460 164.280 ;
        RECT 73.740 163.280 74.000 163.600 ;
        RECT 73.740 162.600 74.000 162.920 ;
        RECT 73.800 159.180 73.940 162.600 ;
        RECT 73.740 158.860 74.000 159.180 ;
        RECT 74.260 158.160 74.400 163.960 ;
        RECT 74.720 163.260 74.860 166.680 ;
        RECT 75.180 166.660 75.320 171.925 ;
        RECT 76.100 169.720 76.240 174.500 ;
        RECT 77.020 172.100 77.160 184.960 ;
        RECT 77.480 184.680 77.620 185.040 ;
        RECT 78.330 184.845 78.610 185.215 ;
        RECT 79.260 185.040 79.520 185.360 ;
        RECT 77.420 184.360 77.680 184.680 ;
        RECT 78.340 184.360 78.600 184.680 ;
        RECT 77.420 181.640 77.680 181.960 ;
        RECT 77.880 181.640 78.140 181.960 ;
        RECT 77.480 179.920 77.620 181.640 ;
        RECT 77.940 179.920 78.080 181.640 ;
        RECT 78.400 180.940 78.540 184.360 ;
        RECT 79.320 183.320 79.460 185.040 ;
        RECT 79.780 184.680 79.920 188.440 ;
        RECT 79.720 184.360 79.980 184.680 ;
        RECT 79.260 183.000 79.520 183.320 ;
        RECT 78.800 182.320 79.060 182.640 ;
        RECT 78.340 180.620 78.600 180.940 ;
        RECT 77.420 179.600 77.680 179.920 ;
        RECT 77.880 179.600 78.140 179.920 ;
        RECT 76.500 171.780 76.760 172.100 ;
        RECT 76.960 171.780 77.220 172.100 ;
        RECT 76.040 169.400 76.300 169.720 ;
        RECT 76.040 166.680 76.300 167.000 ;
        RECT 75.120 166.340 75.380 166.660 ;
        RECT 75.580 166.340 75.840 166.660 ;
        RECT 75.640 164.620 75.780 166.340 ;
        RECT 75.580 164.300 75.840 164.620 ;
        RECT 75.120 163.620 75.380 163.940 ;
        RECT 74.660 162.940 74.920 163.260 ;
        RECT 74.720 161.560 74.860 162.940 ;
        RECT 75.180 161.980 75.320 163.620 ;
        RECT 75.640 163.600 75.780 164.300 ;
        RECT 75.580 163.280 75.840 163.600 ;
        RECT 75.180 161.840 75.780 161.980 ;
        RECT 75.640 161.560 75.780 161.840 ;
        RECT 74.660 161.240 74.920 161.560 ;
        RECT 75.580 161.240 75.840 161.560 ;
        RECT 74.660 160.560 74.920 160.880 ;
        RECT 74.720 160.200 74.860 160.560 ;
        RECT 75.580 160.220 75.840 160.540 ;
        RECT 74.660 159.880 74.920 160.200 ;
        RECT 75.120 159.880 75.380 160.200 ;
        RECT 75.180 159.180 75.320 159.880 ;
        RECT 75.120 158.860 75.380 159.180 ;
        RECT 73.280 157.840 73.540 158.160 ;
        RECT 73.740 157.840 74.000 158.160 ;
        RECT 74.200 157.840 74.460 158.160 ;
        RECT 73.340 155.780 73.480 157.840 ;
        RECT 73.800 157.480 73.940 157.840 ;
        RECT 73.740 157.160 74.000 157.480 ;
        RECT 73.280 155.460 73.540 155.780 ;
        RECT 72.820 155.120 73.080 155.440 ;
        RECT 73.800 155.180 73.940 157.160 ;
        RECT 74.260 156.120 74.400 157.840 ;
        RECT 75.640 157.820 75.780 160.220 ;
        RECT 76.100 159.180 76.240 166.680 ;
        RECT 76.560 161.415 76.700 171.780 ;
        RECT 77.020 168.360 77.160 171.780 ;
        RECT 77.480 171.080 77.620 179.600 ;
        RECT 78.340 178.920 78.600 179.240 ;
        RECT 77.880 174.390 78.140 174.480 ;
        RECT 78.400 174.390 78.540 178.920 ;
        RECT 78.860 177.880 79.000 182.320 ;
        RECT 80.240 178.980 80.380 188.780 ;
        RECT 80.640 187.760 80.900 188.080 ;
        RECT 80.700 183.660 80.840 187.760 ;
        RECT 80.640 183.340 80.900 183.660 ;
        RECT 80.640 182.660 80.900 182.980 ;
        RECT 80.700 180.600 80.840 182.660 ;
        RECT 80.640 180.280 80.900 180.600 ;
        RECT 80.700 179.580 80.840 180.280 ;
        RECT 81.160 179.920 81.300 190.140 ;
        RECT 81.620 189.295 81.760 192.520 ;
        RECT 82.480 191.160 82.740 191.480 ;
        RECT 82.020 190.140 82.280 190.460 ;
        RECT 81.550 188.925 81.830 189.295 ;
        RECT 82.080 189.100 82.220 190.140 ;
        RECT 82.540 189.100 82.680 191.160 ;
        RECT 83.460 190.800 83.600 193.200 ;
        RECT 87.600 191.820 87.740 193.540 ;
        RECT 87.540 191.500 87.800 191.820 ;
        RECT 91.280 191.480 91.420 193.540 ;
        RECT 91.220 191.160 91.480 191.480 ;
        RECT 83.400 190.480 83.660 190.800 ;
        RECT 86.620 190.480 86.880 190.800 ;
        RECT 88.920 190.480 89.180 190.800 ;
        RECT 92.140 190.710 92.400 190.800 ;
        RECT 93.060 190.710 93.320 190.800 ;
        RECT 92.140 190.570 93.320 190.710 ;
        RECT 92.140 190.480 92.400 190.570 ;
        RECT 93.060 190.480 93.320 190.570 ;
        RECT 83.460 189.100 83.600 190.480 ;
        RECT 82.020 188.780 82.280 189.100 ;
        RECT 82.480 188.780 82.740 189.100 ;
        RECT 83.400 188.780 83.660 189.100 ;
        RECT 82.020 188.100 82.280 188.420 ;
        RECT 82.080 186.040 82.220 188.100 ;
        RECT 82.480 187.420 82.740 187.740 ;
        RECT 82.020 185.720 82.280 186.040 ;
        RECT 82.080 184.680 82.220 185.720 ;
        RECT 82.020 184.360 82.280 184.680 ;
        RECT 82.540 181.135 82.680 187.420 ;
        RECT 86.680 187.255 86.820 190.480 ;
        RECT 88.980 189.975 89.120 190.480 ;
        RECT 88.910 189.605 89.190 189.975 ;
        RECT 89.380 189.800 89.640 190.120 ;
        RECT 90.760 189.800 91.020 190.120 ;
        RECT 88.460 188.100 88.720 188.420 ;
        RECT 87.990 187.565 88.270 187.935 ;
        RECT 88.000 187.420 88.260 187.565 ;
        RECT 86.610 186.885 86.890 187.255 ;
        RECT 87.080 187.080 87.340 187.400 ;
        RECT 85.700 186.060 85.960 186.380 ;
        RECT 82.940 184.700 83.200 185.020 ;
        RECT 84.320 184.700 84.580 185.020 ;
        RECT 82.470 180.765 82.750 181.135 ;
        RECT 81.100 179.830 81.360 179.920 ;
        RECT 82.020 179.830 82.280 179.920 ;
        RECT 81.100 179.690 82.280 179.830 ;
        RECT 81.100 179.600 81.360 179.690 ;
        RECT 82.020 179.600 82.280 179.690 ;
        RECT 80.640 179.260 80.900 179.580 ;
        RECT 80.240 178.840 81.300 178.980 ;
        RECT 82.020 178.920 82.280 179.240 ;
        RECT 78.800 177.560 79.060 177.880 ;
        RECT 80.640 177.220 80.900 177.540 ;
        RECT 78.800 176.880 79.060 177.200 ;
        RECT 78.860 174.820 79.000 176.880 ;
        RECT 80.700 176.375 80.840 177.220 ;
        RECT 80.630 176.005 80.910 176.375 ;
        RECT 78.800 174.500 79.060 174.820 ;
        RECT 79.260 174.500 79.520 174.820 ;
        RECT 77.880 174.250 78.540 174.390 ;
        RECT 77.880 174.160 78.140 174.250 ;
        RECT 79.320 174.220 79.460 174.500 ;
        RECT 78.860 174.080 79.460 174.220 ;
        RECT 79.720 174.160 79.980 174.480 ;
        RECT 80.180 174.160 80.440 174.480 ;
        RECT 77.880 171.780 78.140 172.100 ;
        RECT 77.420 170.760 77.680 171.080 ;
        RECT 76.960 168.040 77.220 168.360 ;
        RECT 77.480 166.570 77.620 170.760 ;
        RECT 77.940 170.060 78.080 171.780 ;
        RECT 77.880 169.740 78.140 170.060 ;
        RECT 78.860 169.380 79.000 174.080 ;
        RECT 79.260 173.480 79.520 173.800 ;
        RECT 79.320 172.100 79.460 173.480 ;
        RECT 79.260 171.780 79.520 172.100 ;
        RECT 78.800 169.060 79.060 169.380 ;
        RECT 78.790 168.525 79.070 168.895 ;
        RECT 78.860 166.660 79.000 168.525 ;
        RECT 77.880 166.570 78.140 166.660 ;
        RECT 77.480 166.430 78.140 166.570 ;
        RECT 76.960 166.000 77.220 166.320 ;
        RECT 76.490 161.045 76.770 161.415 ;
        RECT 76.040 158.860 76.300 159.180 ;
        RECT 76.100 158.500 76.240 158.860 ;
        RECT 76.040 158.180 76.300 158.500 ;
        RECT 76.500 158.180 76.760 158.500 ;
        RECT 75.580 157.500 75.840 157.820 ;
        RECT 76.100 157.480 76.240 158.180 ;
        RECT 76.040 157.160 76.300 157.480 ;
        RECT 74.200 155.800 74.460 156.120 ;
        RECT 76.560 155.780 76.700 158.180 ;
        RECT 76.500 155.460 76.760 155.780 ;
        RECT 73.800 155.040 74.860 155.180 ;
        RECT 74.720 154.760 74.860 155.040 ;
        RECT 72.820 154.670 73.080 154.760 ;
        RECT 72.820 154.530 73.480 154.670 ;
        RECT 72.820 154.440 73.080 154.530 ;
        RECT 72.820 153.420 73.080 153.740 ;
        RECT 72.880 152.720 73.020 153.420 ;
        RECT 73.340 153.255 73.480 154.530 ;
        RECT 74.200 154.440 74.460 154.760 ;
        RECT 74.660 154.440 74.920 154.760 ;
        RECT 73.270 152.885 73.550 153.255 ;
        RECT 72.820 152.400 73.080 152.720 ;
        RECT 73.740 152.400 74.000 152.720 ;
        RECT 73.280 151.720 73.540 152.040 ;
        RECT 72.360 150.020 72.620 150.340 ;
        RECT 73.340 146.940 73.480 151.720 ;
        RECT 73.800 151.020 73.940 152.400 ;
        RECT 73.740 150.700 74.000 151.020 ;
        RECT 74.260 147.280 74.400 154.440 ;
        RECT 77.020 153.400 77.160 166.000 ;
        RECT 77.480 162.920 77.620 166.430 ;
        RECT 77.880 166.340 78.140 166.430 ;
        RECT 78.800 166.340 79.060 166.660 ;
        RECT 79.260 165.660 79.520 165.980 ;
        RECT 79.320 164.135 79.460 165.660 ;
        RECT 79.250 163.765 79.530 164.135 ;
        RECT 78.340 162.940 78.600 163.260 ;
        RECT 77.420 162.600 77.680 162.920 ;
        RECT 78.400 161.900 78.540 162.940 ;
        RECT 78.800 162.600 79.060 162.920 ;
        RECT 78.340 161.580 78.600 161.900 ;
        RECT 78.860 160.735 79.000 162.600 ;
        RECT 79.250 162.405 79.530 162.775 ;
        RECT 79.320 160.880 79.460 162.405 ;
        RECT 79.780 161.130 79.920 174.160 ;
        RECT 80.240 171.420 80.380 174.160 ;
        RECT 80.700 172.100 80.840 176.005 ;
        RECT 81.160 174.480 81.300 178.840 ;
        RECT 81.550 174.645 81.830 175.015 ;
        RECT 81.100 174.160 81.360 174.480 ;
        RECT 81.090 173.285 81.370 173.655 ;
        RECT 80.640 171.780 80.900 172.100 ;
        RECT 80.180 171.100 80.440 171.420 ;
        RECT 80.180 168.610 80.440 168.700 ;
        RECT 81.160 168.610 81.300 173.285 ;
        RECT 81.620 172.440 81.760 174.645 ;
        RECT 82.080 174.480 82.220 178.920 ;
        RECT 83.000 177.880 83.140 184.700 ;
        RECT 83.400 184.360 83.660 184.680 ;
        RECT 83.860 184.360 84.120 184.680 ;
        RECT 83.460 180.600 83.600 184.360 ;
        RECT 83.920 180.940 84.060 184.360 ;
        RECT 84.380 182.980 84.520 184.700 ;
        RECT 84.320 182.660 84.580 182.980 ;
        RECT 83.860 180.620 84.120 180.940 ;
        RECT 83.400 180.280 83.660 180.600 ;
        RECT 82.940 177.560 83.200 177.880 ;
        RECT 82.480 177.055 82.740 177.200 ;
        RECT 82.470 176.685 82.750 177.055 ;
        RECT 82.020 174.160 82.280 174.480 ;
        RECT 82.480 174.390 82.740 174.480 ;
        RECT 83.000 174.390 83.140 177.560 ;
        RECT 82.480 174.250 83.140 174.390 ;
        RECT 82.480 174.160 82.740 174.250 ;
        RECT 82.010 172.605 82.290 172.975 ;
        RECT 82.540 172.780 82.680 174.160 ;
        RECT 83.850 173.965 84.130 174.335 ;
        RECT 81.560 172.120 81.820 172.440 ;
        RECT 82.080 171.420 82.220 172.605 ;
        RECT 82.480 172.460 82.740 172.780 ;
        RECT 83.390 172.605 83.670 172.975 ;
        RECT 82.020 171.100 82.280 171.420 ;
        RECT 82.020 168.720 82.280 169.040 ;
        RECT 80.180 168.470 81.300 168.610 ;
        RECT 80.180 168.380 80.440 168.470 ;
        RECT 80.180 166.680 80.440 167.000 ;
        RECT 80.240 164.815 80.380 166.680 ;
        RECT 80.170 164.445 80.450 164.815 ;
        RECT 82.080 164.620 82.220 168.720 ;
        RECT 82.940 168.610 83.200 168.700 ;
        RECT 83.460 168.610 83.600 172.605 ;
        RECT 83.920 169.040 84.060 173.965 ;
        RECT 84.380 171.500 84.520 182.660 ;
        RECT 84.780 181.640 85.040 181.960 ;
        RECT 84.840 179.920 84.980 181.640 ;
        RECT 85.760 179.920 85.900 186.060 ;
        RECT 87.140 185.700 87.280 187.080 ;
        RECT 87.080 185.380 87.340 185.700 ;
        RECT 86.160 184.360 86.420 184.680 ;
        RECT 86.220 183.660 86.360 184.360 ;
        RECT 88.520 183.660 88.660 188.100 ;
        RECT 86.160 183.340 86.420 183.660 ;
        RECT 88.460 183.340 88.720 183.660 ;
        RECT 88.910 182.805 89.190 183.175 ;
        RECT 87.080 181.640 87.340 181.960 ;
        RECT 84.780 179.600 85.040 179.920 ;
        RECT 85.700 179.600 85.960 179.920 ;
        RECT 84.780 175.180 85.040 175.500 ;
        RECT 84.840 174.335 84.980 175.180 ;
        RECT 84.770 173.965 85.050 174.335 ;
        RECT 85.240 173.820 85.500 174.140 ;
        RECT 84.780 173.655 85.040 173.800 ;
        RECT 84.770 173.285 85.050 173.655 ;
        RECT 84.380 171.360 84.980 171.500 ;
        RECT 84.320 170.760 84.580 171.080 ;
        RECT 84.380 169.380 84.520 170.760 ;
        RECT 84.320 169.060 84.580 169.380 ;
        RECT 83.860 168.720 84.120 169.040 ;
        RECT 84.840 168.780 84.980 171.360 ;
        RECT 85.300 170.060 85.440 173.820 ;
        RECT 85.240 169.740 85.500 170.060 ;
        RECT 85.760 169.290 85.900 179.600 ;
        RECT 86.160 174.160 86.420 174.480 ;
        RECT 86.620 174.160 86.880 174.480 ;
        RECT 86.220 172.780 86.360 174.160 ;
        RECT 86.680 173.800 86.820 174.160 ;
        RECT 86.620 173.480 86.880 173.800 ;
        RECT 86.160 172.460 86.420 172.780 ;
        RECT 86.160 171.440 86.420 171.760 ;
        RECT 86.680 171.615 86.820 173.480 ;
        RECT 86.220 169.720 86.360 171.440 ;
        RECT 86.610 171.245 86.890 171.615 ;
        RECT 86.610 169.885 86.890 170.255 ;
        RECT 86.620 169.740 86.880 169.885 ;
        RECT 86.160 169.400 86.420 169.720 ;
        RECT 82.940 168.470 83.600 168.610 ;
        RECT 84.380 168.640 84.980 168.780 ;
        RECT 85.300 169.150 85.900 169.290 ;
        RECT 82.940 168.380 83.200 168.470 ;
        RECT 83.000 168.215 83.140 168.380 ;
        RECT 82.930 167.845 83.210 168.215 ;
        RECT 83.400 165.320 83.660 165.640 ;
        RECT 83.860 165.320 84.120 165.640 ;
        RECT 81.560 164.300 81.820 164.620 ;
        RECT 82.020 164.300 82.280 164.620 ;
        RECT 80.170 163.765 80.450 164.135 ;
        RECT 80.240 163.600 80.380 163.765 ;
        RECT 80.180 163.280 80.440 163.600 ;
        RECT 80.240 162.095 80.380 163.280 ;
        RECT 81.100 162.940 81.360 163.260 ;
        RECT 80.170 161.725 80.450 162.095 ;
        RECT 79.780 160.990 80.380 161.130 ;
        RECT 80.630 161.045 80.910 161.415 ;
        RECT 77.420 160.220 77.680 160.540 ;
        RECT 78.790 160.365 79.070 160.735 ;
        RECT 79.260 160.560 79.520 160.880 ;
        RECT 77.480 160.055 77.620 160.220 ;
        RECT 77.410 159.685 77.690 160.055 ;
        RECT 77.880 159.880 78.140 160.200 ;
        RECT 79.260 159.880 79.520 160.200 ;
        RECT 77.420 157.840 77.680 158.160 ;
        RECT 77.480 155.440 77.620 157.840 ;
        RECT 77.940 155.860 78.080 159.880 ;
        RECT 79.320 158.160 79.460 159.880 ;
        RECT 79.710 159.685 79.990 160.055 ;
        RECT 79.780 158.160 79.920 159.685 ;
        RECT 79.260 157.840 79.520 158.160 ;
        RECT 79.720 157.840 79.980 158.160 ;
        RECT 78.800 157.500 79.060 157.820 ;
        RECT 78.860 156.460 79.000 157.500 ;
        RECT 79.320 156.460 79.460 157.840 ;
        RECT 79.720 157.160 79.980 157.480 ;
        RECT 78.800 156.140 79.060 156.460 ;
        RECT 79.260 156.140 79.520 156.460 ;
        RECT 77.940 155.720 79.000 155.860 ;
        RECT 77.420 155.350 77.680 155.440 ;
        RECT 78.340 155.350 78.600 155.440 ;
        RECT 77.420 155.210 78.600 155.350 ;
        RECT 77.420 155.120 77.680 155.210 ;
        RECT 78.340 155.120 78.600 155.210 ;
        RECT 78.860 154.760 79.000 155.720 ;
        RECT 79.250 155.605 79.530 155.975 ;
        RECT 79.260 155.460 79.520 155.605 ;
        RECT 78.800 154.440 79.060 154.760 ;
        RECT 76.960 153.080 77.220 153.400 ;
        RECT 78.860 152.720 79.000 154.440 ;
        RECT 79.780 152.720 79.920 157.160 ;
        RECT 80.240 155.780 80.380 160.990 ;
        RECT 80.700 160.200 80.840 161.045 ;
        RECT 81.160 160.540 81.300 162.940 ;
        RECT 81.100 160.220 81.360 160.540 ;
        RECT 80.640 159.880 80.900 160.200 ;
        RECT 81.160 159.180 81.300 160.220 ;
        RECT 81.100 158.860 81.360 159.180 ;
        RECT 80.640 157.840 80.900 158.160 ;
        RECT 80.180 155.460 80.440 155.780 ;
        RECT 80.700 154.760 80.840 157.840 ;
        RECT 81.620 157.480 81.760 164.300 ;
        RECT 82.020 163.280 82.280 163.600 ;
        RECT 81.560 157.160 81.820 157.480 ;
        RECT 81.100 156.370 81.360 156.460 ;
        RECT 81.620 156.370 81.760 157.160 ;
        RECT 82.080 156.460 82.220 163.280 ;
        RECT 82.940 162.600 83.200 162.920 ;
        RECT 82.470 161.725 82.750 162.095 ;
        RECT 82.540 158.070 82.680 161.725 ;
        RECT 83.000 160.540 83.140 162.600 ;
        RECT 82.940 160.220 83.200 160.540 ;
        RECT 83.460 159.180 83.600 165.320 ;
        RECT 83.920 164.135 84.060 165.320 ;
        RECT 83.850 163.765 84.130 164.135 ;
        RECT 84.380 163.600 84.520 168.640 ;
        RECT 84.780 168.040 85.040 168.360 ;
        RECT 84.840 166.660 84.980 168.040 ;
        RECT 85.300 167.340 85.440 169.150 ;
        RECT 85.700 168.380 85.960 168.700 ;
        RECT 85.240 167.020 85.500 167.340 ;
        RECT 84.780 166.340 85.040 166.660 ;
        RECT 83.860 163.280 84.120 163.600 ;
        RECT 84.320 163.455 84.580 163.600 ;
        RECT 83.920 162.775 84.060 163.280 ;
        RECT 84.310 163.085 84.590 163.455 ;
        RECT 83.850 162.405 84.130 162.775 ;
        RECT 84.320 162.600 84.580 162.920 ;
        RECT 84.380 161.900 84.520 162.600 ;
        RECT 84.320 161.580 84.580 161.900 ;
        RECT 84.840 161.415 84.980 166.340 ;
        RECT 84.770 161.045 85.050 161.415 ;
        RECT 85.300 161.220 85.440 167.020 ;
        RECT 85.760 165.640 85.900 168.380 ;
        RECT 86.610 167.845 86.890 168.215 ;
        RECT 85.700 165.320 85.960 165.640 ;
        RECT 85.760 162.775 85.900 165.320 ;
        RECT 86.160 163.960 86.420 164.280 ;
        RECT 85.690 162.405 85.970 162.775 ;
        RECT 86.220 161.220 86.360 163.960 ;
        RECT 86.680 163.600 86.820 167.845 ;
        RECT 87.140 165.640 87.280 181.640 ;
        RECT 88.460 176.540 88.720 176.860 ;
        RECT 88.520 174.480 88.660 176.540 ;
        RECT 88.460 174.390 88.720 174.480 ;
        RECT 88.060 174.250 88.720 174.390 ;
        RECT 87.540 173.480 87.800 173.800 ;
        RECT 87.600 170.255 87.740 173.480 ;
        RECT 87.530 169.885 87.810 170.255 ;
        RECT 87.530 169.205 87.810 169.575 ;
        RECT 87.600 168.700 87.740 169.205 ;
        RECT 88.060 169.040 88.200 174.250 ;
        RECT 88.460 174.160 88.720 174.250 ;
        RECT 88.460 171.440 88.720 171.760 ;
        RECT 88.000 168.720 88.260 169.040 ;
        RECT 87.540 168.380 87.800 168.700 ;
        RECT 88.520 167.535 88.660 171.440 ;
        RECT 88.450 167.165 88.730 167.535 ;
        RECT 88.460 166.680 88.720 167.000 ;
        RECT 88.000 166.340 88.260 166.660 ;
        RECT 87.540 165.660 87.800 165.980 ;
        RECT 87.080 165.320 87.340 165.640 ;
        RECT 86.620 163.280 86.880 163.600 ;
        RECT 87.140 161.220 87.280 165.320 ;
        RECT 87.600 163.600 87.740 165.660 ;
        RECT 88.060 165.640 88.200 166.340 ;
        RECT 88.000 165.320 88.260 165.640 ;
        RECT 88.060 164.815 88.200 165.320 ;
        RECT 87.990 164.445 88.270 164.815 ;
        RECT 88.520 164.530 88.660 166.680 ;
        RECT 88.980 165.980 89.120 182.805 ;
        RECT 89.440 179.920 89.580 189.800 ;
        RECT 90.300 188.100 90.560 188.420 ;
        RECT 90.360 183.660 90.500 188.100 ;
        RECT 90.820 185.360 90.960 189.800 ;
        RECT 94.040 188.860 94.180 193.880 ;
        RECT 97.190 193.685 97.470 194.055 ;
        RECT 95.360 192.750 95.620 192.840 ;
        RECT 94.960 192.610 95.620 192.750 ;
        RECT 94.960 191.140 95.100 192.610 ;
        RECT 95.360 192.520 95.620 192.610 ;
        RECT 94.900 190.820 95.160 191.140 ;
        RECT 95.820 189.800 96.080 190.120 ;
        RECT 96.740 190.030 97.000 190.120 ;
        RECT 96.340 189.890 97.000 190.030 ;
        RECT 93.520 188.500 93.780 188.760 ;
        RECT 94.040 188.720 95.100 188.860 ;
        RECT 93.520 188.440 94.180 188.500 ;
        RECT 93.580 188.360 94.180 188.440 ;
        RECT 93.050 186.205 93.330 186.575 ;
        RECT 93.060 186.060 93.320 186.205 ;
        RECT 93.520 186.060 93.780 186.380 ;
        RECT 90.760 185.040 91.020 185.360 ;
        RECT 92.600 185.270 92.860 185.360 ;
        RECT 92.200 185.130 92.860 185.270 ;
        RECT 90.300 183.340 90.560 183.660 ;
        RECT 89.840 182.660 90.100 182.980 ;
        RECT 89.900 180.600 90.040 182.660 ;
        RECT 89.840 180.280 90.100 180.600 ;
        RECT 90.360 180.455 90.500 183.340 ;
        RECT 90.820 182.640 90.960 185.040 ;
        RECT 91.220 184.360 91.480 184.680 ;
        RECT 91.280 183.320 91.420 184.360 ;
        RECT 91.220 183.000 91.480 183.320 ;
        RECT 90.760 182.320 91.020 182.640 ;
        RECT 89.380 179.600 89.640 179.920 ;
        RECT 89.900 179.580 90.040 180.280 ;
        RECT 90.290 180.085 90.570 180.455 ;
        RECT 90.360 179.920 90.500 180.085 ;
        RECT 90.300 179.600 90.560 179.920 ;
        RECT 89.840 179.260 90.100 179.580 ;
        RECT 89.900 178.220 90.040 179.260 ;
        RECT 90.820 179.150 90.960 182.320 ;
        RECT 91.280 179.920 91.420 183.000 ;
        RECT 91.220 179.600 91.480 179.920 ;
        RECT 90.360 179.010 90.960 179.150 ;
        RECT 92.200 179.095 92.340 185.130 ;
        RECT 92.600 185.040 92.860 185.130 ;
        RECT 92.600 182.320 92.860 182.640 ;
        RECT 89.840 177.900 90.100 178.220 ;
        RECT 89.840 174.730 90.100 174.820 ;
        RECT 89.440 174.590 90.100 174.730 ;
        RECT 89.440 166.855 89.580 174.590 ;
        RECT 89.840 174.500 90.100 174.590 ;
        RECT 89.840 173.480 90.100 173.800 ;
        RECT 89.900 168.895 90.040 173.480 ;
        RECT 89.830 168.525 90.110 168.895 ;
        RECT 89.840 168.040 90.100 168.360 ;
        RECT 89.370 166.485 89.650 166.855 ;
        RECT 89.900 165.980 90.040 168.040 ;
        RECT 88.920 165.660 89.180 165.980 ;
        RECT 89.840 165.660 90.100 165.980 ;
        RECT 90.360 165.550 90.500 179.010 ;
        RECT 92.130 178.725 92.410 179.095 ;
        RECT 91.680 177.220 91.940 177.540 ;
        RECT 91.740 174.480 91.880 177.220 ;
        RECT 91.210 173.965 91.490 174.335 ;
        RECT 91.680 174.160 91.940 174.480 ;
        RECT 91.220 173.820 91.480 173.965 ;
        RECT 90.760 173.480 91.020 173.800 ;
        RECT 90.820 169.040 90.960 173.480 ;
        RECT 91.680 171.610 91.940 171.930 ;
        RECT 91.220 169.630 91.480 169.720 ;
        RECT 91.740 169.630 91.880 171.610 ;
        RECT 91.220 169.490 91.880 169.630 ;
        RECT 91.220 169.400 91.480 169.490 ;
        RECT 92.200 169.040 92.340 178.725 ;
        RECT 92.660 178.415 92.800 182.320 ;
        RECT 92.590 178.045 92.870 178.415 ;
        RECT 93.120 177.790 93.260 186.060 ;
        RECT 93.580 185.360 93.720 186.060 ;
        RECT 94.040 186.040 94.180 188.360 ;
        RECT 93.980 185.720 94.240 186.040 ;
        RECT 93.520 185.040 93.780 185.360 ;
        RECT 93.980 185.040 94.240 185.360 ;
        RECT 94.040 182.495 94.180 185.040 ;
        RECT 94.440 182.660 94.700 182.980 ;
        RECT 93.970 182.125 94.250 182.495 ;
        RECT 94.500 182.300 94.640 182.660 ;
        RECT 94.440 181.980 94.700 182.300 ;
        RECT 93.970 180.765 94.250 181.135 ;
        RECT 93.980 180.620 94.240 180.765 ;
        RECT 94.500 180.260 94.640 181.980 ;
        RECT 94.960 180.940 95.100 188.720 ;
        RECT 95.360 188.100 95.620 188.420 ;
        RECT 95.420 186.380 95.560 188.100 ;
        RECT 95.360 186.060 95.620 186.380 ;
        RECT 95.880 185.360 96.020 189.800 ;
        RECT 96.340 188.420 96.480 189.890 ;
        RECT 96.740 189.800 97.000 189.890 ;
        RECT 96.740 188.440 97.000 188.760 ;
        RECT 96.280 188.100 96.540 188.420 ;
        RECT 96.340 185.360 96.480 188.100 ;
        RECT 96.800 187.935 96.940 188.440 ;
        RECT 96.730 187.565 97.010 187.935 ;
        RECT 96.800 186.575 96.940 187.565 ;
        RECT 96.730 186.205 97.010 186.575 ;
        RECT 96.800 185.360 96.940 186.205 ;
        RECT 95.820 185.040 96.080 185.360 ;
        RECT 96.280 185.040 96.540 185.360 ;
        RECT 96.740 185.040 97.000 185.360 ;
        RECT 95.880 184.535 96.020 185.040 ;
        RECT 95.810 184.165 96.090 184.535 ;
        RECT 95.880 182.980 96.020 184.165 ;
        RECT 96.340 183.320 96.480 185.040 ;
        RECT 97.260 183.660 97.400 193.685 ;
        RECT 98.180 193.180 98.320 196.520 ;
        RECT 98.570 195.725 98.850 196.095 ;
        RECT 98.640 194.540 98.780 195.725 ;
        RECT 98.580 194.220 98.840 194.540 ;
        RECT 98.120 192.860 98.380 193.180 ;
        RECT 98.570 189.605 98.850 189.975 ;
        RECT 97.660 188.100 97.920 188.420 ;
        RECT 98.120 188.100 98.380 188.420 ;
        RECT 97.720 184.535 97.860 188.100 ;
        RECT 98.180 186.040 98.320 188.100 ;
        RECT 98.120 185.720 98.380 186.040 ;
        RECT 97.650 184.165 97.930 184.535 ;
        RECT 98.180 183.660 98.320 185.720 ;
        RECT 98.640 185.360 98.780 189.605 ;
        RECT 99.100 186.040 99.240 206.800 ;
        RECT 99.960 195.240 100.220 195.560 ;
        RECT 99.500 188.100 99.760 188.420 ;
        RECT 99.560 186.380 99.700 188.100 ;
        RECT 100.020 186.380 100.160 195.240 ;
        RECT 101.330 194.365 101.610 194.735 ;
        RECT 101.860 194.540 102.000 206.840 ;
        RECT 102.720 195.580 102.980 195.900 ;
        RECT 100.420 193.540 100.680 193.860 ;
        RECT 100.480 191.820 100.620 193.540 ;
        RECT 100.880 192.860 101.140 193.180 ;
        RECT 100.420 191.500 100.680 191.820 ;
        RECT 100.940 191.220 101.080 192.860 ;
        RECT 101.400 192.840 101.540 194.365 ;
        RECT 101.800 194.220 102.060 194.540 ;
        RECT 101.340 192.520 101.600 192.840 ;
        RECT 101.790 192.325 102.070 192.695 ;
        RECT 100.480 191.080 101.080 191.220 ;
        RECT 99.500 186.060 99.760 186.380 ;
        RECT 99.960 186.060 100.220 186.380 ;
        RECT 99.040 185.720 99.300 186.040 ;
        RECT 100.480 185.360 100.620 191.080 ;
        RECT 101.340 188.780 101.600 189.100 ;
        RECT 101.860 188.860 102.000 192.325 ;
        RECT 102.780 190.800 102.920 195.580 ;
        RECT 105.080 194.540 105.220 206.840 ;
        RECT 106.390 201.845 106.670 202.215 ;
        RECT 105.470 195.045 105.750 195.415 ;
        RECT 105.020 194.220 105.280 194.540 ;
        RECT 103.640 193.540 103.900 193.860 ;
        RECT 103.700 193.180 103.840 193.540 ;
        RECT 103.640 192.860 103.900 193.180 ;
        RECT 105.010 193.005 105.290 193.375 ;
        RECT 104.560 191.160 104.820 191.480 ;
        RECT 102.720 190.480 102.980 190.800 ;
        RECT 100.880 187.080 101.140 187.400 ;
        RECT 100.940 185.360 101.080 187.080 ;
        RECT 101.400 186.380 101.540 188.780 ;
        RECT 101.860 188.720 102.920 188.860 ;
        RECT 104.620 188.760 104.760 191.160 ;
        RECT 101.860 188.420 102.000 188.720 ;
        RECT 101.800 188.100 102.060 188.420 ;
        RECT 102.260 188.100 102.520 188.420 ;
        RECT 102.320 187.935 102.460 188.100 ;
        RECT 101.800 187.420 102.060 187.740 ;
        RECT 102.250 187.565 102.530 187.935 ;
        RECT 101.340 186.060 101.600 186.380 ;
        RECT 101.340 185.380 101.600 185.700 ;
        RECT 98.580 185.040 98.840 185.360 ;
        RECT 99.950 184.845 100.230 185.215 ;
        RECT 100.420 185.040 100.680 185.360 ;
        RECT 100.880 185.040 101.140 185.360 ;
        RECT 101.400 185.215 101.540 185.380 ;
        RECT 101.330 184.845 101.610 185.215 ;
        RECT 97.200 183.340 97.460 183.660 ;
        RECT 98.120 183.340 98.380 183.660 ;
        RECT 96.280 183.000 96.540 183.320 ;
        RECT 95.820 182.660 96.080 182.980 ;
        RECT 97.200 182.660 97.460 182.980 ;
        RECT 94.900 180.620 95.160 180.940 ;
        RECT 94.440 179.940 94.700 180.260 ;
        RECT 95.820 179.940 96.080 180.260 ;
        RECT 96.280 179.940 96.540 180.260 ;
        RECT 95.360 179.600 95.620 179.920 ;
        RECT 93.980 177.900 94.240 178.220 ;
        RECT 92.660 177.650 93.260 177.790 ;
        RECT 92.660 172.690 92.800 177.650 ;
        RECT 93.520 177.220 93.780 177.540 ;
        RECT 93.580 176.860 93.720 177.220 ;
        RECT 93.520 176.540 93.780 176.860 ;
        RECT 93.050 176.005 93.330 176.375 ;
        RECT 93.120 174.140 93.260 176.005 ;
        RECT 93.580 175.160 93.720 176.540 ;
        RECT 93.520 174.840 93.780 175.160 ;
        RECT 93.060 173.820 93.320 174.140 ;
        RECT 92.660 172.550 93.260 172.690 ;
        RECT 92.590 171.925 92.870 172.295 ;
        RECT 92.660 169.040 92.800 171.925 ;
        RECT 93.120 169.040 93.260 172.550 ;
        RECT 94.040 172.440 94.180 177.900 ;
        RECT 94.440 177.220 94.700 177.540 ;
        RECT 94.500 175.695 94.640 177.220 ;
        RECT 94.900 176.880 95.160 177.200 ;
        RECT 94.430 175.325 94.710 175.695 ;
        RECT 94.500 174.480 94.640 175.325 ;
        RECT 94.960 175.160 95.100 176.880 ;
        RECT 94.900 174.840 95.160 175.160 ;
        RECT 94.440 174.390 94.700 174.480 ;
        RECT 94.440 174.250 95.100 174.390 ;
        RECT 94.440 174.160 94.700 174.250 ;
        RECT 94.440 173.480 94.700 173.800 ;
        RECT 93.980 172.120 94.240 172.440 ;
        RECT 94.500 172.180 94.640 173.480 ;
        RECT 94.960 172.780 95.100 174.250 ;
        RECT 94.900 172.460 95.160 172.780 ;
        RECT 93.520 171.780 93.780 172.100 ;
        RECT 94.500 172.040 95.100 172.180 ;
        RECT 93.580 171.420 93.720 171.780 ;
        RECT 93.980 171.440 94.240 171.760 ;
        RECT 94.440 171.440 94.700 171.760 ;
        RECT 93.520 171.100 93.780 171.420 ;
        RECT 90.760 168.950 91.020 169.040 ;
        RECT 90.760 168.810 91.880 168.950 ;
        RECT 90.760 168.720 91.020 168.810 ;
        RECT 91.220 166.340 91.480 166.660 ;
        RECT 91.280 166.175 91.420 166.340 ;
        RECT 91.210 165.805 91.490 166.175 ;
        RECT 91.220 165.550 91.480 165.640 ;
        RECT 90.360 165.410 91.480 165.550 ;
        RECT 88.520 164.390 89.580 164.530 ;
        RECT 88.920 163.620 89.180 163.940 ;
        RECT 87.540 163.280 87.800 163.600 ;
        RECT 88.450 163.085 88.730 163.455 ;
        RECT 88.520 162.920 88.660 163.085 ;
        RECT 88.460 162.600 88.720 162.920 ;
        RECT 88.980 161.900 89.120 163.620 ;
        RECT 88.920 161.580 89.180 161.900 ;
        RECT 85.240 160.900 85.500 161.220 ;
        RECT 85.700 160.900 85.960 161.220 ;
        RECT 86.160 160.900 86.420 161.220 ;
        RECT 87.080 161.130 87.340 161.220 ;
        RECT 87.080 160.990 87.740 161.130 ;
        RECT 87.080 160.900 87.340 160.990 ;
        RECT 83.860 160.220 84.120 160.540 ;
        RECT 82.940 158.860 83.200 159.180 ;
        RECT 83.400 158.860 83.660 159.180 ;
        RECT 83.000 158.580 83.140 158.860 ;
        RECT 83.920 158.695 84.060 160.220 ;
        RECT 85.230 159.685 85.510 160.055 ;
        RECT 83.000 158.500 83.600 158.580 ;
        RECT 83.000 158.440 83.660 158.500 ;
        RECT 83.400 158.180 83.660 158.440 ;
        RECT 83.850 158.325 84.130 158.695 ;
        RECT 85.300 158.500 85.440 159.685 ;
        RECT 85.760 159.180 85.900 160.900 ;
        RECT 86.680 159.180 87.280 159.260 ;
        RECT 85.700 158.860 85.960 159.180 ;
        RECT 86.680 159.120 87.340 159.180 ;
        RECT 85.240 158.180 85.500 158.500 ;
        RECT 82.940 158.070 83.200 158.160 ;
        RECT 82.540 157.930 83.200 158.070 ;
        RECT 82.940 157.840 83.200 157.930 ;
        RECT 82.470 156.965 82.750 157.335 ;
        RECT 82.940 157.160 83.200 157.480 ;
        RECT 81.100 156.230 81.760 156.370 ;
        RECT 81.100 156.140 81.360 156.230 ;
        RECT 82.020 156.140 82.280 156.460 ;
        RECT 81.560 155.690 81.820 155.780 ;
        RECT 81.160 155.550 81.820 155.690 ;
        RECT 80.640 154.440 80.900 154.760 ;
        RECT 76.500 152.400 76.760 152.720 ;
        RECT 78.800 152.400 79.060 152.720 ;
        RECT 79.720 152.400 79.980 152.720 ;
        RECT 74.660 151.720 74.920 152.040 ;
        RECT 74.200 146.960 74.460 147.280 ;
        RECT 73.280 146.620 73.540 146.940 ;
        RECT 74.720 145.920 74.860 151.720 ;
        RECT 76.560 150.680 76.700 152.400 ;
        RECT 81.160 152.040 81.300 155.550 ;
        RECT 81.560 155.460 81.820 155.550 ;
        RECT 82.540 152.720 82.680 156.965 ;
        RECT 83.000 154.760 83.140 157.160 ;
        RECT 83.460 155.780 83.600 158.180 ;
        RECT 85.700 157.840 85.960 158.160 ;
        RECT 84.310 156.285 84.590 156.655 ;
        RECT 84.320 156.140 84.580 156.285 ;
        RECT 85.760 156.120 85.900 157.840 ;
        RECT 85.700 155.800 85.960 156.120 ;
        RECT 83.400 155.460 83.660 155.780 ;
        RECT 85.240 155.460 85.500 155.780 ;
        RECT 85.300 155.295 85.440 155.460 ;
        RECT 85.230 154.925 85.510 155.295 ;
        RECT 86.680 154.760 86.820 159.120 ;
        RECT 87.080 158.860 87.340 159.120 ;
        RECT 87.600 157.480 87.740 160.990 ;
        RECT 88.920 160.900 89.180 161.220 ;
        RECT 87.990 157.645 88.270 158.015 ;
        RECT 87.080 157.160 87.340 157.480 ;
        RECT 87.540 157.160 87.800 157.480 ;
        RECT 87.140 155.780 87.280 157.160 ;
        RECT 88.060 155.780 88.200 157.645 ;
        RECT 88.980 155.975 89.120 160.900 ;
        RECT 89.440 158.015 89.580 164.390 ;
        RECT 89.840 164.300 90.100 164.620 ;
        RECT 89.370 157.645 89.650 158.015 ;
        RECT 89.380 157.160 89.640 157.480 ;
        RECT 87.080 155.460 87.340 155.780 ;
        RECT 88.000 155.460 88.260 155.780 ;
        RECT 88.910 155.605 89.190 155.975 ;
        RECT 82.940 154.440 83.200 154.760 ;
        RECT 86.620 154.440 86.880 154.760 ;
        RECT 88.920 154.440 89.180 154.760 ;
        RECT 87.080 153.420 87.340 153.740 ;
        RECT 82.940 153.080 83.200 153.400 ;
        RECT 82.480 152.400 82.740 152.720 ;
        RECT 78.800 151.720 79.060 152.040 ;
        RECT 81.100 151.720 81.360 152.040 ;
        RECT 81.560 151.720 81.820 152.040 ;
        RECT 76.500 150.360 76.760 150.680 ;
        RECT 78.860 146.600 79.000 151.720 ;
        RECT 81.620 148.980 81.760 151.720 ;
        RECT 81.560 148.660 81.820 148.980 ;
        RECT 78.800 146.280 79.060 146.600 ;
        RECT 74.660 145.600 74.920 145.920 ;
        RECT 83.000 145.580 83.140 153.080 ;
        RECT 87.140 152.720 87.280 153.420 ;
        RECT 87.080 152.400 87.340 152.720 ;
        RECT 88.460 152.400 88.720 152.720 ;
        RECT 83.400 152.060 83.660 152.380 ;
        RECT 83.460 149.320 83.600 152.060 ;
        RECT 83.400 149.000 83.660 149.320 ;
        RECT 88.520 148.640 88.660 152.400 ;
        RECT 88.460 148.320 88.720 148.640 ;
        RECT 82.940 145.260 83.200 145.580 ;
        RECT 37.390 140.490 37.670 140.990 ;
        RECT 40.610 140.490 40.890 140.990 ;
        RECT 43.830 140.490 44.110 140.990 ;
        RECT 47.050 140.490 47.330 140.990 ;
        RECT 53.490 140.490 53.770 140.990 ;
        RECT 56.710 140.490 56.990 140.990 ;
        RECT 66.370 140.645 66.650 141.015 ;
        RECT 70.520 140.840 70.780 141.160 ;
        RECT 88.980 140.990 89.120 154.440 ;
        RECT 89.440 152.720 89.580 157.160 ;
        RECT 89.900 155.780 90.040 164.300 ;
        RECT 90.300 163.280 90.560 163.600 ;
        RECT 90.360 161.220 90.500 163.280 ;
        RECT 90.300 160.900 90.560 161.220 ;
        RECT 90.300 160.055 90.560 160.200 ;
        RECT 90.290 159.685 90.570 160.055 ;
        RECT 90.300 157.390 90.560 157.480 ;
        RECT 90.820 157.390 90.960 165.410 ;
        RECT 91.220 165.320 91.480 165.410 ;
        RECT 91.740 163.455 91.880 168.810 ;
        RECT 92.140 168.720 92.400 169.040 ;
        RECT 92.600 168.720 92.860 169.040 ;
        RECT 93.060 168.720 93.320 169.040 ;
        RECT 92.200 166.660 92.340 168.720 ;
        RECT 92.140 166.340 92.400 166.660 ;
        RECT 92.200 164.280 92.340 166.340 ;
        RECT 92.660 166.230 92.800 168.720 ;
        RECT 93.120 166.910 93.260 168.720 ;
        RECT 93.580 168.700 93.720 171.100 ;
        RECT 94.040 170.060 94.180 171.440 ;
        RECT 93.980 169.740 94.240 170.060 ;
        RECT 94.500 169.040 94.640 171.440 ;
        RECT 94.960 169.720 95.100 172.040 ;
        RECT 94.900 169.400 95.160 169.720 ;
        RECT 94.440 168.720 94.700 169.040 ;
        RECT 93.520 168.380 93.780 168.700 ;
        RECT 94.500 167.340 94.640 168.720 ;
        RECT 94.900 168.380 95.160 168.700 ;
        RECT 94.440 167.020 94.700 167.340 ;
        RECT 93.520 166.910 93.780 167.000 ;
        RECT 93.120 166.770 93.780 166.910 ;
        RECT 94.960 166.855 95.100 168.380 ;
        RECT 93.520 166.680 93.780 166.770 ;
        RECT 93.060 166.230 93.320 166.320 ;
        RECT 92.660 166.090 93.320 166.230 ;
        RECT 93.060 166.000 93.320 166.090 ;
        RECT 93.580 165.495 93.720 166.680 ;
        RECT 94.890 166.485 95.170 166.855 ;
        RECT 93.980 166.000 94.240 166.320 ;
        RECT 94.040 165.640 94.180 166.000 ;
        RECT 94.430 165.805 94.710 166.175 ;
        RECT 93.510 165.125 93.790 165.495 ;
        RECT 93.980 165.320 94.240 165.640 ;
        RECT 92.140 163.960 92.400 164.280 ;
        RECT 91.670 163.085 91.950 163.455 ;
        RECT 92.600 162.940 92.860 163.260 ;
        RECT 92.140 162.600 92.400 162.920 ;
        RECT 91.220 159.880 91.480 160.200 ;
        RECT 91.280 158.160 91.420 159.880 ;
        RECT 92.200 158.840 92.340 162.600 ;
        RECT 92.140 158.520 92.400 158.840 ;
        RECT 91.220 157.840 91.480 158.160 ;
        RECT 90.300 157.250 90.960 157.390 ;
        RECT 90.300 157.160 90.560 157.250 ;
        RECT 91.680 157.160 91.940 157.480 ;
        RECT 90.360 156.460 90.500 157.160 ;
        RECT 90.300 156.140 90.560 156.460 ;
        RECT 89.840 155.460 90.100 155.780 ;
        RECT 89.380 152.400 89.640 152.720 ;
        RECT 91.740 150.680 91.880 157.160 ;
        RECT 91.680 150.360 91.940 150.680 ;
        RECT 92.660 150.000 92.800 162.940 ;
        RECT 94.500 161.900 94.640 165.805 ;
        RECT 94.900 165.320 95.160 165.640 ;
        RECT 93.060 161.580 93.320 161.900 ;
        RECT 94.440 161.580 94.700 161.900 ;
        RECT 93.120 158.500 93.260 161.580 ;
        RECT 94.960 161.130 95.100 165.320 ;
        RECT 93.580 160.990 95.100 161.130 ;
        RECT 93.060 158.180 93.320 158.500 ;
        RECT 93.580 157.335 93.720 160.990 ;
        RECT 95.420 160.880 95.560 179.600 ;
        RECT 95.880 178.220 96.020 179.940 ;
        RECT 95.820 177.900 96.080 178.220 ;
        RECT 96.340 177.880 96.480 179.940 ;
        RECT 96.740 178.920 97.000 179.240 ;
        RECT 96.280 177.560 96.540 177.880 ;
        RECT 95.820 177.220 96.080 177.540 ;
        RECT 95.880 173.800 96.020 177.220 ;
        RECT 96.340 173.800 96.480 177.560 ;
        RECT 95.820 173.480 96.080 173.800 ;
        RECT 96.280 173.480 96.540 173.800 ;
        RECT 96.280 171.780 96.540 172.100 ;
        RECT 95.820 171.100 96.080 171.420 ;
        RECT 95.880 167.340 96.020 171.100 ;
        RECT 95.820 167.020 96.080 167.340 ;
        RECT 96.340 166.740 96.480 171.780 ;
        RECT 96.800 167.340 96.940 178.920 ;
        RECT 97.260 175.695 97.400 182.660 ;
        RECT 97.660 179.260 97.920 179.580 ;
        RECT 98.580 179.260 98.840 179.580 ;
        RECT 97.720 179.095 97.860 179.260 ;
        RECT 97.650 178.725 97.930 179.095 ;
        RECT 98.110 176.005 98.390 176.375 ;
        RECT 97.190 175.325 97.470 175.695 ;
        RECT 97.200 174.840 97.460 175.160 ;
        RECT 97.260 171.080 97.400 174.840 ;
        RECT 97.660 174.500 97.920 174.820 ;
        RECT 97.200 170.760 97.460 171.080 ;
        RECT 97.720 170.935 97.860 174.500 ;
        RECT 98.180 171.420 98.320 176.005 ;
        RECT 98.640 172.295 98.780 179.260 ;
        RECT 99.500 178.920 99.760 179.240 ;
        RECT 99.040 176.200 99.300 176.520 ;
        RECT 99.100 174.335 99.240 176.200 ;
        RECT 99.560 175.500 99.700 178.920 ;
        RECT 100.020 176.940 100.160 184.845 ;
        RECT 100.420 182.660 100.680 182.980 ;
        RECT 100.480 181.135 100.620 182.660 ;
        RECT 100.880 182.495 101.140 182.640 ;
        RECT 100.870 182.125 101.150 182.495 ;
        RECT 100.870 181.445 101.150 181.815 ;
        RECT 101.340 181.640 101.600 181.960 ;
        RECT 100.410 180.765 100.690 181.135 ;
        RECT 100.940 179.920 101.080 181.445 ;
        RECT 100.880 179.600 101.140 179.920 ;
        RECT 100.880 177.220 101.140 177.540 ;
        RECT 100.020 176.860 100.620 176.940 ;
        RECT 100.020 176.800 100.680 176.860 ;
        RECT 100.420 176.540 100.680 176.800 ;
        RECT 99.960 176.200 100.220 176.520 ;
        RECT 100.020 175.695 100.160 176.200 ;
        RECT 99.500 175.180 99.760 175.500 ;
        RECT 99.950 175.325 100.230 175.695 ;
        RECT 100.940 175.015 101.080 177.220 ;
        RECT 99.490 174.645 99.770 175.015 ;
        RECT 100.870 174.645 101.150 175.015 ;
        RECT 99.030 173.965 99.310 174.335 ;
        RECT 99.040 173.480 99.300 173.800 ;
        RECT 98.570 171.925 98.850 172.295 ;
        RECT 99.100 172.100 99.240 173.480 ;
        RECT 99.560 172.780 99.700 174.645 ;
        RECT 100.880 174.160 101.140 174.480 ;
        RECT 100.420 173.820 100.680 174.140 ;
        RECT 99.500 172.460 99.760 172.780 ;
        RECT 99.960 172.120 100.220 172.440 ;
        RECT 99.040 171.780 99.300 172.100 ;
        RECT 98.120 171.100 98.380 171.420 ;
        RECT 97.650 170.565 97.930 170.935 ;
        RECT 97.200 169.060 97.460 169.380 ;
        RECT 96.740 167.020 97.000 167.340 ;
        RECT 95.820 166.340 96.080 166.660 ;
        RECT 96.340 166.600 96.940 166.740 ;
        RECT 95.880 163.940 96.020 166.340 ;
        RECT 96.800 166.320 96.940 166.600 ;
        RECT 96.280 166.175 96.540 166.320 ;
        RECT 96.270 165.805 96.550 166.175 ;
        RECT 96.740 166.000 97.000 166.320 ;
        RECT 95.820 163.620 96.080 163.940 ;
        RECT 95.810 161.725 96.090 162.095 ;
        RECT 95.880 160.880 96.020 161.725 ;
        RECT 96.340 161.560 96.480 165.805 ;
        RECT 96.280 161.240 96.540 161.560 ;
        RECT 95.360 160.560 95.620 160.880 ;
        RECT 95.820 160.560 96.080 160.880 ;
        RECT 94.440 160.220 94.700 160.540 ;
        RECT 94.900 160.220 95.160 160.540 ;
        RECT 93.980 158.520 94.240 158.840 ;
        RECT 94.040 158.160 94.180 158.520 ;
        RECT 94.500 158.160 94.640 160.220 ;
        RECT 93.980 157.840 94.240 158.160 ;
        RECT 94.440 157.840 94.700 158.160 ;
        RECT 93.510 156.965 93.790 157.335 ;
        RECT 94.500 153.255 94.640 157.840 ;
        RECT 94.960 156.460 95.100 160.220 ;
        RECT 95.880 158.840 96.020 160.560 ;
        RECT 95.350 158.325 95.630 158.695 ;
        RECT 95.820 158.520 96.080 158.840 ;
        RECT 95.420 158.160 95.560 158.325 ;
        RECT 95.360 157.840 95.620 158.160 ;
        RECT 94.900 156.140 95.160 156.460 ;
        RECT 95.420 156.120 95.560 157.840 ;
        RECT 95.360 155.800 95.620 156.120 ;
        RECT 94.430 152.885 94.710 153.255 ;
        RECT 92.600 149.680 92.860 150.000 ;
        RECT 92.140 148.660 92.400 148.980 ;
        RECT 92.200 140.990 92.340 148.660 ;
        RECT 95.420 148.640 95.560 155.800 ;
        RECT 96.800 152.380 96.940 166.000 ;
        RECT 97.260 161.220 97.400 169.060 ;
        RECT 97.720 169.040 97.860 170.565 ;
        RECT 97.660 168.720 97.920 169.040 ;
        RECT 97.650 166.485 97.930 166.855 ;
        RECT 98.180 166.660 98.320 171.100 ;
        RECT 98.580 170.760 98.840 171.080 ;
        RECT 98.640 169.040 98.780 170.760 ;
        RECT 99.100 169.040 99.240 171.780 ;
        RECT 100.020 170.060 100.160 172.120 ;
        RECT 99.960 169.740 100.220 170.060 ;
        RECT 100.480 169.720 100.620 173.820 ;
        RECT 100.420 169.400 100.680 169.720 ;
        RECT 98.580 168.720 98.840 169.040 ;
        RECT 99.040 168.720 99.300 169.040 ;
        RECT 100.410 168.525 100.690 168.895 ;
        RECT 98.580 168.040 98.840 168.360 ;
        RECT 97.660 166.340 97.920 166.485 ;
        RECT 98.120 166.340 98.380 166.660 ;
        RECT 97.720 164.620 97.860 166.340 ;
        RECT 97.660 164.300 97.920 164.620 ;
        RECT 98.180 163.600 98.320 166.340 ;
        RECT 98.120 163.280 98.380 163.600 ;
        RECT 97.650 161.725 97.930 162.095 ;
        RECT 97.200 160.900 97.460 161.220 ;
        RECT 97.720 160.200 97.860 161.725 ;
        RECT 98.120 160.790 98.380 160.880 ;
        RECT 98.640 160.790 98.780 168.040 ;
        RECT 99.960 167.020 100.220 167.340 ;
        RECT 100.020 164.280 100.160 167.020 ;
        RECT 100.480 164.620 100.620 168.525 ;
        RECT 100.940 166.855 101.080 174.160 ;
        RECT 101.400 173.800 101.540 181.640 ;
        RECT 101.860 180.455 102.000 187.420 ;
        RECT 102.780 185.950 102.920 188.720 ;
        RECT 103.170 188.245 103.450 188.615 ;
        RECT 104.560 188.440 104.820 188.760 ;
        RECT 103.240 188.080 103.380 188.245 ;
        RECT 103.180 187.760 103.440 188.080 ;
        RECT 105.080 187.400 105.220 193.005 ;
        RECT 105.540 188.330 105.680 195.045 ;
        RECT 106.460 193.860 106.600 201.845 ;
        RECT 108.300 200.175 108.440 206.840 ;
        RECT 111.520 200.855 111.660 206.840 ;
        RECT 111.450 200.485 111.730 200.855 ;
        RECT 108.230 199.805 108.510 200.175 ;
        RECT 111.450 198.445 111.730 198.815 ;
        RECT 107.320 193.880 107.580 194.200 ;
        RECT 106.400 193.540 106.660 193.860 ;
        RECT 106.860 193.540 107.120 193.860 ;
        RECT 106.920 191.820 107.060 193.540 ;
        RECT 106.860 191.500 107.120 191.820 ;
        RECT 106.860 190.480 107.120 190.800 ;
        RECT 105.540 188.190 106.140 188.330 ;
        RECT 106.390 188.245 106.670 188.615 ;
        RECT 106.920 188.420 107.060 190.480 ;
        RECT 105.480 187.420 105.740 187.740 ;
        RECT 103.170 186.885 103.450 187.255 ;
        RECT 104.090 186.885 104.370 187.255 ;
        RECT 105.020 187.080 105.280 187.400 ;
        RECT 103.240 186.040 103.380 186.885 ;
        RECT 102.320 185.810 102.920 185.950 ;
        RECT 102.320 185.270 102.460 185.810 ;
        RECT 103.180 185.720 103.440 186.040 ;
        RECT 103.180 185.270 103.440 185.360 ;
        RECT 102.320 185.130 102.920 185.270 ;
        RECT 102.260 184.360 102.520 184.680 ;
        RECT 102.320 183.320 102.460 184.360 ;
        RECT 102.260 183.000 102.520 183.320 ;
        RECT 102.780 182.980 102.920 185.130 ;
        RECT 103.180 185.130 103.840 185.270 ;
        RECT 103.180 185.040 103.440 185.130 ;
        RECT 103.700 183.570 103.840 185.130 ;
        RECT 104.160 183.660 104.300 186.885 ;
        RECT 104.550 186.205 104.830 186.575 ;
        RECT 105.080 186.380 105.220 187.080 ;
        RECT 104.620 186.040 104.760 186.205 ;
        RECT 105.020 186.060 105.280 186.380 ;
        RECT 104.560 185.720 104.820 186.040 ;
        RECT 105.540 185.700 105.680 187.420 ;
        RECT 105.480 185.380 105.740 185.700 ;
        RECT 106.000 185.360 106.140 188.190 ;
        RECT 106.460 186.575 106.600 188.245 ;
        RECT 106.860 188.100 107.120 188.420 ;
        RECT 107.380 188.330 107.520 193.880 ;
        RECT 110.540 193.200 110.800 193.520 ;
        RECT 109.160 192.520 109.420 192.840 ;
        RECT 107.770 190.965 108.050 191.335 ;
        RECT 109.220 191.140 109.360 192.520 ;
        RECT 107.840 188.330 107.980 190.965 ;
        RECT 108.700 190.820 108.960 191.140 ;
        RECT 109.160 190.820 109.420 191.140 ;
        RECT 108.240 190.480 108.500 190.800 ;
        RECT 108.300 188.760 108.440 190.480 ;
        RECT 108.760 189.295 108.900 190.820 ;
        RECT 108.690 188.925 108.970 189.295 ;
        RECT 108.240 188.440 108.500 188.760 ;
        RECT 107.380 188.190 107.980 188.330 ;
        RECT 108.240 187.990 108.500 188.080 ;
        RECT 107.380 187.850 108.500 187.990 ;
        RECT 108.700 187.935 108.960 188.080 ;
        RECT 106.390 186.205 106.670 186.575 ;
        RECT 106.400 186.060 106.660 186.205 ;
        RECT 106.860 185.720 107.120 186.040 ;
        RECT 105.940 185.040 106.200 185.360 ;
        RECT 104.560 184.360 104.820 184.680 ;
        RECT 103.240 183.430 103.840 183.570 ;
        RECT 102.720 182.660 102.980 182.980 ;
        RECT 102.260 181.980 102.520 182.300 ;
        RECT 102.320 181.815 102.460 181.980 ;
        RECT 102.720 181.870 102.980 181.960 ;
        RECT 103.240 181.870 103.380 183.430 ;
        RECT 104.100 183.340 104.360 183.660 ;
        RECT 104.620 182.980 104.760 184.360 ;
        RECT 105.940 183.000 106.200 183.320 ;
        RECT 103.640 182.890 103.900 182.980 ;
        RECT 103.640 182.750 104.300 182.890 ;
        RECT 103.640 182.660 103.900 182.750 ;
        RECT 102.250 181.445 102.530 181.815 ;
        RECT 102.720 181.730 103.380 181.870 ;
        RECT 102.720 181.640 102.980 181.730 ;
        RECT 103.630 181.445 103.910 181.815 ;
        RECT 103.180 180.620 103.440 180.940 ;
        RECT 101.790 180.085 102.070 180.455 ;
        RECT 102.260 179.600 102.520 179.920 ;
        RECT 102.720 179.600 102.980 179.920 ;
        RECT 101.800 176.880 102.060 177.200 ;
        RECT 101.860 175.015 102.000 176.880 ;
        RECT 101.790 174.645 102.070 175.015 ;
        RECT 102.320 174.220 102.460 179.600 ;
        RECT 102.780 174.730 102.920 179.600 ;
        RECT 103.240 177.540 103.380 180.620 ;
        RECT 103.700 179.920 103.840 181.445 ;
        RECT 104.160 180.455 104.300 182.750 ;
        RECT 104.560 182.660 104.820 182.980 ;
        RECT 104.090 180.085 104.370 180.455 ;
        RECT 103.640 179.600 103.900 179.920 ;
        RECT 104.100 179.600 104.360 179.920 ;
        RECT 103.640 178.920 103.900 179.240 ;
        RECT 103.180 177.220 103.440 177.540 ;
        RECT 103.180 176.200 103.440 176.520 ;
        RECT 103.240 175.060 103.380 176.200 ;
        RECT 103.700 175.410 103.840 178.920 ;
        RECT 104.160 177.880 104.300 179.600 ;
        RECT 104.620 179.580 104.760 182.660 ;
        RECT 106.000 182.300 106.140 183.000 ;
        RECT 106.400 182.890 106.660 182.980 ;
        RECT 106.920 182.890 107.060 185.720 ;
        RECT 107.380 185.360 107.520 187.850 ;
        RECT 108.240 187.760 108.500 187.850 ;
        RECT 108.690 187.565 108.970 187.935 ;
        RECT 107.780 187.080 108.040 187.400 ;
        RECT 107.320 185.040 107.580 185.360 ;
        RECT 107.840 184.680 107.980 187.080 ;
        RECT 109.220 185.950 109.360 190.820 ;
        RECT 109.620 190.140 109.880 190.460 ;
        RECT 109.680 186.040 109.820 190.140 ;
        RECT 110.080 187.080 110.340 187.400 ;
        RECT 108.760 185.810 109.360 185.950 ;
        RECT 108.240 185.040 108.500 185.360 ;
        RECT 107.780 184.360 108.040 184.680 ;
        RECT 107.780 183.230 108.040 183.320 ;
        RECT 106.400 182.750 107.060 182.890 ;
        RECT 106.400 182.660 106.660 182.750 ;
        RECT 105.020 182.210 105.280 182.300 ;
        RECT 105.020 182.070 105.680 182.210 ;
        RECT 105.020 181.980 105.280 182.070 ;
        RECT 105.020 179.940 105.280 180.260 ;
        RECT 104.560 179.260 104.820 179.580 ;
        RECT 104.550 178.725 104.830 179.095 ;
        RECT 104.100 177.560 104.360 177.880 ;
        RECT 104.620 177.540 104.760 178.725 ;
        RECT 105.080 178.220 105.220 179.940 ;
        RECT 105.540 179.920 105.680 182.070 ;
        RECT 105.940 181.980 106.200 182.300 ;
        RECT 106.000 180.940 106.140 181.980 ;
        RECT 105.940 180.620 106.200 180.940 ;
        RECT 106.920 180.340 107.060 182.750 ;
        RECT 106.000 180.200 107.060 180.340 ;
        RECT 107.380 183.090 108.040 183.230 ;
        RECT 105.480 179.600 105.740 179.920 ;
        RECT 105.020 177.900 105.280 178.220 ;
        RECT 105.540 177.540 105.680 179.600 ;
        RECT 106.000 179.095 106.140 180.200 ;
        RECT 106.800 179.830 107.060 179.920 ;
        RECT 106.460 179.690 107.060 179.830 ;
        RECT 105.930 178.725 106.210 179.095 ;
        RECT 104.560 177.220 104.820 177.540 ;
        RECT 105.020 177.220 105.280 177.540 ;
        RECT 105.480 177.220 105.740 177.540 ;
        RECT 104.560 176.540 104.820 176.860 ;
        RECT 105.075 176.770 105.215 177.220 ;
        RECT 105.075 176.630 105.220 176.770 ;
        RECT 104.620 175.580 104.760 176.540 ;
        RECT 105.080 176.375 105.220 176.630 ;
        RECT 105.010 176.005 105.290 176.375 ;
        RECT 104.620 175.440 105.220 175.580 ;
        RECT 103.700 175.270 104.300 175.410 ;
        RECT 103.240 174.920 103.840 175.060 ;
        RECT 102.780 174.590 103.380 174.730 ;
        RECT 101.860 174.080 102.460 174.220 ;
        RECT 101.340 173.480 101.600 173.800 ;
        RECT 101.400 167.000 101.540 173.480 ;
        RECT 101.860 171.760 102.000 174.080 ;
        RECT 102.720 173.820 102.980 174.140 ;
        RECT 102.260 173.480 102.520 173.800 ;
        RECT 102.320 172.100 102.460 173.480 ;
        RECT 102.260 171.780 102.520 172.100 ;
        RECT 101.800 171.440 102.060 171.760 ;
        RECT 102.320 170.060 102.460 171.780 ;
        RECT 102.260 169.740 102.520 170.060 ;
        RECT 101.800 169.400 102.060 169.720 ;
        RECT 101.860 169.040 102.000 169.400 ;
        RECT 101.800 168.720 102.060 169.040 ;
        RECT 102.260 168.720 102.520 169.040 ;
        RECT 100.870 166.485 101.150 166.855 ;
        RECT 101.340 166.680 101.600 167.000 ;
        RECT 101.860 166.060 102.000 168.720 ;
        RECT 102.320 166.855 102.460 168.720 ;
        RECT 102.250 166.485 102.530 166.855 ;
        RECT 100.940 165.920 102.000 166.060 ;
        RECT 100.420 164.300 100.680 164.620 ;
        RECT 99.040 163.960 99.300 164.280 ;
        RECT 99.960 163.960 100.220 164.280 ;
        RECT 99.100 163.600 99.240 163.960 ;
        RECT 99.040 163.280 99.300 163.600 ;
        RECT 99.500 163.280 99.760 163.600 ;
        RECT 99.100 161.560 99.240 163.280 ;
        RECT 99.560 162.920 99.700 163.280 ;
        RECT 99.500 162.600 99.760 162.920 ;
        RECT 99.040 161.240 99.300 161.560 ;
        RECT 100.020 161.300 100.160 163.960 ;
        RECT 100.940 163.600 101.080 165.920 ;
        RECT 102.250 165.805 102.530 166.175 ;
        RECT 101.340 165.320 101.600 165.640 ;
        RECT 100.420 163.280 100.680 163.600 ;
        RECT 100.880 163.280 101.140 163.600 ;
        RECT 99.560 161.160 100.160 161.300 ;
        RECT 98.120 160.650 98.780 160.790 ;
        RECT 99.040 160.735 99.300 160.880 ;
        RECT 98.120 160.560 98.380 160.650 ;
        RECT 97.660 159.880 97.920 160.200 ;
        RECT 98.180 159.375 98.320 160.560 ;
        RECT 99.030 160.365 99.310 160.735 ;
        RECT 98.580 159.880 98.840 160.200 ;
        RECT 98.110 159.005 98.390 159.375 ;
        RECT 98.640 157.480 98.780 159.880 ;
        RECT 99.560 158.160 99.700 161.160 ;
        RECT 99.960 160.735 100.220 160.880 ;
        RECT 99.950 160.365 100.230 160.735 ;
        RECT 100.480 158.840 100.620 163.280 ;
        RECT 100.420 158.520 100.680 158.840 ;
        RECT 99.500 157.840 99.760 158.160 ;
        RECT 100.420 157.840 100.680 158.160 ;
        RECT 98.580 157.160 98.840 157.480 ;
        RECT 100.480 153.740 100.620 157.840 ;
        RECT 100.880 154.440 101.140 154.760 ;
        RECT 100.940 153.740 101.080 154.440 ;
        RECT 100.420 153.420 100.680 153.740 ;
        RECT 100.880 153.420 101.140 153.740 ;
        RECT 96.740 152.060 97.000 152.380 ;
        RECT 101.400 149.660 101.540 165.320 ;
        RECT 101.800 162.940 102.060 163.260 ;
        RECT 101.860 161.220 102.000 162.940 ;
        RECT 101.800 160.900 102.060 161.220 ;
        RECT 101.800 158.070 102.060 158.160 ;
        RECT 102.320 158.070 102.460 165.805 ;
        RECT 102.780 164.620 102.920 173.820 ;
        RECT 103.240 172.100 103.380 174.590 ;
        RECT 103.180 171.780 103.440 172.100 ;
        RECT 103.700 169.460 103.840 174.920 ;
        RECT 104.160 174.390 104.300 175.270 ;
        RECT 105.080 174.820 105.220 175.440 ;
        RECT 106.460 175.160 106.600 179.690 ;
        RECT 106.800 179.600 107.060 179.690 ;
        RECT 106.400 174.840 106.660 175.160 ;
        RECT 105.020 174.500 105.280 174.820 ;
        RECT 104.560 174.390 104.820 174.480 ;
        RECT 104.160 174.250 104.820 174.390 ;
        RECT 104.560 174.160 104.820 174.250 ;
        RECT 106.860 174.160 107.120 174.480 ;
        RECT 105.480 173.480 105.740 173.800 ;
        RECT 105.020 169.740 105.280 170.060 ;
        RECT 103.240 169.320 103.840 169.460 ;
        RECT 103.240 166.175 103.380 169.320 ;
        RECT 103.640 168.720 103.900 169.040 ;
        RECT 103.170 165.805 103.450 166.175 ;
        RECT 103.180 165.495 103.440 165.640 ;
        RECT 103.170 165.125 103.450 165.495 ;
        RECT 102.720 164.300 102.980 164.620 ;
        RECT 103.180 163.510 103.440 163.600 ;
        RECT 103.700 163.510 103.840 168.720 ;
        RECT 104.090 168.525 104.370 168.895 ;
        RECT 104.100 168.380 104.360 168.525 ;
        RECT 105.080 166.660 105.220 169.740 ;
        RECT 105.540 166.660 105.680 173.480 ;
        RECT 106.400 171.780 106.660 172.100 ;
        RECT 105.940 170.760 106.200 171.080 ;
        RECT 106.000 169.040 106.140 170.760 ;
        RECT 105.940 168.720 106.200 169.040 ;
        RECT 105.940 166.680 106.200 167.000 ;
        RECT 104.100 166.340 104.360 166.660 ;
        RECT 105.020 166.340 105.280 166.660 ;
        RECT 105.480 166.340 105.740 166.660 ;
        RECT 104.160 163.600 104.300 166.340 ;
        RECT 104.550 163.765 104.830 164.135 ;
        RECT 103.180 163.370 103.840 163.510 ;
        RECT 103.180 163.280 103.440 163.370 ;
        RECT 104.100 163.280 104.360 163.600 ;
        RECT 103.240 161.900 103.380 163.280 ;
        RECT 103.640 162.600 103.900 162.920 ;
        RECT 103.180 161.580 103.440 161.900 ;
        RECT 103.700 160.880 103.840 162.600 ;
        RECT 104.620 161.220 104.760 163.765 ;
        RECT 105.540 162.920 105.680 166.340 ;
        RECT 105.010 162.405 105.290 162.775 ;
        RECT 105.480 162.600 105.740 162.920 ;
        RECT 104.100 160.900 104.360 161.220 ;
        RECT 104.560 160.900 104.820 161.220 ;
        RECT 103.640 160.560 103.900 160.880 ;
        RECT 102.710 159.005 102.990 159.375 ;
        RECT 102.780 158.160 102.920 159.005 ;
        RECT 104.160 158.840 104.300 160.900 ;
        RECT 104.100 158.520 104.360 158.840 ;
        RECT 101.800 157.930 102.460 158.070 ;
        RECT 101.800 157.840 102.060 157.930 ;
        RECT 102.720 157.840 102.980 158.160 ;
        RECT 103.180 157.500 103.440 157.820 ;
        RECT 101.800 156.140 102.060 156.460 ;
        RECT 101.860 151.020 102.000 156.140 ;
        RECT 103.240 155.780 103.380 157.500 ;
        RECT 103.180 155.460 103.440 155.780 ;
        RECT 103.640 155.120 103.900 155.440 ;
        RECT 103.700 152.380 103.840 155.120 ;
        RECT 105.080 154.760 105.220 162.405 ;
        RECT 106.000 157.480 106.140 166.680 ;
        RECT 106.460 165.640 106.600 171.780 ;
        RECT 106.400 165.320 106.660 165.640 ;
        RECT 106.920 158.500 107.060 174.160 ;
        RECT 107.380 173.800 107.520 183.090 ;
        RECT 107.780 183.000 108.040 183.090 ;
        RECT 107.780 181.640 108.040 181.960 ;
        RECT 107.840 180.940 107.980 181.640 ;
        RECT 107.780 180.620 108.040 180.940 ;
        RECT 107.770 180.085 108.050 180.455 ;
        RECT 107.840 179.920 107.980 180.085 ;
        RECT 107.780 179.600 108.040 179.920 ;
        RECT 107.770 178.725 108.050 179.095 ;
        RECT 107.840 175.160 107.980 178.725 ;
        RECT 108.300 178.220 108.440 185.040 ;
        RECT 108.760 182.300 108.900 185.810 ;
        RECT 109.620 185.720 109.880 186.040 ;
        RECT 109.160 185.040 109.420 185.360 ;
        RECT 109.220 184.535 109.360 185.040 ;
        RECT 109.150 184.165 109.430 184.535 ;
        RECT 109.620 183.000 109.880 183.320 ;
        RECT 108.700 181.980 108.960 182.300 ;
        RECT 109.160 181.640 109.420 181.960 ;
        RECT 109.220 180.455 109.360 181.640 ;
        RECT 109.150 180.085 109.430 180.455 ;
        RECT 108.700 178.920 108.960 179.240 ;
        RECT 108.240 177.900 108.500 178.220 ;
        RECT 108.300 175.160 108.440 177.900 ;
        RECT 107.780 174.840 108.040 175.160 ;
        RECT 108.240 174.840 108.500 175.160 ;
        RECT 108.760 174.820 108.900 178.920 ;
        RECT 109.220 177.880 109.360 180.085 ;
        RECT 109.160 177.560 109.420 177.880 ;
        RECT 109.160 176.200 109.420 176.520 ;
        RECT 109.220 174.820 109.360 176.200 ;
        RECT 108.700 174.500 108.960 174.820 ;
        RECT 109.160 174.500 109.420 174.820 ;
        RECT 108.240 174.160 108.500 174.480 ;
        RECT 107.320 173.480 107.580 173.800 ;
        RECT 108.300 172.295 108.440 174.160 ;
        RECT 108.230 171.925 108.510 172.295 ;
        RECT 109.220 172.100 109.360 174.500 ;
        RECT 109.160 171.780 109.420 172.100 ;
        RECT 108.240 170.760 108.500 171.080 ;
        RECT 107.780 168.895 108.040 169.040 ;
        RECT 107.770 168.525 108.050 168.895 ;
        RECT 107.780 166.680 108.040 167.000 ;
        RECT 107.840 163.455 107.980 166.680 ;
        RECT 107.770 163.085 108.050 163.455 ;
        RECT 108.300 160.735 108.440 170.760 ;
        RECT 109.220 169.720 109.360 171.780 ;
        RECT 109.680 170.060 109.820 183.000 ;
        RECT 110.140 174.820 110.280 187.080 ;
        RECT 110.600 186.380 110.740 193.200 ;
        RECT 111.000 192.860 111.260 193.180 ;
        RECT 111.060 190.800 111.200 192.860 ;
        RECT 111.000 190.480 111.260 190.800 ;
        RECT 111.520 188.420 111.660 198.445 ;
        RECT 114.740 194.540 114.880 206.840 ;
        RECT 117.960 206.720 118.560 206.840 ;
        RECT 114.680 194.220 114.940 194.540 ;
        RECT 111.920 193.540 112.180 193.860 ;
        RECT 116.520 193.540 116.780 193.860 ;
        RECT 111.980 190.800 112.120 193.540 ;
        RECT 115.600 192.860 115.860 193.180 ;
        RECT 112.380 192.520 112.640 192.840 ;
        RECT 114.220 192.520 114.480 192.840 ;
        RECT 112.440 191.820 112.580 192.520 ;
        RECT 112.380 191.500 112.640 191.820 ;
        RECT 113.760 190.820 114.020 191.140 ;
        RECT 111.920 190.710 112.180 190.800 ;
        RECT 113.300 190.710 113.560 190.800 ;
        RECT 111.920 190.570 113.560 190.710 ;
        RECT 111.920 190.480 112.180 190.570 ;
        RECT 113.300 190.480 113.560 190.570 ;
        RECT 113.820 189.975 113.960 190.820 ;
        RECT 113.750 189.605 114.030 189.975 ;
        RECT 111.460 188.100 111.720 188.420 ;
        RECT 110.540 186.060 110.800 186.380 ;
        RECT 111.920 185.950 112.180 186.040 ;
        RECT 111.520 185.810 112.180 185.950 ;
        RECT 111.520 185.780 111.660 185.810 ;
        RECT 110.600 185.640 111.660 185.780 ;
        RECT 111.920 185.720 112.180 185.810 ;
        RECT 110.600 183.175 110.740 185.640 ;
        RECT 112.830 185.525 113.110 185.895 ;
        RECT 112.900 185.360 113.040 185.525 ;
        RECT 112.840 185.040 113.100 185.360 ;
        RECT 113.300 185.040 113.560 185.360 ;
        RECT 113.760 185.040 114.020 185.360 ;
        RECT 112.370 184.165 112.650 184.535 ;
        RECT 112.840 184.360 113.100 184.680 ;
        RECT 111.460 183.340 111.720 183.660 ;
        RECT 110.530 182.805 110.810 183.175 ;
        RECT 111.000 182.660 111.260 182.980 ;
        RECT 111.060 182.300 111.200 182.660 ;
        RECT 110.540 181.980 110.800 182.300 ;
        RECT 111.000 181.980 111.260 182.300 ;
        RECT 110.600 180.455 110.740 181.980 ;
        RECT 111.060 180.940 111.200 181.980 ;
        RECT 111.000 180.620 111.260 180.940 ;
        RECT 110.530 180.085 110.810 180.455 ;
        RECT 111.520 179.920 111.660 183.340 ;
        RECT 111.920 180.620 112.180 180.940 ;
        RECT 111.980 179.920 112.120 180.620 ;
        RECT 110.540 179.830 110.800 179.920 ;
        RECT 110.540 179.690 111.200 179.830 ;
        RECT 110.540 179.600 110.800 179.690 ;
        RECT 110.540 178.920 110.800 179.240 ;
        RECT 111.060 179.150 111.200 179.690 ;
        RECT 111.460 179.600 111.720 179.920 ;
        RECT 111.920 179.600 112.180 179.920 ;
        RECT 111.060 179.010 112.120 179.150 ;
        RECT 110.080 174.500 110.340 174.820 ;
        RECT 110.600 172.295 110.740 178.920 ;
        RECT 111.000 176.540 111.260 176.860 ;
        RECT 110.530 171.925 110.810 172.295 ;
        RECT 111.060 170.935 111.200 176.540 ;
        RECT 111.980 174.480 112.120 179.010 ;
        RECT 112.440 176.430 112.580 184.165 ;
        RECT 112.900 183.320 113.040 184.360 ;
        RECT 112.840 183.000 113.100 183.320 ;
        RECT 113.360 180.940 113.500 185.040 ;
        RECT 113.820 180.940 113.960 185.040 ;
        RECT 114.280 184.680 114.420 192.520 ;
        RECT 115.660 190.800 115.800 192.860 ;
        RECT 115.600 190.480 115.860 190.800 ;
        RECT 114.680 188.100 114.940 188.420 ;
        RECT 114.220 184.360 114.480 184.680 ;
        RECT 113.300 180.620 113.560 180.940 ;
        RECT 113.760 180.620 114.020 180.940 ;
        RECT 113.300 180.170 113.560 180.260 ;
        RECT 113.820 180.170 113.960 180.620 ;
        RECT 114.220 180.280 114.480 180.600 ;
        RECT 113.300 180.030 113.960 180.170 ;
        RECT 113.300 179.940 113.560 180.030 ;
        RECT 113.360 177.735 113.500 179.940 ;
        RECT 113.290 177.365 113.570 177.735 ;
        RECT 114.280 176.520 114.420 180.280 ;
        RECT 114.740 179.580 114.880 188.100 ;
        RECT 115.140 185.040 115.400 185.360 ;
        RECT 114.680 179.260 114.940 179.580 ;
        RECT 112.440 176.290 113.500 176.430 ;
        RECT 112.840 174.840 113.100 175.160 ;
        RECT 111.920 174.160 112.180 174.480 ;
        RECT 112.370 171.925 112.650 172.295 ;
        RECT 111.920 170.935 112.180 171.080 ;
        RECT 110.990 170.565 111.270 170.935 ;
        RECT 111.910 170.565 112.190 170.935 ;
        RECT 109.620 169.740 109.880 170.060 ;
        RECT 109.160 169.400 109.420 169.720 ;
        RECT 112.440 169.040 112.580 171.925 ;
        RECT 112.900 169.380 113.040 174.840 ;
        RECT 113.360 174.480 113.500 176.290 ;
        RECT 114.220 176.200 114.480 176.520 ;
        RECT 113.300 174.160 113.560 174.480 ;
        RECT 113.760 174.160 114.020 174.480 ;
        RECT 113.300 173.710 113.560 173.800 ;
        RECT 113.820 173.710 113.960 174.160 ;
        RECT 114.220 173.820 114.480 174.140 ;
        RECT 113.300 173.570 113.960 173.710 ;
        RECT 113.300 173.480 113.560 173.570 ;
        RECT 112.840 169.060 113.100 169.380 ;
        RECT 112.380 168.720 112.640 169.040 ;
        RECT 109.160 168.380 109.420 168.700 ;
        RECT 108.690 167.165 108.970 167.535 ;
        RECT 108.760 166.320 108.900 167.165 ;
        RECT 108.700 166.000 108.960 166.320 ;
        RECT 108.230 160.365 108.510 160.735 ;
        RECT 106.860 158.180 107.120 158.500 ;
        RECT 105.940 157.160 106.200 157.480 ;
        RECT 109.220 156.655 109.360 168.380 ;
        RECT 110.080 166.340 110.340 166.660 ;
        RECT 112.380 166.340 112.640 166.660 ;
        RECT 110.140 160.880 110.280 166.340 ;
        RECT 112.440 165.495 112.580 166.340 ;
        RECT 112.370 165.125 112.650 165.495 ;
        RECT 112.840 165.320 113.100 165.640 ;
        RECT 110.540 163.960 110.800 164.280 ;
        RECT 110.600 160.880 110.740 163.960 ;
        RECT 110.080 160.560 110.340 160.880 ;
        RECT 110.540 160.560 110.800 160.880 ;
        RECT 109.150 156.285 109.430 156.655 ;
        RECT 110.080 156.140 110.340 156.460 ;
        RECT 105.020 154.440 105.280 154.760 ;
        RECT 104.100 153.420 104.360 153.740 ;
        RECT 104.160 152.380 104.300 153.420 ;
        RECT 107.320 153.080 107.580 153.400 ;
        RECT 107.380 152.720 107.520 153.080 ;
        RECT 110.140 152.720 110.280 156.140 ;
        RECT 110.600 155.440 110.740 160.560 ;
        RECT 112.900 158.160 113.040 165.320 ;
        RECT 113.360 160.055 113.500 173.480 ;
        RECT 113.760 171.440 114.020 171.760 ;
        RECT 113.820 161.220 113.960 171.440 ;
        RECT 114.280 165.640 114.420 173.820 ;
        RECT 114.220 165.320 114.480 165.640 ;
        RECT 114.220 162.940 114.480 163.260 ;
        RECT 113.760 160.900 114.020 161.220 ;
        RECT 113.290 159.685 113.570 160.055 ;
        RECT 112.840 157.840 113.100 158.160 ;
        RECT 112.840 157.160 113.100 157.480 ;
        RECT 112.900 156.120 113.040 157.160 ;
        RECT 114.280 156.460 114.420 162.940 ;
        RECT 114.740 158.160 114.880 179.260 ;
        RECT 115.200 174.820 115.340 185.040 ;
        RECT 115.660 180.600 115.800 190.480 ;
        RECT 116.580 186.380 116.720 193.540 ;
        RECT 116.970 191.645 117.250 192.015 ;
        RECT 116.520 186.060 116.780 186.380 ;
        RECT 116.060 185.040 116.320 185.360 ;
        RECT 115.600 180.280 115.860 180.600 ;
        RECT 116.120 179.095 116.260 185.040 ;
        RECT 117.040 185.020 117.180 191.645 ;
        RECT 117.900 190.140 118.160 190.460 ;
        RECT 116.980 184.700 117.240 185.020 ;
        RECT 117.440 184.700 117.700 185.020 ;
        RECT 116.510 182.805 116.790 183.175 ;
        RECT 116.520 182.660 116.780 182.805 ;
        RECT 116.980 182.320 117.240 182.640 ;
        RECT 117.040 179.775 117.180 182.320 ;
        RECT 116.970 179.405 117.250 179.775 ;
        RECT 116.050 178.725 116.330 179.095 ;
        RECT 116.520 177.900 116.780 178.220 ;
        RECT 116.580 177.540 116.720 177.900 ;
        RECT 116.520 177.220 116.780 177.540 ;
        RECT 115.600 175.180 115.860 175.500 ;
        RECT 115.140 174.500 115.400 174.820 ;
        RECT 115.660 170.060 115.800 175.180 ;
        RECT 117.500 172.295 117.640 184.700 ;
        RECT 117.960 172.440 118.100 190.140 ;
        RECT 118.820 189.800 119.080 190.120 ;
        RECT 118.880 188.420 119.020 189.800 ;
        RECT 118.820 188.100 119.080 188.420 ;
        RECT 118.880 182.980 119.020 188.100 ;
        RECT 119.340 184.680 119.480 207.020 ;
        RECT 121.110 206.840 121.390 207.340 ;
        RECT 124.330 206.840 124.610 207.340 ;
        RECT 127.550 206.840 127.830 207.340 ;
        RECT 130.770 206.840 131.050 207.340 ;
        RECT 133.540 206.860 133.800 207.120 ;
        RECT 133.990 206.860 134.270 207.340 ;
        RECT 133.540 206.840 134.270 206.860 ;
        RECT 137.210 206.840 137.490 207.340 ;
        RECT 140.430 206.840 140.710 207.340 ;
        RECT 121.180 195.900 121.320 206.840 ;
        RECT 123.410 200.485 123.690 200.855 ;
        RECT 122.030 199.805 122.310 200.175 ;
        RECT 121.120 195.580 121.380 195.900 ;
        RECT 122.100 193.860 122.240 199.805 ;
        RECT 123.480 193.860 123.620 200.485 ;
        RECT 124.400 196.095 124.540 206.840 ;
        RECT 124.330 195.725 124.610 196.095 ;
        RECT 125.260 195.240 125.520 195.560 ;
        RECT 125.720 195.240 125.980 195.560 ;
        RECT 125.320 193.860 125.460 195.240 ;
        RECT 122.040 193.540 122.300 193.860 ;
        RECT 123.420 193.540 123.680 193.860 ;
        RECT 125.260 193.540 125.520 193.860 ;
        RECT 123.880 193.375 124.140 193.520 ;
        RECT 123.870 193.005 124.150 193.375 ;
        RECT 121.120 192.520 121.380 192.840 ;
        RECT 124.340 192.520 124.600 192.840 ;
        RECT 125.260 192.520 125.520 192.840 ;
        RECT 121.180 191.140 121.320 192.520 ;
        RECT 121.120 190.820 121.380 191.140 ;
        RECT 119.730 190.285 120.010 190.655 ;
        RECT 123.880 190.480 124.140 190.800 ;
        RECT 119.280 184.360 119.540 184.680 ;
        RECT 119.800 182.980 119.940 190.285 ;
        RECT 123.420 190.140 123.680 190.460 ;
        RECT 121.580 188.100 121.840 188.420 ;
        RECT 121.640 186.380 121.780 188.100 ;
        RECT 121.580 186.060 121.840 186.380 ;
        RECT 118.820 182.660 119.080 182.980 ;
        RECT 119.740 182.660 120.000 182.980 ;
        RECT 121.120 180.280 121.380 180.600 ;
        RECT 120.660 179.600 120.920 179.920 ;
        RECT 121.180 179.775 121.320 180.280 ;
        RECT 121.640 180.260 121.780 186.060 ;
        RECT 122.960 185.720 123.220 186.040 ;
        RECT 122.490 183.485 122.770 183.855 ;
        RECT 122.560 183.320 122.700 183.485 ;
        RECT 122.500 183.000 122.760 183.320 ;
        RECT 123.020 182.980 123.160 185.720 ;
        RECT 123.480 183.660 123.620 190.140 ;
        RECT 123.420 183.340 123.680 183.660 ;
        RECT 122.960 182.660 123.220 182.980 ;
        RECT 121.580 179.940 121.840 180.260 ;
        RECT 123.020 180.170 123.160 182.660 ;
        RECT 123.020 180.030 123.620 180.170 ;
        RECT 120.200 176.200 120.460 176.520 ;
        RECT 116.060 171.780 116.320 172.100 ;
        RECT 117.430 171.925 117.710 172.295 ;
        RECT 117.900 172.120 118.160 172.440 ;
        RECT 118.820 172.120 119.080 172.440 ;
        RECT 115.600 169.740 115.860 170.060 ;
        RECT 116.120 160.540 116.260 171.780 ;
        RECT 116.520 161.240 116.780 161.560 ;
        RECT 116.060 160.450 116.320 160.540 ;
        RECT 115.200 160.310 116.320 160.450 ;
        RECT 114.680 157.840 114.940 158.160 ;
        RECT 114.220 156.140 114.480 156.460 ;
        RECT 112.840 155.800 113.100 156.120 ;
        RECT 110.540 155.120 110.800 155.440 ;
        RECT 110.600 152.720 110.740 155.120 ;
        RECT 112.900 152.720 113.040 155.800 ;
        RECT 114.220 155.460 114.480 155.780 ;
        RECT 114.280 153.740 114.420 155.460 ;
        RECT 114.680 154.780 114.940 155.100 ;
        RECT 114.220 153.420 114.480 153.740 ;
        RECT 114.740 153.060 114.880 154.780 ;
        RECT 115.200 153.400 115.340 160.310 ;
        RECT 116.060 160.220 116.320 160.310 ;
        RECT 116.580 159.940 116.720 161.240 ;
        RECT 116.120 159.800 116.720 159.940 ;
        RECT 115.600 157.160 115.860 157.480 ;
        RECT 115.140 153.080 115.400 153.400 ;
        RECT 114.680 152.740 114.940 153.060 ;
        RECT 107.320 152.400 107.580 152.720 ;
        RECT 110.080 152.400 110.340 152.720 ;
        RECT 110.540 152.400 110.800 152.720 ;
        RECT 112.840 152.400 113.100 152.720 ;
        RECT 103.640 152.060 103.900 152.380 ;
        RECT 104.100 152.060 104.360 152.380 ;
        RECT 115.660 152.040 115.800 157.160 ;
        RECT 116.120 154.760 116.260 159.800 ;
        RECT 117.440 157.500 117.700 157.820 ;
        RECT 116.060 154.440 116.320 154.760 ;
        RECT 116.520 154.440 116.780 154.760 ;
        RECT 116.580 152.970 116.720 154.440 ;
        RECT 117.500 153.060 117.640 157.500 ;
        RECT 117.960 156.120 118.100 172.120 ;
        RECT 118.880 167.000 119.020 172.120 ;
        RECT 118.820 166.680 119.080 167.000 ;
        RECT 118.880 159.180 119.020 166.680 ;
        RECT 120.260 160.450 120.400 176.200 ;
        RECT 120.720 170.060 120.860 179.600 ;
        RECT 121.110 179.405 121.390 179.775 ;
        RECT 121.180 177.450 121.320 179.405 ;
        RECT 121.640 178.220 121.780 179.940 ;
        RECT 122.960 179.260 123.220 179.580 ;
        RECT 121.580 177.900 121.840 178.220 ;
        RECT 121.580 177.450 121.840 177.540 ;
        RECT 122.500 177.450 122.760 177.540 ;
        RECT 121.180 177.310 121.840 177.450 ;
        RECT 121.580 177.220 121.840 177.310 ;
        RECT 122.100 177.310 122.760 177.450 ;
        RECT 121.580 176.200 121.840 176.520 ;
        RECT 121.640 173.800 121.780 176.200 ;
        RECT 121.580 173.480 121.840 173.800 ;
        RECT 122.100 173.655 122.240 177.310 ;
        RECT 122.500 177.220 122.760 177.310 ;
        RECT 122.490 173.965 122.770 174.335 ;
        RECT 122.030 173.285 122.310 173.655 ;
        RECT 120.660 169.740 120.920 170.060 ;
        RECT 120.720 163.600 120.860 169.740 ;
        RECT 121.120 169.060 121.380 169.380 ;
        RECT 120.660 163.280 120.920 163.600 ;
        RECT 121.180 160.880 121.320 169.060 ;
        RECT 122.100 167.420 122.240 173.285 ;
        RECT 121.640 167.280 122.240 167.420 ;
        RECT 121.640 166.320 121.780 167.280 ;
        RECT 122.040 166.680 122.300 167.000 ;
        RECT 121.580 166.000 121.840 166.320 ;
        RECT 121.580 164.300 121.840 164.620 ;
        RECT 121.120 160.560 121.380 160.880 ;
        RECT 120.660 160.450 120.920 160.540 ;
        RECT 120.260 160.310 120.920 160.450 ;
        RECT 120.660 160.220 120.920 160.310 ;
        RECT 119.280 159.880 119.540 160.200 ;
        RECT 118.360 158.860 118.620 159.180 ;
        RECT 118.820 158.860 119.080 159.180 ;
        RECT 118.420 158.500 118.560 158.860 ;
        RECT 118.360 158.180 118.620 158.500 ;
        RECT 117.900 155.800 118.160 156.120 ;
        RECT 116.120 152.830 116.720 152.970 ;
        RECT 115.600 151.720 115.860 152.040 ;
        RECT 101.800 150.700 102.060 151.020 ;
        RECT 101.340 149.340 101.600 149.660 ;
        RECT 116.120 149.320 116.260 152.830 ;
        RECT 117.440 152.740 117.700 153.060 ;
        RECT 117.900 152.740 118.160 153.060 ;
        RECT 116.520 152.060 116.780 152.380 ;
        RECT 116.580 150.340 116.720 152.060 ;
        RECT 116.520 150.020 116.780 150.340 ;
        RECT 116.060 149.000 116.320 149.320 ;
        RECT 95.360 148.320 95.620 148.640 ;
        RECT 111.460 146.960 111.720 147.280 ;
        RECT 105.020 146.620 105.280 146.940 ;
        RECT 98.580 146.280 98.840 146.600 ;
        RECT 95.360 145.260 95.620 145.580 ;
        RECT 95.420 140.990 95.560 145.260 ;
        RECT 98.640 140.990 98.780 146.280 ;
        RECT 101.800 145.600 102.060 145.920 ;
        RECT 101.860 140.990 102.000 145.600 ;
        RECT 105.080 140.990 105.220 146.620 ;
        RECT 108.240 145.940 108.500 146.260 ;
        RECT 108.300 140.990 108.440 145.940 ;
        RECT 111.520 140.990 111.660 146.960 ;
        RECT 114.680 140.990 114.940 141.160 ;
        RECT 117.960 140.990 118.100 152.740 ;
        RECT 119.340 152.720 119.480 159.880 ;
        RECT 120.720 157.480 120.860 160.220 ;
        RECT 120.660 157.160 120.920 157.480 ;
        RECT 121.180 155.780 121.320 160.560 ;
        RECT 121.640 157.480 121.780 164.300 ;
        RECT 122.100 160.880 122.240 166.680 ;
        RECT 122.040 160.560 122.300 160.880 ;
        RECT 122.560 159.180 122.700 173.965 ;
        RECT 123.020 172.100 123.160 179.260 ;
        RECT 123.480 179.240 123.620 180.030 ;
        RECT 123.420 178.920 123.680 179.240 ;
        RECT 123.480 177.880 123.620 178.920 ;
        RECT 123.420 177.560 123.680 177.880 ;
        RECT 123.940 176.520 124.080 190.480 ;
        RECT 124.400 190.370 124.540 192.520 ;
        RECT 124.800 190.370 125.060 190.460 ;
        RECT 124.400 190.230 125.060 190.370 ;
        RECT 124.400 188.080 124.540 190.230 ;
        RECT 124.800 190.140 125.060 190.230 ;
        RECT 124.340 187.760 124.600 188.080 ;
        RECT 124.800 184.360 125.060 184.680 ;
        RECT 124.860 183.660 125.000 184.360 ;
        RECT 124.800 183.340 125.060 183.660 ;
        RECT 124.340 183.000 124.600 183.320 ;
        RECT 124.400 182.495 124.540 183.000 ;
        RECT 124.330 182.125 124.610 182.495 ;
        RECT 123.880 176.200 124.140 176.520 ;
        RECT 123.420 174.160 123.680 174.480 ;
        RECT 122.960 171.780 123.220 172.100 ;
        RECT 123.480 167.340 123.620 174.160 ;
        RECT 123.880 173.820 124.140 174.140 ;
        RECT 123.420 167.020 123.680 167.340 ;
        RECT 123.940 166.660 124.080 173.820 ;
        RECT 124.400 166.660 124.540 182.125 ;
        RECT 125.320 177.540 125.460 192.520 ;
        RECT 125.780 191.820 125.920 195.240 ;
        RECT 127.100 193.540 127.360 193.860 ;
        RECT 127.160 192.695 127.300 193.540 ;
        RECT 127.090 192.325 127.370 192.695 ;
        RECT 127.620 191.820 127.760 206.840 ;
        RECT 130.310 194.365 130.590 194.735 ;
        RECT 130.380 194.200 130.520 194.365 ;
        RECT 129.850 193.685 130.130 194.055 ;
        RECT 130.320 193.880 130.580 194.200 ;
        RECT 129.860 193.540 130.120 193.685 ;
        RECT 129.860 192.860 130.120 193.180 ;
        RECT 128.480 192.520 128.740 192.840 ;
        RECT 125.720 191.500 125.980 191.820 ;
        RECT 127.560 191.500 127.820 191.820 ;
        RECT 126.640 187.080 126.900 187.400 ;
        RECT 127.100 187.080 127.360 187.400 ;
        RECT 126.180 183.000 126.440 183.320 ;
        RECT 125.720 182.660 125.980 182.980 ;
        RECT 125.780 178.220 125.920 182.660 ;
        RECT 126.240 181.135 126.380 183.000 ;
        RECT 126.700 182.980 126.840 187.080 ;
        RECT 126.640 182.660 126.900 182.980 ;
        RECT 126.170 180.765 126.450 181.135 ;
        RECT 125.720 177.900 125.980 178.220 ;
        RECT 125.260 177.220 125.520 177.540 ;
        RECT 125.260 176.540 125.520 176.860 ;
        RECT 124.800 171.780 125.060 172.100 ;
        RECT 123.880 166.340 124.140 166.660 ;
        RECT 124.340 166.340 124.600 166.660 ;
        RECT 124.860 164.620 125.000 171.780 ;
        RECT 125.320 169.040 125.460 176.540 ;
        RECT 126.240 171.760 126.380 180.765 ;
        RECT 127.160 174.220 127.300 187.080 ;
        RECT 128.540 185.360 128.680 192.520 ;
        RECT 129.400 187.420 129.660 187.740 ;
        RECT 127.560 185.270 127.820 185.360 ;
        RECT 127.560 185.130 128.220 185.270 ;
        RECT 128.480 185.215 128.740 185.360 ;
        RECT 127.560 185.040 127.820 185.130 ;
        RECT 127.550 182.805 127.830 183.175 ;
        RECT 127.560 182.660 127.820 182.805 ;
        RECT 127.550 175.325 127.830 175.695 ;
        RECT 126.700 174.080 127.300 174.220 ;
        RECT 125.720 171.440 125.980 171.760 ;
        RECT 126.180 171.440 126.440 171.760 ;
        RECT 125.780 169.040 125.920 171.440 ;
        RECT 126.180 170.760 126.440 171.080 ;
        RECT 126.240 169.720 126.380 170.760 ;
        RECT 126.180 169.400 126.440 169.720 ;
        RECT 125.260 168.720 125.520 169.040 ;
        RECT 125.720 168.720 125.980 169.040 ;
        RECT 126.180 167.020 126.440 167.340 ;
        RECT 126.240 166.855 126.380 167.020 ;
        RECT 126.170 166.485 126.450 166.855 ;
        RECT 126.180 166.340 126.440 166.485 ;
        RECT 126.700 166.320 126.840 174.080 ;
        RECT 127.100 173.480 127.360 173.800 ;
        RECT 127.160 172.440 127.300 173.480 ;
        RECT 127.620 172.440 127.760 175.325 ;
        RECT 127.100 172.120 127.360 172.440 ;
        RECT 127.560 172.120 127.820 172.440 ;
        RECT 127.160 166.660 127.300 172.120 ;
        RECT 127.560 171.440 127.820 171.760 ;
        RECT 127.100 166.340 127.360 166.660 ;
        RECT 126.640 166.000 126.900 166.320 ;
        RECT 124.800 164.300 125.060 164.620 ;
        RECT 124.860 161.900 125.000 164.300 ;
        RECT 124.800 161.580 125.060 161.900 ;
        RECT 123.880 160.900 124.140 161.220 ;
        RECT 124.800 160.900 125.060 161.220 ;
        RECT 122.500 158.860 122.760 159.180 ;
        RECT 123.940 158.500 124.080 160.900 ;
        RECT 123.880 158.180 124.140 158.500 ;
        RECT 124.860 158.160 125.000 160.900 ;
        RECT 124.800 157.840 125.060 158.160 ;
        RECT 121.580 157.160 121.840 157.480 ;
        RECT 121.120 155.460 121.380 155.780 ;
        RECT 119.280 152.400 119.540 152.720 ;
        RECT 126.700 152.380 126.840 166.000 ;
        RECT 127.620 165.640 127.760 171.440 ;
        RECT 128.080 165.980 128.220 185.130 ;
        RECT 128.470 184.845 128.750 185.215 ;
        RECT 128.940 184.700 129.200 185.020 ;
        RECT 128.480 177.220 128.740 177.540 ;
        RECT 128.540 175.500 128.680 177.220 ;
        RECT 128.480 175.180 128.740 175.500 ;
        RECT 129.000 174.140 129.140 184.700 ;
        RECT 129.460 182.980 129.600 187.420 ;
        RECT 129.920 185.700 130.060 192.860 ;
        RECT 130.320 189.800 130.580 190.120 ;
        RECT 129.860 185.380 130.120 185.700 ;
        RECT 130.380 185.360 130.520 189.800 ;
        RECT 130.840 188.860 130.980 206.840 ;
        RECT 133.540 206.800 134.200 206.840 ;
        RECT 133.600 206.720 134.200 206.800 ;
        RECT 131.240 195.240 131.500 195.560 ;
        RECT 131.300 193.180 131.440 195.240 ;
        RECT 131.700 193.880 131.960 194.200 ;
        RECT 133.540 193.880 133.800 194.200 ;
        RECT 131.240 192.860 131.500 193.180 ;
        RECT 131.300 190.800 131.440 192.860 ;
        RECT 131.240 190.480 131.500 190.800 ;
        RECT 130.840 188.720 131.440 188.860 ;
        RECT 130.780 188.100 131.040 188.420 ;
        RECT 130.320 185.040 130.580 185.360 ;
        RECT 129.400 182.660 129.660 182.980 ;
        RECT 129.400 180.620 129.660 180.940 ;
        RECT 129.460 177.880 129.600 180.620 ;
        RECT 129.400 177.560 129.660 177.880 ;
        RECT 128.940 173.820 129.200 174.140 ;
        RECT 128.940 171.780 129.200 172.100 ;
        RECT 128.480 170.760 128.740 171.080 ;
        RECT 128.020 165.660 128.280 165.980 ;
        RECT 127.560 165.320 127.820 165.640 ;
        RECT 127.100 158.860 127.360 159.180 ;
        RECT 127.160 156.120 127.300 158.860 ;
        RECT 128.080 156.460 128.220 165.660 ;
        RECT 128.020 156.140 128.280 156.460 ;
        RECT 127.100 155.800 127.360 156.120 ;
        RECT 128.540 155.440 128.680 170.760 ;
        RECT 129.000 160.880 129.140 171.780 ;
        RECT 129.460 163.940 129.600 177.560 ;
        RECT 129.860 177.220 130.120 177.540 ;
        RECT 129.920 177.055 130.060 177.220 ;
        RECT 129.850 176.685 130.130 177.055 ;
        RECT 129.860 176.200 130.120 176.520 ;
        RECT 129.920 165.640 130.060 176.200 ;
        RECT 130.840 175.060 130.980 188.100 ;
        RECT 131.300 187.400 131.440 188.720 ;
        RECT 131.240 187.080 131.500 187.400 ;
        RECT 131.760 185.360 131.900 193.880 ;
        RECT 132.160 192.520 132.420 192.840 ;
        RECT 132.620 192.520 132.880 192.840 ;
        RECT 132.220 189.295 132.360 192.520 ;
        RECT 132.150 188.925 132.430 189.295 ;
        RECT 131.700 185.040 131.960 185.360 ;
        RECT 132.160 184.360 132.420 184.680 ;
        RECT 132.220 182.980 132.360 184.360 ;
        RECT 132.160 182.660 132.420 182.980 ;
        RECT 132.680 182.495 132.820 192.520 ;
        RECT 133.600 190.800 133.740 193.880 ;
        RECT 133.540 190.480 133.800 190.800 ;
        RECT 133.080 188.100 133.340 188.420 ;
        RECT 132.610 182.125 132.890 182.495 ;
        RECT 133.140 180.940 133.280 188.100 ;
        RECT 133.600 186.575 133.740 190.480 ;
        RECT 134.000 189.800 134.260 190.120 ;
        RECT 133.530 186.205 133.810 186.575 ;
        RECT 134.060 183.660 134.200 189.800 ;
        RECT 134.920 187.420 135.180 187.740 ;
        RECT 134.000 183.340 134.260 183.660 ;
        RECT 133.080 180.620 133.340 180.940 ;
        RECT 131.240 178.920 131.500 179.240 ;
        RECT 131.300 177.540 131.440 178.920 ;
        RECT 132.160 177.560 132.420 177.880 ;
        RECT 131.240 177.220 131.500 177.540 ;
        RECT 130.380 174.920 130.980 175.060 ;
        RECT 130.380 167.340 130.520 174.920 ;
        RECT 130.780 173.820 131.040 174.140 ;
        RECT 130.320 167.020 130.580 167.340 ;
        RECT 129.860 165.320 130.120 165.640 ;
        RECT 129.400 163.620 129.660 163.940 ;
        RECT 129.460 161.560 129.600 163.620 ;
        RECT 129.920 161.560 130.060 165.320 ;
        RECT 129.400 161.240 129.660 161.560 ;
        RECT 129.860 161.240 130.120 161.560 ;
        RECT 128.940 160.560 129.200 160.880 ;
        RECT 129.400 160.220 129.660 160.540 ;
        RECT 128.480 155.120 128.740 155.440 ;
        RECT 126.180 152.060 126.440 152.380 ;
        RECT 126.640 152.060 126.900 152.380 ;
        RECT 126.240 151.215 126.380 152.060 ;
        RECT 129.460 152.040 129.600 160.220 ;
        RECT 129.850 156.285 130.130 156.655 ;
        RECT 129.920 155.780 130.060 156.285 ;
        RECT 129.860 155.460 130.120 155.780 ;
        RECT 129.920 153.060 130.060 155.460 ;
        RECT 130.380 153.060 130.520 167.020 ;
        RECT 130.840 163.600 130.980 173.820 ;
        RECT 131.300 171.420 131.440 177.220 ;
        RECT 132.220 174.390 132.360 177.560 ;
        RECT 132.620 177.220 132.880 177.540 ;
        RECT 132.680 175.060 132.820 177.220 ;
        RECT 134.460 176.540 134.720 176.860 ;
        RECT 132.680 174.920 133.280 175.060 ;
        RECT 132.220 174.250 132.820 174.390 ;
        RECT 131.690 171.925 131.970 172.295 ;
        RECT 131.700 171.780 131.960 171.925 ;
        RECT 131.240 171.100 131.500 171.420 ;
        RECT 132.680 169.575 132.820 174.250 ;
        RECT 133.140 172.975 133.280 174.920 ;
        RECT 133.070 172.860 133.350 172.975 ;
        RECT 133.070 172.720 133.740 172.860 ;
        RECT 133.070 172.605 133.350 172.720 ;
        RECT 133.080 171.780 133.340 172.100 ;
        RECT 132.610 169.205 132.890 169.575 ;
        RECT 132.680 166.660 132.820 169.205 ;
        RECT 133.140 167.340 133.280 171.780 ;
        RECT 133.080 167.020 133.340 167.340 ;
        RECT 133.600 166.660 133.740 172.720 ;
        RECT 134.000 170.760 134.260 171.080 ;
        RECT 134.060 169.720 134.200 170.760 ;
        RECT 134.000 169.400 134.260 169.720 ;
        RECT 132.620 166.340 132.880 166.660 ;
        RECT 133.080 166.340 133.340 166.660 ;
        RECT 133.540 166.340 133.800 166.660 ;
        RECT 131.240 165.320 131.500 165.640 ;
        RECT 130.780 163.280 131.040 163.600 ;
        RECT 131.300 161.220 131.440 165.320 ;
        RECT 131.240 160.900 131.500 161.220 ;
        RECT 132.160 160.900 132.420 161.220 ;
        RECT 132.220 156.460 132.360 160.900 ;
        RECT 133.140 156.460 133.280 166.340 ;
        RECT 133.540 163.280 133.800 163.600 ;
        RECT 133.600 158.160 133.740 163.280 ;
        RECT 134.000 162.600 134.260 162.920 ;
        RECT 133.540 157.840 133.800 158.160 ;
        RECT 132.160 156.140 132.420 156.460 ;
        RECT 133.080 156.140 133.340 156.460 ;
        RECT 132.150 153.565 132.430 153.935 ;
        RECT 129.860 152.740 130.120 153.060 ;
        RECT 130.320 152.740 130.580 153.060 ;
        RECT 132.220 152.720 132.360 153.565 ;
        RECT 132.620 153.255 132.880 153.400 ;
        RECT 132.610 152.885 132.890 153.255 ;
        RECT 132.160 152.400 132.420 152.720 ;
        RECT 129.400 151.720 129.660 152.040 ;
        RECT 126.170 150.845 126.450 151.215 ;
        RECT 134.060 144.415 134.200 162.600 ;
        RECT 134.520 153.740 134.660 176.540 ;
        RECT 134.980 156.120 135.120 187.420 ;
        RECT 137.280 186.380 137.420 206.840 ;
        RECT 139.050 205.245 139.330 205.615 ;
        RECT 137.220 186.060 137.480 186.380 ;
        RECT 139.120 182.980 139.260 205.245 ;
        RECT 140.500 188.760 140.640 206.840 ;
        RECT 140.440 188.440 140.700 188.760 ;
        RECT 139.060 182.660 139.320 182.980 ;
        RECT 139.970 181.445 140.250 181.815 ;
        RECT 140.040 175.160 140.180 181.445 ;
        RECT 139.980 174.840 140.240 175.160 ;
        RECT 134.920 155.800 135.180 156.120 ;
        RECT 134.460 153.420 134.720 153.740 ;
        RECT 133.990 144.045 134.270 144.415 ;
        RECT 127.560 143.560 127.820 143.880 ;
        RECT 127.620 140.990 127.760 143.560 ;
        RECT 88.910 140.490 89.190 140.990 ;
        RECT 92.130 140.490 92.410 140.990 ;
        RECT 95.350 140.490 95.630 140.990 ;
        RECT 98.570 140.490 98.850 140.990 ;
        RECT 101.790 140.490 102.070 140.990 ;
        RECT 105.010 140.490 105.290 140.990 ;
        RECT 108.230 140.490 108.510 140.990 ;
        RECT 111.450 140.490 111.730 140.990 ;
        RECT 114.670 140.490 114.950 140.990 ;
        RECT 117.890 140.490 118.170 140.990 ;
        RECT 127.550 140.490 127.830 140.990 ;
        RECT 53.325 59.470 64.870 60.060 ;
        RECT 111.750 59.945 112.295 61.945 ;
        RECT 69.915 59.895 70.565 59.915 ;
        RECT 69.915 59.350 81.855 59.895 ;
        RECT 69.915 59.280 70.565 59.350 ;
        RECT 86.775 59.345 98.425 59.890 ;
        RECT 103.345 59.400 112.295 59.945 ;
        RECT 55.995 58.715 56.590 59.155 ;
        RECT 48.675 58.120 56.590 58.715 ;
        RECT 61.655 58.415 73.225 59.005 ;
        RECT 78.395 58.205 90.005 58.795 ;
        RECT 95.040 58.200 106.720 58.745 ;
        RECT 1.590 48.345 2.085 50.885 ;
        RECT 10.550 48.800 10.995 50.625 ;
        RECT 10.295 48.355 11.245 48.800 ;
        RECT 13.120 48.430 13.900 57.440 ;
        RECT 1.560 47.850 2.115 48.345 ;
        RECT 14.520 46.920 14.795 46.950 ;
        RECT 12.590 46.645 14.795 46.920 ;
        RECT 12.590 44.305 12.865 46.645 ;
        RECT 14.520 46.615 14.795 46.645 ;
        RECT 3.045 40.875 3.365 40.930 ;
        RECT 8.925 40.875 9.245 40.930 ;
        RECT 3.045 40.725 9.245 40.875 ;
        RECT 3.045 40.670 3.365 40.725 ;
        RECT 8.925 40.670 9.245 40.725 ;
        RECT 1.890 39.095 7.495 39.425 ;
        RECT 1.890 23.395 2.220 39.095 ;
        RECT 3.840 37.265 4.160 37.290 ;
        RECT 20.960 37.265 21.280 37.290 ;
        RECT 3.840 37.055 21.280 37.265 ;
        RECT 3.840 37.030 4.160 37.055 ;
        RECT 20.960 37.030 21.280 37.055 ;
        RECT 11.295 36.260 15.800 36.555 ;
        RECT 25.745 32.720 26.120 51.710 ;
        RECT 10.295 32.345 26.120 32.720 ;
        RECT 14.520 30.920 14.795 30.950 ;
        RECT 12.590 30.645 14.795 30.920 ;
        RECT 12.590 28.305 12.865 30.645 ;
        RECT 14.520 30.615 14.795 30.645 ;
        RECT 3.045 24.875 3.365 24.930 ;
        RECT 8.925 24.875 9.245 24.930 ;
        RECT 3.045 24.725 9.245 24.875 ;
        RECT 3.045 24.670 3.365 24.725 ;
        RECT 8.925 24.670 9.245 24.725 ;
        RECT 1.890 23.065 7.525 23.395 ;
        RECT 1.900 7.445 2.230 23.065 ;
        RECT 3.840 21.265 4.160 21.290 ;
        RECT 20.960 21.265 21.280 21.290 ;
        RECT 3.840 21.055 21.280 21.265 ;
        RECT 3.840 21.030 4.160 21.055 ;
        RECT 20.960 21.030 21.280 21.055 ;
        RECT 11.295 20.260 15.800 20.555 ;
        RECT 26.595 16.035 27.000 50.605 ;
        RECT 27.990 39.880 28.240 53.505 ;
        RECT 27.990 39.795 28.490 39.880 ;
        RECT 27.585 39.535 28.490 39.795 ;
        RECT 28.190 39.480 28.490 39.535 ;
        RECT 28.715 39.050 29.060 53.450 ;
        RECT 27.945 38.705 29.060 39.050 ;
        RECT 27.945 23.795 28.290 38.705 ;
        RECT 29.650 38.120 29.930 53.420 ;
        RECT 38.585 48.715 38.960 50.660 ;
        RECT 38.295 48.340 39.245 48.715 ;
        RECT 42.520 46.920 42.795 46.950 ;
        RECT 40.590 46.645 42.795 46.920 ;
        RECT 40.590 44.305 40.865 46.645 ;
        RECT 42.520 46.615 42.795 46.645 ;
        RECT 31.045 40.875 31.365 40.930 ;
        RECT 36.925 40.875 37.245 40.930 ;
        RECT 31.045 40.725 37.245 40.875 ;
        RECT 31.045 40.670 31.365 40.725 ;
        RECT 36.925 40.670 37.245 40.725 ;
        RECT 28.850 37.840 29.930 38.120 ;
        RECT 30.390 39.370 35.500 39.720 ;
        RECT 27.585 23.450 28.645 23.795 ;
        RECT 28.850 23.220 29.130 37.840 ;
        RECT 10.295 15.630 27.000 16.035 ;
        RECT 27.975 22.940 29.130 23.220 ;
        RECT 30.390 23.385 30.740 39.370 ;
        RECT 31.840 37.265 32.160 37.290 ;
        RECT 48.960 37.265 49.280 37.290 ;
        RECT 31.840 37.055 49.280 37.265 ;
        RECT 31.840 37.030 32.160 37.055 ;
        RECT 48.960 37.030 49.280 37.055 ;
        RECT 39.295 36.260 43.800 36.555 ;
        RECT 53.810 32.600 54.210 51.745 ;
        RECT 38.295 32.200 54.210 32.600 ;
        RECT 42.520 30.920 42.795 30.950 ;
        RECT 40.590 30.645 42.795 30.920 ;
        RECT 40.590 28.305 40.865 30.645 ;
        RECT 42.520 30.615 42.795 30.645 ;
        RECT 31.045 24.875 31.365 24.930 ;
        RECT 36.925 24.875 37.245 24.930 ;
        RECT 31.045 24.725 37.245 24.875 ;
        RECT 31.045 24.670 31.365 24.725 ;
        RECT 36.925 24.670 37.245 24.725 ;
        RECT 30.390 23.035 35.495 23.385 ;
        RECT 14.520 14.920 14.795 14.950 ;
        RECT 12.590 14.645 14.795 14.920 ;
        RECT 12.590 12.305 12.865 14.645 ;
        RECT 14.520 14.615 14.795 14.645 ;
        RECT 3.045 8.875 3.365 8.930 ;
        RECT 8.925 8.875 9.245 8.930 ;
        RECT 3.045 8.725 9.245 8.875 ;
        RECT 3.045 8.670 3.365 8.725 ;
        RECT 8.925 8.670 9.245 8.725 ;
        RECT 27.975 7.795 28.255 22.940 ;
        RECT 27.585 7.515 28.645 7.795 ;
        RECT 1.900 7.115 7.750 7.445 ;
        RECT 30.390 7.420 30.740 23.035 ;
        RECT 31.840 21.265 32.160 21.290 ;
        RECT 48.960 21.265 49.280 21.290 ;
        RECT 31.840 21.055 49.280 21.265 ;
        RECT 31.840 21.030 32.160 21.055 ;
        RECT 48.960 21.030 49.280 21.055 ;
        RECT 39.295 20.260 43.800 20.555 ;
        RECT 54.695 16.730 55.100 50.710 ;
        RECT 55.615 38.765 55.890 53.615 ;
        RECT 56.365 38.100 56.610 53.600 ;
        RECT 55.625 37.855 56.610 38.100 ;
        RECT 55.625 23.825 55.870 37.855 ;
        RECT 57.025 37.140 57.350 53.540 ;
        RECT 66.595 48.470 66.945 50.685 ;
        RECT 79.480 50.170 80.050 50.690 ;
        RECT 68.565 48.855 70.130 49.935 ;
        RECT 66.295 48.120 67.245 48.470 ;
        RECT 70.520 46.920 70.795 46.950 ;
        RECT 68.590 46.645 70.795 46.920 ;
        RECT 68.590 44.305 68.865 46.645 ;
        RECT 70.520 46.615 70.795 46.645 ;
        RECT 59.045 40.875 59.365 40.930 ;
        RECT 64.925 40.875 65.245 40.930 ;
        RECT 59.045 40.725 65.245 40.875 ;
        RECT 59.045 40.670 59.365 40.725 ;
        RECT 64.925 40.670 65.245 40.725 ;
        RECT 56.290 36.815 57.350 37.140 ;
        RECT 57.605 39.260 63.490 39.605 ;
        RECT 55.615 22.765 55.875 23.825 ;
        RECT 38.295 16.325 55.100 16.730 ;
        RECT 42.520 14.920 42.795 14.950 ;
        RECT 40.590 14.645 42.795 14.920 ;
        RECT 40.590 12.305 40.865 14.645 ;
        RECT 42.520 14.615 42.795 14.645 ;
        RECT 31.045 8.875 31.365 8.930 ;
        RECT 36.925 8.875 37.245 8.930 ;
        RECT 31.045 8.725 37.245 8.875 ;
        RECT 31.045 8.670 31.365 8.725 ;
        RECT 36.925 8.670 37.245 8.725 ;
        RECT 35.680 7.445 35.960 7.465 ;
        RECT 35.205 7.420 35.985 7.445 ;
        RECT 30.390 7.115 35.985 7.420 ;
        RECT 30.390 7.095 35.960 7.115 ;
        RECT 30.390 7.070 35.805 7.095 ;
        RECT 35.365 7.065 35.805 7.070 ;
        RECT 56.290 6.765 56.615 36.815 ;
        RECT 57.605 23.425 57.950 39.260 ;
        RECT 59.840 37.265 60.160 37.290 ;
        RECT 76.960 37.265 77.280 37.290 ;
        RECT 59.840 37.055 77.280 37.265 ;
        RECT 59.840 37.030 60.160 37.055 ;
        RECT 76.960 37.030 77.280 37.055 ;
        RECT 67.295 36.260 71.800 36.555 ;
        RECT 79.805 34.570 81.180 36.025 ;
        RECT 68.645 33.350 69.995 34.205 ;
        RECT 68.690 33.320 69.950 33.350 ;
        RECT 81.780 32.540 82.120 50.765 ;
        RECT 82.740 37.785 83.135 50.785 ;
        RECT 83.635 39.825 83.855 53.395 ;
        RECT 83.615 38.765 83.875 39.825 ;
        RECT 82.740 37.390 83.865 37.785 ;
        RECT 66.295 32.200 82.120 32.540 ;
        RECT 70.520 30.920 70.795 30.950 ;
        RECT 68.590 30.645 70.795 30.920 ;
        RECT 68.590 28.305 68.865 30.645 ;
        RECT 70.520 30.615 70.795 30.645 ;
        RECT 59.045 24.875 59.365 24.930 ;
        RECT 64.925 24.875 65.245 24.930 ;
        RECT 59.045 24.725 65.245 24.875 ;
        RECT 59.045 24.670 59.365 24.725 ;
        RECT 64.925 24.670 65.245 24.725 ;
        RECT 57.605 23.080 63.540 23.425 ;
        RECT 57.625 7.465 57.970 23.080 ;
        RECT 59.840 21.265 60.160 21.290 ;
        RECT 76.960 21.265 77.280 21.290 ;
        RECT 59.840 21.055 77.280 21.265 ;
        RECT 59.840 21.030 60.160 21.055 ;
        RECT 76.960 21.030 77.280 21.055 ;
        RECT 67.295 20.260 71.800 20.555 ;
        RECT 80.460 18.535 81.835 19.990 ;
        RECT 68.745 16.870 69.890 18.105 ;
        RECT 83.470 16.550 83.865 37.390 ;
        RECT 84.315 22.765 84.615 53.320 ;
        RECT 85.115 52.855 85.480 53.355 ;
        RECT 85.110 22.360 85.480 52.855 ;
        RECT 85.895 47.895 86.200 53.345 ;
        RECT 86.535 48.445 86.860 53.330 ;
        RECT 87.210 49.015 87.515 53.345 ;
        RECT 87.860 49.660 88.205 53.340 ;
        RECT 88.565 50.245 88.915 53.325 ;
        RECT 89.320 51.020 89.710 53.215 ;
        RECT 89.320 50.630 141.315 51.020 ;
        RECT 88.565 49.895 140.615 50.245 ;
        RECT 87.860 49.315 139.960 49.660 ;
        RECT 87.210 48.710 113.130 49.015 ;
        RECT 86.535 48.120 112.540 48.445 ;
        RECT 85.895 47.620 111.920 47.895 ;
        RECT 85.895 47.590 107.810 47.620 ;
        RECT 108.860 47.590 111.920 47.620 ;
        RECT 98.520 46.920 98.795 46.950 ;
        RECT 94.475 46.100 95.240 46.800 ;
        RECT 96.590 46.645 98.795 46.920 ;
        RECT 96.590 44.305 96.865 46.645 ;
        RECT 98.520 46.615 98.795 46.645 ;
        RECT 87.045 40.875 87.365 40.930 ;
        RECT 92.925 40.875 93.245 40.930 ;
        RECT 87.045 40.725 93.245 40.875 ;
        RECT 87.045 40.670 87.365 40.725 ;
        RECT 92.925 40.670 93.245 40.725 ;
        RECT 85.980 39.200 91.525 39.600 ;
        RECT 66.295 16.155 83.865 16.550 ;
        RECT 84.245 21.990 85.480 22.360 ;
        RECT 86.010 23.410 86.410 39.200 ;
        RECT 111.615 38.765 111.920 47.590 ;
        RECT 112.215 37.960 112.540 48.120 ;
        RECT 111.615 37.635 112.540 37.960 ;
        RECT 87.840 37.265 88.160 37.290 ;
        RECT 104.960 37.265 105.280 37.290 ;
        RECT 87.840 37.055 105.280 37.265 ;
        RECT 87.840 37.030 88.160 37.055 ;
        RECT 104.960 37.030 105.280 37.055 ;
        RECT 95.295 36.260 99.800 36.555 ;
        RECT 94.605 31.765 95.370 32.465 ;
        RECT 98.520 30.920 98.795 30.950 ;
        RECT 96.590 30.645 98.795 30.920 ;
        RECT 96.590 28.305 96.865 30.645 ;
        RECT 98.520 30.615 98.795 30.645 ;
        RECT 87.045 24.875 87.365 24.930 ;
        RECT 92.925 24.875 93.245 24.930 ;
        RECT 87.045 24.725 93.245 24.875 ;
        RECT 87.045 24.670 87.365 24.725 ;
        RECT 92.925 24.670 93.245 24.725 ;
        RECT 86.010 23.010 91.555 23.410 ;
        RECT 70.520 14.920 70.795 14.950 ;
        RECT 68.590 14.645 70.795 14.920 ;
        RECT 68.590 12.305 68.865 14.645 ;
        RECT 70.520 14.615 70.795 14.645 ;
        RECT 59.045 8.875 59.365 8.930 ;
        RECT 64.925 8.875 65.245 8.930 ;
        RECT 59.045 8.725 65.245 8.875 ;
        RECT 59.045 8.670 59.365 8.725 ;
        RECT 64.925 8.670 65.245 8.725 ;
        RECT 57.625 7.120 63.500 7.465 ;
        RECT 58.505 7.115 59.265 7.120 ;
        RECT 58.530 7.095 58.810 7.115 ;
        RECT 84.245 6.765 84.615 21.990 ;
        RECT 86.010 7.405 86.410 23.010 ;
        RECT 111.615 22.765 111.940 37.635 ;
        RECT 112.825 37.195 113.130 48.710 ;
        RECT 126.520 46.920 126.795 46.950 ;
        RECT 124.590 46.645 126.795 46.920 ;
        RECT 124.590 44.305 124.865 46.645 ;
        RECT 126.520 46.615 126.795 46.645 ;
        RECT 122.420 43.515 123.095 44.300 ;
        RECT 115.045 40.875 115.365 40.930 ;
        RECT 120.925 40.875 121.245 40.930 ;
        RECT 115.045 40.725 121.245 40.875 ;
        RECT 115.045 40.670 115.365 40.725 ;
        RECT 120.925 40.670 121.245 40.725 ;
        RECT 112.255 36.890 113.130 37.195 ;
        RECT 114.105 39.165 119.460 39.450 ;
        RECT 87.840 21.265 88.160 21.290 ;
        RECT 104.960 21.265 105.280 21.290 ;
        RECT 87.840 21.055 105.280 21.265 ;
        RECT 87.840 21.030 88.160 21.055 ;
        RECT 104.960 21.030 105.280 21.055 ;
        RECT 95.295 20.260 99.800 20.555 ;
        RECT 94.375 15.590 95.140 16.290 ;
        RECT 98.520 14.920 98.795 14.950 ;
        RECT 96.590 14.645 98.795 14.920 ;
        RECT 96.590 12.305 96.865 14.645 ;
        RECT 98.520 14.615 98.795 14.645 ;
        RECT 87.045 8.875 87.365 8.930 ;
        RECT 92.925 8.875 93.245 8.930 ;
        RECT 87.045 8.725 93.245 8.875 ;
        RECT 87.045 8.670 87.365 8.725 ;
        RECT 92.925 8.670 93.245 8.725 ;
        RECT 112.255 7.825 112.560 36.890 ;
        RECT 114.105 23.430 114.390 39.165 ;
        RECT 139.615 38.765 139.960 49.315 ;
        RECT 115.840 37.265 116.160 37.290 ;
        RECT 132.960 37.265 133.280 37.290 ;
        RECT 115.840 37.055 133.280 37.265 ;
        RECT 115.840 37.030 116.160 37.055 ;
        RECT 132.960 37.030 133.280 37.055 ;
        RECT 123.295 36.260 127.800 36.555 ;
        RECT 126.520 30.920 126.795 30.950 ;
        RECT 124.590 30.645 126.795 30.920 ;
        RECT 124.590 28.305 124.865 30.645 ;
        RECT 126.520 30.615 126.795 30.645 ;
        RECT 122.505 27.090 123.180 27.875 ;
        RECT 115.045 24.875 115.365 24.930 ;
        RECT 120.925 24.875 121.245 24.930 ;
        RECT 115.045 24.725 121.245 24.875 ;
        RECT 115.045 24.670 115.365 24.725 ;
        RECT 120.925 24.670 121.245 24.725 ;
        RECT 114.105 23.145 119.475 23.430 ;
        RECT 86.865 7.445 87.145 7.465 ;
        RECT 86.840 7.405 87.740 7.445 ;
        RECT 86.010 7.005 91.525 7.405 ;
        RECT 112.200 6.765 112.615 7.825 ;
        RECT 114.105 7.470 114.390 23.145 ;
        RECT 140.265 22.765 140.615 49.895 ;
        RECT 140.925 22.085 141.315 50.630 ;
        RECT 146.890 48.490 147.295 49.315 ;
        RECT 146.490 48.085 147.295 48.490 ;
        RECT 144.190 46.565 144.620 47.380 ;
        RECT 146.890 47.255 147.295 48.085 ;
        RECT 143.565 46.135 144.620 46.565 ;
        RECT 144.190 45.320 144.620 46.135 ;
        RECT 150.770 45.100 151.535 45.800 ;
        RECT 148.940 43.595 149.955 44.095 ;
        RECT 141.820 42.945 142.260 42.975 ;
        RECT 141.525 42.475 142.260 42.945 ;
        RECT 141.525 27.170 141.965 42.475 ;
        RECT 140.225 21.695 141.315 22.085 ;
        RECT 115.840 21.265 116.160 21.290 ;
        RECT 132.960 21.265 133.280 21.290 ;
        RECT 115.840 21.055 133.280 21.265 ;
        RECT 115.840 21.030 116.160 21.055 ;
        RECT 132.960 21.030 133.280 21.055 ;
        RECT 123.295 20.260 127.800 20.555 ;
        RECT 126.520 14.920 126.795 14.950 ;
        RECT 124.590 14.645 126.795 14.920 ;
        RECT 122.465 13.335 123.140 14.120 ;
        RECT 124.590 12.305 124.865 14.645 ;
        RECT 126.520 14.615 126.795 14.645 ;
        RECT 115.045 8.875 115.365 8.930 ;
        RECT 120.925 8.875 121.245 8.930 ;
        RECT 115.045 8.725 121.245 8.875 ;
        RECT 115.045 8.670 115.365 8.725 ;
        RECT 120.925 8.670 121.245 8.725 ;
        RECT 114.105 7.185 119.465 7.470 ;
        RECT 114.800 7.115 115.590 7.185 ;
        RECT 114.825 7.095 115.105 7.115 ;
        RECT 140.225 6.765 140.615 21.695 ;
        RECT 142.380 13.435 142.880 41.065 ;
        RECT 3.840 5.265 4.160 5.290 ;
        RECT 20.960 5.265 21.280 5.290 ;
        RECT 3.840 5.055 21.280 5.265 ;
        RECT 3.840 5.030 4.160 5.055 ;
        RECT 20.960 5.030 21.280 5.055 ;
        RECT 31.840 5.265 32.160 5.290 ;
        RECT 48.960 5.265 49.280 5.290 ;
        RECT 31.840 5.055 49.280 5.265 ;
        RECT 31.840 5.030 32.160 5.055 ;
        RECT 48.960 5.030 49.280 5.055 ;
        RECT 59.840 5.265 60.160 5.290 ;
        RECT 76.960 5.265 77.280 5.290 ;
        RECT 59.840 5.055 77.280 5.265 ;
        RECT 59.840 5.030 60.160 5.055 ;
        RECT 76.960 5.030 77.280 5.055 ;
        RECT 87.840 5.265 88.160 5.290 ;
        RECT 104.960 5.265 105.280 5.290 ;
        RECT 87.840 5.055 105.280 5.265 ;
        RECT 87.840 5.030 88.160 5.055 ;
        RECT 104.960 5.030 105.280 5.055 ;
        RECT 115.840 5.265 116.160 5.290 ;
        RECT 132.960 5.265 133.280 5.290 ;
        RECT 115.840 5.055 133.280 5.265 ;
        RECT 115.840 5.030 116.160 5.055 ;
        RECT 132.960 5.030 133.280 5.055 ;
        RECT 11.295 4.260 15.800 4.555 ;
        RECT 39.295 4.260 43.800 4.555 ;
        RECT 67.295 4.260 71.800 4.555 ;
        RECT 80.415 2.885 81.790 4.340 ;
        RECT 95.295 4.260 99.800 4.555 ;
        RECT 123.295 4.260 127.800 4.555 ;
      LAYER met3 ;
        RECT 139.025 205.580 139.355 205.595 ;
        RECT 141.240 205.580 141.740 205.730 ;
        RECT 139.025 205.280 141.740 205.580 ;
        RECT 139.025 205.265 139.355 205.280 ;
        RECT 141.240 205.130 141.740 205.280 ;
        RECT 106.365 202.180 106.695 202.195 ;
        RECT 141.240 202.180 141.740 202.330 ;
        RECT 106.365 201.880 141.740 202.180 ;
        RECT 106.365 201.865 106.695 201.880 ;
        RECT 141.240 201.730 141.740 201.880 ;
        RECT 111.425 200.820 111.755 200.835 ;
        RECT 123.385 200.820 123.715 200.835 ;
        RECT 111.425 200.520 123.715 200.820 ;
        RECT 111.425 200.505 111.755 200.520 ;
        RECT 123.385 200.505 123.715 200.520 ;
        RECT 108.205 200.140 108.535 200.155 ;
        RECT 122.005 200.140 122.335 200.155 ;
        RECT 108.205 199.840 122.335 200.140 ;
        RECT 108.205 199.825 108.535 199.840 ;
        RECT 122.005 199.825 122.335 199.840 ;
        RECT 111.425 198.780 111.755 198.795 ;
        RECT 141.240 198.780 141.740 198.930 ;
        RECT 111.425 198.480 141.740 198.780 ;
        RECT 111.425 198.465 111.755 198.480 ;
        RECT 141.240 198.330 141.740 198.480 ;
        RECT 98.545 196.060 98.875 196.075 ;
        RECT 124.305 196.060 124.635 196.075 ;
        RECT 98.545 195.760 124.635 196.060 ;
        RECT 98.545 195.745 98.875 195.760 ;
        RECT 124.305 195.745 124.635 195.760 ;
        RECT 17.980 195.380 18.480 195.530 ;
        RECT 24.485 195.380 24.815 195.395 ;
        RECT 17.980 195.080 24.815 195.380 ;
        RECT 17.980 194.930 18.480 195.080 ;
        RECT 24.485 195.065 24.815 195.080 ;
        RECT 105.445 195.380 105.775 195.395 ;
        RECT 141.240 195.380 141.740 195.530 ;
        RECT 105.445 195.080 141.740 195.380 ;
        RECT 105.445 195.065 105.775 195.080 ;
        RECT 42.330 194.725 43.910 195.055 ;
        RECT 141.240 194.930 141.740 195.080 ;
        RECT 101.305 194.700 101.635 194.715 ;
        RECT 130.285 194.700 130.615 194.715 ;
        RECT 101.305 194.400 130.615 194.700 ;
        RECT 101.305 194.385 101.635 194.400 ;
        RECT 130.285 194.385 130.615 194.400 ;
        RECT 97.165 194.020 97.495 194.035 ;
        RECT 129.825 194.020 130.155 194.035 ;
        RECT 97.165 193.720 130.155 194.020 ;
        RECT 97.165 193.705 97.495 193.720 ;
        RECT 129.825 193.705 130.155 193.720 ;
        RECT 104.985 193.340 105.315 193.355 ;
        RECT 123.845 193.340 124.175 193.355 ;
        RECT 104.985 193.040 124.175 193.340 ;
        RECT 104.985 193.025 105.315 193.040 ;
        RECT 123.845 193.025 124.175 193.040 ;
        RECT 101.765 192.660 102.095 192.675 ;
        RECT 127.065 192.660 127.395 192.675 ;
        RECT 101.765 192.360 127.395 192.660 ;
        RECT 101.765 192.345 102.095 192.360 ;
        RECT 127.065 192.345 127.395 192.360 ;
        RECT 17.980 191.980 18.480 192.130 ;
        RECT 39.030 192.005 40.610 192.335 ;
        RECT 19.885 191.980 20.215 191.995 ;
        RECT 17.980 191.680 20.215 191.980 ;
        RECT 17.980 191.530 18.480 191.680 ;
        RECT 19.885 191.665 20.215 191.680 ;
        RECT 116.945 191.980 117.275 191.995 ;
        RECT 141.240 191.980 141.740 192.130 ;
        RECT 116.945 191.680 141.740 191.980 ;
        RECT 116.945 191.665 117.275 191.680 ;
        RECT 141.240 191.530 141.740 191.680 ;
        RECT 107.745 191.300 108.075 191.315 ;
        RECT 112.090 191.300 112.470 191.310 ;
        RECT 107.745 191.000 112.470 191.300 ;
        RECT 107.745 190.985 108.075 191.000 ;
        RECT 112.090 190.990 112.470 191.000 ;
        RECT 71.405 190.620 71.735 190.635 ;
        RECT 119.705 190.620 120.035 190.635 ;
        RECT 71.405 190.320 120.035 190.620 ;
        RECT 71.405 190.305 71.735 190.320 ;
        RECT 119.705 190.305 120.035 190.320 ;
        RECT 66.805 189.940 67.135 189.955 ;
        RECT 88.885 189.940 89.215 189.955 ;
        RECT 66.805 189.640 89.215 189.940 ;
        RECT 66.805 189.625 67.135 189.640 ;
        RECT 88.885 189.625 89.215 189.640 ;
        RECT 98.545 189.940 98.875 189.955 ;
        RECT 113.725 189.940 114.055 189.955 ;
        RECT 98.545 189.640 114.055 189.940 ;
        RECT 98.545 189.625 98.875 189.640 ;
        RECT 113.725 189.625 114.055 189.640 ;
        RECT 42.330 189.285 43.910 189.615 ;
        RECT 81.525 189.260 81.855 189.275 ;
        RECT 108.665 189.260 108.995 189.275 ;
        RECT 110.250 189.260 110.630 189.270 ;
        RECT 81.525 188.960 107.830 189.260 ;
        RECT 81.525 188.945 81.855 188.960 ;
        RECT 17.980 188.580 18.480 188.730 ;
        RECT 19.885 188.580 20.215 188.595 ;
        RECT 17.980 188.280 20.215 188.580 ;
        RECT 17.980 188.130 18.480 188.280 ;
        RECT 19.885 188.265 20.215 188.280 ;
        RECT 64.250 188.580 64.630 188.590 ;
        RECT 103.145 188.580 103.475 188.595 ;
        RECT 106.365 188.580 106.695 188.595 ;
        RECT 64.250 188.280 103.475 188.580 ;
        RECT 64.250 188.270 64.630 188.280 ;
        RECT 103.145 188.265 103.475 188.280 ;
        RECT 103.850 188.280 106.695 188.580 ;
        RECT 107.530 188.580 107.830 188.960 ;
        RECT 108.665 188.960 110.630 189.260 ;
        RECT 108.665 188.945 108.995 188.960 ;
        RECT 110.250 188.950 110.630 188.960 ;
        RECT 127.730 189.260 128.110 189.270 ;
        RECT 132.125 189.260 132.455 189.275 ;
        RECT 127.730 188.960 132.455 189.260 ;
        RECT 127.730 188.950 128.110 188.960 ;
        RECT 132.125 188.945 132.455 188.960 ;
        RECT 141.240 188.580 141.740 188.730 ;
        RECT 107.530 188.280 141.740 188.580 ;
        RECT 78.305 187.900 78.635 187.915 ;
        RECT 87.965 187.900 88.295 187.915 ;
        RECT 78.305 187.600 88.295 187.900 ;
        RECT 78.305 187.585 78.635 187.600 ;
        RECT 87.965 187.585 88.295 187.600 ;
        RECT 96.705 187.900 97.035 187.915 ;
        RECT 102.225 187.900 102.555 187.915 ;
        RECT 103.850 187.900 104.150 188.280 ;
        RECT 106.365 188.265 106.695 188.280 ;
        RECT 141.240 188.130 141.740 188.280 ;
        RECT 96.705 187.600 102.555 187.900 ;
        RECT 96.705 187.585 97.035 187.600 ;
        RECT 102.225 187.585 102.555 187.600 ;
        RECT 103.160 187.600 104.150 187.900 ;
        RECT 104.730 187.900 105.110 187.910 ;
        RECT 108.665 187.900 108.995 187.915 ;
        RECT 104.730 187.600 108.995 187.900 ;
        RECT 103.160 187.235 103.460 187.600 ;
        RECT 104.730 187.590 105.110 187.600 ;
        RECT 108.665 187.585 108.995 187.600 ;
        RECT 86.585 187.220 86.915 187.235 ;
        RECT 101.050 187.220 101.430 187.230 ;
        RECT 86.585 186.920 101.430 187.220 ;
        RECT 86.585 186.905 86.915 186.920 ;
        RECT 101.050 186.910 101.430 186.920 ;
        RECT 103.145 186.905 103.475 187.235 ;
        RECT 104.065 187.220 104.395 187.235 ;
        RECT 104.065 186.920 135.430 187.220 ;
        RECT 104.065 186.905 104.395 186.920 ;
        RECT 39.030 186.565 40.610 186.895 ;
        RECT 64.045 186.540 64.375 186.555 ;
        RECT 93.025 186.540 93.355 186.555 ;
        RECT 96.705 186.540 97.035 186.555 ;
        RECT 104.525 186.550 104.855 186.555 ;
        RECT 104.525 186.540 105.110 186.550 ;
        RECT 64.045 186.240 97.035 186.540 ;
        RECT 104.300 186.240 105.110 186.540 ;
        RECT 64.045 186.225 64.375 186.240 ;
        RECT 93.025 186.225 93.355 186.240 ;
        RECT 96.705 186.225 97.035 186.240 ;
        RECT 104.525 186.230 105.110 186.240 ;
        RECT 106.365 186.540 106.695 186.555 ;
        RECT 133.505 186.540 133.835 186.555 ;
        RECT 106.365 186.240 133.835 186.540 ;
        RECT 104.525 186.225 104.855 186.230 ;
        RECT 106.365 186.225 106.695 186.240 ;
        RECT 133.505 186.225 133.835 186.240 ;
        RECT 68.185 185.860 68.515 185.875 ;
        RECT 112.805 185.860 113.135 185.875 ;
        RECT 68.185 185.560 113.135 185.860 ;
        RECT 68.185 185.545 68.515 185.560 ;
        RECT 112.805 185.545 113.135 185.560 ;
        RECT 34.605 185.180 34.935 185.195 ;
        RECT 47.945 185.180 48.275 185.195 ;
        RECT 34.605 184.880 48.275 185.180 ;
        RECT 34.605 184.865 34.935 184.880 ;
        RECT 47.945 184.865 48.275 184.880 ;
        RECT 70.945 185.180 71.275 185.195 ;
        RECT 78.305 185.180 78.635 185.195 ;
        RECT 99.925 185.180 100.255 185.195 ;
        RECT 101.305 185.190 101.635 185.195 ;
        RECT 101.050 185.180 101.635 185.190 ;
        RECT 70.945 184.880 100.255 185.180 ;
        RECT 100.850 184.880 101.635 185.180 ;
        RECT 70.945 184.865 71.275 184.880 ;
        RECT 78.305 184.865 78.635 184.880 ;
        RECT 99.925 184.865 100.255 184.880 ;
        RECT 101.050 184.870 101.635 184.880 ;
        RECT 102.890 185.180 103.270 185.190 ;
        RECT 128.445 185.180 128.775 185.195 ;
        RECT 102.890 184.880 128.775 185.180 ;
        RECT 135.130 185.180 135.430 186.920 ;
        RECT 141.240 185.180 141.740 185.330 ;
        RECT 135.130 184.880 141.740 185.180 ;
        RECT 102.890 184.870 103.270 184.880 ;
        RECT 101.305 184.865 101.635 184.870 ;
        RECT 128.445 184.865 128.775 184.880 ;
        RECT 141.240 184.730 141.740 184.880 ;
        RECT 95.785 184.500 96.115 184.515 ;
        RECT 97.625 184.500 97.955 184.515 ;
        RECT 109.125 184.500 109.455 184.515 ;
        RECT 112.345 184.500 112.675 184.515 ;
        RECT 95.785 184.200 112.675 184.500 ;
        RECT 95.785 184.185 96.115 184.200 ;
        RECT 97.625 184.185 97.955 184.200 ;
        RECT 109.125 184.185 109.455 184.200 ;
        RECT 112.345 184.185 112.675 184.200 ;
        RECT 42.330 183.845 43.910 184.175 ;
        RECT 89.090 183.820 89.470 183.830 ;
        RECT 122.465 183.820 122.795 183.835 ;
        RECT 89.090 183.520 122.795 183.820 ;
        RECT 89.090 183.510 89.470 183.520 ;
        RECT 122.465 183.505 122.795 183.520 ;
        RECT 88.885 183.140 89.215 183.155 ;
        RECT 110.505 183.140 110.835 183.155 ;
        RECT 88.885 182.840 110.835 183.140 ;
        RECT 88.885 182.825 89.215 182.840 ;
        RECT 110.505 182.825 110.835 182.840 ;
        RECT 116.485 183.140 116.815 183.155 ;
        RECT 127.525 183.140 127.855 183.155 ;
        RECT 116.485 182.840 127.855 183.140 ;
        RECT 116.485 182.825 116.815 182.840 ;
        RECT 127.525 182.825 127.855 182.840 ;
        RECT 91.850 182.460 92.230 182.470 ;
        RECT 93.945 182.460 94.275 182.475 ;
        RECT 91.850 182.160 94.275 182.460 ;
        RECT 91.850 182.150 92.230 182.160 ;
        RECT 93.945 182.145 94.275 182.160 ;
        RECT 100.845 182.460 101.175 182.475 ;
        RECT 124.305 182.460 124.635 182.475 ;
        RECT 132.585 182.460 132.915 182.475 ;
        RECT 100.845 182.160 124.635 182.460 ;
        RECT 100.845 182.145 101.175 182.160 ;
        RECT 124.305 182.145 124.635 182.160 ;
        RECT 128.230 182.160 132.915 182.460 ;
        RECT 86.330 181.780 86.710 181.790 ;
        RECT 100.845 181.780 101.175 181.795 ;
        RECT 86.330 181.480 101.175 181.780 ;
        RECT 86.330 181.470 86.710 181.480 ;
        RECT 100.845 181.465 101.175 181.480 ;
        RECT 102.225 181.780 102.555 181.795 ;
        RECT 102.890 181.780 103.270 181.790 ;
        RECT 102.225 181.480 103.270 181.780 ;
        RECT 102.225 181.465 102.555 181.480 ;
        RECT 102.890 181.470 103.270 181.480 ;
        RECT 103.605 181.780 103.935 181.795 ;
        RECT 128.230 181.780 128.530 182.160 ;
        RECT 132.585 182.145 132.915 182.160 ;
        RECT 103.605 181.480 128.530 181.780 ;
        RECT 139.945 181.780 140.275 181.795 ;
        RECT 141.240 181.780 141.740 181.930 ;
        RECT 139.945 181.480 141.740 181.780 ;
        RECT 103.605 181.465 103.935 181.480 ;
        RECT 139.945 181.465 140.275 181.480 ;
        RECT 39.030 181.125 40.610 181.455 ;
        RECT 141.240 181.330 141.740 181.480 ;
        RECT 71.865 181.100 72.195 181.115 ;
        RECT 82.445 181.100 82.775 181.115 ;
        RECT 93.945 181.100 94.275 181.115 ;
        RECT 100.385 181.100 100.715 181.115 ;
        RECT 126.145 181.100 126.475 181.115 ;
        RECT 71.865 180.800 93.110 181.100 ;
        RECT 71.865 180.785 72.195 180.800 ;
        RECT 82.445 180.785 82.775 180.800 ;
        RECT 63.125 180.420 63.455 180.435 ;
        RECT 65.885 180.420 66.215 180.435 ;
        RECT 63.125 180.120 66.215 180.420 ;
        RECT 63.125 180.105 63.455 180.120 ;
        RECT 65.885 180.105 66.215 180.120 ;
        RECT 68.645 180.420 68.975 180.435 ;
        RECT 90.265 180.420 90.595 180.435 ;
        RECT 92.810 180.430 93.110 180.800 ;
        RECT 93.945 180.800 126.475 181.100 ;
        RECT 93.945 180.785 94.275 180.800 ;
        RECT 100.385 180.785 100.715 180.800 ;
        RECT 126.145 180.785 126.475 180.800 ;
        RECT 68.645 180.120 90.595 180.420 ;
        RECT 68.645 180.105 68.975 180.120 ;
        RECT 90.265 180.105 90.595 180.120 ;
        RECT 92.770 180.420 93.150 180.430 ;
        RECT 101.765 180.420 102.095 180.435 ;
        RECT 92.770 180.120 102.095 180.420 ;
        RECT 92.770 180.110 93.150 180.120 ;
        RECT 101.765 180.105 102.095 180.120 ;
        RECT 104.065 180.420 104.395 180.435 ;
        RECT 107.745 180.420 108.075 180.435 ;
        RECT 109.125 180.420 109.455 180.435 ;
        RECT 104.065 180.120 109.455 180.420 ;
        RECT 104.065 180.105 104.395 180.120 ;
        RECT 107.745 180.105 108.075 180.120 ;
        RECT 109.125 180.105 109.455 180.120 ;
        RECT 110.505 180.420 110.835 180.435 ;
        RECT 111.170 180.420 111.550 180.430 ;
        RECT 110.505 180.120 111.550 180.420 ;
        RECT 110.505 180.105 110.835 180.120 ;
        RECT 111.170 180.110 111.550 180.120 ;
        RECT 41.045 179.740 41.375 179.755 ;
        RECT 44.265 179.740 44.595 179.755 ;
        RECT 116.945 179.740 117.275 179.755 ;
        RECT 121.085 179.740 121.415 179.755 ;
        RECT 41.045 179.440 121.415 179.740 ;
        RECT 41.045 179.425 41.375 179.440 ;
        RECT 44.265 179.425 44.595 179.440 ;
        RECT 116.945 179.425 117.275 179.440 ;
        RECT 121.085 179.425 121.415 179.440 ;
        RECT 68.185 179.060 68.515 179.075 ;
        RECT 92.105 179.060 92.435 179.075 ;
        RECT 97.625 179.070 97.955 179.075 ;
        RECT 68.185 178.760 92.435 179.060 ;
        RECT 68.185 178.745 68.515 178.760 ;
        RECT 92.105 178.745 92.435 178.760 ;
        RECT 97.370 179.060 97.955 179.070 ;
        RECT 104.525 179.060 104.855 179.075 ;
        RECT 105.905 179.060 106.235 179.075 ;
        RECT 97.370 178.760 98.180 179.060 ;
        RECT 104.525 178.760 106.235 179.060 ;
        RECT 97.370 178.750 97.955 178.760 ;
        RECT 97.625 178.745 97.955 178.750 ;
        RECT 104.525 178.745 104.855 178.760 ;
        RECT 105.905 178.745 106.235 178.760 ;
        RECT 107.745 179.060 108.075 179.075 ;
        RECT 116.025 179.060 116.355 179.075 ;
        RECT 107.745 178.760 116.355 179.060 ;
        RECT 107.745 178.745 108.075 178.760 ;
        RECT 116.025 178.745 116.355 178.760 ;
        RECT 17.980 178.380 18.480 178.530 ;
        RECT 42.330 178.405 43.910 178.735 ;
        RECT 19.885 178.380 20.215 178.395 ;
        RECT 17.980 178.080 20.215 178.380 ;
        RECT 17.980 177.930 18.480 178.080 ;
        RECT 19.885 178.065 20.215 178.080 ;
        RECT 92.565 178.380 92.895 178.395 ;
        RECT 141.240 178.380 141.740 178.530 ;
        RECT 92.565 178.080 141.740 178.380 ;
        RECT 92.565 178.065 92.895 178.080 ;
        RECT 141.240 177.930 141.740 178.080 ;
        RECT 62.205 177.700 62.535 177.715 ;
        RECT 64.965 177.700 65.295 177.715 ;
        RECT 62.205 177.400 65.295 177.700 ;
        RECT 62.205 177.385 62.535 177.400 ;
        RECT 64.965 177.385 65.295 177.400 ;
        RECT 72.785 177.700 73.115 177.715 ;
        RECT 113.265 177.700 113.595 177.715 ;
        RECT 72.785 177.400 113.595 177.700 ;
        RECT 72.785 177.385 73.115 177.400 ;
        RECT 113.265 177.385 113.595 177.400 ;
        RECT 82.445 177.020 82.775 177.035 ;
        RECT 129.825 177.020 130.155 177.035 ;
        RECT 82.445 176.720 130.155 177.020 ;
        RECT 82.445 176.705 82.775 176.720 ;
        RECT 129.825 176.705 130.155 176.720 ;
        RECT 80.605 176.340 80.935 176.355 ;
        RECT 93.025 176.340 93.355 176.355 ;
        RECT 80.605 176.040 93.355 176.340 ;
        RECT 80.605 176.025 80.935 176.040 ;
        RECT 93.025 176.025 93.355 176.040 ;
        RECT 98.085 176.340 98.415 176.355 ;
        RECT 104.985 176.340 105.315 176.355 ;
        RECT 98.085 176.040 105.315 176.340 ;
        RECT 98.085 176.025 98.415 176.040 ;
        RECT 104.985 176.025 105.315 176.040 ;
        RECT 39.030 175.685 40.610 176.015 ;
        RECT 76.465 175.660 76.795 175.675 ;
        RECT 94.405 175.660 94.735 175.675 ;
        RECT 76.465 175.360 94.735 175.660 ;
        RECT 76.465 175.345 76.795 175.360 ;
        RECT 94.405 175.345 94.735 175.360 ;
        RECT 95.530 175.660 95.910 175.670 ;
        RECT 97.165 175.660 97.495 175.675 ;
        RECT 95.530 175.360 97.495 175.660 ;
        RECT 95.530 175.350 95.910 175.360 ;
        RECT 97.165 175.345 97.495 175.360 ;
        RECT 99.925 175.660 100.255 175.675 ;
        RECT 127.525 175.660 127.855 175.675 ;
        RECT 99.925 175.360 127.855 175.660 ;
        RECT 99.925 175.345 100.255 175.360 ;
        RECT 127.525 175.345 127.855 175.360 ;
        RECT 17.980 174.980 18.480 175.130 ;
        RECT 18.965 174.980 19.295 174.995 ;
        RECT 17.980 174.680 19.295 174.980 ;
        RECT 17.980 174.530 18.480 174.680 ;
        RECT 18.965 174.665 19.295 174.680 ;
        RECT 81.525 174.980 81.855 174.995 ;
        RECT 99.465 174.980 99.795 174.995 ;
        RECT 100.845 174.990 101.175 174.995 ;
        RECT 100.845 174.980 101.430 174.990 ;
        RECT 81.525 174.680 99.795 174.980 ;
        RECT 100.620 174.680 101.430 174.980 ;
        RECT 81.525 174.665 81.855 174.680 ;
        RECT 99.465 174.665 99.795 174.680 ;
        RECT 100.845 174.670 101.430 174.680 ;
        RECT 101.765 174.980 102.095 174.995 ;
        RECT 141.240 174.980 141.740 175.130 ;
        RECT 101.765 174.680 141.740 174.980 ;
        RECT 100.845 174.665 101.175 174.670 ;
        RECT 101.765 174.665 102.095 174.680 ;
        RECT 141.240 174.530 141.740 174.680 ;
        RECT 83.825 174.300 84.155 174.315 ;
        RECT 84.745 174.300 85.075 174.315 ;
        RECT 83.825 174.000 85.075 174.300 ;
        RECT 83.825 173.985 84.155 174.000 ;
        RECT 84.745 173.985 85.075 174.000 ;
        RECT 88.170 174.300 88.550 174.310 ;
        RECT 91.185 174.300 91.515 174.315 ;
        RECT 88.170 174.000 91.515 174.300 ;
        RECT 88.170 173.990 88.550 174.000 ;
        RECT 91.185 173.985 91.515 174.000 ;
        RECT 99.005 174.300 99.335 174.315 ;
        RECT 122.465 174.300 122.795 174.315 ;
        RECT 99.005 174.000 122.795 174.300 ;
        RECT 99.005 173.985 99.335 174.000 ;
        RECT 122.465 173.985 122.795 174.000 ;
        RECT 65.425 173.620 65.755 173.635 ;
        RECT 73.245 173.620 73.575 173.635 ;
        RECT 65.425 173.320 73.575 173.620 ;
        RECT 65.425 173.305 65.755 173.320 ;
        RECT 73.245 173.305 73.575 173.320 ;
        RECT 81.065 173.620 81.395 173.635 ;
        RECT 84.745 173.620 85.075 173.635 ;
        RECT 122.005 173.620 122.335 173.635 ;
        RECT 81.065 173.320 122.335 173.620 ;
        RECT 81.065 173.305 81.395 173.320 ;
        RECT 84.745 173.305 85.075 173.320 ;
        RECT 122.005 173.305 122.335 173.320 ;
        RECT 42.330 172.965 43.910 173.295 ;
        RECT 70.485 172.940 70.815 172.955 ;
        RECT 72.325 172.940 72.655 172.955 ;
        RECT 70.485 172.640 72.655 172.940 ;
        RECT 70.485 172.625 70.815 172.640 ;
        RECT 72.325 172.625 72.655 172.640 ;
        RECT 74.625 172.940 74.955 172.955 ;
        RECT 81.985 172.940 82.315 172.955 ;
        RECT 74.625 172.640 82.315 172.940 ;
        RECT 74.625 172.625 74.955 172.640 ;
        RECT 81.985 172.625 82.315 172.640 ;
        RECT 83.365 172.940 83.695 172.955 ;
        RECT 133.045 172.940 133.375 172.955 ;
        RECT 83.365 172.640 133.375 172.940 ;
        RECT 83.365 172.625 83.695 172.640 ;
        RECT 133.045 172.625 133.375 172.640 ;
        RECT 33.225 172.260 33.555 172.275 ;
        RECT 36.905 172.260 37.235 172.275 ;
        RECT 75.085 172.260 75.415 172.275 ;
        RECT 92.565 172.270 92.895 172.275 ;
        RECT 92.565 172.260 93.150 172.270 ;
        RECT 33.225 171.960 75.415 172.260 ;
        RECT 92.340 171.960 93.150 172.260 ;
        RECT 33.225 171.945 33.555 171.960 ;
        RECT 36.905 171.945 37.235 171.960 ;
        RECT 75.085 171.945 75.415 171.960 ;
        RECT 92.565 171.950 93.150 171.960 ;
        RECT 96.450 172.260 96.830 172.270 ;
        RECT 98.545 172.260 98.875 172.275 ;
        RECT 96.450 171.960 98.875 172.260 ;
        RECT 96.450 171.950 96.830 171.960 ;
        RECT 92.565 171.945 92.895 171.950 ;
        RECT 98.545 171.945 98.875 171.960 ;
        RECT 108.205 172.260 108.535 172.275 ;
        RECT 110.505 172.260 110.835 172.275 ;
        RECT 112.345 172.260 112.675 172.275 ;
        RECT 108.205 171.960 112.675 172.260 ;
        RECT 108.205 171.945 108.535 171.960 ;
        RECT 110.505 171.945 110.835 171.960 ;
        RECT 112.345 171.945 112.675 171.960 ;
        RECT 117.405 172.260 117.735 172.275 ;
        RECT 131.665 172.260 131.995 172.275 ;
        RECT 117.405 171.960 131.995 172.260 ;
        RECT 117.405 171.945 117.735 171.960 ;
        RECT 131.665 171.945 131.995 171.960 ;
        RECT 17.980 171.580 18.480 171.730 ;
        RECT 21.725 171.580 22.055 171.595 ;
        RECT 17.980 171.280 22.055 171.580 ;
        RECT 17.980 171.130 18.480 171.280 ;
        RECT 21.725 171.265 22.055 171.280 ;
        RECT 86.585 171.580 86.915 171.595 ;
        RECT 141.240 171.580 141.740 171.730 ;
        RECT 86.585 171.280 141.740 171.580 ;
        RECT 86.585 171.265 86.915 171.280 ;
        RECT 141.240 171.130 141.740 171.280 ;
        RECT 60.365 170.900 60.695 170.915 ;
        RECT 97.625 170.900 97.955 170.915 ;
        RECT 60.365 170.600 97.955 170.900 ;
        RECT 60.365 170.585 60.695 170.600 ;
        RECT 97.625 170.585 97.955 170.600 ;
        RECT 101.050 170.900 101.430 170.910 ;
        RECT 110.965 170.900 111.295 170.915 ;
        RECT 101.050 170.600 111.295 170.900 ;
        RECT 101.050 170.590 101.430 170.600 ;
        RECT 110.965 170.585 111.295 170.600 ;
        RECT 111.885 170.910 112.215 170.915 ;
        RECT 111.885 170.900 112.470 170.910 ;
        RECT 111.885 170.600 112.670 170.900 ;
        RECT 111.885 170.590 112.470 170.600 ;
        RECT 111.885 170.585 112.215 170.590 ;
        RECT 39.030 170.245 40.610 170.575 ;
        RECT 46.105 170.220 46.435 170.235 ;
        RECT 72.325 170.220 72.655 170.235 ;
        RECT 86.585 170.230 86.915 170.235 ;
        RECT 86.330 170.220 86.915 170.230 ;
        RECT 46.105 169.920 72.655 170.220 ;
        RECT 86.130 169.920 86.915 170.220 ;
        RECT 46.105 169.905 46.435 169.920 ;
        RECT 72.325 169.905 72.655 169.920 ;
        RECT 86.330 169.910 86.915 169.920 ;
        RECT 86.585 169.905 86.915 169.910 ;
        RECT 87.505 170.220 87.835 170.235 ;
        RECT 107.490 170.220 107.870 170.230 ;
        RECT 87.505 169.920 107.870 170.220 ;
        RECT 87.505 169.905 87.835 169.920 ;
        RECT 107.490 169.910 107.870 169.920 ;
        RECT 71.405 169.540 71.735 169.555 ;
        RECT 87.505 169.540 87.835 169.555 ;
        RECT 132.585 169.540 132.915 169.555 ;
        RECT 71.405 169.240 132.915 169.540 ;
        RECT 71.405 169.225 71.735 169.240 ;
        RECT 87.505 169.225 87.835 169.240 ;
        RECT 132.585 169.225 132.915 169.240 ;
        RECT 54.385 168.860 54.715 168.875 ;
        RECT 78.765 168.860 79.095 168.875 ;
        RECT 88.170 168.860 88.550 168.870 ;
        RECT 54.385 168.560 88.550 168.860 ;
        RECT 54.385 168.545 54.715 168.560 ;
        RECT 78.765 168.545 79.095 168.560 ;
        RECT 88.170 168.550 88.550 168.560 ;
        RECT 89.805 168.860 90.135 168.875 ;
        RECT 93.690 168.860 94.070 168.870 ;
        RECT 89.805 168.560 94.070 168.860 ;
        RECT 89.805 168.545 90.135 168.560 ;
        RECT 93.690 168.550 94.070 168.560 ;
        RECT 100.385 168.860 100.715 168.875 ;
        RECT 104.065 168.860 104.395 168.875 ;
        RECT 100.385 168.560 104.395 168.860 ;
        RECT 100.385 168.545 100.715 168.560 ;
        RECT 104.065 168.545 104.395 168.560 ;
        RECT 107.745 168.860 108.075 168.875 ;
        RECT 110.250 168.860 110.630 168.870 ;
        RECT 107.745 168.560 110.630 168.860 ;
        RECT 107.745 168.545 108.075 168.560 ;
        RECT 110.250 168.550 110.630 168.560 ;
        RECT 17.980 168.180 18.480 168.330 ;
        RECT 21.725 168.180 22.055 168.195 ;
        RECT 17.980 167.880 22.055 168.180 ;
        RECT 17.980 167.730 18.480 167.880 ;
        RECT 21.725 167.865 22.055 167.880 ;
        RECT 44.725 168.180 45.055 168.195 ;
        RECT 53.005 168.180 53.335 168.195 ;
        RECT 44.725 167.880 53.335 168.180 ;
        RECT 44.725 167.865 45.055 167.880 ;
        RECT 53.005 167.865 53.335 167.880 ;
        RECT 68.645 168.180 68.975 168.195 ;
        RECT 82.905 168.180 83.235 168.195 ;
        RECT 68.645 167.880 83.235 168.180 ;
        RECT 68.645 167.865 68.975 167.880 ;
        RECT 82.905 167.865 83.235 167.880 ;
        RECT 86.585 168.180 86.915 168.195 ;
        RECT 141.240 168.180 141.740 168.330 ;
        RECT 86.585 167.880 141.740 168.180 ;
        RECT 86.585 167.865 86.915 167.880 ;
        RECT 42.330 167.525 43.910 167.855 ;
        RECT 141.240 167.730 141.740 167.880 ;
        RECT 50.245 167.500 50.575 167.515 ;
        RECT 57.145 167.500 57.475 167.515 ;
        RECT 50.245 167.200 57.475 167.500 ;
        RECT 50.245 167.185 50.575 167.200 ;
        RECT 57.145 167.185 57.475 167.200 ;
        RECT 74.165 167.500 74.495 167.515 ;
        RECT 88.425 167.500 88.755 167.515 ;
        RECT 108.665 167.500 108.995 167.515 ;
        RECT 74.165 167.200 108.995 167.500 ;
        RECT 74.165 167.185 74.495 167.200 ;
        RECT 88.425 167.185 88.755 167.200 ;
        RECT 108.665 167.185 108.995 167.200 ;
        RECT 37.825 166.820 38.155 166.835 ;
        RECT 47.485 166.820 47.815 166.835 ;
        RECT 53.005 166.820 53.335 166.835 ;
        RECT 37.825 166.520 53.335 166.820 ;
        RECT 37.825 166.505 38.155 166.520 ;
        RECT 47.485 166.505 47.815 166.520 ;
        RECT 53.005 166.505 53.335 166.520 ;
        RECT 54.845 166.820 55.175 166.835 ;
        RECT 58.985 166.820 59.315 166.835 ;
        RECT 54.845 166.520 59.315 166.820 ;
        RECT 54.845 166.505 55.175 166.520 ;
        RECT 58.985 166.505 59.315 166.520 ;
        RECT 73.705 166.820 74.035 166.835 ;
        RECT 89.345 166.820 89.675 166.835 ;
        RECT 94.865 166.820 95.195 166.835 ;
        RECT 73.705 166.520 95.195 166.820 ;
        RECT 73.705 166.505 74.035 166.520 ;
        RECT 89.345 166.505 89.675 166.520 ;
        RECT 94.865 166.505 95.195 166.520 ;
        RECT 97.625 166.820 97.955 166.835 ;
        RECT 100.845 166.820 101.175 166.835 ;
        RECT 102.225 166.820 102.555 166.835 ;
        RECT 97.625 166.520 102.555 166.820 ;
        RECT 97.625 166.505 97.955 166.520 ;
        RECT 100.845 166.505 101.175 166.520 ;
        RECT 102.225 166.505 102.555 166.520 ;
        RECT 107.490 166.820 107.870 166.830 ;
        RECT 126.145 166.820 126.475 166.835 ;
        RECT 107.490 166.520 126.475 166.820 ;
        RECT 107.490 166.510 107.870 166.520 ;
        RECT 126.145 166.505 126.475 166.520 ;
        RECT 53.005 166.140 53.335 166.155 ;
        RECT 53.925 166.140 54.255 166.155 ;
        RECT 53.005 165.840 54.255 166.140 ;
        RECT 53.005 165.825 53.335 165.840 ;
        RECT 53.925 165.825 54.255 165.840 ;
        RECT 91.185 166.140 91.515 166.155 ;
        RECT 91.850 166.140 92.230 166.150 ;
        RECT 94.405 166.140 94.735 166.155 ;
        RECT 91.185 165.840 94.735 166.140 ;
        RECT 91.185 165.825 91.515 165.840 ;
        RECT 91.850 165.830 92.230 165.840 ;
        RECT 94.405 165.825 94.735 165.840 ;
        RECT 96.245 166.140 96.575 166.155 ;
        RECT 102.225 166.140 102.555 166.155 ;
        RECT 103.145 166.140 103.475 166.155 ;
        RECT 96.245 165.840 103.475 166.140 ;
        RECT 96.245 165.825 96.575 165.840 ;
        RECT 102.225 165.825 102.555 165.840 ;
        RECT 103.145 165.825 103.475 165.840 ;
        RECT 53.925 165.460 54.255 165.475 ;
        RECT 61.745 165.460 62.075 165.475 ;
        RECT 53.925 165.160 62.075 165.460 ;
        RECT 53.925 165.145 54.255 165.160 ;
        RECT 61.745 165.145 62.075 165.160 ;
        RECT 93.485 165.460 93.815 165.475 ;
        RECT 103.145 165.460 103.475 165.475 ;
        RECT 112.345 165.460 112.675 165.475 ;
        RECT 93.485 165.160 112.675 165.460 ;
        RECT 93.485 165.145 93.815 165.160 ;
        RECT 103.145 165.145 103.475 165.160 ;
        RECT 112.345 165.145 112.675 165.160 ;
        RECT 17.980 164.780 18.480 164.930 ;
        RECT 39.030 164.805 40.610 165.135 ;
        RECT 20.805 164.780 21.135 164.795 ;
        RECT 17.980 164.480 21.135 164.780 ;
        RECT 17.980 164.330 18.480 164.480 ;
        RECT 20.805 164.465 21.135 164.480 ;
        RECT 46.105 164.780 46.435 164.795 ;
        RECT 80.145 164.780 80.475 164.795 ;
        RECT 46.105 164.480 80.475 164.780 ;
        RECT 46.105 164.465 46.435 164.480 ;
        RECT 80.145 164.465 80.475 164.480 ;
        RECT 87.965 164.780 88.295 164.795 ;
        RECT 141.240 164.780 141.740 164.930 ;
        RECT 87.965 164.480 141.740 164.780 ;
        RECT 87.965 164.465 88.295 164.480 ;
        RECT 141.240 164.330 141.740 164.480 ;
        RECT 57.145 164.100 57.475 164.115 ;
        RECT 64.045 164.110 64.375 164.115 ;
        RECT 64.045 164.100 64.630 164.110 ;
        RECT 57.145 163.800 64.630 164.100 ;
        RECT 57.145 163.785 57.475 163.800 ;
        RECT 64.045 163.790 64.630 163.800 ;
        RECT 79.225 164.100 79.555 164.115 ;
        RECT 80.145 164.100 80.475 164.115 ;
        RECT 79.225 163.800 80.475 164.100 ;
        RECT 64.045 163.785 64.375 163.790 ;
        RECT 79.225 163.785 79.555 163.800 ;
        RECT 80.145 163.785 80.475 163.800 ;
        RECT 83.825 164.100 84.155 164.115 ;
        RECT 104.525 164.100 104.855 164.115 ;
        RECT 83.825 163.800 104.855 164.100 ;
        RECT 83.825 163.785 84.155 163.800 ;
        RECT 104.525 163.785 104.855 163.800 ;
        RECT 43.805 163.420 44.135 163.435 ;
        RECT 84.285 163.420 84.615 163.435 ;
        RECT 43.805 163.120 84.615 163.420 ;
        RECT 43.805 163.105 44.135 163.120 ;
        RECT 84.285 163.105 84.615 163.120 ;
        RECT 88.425 163.420 88.755 163.435 ;
        RECT 89.090 163.420 89.470 163.430 ;
        RECT 88.425 163.120 89.470 163.420 ;
        RECT 88.425 163.105 88.755 163.120 ;
        RECT 89.090 163.110 89.470 163.120 ;
        RECT 91.645 163.420 91.975 163.435 ;
        RECT 107.745 163.420 108.075 163.435 ;
        RECT 91.645 163.120 108.075 163.420 ;
        RECT 91.645 163.105 91.975 163.120 ;
        RECT 107.745 163.105 108.075 163.120 ;
        RECT 79.225 162.740 79.555 162.755 ;
        RECT 83.825 162.740 84.155 162.755 ;
        RECT 79.225 162.440 84.155 162.740 ;
        RECT 79.225 162.425 79.555 162.440 ;
        RECT 83.825 162.425 84.155 162.440 ;
        RECT 85.665 162.740 85.995 162.755 ;
        RECT 104.985 162.740 105.315 162.755 ;
        RECT 85.665 162.440 105.315 162.740 ;
        RECT 85.665 162.425 85.995 162.440 ;
        RECT 104.985 162.425 105.315 162.440 ;
        RECT 42.330 162.085 43.910 162.415 ;
        RECT 80.145 162.060 80.475 162.075 ;
        RECT 82.445 162.060 82.775 162.075 ;
        RECT 80.145 161.760 82.775 162.060 ;
        RECT 80.145 161.745 80.475 161.760 ;
        RECT 82.445 161.745 82.775 161.760 ;
        RECT 95.785 162.060 96.115 162.075 ;
        RECT 97.625 162.070 97.955 162.075 ;
        RECT 96.450 162.060 96.830 162.070 ;
        RECT 95.785 161.760 96.830 162.060 ;
        RECT 95.785 161.745 96.115 161.760 ;
        RECT 96.450 161.750 96.830 161.760 ;
        RECT 97.370 162.060 97.955 162.070 ;
        RECT 97.370 161.760 98.180 162.060 ;
        RECT 97.370 161.750 97.955 161.760 ;
        RECT 97.625 161.745 97.955 161.750 ;
        RECT 76.465 161.380 76.795 161.395 ;
        RECT 80.605 161.380 80.935 161.395 ;
        RECT 76.465 161.080 80.935 161.380 ;
        RECT 76.465 161.065 76.795 161.080 ;
        RECT 80.605 161.065 80.935 161.080 ;
        RECT 84.745 161.380 85.075 161.395 ;
        RECT 141.240 161.380 141.740 161.530 ;
        RECT 84.745 161.080 141.740 161.380 ;
        RECT 84.745 161.065 85.075 161.080 ;
        RECT 141.240 160.930 141.740 161.080 ;
        RECT 58.065 160.700 58.395 160.715 ;
        RECT 64.505 160.700 64.835 160.715 ;
        RECT 58.065 160.400 64.835 160.700 ;
        RECT 58.065 160.385 58.395 160.400 ;
        RECT 64.505 160.385 64.835 160.400 ;
        RECT 78.765 160.700 79.095 160.715 ;
        RECT 99.005 160.700 99.335 160.715 ;
        RECT 78.765 160.400 99.335 160.700 ;
        RECT 78.765 160.385 79.095 160.400 ;
        RECT 99.005 160.385 99.335 160.400 ;
        RECT 99.925 160.700 100.255 160.715 ;
        RECT 108.205 160.700 108.535 160.715 ;
        RECT 99.925 160.400 108.535 160.700 ;
        RECT 99.925 160.385 100.255 160.400 ;
        RECT 108.205 160.385 108.535 160.400 ;
        RECT 77.385 160.020 77.715 160.035 ;
        RECT 79.685 160.020 80.015 160.035 ;
        RECT 85.205 160.020 85.535 160.035 ;
        RECT 77.385 159.720 85.535 160.020 ;
        RECT 77.385 159.705 77.715 159.720 ;
        RECT 79.685 159.705 80.015 159.720 ;
        RECT 85.205 159.705 85.535 159.720 ;
        RECT 90.265 160.020 90.595 160.035 ;
        RECT 113.265 160.020 113.595 160.035 ;
        RECT 90.265 159.720 113.595 160.020 ;
        RECT 90.265 159.705 90.595 159.720 ;
        RECT 113.265 159.705 113.595 159.720 ;
        RECT 39.030 159.365 40.610 159.695 ;
        RECT 64.045 159.340 64.375 159.355 ;
        RECT 67.265 159.340 67.595 159.355 ;
        RECT 98.085 159.340 98.415 159.355 ;
        RECT 102.685 159.340 103.015 159.355 ;
        RECT 64.045 159.040 103.015 159.340 ;
        RECT 64.045 159.025 64.375 159.040 ;
        RECT 67.265 159.025 67.595 159.040 ;
        RECT 98.085 159.025 98.415 159.040 ;
        RECT 102.685 159.025 103.015 159.040 ;
        RECT 68.185 158.660 68.515 158.675 ;
        RECT 83.825 158.660 84.155 158.675 ;
        RECT 95.325 158.670 95.655 158.675 ;
        RECT 95.325 158.660 95.910 158.670 ;
        RECT 68.185 158.360 84.155 158.660 ;
        RECT 95.100 158.360 95.910 158.660 ;
        RECT 68.185 158.345 68.515 158.360 ;
        RECT 83.825 158.345 84.155 158.360 ;
        RECT 95.325 158.350 95.910 158.360 ;
        RECT 95.325 158.345 95.655 158.350 ;
        RECT 41.045 157.980 41.375 157.995 ;
        RECT 87.965 157.980 88.295 157.995 ;
        RECT 41.045 157.680 88.295 157.980 ;
        RECT 41.045 157.665 41.375 157.680 ;
        RECT 87.965 157.665 88.295 157.680 ;
        RECT 89.345 157.980 89.675 157.995 ;
        RECT 141.240 157.980 141.740 158.130 ;
        RECT 89.345 157.680 141.740 157.980 ;
        RECT 89.345 157.665 89.675 157.680 ;
        RECT 141.240 157.530 141.740 157.680 ;
        RECT 82.445 157.300 82.775 157.315 ;
        RECT 93.485 157.300 93.815 157.315 ;
        RECT 82.445 157.000 93.815 157.300 ;
        RECT 82.445 156.985 82.775 157.000 ;
        RECT 93.485 156.985 93.815 157.000 ;
        RECT 42.330 156.645 43.910 156.975 ;
        RECT 84.285 156.620 84.615 156.635 ;
        RECT 109.125 156.620 109.455 156.635 ;
        RECT 129.825 156.620 130.155 156.635 ;
        RECT 84.285 156.320 109.455 156.620 ;
        RECT 84.285 156.305 84.615 156.320 ;
        RECT 109.125 156.305 109.455 156.320 ;
        RECT 128.230 156.320 130.155 156.620 ;
        RECT 55.765 155.940 56.095 155.955 ;
        RECT 60.825 155.940 61.155 155.955 ;
        RECT 55.765 155.640 61.155 155.940 ;
        RECT 55.765 155.625 56.095 155.640 ;
        RECT 60.825 155.625 61.155 155.640 ;
        RECT 79.225 155.940 79.555 155.955 ;
        RECT 88.885 155.940 89.215 155.955 ;
        RECT 79.225 155.640 89.215 155.940 ;
        RECT 79.225 155.625 79.555 155.640 ;
        RECT 88.885 155.625 89.215 155.640 ;
        RECT 71.865 155.260 72.195 155.275 ;
        RECT 85.205 155.260 85.535 155.275 ;
        RECT 111.170 155.260 111.550 155.270 ;
        RECT 128.230 155.260 128.530 156.320 ;
        RECT 129.825 156.305 130.155 156.320 ;
        RECT 71.865 154.960 128.530 155.260 ;
        RECT 71.865 154.945 72.195 154.960 ;
        RECT 85.205 154.945 85.535 154.960 ;
        RECT 111.170 154.950 111.550 154.960 ;
        RECT 17.980 154.580 18.480 154.730 ;
        RECT 21.725 154.580 22.055 154.595 ;
        RECT 17.980 154.280 22.055 154.580 ;
        RECT 17.980 154.130 18.480 154.280 ;
        RECT 21.725 154.265 22.055 154.280 ;
        RECT 69.565 154.580 69.895 154.595 ;
        RECT 141.240 154.580 141.740 154.730 ;
        RECT 69.565 154.280 141.740 154.580 ;
        RECT 69.565 154.265 69.895 154.280 ;
        RECT 39.030 153.925 40.610 154.255 ;
        RECT 141.240 154.130 141.740 154.280 ;
        RECT 61.745 153.900 62.075 153.915 ;
        RECT 68.645 153.900 68.975 153.915 ;
        RECT 61.745 153.600 68.975 153.900 ;
        RECT 61.745 153.585 62.075 153.600 ;
        RECT 68.645 153.585 68.975 153.600 ;
        RECT 93.690 153.900 94.070 153.910 ;
        RECT 132.125 153.900 132.455 153.915 ;
        RECT 93.690 153.600 132.455 153.900 ;
        RECT 93.690 153.590 94.070 153.600 ;
        RECT 132.125 153.585 132.455 153.600 ;
        RECT 73.245 153.220 73.575 153.235 ;
        RECT 94.405 153.220 94.735 153.235 ;
        RECT 73.245 152.920 94.735 153.220 ;
        RECT 73.245 152.905 73.575 152.920 ;
        RECT 94.405 152.905 94.735 152.920 ;
        RECT 127.730 153.220 128.110 153.230 ;
        RECT 132.585 153.220 132.915 153.235 ;
        RECT 127.730 152.920 132.915 153.220 ;
        RECT 127.730 152.910 128.110 152.920 ;
        RECT 132.585 152.905 132.915 152.920 ;
        RECT 42.330 151.205 43.910 151.535 ;
        RECT 126.145 151.180 126.475 151.195 ;
        RECT 141.240 151.180 141.740 151.330 ;
        RECT 126.145 150.880 141.740 151.180 ;
        RECT 126.145 150.865 126.475 150.880 ;
        RECT 141.240 150.730 141.740 150.880 ;
        RECT 60.365 149.820 60.695 149.835 ;
        RECT 60.365 149.520 128.530 149.820 ;
        RECT 60.365 149.505 60.695 149.520 ;
        RECT 128.230 147.780 128.530 149.520 ;
        RECT 141.240 147.780 141.740 147.930 ;
        RECT 128.230 147.480 141.740 147.780 ;
        RECT 141.240 147.330 141.740 147.480 ;
        RECT 133.965 144.380 134.295 144.395 ;
        RECT 141.240 144.380 141.740 144.530 ;
        RECT 133.965 144.080 141.740 144.380 ;
        RECT 133.965 144.065 134.295 144.080 ;
        RECT 141.240 143.930 141.740 144.080 ;
        RECT 66.345 140.980 66.675 140.995 ;
        RECT 141.240 140.980 141.740 141.130 ;
        RECT 66.345 140.680 141.740 140.980 ;
        RECT 66.345 140.665 66.675 140.680 ;
        RECT 141.240 140.530 141.740 140.680 ;
        RECT 79.480 50.170 80.050 50.690 ;
        RECT 68.665 49.870 69.975 49.875 ;
        RECT 68.635 48.950 70.005 49.870 ;
        RECT 68.665 48.945 69.975 48.950 ;
        RECT 146.510 48.490 146.965 48.515 ;
        RECT 94.645 48.085 146.965 48.490 ;
        RECT 94.645 46.215 95.050 48.085 ;
        RECT 146.510 48.060 146.965 48.085 ;
        RECT 143.585 46.565 144.065 46.590 ;
        RECT 95.565 46.470 107.495 46.565 ;
        RECT 109.175 46.470 144.065 46.565 ;
        RECT 95.565 46.135 144.065 46.470 ;
        RECT 79.805 34.570 81.180 36.025 ;
        RECT 68.665 34.225 69.975 34.230 ;
        RECT 68.635 33.330 70.005 34.225 ;
        RECT 68.665 33.325 69.975 33.330 ;
        RECT 95.565 32.295 95.995 46.135 ;
        RECT 143.585 46.110 144.065 46.135 ;
        RECT 150.825 45.680 151.375 45.705 ;
        RECT 94.695 31.865 95.995 32.295 ;
        RECT 96.770 45.180 151.375 45.680 ;
        RECT 80.460 18.535 81.835 19.990 ;
        RECT 68.660 16.800 69.980 18.180 ;
        RECT 96.770 16.190 97.270 45.180 ;
        RECT 150.825 45.155 151.375 45.180 ;
        RECT 148.960 44.095 149.510 44.120 ;
        RECT 122.495 43.595 149.510 44.095 ;
        RECT 148.960 43.570 149.510 43.595 ;
        RECT 141.500 27.655 141.990 27.680 ;
        RECT 122.590 27.215 141.990 27.655 ;
        RECT 141.500 27.190 141.990 27.215 ;
        RECT 94.530 15.690 97.270 16.190 ;
        RECT 142.355 13.980 142.905 14.005 ;
        RECT 122.560 13.480 142.905 13.980 ;
        RECT 142.355 13.455 142.905 13.480 ;
        RECT 7.350 7.445 7.730 7.470 ;
        RECT 7.350 7.115 142.905 7.445 ;
        RECT 7.350 7.090 7.730 7.115 ;
        RECT 80.415 2.885 81.790 4.340 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 39.020 151.130 40.620 195.130 ;
        RECT 42.320 151.130 43.920 195.130 ;
        RECT 112.115 190.985 112.445 191.315 ;
        RECT 110.275 188.945 110.605 189.275 ;
        RECT 64.275 188.265 64.605 188.595 ;
        RECT 64.290 164.115 64.590 188.265 ;
        RECT 104.755 187.585 105.085 187.915 ;
        RECT 101.075 186.905 101.405 187.235 ;
        RECT 101.090 185.195 101.390 186.905 ;
        RECT 104.770 186.555 105.070 187.585 ;
        RECT 104.755 186.225 105.085 186.555 ;
        RECT 101.075 184.865 101.405 185.195 ;
        RECT 102.915 184.865 103.245 185.195 ;
        RECT 89.115 183.505 89.445 183.835 ;
        RECT 86.355 181.465 86.685 181.795 ;
        RECT 86.370 170.235 86.670 181.465 ;
        RECT 88.195 173.985 88.525 174.315 ;
        RECT 86.355 169.905 86.685 170.235 ;
        RECT 88.210 168.875 88.510 173.985 ;
        RECT 88.195 168.545 88.525 168.875 ;
        RECT 64.275 163.785 64.605 164.115 ;
        RECT 89.130 163.435 89.430 183.505 ;
        RECT 91.875 182.145 92.205 182.475 ;
        RECT 91.890 166.155 92.190 182.145 ;
        RECT 102.930 181.795 103.230 184.865 ;
        RECT 102.915 181.465 103.245 181.795 ;
        RECT 92.795 180.105 93.125 180.435 ;
        RECT 92.810 172.275 93.110 180.105 ;
        RECT 97.395 178.745 97.725 179.075 ;
        RECT 95.555 175.345 95.885 175.675 ;
        RECT 92.795 171.945 93.125 172.275 ;
        RECT 93.715 168.545 94.045 168.875 ;
        RECT 91.875 165.825 92.205 166.155 ;
        RECT 89.115 163.105 89.445 163.435 ;
        RECT 93.730 153.915 94.030 168.545 ;
        RECT 95.570 158.675 95.870 175.345 ;
        RECT 96.475 171.945 96.805 172.275 ;
        RECT 96.490 162.075 96.790 171.945 ;
        RECT 97.410 162.075 97.710 178.745 ;
        RECT 101.075 174.665 101.405 174.995 ;
        RECT 101.090 170.915 101.390 174.665 ;
        RECT 101.075 170.585 101.405 170.915 ;
        RECT 107.515 169.905 107.845 170.235 ;
        RECT 107.530 166.835 107.830 169.905 ;
        RECT 110.290 168.875 110.590 188.945 ;
        RECT 111.195 180.105 111.525 180.435 ;
        RECT 110.275 168.545 110.605 168.875 ;
        RECT 107.515 166.505 107.845 166.835 ;
        RECT 96.475 161.745 96.805 162.075 ;
        RECT 97.395 161.745 97.725 162.075 ;
        RECT 95.555 158.345 95.885 158.675 ;
        RECT 111.210 155.275 111.510 180.105 ;
        RECT 112.130 170.915 112.430 190.985 ;
        RECT 127.755 188.945 128.085 189.275 ;
        RECT 112.115 170.585 112.445 170.915 ;
        RECT 111.195 154.945 111.525 155.275 ;
        RECT 93.715 153.585 94.045 153.915 ;
        RECT 127.770 153.235 128.070 188.945 ;
        RECT 127.755 152.905 128.085 153.235 ;
        RECT 80.525 50.625 81.705 50.740 ;
        RECT 79.535 50.230 81.705 50.625 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 68.660 18.155 69.980 49.875 ;
        RECT 80.525 35.855 81.705 50.230 ;
        RECT 79.870 34.675 81.705 35.855 ;
        RECT 68.655 16.825 69.985 18.155 ;
        RECT 80.525 4.270 81.705 34.675 ;
        RECT 80.495 3.030 81.735 4.270 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

