magic
tech sky130A
magscale 1 2
timestamp 1757923025
<< nwell >>
rect -12800 1806 -12300 3900
rect -12770 1805 -12300 1806
rect -12749 1802 -12300 1805
rect -7100 1800 -6600 3900
rect -1600 1813 -1100 3900
rect -1620 1806 -1100 1813
rect -1402 1805 -1100 1806
rect -1288 1800 -1100 1805
rect 4100 1800 4600 3900
rect -12800 -1394 -12300 700
rect -7200 -1394 -6700 700
rect -12507 -1400 -12300 -1394
rect -6890 -1400 -6700 -1394
rect -1500 -1400 -1000 700
rect 4100 -1400 4600 700
rect -12700 -4600 -12200 -2500
rect -7200 -4591 -6700 -2500
rect -7206 -4594 -6700 -4591
rect -7159 -4595 -6700 -4594
rect -6835 -4596 -6700 -4595
rect -1500 -4600 -1000 -2500
rect 4100 -4600 4600 -2500
<< locali >>
rect -5972 4422 -4724 4432
rect -5972 4350 -5962 4422
rect -4738 4350 -4724 4422
rect -5972 4342 -4724 4350
rect -17941 4089 -16266 4095
rect -17941 4074 -16360 4089
rect -17941 4012 -17916 4074
rect -17941 4002 -16360 4012
rect -16273 4002 -16266 4089
rect -17941 3996 -16266 4002
rect -2700 4044 -2186 4062
rect -2700 3974 -2684 4044
rect -2202 3974 -2186 4044
rect -2700 3958 -2186 3974
rect 11898 2072 12610 2084
rect 11898 1996 11920 2072
rect 12594 1996 12610 2072
rect 11898 1974 12610 1996
<< viali >>
rect -5962 4350 -4738 4422
rect -16360 4074 -16273 4089
rect -17916 4012 -16273 4074
rect -16360 4002 -16273 4012
rect -2684 3974 -2202 4044
rect 11920 1996 12594 2072
<< metal1 >>
rect -17840 4900 -17460 5380
rect -17280 5260 -16220 5380
rect -16064 5250 -15634 5406
rect -15478 5250 -15472 5406
rect -17280 4900 -16220 5020
rect -17800 4180 -17420 4660
rect -17280 4540 -16220 4660
rect -16080 4540 -15700 5020
rect -5974 4432 -5932 4438
rect -5974 4422 -4724 4432
rect -5974 4350 -5962 4422
rect -4738 4350 -4724 4422
rect -5974 4342 -4724 4350
rect -5974 4336 -5932 4342
rect -16080 4299 -15615 4300
rect -17280 4160 -16220 4280
rect -16080 4160 -15022 4299
rect -14890 4175 -13826 4294
rect -13109 4286 -13034 4313
rect -10045 4299 -9020 4300
rect -13696 4260 -12632 4286
rect -13696 4185 -13109 4260
rect -13034 4185 -12632 4260
rect -15714 4158 -15022 4160
rect -17946 3996 -17940 4095
rect -17841 4089 -16261 4095
rect -17841 4074 -16360 4089
rect -17841 4002 -16360 4012
rect -16273 4002 -16261 4089
rect -17841 3996 -16261 4002
rect -16154 3954 -16148 4043
rect -16059 4024 -16053 4043
rect -14852 4024 -14801 4175
rect -13696 4167 -12632 4185
rect -12494 4178 -9020 4299
rect -8880 4180 -7820 4320
rect -7680 4267 -6620 4300
rect -7680 4187 -7496 4267
rect -7416 4187 -6620 4267
rect -12487 4039 -12406 4178
rect -10045 4160 -9020 4178
rect -8831 4050 -8756 4180
rect -7680 4160 -6620 4187
rect -6480 4160 -4200 4300
rect -4080 4160 -3020 4300
rect -2880 4180 -1820 4300
rect -1632 4244 -1553 4283
rect -6445 4060 -6364 4160
rect -16059 3973 -14801 4024
rect -16059 3954 -16053 3973
rect -12945 3958 -12939 4039
rect -12858 3958 -12406 4039
rect -10547 3975 -10541 4050
rect -10466 3975 -8756 4050
rect -7325 3979 -7319 4060
rect -7238 3979 -6364 4060
rect -4055 4055 -3985 4160
rect -1902 4071 -1834 4180
rect -1664 4156 -1276 4244
rect -1632 4075 -1553 4156
rect -4945 3985 -4939 4055
rect -4869 3985 -3985 4055
rect -2700 4051 -2186 4062
rect -2700 4044 -2353 4051
rect -2270 4044 -2186 4051
rect -2700 3974 -2684 4044
rect -2202 3974 -2186 4044
rect -1908 4003 -1902 4071
rect -1834 4003 -1828 4071
rect -1716 3996 -1710 4075
rect -1631 3996 -1553 4075
rect -1364 4144 -1276 4156
rect 10580 4144 10980 4160
rect -1364 4056 10980 4144
rect -2700 3968 -2353 3974
rect -2270 3968 -2186 3974
rect -2700 3958 -2186 3968
rect -12760 3780 -12220 3920
rect -7180 3780 -6640 3920
rect -16193 3684 -16015 3690
rect -17940 3593 -17841 3599
rect -15640 3616 -15634 3772
rect -15478 3616 -15472 3772
rect -1560 3780 -1100 3920
rect 4060 3780 4520 3920
rect 10580 3680 10980 4056
rect -10593 3667 -10415 3673
rect -16193 3589 -16015 3595
rect -10593 3586 -10415 3592
rect -4993 3618 -4815 3624
rect -4993 3542 -4815 3548
rect -17940 1900 -17841 3494
rect 10580 3394 10980 3420
rect 10574 2994 10580 3394
rect 10666 2994 10980 3394
rect 11114 3381 11120 3781
rect 11201 3780 11207 3781
rect 11201 3381 11520 3780
rect 11120 3300 11520 3381
rect 10580 2940 10980 2994
rect 11120 2960 11912 3060
rect 12012 2960 12720 3060
rect 11627 2743 11727 2749
rect 10580 2513 10980 2700
rect 11120 2643 11627 2680
rect 11727 2643 12180 2680
rect 11120 2580 12180 2643
rect 12320 2580 12720 2960
rect 10100 2425 10106 2513
rect 10194 2425 10980 2513
rect -16831 1809 -16765 2241
rect -12735 1883 -12535 1889
rect -12580 1831 -12535 1883
rect -12735 1825 -12535 1831
rect -11234 1868 -11164 2397
rect -11234 1792 -11164 1798
rect -16831 1737 -16765 1743
rect -7141 1683 -7135 1883
rect -7080 1683 -7074 1883
rect -5635 1845 -5566 2275
rect -5635 1770 -5566 1776
rect -1541 1683 -1535 1883
rect -1483 1683 -1477 1883
rect -39 1844 41 2371
rect 10580 2220 10980 2425
rect 12455 2320 12613 2325
rect 11120 2220 12180 2320
rect 12320 2220 12662 2320
rect -39 1758 41 1764
rect 4059 1683 4065 1883
rect 4126 1683 4132 1883
rect 5571 1814 5628 2208
rect 11648 2172 11804 2220
rect 11648 2131 11748 2172
rect 10212 2031 10218 2131
rect 10318 2031 11748 2131
rect 12455 2123 12613 2220
rect 11899 2072 12613 2123
rect 11899 1996 11920 2072
rect 12594 1996 12613 2072
rect 11899 1965 12613 1996
rect 11899 1935 12057 1965
rect 5571 1751 5628 1757
rect 9659 1683 9665 1883
rect 9734 1683 9740 1883
rect 9963 1777 12057 1935
rect -2292 1097 -2276 1116
rect -2292 1095 -2280 1097
rect -2292 1081 -2284 1095
rect -12660 800 -12300 980
rect -7140 800 -6660 980
rect 9215 991 9373 1133
rect 9963 991 10121 1777
rect -1540 800 -1060 980
rect 4040 800 4580 980
rect 9215 833 10121 991
rect -12700 580 -12160 720
rect -7180 560 -6660 720
rect -4526 594 -4520 694
rect -4268 594 -4262 694
rect -1580 580 -1000 720
rect 3980 580 4580 720
rect -16193 468 -16015 474
rect -16193 387 -16015 393
rect -10593 444 -10415 450
rect -10593 358 -10415 364
rect -4993 432 -4815 438
rect -4993 358 -4815 364
rect -16825 -1397 -16759 -934
rect -12735 -1317 -12535 -1311
rect -12735 -1392 -12535 -1386
rect -16825 -1469 -16759 -1463
rect -11235 -1399 -11165 -1021
rect -11235 -1475 -11165 -1469
rect -7141 -1517 -7135 -1317
rect -7083 -1517 -7077 -1317
rect -5625 -1391 -5556 -922
rect -5625 -1466 -5556 -1460
rect -1401 -1517 -1395 -1317
rect -1335 -1517 -1329 -1317
rect -33 -1394 47 -1031
rect -33 -1480 47 -1474
rect 4059 -1517 4065 -1317
rect 4130 -1517 4136 -1317
rect 5574 -1390 5631 -989
rect 5574 -1453 5631 -1447
rect 9789 -1517 9795 -1317
rect 9865 -1517 9871 -1317
rect -12680 -2400 -12260 -2220
rect -7160 -2400 -6660 -2220
rect -1500 -2400 -1080 -2220
rect -12700 -2620 -12120 -2480
rect -7180 -2620 -6680 -2480
rect -4489 -2485 -4301 -2479
rect -1520 -2620 -1020 -2480
rect -4489 -2679 -4301 -2673
rect -10593 -2730 -10415 -2724
rect -10593 -2817 -10415 -2811
rect -4993 -2766 -4815 -2760
rect -4993 -2851 -4815 -2845
rect -16193 -2869 -16015 -2863
rect -16193 -2956 -16015 -2950
rect -4426 -2873 -4364 -2679
rect -4426 -2935 -3804 -2873
rect -4426 -3147 -4364 -2935
rect -3866 -3014 -3804 -2935
rect -16832 -4587 -16766 -3932
rect -12735 -4517 -12535 -4511
rect -12735 -4579 -12535 -4573
rect -16832 -4659 -16766 -4653
rect -11216 -4592 -11146 -4203
rect -11216 -4668 -11146 -4662
rect -7006 -4717 -7000 -4517
rect -6935 -4717 -6929 -4517
rect -5633 -4583 -5564 -4010
rect -5633 -4658 -5564 -4652
rect -1415 -4717 -1409 -4517
rect -1335 -4717 -1329 -4517
rect -39 -4595 41 -4198
rect -39 -4681 41 -4675
rect 4176 -4717 4182 -4517
rect 4265 -4717 4271 -4517
rect 5572 -4582 5629 -4106
rect 5572 -4645 5629 -4639
rect 9781 -4717 9787 -4517
rect 9865 -4717 9871 -4517
rect -12660 -5600 -12240 -5420
rect -7100 -5600 -6680 -5420
rect -2159 -5464 -2153 -5228
rect -1917 -5464 -1911 -5228
rect -1480 -5600 -1060 -5420
rect 4060 -5600 4480 -5420
<< via1 >>
rect -15634 5250 -15478 5406
rect -13109 4185 -13034 4260
rect -17940 4074 -17841 4095
rect -17940 4012 -17916 4074
rect -17916 4012 -17841 4074
rect -17940 3996 -17841 4012
rect -16148 3954 -16059 4043
rect -7496 4187 -7416 4267
rect -12939 3958 -12858 4039
rect -10541 3975 -10466 4050
rect -7319 3979 -7238 4060
rect -4939 3985 -4869 4055
rect -2353 4044 -2270 4051
rect -2353 3974 -2270 4044
rect -1902 4003 -1834 4071
rect -1710 3996 -1631 4075
rect -2353 3968 -2270 3974
rect -17940 3494 -17841 3593
rect -16193 3595 -16015 3684
rect -15634 3616 -15478 3772
rect -4520 3713 -4268 3899
rect -10593 3592 -10415 3667
rect -4993 3548 -4815 3618
rect 671 3167 752 3248
rect 10580 2994 10666 3394
rect 11120 3381 11201 3781
rect 11912 2960 12012 3060
rect 6241 2643 6341 2743
rect 11627 2643 11727 2743
rect 10106 2425 10194 2513
rect -12735 1831 -12580 1883
rect -16831 1743 -16765 1809
rect -11234 1798 -11164 1868
rect -7135 1683 -7080 1883
rect -5635 1776 -5566 1845
rect -1535 1683 -1483 1883
rect -39 1764 41 1844
rect 4065 1683 4126 1883
rect 10218 2031 10318 2131
rect 5571 1757 5628 1814
rect 9665 1683 9734 1883
rect -2284 859 -2048 1095
rect -4520 594 -4268 694
rect -16193 393 -16015 468
rect -10593 364 -10415 444
rect -4993 364 -4815 432
rect 681 297 767 383
rect 6260 -633 6348 -545
rect -12735 -1386 -12535 -1317
rect -16825 -1463 -16759 -1397
rect -11235 -1469 -11165 -1399
rect -7135 -1517 -7083 -1317
rect -5625 -1460 -5556 -1391
rect -1395 -1517 -1335 -1317
rect -33 -1474 47 -1394
rect 4065 -1517 4130 -1317
rect 5574 -1447 5631 -1390
rect 9795 -1517 9865 -1317
rect -2153 -2349 -1917 -2113
rect -4489 -2673 -4301 -2485
rect -10593 -2811 -10415 -2730
rect -4993 -2845 -4815 -2766
rect -16193 -2950 -16015 -2869
rect 648 -2938 748 -2838
rect 6254 -3380 6354 -3280
rect -12735 -4573 -12535 -4517
rect -16832 -4653 -16766 -4587
rect -11216 -4662 -11146 -4592
rect -7000 -4717 -6935 -4517
rect -5633 -4652 -5564 -4583
rect -1409 -4717 -1335 -4517
rect -39 -4675 41 -4595
rect 4182 -4717 4265 -4517
rect 5572 -4639 5629 -4582
rect 9787 -4717 9865 -4517
rect -2153 -5464 -1917 -5228
<< metal2 >>
rect -15634 5406 -15478 5412
rect -17940 4095 -17841 4101
rect -17940 3593 -17841 3996
rect -16148 4043 -16059 4049
rect -16148 3684 -16059 3954
rect -15634 3772 -15478 5250
rect -16199 3595 -16193 3684
rect -16015 3595 -16009 3684
rect -15634 3610 -15478 3616
rect -13109 4260 -13034 4266
rect -17946 3494 -17940 3593
rect -17841 3494 -17835 3593
rect -17880 1743 -16831 1809
rect -16765 1743 -16759 1809
rect -17880 -1397 -17814 1743
rect -13109 468 -13034 4185
rect -16199 393 -16193 468
rect -16015 393 -13034 468
rect -12939 4039 -12858 4045
rect -17880 -1463 -16825 -1397
rect -16759 -1463 -16753 -1397
rect -17878 -4587 -17812 -1463
rect -12939 -2869 -12858 3958
rect -12660 1900 -12610 4625
rect -12660 1883 -12560 1900
rect -12741 1831 -12735 1883
rect -12580 1831 -12560 1883
rect -12620 1820 -12560 1831
rect -12515 1734 -12446 4614
rect -12669 1665 -12446 1734
rect -12669 -1317 -12600 1665
rect -12328 1548 -12272 4608
rect -7496 4267 -7416 4273
rect -10541 4050 -10466 4056
rect -10541 3667 -10466 3975
rect -10599 3592 -10593 3667
rect -10415 3592 -10409 3667
rect -12488 1492 -12272 1548
rect -12180 1798 -11234 1868
rect -11164 1798 -11158 1868
rect -12741 -1386 -12735 -1317
rect -12535 -1386 -12529 -1317
rect -12488 -1432 -12432 1492
rect -16199 -2950 -16193 -2869
rect -16015 -2950 -12858 -2869
rect -12663 -1488 -12432 -1432
rect -12180 -1399 -12110 1798
rect -7496 444 -7416 4187
rect -10599 364 -10593 444
rect -10415 364 -7416 444
rect -7319 4060 -7238 4066
rect -12180 -1469 -11235 -1399
rect -11165 -1469 -11159 -1399
rect -12663 -4517 -12607 -1488
rect -12741 -4573 -12735 -4517
rect -12535 -4573 -12529 -4517
rect -17878 -4653 -16832 -4587
rect -16717 -4653 -16708 -4587
rect -12180 -4592 -12110 -1469
rect -7319 -2730 -7238 3979
rect -7135 1883 -7080 4647
rect -7135 1677 -7080 1683
rect -6985 1544 -6936 4644
rect -7133 1495 -6936 1544
rect -7133 -1311 -7084 1495
rect -6853 1352 -6788 4632
rect -1902 4071 -1834 4077
rect -4939 4055 -4869 4061
rect -4939 3618 -4869 3985
rect -2362 4051 -2248 4062
rect -2362 3968 -2353 4051
rect -2270 3968 -2248 4051
rect -2362 3958 -2248 3968
rect -4545 3899 -4232 3911
rect -4545 3713 -4520 3899
rect -4268 3713 -4232 3899
rect -4545 3695 -4232 3713
rect -4999 3548 -4993 3618
rect -4815 3548 -4809 3618
rect -7000 1287 -6788 1352
rect -6737 1776 -5635 1845
rect -5566 1776 -5560 1845
rect -7135 -1317 -7083 -1311
rect -7135 -1523 -7083 -1517
rect -10599 -2811 -10593 -2730
rect -10415 -2811 -7238 -2730
rect -7000 -4517 -6935 1287
rect -6737 -1391 -6668 1776
rect -2297 1095 -2022 1129
rect -2297 859 -2284 1095
rect -2048 859 -2022 1095
rect -2297 838 -2022 859
rect -4529 594 -4520 765
rect -4268 594 -4259 765
rect -4520 588 -4268 594
rect -1902 432 -1834 4003
rect -1710 4075 -1631 4081
rect -1710 1481 -1631 3996
rect -1531 1889 -1487 4603
rect -1535 1883 -1483 1889
rect -1535 1677 -1483 1683
rect -1710 1402 -1485 1481
rect -4999 364 -4993 432
rect -4815 364 -1834 432
rect -6737 -1460 -5625 -1391
rect -5556 -1460 -5550 -1391
rect -11122 -4587 -11066 -4583
rect -11217 -4592 -11061 -4587
rect -12180 -4662 -11216 -4592
rect -11146 -4648 -11122 -4592
rect -11066 -4648 -11061 -4592
rect -11146 -4653 -11061 -4648
rect -11146 -4657 -11066 -4653
rect -11146 -4662 -11097 -4657
rect -11185 -4663 -11097 -4662
rect -6733 -4583 -6664 -1460
rect -2166 -2113 -1891 -2078
rect -2166 -2349 -2153 -2113
rect -1917 -2349 -1891 -2113
rect -2166 -2369 -1891 -2349
rect -4509 -2464 -4280 -2455
rect -4509 -2702 -4280 -2693
rect -1564 -2766 -1485 1402
rect -1395 -1317 -1335 4588
rect -1235 4495 -1162 4595
rect -1395 -1523 -1335 -1517
rect -1236 -1604 -1162 4495
rect -1079 3503 -1018 4593
rect -951 3613 -886 4590
rect -816 3727 -755 4593
rect -686 3856 -617 4592
rect -545 3973 -475 4589
rect -394 4128 -316 4567
rect -394 4050 10005 4128
rect -545 3903 9865 3973
rect -686 3787 9734 3856
rect -816 3666 4368 3727
rect -951 3548 4250 3613
rect -1079 3448 4126 3503
rect -1079 3442 3304 3448
rect 3514 3442 4126 3448
rect 637 3248 790 3284
rect 637 3167 671 3248
rect 752 3167 790 3248
rect 637 3144 790 3167
rect 4065 1883 4126 3442
rect -1062 1764 -39 1844
rect 41 1764 47 1844
rect -4999 -2845 -4993 -2766
rect -4815 -2845 -1485 -2766
rect -1409 -1678 -1162 -1604
rect -1056 -1394 -976 1764
rect 4065 1677 4126 1683
rect 4185 1516 4250 3548
rect 4065 1451 4250 1516
rect 663 383 816 417
rect 663 297 681 383
rect 767 297 816 383
rect 663 277 816 297
rect 4065 -1317 4130 1451
rect 4307 1363 4368 3666
rect 6226 2743 6361 2784
rect 6226 2643 6241 2743
rect 6341 2643 6361 2743
rect 6226 2627 6361 2643
rect 9665 1883 9734 3787
rect -1056 -1474 -33 -1394
rect 47 -1474 53 -1394
rect -1409 -4517 -1335 -1678
rect -6733 -4592 -5633 -4583
rect -6733 -4648 -6552 -4592
rect -6496 -4648 -5633 -4592
rect -6733 -4652 -5633 -4648
rect -5564 -4652 -5558 -4583
rect -6557 -4653 -6405 -4652
rect -6552 -4657 -6496 -4653
rect -7000 -4723 -6935 -4717
rect -1056 -4595 -976 -1474
rect 4065 -1523 4130 -1517
rect 4193 1302 4368 1363
rect 4563 1757 5571 1814
rect 5628 1757 5634 1814
rect 617 -2838 770 -2818
rect 617 -2938 648 -2838
rect 748 -2938 770 -2838
rect 617 -2958 770 -2938
rect 4193 -4511 4254 1302
rect 4563 -1390 4620 1757
rect 9665 1677 9734 1683
rect 6243 -545 6378 -501
rect 6243 -633 6260 -545
rect 6348 -633 6378 -545
rect 6243 -658 6378 -633
rect 9795 -1317 9865 3903
rect 4563 -1447 5574 -1390
rect 5631 -1447 5637 -1390
rect 4182 -4517 4265 -4511
rect -885 -4587 -829 -4583
rect -890 -4592 -710 -4587
rect -890 -4595 -885 -4592
rect -1056 -4648 -885 -4595
rect -829 -4595 -710 -4592
rect -829 -4648 -39 -4595
rect -1056 -4675 -39 -4648
rect 41 -4675 47 -4595
rect -1409 -4723 -1335 -4717
rect 4563 -4582 4620 -1447
rect 9795 -1523 9865 -1517
rect 9927 -1659 10005 4050
rect 11120 3781 11201 3787
rect 11040 3541 11049 3622
rect 10580 3394 10666 3400
rect 10455 3151 10464 3237
rect 10550 3151 10580 3237
rect 11120 3375 11201 3381
rect 10580 2988 10666 2994
rect 11896 3060 12049 3084
rect 11896 2960 11912 3060
rect 12012 2960 12049 3060
rect 11896 2944 12049 2960
rect 11530 2643 11539 2743
rect 11727 2643 11733 2743
rect 10106 2513 10194 2519
rect 10047 2425 10106 2513
rect 10047 2419 10194 2425
rect 10047 -545 10135 2419
rect 10047 -642 10135 -633
rect 10218 2131 10318 2137
rect 9787 -1737 10005 -1659
rect 6235 -3280 6370 -3252
rect 6235 -3380 6254 -3280
rect 6354 -3380 6370 -3280
rect 6235 -3409 6370 -3380
rect 9787 -4517 9865 -1737
rect 10218 -3280 10318 2031
rect 10218 -3389 10318 -3380
rect 4563 -4592 5572 -4582
rect 4563 -4639 4707 -4592
rect 4702 -4648 4707 -4639
rect 4763 -4639 5572 -4592
rect 5629 -4639 5635 -4582
rect 4763 -4648 4860 -4639
rect 4702 -4653 4860 -4648
rect 4707 -4657 4763 -4653
rect 4182 -4723 4265 -4717
rect 9787 -4723 9865 -4717
rect -2175 -5228 -1900 -5208
rect -2175 -5464 -2153 -5228
rect -1917 -5464 -1900 -5228
rect -2175 -5499 -1900 -5464
<< via2 >>
rect -16783 -4653 -16766 -4587
rect -16766 -4653 -16717 -4587
rect -2348 3973 -2275 4046
rect -4520 3718 -4268 3894
rect -2279 864 -2053 1090
rect -4520 694 -4268 765
rect -4520 594 -4268 694
rect -11122 -4648 -11066 -4592
rect -2148 -2344 -1922 -2118
rect -4509 -2485 -4280 -2464
rect -4509 -2673 -4489 -2485
rect -4489 -2673 -4301 -2485
rect -4301 -2673 -4280 -2485
rect -4509 -2693 -4280 -2673
rect 676 3172 747 3243
rect 686 302 762 378
rect 6246 2648 6336 2738
rect -6552 -4648 -6496 -4592
rect 653 -2933 743 -2843
rect 6265 -628 6343 -550
rect -885 -4648 -829 -4592
rect 11049 3541 11120 3622
rect 11120 3541 11130 3622
rect 10464 3151 10550 3237
rect 11912 2960 12012 3060
rect 11539 2643 11627 2743
rect 11627 2643 11639 2743
rect 10047 -633 10135 -545
rect 6259 -3375 6349 -3285
rect 10218 -3380 10318 -3280
rect 4707 -4648 4763 -4592
rect -2153 -5464 -1917 -5228
<< metal3 >>
rect -2362 4048 -2248 4062
rect -2362 3971 -2350 4048
rect -2273 3971 -2248 4048
rect -2362 3958 -2248 3971
rect -4525 3898 -4263 3899
rect -4531 3714 -4525 3898
rect -4263 3714 -4257 3898
rect -4525 3713 -4263 3714
rect 11044 3622 11135 3627
rect 671 3541 11049 3622
rect 11130 3541 11135 3622
rect 671 3243 752 3541
rect 11044 3536 11135 3541
rect 671 3172 676 3243
rect 747 3172 752 3243
rect 10459 3237 10555 3242
rect 671 3167 752 3172
rect 855 3218 3241 3237
rect 3577 3218 10464 3237
rect 855 3151 10464 3218
rect 10550 3151 10555 3237
rect -2297 1094 -2022 1129
rect -2297 860 -2283 1094
rect -2049 860 -2022 1094
rect -2297 838 -2022 860
rect -4525 769 -4263 770
rect -4531 590 -4525 769
rect -4263 590 -4257 769
rect -4525 589 -4263 590
rect 855 383 941 3151
rect 10459 3146 10555 3151
rect 11907 3060 12017 3065
rect 681 378 941 383
rect 681 302 686 378
rect 762 302 941 378
rect 681 297 941 302
rect 1096 2960 11912 3060
rect 12012 2960 12017 3060
rect -2166 -2114 -1891 -2078
rect -2166 -2348 -2152 -2114
rect -1918 -2348 -1891 -2114
rect -2166 -2369 -1891 -2348
rect -4526 -2446 -4262 -2440
rect -4526 -2716 -4262 -2710
rect 1096 -2838 1196 2960
rect 11907 2955 12017 2960
rect 11534 2743 11644 2748
rect 6241 2738 11539 2743
rect 6241 2648 6246 2738
rect 6336 2648 11539 2738
rect 6241 2643 11539 2648
rect 11639 2643 11644 2743
rect 11534 2638 11644 2643
rect 10042 -545 10140 -540
rect 6260 -550 10047 -545
rect 6260 -628 6265 -550
rect 6343 -628 10047 -550
rect 6260 -633 10047 -628
rect 10135 -633 10140 -545
rect 10042 -638 10140 -633
rect 648 -2843 1196 -2838
rect 648 -2933 653 -2843
rect 743 -2933 1196 -2843
rect 648 -2938 1196 -2933
rect 10213 -3280 10323 -3275
rect 6254 -3285 10218 -3280
rect 6254 -3375 6259 -3285
rect 6349 -3375 10218 -3285
rect 6254 -3380 10218 -3375
rect 10318 -3380 10323 -3280
rect 10213 -3385 10323 -3380
rect -16788 -4587 -16712 -4582
rect -16788 -4653 -16783 -4587
rect -16717 -4592 10323 -4587
rect -16717 -4648 -11122 -4592
rect -11066 -4648 -6552 -4592
rect -6496 -4648 -885 -4592
rect -829 -4648 4707 -4592
rect 4763 -4648 10323 -4592
rect -16717 -4653 10323 -4648
rect -16788 -4658 -16712 -4653
rect -2175 -5223 -1900 -5208
rect -2175 -5469 -2158 -5223
rect -1912 -5469 -1900 -5223
rect -2175 -5499 -1900 -5469
<< via3 >>
rect -2350 4046 -2273 4048
rect -2350 3973 -2348 4046
rect -2348 3973 -2275 4046
rect -2275 3973 -2273 4046
rect -2350 3971 -2273 3973
rect -4525 3894 -4263 3898
rect -4525 3718 -4520 3894
rect -4520 3718 -4268 3894
rect -4268 3718 -4263 3894
rect -4525 3714 -4263 3718
rect -2283 1090 -2049 1094
rect -2283 864 -2279 1090
rect -2279 864 -2053 1090
rect -2053 864 -2049 1090
rect -2283 860 -2049 864
rect -4525 765 -4263 769
rect -4525 594 -4520 765
rect -4520 594 -4268 765
rect -4268 594 -4263 765
rect -4525 590 -4263 594
rect -2152 -2118 -1918 -2114
rect -2152 -2344 -2148 -2118
rect -2148 -2344 -1922 -2118
rect -1922 -2344 -1918 -2118
rect -2152 -2348 -1918 -2344
rect -4526 -2464 -4262 -2446
rect -4526 -2693 -4509 -2464
rect -4509 -2693 -4280 -2464
rect -4280 -2693 -4262 -2464
rect -4526 -2710 -4262 -2693
rect -2158 -5228 -1912 -5223
rect -2158 -5464 -2153 -5228
rect -2153 -5464 -1917 -5228
rect -1917 -5464 -1912 -5228
rect -2158 -5469 -1912 -5464
<< metal4 >>
rect -2153 4049 -1917 4072
rect -2351 4048 -1917 4049
rect -2351 3971 -2350 4048
rect -2273 3971 -1917 4048
rect -2351 3970 -1917 3971
rect -4526 3898 -4262 3899
rect -4526 3714 -4525 3898
rect -4263 3714 -4262 3898
rect -4526 769 -4262 3714
rect -2153 1095 -1917 3970
rect -2284 1094 -1917 1095
rect -2284 860 -2283 1094
rect -2049 860 -1917 1094
rect -2284 859 -1917 860
rect -4526 590 -4525 769
rect -4263 590 -4262 769
rect -4526 -2445 -4262 590
rect -2153 -2114 -1917 859
rect -2153 -2348 -2152 -2114
rect -1918 -2348 -1917 -2114
rect -4527 -2446 -4261 -2445
rect -4527 -2710 -4526 -2446
rect -4262 -2710 -4261 -2446
rect -4527 -2711 -4261 -2710
rect -2153 -5222 -1917 -2348
rect -2159 -5223 -1911 -5222
rect -2159 -5469 -2158 -5223
rect -1912 -5469 -1911 -5223
rect -2159 -5470 -1911 -5469
use compr  compr_0
timestamp 1757923025
transform 1 0 3890 0 1 -4197
box 510 -1403 5975 1713
use compr  compr_1
timestamp 1757923025
transform 1 0 -1710 0 1 -4197
box 510 -1403 5975 1713
use compr  compr_2
timestamp 1757923025
transform 1 0 -7310 0 1 -4197
box 510 -1403 5975 1713
use compr  compr_3
timestamp 1757923025
transform 1 0 -12910 0 1 -4197
box 510 -1403 5975 1713
use compr  compr_4
timestamp 1757923025
transform 1 0 -18510 0 1 -4197
box 510 -1403 5975 1713
use compr  compr_5
timestamp 1757923025
transform 1 0 3890 0 1 -997
box 510 -1403 5975 1713
use compr  compr_6
timestamp 1757923025
transform 1 0 -1710 0 1 -997
box 510 -1403 5975 1713
use compr  compr_7
timestamp 1757923025
transform 1 0 -7310 0 1 -997
box 510 -1403 5975 1713
use compr  compr_8
timestamp 1757923025
transform 1 0 -12910 0 1 -997
box 510 -1403 5975 1713
use compr  compr_9
timestamp 1757923025
transform 1 0 -18510 0 1 -997
box 510 -1403 5975 1713
use compr  compr_10
timestamp 1757923025
transform 1 0 3890 0 1 2203
box 510 -1403 5975 1713
use compr  compr_11
timestamp 1757923025
transform 1 0 -1710 0 1 2203
box 510 -1403 5975 1713
use compr  compr_12
timestamp 1757923025
transform 1 0 -7310 0 1 2203
box 510 -1403 5975 1713
use compr  compr_13
timestamp 1757923025
transform 1 0 -12910 0 1 2203
box 510 -1403 5975 1713
use compr  compr_14
timestamp 1757923025
transform 1 0 -18510 0 1 2203
box 510 -1403 5975 1713
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_0
timestamp 1757903622
transform 0 1 -1753 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_1
timestamp 1757903622
transform 0 -1 11051 1 0 2271
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_2
timestamp 1757903622
transform 0 1 11051 -1 0 2635
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_3
timestamp 1757903622
transform 0 1 -2949 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_4
timestamp 1757903622
transform 0 1 11051 -1 0 2999
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_5
timestamp 1757903622
transform 0 1 -4145 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_6
timestamp 1757903622
transform 0 1 -17349 -1 0 5327
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_7
timestamp 1757903622
transform 0 1 -6553 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_8
timestamp 1757903622
transform 0 1 11051 -1 0 3363
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_9
timestamp 1757903622
transform 0 1 11051 -1 0 3727
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_10
timestamp 1757903622
transform 0 1 -8945 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_11
timestamp 1757903622
transform 0 1 -7749 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_12
timestamp 1757903622
transform 0 1 -16153 -1 0 5327
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_13
timestamp 1757903622
transform 0 1 12247 -1 0 2635
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_14
timestamp 1757903622
transform 0 1 12247 -1 0 2271
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_15
timestamp 1757903622
transform 0 1 -17349 -1 0 4963
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_16
timestamp 1757903622
transform 0 1 -16153 -1 0 4599
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_17
timestamp 1757903622
transform 0 1 -17349 -1 0 4599
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_18
timestamp 1757903622
transform 0 1 -12565 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_19
timestamp 1757903622
transform 0 1 -13761 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_20
timestamp 1757903622
transform 0 1 -14957 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_21
timestamp 1757903622
transform 0 1 -16153 -1 0 4963
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_22
timestamp 1757903622
transform 0 1 -16153 -1 0 4235
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  sky130_fd_pr__res_high_po_0p69_ZKG2N9_23
timestamp 1757903622
transform 0 1 -17349 -1 0 4235
box -235 -651 235 651
<< labels >>
rlabel metal2 -12652 4551 -12615 4615 1 AF14
port 1 n
rlabel metal2 -7121 4505 -7086 4628 1 AF13
port 2 n
rlabel metal2 -1529 4460 -1494 4583 1 AF12
port 3 n
rlabel metal2 -1066 4460 -1031 4583 1 AF11
port 4 n
rlabel metal2 -670 4449 -635 4572 1 AF10
port 5 n
rlabel metal2 -379 4225 -327 4365 1 AF0
port 6 n
rlabel metal2 -810 4425 -758 4565 1 AF1
port 7 n
rlabel metal2 -1234 4452 -1182 4592 1 AF2
port 8 n
rlabel metal2 -6846 4476 -6794 4616 1 AF3
port 9 n
rlabel metal2 -12328 4461 -12276 4601 1 AF4
port 10 n
rlabel metal2 -536 4422 -484 4562 1 AF5
port 11 n
rlabel metal2 -946 4402 -894 4542 1 AF6
port 12 n
rlabel space -1385 4393 -1333 4533 1 AF7
port 13 n
rlabel space -6987 4495 -6935 4635 1 AF8
port 14 n
rlabel metal2 -12506 4446 -12454 4586 1 AF9
port 15 n
rlabel metal4 -2134 -59 -1920 275 1 VSS
port 16 n
rlabel metal4 -4500 629 -4286 963 1 VDD
port 17 n
rlabel metal3 9910 -4650 10320 -4590 1 A0
port 18 n
<< end >>
