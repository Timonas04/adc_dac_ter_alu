magic
tech sky130A
magscale 1 2
timestamp 1757965112
<< pwell >>
rect 8367 -3739 9064 -3591
rect 1420 -5416 1508 -4264
rect 8916 -5304 9064 -3739
rect 8916 -5452 12848 -5304
rect 12854 -5940 12970 -5932
rect 1858 -5998 12992 -5940
rect 12854 -6064 12970 -5998
<< locali >>
rect 7106 -3289 7540 -3186
rect 7780 -3208 8632 -3088
rect 7106 -3392 7226 -3289
rect 7329 -3392 7540 -3289
rect 7106 -3460 7540 -3392
rect 1382 -4286 1766 -4228
rect -3605 -4668 -3498 -4583
rect -3605 -4698 -3542 -4668
rect -3383 -4698 -3362 -4614
rect -3586 -5766 -3542 -4698
rect -3392 -5766 -3362 -4698
rect 1382 -5396 1470 -4286
rect 1704 -5396 1766 -4286
rect 5746 -5108 6712 -4990
rect 6884 -5064 7376 -4774
rect 6884 -5088 8450 -5064
rect 6884 -5106 7834 -5088
rect 6888 -5112 7834 -5106
rect 5772 -5174 7834 -5112
rect 8356 -5174 8450 -5088
rect 5772 -5234 8450 -5174
rect 5772 -5242 8212 -5234
rect 1382 -5446 1766 -5396
rect -3586 -5806 -3362 -5766
rect -9510 -5880 -7416 -5806
rect -9510 -6138 -9460 -5880
rect -7460 -6138 -7416 -5880
rect 1888 -5968 12912 -5966
rect 1888 -6004 12978 -5968
rect -9510 -6186 -7416 -6138
rect -4040 -6082 -3398 -6032
rect 1888 -6054 12912 -6004
rect -4040 -6338 -3964 -6082
rect -3464 -6330 -3398 -6082
rect -2822 -6268 2144 -6266
rect -2950 -6330 2144 -6268
rect -4040 -6382 -3514 -6338
rect -3462 -6376 2144 -6330
rect -3462 -6382 -1510 -6376
rect -4040 -6390 -2770 -6382
rect -4026 -7080 -4006 -6978
rect -3464 -7080 -3438 -6978
rect -4026 -7096 -3438 -7080
<< viali >>
rect 7226 -3392 7329 -3289
rect -3498 -4668 -3383 -4583
rect -3542 -4698 -3383 -4668
rect -3542 -5766 -3392 -4698
rect 1470 -5396 1704 -4286
rect 7834 -5174 8356 -5088
rect -9460 -6138 -7460 -5880
rect -3964 -6330 -3464 -6082
rect -3964 -6338 -3462 -6330
rect -3514 -6382 -3462 -6338
rect -4006 -7080 -3464 -6938
<< metal1 >>
rect 7356 -3102 7907 -3037
rect 7356 -3152 8597 -3102
rect 7356 -3283 7471 -3152
rect 7792 -3217 8597 -3152
rect 7588 -3255 7662 -3220
rect 6604 -3289 7471 -3283
rect 6604 -3392 7226 -3289
rect 7329 -3392 7471 -3289
rect 6604 -3398 7471 -3392
rect 6180 -3573 6295 -3567
rect 6604 -3573 6719 -3398
rect 5795 -3688 6180 -3575
rect 6295 -3688 6779 -3573
rect 5795 -3755 6779 -3688
rect 7581 -3830 7664 -3255
rect 8744 -3312 8818 -3212
rect 7776 -3430 8622 -3324
rect 5403 -3913 7664 -3830
rect -3886 -4296 -3686 -4280
rect -1150 -4296 -1046 -4232
rect -9512 -4506 -9000 -4428
rect -7521 -4506 -7515 -4460
rect -9512 -4583 -7515 -4506
rect -7392 -4506 -7386 -4460
rect -6868 -4482 -6853 -4296
rect -6730 -4318 -1584 -4296
rect -6730 -4324 -1577 -4318
rect -6730 -4453 -1706 -4324
rect -6730 -4459 -1577 -4453
rect -6730 -4482 -1584 -4459
rect -1270 -4482 -1264 -4296
rect -1135 -4482 -1046 -4296
rect -7392 -4583 -7382 -4506
rect -9512 -4688 -7382 -4583
rect -3504 -4577 -3377 -4571
rect -6348 -4600 -4382 -4596
rect -7024 -4844 -3844 -4600
rect -3586 -4668 -3504 -4626
rect -3586 -4734 -3542 -4668
rect -3377 -4630 -3344 -4626
rect -3377 -4704 -2066 -4630
rect -9612 -5246 -7294 -5116
rect -7024 -5246 -6780 -4844
rect -6348 -4994 -4382 -4844
rect -4062 -5114 -3846 -4844
rect -3644 -4934 -3542 -4734
rect -9612 -5490 -6780 -5246
rect -6432 -5292 -4314 -5134
rect -6432 -5375 -4585 -5292
rect -4502 -5375 -4314 -5292
rect -9612 -5574 -7294 -5490
rect -6432 -5628 -4314 -5375
rect -4062 -5330 -3840 -5114
rect -9510 -5880 -7420 -5808
rect -9510 -6138 -9460 -5880
rect -7460 -6052 -7420 -5880
rect -4062 -5979 -3846 -5330
rect -3586 -5766 -3542 -4934
rect -3392 -4734 -2066 -4704
rect -3392 -4836 -1587 -4734
rect -3392 -4892 -2066 -4836
rect -3392 -5766 -3344 -4892
rect -3020 -5010 -2070 -4892
rect -2501 -5068 -2418 -5062
rect -3116 -5151 -2501 -5088
rect -2418 -5151 -1960 -5088
rect -3116 -5212 -1960 -5151
rect -3586 -5804 -3344 -5766
rect -3036 -5710 -2064 -5462
rect -1689 -5515 -1587 -4836
rect -1150 -5462 -1046 -4482
rect -294 -5515 710 -4148
rect 1376 -4286 1758 -4246
rect 1376 -5396 1470 -4286
rect 1704 -5396 1758 -4286
rect 2296 -4832 2496 -4756
rect 5403 -4832 5486 -3913
rect 5780 -4232 6770 -4210
rect 5780 -4296 5810 -4232
rect 6746 -4296 6770 -4232
rect 5780 -4316 6770 -4296
rect 7581 -4353 7664 -3913
rect 7726 -3452 8622 -3430
rect 7726 -3553 8664 -3452
rect 7726 -3741 9058 -3553
rect 7726 -3970 8664 -3741
rect 7579 -4372 7664 -4353
rect 7579 -4444 8768 -4372
rect 7577 -4534 8768 -4444
rect 7579 -4606 8768 -4534
rect 2296 -4915 2731 -4832
rect 2814 -4915 5486 -4832
rect 5764 -4714 6170 -4708
rect 5764 -4756 6674 -4714
rect 5764 -4808 5786 -4756
rect 6632 -4808 6674 -4756
rect 5764 -4894 6674 -4808
rect 2296 -4956 2496 -4915
rect 5626 -5000 5700 -4900
rect 6766 -4927 6840 -4910
rect 7579 -4916 7653 -4606
rect 7579 -4927 7588 -4916
rect 6766 -4968 7588 -4927
rect 7640 -4968 7653 -4916
rect 6766 -5001 7653 -4968
rect 6766 -5010 6840 -5001
rect 7808 -5075 8692 -4706
rect 1987 -5181 1993 -5075
rect 2099 -5088 8692 -5075
rect 2099 -5174 7834 -5088
rect 8356 -5174 8692 -5088
rect 2099 -5181 8692 -5174
rect 7808 -5198 8692 -5181
rect 8870 -5278 9058 -3741
rect 1376 -5432 1758 -5396
rect -1689 -5542 710 -5515
rect -1689 -5617 -167 -5542
rect 1492 -5710 1630 -5432
rect -3036 -5832 1630 -5710
rect 2052 -5804 2416 -5380
rect 8870 -5466 12838 -5278
rect 12586 -5724 12702 -5718
rect -3036 -5882 1610 -5832
rect 12702 -5840 12806 -5724
rect 12586 -5846 12702 -5840
rect -3036 -5930 -2064 -5882
rect -3166 -5968 -2064 -5930
rect -3612 -5979 -3509 -5978
rect -7460 -6138 -7118 -6052
rect -9510 -6168 -7118 -6138
rect -6366 -6168 -4382 -6002
rect -9510 -6186 -4382 -6168
rect -7772 -6364 -4382 -6186
rect -7772 -6392 -7118 -6364
rect -6366 -6722 -4382 -6364
rect -4062 -6082 -3451 -5979
rect -4062 -6338 -3964 -6082
rect -3464 -6085 -3451 -6082
rect -3345 -6085 -3339 -5979
rect -3166 -5984 -1780 -5968
rect -3214 -5996 -1780 -5984
rect -3214 -6006 -1632 -5996
rect -3214 -6012 -3010 -6006
rect -3464 -6322 -3406 -6085
rect -3214 -6156 -3066 -6012
rect -2102 -6028 -1632 -6006
rect -1886 -6154 -1632 -6028
rect 12788 -6168 12912 -6114
rect -3364 -6258 -3300 -6170
rect 12778 -6172 12912 -6168
rect 698 -6276 1976 -6244
rect 12778 -6256 12788 -6172
rect -2770 -6322 1976 -6276
rect 12782 -6296 12788 -6256
rect 12845 -6296 12912 -6172
rect -3464 -6328 1976 -6322
rect -3464 -6330 750 -6328
rect -4062 -6382 -3514 -6338
rect -3462 -6374 750 -6330
rect -3462 -6382 -2718 -6374
rect -4062 -6388 -3406 -6382
rect -3612 -6394 -3456 -6388
rect -3612 -6395 -3509 -6394
rect 12830 -6708 12902 -6296
rect -11346 -6820 -11314 -6746
rect -11252 -6938 12714 -6856
rect 12796 -6890 12920 -6708
rect -11252 -7014 -4006 -6938
rect -4024 -7080 -4006 -7014
rect -3464 -7014 12714 -6938
rect -3464 -7080 -3438 -7014
rect -4024 -7100 -3438 -7080
rect -3677 -7133 -3439 -7100
<< via1 >>
rect 6180 -3688 6295 -3573
rect -7515 -4583 -7392 -4460
rect -6853 -4482 -6730 -4296
rect -1706 -4453 -1577 -4324
rect -1264 -4482 -1135 -4296
rect -3504 -4583 -3377 -4577
rect -3504 -4668 -3498 -4583
rect -3498 -4668 -3383 -4583
rect -3504 -4698 -3383 -4668
rect -3383 -4698 -3377 -4583
rect -3504 -4704 -3392 -4698
rect -3392 -4704 -3377 -4698
rect -4585 -5375 -4502 -5292
rect -3519 -5711 -3433 -5625
rect -2501 -5151 -2418 -5068
rect 5810 -4296 6746 -4232
rect 2731 -4915 2814 -4832
rect 5786 -4808 6632 -4756
rect 7588 -4968 7640 -4916
rect 1993 -5181 2099 -5075
rect 12586 -5840 12702 -5724
rect -3451 -6085 -3345 -5979
rect 12788 -6296 12845 -6172
rect -3677 -7071 -3591 -6985
<< metal2 >>
rect 5320 -3688 6180 -3573
rect 6295 -3688 6301 -3573
rect -6853 -4296 -6730 -4290
rect -7515 -4450 -6853 -4327
rect -7515 -4460 -7392 -4450
rect -1264 -4296 -1135 -4290
rect -6730 -4450 -6729 -4327
rect -1712 -4453 -1706 -4324
rect -1577 -4453 -1264 -4324
rect -6853 -4488 -6730 -4482
rect -1135 -4453 -1134 -4324
rect -1264 -4488 -1135 -4482
rect -7515 -4589 -7392 -4583
rect -3514 -4577 -3366 -4564
rect -3514 -4704 -3504 -4577
rect -3377 -4582 -3366 -4577
rect 5320 -4582 5435 -3688
rect -3377 -4697 5435 -4582
rect 5768 -4232 6770 -4200
rect 5768 -4296 5810 -4232
rect 6746 -4296 6770 -4232
rect -3377 -4704 -3366 -4697
rect -3514 -4714 -3366 -4704
rect 5768 -4756 6770 -4296
rect 5768 -4808 5786 -4756
rect 6632 -4808 6770 -4756
rect 2731 -4832 2814 -4826
rect 5768 -4832 6770 -4808
rect -1843 -4915 2731 -4832
rect -1843 -5068 -1760 -4915
rect 2731 -4921 2814 -4915
rect -4445 -5151 -2501 -5068
rect -2418 -5151 -1760 -5068
rect 1993 -5075 2099 -5069
rect -4445 -5292 -4362 -5151
rect -4591 -5375 -4585 -5292
rect -4502 -5375 -4362 -5292
rect -1579 -5181 1993 -5075
rect -3677 -5711 -3519 -5625
rect -3433 -5711 -3427 -5625
rect -3677 -6985 -3591 -5711
rect -1579 -5847 -1473 -5181
rect 1993 -5187 2099 -5181
rect 6482 -5724 6598 -4832
rect 7588 -4916 7640 -4910
rect 7588 -5724 7640 -4968
rect 6482 -5840 12586 -5724
rect 12702 -5840 12708 -5724
rect -3451 -5953 -1473 -5847
rect -3451 -5979 -3345 -5953
rect -3451 -6091 -3345 -6085
rect 7588 -6208 7640 -5840
rect 12788 -6172 12845 -6166
rect 7588 -6260 12788 -6208
rect 12788 -6302 12845 -6296
rect -3683 -7071 -3677 -6985
rect -3591 -7071 -3585 -6985
use sky130_fd_pr__pfet_g5v0d16v0_KV2QNB  XM2
timestamp 1757939962
transform 0 -1 -2542 1 0 -5236
box -694 -928 694 928
use sky130_fd_pr__nfet_g5v0d16v0_KC9U4L  XM3
timestamp 1757939962
transform 0 1 8204 -1 0 -4331
box -799 -898 799 898
use sky130_fd_pr__nfet_01v8_lvt_BBNS5X  XM4
timestamp 1757939962
transform 0 1 6234 -1 0 -4951
box -211 -710 211 710
use sky130_fd_pr__pfet_01v8_lvt_4QXYT3  XM5
timestamp 1757939962
transform 0 1 8199 -1 0 -3267
box -231 -719 231 719
use sky130_fd_pr__pfet_g5v0d16v0_KV2QNB  XM6
timestamp 1757939962
transform 0 -1 6276 1 0 -3978
box -694 -928 694 928
use sky130_fd_pr__nfet_g5v0d16v0_H7ZMNC  XM7
timestamp 1757939962
transform 1 0 167 0 1 -4846
box -1649 -1028 1649 1028
use sky130_fd_pr__nfet_01v8_lvt_NFLWKG  XM11
timestamp 1757939962
transform 0 1 4738 -1 0 -6214
box -216 -8210 216 8210
use sky130_fd_pr__pfet_g5v0d16v0_DCHRLX  XM12
timestamp 1757939962
transform 0 1 -8454 -1 0 -5251
box -1019 -1508 1019 1508
use sky130_fd_pr__nfet_g5v0d16v0_D75ULX  XM13
timestamp 1757939962
transform 0 -1 -5376 1 0 -5493
box -949 -1398 949 1398
use sky130_fd_pr__pfet_01v8_lvt_X35DX6  XM14
timestamp 1757939962
transform 0 1 737 -1 0 -6784
box -246 -12219 246 12219
use sky130_fd_pr__res_xhigh_po_0p69_M8H66P  XR1
timestamp 1757939962
transform 0 1 7436 -1 0 -5777
box -235 -5582 235 5582
use sky130_fd_pr__res_xhigh_po_0p69_M8H66P  XR3
timestamp 1757939962
transform 0 1 7436 -1 0 -5413
box -235 -5582 235 5582
<< labels >>
flabel metal1 -3802 -6388 -3602 -6188 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 -3644 -4934 -3444 -4734 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -3886 -4480 -3686 -4280 0 FreeSans 256 0 0 0 O_STI_NR
port 4 nsew
flabel metal1 2094 -5712 2294 -5512 0 FreeSans 256 0 0 0 O_STI
port 3 nsew
flabel metal1 2296 -4956 2496 -4756 0 FreeSans 256 0 0 0 IN
port 1 nsew
<< end >>
