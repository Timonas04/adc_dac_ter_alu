VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.405 212.675 14.575 212.865 ;
        RECT 15.785 212.675 15.955 212.865 ;
        RECT 23.170 212.695 23.340 212.865 ;
        RECT 23.170 212.675 23.280 212.695 ;
        RECT 24.065 212.675 24.235 212.865 ;
        RECT 33.270 212.695 33.440 212.865 ;
        RECT 33.295 212.675 33.440 212.695 ;
        RECT 36.950 212.675 37.120 212.865 ;
        RECT 40.165 212.675 40.335 212.865 ;
        RECT 49.825 212.675 49.995 212.865 ;
        RECT 59.030 212.675 59.200 212.865 ;
        RECT 62.705 212.675 62.875 212.865 ;
        RECT 65.470 212.675 65.640 212.865 ;
        RECT 67.765 212.675 67.935 212.865 ;
        RECT 69.660 212.725 69.780 212.835 ;
        RECT 70.070 212.675 70.240 212.865 ;
        RECT 72.355 212.675 72.525 212.865 ;
        RECT 73.735 212.675 73.905 212.865 ;
        RECT 74.665 212.720 74.825 212.830 ;
        RECT 76.495 212.675 76.665 212.865 ;
        RECT 77.875 212.675 78.045 212.865 ;
        RECT 78.350 212.675 78.520 212.865 ;
        RECT 82.015 212.675 82.185 212.865 ;
        RECT 82.485 212.695 82.655 212.865 ;
        RECT 84.775 212.675 84.945 212.865 ;
        RECT 86.625 212.675 86.795 212.865 ;
        RECT 87.545 212.720 87.705 212.830 ;
        RECT 89.375 212.675 89.545 212.865 ;
        RECT 89.845 212.715 90.015 212.865 ;
        RECT 91.225 212.720 91.385 212.830 ;
        RECT 14.265 211.865 15.635 212.675 ;
        RECT 15.725 211.765 18.725 212.675 ;
        RECT 18.865 211.995 23.280 212.675 ;
        RECT 18.865 211.765 22.795 211.995 ;
        RECT 23.475 211.805 23.905 212.590 ;
        RECT 23.925 211.995 33.030 212.675 ;
        RECT 33.295 211.765 36.335 212.675 ;
        RECT 36.355 211.805 36.785 212.590 ;
        RECT 36.950 212.445 40.005 212.675 ;
        RECT 36.805 211.765 40.005 212.445 ;
        RECT 40.025 211.995 49.130 212.675 ;
        RECT 49.235 211.805 49.665 212.590 ;
        RECT 49.685 211.995 58.790 212.675 ;
        RECT 59.030 212.445 62.085 212.675 ;
        RECT 58.885 211.765 62.085 212.445 ;
        RECT 62.115 211.805 62.545 212.590 ;
        RECT 62.565 211.995 65.305 212.675 ;
        RECT 65.325 211.765 67.535 212.675 ;
        RECT 67.625 211.995 69.455 212.675 ;
        RECT 68.110 211.765 69.455 211.995 ;
        RECT 69.925 211.765 71.275 212.675 ;
        RECT 71.305 211.895 72.675 212.675 ;
        RECT 72.685 211.895 74.055 212.675 ;
        RECT 74.995 211.805 75.425 212.590 ;
        RECT 75.445 211.895 76.815 212.675 ;
        RECT 76.825 211.895 78.195 212.675 ;
        RECT 78.205 211.765 80.815 212.675 ;
        RECT 80.965 211.895 82.335 212.675 ;
        RECT 83.725 211.895 85.095 212.675 ;
        RECT 85.105 211.995 86.935 212.675 ;
        RECT 85.105 211.765 86.450 211.995 ;
        RECT 87.875 211.805 88.305 212.590 ;
        RECT 88.325 211.895 89.695 212.675 ;
        RECT 89.725 211.765 90.615 212.715 ;
        RECT 92.595 212.675 92.765 212.865 ;
        RECT 94.445 212.675 94.615 212.865 ;
        RECT 91.545 211.895 92.915 212.675 ;
        RECT 92.925 211.995 94.755 212.675 ;
        RECT 94.765 212.445 97.475 212.675 ;
        RECT 98.585 212.445 98.755 212.865 ;
        RECT 100.425 212.675 100.595 212.865 ;
        RECT 101.400 212.725 101.520 212.835 ;
        RECT 102.715 212.675 102.885 212.865 ;
        RECT 104.105 212.675 104.275 212.865 ;
        RECT 105.945 212.675 106.115 212.865 ;
        RECT 107.785 212.675 107.955 212.865 ;
        RECT 109.165 212.675 109.335 212.865 ;
        RECT 111.005 212.675 111.175 212.865 ;
        RECT 112.375 212.675 112.545 212.865 ;
        RECT 113.305 212.720 113.465 212.830 ;
        RECT 114.280 212.725 114.400 212.835 ;
        RECT 119.745 212.675 119.915 212.865 ;
        RECT 125.265 212.675 125.435 212.865 ;
        RECT 126.645 212.675 126.815 212.865 ;
        RECT 94.765 211.995 98.860 212.445 ;
        RECT 94.765 211.765 95.715 211.995 ;
        RECT 97.485 211.765 98.860 211.995 ;
        RECT 98.905 211.865 100.735 212.675 ;
        RECT 100.755 211.805 101.185 212.590 ;
        RECT 101.665 211.895 103.035 212.675 ;
        RECT 103.045 211.865 104.415 212.675 ;
        RECT 104.425 211.995 106.255 212.675 ;
        RECT 104.425 211.765 105.770 211.995 ;
        RECT 106.265 211.865 108.095 212.675 ;
        RECT 108.105 211.895 109.475 212.675 ;
        RECT 109.485 211.865 111.315 212.675 ;
        RECT 111.325 211.895 112.695 212.675 ;
        RECT 113.635 211.805 114.065 212.590 ;
        RECT 114.545 211.865 120.055 212.675 ;
        RECT 120.065 211.865 125.575 212.675 ;
        RECT 125.585 211.865 126.955 212.675 ;
      LAYER nwell ;
        RECT 14.070 208.645 127.150 211.475 ;
      LAYER pwell ;
        RECT 14.265 207.445 15.635 208.255 ;
        RECT 16.185 207.445 19.635 208.355 ;
        RECT 20.245 207.445 23.455 208.355 ;
        RECT 23.475 207.530 23.905 208.315 ;
        RECT 33.125 208.155 34.535 208.355 ;
        RECT 24.010 207.445 33.115 208.125 ;
        RECT 33.125 207.475 35.860 208.155 ;
        RECT 33.125 207.445 34.520 207.475 ;
        RECT 14.405 207.235 14.575 207.445 ;
        RECT 15.840 207.285 15.960 207.395 ;
        RECT 16.245 207.255 16.415 207.445 ;
        RECT 17.620 207.235 17.790 207.425 ;
        RECT 19.980 207.285 20.100 207.395 ;
        RECT 23.145 207.255 23.315 207.445 ;
        RECT 26.825 207.235 26.995 207.425 ;
        RECT 32.805 207.255 32.975 207.445 ;
        RECT 35.565 207.255 35.735 207.475 ;
        RECT 35.885 207.445 44.990 208.125 ;
        RECT 45.625 207.445 49.210 208.355 ;
        RECT 49.235 207.530 49.665 208.315 ;
        RECT 58.885 208.125 60.230 208.355 ;
        RECT 49.685 207.445 58.790 208.125 ;
        RECT 58.885 207.445 60.715 208.125 ;
        RECT 60.990 207.445 63.925 208.355 ;
        RECT 65.095 208.265 66.685 208.355 ;
        RECT 64.115 207.445 66.685 208.265 ;
        RECT 68.040 208.155 68.995 208.355 ;
        RECT 66.715 207.475 68.995 208.155 ;
        RECT 36.025 207.235 36.195 207.445 ;
        RECT 37.000 207.285 37.120 207.395 ;
        RECT 37.405 207.235 37.575 207.425 ;
        RECT 45.280 207.285 45.400 207.395 ;
        RECT 48.900 207.255 49.070 207.445 ;
        RECT 49.825 207.425 49.995 207.445 ;
        RECT 49.820 207.255 49.995 207.425 ;
        RECT 50.340 207.285 50.460 207.395 ;
        RECT 49.820 207.235 49.990 207.255 ;
        RECT 54.880 207.235 55.050 207.425 ;
        RECT 58.100 207.235 58.270 207.425 ;
        RECT 58.620 207.285 58.740 207.395 ;
        RECT 59.025 207.255 59.195 207.425 ;
        RECT 60.405 207.255 60.575 207.445 ;
        RECT 60.990 207.425 61.035 207.445 ;
        RECT 64.115 207.425 64.255 207.445 ;
        RECT 60.865 207.255 61.035 207.425 ;
        RECT 63.165 207.280 63.325 207.390 ;
        RECT 14.265 206.425 15.635 207.235 ;
        RECT 15.725 206.325 17.935 207.235 ;
        RECT 18.030 206.555 27.135 207.235 ;
        RECT 27.230 206.555 36.335 207.235 ;
        RECT 36.355 206.365 36.785 207.150 ;
        RECT 37.265 206.555 46.370 207.235 ;
        RECT 46.480 206.325 50.135 207.235 ;
        RECT 50.605 206.555 55.195 207.235 ;
        RECT 55.215 207.005 58.270 207.235 ;
        RECT 59.150 207.235 59.195 207.255 ;
        RECT 63.625 207.235 63.795 207.425 ;
        RECT 64.085 207.255 64.255 207.425 ;
        RECT 66.840 207.425 67.010 207.475 ;
        RECT 68.040 207.445 68.995 207.475 ;
        RECT 69.015 207.445 70.365 208.355 ;
        RECT 71.385 207.445 74.835 208.355 ;
        RECT 74.995 207.530 75.425 208.315 ;
        RECT 75.445 207.445 76.795 208.355 ;
        RECT 76.825 207.445 78.195 208.225 ;
        RECT 78.215 207.445 79.565 208.355 ;
        RECT 79.585 207.445 80.955 208.225 ;
        RECT 81.910 208.125 85.520 208.355 ;
        RECT 81.425 207.445 85.520 208.125 ;
        RECT 85.570 208.125 86.950 208.355 ;
        RECT 88.740 208.125 90.115 208.355 ;
        RECT 90.650 208.125 91.995 208.355 ;
        RECT 92.490 208.125 93.835 208.355 ;
        RECT 85.570 207.675 90.115 208.125 ;
        RECT 85.570 207.445 88.730 207.675 ;
        RECT 66.840 207.255 67.015 207.425 ;
        RECT 69.145 207.255 69.315 207.445 ;
        RECT 70.985 207.290 71.145 207.400 ;
        RECT 71.445 207.255 71.615 207.445 ;
        RECT 66.845 207.235 67.015 207.255 ;
        RECT 53.370 206.325 54.710 206.555 ;
        RECT 55.215 206.325 58.415 207.005 ;
        RECT 59.150 206.325 62.085 207.235 ;
        RECT 62.115 206.365 62.545 207.150 ;
        RECT 63.565 206.325 66.565 207.235 ;
        RECT 66.785 206.325 70.235 207.235 ;
        RECT 70.385 207.205 71.340 207.235 ;
        RECT 72.370 207.205 72.540 207.425 ;
        RECT 74.665 207.235 74.835 207.425 ;
        RECT 75.125 207.235 75.295 207.425 ;
        RECT 75.590 207.255 75.760 207.445 ;
        RECT 77.875 207.255 78.045 207.445 ;
        RECT 78.345 207.255 78.515 207.445 ;
        RECT 80.185 207.235 80.355 207.425 ;
        RECT 80.635 207.255 80.805 207.445 ;
        RECT 81.570 207.425 81.740 207.445 ;
        RECT 81.160 207.285 81.280 207.395 ;
        RECT 81.565 207.255 81.740 207.425 ;
        RECT 81.565 207.235 81.735 207.255 ;
        RECT 82.025 207.235 82.195 207.425 ;
        RECT 84.785 207.235 84.955 207.425 ;
        RECT 88.465 207.235 88.635 207.425 ;
        RECT 89.840 207.255 90.010 207.675 ;
        RECT 90.165 207.445 91.995 208.125 ;
        RECT 92.005 207.445 93.835 208.125 ;
        RECT 93.880 208.125 97.490 208.355 ;
        RECT 98.470 208.125 99.815 208.355 ;
        RECT 93.880 207.445 97.975 208.125 ;
        RECT 97.985 207.445 99.815 208.125 ;
        RECT 100.755 207.530 101.185 208.315 ;
        RECT 102.125 207.445 107.635 208.255 ;
        RECT 107.645 207.445 113.155 208.255 ;
        RECT 113.165 207.445 118.675 208.255 ;
        RECT 118.685 207.445 124.195 208.255 ;
        RECT 125.585 207.445 126.955 208.255 ;
        RECT 90.305 207.255 90.475 207.445 ;
        RECT 92.145 207.255 92.315 207.445 ;
        RECT 92.605 207.235 92.775 207.425 ;
        RECT 95.365 207.235 95.535 207.425 ;
        RECT 97.660 207.255 97.830 207.445 ;
        RECT 98.125 207.255 98.295 207.445 ;
        RECT 100.425 207.290 100.585 207.400 ;
        RECT 101.805 207.290 101.965 207.400 ;
        RECT 102.265 207.235 102.435 207.425 ;
        RECT 107.325 207.255 107.495 207.445 ;
        RECT 107.785 207.235 107.955 207.425 ;
        RECT 112.845 207.255 113.015 207.445 ;
        RECT 113.305 207.235 113.475 207.425 ;
        RECT 114.280 207.285 114.400 207.395 ;
        RECT 118.365 207.255 118.535 207.445 ;
        RECT 119.745 207.235 119.915 207.425 ;
        RECT 123.885 207.255 124.055 207.445 ;
        RECT 124.345 207.255 124.515 207.425 ;
        RECT 125.265 207.235 125.435 207.425 ;
        RECT 126.645 207.235 126.815 207.445 ;
        RECT 70.385 206.525 72.665 207.205 ;
        RECT 72.685 206.555 74.975 207.235 ;
        RECT 70.385 206.325 71.340 206.525 ;
        RECT 72.685 206.325 73.605 206.555 ;
        RECT 74.985 206.325 78.195 207.235 ;
        RECT 78.205 206.555 80.495 207.235 ;
        RECT 78.205 206.325 79.125 206.555 ;
        RECT 80.515 206.325 81.865 207.235 ;
        RECT 81.895 206.325 84.625 207.235 ;
        RECT 84.645 206.325 87.855 207.235 ;
        RECT 87.875 206.365 88.305 207.150 ;
        RECT 88.325 206.325 91.535 207.235 ;
        RECT 92.475 206.325 95.205 207.235 ;
        RECT 95.240 206.325 97.055 207.235 ;
        RECT 97.065 206.425 102.575 207.235 ;
        RECT 102.585 206.425 108.095 207.235 ;
        RECT 108.105 206.425 113.615 207.235 ;
        RECT 113.635 206.365 114.065 207.150 ;
        RECT 114.545 206.425 120.055 207.235 ;
        RECT 120.065 206.425 125.575 207.235 ;
        RECT 125.585 206.425 126.955 207.235 ;
      LAYER nwell ;
        RECT 14.070 203.205 127.150 206.035 ;
      LAYER pwell ;
        RECT 14.265 202.005 15.635 202.815 ;
        RECT 15.655 202.005 17.005 202.915 ;
        RECT 17.225 202.005 22.535 202.915 ;
        RECT 23.475 202.090 23.905 202.875 ;
        RECT 23.930 202.005 27.595 202.915 ;
        RECT 27.605 202.005 31.735 202.915 ;
        RECT 31.830 202.005 40.935 202.685 ;
        RECT 40.955 202.235 44.155 202.915 ;
        RECT 40.955 202.005 44.010 202.235 ;
        RECT 44.260 202.005 49.215 202.915 ;
        RECT 49.235 202.090 49.665 202.875 ;
        RECT 49.685 202.005 53.815 202.915 ;
        RECT 55.645 202.685 56.575 202.915 ;
        RECT 53.825 202.005 56.575 202.685 ;
        RECT 56.595 202.235 59.795 202.915 ;
        RECT 59.805 202.685 60.735 202.915 ;
        RECT 56.595 202.005 59.650 202.235 ;
        RECT 59.805 202.005 62.555 202.685 ;
        RECT 62.565 202.005 63.935 202.815 ;
        RECT 63.945 202.005 67.155 202.915 ;
        RECT 67.180 202.005 68.995 202.915 ;
        RECT 69.005 202.005 70.375 202.815 ;
        RECT 70.385 202.685 71.305 202.915 ;
        RECT 72.685 202.685 73.605 202.915 ;
        RECT 70.385 202.005 72.675 202.685 ;
        RECT 72.685 202.005 74.975 202.685 ;
        RECT 74.995 202.090 75.425 202.875 ;
        RECT 75.445 202.715 76.390 202.915 ;
        RECT 75.445 202.035 78.195 202.715 ;
        RECT 75.445 202.005 76.390 202.035 ;
        RECT 14.405 201.795 14.575 202.005 ;
        RECT 16.705 201.815 16.875 202.005 ;
        RECT 17.165 201.795 17.335 201.985 ;
        RECT 17.680 201.845 17.800 201.955 ;
        RECT 18.085 201.795 18.255 201.985 ;
        RECT 22.225 201.815 22.395 202.005 ;
        RECT 23.145 201.850 23.305 201.960 ;
        RECT 27.280 201.815 27.450 202.005 ;
        RECT 31.420 201.815 31.590 202.005 ;
        RECT 36.025 201.795 36.195 201.985 ;
        RECT 36.945 201.795 37.115 201.985 ;
        RECT 40.625 201.815 40.795 202.005 ;
        RECT 43.840 201.815 44.010 202.005 ;
        RECT 48.900 201.815 49.070 202.005 ;
        RECT 49.365 201.815 49.535 201.985 ;
        RECT 49.335 201.795 49.535 201.815 ;
        RECT 52.580 201.795 52.750 201.985 ;
        RECT 53.045 201.795 53.215 201.985 ;
        RECT 53.500 201.815 53.670 202.005 ;
        RECT 53.965 201.815 54.135 202.005 ;
        RECT 55.810 201.795 55.980 201.985 ;
        RECT 58.565 201.840 58.725 201.950 ;
        RECT 59.480 201.815 59.650 202.005 ;
        RECT 60.860 201.795 61.030 201.985 ;
        RECT 61.785 201.840 61.945 201.950 ;
        RECT 62.245 201.815 62.415 202.005 ;
        RECT 63.625 201.795 63.795 202.005 ;
        RECT 64.085 201.835 64.255 201.985 ;
        RECT 14.265 200.985 15.635 201.795 ;
        RECT 15.645 201.115 17.475 201.795 ;
        RECT 17.945 201.115 27.050 201.795 ;
        RECT 27.230 201.115 36.335 201.795 ;
        RECT 15.645 200.885 16.990 201.115 ;
        RECT 36.355 200.925 36.785 201.710 ;
        RECT 36.805 201.115 45.910 201.795 ;
        RECT 46.005 201.115 49.535 201.795 ;
        RECT 46.005 200.885 48.830 201.115 ;
        RECT 49.685 200.885 52.895 201.795 ;
        RECT 52.905 201.115 55.645 201.795 ;
        RECT 55.665 200.885 57.875 201.795 ;
        RECT 59.340 201.565 61.030 201.795 ;
        RECT 59.340 200.885 61.175 201.565 ;
        RECT 62.115 200.925 62.545 201.710 ;
        RECT 62.565 201.015 63.935 201.795 ;
        RECT 63.965 200.885 64.855 201.835 ;
        RECT 65.005 201.795 65.175 201.985 ;
        RECT 66.855 201.815 67.025 202.005 ;
        RECT 67.305 201.815 67.475 202.005 ;
        RECT 70.065 201.815 70.235 202.005 ;
        RECT 70.520 201.795 70.690 201.985 ;
        RECT 70.985 201.795 71.155 201.985 ;
        RECT 72.365 201.815 72.535 202.005 ;
        RECT 73.285 201.795 73.455 201.985 ;
        RECT 74.205 201.840 74.365 201.950 ;
        RECT 74.665 201.815 74.835 202.005 ;
        RECT 76.045 201.795 76.215 201.985 ;
        RECT 77.880 201.815 78.050 202.035 ;
        RECT 78.205 202.005 83.715 202.815 ;
        RECT 83.725 202.005 85.075 202.915 ;
        RECT 85.105 202.005 86.920 202.915 ;
        RECT 87.995 202.685 88.925 202.915 ;
        RECT 87.090 202.005 88.925 202.685 ;
        RECT 89.245 202.005 92.915 202.915 ;
        RECT 93.405 202.005 94.755 202.915 ;
        RECT 95.225 202.005 100.735 202.815 ;
        RECT 100.755 202.090 101.185 202.875 ;
        RECT 106.485 202.825 107.435 202.915 ;
        RECT 101.665 202.005 103.495 202.815 ;
        RECT 103.505 202.005 105.335 202.685 ;
        RECT 105.505 202.005 107.435 202.825 ;
        RECT 107.645 202.005 110.395 202.815 ;
        RECT 110.405 202.005 112.235 202.685 ;
        RECT 112.705 202.005 114.535 202.815 ;
        RECT 114.545 202.005 120.055 202.815 ;
        RECT 120.065 202.005 125.575 202.815 ;
        RECT 125.585 202.005 126.955 202.815 ;
        RECT 78.805 201.795 78.975 201.985 ;
        RECT 80.185 201.795 80.355 201.985 ;
        RECT 83.405 201.815 83.575 202.005 ;
        RECT 84.790 201.815 84.960 202.005 ;
        RECT 85.705 201.795 85.875 201.985 ;
        RECT 86.165 201.795 86.335 201.985 ;
        RECT 86.625 201.815 86.795 202.005 ;
        RECT 87.090 201.985 87.255 202.005 ;
        RECT 87.085 201.815 87.255 201.985 ;
        RECT 88.520 201.845 88.640 201.955 ;
        RECT 88.925 201.795 89.095 201.985 ;
        RECT 92.605 201.955 92.775 202.005 ;
        RECT 92.605 201.845 92.780 201.955 ;
        RECT 93.120 201.845 93.240 201.955 ;
        RECT 92.605 201.815 92.775 201.845 ;
        RECT 93.520 201.815 93.690 202.005 ;
        RECT 94.900 201.955 95.070 201.985 ;
        RECT 94.900 201.845 95.080 201.955 ;
        RECT 94.900 201.795 95.070 201.845 ;
        RECT 95.370 201.795 95.540 201.985 ;
        RECT 96.800 201.845 96.920 201.955 ;
        RECT 99.505 201.795 99.675 201.985 ;
        RECT 99.955 201.795 100.125 201.985 ;
        RECT 100.425 201.815 100.595 202.005 ;
        RECT 103.185 201.955 103.355 202.005 ;
        RECT 101.400 201.845 101.520 201.955 ;
        RECT 103.185 201.845 103.360 201.955 ;
        RECT 103.185 201.815 103.355 201.845 ;
        RECT 103.645 201.815 103.815 202.005 ;
        RECT 105.505 201.985 105.655 202.005 ;
        RECT 105.485 201.815 105.655 201.985 ;
        RECT 105.945 201.795 106.115 201.985 ;
        RECT 108.705 201.795 108.875 201.985 ;
        RECT 110.085 201.815 110.255 202.005 ;
        RECT 110.545 201.815 110.715 202.005 ;
        RECT 111.920 201.795 112.090 201.985 ;
        RECT 112.440 201.845 112.560 201.955 ;
        RECT 113.305 201.795 113.475 201.985 ;
        RECT 114.225 201.955 114.395 202.005 ;
        RECT 114.225 201.845 114.400 201.955 ;
        RECT 114.225 201.815 114.395 201.845 ;
        RECT 119.745 201.795 119.915 202.005 ;
        RECT 125.265 201.795 125.435 202.005 ;
        RECT 126.645 201.795 126.815 202.005 ;
        RECT 64.880 200.885 66.695 201.795 ;
        RECT 67.180 200.885 70.835 201.795 ;
        RECT 70.855 200.885 72.205 201.795 ;
        RECT 72.225 201.015 73.595 201.795 ;
        RECT 74.525 200.885 76.340 201.795 ;
        RECT 76.375 200.885 79.105 201.795 ;
        RECT 79.125 200.985 80.495 201.795 ;
        RECT 80.505 200.985 86.015 201.795 ;
        RECT 86.025 201.115 87.855 201.795 ;
        RECT 86.510 200.885 87.855 201.115 ;
        RECT 87.875 200.925 88.305 201.710 ;
        RECT 88.785 200.885 92.455 201.795 ;
        RECT 93.380 201.565 95.070 201.795 ;
        RECT 93.380 200.885 95.215 201.565 ;
        RECT 95.225 200.885 96.575 201.795 ;
        RECT 97.065 200.985 99.815 201.795 ;
        RECT 99.825 200.885 103.035 201.795 ;
        RECT 103.505 200.985 106.255 201.795 ;
        RECT 106.265 201.115 109.015 201.795 ;
        RECT 109.025 201.115 112.235 201.795 ;
        RECT 106.265 200.885 107.195 201.115 ;
        RECT 109.025 200.885 110.390 201.115 ;
        RECT 112.245 200.985 113.615 201.795 ;
        RECT 113.635 200.925 114.065 201.710 ;
        RECT 114.545 200.985 120.055 201.795 ;
        RECT 120.065 200.985 125.575 201.795 ;
        RECT 125.585 200.985 126.955 201.795 ;
      LAYER nwell ;
        RECT 14.070 197.765 127.150 200.595 ;
      LAYER pwell ;
        RECT 14.265 196.565 15.635 197.375 ;
        RECT 15.645 196.795 18.395 197.475 ;
        RECT 15.785 196.565 18.395 196.795 ;
        RECT 18.410 196.795 23.455 197.475 ;
        RECT 18.410 196.565 23.315 196.795 ;
        RECT 23.475 196.650 23.905 197.435 ;
        RECT 25.730 197.275 26.675 197.475 ;
        RECT 23.925 196.595 26.675 197.275 ;
        RECT 14.405 196.355 14.575 196.565 ;
        RECT 15.785 196.375 15.955 196.565 ;
        RECT 23.145 196.375 23.315 196.565 ;
        RECT 24.070 196.375 24.240 196.595 ;
        RECT 25.730 196.565 26.675 196.595 ;
        RECT 26.920 196.565 31.735 197.245 ;
        RECT 31.830 196.565 40.935 197.245 ;
        RECT 40.965 196.565 42.315 197.475 ;
        RECT 42.325 196.565 46.400 197.475 ;
        RECT 47.805 197.275 49.215 197.475 ;
        RECT 46.480 196.595 49.215 197.275 ;
        RECT 49.235 196.650 49.665 197.435 ;
        RECT 24.525 196.355 24.695 196.545 ;
        RECT 24.985 196.355 25.155 196.545 ;
        RECT 26.825 196.400 26.985 196.510 ;
        RECT 31.425 196.375 31.595 196.565 ;
        RECT 36.025 196.355 36.195 196.545 ;
        RECT 37.865 196.355 38.035 196.545 ;
        RECT 40.625 196.375 40.795 196.565 ;
        RECT 41.080 196.375 41.250 196.565 ;
        RECT 45.225 196.355 45.395 196.545 ;
        RECT 46.170 196.510 46.340 196.565 ;
        RECT 46.145 196.400 46.340 196.510 ;
        RECT 46.170 196.375 46.340 196.400 ;
        RECT 46.605 196.375 46.775 196.595 ;
        RECT 47.820 196.565 49.215 196.595 ;
        RECT 49.685 196.565 51.055 197.345 ;
        RECT 51.065 196.565 54.275 197.475 ;
        RECT 54.295 196.565 55.645 197.475 ;
        RECT 55.665 196.565 58.875 197.475 ;
        RECT 49.825 196.545 49.995 196.565 ;
        RECT 49.820 196.375 49.995 196.545 ;
        RECT 49.820 196.355 49.990 196.375 ;
        RECT 50.285 196.355 50.455 196.545 ;
        RECT 51.205 196.375 51.375 196.565 ;
        RECT 52.180 196.405 52.300 196.515 ;
        RECT 54.425 196.375 54.595 196.565 ;
        RECT 55.805 196.545 55.975 196.565 ;
        RECT 55.800 196.375 55.975 196.545 ;
        RECT 55.800 196.355 55.970 196.375 ;
        RECT 56.265 196.355 56.435 196.545 ;
        RECT 58.885 196.525 59.775 197.475 ;
        RECT 60.290 197.245 61.635 197.475 ;
        RECT 59.805 196.565 61.635 197.245 ;
        RECT 61.645 196.565 63.015 197.345 ;
        RECT 63.025 196.565 64.395 197.345 ;
        RECT 64.405 196.565 65.775 197.345 ;
        RECT 66.245 196.565 67.615 197.345 ;
        RECT 67.625 196.565 69.455 197.245 ;
        RECT 70.585 196.565 74.975 197.475 ;
        RECT 74.995 196.650 75.425 197.435 ;
        RECT 75.445 196.565 77.275 197.245 ;
        RECT 78.205 196.565 83.715 197.375 ;
        RECT 83.725 196.565 89.235 197.375 ;
        RECT 89.265 196.565 90.615 197.475 ;
        RECT 92.470 197.245 93.835 197.475 ;
        RECT 90.625 196.565 93.835 197.245 ;
        RECT 93.845 196.565 97.055 197.475 ;
        RECT 97.065 196.565 100.735 197.475 ;
        RECT 100.755 196.650 101.185 197.435 ;
        RECT 102.450 196.565 106.105 197.475 ;
        RECT 107.185 196.565 110.395 197.475 ;
        RECT 110.415 196.565 113.145 197.475 ;
        RECT 113.165 196.565 114.535 197.375 ;
        RECT 114.545 196.565 118.215 197.375 ;
        RECT 118.225 196.565 123.735 197.375 ;
        RECT 123.745 196.565 125.575 197.245 ;
        RECT 125.585 196.565 126.955 197.375 ;
        RECT 59.485 196.375 59.660 196.525 ;
        RECT 59.945 196.375 60.115 196.565 ;
        RECT 62.705 196.375 62.875 196.565 ;
        RECT 64.075 196.375 64.245 196.565 ;
        RECT 59.490 196.355 59.660 196.375 ;
        RECT 14.265 195.545 15.635 196.355 ;
        RECT 15.730 195.675 24.835 196.355 ;
        RECT 24.855 195.445 26.205 196.355 ;
        RECT 27.230 195.675 36.335 196.355 ;
        RECT 36.355 195.485 36.785 196.270 ;
        RECT 36.815 195.445 38.165 196.355 ;
        RECT 38.625 195.445 45.535 196.355 ;
        RECT 46.660 195.445 50.135 196.355 ;
        RECT 50.160 195.445 51.975 196.355 ;
        RECT 52.530 195.675 56.115 196.355 ;
        RECT 55.195 195.445 56.115 195.675 ;
        RECT 56.125 195.445 59.335 196.355 ;
        RECT 59.345 195.445 62.095 196.355 ;
        RECT 62.565 196.325 63.510 196.355 ;
        RECT 65.000 196.325 65.170 196.545 ;
        RECT 65.455 196.515 65.625 196.565 ;
        RECT 65.925 196.515 66.095 196.545 ;
        RECT 65.455 196.405 65.640 196.515 ;
        RECT 65.925 196.405 66.100 196.515 ;
        RECT 65.455 196.375 65.625 196.405 ;
        RECT 65.925 196.395 66.095 196.405 ;
        RECT 62.115 195.485 62.545 196.270 ;
        RECT 62.565 195.645 65.315 196.325 ;
        RECT 62.565 195.445 63.510 195.645 ;
        RECT 65.805 195.445 66.695 196.395 ;
        RECT 66.845 196.355 67.015 196.545 ;
        RECT 67.295 196.375 67.465 196.565 ;
        RECT 68.740 196.405 68.860 196.515 ;
        RECT 69.145 196.375 69.315 196.565 ;
        RECT 70.065 196.410 70.225 196.520 ;
        RECT 70.525 196.355 70.695 196.545 ;
        RECT 71.445 196.400 71.605 196.510 ;
        RECT 74.660 196.375 74.830 196.565 ;
        RECT 75.125 196.355 75.295 196.545 ;
        RECT 76.965 196.375 77.135 196.565 ;
        RECT 77.425 196.375 77.595 196.545 ;
        RECT 77.885 196.410 78.045 196.520 ;
        RECT 77.425 196.355 77.590 196.375 ;
        RECT 80.645 196.355 80.815 196.545 ;
        RECT 83.405 196.375 83.575 196.565 ;
        RECT 84.320 196.355 84.490 196.545 ;
        RECT 84.840 196.405 84.960 196.515 ;
        RECT 87.545 196.355 87.715 196.545 ;
        RECT 88.925 196.375 89.095 196.565 ;
        RECT 89.385 196.355 89.555 196.545 ;
        RECT 90.300 196.375 90.470 196.565 ;
        RECT 90.770 196.355 90.940 196.565 ;
        RECT 91.280 196.405 91.400 196.515 ;
        RECT 93.985 196.375 94.155 196.565 ;
        RECT 94.440 196.355 94.610 196.545 ;
        RECT 94.960 196.405 95.080 196.515 ;
        RECT 96.745 196.355 96.915 196.545 ;
        RECT 100.420 196.375 100.590 196.565 ;
        RECT 105.945 196.545 106.105 196.565 ;
        RECT 101.805 196.410 101.965 196.520 ;
        RECT 102.265 196.355 102.435 196.545 ;
        RECT 104.565 196.375 104.735 196.545 ;
        RECT 105.945 196.375 106.115 196.545 ;
        RECT 104.565 196.355 104.730 196.375 ;
        RECT 106.405 196.355 106.575 196.545 ;
        RECT 106.865 196.410 107.025 196.520 ;
        RECT 107.315 196.375 107.485 196.565 ;
        RECT 109.165 196.355 109.335 196.545 ;
        RECT 110.545 196.375 110.715 196.565 ;
        RECT 111.465 196.375 111.635 196.545 ;
        RECT 111.465 196.355 111.615 196.375 ;
        RECT 113.305 196.355 113.475 196.545 ;
        RECT 114.225 196.375 114.395 196.565 ;
        RECT 115.605 196.355 115.775 196.545 ;
        RECT 117.905 196.375 118.075 196.565 ;
        RECT 121.125 196.355 121.295 196.545 ;
        RECT 121.585 196.355 121.755 196.545 ;
        RECT 123.425 196.375 123.595 196.565 ;
        RECT 123.885 196.355 124.055 196.545 ;
        RECT 125.265 196.375 125.435 196.565 ;
        RECT 126.645 196.355 126.815 196.565 ;
        RECT 66.720 195.445 68.535 196.355 ;
        RECT 69.005 195.445 70.820 196.355 ;
        RECT 71.765 195.545 75.435 196.355 ;
        RECT 75.755 195.675 77.590 196.355 ;
        RECT 75.755 195.445 76.685 195.675 ;
        RECT 78.175 195.445 80.955 196.355 ;
        RECT 81.160 195.445 84.635 196.355 ;
        RECT 85.105 195.545 87.855 196.355 ;
        RECT 87.875 195.485 88.305 196.270 ;
        RECT 88.325 195.545 89.695 196.355 ;
        RECT 89.705 195.445 91.055 196.355 ;
        RECT 91.555 196.125 94.610 196.355 ;
        RECT 91.555 195.445 94.755 196.125 ;
        RECT 95.225 195.545 97.055 196.355 ;
        RECT 97.065 195.545 102.575 196.355 ;
        RECT 102.895 195.675 104.730 196.355 ;
        RECT 104.885 195.675 106.715 196.355 ;
        RECT 102.895 195.445 103.825 195.675 ;
        RECT 104.885 195.445 106.230 195.675 ;
        RECT 106.725 195.445 109.475 196.355 ;
        RECT 109.685 195.535 111.615 196.355 ;
        RECT 111.785 195.545 113.615 196.355 ;
        RECT 109.685 195.445 110.635 195.535 ;
        RECT 113.635 195.485 114.065 196.270 ;
        RECT 114.085 195.545 115.915 196.355 ;
        RECT 115.925 195.545 121.435 196.355 ;
        RECT 121.445 195.575 122.815 196.355 ;
        RECT 123.745 195.675 125.575 196.355 ;
        RECT 124.230 195.445 125.575 195.675 ;
        RECT 125.585 195.545 126.955 196.355 ;
      LAYER nwell ;
        RECT 14.070 192.325 127.150 195.155 ;
      LAYER pwell ;
        RECT 14.265 191.125 15.635 191.935 ;
        RECT 15.645 191.125 19.315 192.035 ;
        RECT 19.335 191.805 20.680 192.035 ;
        RECT 19.335 191.125 23.360 191.805 ;
        RECT 23.475 191.210 23.905 191.995 ;
        RECT 24.845 191.125 28.715 192.035 ;
        RECT 28.985 191.125 32.100 192.035 ;
        RECT 32.665 191.125 35.415 191.935 ;
        RECT 35.425 191.125 44.530 191.805 ;
        RECT 44.625 191.125 47.835 192.035 ;
        RECT 47.855 191.125 49.205 192.035 ;
        RECT 49.235 191.210 49.665 191.995 ;
        RECT 49.685 191.125 51.035 192.035 ;
        RECT 51.390 191.125 55.045 192.035 ;
        RECT 55.665 191.125 58.415 192.035 ;
        RECT 58.445 191.125 59.795 192.035 ;
        RECT 60.265 191.805 63.090 192.035 ;
        RECT 63.945 191.805 66.770 192.035 ;
        RECT 60.265 191.125 63.795 191.805 ;
        RECT 63.945 191.125 67.475 191.805 ;
        RECT 68.560 191.125 72.215 192.035 ;
        RECT 72.240 191.125 74.055 192.035 ;
        RECT 74.995 191.210 75.425 191.995 ;
        RECT 76.655 191.125 79.575 192.035 ;
        RECT 79.585 191.835 80.530 192.035 ;
        RECT 81.865 191.835 82.795 192.035 ;
        RECT 79.585 191.355 82.795 191.835 ;
        RECT 83.265 191.805 84.190 192.035 ;
        RECT 79.585 191.155 82.655 191.355 ;
        RECT 79.585 191.125 80.530 191.155 ;
        RECT 14.405 190.915 14.575 191.125 ;
        RECT 15.790 190.935 15.960 191.125 ;
        RECT 17.165 190.915 17.335 191.105 ;
        RECT 17.680 190.965 17.800 191.075 ;
        RECT 19.445 190.935 19.615 191.125 ;
        RECT 24.525 190.970 24.685 191.080 ;
        RECT 24.990 190.935 25.160 191.125 ;
        RECT 26.825 190.915 26.995 191.105 ;
        RECT 29.130 190.935 29.300 191.125 ;
        RECT 32.400 190.965 32.520 191.075 ;
        RECT 35.105 190.935 35.275 191.125 ;
        RECT 35.565 190.935 35.735 191.125 ;
        RECT 36.025 190.915 36.195 191.105 ;
        RECT 37.870 190.915 38.040 191.105 ;
        RECT 38.330 190.915 38.500 191.105 ;
        RECT 44.770 190.935 44.940 191.125 ;
        RECT 45.685 190.915 45.855 191.105 ;
        RECT 46.150 190.915 46.320 191.105 ;
        RECT 47.525 190.915 47.695 191.105 ;
        RECT 47.985 190.935 48.155 191.125 ;
        RECT 49.830 190.935 50.000 191.125 ;
        RECT 54.885 191.105 55.045 191.125 ;
        RECT 54.885 190.935 55.055 191.105 ;
        RECT 55.400 190.965 55.520 191.075 ;
        RECT 55.810 190.935 55.980 191.125 ;
        RECT 56.725 190.915 56.895 191.105 ;
        RECT 58.560 190.935 58.730 191.125 ;
        RECT 63.595 191.105 63.795 191.125 ;
        RECT 67.275 191.105 67.475 191.125 ;
        RECT 71.900 191.105 72.070 191.125 ;
        RECT 59.950 190.915 60.120 191.105 ;
        RECT 61.785 190.960 61.945 191.070 ;
        RECT 63.625 190.915 63.795 191.105 ;
        RECT 64.085 190.955 64.255 191.105 ;
        RECT 65.465 190.960 65.625 191.070 ;
        RECT 14.265 190.105 15.635 190.915 ;
        RECT 15.645 190.235 17.475 190.915 ;
        RECT 18.030 190.235 27.135 190.915 ;
        RECT 27.230 190.235 36.335 190.915 ;
        RECT 15.645 190.005 16.990 190.235 ;
        RECT 36.355 190.045 36.785 190.830 ;
        RECT 36.805 190.005 38.155 190.915 ;
        RECT 38.185 190.005 42.315 190.915 ;
        RECT 42.325 190.105 45.995 190.915 ;
        RECT 46.005 190.005 47.355 190.915 ;
        RECT 47.385 190.235 56.490 190.915 ;
        RECT 56.585 190.005 59.795 190.915 ;
        RECT 59.805 190.005 61.155 190.915 ;
        RECT 62.115 190.045 62.545 190.830 ;
        RECT 62.565 190.135 63.935 190.915 ;
        RECT 63.965 190.005 64.855 190.955 ;
        RECT 67.305 190.915 67.475 191.105 ;
        RECT 67.740 190.915 67.910 191.105 ;
        RECT 68.225 190.970 68.385 191.080 ;
        RECT 71.900 190.935 72.075 191.105 ;
        RECT 72.365 190.935 72.535 191.125 ;
        RECT 74.665 190.970 74.825 191.080 ;
        RECT 76.045 190.970 76.205 191.080 ;
        RECT 71.905 190.915 72.075 190.935 ;
        RECT 76.505 190.915 76.675 191.105 ;
        RECT 76.960 190.915 77.130 191.105 ;
        RECT 78.345 190.915 78.515 191.105 ;
        RECT 79.260 190.935 79.430 191.125 ;
        RECT 82.485 190.935 82.655 191.155 ;
        RECT 83.265 191.125 86.935 191.805 ;
        RECT 86.945 191.125 89.695 191.935 ;
        RECT 89.705 191.125 95.215 191.935 ;
        RECT 95.225 191.125 100.735 191.935 ;
        RECT 100.755 191.210 101.185 191.995 ;
        RECT 105.545 191.945 106.495 192.035 ;
        RECT 101.665 191.125 105.335 191.935 ;
        RECT 105.545 191.125 107.475 191.945 ;
        RECT 107.645 191.835 108.575 192.035 ;
        RECT 109.905 191.835 110.855 192.035 ;
        RECT 107.645 191.355 110.855 191.835 ;
        RECT 113.630 191.805 114.970 192.035 ;
        RECT 83.000 190.965 83.120 191.075 ;
        RECT 83.410 190.935 83.580 191.125 ;
        RECT 65.785 190.005 67.600 190.915 ;
        RECT 67.680 190.005 71.755 190.915 ;
        RECT 71.765 190.005 74.975 190.915 ;
        RECT 74.985 190.105 76.815 190.915 ;
        RECT 76.845 190.005 78.195 190.915 ;
        RECT 78.215 190.005 80.945 190.915 ;
        RECT 80.965 190.885 81.910 190.915 ;
        RECT 83.865 190.885 84.035 191.105 ;
        RECT 84.785 190.960 84.945 191.070 ;
        RECT 87.545 190.915 87.715 191.105 ;
        RECT 88.520 190.965 88.640 191.075 ;
        RECT 89.385 190.935 89.555 191.125 ;
        RECT 92.145 190.915 92.315 191.105 ;
        RECT 93.525 190.915 93.695 191.105 ;
        RECT 94.040 190.965 94.160 191.075 ;
        RECT 94.905 190.935 95.075 191.125 ;
        RECT 99.505 190.915 99.675 191.105 ;
        RECT 99.965 190.915 100.135 191.105 ;
        RECT 100.425 190.935 100.595 191.125 ;
        RECT 101.400 190.965 101.520 191.075 ;
        RECT 102.265 190.960 102.425 191.070 ;
        RECT 102.725 190.915 102.895 191.105 ;
        RECT 105.025 190.935 105.195 191.125 ;
        RECT 107.325 191.105 107.475 191.125 ;
        RECT 107.790 191.155 110.855 191.355 ;
        RECT 107.325 190.935 107.495 191.105 ;
        RECT 107.790 190.935 107.960 191.155 ;
        RECT 109.920 191.125 110.855 191.155 ;
        RECT 110.865 191.125 115.455 191.805 ;
        RECT 115.925 191.125 121.435 191.935 ;
        RECT 121.445 191.125 122.815 191.905 ;
        RECT 123.745 191.125 125.575 191.805 ;
        RECT 125.585 191.125 126.955 191.935 ;
        RECT 109.625 190.915 109.795 191.105 ;
        RECT 113.305 190.915 113.475 191.105 ;
        RECT 115.140 190.935 115.310 191.125 ;
        RECT 115.660 190.965 115.780 191.075 ;
        RECT 116.525 190.935 116.695 191.105 ;
        RECT 116.525 190.915 116.665 190.935 ;
        RECT 119.285 190.915 119.455 191.105 ;
        RECT 121.125 190.935 121.295 191.125 ;
        RECT 121.585 190.935 121.755 191.125 ;
        RECT 122.500 190.915 122.670 191.105 ;
        RECT 123.425 190.970 123.585 191.080 ;
        RECT 123.885 190.915 124.055 191.105 ;
        RECT 125.265 190.915 125.435 191.125 ;
        RECT 126.645 190.915 126.815 191.125 ;
        RECT 80.965 190.685 84.035 190.885 ;
        RECT 80.965 190.205 84.175 190.685 ;
        RECT 80.965 190.005 81.910 190.205 ;
        RECT 83.245 190.005 84.175 190.205 ;
        RECT 85.105 190.235 87.855 190.915 ;
        RECT 85.105 190.005 86.035 190.235 ;
        RECT 87.875 190.045 88.305 190.830 ;
        RECT 88.785 190.105 92.455 190.915 ;
        RECT 92.475 190.005 93.825 190.915 ;
        RECT 94.305 190.105 99.815 190.915 ;
        RECT 99.840 190.005 101.655 190.915 ;
        RECT 102.665 190.005 106.115 190.915 ;
        RECT 106.265 190.105 109.935 190.915 ;
        RECT 109.945 190.235 113.615 190.915 ;
        RECT 109.945 190.005 110.875 190.235 ;
        RECT 113.635 190.045 114.065 190.830 ;
        RECT 114.095 190.095 116.665 190.915 ;
        RECT 116.845 190.235 119.595 190.915 ;
        RECT 119.605 190.235 122.815 190.915 ;
        RECT 114.095 190.005 115.685 190.095 ;
        RECT 116.845 190.005 117.775 190.235 ;
        RECT 119.605 190.005 120.970 190.235 ;
        RECT 122.835 190.005 124.185 190.915 ;
        RECT 124.205 190.105 125.575 190.915 ;
        RECT 125.585 190.105 126.955 190.915 ;
      LAYER nwell ;
        RECT 14.070 186.885 127.150 189.715 ;
      LAYER pwell ;
        RECT 14.265 185.685 15.635 186.495 ;
        RECT 15.645 185.685 19.190 186.595 ;
        RECT 19.325 185.685 23.455 186.595 ;
        RECT 23.475 185.770 23.905 186.555 ;
        RECT 23.935 185.685 26.675 186.365 ;
        RECT 26.685 185.685 28.055 186.465 ;
        RECT 28.065 185.685 29.415 186.595 ;
        RECT 29.905 185.685 33.575 186.495 ;
        RECT 33.585 185.685 34.935 186.595 ;
        RECT 35.050 185.685 44.155 186.365 ;
        RECT 44.165 185.685 47.375 186.595 ;
        RECT 47.385 185.685 49.215 186.365 ;
        RECT 49.235 185.770 49.665 186.555 ;
        RECT 49.695 185.685 51.045 186.595 ;
        RECT 51.065 185.685 52.435 186.465 ;
        RECT 53.495 186.365 54.425 186.595 ;
        RECT 52.590 185.685 54.425 186.365 ;
        RECT 54.745 185.685 57.955 186.595 ;
        RECT 57.965 185.685 67.070 186.365 ;
        RECT 67.165 185.685 70.375 186.595 ;
        RECT 71.305 185.685 74.975 186.495 ;
        RECT 74.995 185.770 75.425 186.555 ;
        RECT 75.905 185.685 77.735 186.495 ;
        RECT 77.745 185.685 83.255 186.495 ;
        RECT 86.015 186.365 86.935 186.595 ;
        RECT 83.350 185.685 86.935 186.365 ;
        RECT 86.945 186.365 87.875 186.595 ;
        RECT 86.945 185.685 89.695 186.365 ;
        RECT 90.165 185.685 91.995 186.495 ;
        RECT 92.005 185.685 97.515 186.495 ;
        RECT 97.545 185.685 98.895 186.595 ;
        RECT 98.905 185.685 100.720 186.595 ;
        RECT 100.755 185.770 101.185 186.555 ;
        RECT 101.205 185.685 105.325 186.595 ;
        RECT 105.360 185.685 107.175 186.595 ;
        RECT 107.185 185.685 109.935 186.495 ;
        RECT 109.945 185.685 111.295 186.595 ;
        RECT 111.325 186.395 112.275 186.595 ;
        RECT 113.605 186.395 114.535 186.595 ;
        RECT 111.325 185.915 114.535 186.395 ;
        RECT 111.325 185.715 114.390 185.915 ;
        RECT 111.325 185.685 112.260 185.715 ;
        RECT 14.405 185.475 14.575 185.685 ;
        RECT 15.790 185.495 15.960 185.685 ;
        RECT 16.245 185.475 16.415 185.665 ;
        RECT 17.680 185.525 17.800 185.635 ;
        RECT 23.140 185.495 23.310 185.685 ;
        RECT 26.365 185.495 26.535 185.685 ;
        RECT 26.825 185.475 26.995 185.665 ;
        RECT 27.285 185.475 27.455 185.665 ;
        RECT 27.745 185.495 27.915 185.685 ;
        RECT 29.130 185.495 29.300 185.685 ;
        RECT 29.640 185.525 29.760 185.635 ;
        RECT 33.265 185.495 33.435 185.685 ;
        RECT 33.730 185.495 33.900 185.685 ;
        RECT 40.160 185.475 40.330 185.665 ;
        RECT 43.385 185.475 43.555 185.665 ;
        RECT 43.845 185.475 44.015 185.685 ;
        RECT 44.305 185.495 44.475 185.685 ;
        RECT 47.525 185.495 47.695 185.685 ;
        RECT 48.905 185.475 49.075 185.665 ;
        RECT 49.825 185.495 49.995 185.685 ;
        RECT 50.285 185.495 50.455 185.665 ;
        RECT 51.215 185.495 51.385 185.685 ;
        RECT 52.590 185.665 52.755 185.685 ;
        RECT 14.265 184.665 15.635 185.475 ;
        RECT 16.105 184.695 17.475 185.475 ;
        RECT 18.030 184.795 27.135 185.475 ;
        RECT 27.145 184.795 36.250 185.475 ;
        RECT 36.355 184.605 36.785 185.390 ;
        RECT 36.805 184.795 40.475 185.475 ;
        RECT 36.805 184.565 38.395 184.795 ;
        RECT 40.485 184.565 43.695 185.475 ;
        RECT 43.705 184.795 46.445 185.475 ;
        RECT 46.465 185.245 49.075 185.475 ;
        RECT 50.305 185.475 50.455 185.495 ;
        RECT 46.465 184.565 49.215 185.245 ;
        RECT 50.305 184.655 52.235 185.475 ;
        RECT 52.585 185.445 52.755 185.665 ;
        RECT 54.885 185.495 55.055 185.685 ;
        RECT 57.185 185.475 57.355 185.665 ;
        RECT 57.645 185.515 57.815 185.665 ;
        RECT 58.105 185.515 58.275 185.685 ;
        RECT 54.745 185.445 56.115 185.475 ;
        RECT 52.445 184.765 56.115 185.445 ;
        RECT 51.285 184.565 52.235 184.655 ;
        RECT 54.730 184.565 56.115 184.765 ;
        RECT 56.125 184.695 57.495 185.475 ;
        RECT 57.525 184.565 58.415 185.515 ;
        RECT 61.780 185.475 61.950 185.665 ;
        RECT 63.165 185.520 63.325 185.630 ;
        RECT 63.620 185.475 63.790 185.665 ;
        RECT 67.310 185.495 67.480 185.685 ;
        RECT 67.765 185.475 67.935 185.665 ;
        RECT 70.985 185.475 71.155 185.665 ;
        RECT 72.820 185.475 72.990 185.665 ;
        RECT 74.665 185.475 74.835 185.685 ;
        RECT 75.640 185.525 75.760 185.635 ;
        RECT 77.425 185.495 77.595 185.685 ;
        RECT 80.185 185.475 80.355 185.665 ;
        RECT 80.650 185.475 80.820 185.665 ;
        RECT 82.945 185.495 83.115 185.685 ;
        RECT 86.620 185.495 86.790 185.685 ;
        RECT 87.540 185.475 87.710 185.665 ;
        RECT 88.465 185.475 88.635 185.665 ;
        RECT 89.385 185.495 89.555 185.685 ;
        RECT 89.900 185.525 90.020 185.635 ;
        RECT 90.310 185.475 90.480 185.665 ;
        RECT 91.685 185.495 91.855 185.685 ;
        RECT 97.205 185.665 97.375 185.685 ;
        RECT 93.980 185.475 94.150 185.665 ;
        RECT 94.445 185.495 94.615 185.665 ;
        RECT 96.800 185.525 96.920 185.635 ;
        RECT 94.465 185.475 94.615 185.495 ;
        RECT 97.200 185.495 97.375 185.665 ;
        RECT 98.580 185.495 98.750 185.685 ;
        RECT 100.425 185.495 100.595 185.685 ;
        RECT 101.345 185.495 101.515 185.685 ;
        RECT 101.810 185.495 101.980 185.665 ;
        RECT 103.185 185.495 103.355 185.685 ;
        RECT 105.485 185.665 105.655 185.685 ;
        RECT 105.485 185.495 105.670 185.665 ;
        RECT 97.200 185.475 97.370 185.495 ;
        RECT 101.810 185.475 101.945 185.495 ;
        RECT 105.500 185.475 105.670 185.495 ;
        RECT 108.245 185.475 108.415 185.665 ;
        RECT 109.625 185.475 109.795 185.685 ;
        RECT 110.090 185.495 110.260 185.685 ;
        RECT 111.460 185.475 111.630 185.665 ;
        RECT 113.305 185.475 113.475 185.665 ;
        RECT 114.220 185.495 114.390 185.715 ;
        RECT 114.545 185.685 118.215 186.495 ;
        RECT 118.225 185.685 123.735 186.495 ;
        RECT 124.230 186.365 125.575 186.595 ;
        RECT 123.745 185.685 125.575 186.365 ;
        RECT 125.585 185.685 126.955 186.495 ;
        RECT 115.600 185.475 115.770 185.665 ;
        RECT 116.985 185.475 117.155 185.665 ;
        RECT 117.905 185.495 118.075 185.685 ;
        RECT 120.665 185.475 120.835 185.665 ;
        RECT 123.425 185.495 123.595 185.685 ;
        RECT 123.885 185.495 124.055 185.685 ;
        RECT 125.290 185.495 125.460 185.665 ;
        RECT 125.290 185.475 125.400 185.495 ;
        RECT 126.645 185.475 126.815 185.685 ;
        RECT 58.425 184.565 62.095 185.475 ;
        RECT 62.115 184.605 62.545 185.390 ;
        RECT 63.505 184.565 64.855 185.475 ;
        RECT 64.995 184.565 67.995 185.475 ;
        RECT 68.215 184.565 71.215 185.475 ;
        RECT 71.305 184.565 73.135 185.475 ;
        RECT 73.145 184.665 74.975 185.475 ;
        RECT 74.985 184.665 80.495 185.475 ;
        RECT 80.505 184.565 84.160 185.475 ;
        RECT 84.185 184.565 87.855 185.475 ;
        RECT 87.875 184.605 88.305 185.390 ;
        RECT 88.340 184.565 90.155 185.475 ;
        RECT 90.165 184.795 92.440 185.475 ;
        RECT 91.070 184.565 92.440 184.795 ;
        RECT 92.465 184.565 94.295 185.475 ;
        RECT 94.465 184.655 96.395 185.475 ;
        RECT 95.445 184.565 96.395 184.655 ;
        RECT 97.085 184.565 98.435 185.475 ;
        RECT 98.445 184.565 101.945 185.475 ;
        RECT 102.125 184.565 105.785 185.475 ;
        RECT 105.805 184.665 108.555 185.475 ;
        RECT 108.575 184.565 109.925 185.475 ;
        RECT 109.945 184.565 111.775 185.475 ;
        RECT 111.785 184.795 113.615 185.475 ;
        RECT 111.785 184.565 113.130 184.795 ;
        RECT 113.635 184.605 114.065 185.390 ;
        RECT 114.085 184.565 115.915 185.475 ;
        RECT 115.925 184.665 117.295 185.475 ;
        RECT 117.305 184.665 120.975 185.475 ;
        RECT 120.985 184.795 125.400 185.475 ;
        RECT 120.985 184.565 124.915 184.795 ;
        RECT 125.585 184.665 126.955 185.475 ;
      LAYER nwell ;
        RECT 14.070 181.445 127.150 184.275 ;
      LAYER pwell ;
        RECT 14.265 180.245 15.635 181.055 ;
        RECT 16.105 180.245 17.475 181.025 ;
        RECT 17.625 180.245 21.075 181.155 ;
        RECT 21.245 180.245 23.455 181.155 ;
        RECT 23.475 180.330 23.905 181.115 ;
        RECT 24.385 180.245 25.755 181.025 ;
        RECT 25.795 180.245 29.895 181.155 ;
        RECT 29.905 180.475 35.380 181.155 ;
        RECT 29.905 180.245 33.995 180.475 ;
        RECT 14.405 180.035 14.575 180.245 ;
        RECT 15.840 180.085 15.960 180.195 ;
        RECT 16.245 180.055 16.415 180.245 ;
        RECT 17.155 180.035 17.325 180.225 ;
        RECT 17.625 180.035 17.795 180.225 ;
        RECT 20.845 180.055 21.015 180.245 ;
        RECT 21.765 180.080 21.925 180.190 ;
        RECT 22.225 180.035 22.395 180.225 ;
        RECT 23.140 180.055 23.310 180.245 ;
        RECT 24.120 180.085 24.240 180.195 ;
        RECT 24.535 180.055 24.705 180.245 ;
        RECT 29.580 180.055 29.750 180.245 ;
        RECT 31.425 180.035 31.595 180.225 ;
        RECT 35.105 180.055 35.275 180.475 ;
        RECT 35.425 180.245 38.635 181.155 ;
        RECT 38.645 180.245 41.855 181.155 ;
        RECT 41.865 180.245 45.075 181.155 ;
        RECT 45.105 180.245 46.455 181.155 ;
        RECT 46.485 180.245 47.835 181.155 ;
        RECT 47.845 180.245 49.215 181.025 ;
        RECT 49.235 180.330 49.665 181.115 ;
        RECT 49.685 180.245 51.035 181.155 ;
        RECT 52.310 180.245 55.965 181.155 ;
        RECT 56.125 180.245 57.495 181.025 ;
        RECT 35.565 180.055 35.735 180.245 ;
        RECT 36.020 180.035 36.190 180.225 ;
        RECT 38.790 180.055 38.960 180.245 ;
        RECT 40.160 180.035 40.330 180.225 ;
        RECT 42.465 180.055 42.635 180.225 ;
        RECT 42.465 180.035 42.630 180.055 ;
        RECT 42.935 180.035 43.105 180.225 ;
        RECT 44.315 180.035 44.485 180.225 ;
        RECT 44.765 180.055 44.935 180.245 ;
        RECT 45.220 180.055 45.390 180.245 ;
        RECT 46.600 180.225 46.770 180.245 ;
        RECT 46.600 180.055 46.775 180.225 ;
        RECT 46.605 180.035 46.775 180.055 ;
        RECT 47.065 180.035 47.235 180.225 ;
        RECT 48.445 180.035 48.615 180.225 ;
        RECT 48.895 180.055 49.065 180.245 ;
        RECT 49.830 180.035 50.000 180.245 ;
        RECT 55.805 180.225 55.965 180.245 ;
        RECT 51.665 180.090 51.825 180.200 ;
        RECT 52.115 180.035 52.285 180.225 ;
        RECT 55.345 180.035 55.515 180.225 ;
        RECT 55.805 180.055 55.975 180.225 ;
        RECT 56.265 180.080 56.425 180.190 ;
        RECT 57.175 180.055 57.345 180.245 ;
        RECT 57.525 180.205 58.415 181.155 ;
        RECT 58.425 180.245 62.095 181.155 ;
        RECT 62.565 180.245 68.075 181.055 ;
        RECT 68.085 180.245 69.435 181.155 ;
        RECT 69.465 180.245 71.295 181.055 ;
        RECT 71.305 180.245 73.135 181.155 ;
        RECT 73.605 180.245 74.955 181.155 ;
        RECT 74.995 180.330 75.425 181.115 ;
        RECT 75.445 180.245 76.815 181.055 ;
        RECT 76.825 180.245 82.335 181.055 ;
        RECT 82.375 180.245 85.095 181.155 ;
        RECT 85.105 180.925 86.240 181.155 ;
        RECT 85.105 180.245 88.315 180.925 ;
        RECT 88.325 180.245 89.695 181.055 ;
        RECT 89.705 180.245 93.375 181.055 ;
        RECT 93.385 180.245 98.895 181.055 ;
        RECT 98.925 180.245 100.275 181.155 ;
        RECT 100.755 180.330 101.185 181.115 ;
        RECT 101.675 180.245 103.025 181.155 ;
        RECT 103.965 180.245 107.635 181.055 ;
        RECT 107.655 180.245 109.005 181.155 ;
        RECT 109.025 180.475 110.860 181.155 ;
        RECT 114.525 180.925 115.455 181.155 ;
        RECT 109.170 180.245 110.860 180.475 ;
        RECT 111.555 180.245 115.455 180.925 ;
        RECT 116.385 180.245 120.055 181.055 ;
        RECT 120.065 180.245 125.575 181.055 ;
        RECT 125.585 180.245 126.955 181.055 ;
        RECT 61.780 180.225 61.950 180.245 ;
        RECT 57.645 180.055 57.815 180.205 ;
        RECT 59.025 180.035 59.195 180.225 ;
        RECT 61.780 180.055 61.955 180.225 ;
        RECT 62.300 180.085 62.420 180.195 ;
        RECT 61.785 180.035 61.955 180.055 ;
        RECT 66.110 180.035 66.280 180.225 ;
        RECT 67.120 180.035 67.290 180.225 ;
        RECT 67.765 180.055 67.935 180.245 ;
        RECT 69.150 180.055 69.320 180.245 ;
        RECT 70.985 180.055 71.155 180.245 ;
        RECT 72.820 180.225 72.990 180.245 ;
        RECT 71.445 180.080 71.605 180.190 ;
        RECT 72.820 180.055 73.000 180.225 ;
        RECT 73.340 180.085 73.460 180.195 ;
        RECT 74.670 180.055 74.840 180.245 ;
        RECT 76.505 180.225 76.675 180.245 ;
        RECT 76.500 180.055 76.675 180.225 ;
        RECT 77.020 180.085 77.140 180.195 ;
        RECT 72.830 180.035 73.000 180.055 ;
        RECT 76.500 180.035 76.670 180.055 ;
        RECT 81.130 180.035 81.300 180.225 ;
        RECT 81.620 180.085 81.740 180.195 ;
        RECT 82.025 180.055 82.195 180.245 ;
        RECT 84.785 180.225 84.955 180.245 ;
        RECT 84.325 180.035 84.495 180.225 ;
        RECT 84.785 180.055 84.960 180.225 ;
        RECT 88.005 180.055 88.175 180.245 ;
        RECT 89.385 180.225 89.555 180.245 ;
        RECT 88.925 180.080 89.085 180.190 ;
        RECT 89.380 180.055 89.555 180.225 ;
        RECT 84.790 180.035 84.960 180.055 ;
        RECT 89.380 180.035 89.550 180.055 ;
        RECT 92.145 180.035 92.315 180.225 ;
        RECT 93.065 180.055 93.235 180.245 ;
        RECT 96.010 180.035 96.180 180.225 ;
        RECT 97.665 180.035 97.835 180.225 ;
        RECT 98.125 180.035 98.295 180.225 ;
        RECT 98.585 180.055 98.755 180.245 ;
        RECT 99.040 180.055 99.210 180.245 ;
        RECT 100.480 180.085 100.600 180.195 ;
        RECT 100.885 180.035 101.055 180.225 ;
        RECT 101.400 180.085 101.520 180.195 ;
        RECT 102.725 180.055 102.895 180.245 ;
        RECT 103.185 180.080 103.345 180.190 ;
        RECT 103.640 180.035 103.810 180.225 ;
        RECT 105.080 180.085 105.200 180.195 ;
        RECT 106.410 180.035 106.580 180.225 ;
        RECT 107.325 180.055 107.495 180.245 ;
        RECT 107.785 180.055 107.955 180.245 ;
        RECT 109.170 180.225 109.340 180.245 ;
        RECT 109.165 180.055 109.340 180.225 ;
        RECT 109.165 180.035 109.305 180.055 ;
        RECT 113.030 180.035 113.200 180.225 ;
        RECT 114.870 180.055 115.040 180.245 ;
        RECT 116.065 180.090 116.225 180.200 ;
        RECT 116.985 180.035 117.155 180.225 ;
        RECT 119.745 180.035 119.915 180.245 ;
        RECT 125.265 180.035 125.435 180.245 ;
        RECT 126.645 180.035 126.815 180.245 ;
        RECT 14.265 179.225 15.635 180.035 ;
        RECT 16.105 179.255 17.475 180.035 ;
        RECT 17.565 179.125 21.015 180.035 ;
        RECT 22.085 179.355 31.190 180.035 ;
        RECT 31.285 179.255 32.655 180.035 ;
        RECT 32.680 179.125 36.335 180.035 ;
        RECT 36.355 179.165 36.785 179.950 ;
        RECT 36.805 179.125 40.475 180.035 ;
        RECT 40.795 179.355 42.630 180.035 ;
        RECT 40.795 179.125 41.725 179.355 ;
        RECT 42.785 179.255 44.155 180.035 ;
        RECT 44.165 179.255 45.535 180.035 ;
        RECT 45.545 179.255 46.915 180.035 ;
        RECT 46.935 179.125 48.285 180.035 ;
        RECT 48.315 179.125 49.665 180.035 ;
        RECT 49.685 179.125 51.035 180.035 ;
        RECT 51.065 179.255 52.435 180.035 ;
        RECT 52.445 179.125 55.655 180.035 ;
        RECT 56.585 179.125 59.335 180.035 ;
        RECT 59.345 179.225 62.095 180.035 ;
        RECT 62.115 179.165 62.545 179.950 ;
        RECT 62.795 179.355 66.695 180.035 ;
        RECT 65.765 179.125 66.695 179.355 ;
        RECT 66.705 179.355 70.605 180.035 ;
        RECT 66.705 179.125 67.635 179.355 ;
        RECT 71.765 179.125 73.115 180.035 ;
        RECT 73.145 179.355 76.815 180.035 ;
        RECT 75.890 179.125 76.815 179.355 ;
        RECT 77.285 179.125 81.360 180.035 ;
        RECT 81.885 179.225 84.635 180.035 ;
        RECT 84.645 179.125 87.565 180.035 ;
        RECT 87.875 179.165 88.305 179.950 ;
        RECT 89.265 179.125 90.615 180.035 ;
        RECT 90.625 179.225 92.455 180.035 ;
        RECT 92.695 179.355 96.595 180.035 ;
        RECT 95.665 179.125 96.595 179.355 ;
        RECT 96.605 179.225 97.975 180.035 ;
        RECT 97.995 179.125 100.725 180.035 ;
        RECT 100.760 179.125 102.575 180.035 ;
        RECT 103.525 179.125 104.875 180.035 ;
        RECT 105.345 179.125 106.695 180.035 ;
        RECT 106.735 179.215 109.305 180.035 ;
        RECT 109.715 179.355 113.615 180.035 ;
        RECT 106.735 179.125 108.325 179.215 ;
        RECT 112.685 179.125 113.615 179.355 ;
        RECT 113.635 179.165 114.065 179.950 ;
        RECT 114.085 179.125 117.295 180.035 ;
        RECT 117.305 179.225 120.055 180.035 ;
        RECT 120.065 179.225 125.575 180.035 ;
        RECT 125.585 179.225 126.955 180.035 ;
      LAYER nwell ;
        RECT 14.070 176.005 127.150 178.835 ;
      LAYER pwell ;
        RECT 14.265 174.805 15.635 175.615 ;
        RECT 15.645 175.485 16.990 175.715 ;
        RECT 15.645 174.805 17.475 175.485 ;
        RECT 17.565 174.805 21.015 175.715 ;
        RECT 22.085 174.805 23.455 175.585 ;
        RECT 23.475 174.890 23.905 175.675 ;
        RECT 25.260 174.805 26.215 175.485 ;
        RECT 26.585 174.805 32.655 175.715 ;
        RECT 33.125 174.805 42.230 175.485 ;
        RECT 42.345 174.805 43.695 175.715 ;
        RECT 43.705 174.805 47.375 175.715 ;
        RECT 47.855 174.805 49.205 175.715 ;
        RECT 49.235 174.890 49.665 175.675 ;
        RECT 50.605 174.805 52.420 175.715 ;
        RECT 52.445 174.805 55.655 175.715 ;
        RECT 56.600 174.805 58.415 175.715 ;
        RECT 59.355 174.805 62.085 175.715 ;
        RECT 62.105 174.805 63.935 175.615 ;
        RECT 67.145 175.485 68.075 175.715 ;
        RECT 71.285 175.485 72.215 175.715 ;
        RECT 64.175 174.805 68.075 175.485 ;
        RECT 68.315 174.805 72.215 175.485 ;
        RECT 72.225 174.805 74.975 175.615 ;
        RECT 74.995 174.890 75.425 175.675 ;
        RECT 75.445 174.805 78.195 175.615 ;
        RECT 78.495 174.805 82.795 175.715 ;
        RECT 82.815 174.805 85.545 175.715 ;
        RECT 86.505 174.805 87.855 175.715 ;
        RECT 91.525 175.485 92.455 175.715 ;
        RECT 95.665 175.485 96.595 175.715 ;
        RECT 88.555 174.805 92.455 175.485 ;
        RECT 92.695 174.805 96.595 175.485 ;
        RECT 96.605 174.805 99.815 175.715 ;
        RECT 100.755 174.890 101.185 175.675 ;
        RECT 101.515 175.485 102.445 175.715 ;
        RECT 103.815 175.485 104.745 175.715 ;
        RECT 101.515 174.805 103.350 175.485 ;
        RECT 103.815 174.805 105.650 175.485 ;
        RECT 105.805 174.805 108.555 175.615 ;
        RECT 111.765 175.485 112.695 175.715 ;
        RECT 108.795 174.805 112.695 175.485 ;
        RECT 113.165 174.805 115.915 175.615 ;
        RECT 115.925 174.805 121.435 175.615 ;
        RECT 121.445 174.805 122.815 175.585 ;
        RECT 122.825 174.805 125.575 175.615 ;
        RECT 125.585 174.805 126.955 175.615 ;
        RECT 14.405 174.595 14.575 174.805 ;
        RECT 17.165 174.595 17.335 174.805 ;
        RECT 17.625 174.615 17.795 174.805 ;
        RECT 20.845 174.595 21.015 174.785 ;
        RECT 21.765 174.650 21.925 174.760 ;
        RECT 22.235 174.615 22.405 174.805 ;
        RECT 32.340 174.785 32.510 174.805 ;
        RECT 22.685 174.595 22.855 174.785 ;
        RECT 23.200 174.645 23.320 174.755 ;
        RECT 24.525 174.650 24.685 174.760 ;
        RECT 24.985 174.615 25.155 174.785 ;
        RECT 32.340 174.615 32.515 174.785 ;
        RECT 32.860 174.645 32.980 174.755 ;
        RECT 33.265 174.615 33.435 174.805 ;
        RECT 43.380 174.785 43.550 174.805 ;
        RECT 33.725 174.615 33.895 174.785 ;
        RECT 37.000 174.645 37.120 174.755 ;
        RECT 32.345 174.595 32.515 174.615 ;
        RECT 33.755 174.595 33.895 174.615 ;
        RECT 37.405 174.595 37.575 174.785 ;
        RECT 38.785 174.615 38.955 174.785 ;
        RECT 38.805 174.595 38.955 174.615 ;
        RECT 42.920 174.595 43.090 174.785 ;
        RECT 43.380 174.615 43.560 174.785 ;
        RECT 43.850 174.615 44.020 174.805 ;
        RECT 47.580 174.645 47.700 174.755 ;
        RECT 48.905 174.615 49.075 174.805 ;
        RECT 49.365 174.640 49.525 174.750 ;
        RECT 50.285 174.650 50.445 174.760 ;
        RECT 43.390 174.595 43.560 174.615 ;
        RECT 50.745 174.595 50.915 174.785 ;
        RECT 51.210 174.595 51.380 174.785 ;
        RECT 52.125 174.615 52.295 174.805 ;
        RECT 52.585 174.615 52.755 174.805 ;
        RECT 53.505 174.595 53.675 174.785 ;
        RECT 55.805 174.615 55.975 174.785 ;
        RECT 56.265 174.755 56.425 174.760 ;
        RECT 56.265 174.650 56.440 174.755 ;
        RECT 56.320 174.645 56.440 174.650 ;
        RECT 56.725 174.615 56.895 174.805 ;
        RECT 59.025 174.650 59.185 174.760 ;
        RECT 55.805 174.595 55.955 174.615 ;
        RECT 14.265 173.785 15.635 174.595 ;
        RECT 15.645 173.685 17.460 174.595 ;
        RECT 17.625 173.685 21.075 174.595 ;
        RECT 21.165 173.915 22.995 174.595 ;
        RECT 23.550 173.915 32.655 174.595 ;
        RECT 21.165 173.685 22.510 173.915 ;
        RECT 33.755 173.775 36.325 174.595 ;
        RECT 34.735 173.685 36.325 173.775 ;
        RECT 36.355 173.725 36.785 174.510 ;
        RECT 37.265 173.815 38.635 174.595 ;
        RECT 38.805 173.775 40.735 174.595 ;
        RECT 39.785 173.685 40.735 173.775 ;
        RECT 41.045 173.685 43.235 174.595 ;
        RECT 43.245 173.685 48.375 174.595 ;
        RECT 49.685 173.815 51.055 174.595 ;
        RECT 51.065 173.685 52.415 174.595 ;
        RECT 52.455 173.685 53.805 174.595 ;
        RECT 54.025 173.775 55.955 174.595 ;
        RECT 56.730 174.595 56.895 174.615 ;
        RECT 60.865 174.615 61.035 174.785 ;
        RECT 61.785 174.615 61.955 174.805 ;
        RECT 60.865 174.595 61.015 174.615 ;
        RECT 63.625 174.595 63.795 174.805 ;
        RECT 65.005 174.595 65.175 174.785 ;
        RECT 65.520 174.645 65.640 174.755 ;
        RECT 65.930 174.595 66.100 174.785 ;
        RECT 67.490 174.615 67.660 174.805 ;
        RECT 70.525 174.595 70.695 174.785 ;
        RECT 70.985 174.615 71.155 174.785 ;
        RECT 71.630 174.615 71.800 174.805 ;
        RECT 74.665 174.615 74.835 174.805 ;
        RECT 70.990 174.595 71.155 174.615 ;
        RECT 76.500 174.595 76.670 174.785 ;
        RECT 77.885 174.595 78.055 174.805 ;
        RECT 78.350 174.595 78.520 174.785 ;
        RECT 81.565 174.595 81.735 174.785 ;
        RECT 82.480 174.615 82.650 174.805 ;
        RECT 82.945 174.595 83.115 174.805 ;
        RECT 84.785 174.595 84.955 174.785 ;
        RECT 86.165 174.650 86.325 174.760 ;
        RECT 86.620 174.615 86.790 174.805 ;
        RECT 87.545 174.595 87.715 174.785 ;
        RECT 88.060 174.645 88.180 174.755 ;
        RECT 88.520 174.645 88.640 174.755 ;
        RECT 90.305 174.595 90.475 174.785 ;
        RECT 90.765 174.595 90.935 174.785 ;
        RECT 91.870 174.615 92.040 174.805 ;
        RECT 96.010 174.595 96.180 174.805 ;
        RECT 99.505 174.595 99.675 174.805 ;
        RECT 103.185 174.785 103.350 174.805 ;
        RECT 105.485 174.785 105.650 174.805 ;
        RECT 100.425 174.650 100.585 174.760 ;
        RECT 101.345 174.595 101.515 174.785 ;
        RECT 101.805 174.595 101.975 174.785 ;
        RECT 103.185 174.615 103.355 174.785 ;
        RECT 103.700 174.645 103.820 174.755 ;
        RECT 105.485 174.595 105.655 174.785 ;
        RECT 105.945 174.615 106.115 174.785 ;
        RECT 108.245 174.615 108.415 174.805 ;
        RECT 105.950 174.595 106.115 174.615 ;
        RECT 111.650 174.595 111.820 174.785 ;
        RECT 112.110 174.615 112.280 174.805 ;
        RECT 112.900 174.645 113.020 174.755 ;
        RECT 113.305 174.595 113.475 174.785 ;
        RECT 115.605 174.595 115.775 174.805 ;
        RECT 121.125 174.595 121.295 174.805 ;
        RECT 121.585 174.595 121.755 174.805 ;
        RECT 123.425 174.640 123.585 174.750 ;
        RECT 123.885 174.595 124.055 174.785 ;
        RECT 125.265 174.615 125.435 174.805 ;
        RECT 126.645 174.595 126.815 174.805 ;
        RECT 56.730 173.915 58.565 174.595 ;
        RECT 54.025 173.685 54.975 173.775 ;
        RECT 57.635 173.685 58.565 173.915 ;
        RECT 59.085 173.775 61.015 174.595 ;
        RECT 59.085 173.685 60.035 173.775 ;
        RECT 62.115 173.725 62.545 174.510 ;
        RECT 62.565 173.815 63.935 174.595 ;
        RECT 63.955 173.685 65.305 174.595 ;
        RECT 65.785 173.685 67.975 174.595 ;
        RECT 68.085 173.785 70.835 174.595 ;
        RECT 70.990 173.915 72.825 174.595 ;
        RECT 73.145 173.915 76.815 174.595 ;
        RECT 71.895 173.685 72.825 173.915 ;
        RECT 75.890 173.685 76.815 173.915 ;
        RECT 76.825 173.785 78.195 174.595 ;
        RECT 78.205 173.685 81.415 174.595 ;
        RECT 81.425 173.815 82.795 174.595 ;
        RECT 82.820 173.685 84.635 174.595 ;
        RECT 84.645 173.915 86.475 174.595 ;
        RECT 85.130 173.685 86.475 173.915 ;
        RECT 86.485 173.785 87.855 174.595 ;
        RECT 87.875 173.725 88.305 174.510 ;
        RECT 88.785 173.785 90.615 174.595 ;
        RECT 90.625 173.915 92.455 174.595 ;
        RECT 92.695 173.915 96.595 174.595 ;
        RECT 95.665 173.685 96.595 173.915 ;
        RECT 96.605 173.685 99.815 174.595 ;
        RECT 99.825 173.685 101.640 174.595 ;
        RECT 101.680 173.685 103.495 174.595 ;
        RECT 103.965 173.785 105.795 174.595 ;
        RECT 105.950 173.915 107.785 174.595 ;
        RECT 108.335 173.915 112.235 174.595 ;
        RECT 106.855 173.685 107.785 173.915 ;
        RECT 111.305 173.685 112.235 173.915 ;
        RECT 112.245 173.785 113.615 174.595 ;
        RECT 113.635 173.725 114.065 174.510 ;
        RECT 114.085 173.785 115.915 174.595 ;
        RECT 115.925 173.785 121.435 174.595 ;
        RECT 121.445 173.815 122.815 174.595 ;
        RECT 123.745 173.915 125.575 174.595 ;
        RECT 124.230 173.685 125.575 173.915 ;
        RECT 125.585 173.785 126.955 174.595 ;
      LAYER nwell ;
        RECT 14.070 170.565 127.150 173.395 ;
      LAYER pwell ;
        RECT 14.265 169.365 15.635 170.175 ;
        RECT 15.645 169.365 17.935 170.275 ;
        RECT 18.025 169.365 21.025 170.275 ;
        RECT 21.625 170.045 22.970 170.275 ;
        RECT 21.625 169.365 23.455 170.045 ;
        RECT 23.475 169.450 23.905 170.235 ;
        RECT 23.925 169.365 26.675 170.275 ;
        RECT 26.685 169.365 28.055 170.145 ;
        RECT 28.065 169.365 29.435 170.145 ;
        RECT 29.455 169.365 30.805 170.275 ;
        RECT 30.835 170.185 32.425 170.275 ;
        RECT 30.835 169.365 33.405 170.185 ;
        RECT 34.070 170.045 35.415 170.275 ;
        RECT 33.585 169.365 35.415 170.045 ;
        RECT 36.355 169.450 36.785 170.235 ;
        RECT 37.005 170.185 37.955 170.275 ;
        RECT 37.005 169.365 38.935 170.185 ;
        RECT 40.155 170.045 41.085 170.275 ;
        RECT 14.405 169.175 14.575 169.365 ;
        RECT 17.625 169.175 17.795 169.365 ;
        RECT 18.085 169.175 18.255 169.365 ;
        RECT 21.360 169.205 21.480 169.315 ;
        RECT 23.145 169.175 23.315 169.365 ;
        RECT 24.065 169.175 24.235 169.365 ;
        RECT 26.835 169.175 27.005 169.365 ;
        RECT 28.205 169.175 28.375 169.365 ;
        RECT 29.585 169.175 29.755 169.365 ;
        RECT 33.265 169.345 33.405 169.365 ;
        RECT 33.265 169.175 33.435 169.345 ;
        RECT 33.725 169.175 33.895 169.365 ;
        RECT 38.785 169.345 38.935 169.365 ;
        RECT 39.250 169.365 41.085 170.045 ;
        RECT 41.865 169.365 43.235 170.145 ;
        RECT 43.730 170.045 45.075 170.275 ;
        RECT 43.245 169.365 45.075 170.045 ;
        RECT 45.085 169.365 46.455 170.145 ;
        RECT 46.950 170.045 48.295 170.275 ;
        RECT 46.465 169.365 48.295 170.045 ;
        RECT 49.235 169.450 49.665 170.235 ;
        RECT 50.170 170.045 51.515 170.275 ;
        RECT 49.685 169.365 51.515 170.045 ;
        RECT 51.525 169.365 52.895 170.145 ;
        RECT 53.365 169.365 54.735 170.145 ;
        RECT 54.745 169.365 56.115 170.145 ;
        RECT 56.125 170.045 57.470 170.275 ;
        RECT 56.125 169.365 57.955 170.045 ;
        RECT 57.965 169.365 59.335 170.145 ;
        RECT 60.265 170.045 61.610 170.275 ;
        RECT 60.265 169.365 62.095 170.045 ;
        RECT 62.115 169.450 62.545 170.235 ;
        RECT 63.025 170.045 66.955 170.275 ;
        RECT 63.025 169.365 67.440 170.045 ;
        RECT 67.625 169.365 68.995 170.145 ;
        RECT 39.250 169.345 39.415 169.365 ;
        RECT 36.025 169.210 36.185 169.320 ;
        RECT 38.785 169.175 38.955 169.345 ;
        RECT 39.245 169.175 39.415 169.345 ;
        RECT 41.600 169.205 41.720 169.315 ;
        RECT 42.005 169.175 42.175 169.365 ;
        RECT 43.385 169.175 43.555 169.365 ;
        RECT 45.235 169.175 45.405 169.365 ;
        RECT 46.605 169.175 46.775 169.365 ;
        RECT 48.905 169.210 49.065 169.320 ;
        RECT 49.825 169.175 49.995 169.365 ;
        RECT 52.575 169.175 52.745 169.365 ;
        RECT 53.100 169.205 53.220 169.315 ;
        RECT 53.515 169.175 53.685 169.365 ;
        RECT 55.795 169.175 55.965 169.365 ;
        RECT 57.645 169.175 57.815 169.365 ;
        RECT 59.025 169.175 59.195 169.365 ;
        RECT 59.945 169.210 60.105 169.320 ;
        RECT 61.785 169.175 61.955 169.365 ;
        RECT 67.330 169.345 67.440 169.365 ;
        RECT 62.760 169.205 62.880 169.315 ;
        RECT 67.330 169.175 67.500 169.345 ;
        RECT 68.675 169.175 68.845 169.365 ;
        RECT 69.025 169.325 69.915 170.275 ;
        RECT 69.925 169.365 71.295 170.145 ;
        RECT 71.305 169.365 72.675 170.175 ;
        RECT 72.685 169.365 74.055 170.145 ;
        RECT 74.995 169.450 75.425 170.235 ;
        RECT 75.905 169.365 77.275 170.145 ;
        RECT 78.205 169.365 81.875 170.175 ;
        RECT 82.370 170.045 83.715 170.275 ;
        RECT 81.885 169.365 83.715 170.045 ;
        RECT 83.725 169.365 85.555 170.175 ;
        RECT 85.565 169.365 86.935 170.145 ;
        RECT 87.875 169.450 88.305 170.235 ;
        RECT 88.325 169.365 89.695 170.175 ;
        RECT 89.705 169.365 95.215 170.175 ;
        RECT 95.225 169.365 100.735 170.175 ;
        RECT 100.755 169.450 101.185 170.235 ;
        RECT 101.665 169.365 104.415 170.175 ;
        RECT 104.425 169.365 109.935 170.175 ;
        RECT 109.945 169.365 113.155 170.275 ;
        RECT 113.635 169.450 114.065 170.235 ;
        RECT 114.085 169.365 116.835 170.175 ;
        RECT 116.845 169.365 122.355 170.175 ;
        RECT 124.230 170.045 125.575 170.275 ;
        RECT 123.745 169.365 125.575 170.045 ;
        RECT 125.585 169.365 126.955 170.175 ;
        RECT 69.145 169.175 69.315 169.325 ;
        RECT 70.975 169.175 71.145 169.365 ;
        RECT 72.365 169.175 72.535 169.365 ;
        RECT 72.835 169.175 73.005 169.365 ;
        RECT 74.665 169.210 74.825 169.320 ;
        RECT 75.640 169.205 75.760 169.315 ;
        RECT 76.955 169.175 77.125 169.365 ;
        RECT 77.885 169.210 78.045 169.320 ;
        RECT 81.565 169.175 81.735 169.365 ;
        RECT 82.025 169.175 82.195 169.365 ;
        RECT 85.245 169.175 85.415 169.365 ;
        RECT 86.615 169.175 86.785 169.365 ;
        RECT 87.545 169.210 87.705 169.320 ;
        RECT 89.385 169.175 89.555 169.365 ;
        RECT 94.905 169.175 95.075 169.365 ;
        RECT 100.425 169.175 100.595 169.365 ;
        RECT 101.400 169.205 101.520 169.315 ;
        RECT 104.105 169.175 104.275 169.365 ;
        RECT 109.625 169.175 109.795 169.365 ;
        RECT 110.085 169.175 110.255 169.365 ;
        RECT 113.360 169.205 113.480 169.315 ;
        RECT 116.525 169.175 116.695 169.365 ;
        RECT 122.045 169.175 122.215 169.365 ;
        RECT 122.505 169.175 122.675 169.345 ;
        RECT 123.885 169.175 124.055 169.365 ;
        RECT 126.645 169.175 126.815 169.365 ;
        RECT 1.290 52.730 13.780 58.190 ;
        RECT 46.010 57.320 50.180 69.810 ;
      LAYER nwell ;
        RECT 50.300 61.620 52.410 69.810 ;
      LAYER pwell ;
        RECT 50.280 57.325 52.390 61.425 ;
        RECT 52.475 57.335 58.465 69.825 ;
      LAYER nwell ;
        RECT 58.595 61.635 60.705 69.825 ;
      LAYER pwell ;
        RECT 58.585 57.325 60.695 61.425 ;
        RECT 60.805 57.325 66.795 69.815 ;
      LAYER nwell ;
        RECT 66.910 61.625 69.020 69.815 ;
      LAYER pwell ;
        RECT 66.845 57.325 68.955 61.425 ;
        RECT 69.100 57.315 75.090 69.805 ;
      LAYER nwell ;
        RECT 75.290 61.725 77.400 69.915 ;
      LAYER pwell ;
        RECT 75.265 57.345 77.375 61.445 ;
        RECT 77.545 57.330 83.535 69.820 ;
      LAYER nwell ;
        RECT 83.680 61.650 85.790 69.840 ;
      LAYER pwell ;
        RECT 83.615 57.325 85.725 61.425 ;
        RECT 85.875 57.330 91.865 69.820 ;
      LAYER nwell ;
        RECT 92.010 61.675 94.120 69.865 ;
      LAYER pwell ;
        RECT 92.000 57.320 94.110 61.420 ;
        RECT 94.205 57.330 100.195 69.820 ;
      LAYER nwell ;
        RECT 100.305 61.690 102.415 69.880 ;
      LAYER pwell ;
        RECT 100.240 57.330 102.350 61.430 ;
        RECT 102.510 57.325 108.500 69.815 ;
      LAYER nwell ;
        RECT 108.605 61.670 110.715 69.860 ;
      LAYER pwell ;
        RECT 108.605 57.330 110.715 61.430 ;
        RECT 110.810 57.335 114.980 69.825 ;
      LAYER nwell ;
        RECT 128.225 66.205 135.075 75.125 ;
        RECT 126.190 63.015 135.075 66.205 ;
        RECT 128.225 62.935 135.075 63.015 ;
      LAYER pwell ;
        RECT 128.225 62.895 135.075 62.900 ;
        RECT 126.190 59.795 135.075 62.895 ;
        RECT 128.225 56.800 135.075 59.795 ;
        RECT 1.290 50.380 31.720 52.730 ;
        RECT 43.310 50.380 61.780 52.730 ;
        RECT 67.310 50.380 85.780 52.730 ;
      LAYER nwell ;
        RECT 27.290 49.600 29.790 49.880 ;
        RECT 55.790 49.600 58.290 49.880 ;
        RECT 83.290 49.600 85.790 49.880 ;
        RECT 111.790 49.600 114.290 49.880 ;
        RECT 5.410 49.355 12.800 49.585 ;
        RECT 1.290 47.890 12.800 49.355 ;
        RECT 26.050 49.355 29.790 49.600 ;
        RECT 33.410 49.355 40.800 49.585 ;
        RECT 26.050 47.890 40.800 49.355 ;
        RECT 54.050 49.355 58.290 49.600 ;
        RECT 61.410 49.355 68.800 49.585 ;
        RECT 54.050 47.890 68.800 49.355 ;
        RECT 82.050 49.355 85.790 49.600 ;
        RECT 89.410 49.355 96.800 49.585 ;
        RECT 82.050 47.890 96.800 49.355 ;
        RECT 110.050 49.355 114.290 49.600 ;
        RECT 117.410 49.355 124.800 49.585 ;
        RECT 110.050 47.890 124.800 49.355 ;
        RECT 1.290 45.580 21.135 47.890 ;
        RECT 26.050 45.595 49.135 47.890 ;
        RECT 54.050 45.595 77.135 47.890 ;
        RECT 82.050 45.595 105.135 47.890 ;
        RECT 110.050 45.595 133.135 47.890 ;
        RECT 138.050 45.595 140.160 49.600 ;
        RECT 24.025 45.580 49.135 45.595 ;
        RECT 52.025 45.580 77.135 45.595 ;
        RECT 80.025 45.580 105.135 45.595 ;
        RECT 108.025 45.580 133.135 45.595 ;
        RECT 136.025 45.580 140.160 45.595 ;
        RECT 1.290 39.410 140.160 45.580 ;
      LAYER pwell ;
        RECT 143.290 44.730 149.800 50.190 ;
        RECT 143.290 40.560 155.780 44.730 ;
      LAYER nwell ;
        RECT 1.290 39.405 26.135 39.410 ;
        RECT 27.440 39.405 54.135 39.410 ;
        RECT 55.790 39.405 82.135 39.410 ;
        RECT 84.280 39.405 110.135 39.410 ;
        RECT 111.790 39.405 138.135 39.410 ;
        RECT 1.290 39.395 24.110 39.405 ;
        RECT 12.720 39.390 24.110 39.395 ;
        RECT 27.545 39.395 52.110 39.405 ;
        RECT 27.545 39.390 29.790 39.395 ;
        RECT 40.720 39.390 52.110 39.395 ;
        RECT 55.790 39.395 80.110 39.405 ;
        RECT 55.790 39.380 58.290 39.395 ;
        RECT 68.720 39.390 80.110 39.395 ;
        RECT 84.850 39.395 108.110 39.405 ;
        RECT 84.850 39.380 85.790 39.395 ;
        RECT 96.720 39.390 108.110 39.395 ;
        RECT 111.790 39.395 136.110 39.405 ;
        RECT 111.790 39.380 114.290 39.395 ;
        RECT 124.720 39.390 136.110 39.395 ;
      LAYER pwell ;
        RECT 26.135 39.020 28.245 39.025 ;
        RECT 54.135 39.020 56.245 39.025 ;
        RECT 82.135 39.020 84.245 39.025 ;
        RECT 110.135 39.020 112.245 39.025 ;
        RECT 138.135 39.020 140.245 39.025 ;
        RECT 24.110 39.015 28.245 39.020 ;
        RECT 52.110 39.015 56.245 39.020 ;
        RECT 80.110 39.015 84.245 39.020 ;
        RECT 108.110 39.015 112.245 39.020 ;
        RECT 136.110 39.015 140.245 39.020 ;
        RECT 1.950 35.920 28.245 39.015 ;
        RECT 1.950 34.915 24.200 35.920 ;
        RECT 26.135 34.925 28.245 35.920 ;
        RECT 29.950 35.920 56.245 39.015 ;
        RECT 29.950 34.915 52.200 35.920 ;
        RECT 54.135 34.925 56.245 35.920 ;
        RECT 57.950 35.920 84.245 39.015 ;
        RECT 57.950 34.915 80.200 35.920 ;
        RECT 82.135 34.925 84.245 35.920 ;
        RECT 85.950 35.920 112.245 39.015 ;
        RECT 85.950 34.915 108.200 35.920 ;
        RECT 110.135 34.925 112.245 35.920 ;
        RECT 113.950 35.920 140.245 39.015 ;
        RECT 113.950 34.915 136.200 35.920 ;
        RECT 138.135 34.925 140.245 35.920 ;
      LAYER nwell ;
        RECT 27.290 33.600 29.790 33.880 ;
        RECT 55.290 33.600 57.790 33.880 ;
        RECT 83.790 33.600 86.290 33.880 ;
        RECT 111.790 33.600 114.290 33.880 ;
        RECT 5.410 33.355 12.800 33.585 ;
        RECT 1.290 31.890 12.800 33.355 ;
        RECT 26.050 33.355 29.790 33.600 ;
        RECT 33.410 33.355 40.800 33.585 ;
        RECT 26.050 31.890 40.800 33.355 ;
        RECT 54.050 33.355 57.790 33.600 ;
        RECT 61.410 33.355 68.800 33.585 ;
        RECT 54.050 31.890 68.800 33.355 ;
        RECT 82.050 33.355 86.290 33.600 ;
        RECT 89.410 33.355 96.800 33.585 ;
        RECT 82.050 31.890 96.800 33.355 ;
        RECT 110.050 33.355 114.290 33.600 ;
        RECT 117.410 33.355 124.800 33.585 ;
        RECT 110.050 31.890 124.800 33.355 ;
        RECT 1.290 29.580 21.135 31.890 ;
        RECT 26.050 29.595 49.135 31.890 ;
        RECT 54.050 29.595 77.135 31.890 ;
        RECT 82.050 29.595 105.135 31.890 ;
        RECT 110.050 29.595 133.135 31.890 ;
        RECT 138.050 29.595 140.160 33.600 ;
        RECT 24.025 29.580 49.135 29.595 ;
        RECT 52.025 29.580 77.135 29.595 ;
        RECT 80.025 29.580 105.135 29.595 ;
        RECT 108.025 29.580 133.135 29.595 ;
        RECT 136.025 29.580 140.160 29.595 ;
        RECT 1.290 23.410 140.160 29.580 ;
        RECT 1.290 23.405 26.135 23.410 ;
        RECT 28.755 23.405 54.135 23.410 ;
        RECT 56.840 23.405 82.135 23.410 ;
        RECT 83.790 23.405 110.135 23.410 ;
        RECT 111.790 23.405 138.135 23.410 ;
        RECT 1.290 23.395 24.110 23.405 ;
        RECT 12.720 23.390 24.110 23.395 ;
        RECT 28.755 23.395 52.110 23.405 ;
        RECT 28.755 23.380 29.790 23.395 ;
        RECT 40.720 23.390 52.110 23.395 ;
        RECT 56.840 23.395 80.110 23.405 ;
        RECT 56.840 23.380 57.790 23.395 ;
        RECT 68.720 23.390 80.110 23.395 ;
        RECT 83.790 23.395 108.110 23.405 ;
        RECT 83.790 23.380 86.290 23.395 ;
        RECT 96.720 23.390 108.110 23.395 ;
        RECT 111.790 23.395 136.110 23.405 ;
        RECT 111.790 23.380 114.290 23.395 ;
        RECT 124.720 23.390 136.110 23.395 ;
      LAYER pwell ;
        RECT 26.135 23.020 28.245 23.025 ;
        RECT 54.135 23.020 56.245 23.025 ;
        RECT 82.135 23.020 84.245 23.025 ;
        RECT 110.135 23.020 112.245 23.025 ;
        RECT 138.135 23.020 140.245 23.025 ;
        RECT 24.110 23.015 28.245 23.020 ;
        RECT 52.110 23.015 56.245 23.020 ;
        RECT 80.110 23.015 84.245 23.020 ;
        RECT 108.110 23.015 112.245 23.020 ;
        RECT 136.110 23.015 140.245 23.020 ;
        RECT 1.950 19.920 28.245 23.015 ;
        RECT 1.950 18.915 24.200 19.920 ;
        RECT 26.135 18.925 28.245 19.920 ;
        RECT 29.950 19.920 56.245 23.015 ;
        RECT 29.950 18.915 52.200 19.920 ;
        RECT 54.135 18.925 56.245 19.920 ;
        RECT 57.950 19.920 84.245 23.015 ;
        RECT 57.950 18.915 80.200 19.920 ;
        RECT 82.135 18.925 84.245 19.920 ;
        RECT 85.950 19.920 112.245 23.015 ;
        RECT 85.950 18.915 108.200 19.920 ;
        RECT 110.135 18.925 112.245 19.920 ;
        RECT 113.950 19.920 140.245 23.015 ;
        RECT 113.950 18.915 136.200 19.920 ;
        RECT 138.135 18.925 140.245 19.920 ;
      LAYER nwell ;
        RECT 27.790 17.600 30.290 17.880 ;
        RECT 55.290 17.600 57.790 17.880 ;
        RECT 83.790 17.600 86.290 17.880 ;
        RECT 111.790 17.600 114.290 17.880 ;
        RECT 5.410 17.355 12.800 17.585 ;
        RECT 1.290 15.890 12.800 17.355 ;
        RECT 26.050 17.355 30.290 17.600 ;
        RECT 33.410 17.355 40.800 17.585 ;
        RECT 26.050 15.890 40.800 17.355 ;
        RECT 54.050 17.355 57.790 17.600 ;
        RECT 61.410 17.355 68.800 17.585 ;
        RECT 54.050 15.890 68.800 17.355 ;
        RECT 82.050 17.355 86.290 17.600 ;
        RECT 89.410 17.355 96.800 17.585 ;
        RECT 82.050 15.890 96.800 17.355 ;
        RECT 110.050 17.355 114.290 17.600 ;
        RECT 117.410 17.355 124.800 17.585 ;
        RECT 110.050 15.890 124.800 17.355 ;
        RECT 1.290 13.580 21.135 15.890 ;
        RECT 26.050 13.595 49.135 15.890 ;
        RECT 54.050 13.595 77.135 15.890 ;
        RECT 82.050 13.595 105.135 15.890 ;
        RECT 110.050 13.595 133.135 15.890 ;
        RECT 138.050 13.595 140.160 17.600 ;
        RECT 24.025 13.580 49.135 13.595 ;
        RECT 52.025 13.580 77.135 13.595 ;
        RECT 80.025 13.580 105.135 13.595 ;
        RECT 108.025 13.580 133.135 13.595 ;
        RECT 136.025 13.580 140.160 13.595 ;
        RECT 1.290 7.410 140.160 13.580 ;
        RECT 1.290 7.405 26.135 7.410 ;
        RECT 27.790 7.405 54.135 7.410 ;
        RECT 55.495 7.405 82.135 7.410 ;
        RECT 83.790 7.405 110.135 7.410 ;
        RECT 111.790 7.405 138.135 7.410 ;
        RECT 1.290 7.395 24.110 7.405 ;
        RECT 12.720 7.390 24.110 7.395 ;
        RECT 27.790 7.395 52.110 7.405 ;
        RECT 57.115 7.400 80.110 7.405 ;
        RECT 57.290 7.395 80.110 7.400 ;
        RECT 27.790 7.380 30.290 7.395 ;
        RECT 40.720 7.390 52.110 7.395 ;
        RECT 68.720 7.390 80.110 7.395 ;
        RECT 83.790 7.395 108.110 7.405 ;
        RECT 83.790 7.380 86.290 7.395 ;
        RECT 96.720 7.390 108.110 7.395 ;
        RECT 111.790 7.395 136.110 7.405 ;
        RECT 111.790 7.380 114.290 7.395 ;
        RECT 124.720 7.390 136.110 7.395 ;
      LAYER pwell ;
        RECT 26.135 7.020 28.245 7.025 ;
        RECT 54.135 7.020 56.245 7.025 ;
        RECT 82.135 7.020 84.245 7.025 ;
        RECT 110.135 7.020 112.245 7.025 ;
        RECT 138.135 7.020 140.245 7.025 ;
        RECT 24.110 7.015 28.245 7.020 ;
        RECT 52.110 7.015 56.245 7.020 ;
        RECT 80.110 7.015 84.245 7.020 ;
        RECT 108.110 7.015 112.245 7.020 ;
        RECT 136.110 7.015 140.245 7.020 ;
        RECT 1.950 3.920 28.245 7.015 ;
        RECT 1.950 2.915 24.200 3.920 ;
        RECT 26.135 2.925 28.245 3.920 ;
        RECT 29.950 3.920 56.245 7.015 ;
        RECT 29.950 2.915 52.200 3.920 ;
        RECT 54.135 2.925 56.245 3.920 ;
        RECT 57.950 3.920 84.245 7.015 ;
        RECT 57.950 2.915 80.200 3.920 ;
        RECT 82.135 2.925 84.245 3.920 ;
        RECT 85.950 3.920 112.245 7.015 ;
        RECT 85.950 2.915 108.200 3.920 ;
        RECT 110.135 2.925 112.245 3.920 ;
        RECT 113.950 3.920 140.245 7.015 ;
        RECT 113.950 2.915 136.200 3.920 ;
        RECT 138.135 2.925 140.245 3.920 ;
      LAYER li1 ;
        RECT 14.260 212.695 126.960 212.865 ;
        RECT 14.345 211.945 15.555 212.695 ;
        RECT 15.725 211.955 16.165 212.515 ;
        RECT 16.335 211.955 16.785 212.695 ;
        RECT 16.955 212.125 17.125 212.525 ;
        RECT 17.295 212.295 17.715 212.695 ;
        RECT 17.885 212.125 18.115 212.525 ;
        RECT 16.955 211.955 18.115 212.125 ;
        RECT 18.285 211.955 18.775 212.525 ;
        RECT 14.345 211.405 14.865 211.945 ;
        RECT 15.035 211.235 15.555 211.775 ;
        RECT 14.345 210.145 15.555 211.235 ;
        RECT 15.725 210.945 16.035 211.955 ;
        RECT 16.205 211.335 16.375 211.785 ;
        RECT 16.545 211.505 16.935 211.785 ;
        RECT 17.120 211.455 17.365 211.785 ;
        RECT 16.205 211.165 16.995 211.335 ;
        RECT 15.725 210.315 16.165 210.945 ;
        RECT 16.340 210.145 16.655 210.995 ;
        RECT 16.825 210.485 16.995 211.165 ;
        RECT 17.165 210.655 17.365 211.455 ;
        RECT 17.565 210.655 17.815 211.785 ;
        RECT 18.030 211.455 18.435 211.785 ;
        RECT 18.605 211.285 18.775 211.955 ;
        RECT 18.005 211.115 18.775 211.285 ;
        RECT 18.945 211.955 19.205 212.525 ;
        RECT 19.375 212.295 19.760 212.695 ;
        RECT 19.930 212.125 20.185 212.525 ;
        RECT 19.375 211.955 20.185 212.125 ;
        RECT 20.375 211.955 20.620 212.525 ;
        RECT 20.790 212.295 21.175 212.695 ;
        RECT 21.345 212.125 21.600 212.525 ;
        RECT 20.790 211.955 21.600 212.125 ;
        RECT 21.790 211.955 22.215 212.525 ;
        RECT 22.385 212.295 22.770 212.695 ;
        RECT 22.940 212.125 23.375 212.525 ;
        RECT 22.385 211.955 23.375 212.125 ;
        RECT 23.545 211.970 23.835 212.695 ;
        RECT 24.005 212.185 24.310 212.695 ;
        RECT 18.945 211.285 19.130 211.955 ;
        RECT 19.375 211.785 19.725 211.955 ;
        RECT 20.375 211.785 20.545 211.955 ;
        RECT 20.790 211.785 21.140 211.955 ;
        RECT 21.790 211.785 22.140 211.955 ;
        RECT 22.385 211.785 22.720 211.955 ;
        RECT 19.300 211.455 19.725 211.785 ;
        RECT 18.005 210.485 18.255 211.115 ;
        RECT 16.825 210.315 18.255 210.485 ;
        RECT 18.435 210.145 18.765 210.945 ;
        RECT 18.945 210.315 19.205 211.285 ;
        RECT 19.375 210.935 19.725 211.455 ;
        RECT 19.895 211.285 20.545 211.785 ;
        RECT 20.715 211.455 21.140 211.785 ;
        RECT 19.895 211.105 20.620 211.285 ;
        RECT 19.375 210.740 20.185 210.935 ;
        RECT 19.375 210.145 19.760 210.570 ;
        RECT 19.930 210.315 20.185 210.740 ;
        RECT 20.375 210.315 20.620 211.105 ;
        RECT 20.790 210.935 21.140 211.455 ;
        RECT 21.310 211.285 22.140 211.785 ;
        RECT 22.310 211.455 22.720 211.785 ;
        RECT 21.310 211.105 22.215 211.285 ;
        RECT 20.790 210.740 21.620 210.935 ;
        RECT 20.790 210.145 21.175 210.570 ;
        RECT 21.345 210.315 21.620 210.740 ;
        RECT 21.790 210.315 22.215 211.105 ;
        RECT 22.385 210.910 22.720 211.455 ;
        RECT 22.890 211.080 23.375 211.785 ;
        RECT 24.005 211.455 24.320 212.015 ;
        RECT 24.490 211.705 24.740 212.515 ;
        RECT 24.910 212.170 25.170 212.695 ;
        RECT 25.350 211.705 25.600 212.515 ;
        RECT 25.770 212.135 26.030 212.695 ;
        RECT 26.200 212.045 26.460 212.500 ;
        RECT 26.630 212.215 26.890 212.695 ;
        RECT 27.060 212.045 27.320 212.500 ;
        RECT 27.490 212.215 27.750 212.695 ;
        RECT 27.920 212.045 28.180 212.500 ;
        RECT 28.350 212.215 28.595 212.695 ;
        RECT 28.765 212.045 29.040 212.500 ;
        RECT 29.210 212.215 29.455 212.695 ;
        RECT 29.625 212.045 29.885 212.500 ;
        RECT 30.065 212.215 30.315 212.695 ;
        RECT 30.485 212.045 30.745 212.500 ;
        RECT 30.925 212.215 31.175 212.695 ;
        RECT 31.345 212.045 31.605 212.500 ;
        RECT 31.785 212.215 32.045 212.695 ;
        RECT 32.215 212.045 32.475 212.500 ;
        RECT 32.645 212.215 32.945 212.695 ;
        RECT 33.385 212.315 33.715 212.695 ;
        RECT 33.885 212.145 34.075 212.525 ;
        RECT 34.245 212.335 34.575 212.695 ;
        RECT 26.200 211.875 32.945 212.045 ;
        RECT 24.490 211.455 31.610 211.705 ;
        RECT 22.385 210.740 23.375 210.910 ;
        RECT 22.385 210.145 22.770 210.570 ;
        RECT 22.940 210.315 23.375 210.740 ;
        RECT 23.545 210.145 23.835 211.310 ;
        RECT 24.015 210.145 24.310 210.955 ;
        RECT 24.490 210.315 24.735 211.455 ;
        RECT 24.910 210.145 25.170 210.955 ;
        RECT 25.350 210.320 25.600 211.455 ;
        RECT 31.780 211.335 32.945 211.875 ;
        RECT 33.675 211.955 34.075 212.145 ;
        RECT 34.795 212.125 34.985 212.525 ;
        RECT 34.245 211.955 34.985 212.125 ;
        RECT 31.780 211.285 32.975 211.335 ;
        RECT 26.200 211.165 32.975 211.285 ;
        RECT 26.200 211.060 32.945 211.165 ;
        RECT 26.200 211.045 31.605 211.060 ;
        RECT 25.770 210.150 26.030 210.945 ;
        RECT 26.200 210.320 26.460 211.045 ;
        RECT 26.630 210.150 26.890 210.875 ;
        RECT 27.060 210.320 27.320 211.045 ;
        RECT 27.490 210.150 27.750 210.875 ;
        RECT 27.920 210.320 28.180 211.045 ;
        RECT 28.350 210.150 28.610 210.875 ;
        RECT 28.780 210.320 29.040 211.045 ;
        RECT 29.210 210.150 29.455 210.875 ;
        RECT 29.625 210.320 29.885 211.045 ;
        RECT 30.070 210.150 30.315 210.875 ;
        RECT 30.485 210.320 30.745 211.045 ;
        RECT 30.930 210.150 31.175 210.875 ;
        RECT 31.345 210.320 31.605 211.045 ;
        RECT 31.790 210.150 32.045 210.875 ;
        RECT 32.215 210.320 32.505 211.060 ;
        RECT 25.770 210.145 32.045 210.150 ;
        RECT 32.675 210.145 32.945 210.890 ;
        RECT 33.215 210.145 33.505 211.115 ;
        RECT 33.675 210.315 33.905 211.955 ;
        RECT 34.245 211.785 34.415 211.955 ;
        RECT 34.075 211.090 34.415 211.785 ;
        RECT 34.585 211.370 34.910 211.785 ;
        RECT 35.360 211.455 35.740 212.415 ;
        RECT 35.925 212.215 36.255 212.695 ;
        RECT 35.930 211.455 36.245 212.030 ;
        RECT 36.425 211.970 36.715 212.695 ;
        RECT 36.910 211.940 37.145 212.270 ;
        RECT 37.315 211.955 37.645 212.695 ;
        RECT 37.880 212.315 39.075 212.525 ;
        RECT 34.075 210.860 34.910 211.090 ;
        RECT 34.075 210.145 34.405 210.560 ;
        RECT 34.595 210.315 34.910 210.860 ;
        RECT 35.080 210.845 36.195 211.110 ;
        RECT 35.080 210.315 35.305 210.845 ;
        RECT 35.475 210.145 35.805 210.655 ;
        RECT 35.975 210.315 36.195 210.845 ;
        RECT 36.425 210.145 36.715 211.310 ;
        RECT 36.910 211.285 37.080 211.940 ;
        RECT 37.880 211.875 38.155 212.315 ;
        RECT 38.325 211.975 38.655 212.145 ;
        RECT 38.330 211.875 38.655 211.975 ;
        RECT 38.825 212.085 39.075 212.315 ;
        RECT 39.245 212.255 39.415 212.695 ;
        RECT 39.585 212.085 39.935 212.525 ;
        RECT 40.105 212.185 40.410 212.695 ;
        RECT 38.825 211.875 39.935 212.085 ;
        RECT 37.255 211.455 37.600 211.785 ;
        RECT 37.830 211.285 38.160 211.705 ;
        RECT 36.910 211.115 38.160 211.285 ;
        RECT 36.910 210.920 37.210 211.115 ;
        RECT 38.330 210.945 38.610 211.875 ;
        RECT 38.790 211.505 39.935 211.705 ;
        RECT 38.790 211.125 38.980 211.505 ;
        RECT 40.105 211.455 40.420 212.015 ;
        RECT 40.590 211.705 40.840 212.515 ;
        RECT 41.010 212.170 41.270 212.695 ;
        RECT 41.450 211.705 41.700 212.515 ;
        RECT 41.870 212.135 42.130 212.695 ;
        RECT 42.300 212.045 42.560 212.500 ;
        RECT 42.730 212.215 42.990 212.695 ;
        RECT 43.160 212.045 43.420 212.500 ;
        RECT 43.590 212.215 43.850 212.695 ;
        RECT 44.020 212.045 44.280 212.500 ;
        RECT 44.450 212.215 44.695 212.695 ;
        RECT 44.865 212.045 45.140 212.500 ;
        RECT 45.310 212.215 45.555 212.695 ;
        RECT 45.725 212.045 45.985 212.500 ;
        RECT 46.165 212.215 46.415 212.695 ;
        RECT 46.585 212.045 46.845 212.500 ;
        RECT 47.025 212.215 47.275 212.695 ;
        RECT 47.445 212.045 47.705 212.500 ;
        RECT 47.885 212.215 48.145 212.695 ;
        RECT 48.315 212.045 48.575 212.500 ;
        RECT 48.745 212.215 49.045 212.695 ;
        RECT 42.300 212.015 49.045 212.045 ;
        RECT 42.300 211.875 49.075 212.015 ;
        RECT 49.305 211.970 49.595 212.695 ;
        RECT 49.765 212.185 50.070 212.695 ;
        RECT 47.880 211.845 49.075 211.875 ;
        RECT 40.590 211.455 47.710 211.705 ;
        RECT 39.160 210.945 39.435 211.285 ;
        RECT 37.380 210.145 37.635 210.945 ;
        RECT 37.835 210.775 39.435 210.945 ;
        RECT 37.835 210.315 38.165 210.775 ;
        RECT 38.335 210.145 38.910 210.605 ;
        RECT 39.080 210.315 39.435 210.775 ;
        RECT 39.605 210.145 39.935 211.285 ;
        RECT 40.115 210.145 40.410 210.955 ;
        RECT 40.590 210.315 40.835 211.455 ;
        RECT 41.010 210.145 41.270 210.955 ;
        RECT 41.450 210.320 41.700 211.455 ;
        RECT 47.880 211.285 49.045 211.845 ;
        RECT 49.765 211.455 50.080 212.015 ;
        RECT 50.250 211.705 50.500 212.515 ;
        RECT 50.670 212.170 50.930 212.695 ;
        RECT 51.110 211.705 51.360 212.515 ;
        RECT 51.530 212.135 51.790 212.695 ;
        RECT 51.960 212.045 52.220 212.500 ;
        RECT 52.390 212.215 52.650 212.695 ;
        RECT 52.820 212.045 53.080 212.500 ;
        RECT 53.250 212.215 53.510 212.695 ;
        RECT 53.680 212.045 53.940 212.500 ;
        RECT 54.110 212.215 54.355 212.695 ;
        RECT 54.525 212.045 54.800 212.500 ;
        RECT 54.970 212.215 55.215 212.695 ;
        RECT 55.385 212.045 55.645 212.500 ;
        RECT 55.825 212.215 56.075 212.695 ;
        RECT 56.245 212.045 56.505 212.500 ;
        RECT 56.685 212.215 56.935 212.695 ;
        RECT 57.105 212.045 57.365 212.500 ;
        RECT 57.545 212.215 57.805 212.695 ;
        RECT 57.975 212.045 58.235 212.500 ;
        RECT 58.405 212.215 58.705 212.695 ;
        RECT 51.960 211.875 58.705 212.045 ;
        RECT 50.250 211.455 57.370 211.705 ;
        RECT 42.300 211.060 49.045 211.285 ;
        RECT 42.300 211.045 47.705 211.060 ;
        RECT 41.870 210.150 42.130 210.945 ;
        RECT 42.300 210.320 42.560 211.045 ;
        RECT 42.730 210.150 42.990 210.875 ;
        RECT 43.160 210.320 43.420 211.045 ;
        RECT 43.590 210.150 43.850 210.875 ;
        RECT 44.020 210.320 44.280 211.045 ;
        RECT 44.450 210.150 44.710 210.875 ;
        RECT 44.880 210.320 45.140 211.045 ;
        RECT 45.310 210.150 45.555 210.875 ;
        RECT 45.725 210.320 45.985 211.045 ;
        RECT 46.170 210.150 46.415 210.875 ;
        RECT 46.585 210.320 46.845 211.045 ;
        RECT 47.030 210.150 47.275 210.875 ;
        RECT 47.445 210.320 47.705 211.045 ;
        RECT 47.890 210.150 48.145 210.875 ;
        RECT 48.315 210.320 48.605 211.060 ;
        RECT 41.870 210.145 48.145 210.150 ;
        RECT 48.775 210.145 49.045 210.890 ;
        RECT 49.305 210.145 49.595 211.310 ;
        RECT 49.775 210.145 50.070 210.955 ;
        RECT 50.250 210.315 50.495 211.455 ;
        RECT 50.670 210.145 50.930 210.955 ;
        RECT 51.110 210.320 51.360 211.455 ;
        RECT 57.540 211.285 58.705 211.875 ;
        RECT 51.960 211.060 58.705 211.285 ;
        RECT 58.990 211.940 59.225 212.270 ;
        RECT 59.395 211.955 59.725 212.695 ;
        RECT 59.960 212.315 61.155 212.525 ;
        RECT 58.990 211.285 59.160 211.940 ;
        RECT 59.960 211.875 60.235 212.315 ;
        RECT 60.405 211.875 60.735 212.145 ;
        RECT 60.905 212.085 61.155 212.315 ;
        RECT 61.325 212.255 61.495 212.695 ;
        RECT 61.665 212.085 62.015 212.525 ;
        RECT 60.905 211.875 62.015 212.085 ;
        RECT 62.185 211.970 62.475 212.695 ;
        RECT 62.645 212.195 62.945 212.525 ;
        RECT 63.115 212.215 63.390 212.695 ;
        RECT 60.405 211.845 60.690 211.875 ;
        RECT 59.335 211.455 59.680 211.785 ;
        RECT 59.910 211.285 60.240 211.705 ;
        RECT 58.990 211.115 60.240 211.285 ;
        RECT 51.960 211.045 57.365 211.060 ;
        RECT 51.530 210.150 51.790 210.945 ;
        RECT 51.960 210.320 52.220 211.045 ;
        RECT 52.390 210.150 52.650 210.875 ;
        RECT 52.820 210.320 53.080 211.045 ;
        RECT 53.250 210.150 53.510 210.875 ;
        RECT 53.680 210.320 53.940 211.045 ;
        RECT 54.110 210.150 54.370 210.875 ;
        RECT 54.540 210.320 54.800 211.045 ;
        RECT 54.970 210.150 55.215 210.875 ;
        RECT 55.385 210.320 55.645 211.045 ;
        RECT 55.830 210.150 56.075 210.875 ;
        RECT 56.245 210.320 56.505 211.045 ;
        RECT 56.690 210.150 56.935 210.875 ;
        RECT 57.105 210.320 57.365 211.045 ;
        RECT 57.550 210.150 57.805 210.875 ;
        RECT 57.975 210.320 58.265 211.060 ;
        RECT 58.990 210.920 59.290 211.115 ;
        RECT 60.410 210.945 60.690 211.845 ;
        RECT 60.870 211.505 62.015 211.705 ;
        RECT 60.870 211.125 61.060 211.505 ;
        RECT 61.240 210.945 61.515 211.285 ;
        RECT 51.530 210.145 57.805 210.150 ;
        RECT 58.435 210.145 58.705 210.890 ;
        RECT 59.460 210.145 59.715 210.945 ;
        RECT 59.915 210.775 61.515 210.945 ;
        RECT 59.915 210.315 60.245 210.775 ;
        RECT 60.415 210.145 60.990 210.605 ;
        RECT 61.160 210.315 61.515 210.775 ;
        RECT 61.685 210.145 62.015 211.285 ;
        RECT 62.185 210.145 62.475 211.310 ;
        RECT 62.645 211.285 62.815 212.195 ;
        RECT 63.570 212.045 63.865 212.435 ;
        RECT 64.035 212.215 64.290 212.695 ;
        RECT 64.465 212.045 64.725 212.435 ;
        RECT 64.895 212.215 65.175 212.695 ;
        RECT 62.985 211.455 63.335 212.025 ;
        RECT 63.570 211.875 65.220 212.045 ;
        RECT 65.410 211.875 65.685 212.695 ;
        RECT 65.855 212.055 66.185 212.525 ;
        RECT 66.355 212.225 66.525 212.695 ;
        RECT 66.695 212.055 67.025 212.525 ;
        RECT 67.195 212.225 67.485 212.695 ;
        RECT 65.855 212.045 67.025 212.055 ;
        RECT 67.795 212.145 67.965 212.525 ;
        RECT 68.180 212.315 68.510 212.695 ;
        RECT 65.855 211.875 67.455 212.045 ;
        RECT 67.795 211.975 68.510 212.145 ;
        RECT 63.505 211.535 64.645 211.705 ;
        RECT 63.505 211.285 63.675 211.535 ;
        RECT 64.815 211.365 65.220 211.875 ;
        RECT 65.410 211.505 66.130 211.705 ;
        RECT 66.300 211.505 67.070 211.705 ;
        RECT 62.645 211.115 63.675 211.285 ;
        RECT 64.465 211.195 65.220 211.365 ;
        RECT 67.240 211.335 67.455 211.875 ;
        RECT 67.705 211.425 68.060 211.795 ;
        RECT 68.340 211.785 68.510 211.975 ;
        RECT 68.680 211.950 68.935 212.525 ;
        RECT 68.340 211.455 68.595 211.785 ;
        RECT 62.645 210.315 62.955 211.115 ;
        RECT 64.465 210.945 64.725 211.195 ;
        RECT 65.410 211.115 66.525 211.325 ;
        RECT 63.125 210.145 63.435 210.945 ;
        RECT 63.605 210.775 64.725 210.945 ;
        RECT 63.605 210.315 63.865 210.775 ;
        RECT 64.035 210.145 64.290 210.605 ;
        RECT 64.465 210.315 64.725 210.775 ;
        RECT 64.895 210.145 65.180 211.015 ;
        RECT 65.410 210.315 65.685 211.115 ;
        RECT 65.855 210.145 66.185 210.945 ;
        RECT 66.355 210.485 66.525 211.115 ;
        RECT 66.695 211.115 67.455 211.335 ;
        RECT 68.340 211.245 68.510 211.455 ;
        RECT 66.695 210.655 67.025 211.115 ;
        RECT 67.795 211.075 68.510 211.245 ;
        RECT 68.765 211.220 68.935 211.950 ;
        RECT 69.110 211.855 69.370 212.695 ;
        RECT 70.025 211.885 70.265 212.695 ;
        RECT 70.435 211.885 70.765 212.525 ;
        RECT 70.935 211.885 71.205 212.695 ;
        RECT 71.385 212.020 71.645 212.525 ;
        RECT 71.825 212.315 72.155 212.695 ;
        RECT 72.335 212.145 72.505 212.525 ;
        RECT 70.005 211.455 70.355 211.705 ;
        RECT 67.195 210.485 67.495 210.945 ;
        RECT 66.355 210.315 67.495 210.485 ;
        RECT 67.795 210.315 67.965 211.075 ;
        RECT 68.180 210.145 68.510 210.905 ;
        RECT 68.680 210.315 68.935 211.220 ;
        RECT 69.110 210.145 69.370 211.295 ;
        RECT 70.525 211.285 70.695 211.885 ;
        RECT 70.865 211.455 71.215 211.705 ;
        RECT 70.015 211.115 70.695 211.285 ;
        RECT 70.015 210.330 70.345 211.115 ;
        RECT 70.875 210.145 71.205 211.285 ;
        RECT 71.385 211.220 71.565 212.020 ;
        RECT 71.840 211.975 72.505 212.145 ;
        RECT 72.765 212.020 73.025 212.525 ;
        RECT 73.205 212.315 73.535 212.695 ;
        RECT 73.715 212.145 73.885 212.525 ;
        RECT 71.840 211.720 72.010 211.975 ;
        RECT 71.735 211.390 72.010 211.720 ;
        RECT 72.235 211.425 72.575 211.795 ;
        RECT 71.840 211.245 72.010 211.390 ;
        RECT 71.385 210.315 71.655 211.220 ;
        RECT 71.840 211.075 72.515 211.245 ;
        RECT 71.825 210.145 72.155 210.905 ;
        RECT 72.335 210.315 72.515 211.075 ;
        RECT 72.765 211.220 72.945 212.020 ;
        RECT 73.220 211.975 73.885 212.145 ;
        RECT 73.220 211.720 73.390 211.975 ;
        RECT 75.065 211.970 75.355 212.695 ;
        RECT 75.525 212.020 75.785 212.525 ;
        RECT 75.965 212.315 76.295 212.695 ;
        RECT 76.475 212.145 76.645 212.525 ;
        RECT 73.115 211.390 73.390 211.720 ;
        RECT 73.615 211.425 73.955 211.795 ;
        RECT 73.220 211.245 73.390 211.390 ;
        RECT 72.765 210.315 73.035 211.220 ;
        RECT 73.220 211.075 73.895 211.245 ;
        RECT 73.205 210.145 73.535 210.905 ;
        RECT 73.715 210.315 73.895 211.075 ;
        RECT 75.065 210.145 75.355 211.310 ;
        RECT 75.525 211.220 75.705 212.020 ;
        RECT 75.980 211.975 76.645 212.145 ;
        RECT 76.905 212.020 77.165 212.525 ;
        RECT 77.345 212.315 77.675 212.695 ;
        RECT 77.855 212.145 78.025 212.525 ;
        RECT 75.980 211.720 76.150 211.975 ;
        RECT 75.875 211.390 76.150 211.720 ;
        RECT 76.375 211.425 76.715 211.795 ;
        RECT 75.980 211.245 76.150 211.390 ;
        RECT 75.525 210.315 75.795 211.220 ;
        RECT 75.980 211.075 76.655 211.245 ;
        RECT 75.965 210.145 76.295 210.905 ;
        RECT 76.475 210.315 76.655 211.075 ;
        RECT 76.905 211.220 77.085 212.020 ;
        RECT 77.360 211.975 78.025 212.145 ;
        RECT 78.375 212.045 78.545 212.525 ;
        RECT 78.725 212.215 78.965 212.695 ;
        RECT 79.215 212.045 79.385 212.525 ;
        RECT 79.555 212.215 79.885 212.695 ;
        RECT 80.055 212.045 80.225 212.525 ;
        RECT 77.360 211.720 77.530 211.975 ;
        RECT 78.375 211.875 79.010 212.045 ;
        RECT 79.215 211.875 80.225 212.045 ;
        RECT 80.395 211.895 80.725 212.695 ;
        RECT 81.045 212.020 81.305 212.525 ;
        RECT 81.485 212.315 81.815 212.695 ;
        RECT 81.995 212.145 82.165 212.525 ;
        RECT 77.255 211.390 77.530 211.720 ;
        RECT 77.755 211.425 78.095 211.795 ;
        RECT 78.840 211.705 79.010 211.875 ;
        RECT 79.725 211.845 80.225 211.875 ;
        RECT 78.290 211.465 78.670 211.705 ;
        RECT 78.840 211.535 79.340 211.705 ;
        RECT 77.360 211.245 77.530 211.390 ;
        RECT 78.840 211.295 79.010 211.535 ;
        RECT 79.730 211.335 80.225 211.845 ;
        RECT 76.905 210.315 77.175 211.220 ;
        RECT 77.360 211.075 78.035 211.245 ;
        RECT 77.345 210.145 77.675 210.905 ;
        RECT 77.855 210.315 78.035 211.075 ;
        RECT 78.295 211.125 79.010 211.295 ;
        RECT 79.215 211.165 80.225 211.335 ;
        RECT 78.295 210.315 78.625 211.125 ;
        RECT 78.795 210.145 79.035 210.945 ;
        RECT 79.215 210.315 79.385 211.165 ;
        RECT 79.555 210.145 79.885 210.945 ;
        RECT 80.055 210.315 80.225 211.165 ;
        RECT 80.395 210.145 80.725 211.295 ;
        RECT 81.045 211.220 81.225 212.020 ;
        RECT 81.500 211.975 82.165 212.145 ;
        RECT 81.500 211.720 81.670 211.975 ;
        RECT 81.395 211.390 81.670 211.720 ;
        RECT 81.895 211.425 82.235 211.795 ;
        RECT 81.500 211.245 81.670 211.390 ;
        RECT 81.045 210.315 81.315 211.220 ;
        RECT 81.500 211.075 82.175 211.245 ;
        RECT 81.485 210.145 81.815 210.905 ;
        RECT 81.995 210.315 82.175 211.075 ;
        RECT 82.425 211.040 82.945 212.525 ;
        RECT 83.115 212.035 83.455 212.695 ;
        RECT 83.805 212.020 84.065 212.525 ;
        RECT 84.245 212.315 84.575 212.695 ;
        RECT 84.755 212.145 84.925 212.525 ;
        RECT 82.615 210.145 82.945 210.870 ;
        RECT 83.115 210.315 83.635 211.865 ;
        RECT 83.805 211.220 83.985 212.020 ;
        RECT 84.260 211.975 84.925 212.145 ;
        RECT 84.260 211.720 84.430 211.975 ;
        RECT 85.190 211.855 85.450 212.695 ;
        RECT 85.625 211.950 85.880 212.525 ;
        RECT 86.050 212.315 86.380 212.695 ;
        RECT 86.595 212.145 86.765 212.525 ;
        RECT 86.050 211.975 86.765 212.145 ;
        RECT 84.155 211.390 84.430 211.720 ;
        RECT 84.655 211.425 84.995 211.795 ;
        RECT 84.260 211.245 84.430 211.390 ;
        RECT 83.805 210.315 84.075 211.220 ;
        RECT 84.260 211.075 84.935 211.245 ;
        RECT 84.245 210.145 84.575 210.905 ;
        RECT 84.755 210.315 84.935 211.075 ;
        RECT 85.190 210.145 85.450 211.295 ;
        RECT 85.625 211.220 85.795 211.950 ;
        RECT 86.050 211.785 86.220 211.975 ;
        RECT 87.945 211.970 88.235 212.695 ;
        RECT 88.405 212.020 88.665 212.525 ;
        RECT 88.845 212.315 89.175 212.695 ;
        RECT 89.355 212.145 89.525 212.525 ;
        RECT 85.965 211.455 86.220 211.785 ;
        RECT 86.050 211.245 86.220 211.455 ;
        RECT 86.500 211.425 86.855 211.795 ;
        RECT 85.625 210.315 85.880 211.220 ;
        RECT 86.050 211.075 86.765 211.245 ;
        RECT 86.050 210.145 86.380 210.905 ;
        RECT 86.595 210.315 86.765 211.075 ;
        RECT 87.945 210.145 88.235 211.310 ;
        RECT 88.405 211.220 88.585 212.020 ;
        RECT 88.860 211.975 89.525 212.145 ;
        RECT 88.860 211.720 89.030 211.975 ;
        RECT 88.755 211.390 89.030 211.720 ;
        RECT 89.255 211.425 89.595 211.795 ;
        RECT 88.860 211.245 89.030 211.390 ;
        RECT 88.405 210.315 88.675 211.220 ;
        RECT 88.860 211.075 89.535 211.245 ;
        RECT 88.845 210.145 89.175 210.905 ;
        RECT 89.355 210.315 89.535 211.075 ;
        RECT 89.785 210.315 90.535 212.525 ;
        RECT 91.625 212.020 91.885 212.525 ;
        RECT 92.065 212.315 92.395 212.695 ;
        RECT 92.575 212.145 92.745 212.525 ;
        RECT 93.010 212.295 93.345 212.695 ;
        RECT 91.625 211.220 91.805 212.020 ;
        RECT 92.080 211.975 92.745 212.145 ;
        RECT 93.515 212.125 93.720 212.525 ;
        RECT 93.930 212.215 94.205 212.695 ;
        RECT 94.415 212.195 94.675 212.525 ;
        RECT 92.080 211.720 92.250 211.975 ;
        RECT 93.035 211.955 93.720 212.125 ;
        RECT 91.975 211.390 92.250 211.720 ;
        RECT 92.475 211.425 92.815 211.795 ;
        RECT 92.080 211.245 92.250 211.390 ;
        RECT 91.625 210.315 91.895 211.220 ;
        RECT 92.080 211.075 92.755 211.245 ;
        RECT 92.065 210.145 92.395 210.905 ;
        RECT 92.575 210.315 92.755 211.075 ;
        RECT 93.035 210.925 93.375 211.955 ;
        RECT 93.545 211.285 93.795 211.785 ;
        RECT 93.975 211.455 94.335 212.035 ;
        RECT 94.505 211.285 94.675 212.195 ;
        RECT 93.545 211.115 94.675 211.285 ;
        RECT 93.035 210.750 93.700 210.925 ;
        RECT 93.010 210.145 93.345 210.570 ;
        RECT 93.515 210.345 93.700 210.750 ;
        RECT 93.905 210.145 94.235 210.925 ;
        RECT 94.405 210.345 94.675 211.115 ;
        RECT 94.845 212.020 95.120 212.365 ;
        RECT 95.310 212.295 95.690 212.695 ;
        RECT 95.860 212.125 96.030 212.475 ;
        RECT 96.200 212.295 96.530 212.695 ;
        RECT 96.715 212.125 96.885 212.475 ;
        RECT 97.055 212.295 97.430 212.695 ;
        RECT 97.655 212.125 97.825 212.330 ;
        RECT 94.845 211.285 95.015 212.020 ;
        RECT 95.290 211.955 96.885 212.125 ;
        RECT 97.325 211.955 97.825 212.125 ;
        RECT 98.075 211.955 98.245 212.695 ;
        RECT 98.500 211.955 98.815 212.330 ;
        RECT 95.290 211.785 95.460 211.955 ;
        RECT 95.185 211.455 95.460 211.785 ;
        RECT 95.630 211.455 96.285 211.785 ;
        RECT 95.290 211.285 95.460 211.455 ;
        RECT 96.505 211.365 96.675 211.785 ;
        RECT 97.325 211.705 97.495 211.955 ;
        RECT 97.070 211.535 97.495 211.705 ;
        RECT 94.845 210.315 95.120 211.285 ;
        RECT 95.290 211.115 95.950 211.285 ;
        RECT 96.505 211.195 97.155 211.365 ;
        RECT 95.780 210.995 95.950 211.115 ;
        RECT 95.330 210.145 95.610 210.945 ;
        RECT 95.780 210.825 96.815 210.995 ;
        RECT 95.780 210.325 96.420 210.655 ;
        RECT 96.645 210.575 96.815 210.825 ;
        RECT 96.985 210.915 97.155 211.195 ;
        RECT 97.325 211.255 97.495 211.535 ;
        RECT 97.665 211.455 97.955 211.785 ;
        RECT 97.325 211.085 97.910 211.255 ;
        RECT 98.125 211.085 98.475 211.785 ;
        RECT 98.645 210.915 98.815 211.955 ;
        RECT 98.985 211.925 100.655 212.695 ;
        RECT 100.825 211.970 101.115 212.695 ;
        RECT 101.745 212.020 102.005 212.525 ;
        RECT 102.185 212.315 102.515 212.695 ;
        RECT 102.695 212.145 102.865 212.525 ;
        RECT 96.985 210.745 98.815 210.915 ;
        RECT 96.645 210.405 97.390 210.575 ;
        RECT 98.055 210.145 98.385 210.575 ;
        RECT 98.555 210.325 98.815 210.745 ;
        RECT 98.985 211.235 99.735 211.755 ;
        RECT 99.905 211.405 100.655 211.925 ;
        RECT 98.985 210.145 100.655 211.235 ;
        RECT 100.825 210.145 101.115 211.310 ;
        RECT 101.745 211.220 101.925 212.020 ;
        RECT 102.200 211.975 102.865 212.145 ;
        RECT 102.200 211.720 102.370 211.975 ;
        RECT 103.125 211.945 104.335 212.695 ;
        RECT 102.095 211.390 102.370 211.720 ;
        RECT 102.595 211.425 102.935 211.795 ;
        RECT 102.200 211.245 102.370 211.390 ;
        RECT 101.745 210.315 102.015 211.220 ;
        RECT 102.200 211.075 102.875 211.245 ;
        RECT 102.185 210.145 102.515 210.905 ;
        RECT 102.695 210.315 102.875 211.075 ;
        RECT 103.125 211.235 103.645 211.775 ;
        RECT 103.815 211.405 104.335 211.945 ;
        RECT 104.510 211.855 104.770 212.695 ;
        RECT 104.945 211.950 105.200 212.525 ;
        RECT 105.370 212.315 105.700 212.695 ;
        RECT 105.915 212.145 106.085 212.525 ;
        RECT 105.370 211.975 106.085 212.145 ;
        RECT 103.125 210.145 104.335 211.235 ;
        RECT 104.510 210.145 104.770 211.295 ;
        RECT 104.945 211.220 105.115 211.950 ;
        RECT 105.370 211.785 105.540 211.975 ;
        RECT 106.345 211.925 108.015 212.695 ;
        RECT 105.285 211.455 105.540 211.785 ;
        RECT 105.370 211.245 105.540 211.455 ;
        RECT 105.820 211.425 106.175 211.795 ;
        RECT 104.945 210.315 105.200 211.220 ;
        RECT 105.370 211.075 106.085 211.245 ;
        RECT 105.370 210.145 105.700 210.905 ;
        RECT 105.915 210.315 106.085 211.075 ;
        RECT 106.345 211.235 107.095 211.755 ;
        RECT 107.265 211.405 108.015 211.925 ;
        RECT 108.185 212.020 108.445 212.525 ;
        RECT 108.625 212.315 108.955 212.695 ;
        RECT 109.135 212.145 109.305 212.525 ;
        RECT 106.345 210.145 108.015 211.235 ;
        RECT 108.185 211.220 108.355 212.020 ;
        RECT 108.640 211.975 109.305 212.145 ;
        RECT 108.640 211.720 108.810 211.975 ;
        RECT 109.565 211.925 111.235 212.695 ;
        RECT 108.525 211.390 108.810 211.720 ;
        RECT 109.045 211.425 109.375 211.795 ;
        RECT 108.640 211.245 108.810 211.390 ;
        RECT 108.185 210.315 108.455 211.220 ;
        RECT 108.640 211.075 109.305 211.245 ;
        RECT 108.625 210.145 108.955 210.905 ;
        RECT 109.135 210.315 109.305 211.075 ;
        RECT 109.565 211.235 110.315 211.755 ;
        RECT 110.485 211.405 111.235 211.925 ;
        RECT 111.405 212.020 111.665 212.525 ;
        RECT 111.845 212.315 112.175 212.695 ;
        RECT 112.355 212.145 112.525 212.525 ;
        RECT 109.565 210.145 111.235 211.235 ;
        RECT 111.405 211.220 111.585 212.020 ;
        RECT 111.860 211.975 112.525 212.145 ;
        RECT 111.860 211.720 112.030 211.975 ;
        RECT 113.705 211.970 113.995 212.695 ;
        RECT 114.630 212.150 119.975 212.695 ;
        RECT 120.150 212.150 125.495 212.695 ;
        RECT 111.755 211.390 112.030 211.720 ;
        RECT 112.255 211.425 112.595 211.795 ;
        RECT 111.860 211.245 112.030 211.390 ;
        RECT 111.405 210.315 111.675 211.220 ;
        RECT 111.860 211.075 112.535 211.245 ;
        RECT 111.845 210.145 112.175 210.905 ;
        RECT 112.355 210.315 112.535 211.075 ;
        RECT 113.705 210.145 113.995 211.310 ;
        RECT 116.220 210.580 116.570 211.830 ;
        RECT 118.050 211.320 118.390 212.150 ;
        RECT 121.740 210.580 122.090 211.830 ;
        RECT 123.570 211.320 123.910 212.150 ;
        RECT 125.665 211.945 126.875 212.695 ;
        RECT 125.665 211.235 126.185 211.775 ;
        RECT 126.355 211.405 126.875 211.945 ;
        RECT 114.630 210.145 119.975 210.580 ;
        RECT 120.150 210.145 125.495 210.580 ;
        RECT 125.665 210.145 126.875 211.235 ;
        RECT 14.260 209.975 126.960 210.145 ;
        RECT 14.345 208.885 15.555 209.975 ;
        RECT 14.345 208.175 14.865 208.715 ;
        RECT 15.035 208.345 15.555 208.885 ;
        RECT 16.185 208.820 16.525 209.805 ;
        RECT 16.695 209.545 17.105 209.975 ;
        RECT 17.850 209.555 18.180 209.975 ;
        RECT 18.350 209.375 18.675 209.805 ;
        RECT 16.695 209.205 18.675 209.375 ;
        RECT 14.345 207.425 15.555 208.175 ;
        RECT 16.185 208.165 16.440 208.820 ;
        RECT 16.695 208.665 16.960 209.205 ;
        RECT 17.175 208.865 17.800 209.035 ;
        RECT 16.610 208.335 16.960 208.665 ;
        RECT 17.130 208.335 17.460 208.665 ;
        RECT 17.630 208.165 17.800 208.865 ;
        RECT 16.185 207.790 16.545 208.165 ;
        RECT 16.245 207.765 16.415 207.790 ;
        RECT 16.810 207.425 16.980 208.165 ;
        RECT 17.260 207.995 17.800 208.165 ;
        RECT 17.970 208.795 18.675 209.205 ;
        RECT 19.150 208.875 19.480 209.975 ;
        RECT 20.370 209.625 21.645 209.805 ;
        RECT 20.370 209.135 20.675 209.625 ;
        RECT 17.260 207.790 17.430 207.995 ;
        RECT 17.970 207.595 18.140 208.795 ;
        RECT 18.310 208.415 18.880 208.625 ;
        RECT 19.050 208.415 19.695 208.625 ;
        RECT 20.385 208.335 20.660 208.965 ;
        RECT 18.370 208.075 19.540 208.245 ;
        RECT 18.370 207.595 18.700 208.075 ;
        RECT 18.870 207.425 19.040 207.895 ;
        RECT 19.210 207.610 19.540 208.075 ;
        RECT 20.335 207.425 20.665 208.165 ;
        RECT 20.845 208.125 21.145 209.455 ;
        RECT 21.315 209.365 21.645 209.625 ;
        RECT 21.815 209.535 21.985 209.975 ;
        RECT 22.240 209.445 22.410 209.805 ;
        RECT 22.590 209.615 22.920 209.975 ;
        RECT 23.090 209.445 23.350 209.805 ;
        RECT 22.240 209.365 23.350 209.445 ;
        RECT 21.315 209.195 23.350 209.365 ;
        RECT 21.530 208.835 23.315 209.015 ;
        RECT 21.530 208.585 21.855 208.835 ;
        RECT 21.525 208.415 21.855 208.585 ;
        RECT 22.035 208.335 22.645 208.665 ;
        RECT 22.815 208.375 23.315 208.835 ;
        RECT 23.545 208.810 23.835 209.975 ;
        RECT 24.095 209.230 24.365 209.975 ;
        RECT 24.995 209.970 31.270 209.975 ;
        RECT 24.535 209.060 24.825 209.800 ;
        RECT 24.995 209.245 25.250 209.970 ;
        RECT 25.435 209.075 25.695 209.800 ;
        RECT 25.865 209.245 26.110 209.970 ;
        RECT 26.295 209.075 26.555 209.800 ;
        RECT 26.725 209.245 26.970 209.970 ;
        RECT 27.155 209.075 27.415 209.800 ;
        RECT 27.585 209.245 27.830 209.970 ;
        RECT 28.000 209.075 28.260 209.800 ;
        RECT 28.430 209.245 28.690 209.970 ;
        RECT 28.860 209.075 29.120 209.800 ;
        RECT 29.290 209.245 29.550 209.970 ;
        RECT 29.720 209.075 29.980 209.800 ;
        RECT 30.150 209.245 30.410 209.970 ;
        RECT 30.580 209.075 30.840 209.800 ;
        RECT 31.010 209.175 31.270 209.970 ;
        RECT 25.435 209.060 30.840 209.075 ;
        RECT 24.095 208.835 30.840 209.060 ;
        RECT 24.095 208.275 25.260 208.835 ;
        RECT 31.440 208.665 31.690 209.800 ;
        RECT 31.870 209.165 32.130 209.975 ;
        RECT 32.305 208.665 32.550 209.805 ;
        RECT 32.730 209.165 33.025 209.975 ;
        RECT 33.205 208.965 33.465 209.975 ;
        RECT 33.635 209.135 33.910 209.805 ;
        RECT 33.635 208.785 33.805 209.135 ;
        RECT 34.110 209.130 34.325 209.975 ;
        RECT 34.510 209.465 34.985 209.805 ;
        RECT 35.165 209.470 35.795 209.975 ;
        RECT 35.165 209.295 35.355 209.470 ;
        RECT 34.550 208.935 34.800 209.230 ;
        RECT 35.025 209.105 35.355 209.295 ;
        RECT 35.525 208.935 35.780 209.300 ;
        RECT 35.975 209.165 36.270 209.975 ;
        RECT 25.430 208.415 32.550 208.665 ;
        RECT 24.065 208.245 25.260 208.275 ;
        RECT 20.845 207.955 22.505 208.125 ;
        RECT 20.845 207.595 21.165 207.955 ;
        RECT 21.370 207.425 21.700 207.785 ;
        RECT 22.160 207.595 22.505 207.955 ;
        RECT 23.065 207.425 23.360 208.205 ;
        RECT 23.545 207.425 23.835 208.150 ;
        RECT 24.065 208.105 30.840 208.245 ;
        RECT 24.095 208.075 30.840 208.105 ;
        RECT 24.095 207.425 24.395 207.905 ;
        RECT 24.565 207.620 24.825 208.075 ;
        RECT 24.995 207.425 25.255 207.905 ;
        RECT 25.435 207.620 25.695 208.075 ;
        RECT 25.865 207.425 26.115 207.905 ;
        RECT 26.295 207.620 26.555 208.075 ;
        RECT 26.725 207.425 26.975 207.905 ;
        RECT 27.155 207.620 27.415 208.075 ;
        RECT 27.585 207.425 27.830 207.905 ;
        RECT 28.000 207.620 28.275 208.075 ;
        RECT 28.445 207.425 28.690 207.905 ;
        RECT 28.860 207.620 29.120 208.075 ;
        RECT 29.290 207.425 29.550 207.905 ;
        RECT 29.720 207.620 29.980 208.075 ;
        RECT 30.150 207.425 30.410 207.905 ;
        RECT 30.580 207.620 30.840 208.075 ;
        RECT 31.010 207.425 31.270 207.985 ;
        RECT 31.440 207.605 31.690 208.415 ;
        RECT 31.870 207.425 32.130 207.950 ;
        RECT 32.300 207.605 32.550 208.415 ;
        RECT 32.720 208.105 33.035 208.665 ;
        RECT 33.205 208.265 33.820 208.785 ;
        RECT 33.990 208.765 35.780 208.935 ;
        RECT 33.990 208.335 34.220 208.765 ;
        RECT 32.730 207.425 33.035 207.935 ;
        RECT 33.205 207.425 33.480 208.085 ;
        RECT 33.650 208.055 33.820 208.265 ;
        RECT 34.405 208.090 34.815 208.585 ;
        RECT 33.650 207.595 33.900 208.055 ;
        RECT 34.075 207.425 34.405 207.920 ;
        RECT 34.585 207.645 34.815 208.090 ;
        RECT 34.985 207.910 35.240 208.765 ;
        RECT 36.450 208.665 36.695 209.805 ;
        RECT 36.870 209.165 37.130 209.975 ;
        RECT 37.730 209.970 44.005 209.975 ;
        RECT 37.310 208.665 37.560 209.800 ;
        RECT 37.730 209.175 37.990 209.970 ;
        RECT 38.160 209.075 38.420 209.800 ;
        RECT 38.590 209.245 38.850 209.970 ;
        RECT 39.020 209.075 39.280 209.800 ;
        RECT 39.450 209.245 39.710 209.970 ;
        RECT 39.880 209.075 40.140 209.800 ;
        RECT 40.310 209.245 40.570 209.970 ;
        RECT 40.740 209.075 41.000 209.800 ;
        RECT 41.170 209.245 41.415 209.970 ;
        RECT 41.585 209.075 41.845 209.800 ;
        RECT 42.030 209.245 42.275 209.970 ;
        RECT 42.445 209.075 42.705 209.800 ;
        RECT 42.890 209.245 43.135 209.970 ;
        RECT 43.305 209.075 43.565 209.800 ;
        RECT 43.750 209.245 44.005 209.970 ;
        RECT 38.160 209.060 43.565 209.075 ;
        RECT 44.175 209.060 44.465 209.800 ;
        RECT 44.635 209.230 44.905 209.975 ;
        RECT 45.755 209.635 47.805 209.805 ;
        RECT 45.755 209.135 46.005 209.635 ;
        RECT 38.160 208.835 44.905 209.060 ;
        RECT 46.175 208.965 46.385 209.465 ;
        RECT 46.595 209.135 46.805 209.635 ;
        RECT 47.135 208.965 47.385 209.465 ;
        RECT 47.555 209.135 47.805 209.635 ;
        RECT 47.975 208.965 48.225 209.805 ;
        RECT 48.395 209.135 48.645 209.975 ;
        RECT 48.815 208.965 49.070 209.805 ;
        RECT 35.410 208.105 35.795 208.585 ;
        RECT 35.965 208.105 36.280 208.665 ;
        RECT 36.450 208.415 43.570 208.665 ;
        RECT 34.985 207.645 35.775 207.910 ;
        RECT 35.965 207.425 36.270 207.935 ;
        RECT 36.450 207.605 36.700 208.415 ;
        RECT 36.870 207.425 37.130 207.950 ;
        RECT 37.310 207.605 37.560 208.415 ;
        RECT 43.740 208.245 44.905 208.835 ;
        RECT 38.160 208.075 44.905 208.245 ;
        RECT 45.625 208.795 46.385 208.965 ;
        RECT 45.625 208.245 46.085 208.795 ;
        RECT 46.580 208.625 46.845 208.965 ;
        RECT 47.135 208.795 49.070 208.965 ;
        RECT 49.305 208.810 49.595 209.975 ;
        RECT 49.775 209.165 50.070 209.975 ;
        RECT 50.250 208.665 50.495 209.805 ;
        RECT 50.670 209.165 50.930 209.975 ;
        RECT 51.530 209.970 57.805 209.975 ;
        RECT 51.110 208.665 51.360 209.800 ;
        RECT 51.530 209.175 51.790 209.970 ;
        RECT 51.960 209.075 52.220 209.800 ;
        RECT 52.390 209.245 52.650 209.970 ;
        RECT 52.820 209.075 53.080 209.800 ;
        RECT 53.250 209.245 53.510 209.970 ;
        RECT 53.680 209.075 53.940 209.800 ;
        RECT 54.110 209.245 54.370 209.970 ;
        RECT 54.540 209.075 54.800 209.800 ;
        RECT 54.970 209.245 55.215 209.970 ;
        RECT 55.385 209.075 55.645 209.800 ;
        RECT 55.830 209.245 56.075 209.970 ;
        RECT 56.245 209.075 56.505 209.800 ;
        RECT 56.690 209.245 56.935 209.970 ;
        RECT 57.105 209.075 57.365 209.800 ;
        RECT 57.550 209.245 57.805 209.970 ;
        RECT 51.960 209.060 57.365 209.075 ;
        RECT 57.975 209.060 58.265 209.800 ;
        RECT 58.435 209.230 58.705 209.975 ;
        RECT 51.960 208.835 58.705 209.060 ;
        RECT 46.255 208.415 46.845 208.625 ;
        RECT 47.035 208.415 48.085 208.625 ;
        RECT 48.255 208.415 49.085 208.625 ;
        RECT 37.730 207.425 37.990 207.985 ;
        RECT 38.160 207.620 38.420 208.075 ;
        RECT 38.590 207.425 38.850 207.905 ;
        RECT 39.020 207.620 39.280 208.075 ;
        RECT 39.450 207.425 39.710 207.905 ;
        RECT 39.880 207.620 40.140 208.075 ;
        RECT 40.310 207.425 40.555 207.905 ;
        RECT 40.725 207.620 41.000 208.075 ;
        RECT 41.170 207.425 41.415 207.905 ;
        RECT 41.585 207.620 41.845 208.075 ;
        RECT 42.025 207.425 42.275 207.905 ;
        RECT 42.445 207.620 42.705 208.075 ;
        RECT 42.885 207.425 43.135 207.905 ;
        RECT 43.305 207.620 43.565 208.075 ;
        RECT 43.745 207.425 44.005 207.905 ;
        RECT 44.175 207.620 44.435 208.075 ;
        RECT 45.625 208.065 48.685 208.245 ;
        RECT 44.605 207.425 44.905 207.905 ;
        RECT 45.675 207.425 45.965 207.895 ;
        RECT 46.135 207.595 46.465 208.065 ;
        RECT 46.635 207.425 47.345 207.895 ;
        RECT 47.515 207.595 47.845 208.065 ;
        RECT 48.015 207.425 48.185 207.895 ;
        RECT 48.355 207.595 48.685 208.065 ;
        RECT 48.855 207.425 49.130 208.245 ;
        RECT 49.305 207.425 49.595 208.150 ;
        RECT 49.765 208.105 50.080 208.665 ;
        RECT 50.250 208.415 57.370 208.665 ;
        RECT 49.765 207.425 50.070 207.935 ;
        RECT 50.250 207.605 50.500 208.415 ;
        RECT 50.670 207.425 50.930 207.950 ;
        RECT 51.110 207.605 51.360 208.415 ;
        RECT 57.540 208.245 58.705 208.835 ;
        RECT 58.970 208.825 59.230 209.975 ;
        RECT 59.405 208.900 59.660 209.805 ;
        RECT 59.830 209.215 60.160 209.975 ;
        RECT 60.375 209.045 60.545 209.805 ;
        RECT 61.010 209.535 61.340 209.975 ;
        RECT 61.510 209.365 61.745 209.805 ;
        RECT 61.930 209.595 62.260 209.975 ;
        RECT 62.470 209.365 62.815 209.805 ;
        RECT 51.960 208.075 58.705 208.245 ;
        RECT 51.530 207.425 51.790 207.985 ;
        RECT 51.960 207.620 52.220 208.075 ;
        RECT 52.390 207.425 52.650 207.905 ;
        RECT 52.820 207.620 53.080 208.075 ;
        RECT 53.250 207.425 53.510 207.905 ;
        RECT 53.680 207.620 53.940 208.075 ;
        RECT 54.110 207.425 54.355 207.905 ;
        RECT 54.525 207.620 54.800 208.075 ;
        RECT 54.970 207.425 55.215 207.905 ;
        RECT 55.385 207.620 55.645 208.075 ;
        RECT 55.825 207.425 56.075 207.905 ;
        RECT 56.245 207.620 56.505 208.075 ;
        RECT 56.685 207.425 56.935 207.905 ;
        RECT 57.105 207.620 57.365 208.075 ;
        RECT 57.545 207.425 57.805 207.905 ;
        RECT 57.975 207.620 58.235 208.075 ;
        RECT 58.405 207.425 58.705 207.905 ;
        RECT 58.970 207.425 59.230 208.265 ;
        RECT 59.405 208.170 59.575 208.900 ;
        RECT 59.830 208.875 60.545 209.045 ;
        RECT 60.805 209.125 62.815 209.365 ;
        RECT 59.830 208.665 60.000 208.875 ;
        RECT 59.745 208.335 60.000 208.665 ;
        RECT 59.405 207.595 59.660 208.170 ;
        RECT 59.830 208.145 60.000 208.335 ;
        RECT 60.280 208.325 60.635 208.695 ;
        RECT 60.805 208.225 61.035 209.125 ;
        RECT 62.990 208.955 63.335 209.710 ;
        RECT 63.505 209.135 63.835 209.975 ;
        RECT 64.225 209.305 64.505 209.975 ;
        RECT 61.205 208.415 61.535 208.955 ;
        RECT 59.830 207.975 60.545 208.145 ;
        RECT 59.830 207.425 60.160 207.805 ;
        RECT 60.375 207.595 60.545 207.975 ;
        RECT 60.805 207.595 61.410 208.225 ;
        RECT 61.745 207.595 62.075 208.955 ;
        RECT 62.245 208.335 62.535 208.955 ;
        RECT 62.705 208.335 63.335 208.955 ;
        RECT 63.505 208.345 63.835 208.955 ;
        RECT 64.025 208.665 64.340 209.105 ;
        RECT 64.675 209.085 64.975 209.635 ;
        RECT 65.185 209.255 65.515 209.975 ;
        RECT 65.705 209.255 66.155 209.805 ;
        RECT 64.675 208.915 65.615 209.085 ;
        RECT 65.445 208.665 65.615 208.915 ;
        RECT 64.025 208.415 64.715 208.665 ;
        RECT 64.945 208.415 65.275 208.665 ;
        RECT 65.445 208.335 65.735 208.665 ;
        RECT 65.445 208.245 65.615 208.335 ;
        RECT 62.470 207.965 63.835 208.165 ;
        RECT 62.470 207.595 62.815 207.965 ;
        RECT 63.005 207.425 63.335 207.795 ;
        RECT 63.505 207.595 63.835 207.965 ;
        RECT 64.225 208.055 65.615 208.245 ;
        RECT 64.225 207.695 64.555 208.055 ;
        RECT 65.905 207.885 66.155 209.255 ;
        RECT 66.325 208.835 66.615 209.975 ;
        RECT 66.785 209.465 67.975 209.755 ;
        RECT 66.805 209.125 67.975 209.295 ;
        RECT 68.145 209.175 68.425 209.975 ;
        RECT 66.805 208.835 67.130 209.125 ;
        RECT 67.805 209.005 67.975 209.125 ;
        RECT 67.300 208.665 67.495 208.955 ;
        RECT 67.805 208.835 68.465 209.005 ;
        RECT 68.635 208.835 68.910 209.805 ;
        RECT 69.125 208.835 69.355 209.975 ;
        RECT 68.295 208.665 68.465 208.835 ;
        RECT 66.785 208.335 67.130 208.665 ;
        RECT 67.300 208.335 68.125 208.665 ;
        RECT 68.295 208.335 68.570 208.665 ;
        RECT 65.185 207.425 65.435 207.885 ;
        RECT 65.605 207.595 66.155 207.885 ;
        RECT 66.325 207.425 66.615 208.225 ;
        RECT 68.295 208.165 68.465 208.335 ;
        RECT 66.800 207.995 68.465 208.165 ;
        RECT 68.740 208.100 68.910 208.835 ;
        RECT 69.525 208.825 69.855 209.805 ;
        RECT 70.025 208.835 70.235 209.975 ;
        RECT 69.105 208.415 69.435 208.665 ;
        RECT 66.800 207.645 67.055 207.995 ;
        RECT 67.225 207.425 67.555 207.825 ;
        RECT 67.725 207.645 67.895 207.995 ;
        RECT 68.065 207.425 68.445 207.825 ;
        RECT 68.635 207.755 68.910 208.100 ;
        RECT 69.125 207.425 69.355 208.245 ;
        RECT 69.605 208.225 69.855 208.825 ;
        RECT 71.385 208.820 71.725 209.805 ;
        RECT 71.895 209.545 72.305 209.975 ;
        RECT 73.050 209.555 73.380 209.975 ;
        RECT 73.550 209.375 73.875 209.805 ;
        RECT 71.895 209.205 73.875 209.375 ;
        RECT 69.525 207.595 69.855 208.225 ;
        RECT 70.025 207.425 70.235 208.245 ;
        RECT 71.385 208.165 71.640 208.820 ;
        RECT 71.895 208.665 72.160 209.205 ;
        RECT 72.375 208.865 73.000 209.035 ;
        RECT 71.810 208.335 72.160 208.665 ;
        RECT 72.330 208.335 72.660 208.665 ;
        RECT 72.830 208.165 73.000 208.865 ;
        RECT 71.385 207.790 71.745 208.165 ;
        RECT 71.445 207.765 71.615 207.790 ;
        RECT 72.010 207.425 72.180 208.165 ;
        RECT 72.460 207.995 73.000 208.165 ;
        RECT 73.170 208.795 73.875 209.205 ;
        RECT 74.350 208.875 74.680 209.975 ;
        RECT 75.065 208.810 75.355 209.975 ;
        RECT 75.535 209.005 75.865 209.790 ;
        RECT 75.535 208.835 76.215 209.005 ;
        RECT 76.395 208.835 76.725 209.975 ;
        RECT 76.905 208.900 77.175 209.805 ;
        RECT 77.345 209.215 77.675 209.975 ;
        RECT 77.855 209.045 78.035 209.805 ;
        RECT 72.460 207.790 72.630 207.995 ;
        RECT 73.170 207.595 73.340 208.795 ;
        RECT 73.510 208.415 74.080 208.625 ;
        RECT 74.250 208.415 74.895 208.625 ;
        RECT 75.525 208.415 75.875 208.665 ;
        RECT 73.570 208.075 74.740 208.245 ;
        RECT 76.045 208.235 76.215 208.835 ;
        RECT 76.385 208.415 76.735 208.665 ;
        RECT 73.570 207.595 73.900 208.075 ;
        RECT 74.070 207.425 74.240 207.895 ;
        RECT 74.410 207.610 74.740 208.075 ;
        RECT 75.065 207.425 75.355 208.150 ;
        RECT 75.545 207.425 75.785 208.235 ;
        RECT 75.955 207.595 76.285 208.235 ;
        RECT 76.455 207.425 76.725 208.235 ;
        RECT 76.905 208.100 77.085 208.900 ;
        RECT 77.360 208.875 78.035 209.045 ;
        RECT 77.360 208.730 77.530 208.875 ;
        RECT 78.325 208.835 78.555 209.975 ;
        RECT 78.725 208.825 79.055 209.805 ;
        RECT 79.225 208.835 79.435 209.975 ;
        RECT 79.665 208.900 79.935 209.805 ;
        RECT 80.105 209.215 80.435 209.975 ;
        RECT 80.615 209.045 80.795 209.805 ;
        RECT 77.255 208.400 77.530 208.730 ;
        RECT 77.360 208.145 77.530 208.400 ;
        RECT 77.755 208.325 78.095 208.695 ;
        RECT 78.305 208.415 78.635 208.665 ;
        RECT 76.905 207.595 77.165 208.100 ;
        RECT 77.360 207.975 78.025 208.145 ;
        RECT 77.345 207.425 77.675 207.805 ;
        RECT 77.855 207.595 78.025 207.975 ;
        RECT 78.325 207.425 78.555 208.245 ;
        RECT 78.805 208.225 79.055 208.825 ;
        RECT 78.725 207.595 79.055 208.225 ;
        RECT 79.225 207.425 79.435 208.245 ;
        RECT 79.665 208.100 79.845 208.900 ;
        RECT 80.120 208.875 80.795 209.045 ;
        RECT 81.510 209.405 81.830 209.805 ;
        RECT 81.510 208.955 81.680 209.405 ;
        RECT 82.000 209.175 82.310 209.975 ;
        RECT 82.480 209.345 82.810 209.805 ;
        RECT 82.980 209.515 83.150 209.975 ;
        RECT 83.320 209.345 83.650 209.805 ;
        RECT 83.820 209.515 84.070 209.975 ;
        RECT 84.260 209.515 84.510 209.975 ;
        RECT 82.480 209.295 83.650 209.345 ;
        RECT 84.680 209.345 84.930 209.805 ;
        RECT 85.180 209.515 85.470 209.975 ;
        RECT 84.680 209.295 85.470 209.345 ;
        RECT 82.480 209.125 85.470 209.295 ;
        RECT 80.120 208.730 80.290 208.875 ;
        RECT 80.015 208.400 80.290 208.730 ;
        RECT 81.510 208.785 85.070 208.955 ;
        RECT 80.120 208.145 80.290 208.400 ;
        RECT 80.515 208.325 80.855 208.695 ;
        RECT 79.665 207.595 79.925 208.100 ;
        RECT 80.120 207.975 80.785 208.145 ;
        RECT 80.105 207.425 80.435 207.805 ;
        RECT 80.615 207.595 80.785 207.975 ;
        RECT 81.510 207.995 81.680 208.785 ;
        RECT 81.850 208.415 82.200 208.615 ;
        RECT 82.480 208.415 83.160 208.615 ;
        RECT 83.370 208.415 84.560 208.615 ;
        RECT 84.740 208.415 85.070 208.785 ;
        RECT 85.270 208.275 85.470 209.125 ;
        RECT 85.740 208.780 85.910 209.975 ;
        RECT 86.080 208.835 86.355 209.805 ;
        RECT 86.565 209.175 86.845 209.975 ;
        RECT 87.015 209.465 87.655 209.795 ;
        RECT 87.880 209.545 88.625 209.715 ;
        RECT 89.315 209.545 89.645 209.975 ;
        RECT 87.880 209.295 88.050 209.545 ;
        RECT 89.815 209.375 90.075 209.795 ;
        RECT 87.015 209.125 88.050 209.295 ;
        RECT 88.220 209.205 90.075 209.375 ;
        RECT 87.015 209.005 87.185 209.125 ;
        RECT 86.525 208.835 87.185 209.005 ;
        RECT 88.220 208.925 88.390 209.205 ;
        RECT 85.245 208.245 85.470 208.275 ;
        RECT 81.510 207.595 81.830 207.995 ;
        RECT 82.000 207.425 82.310 208.245 ;
        RECT 82.480 208.055 84.170 208.245 ;
        RECT 82.480 207.595 82.810 208.055 ;
        RECT 83.420 207.975 84.170 208.055 ;
        RECT 82.980 207.425 83.230 207.885 ;
        RECT 84.340 207.805 84.510 208.245 ;
        RECT 84.680 207.975 85.470 208.245 ;
        RECT 83.420 207.595 85.470 207.805 ;
        RECT 85.740 207.425 85.910 208.365 ;
        RECT 86.080 208.100 86.250 208.835 ;
        RECT 86.525 208.665 86.695 208.835 ;
        RECT 87.740 208.755 88.390 208.925 ;
        RECT 88.560 208.865 89.165 209.035 ;
        RECT 86.420 208.335 86.695 208.665 ;
        RECT 86.865 208.335 87.520 208.665 ;
        RECT 87.740 208.335 87.910 208.755 ;
        RECT 88.560 208.585 88.750 208.865 ;
        RECT 88.305 208.415 88.750 208.585 ;
        RECT 86.525 208.165 86.695 208.335 ;
        RECT 88.560 208.165 88.750 208.415 ;
        RECT 88.920 208.335 89.210 208.665 ;
        RECT 89.380 208.335 89.730 209.035 ;
        RECT 89.900 208.165 90.075 209.205 ;
        RECT 90.335 209.045 90.505 209.805 ;
        RECT 90.720 209.215 91.050 209.975 ;
        RECT 90.335 208.875 91.050 209.045 ;
        RECT 91.220 208.900 91.475 209.805 ;
        RECT 90.245 208.325 90.600 208.695 ;
        RECT 90.880 208.665 91.050 208.875 ;
        RECT 90.880 208.335 91.135 208.665 ;
        RECT 86.080 207.755 86.355 208.100 ;
        RECT 86.525 207.995 88.135 208.165 ;
        RECT 88.560 207.995 89.080 208.165 ;
        RECT 86.545 207.425 86.925 207.825 ;
        RECT 87.095 207.645 87.265 207.995 ;
        RECT 87.435 207.425 87.765 207.825 ;
        RECT 87.965 207.645 88.135 207.995 ;
        RECT 88.310 207.425 88.665 207.825 ;
        RECT 88.910 207.790 89.080 207.995 ;
        RECT 89.330 207.425 89.500 208.165 ;
        RECT 89.755 207.790 90.075 208.165 ;
        RECT 90.880 208.145 91.050 208.335 ;
        RECT 91.305 208.170 91.475 208.900 ;
        RECT 91.650 208.825 91.910 209.975 ;
        RECT 92.175 209.045 92.345 209.805 ;
        RECT 92.560 209.215 92.890 209.975 ;
        RECT 92.175 208.875 92.890 209.045 ;
        RECT 93.060 208.900 93.315 209.805 ;
        RECT 92.085 208.325 92.440 208.695 ;
        RECT 92.720 208.665 92.890 208.875 ;
        RECT 92.720 208.335 92.975 208.665 ;
        RECT 90.335 207.975 91.050 208.145 ;
        RECT 90.335 207.595 90.505 207.975 ;
        RECT 90.720 207.425 91.050 207.805 ;
        RECT 91.220 207.595 91.475 208.170 ;
        RECT 91.650 207.425 91.910 208.265 ;
        RECT 92.720 208.145 92.890 208.335 ;
        RECT 93.145 208.170 93.315 208.900 ;
        RECT 93.490 208.825 93.750 209.975 ;
        RECT 93.930 209.515 94.220 209.975 ;
        RECT 94.470 209.345 94.720 209.805 ;
        RECT 94.890 209.515 95.140 209.975 ;
        RECT 95.330 209.515 95.580 209.975 ;
        RECT 93.930 209.295 94.720 209.345 ;
        RECT 95.750 209.345 96.080 209.805 ;
        RECT 96.250 209.515 96.420 209.975 ;
        RECT 96.590 209.345 96.920 209.805 ;
        RECT 95.750 209.295 96.920 209.345 ;
        RECT 93.930 209.125 96.920 209.295 ;
        RECT 97.090 209.175 97.400 209.975 ;
        RECT 97.570 209.405 97.890 209.805 ;
        RECT 93.930 208.275 94.130 209.125 ;
        RECT 97.720 208.955 97.890 209.405 ;
        RECT 94.330 208.785 97.890 208.955 ;
        RECT 98.155 209.045 98.325 209.805 ;
        RECT 98.540 209.215 98.870 209.975 ;
        RECT 98.155 208.875 98.870 209.045 ;
        RECT 99.040 208.900 99.295 209.805 ;
        RECT 94.330 208.415 94.660 208.785 ;
        RECT 94.840 208.415 96.030 208.615 ;
        RECT 96.240 208.415 96.920 208.615 ;
        RECT 97.200 208.415 97.550 208.615 ;
        RECT 92.175 207.975 92.890 208.145 ;
        RECT 92.175 207.595 92.345 207.975 ;
        RECT 92.560 207.425 92.890 207.805 ;
        RECT 93.060 207.595 93.315 208.170 ;
        RECT 93.490 207.425 93.750 208.265 ;
        RECT 93.930 208.245 94.155 208.275 ;
        RECT 93.930 207.975 94.720 208.245 ;
        RECT 94.890 207.805 95.060 208.245 ;
        RECT 95.230 208.055 96.920 208.245 ;
        RECT 95.230 207.975 95.980 208.055 ;
        RECT 93.930 207.595 95.980 207.805 ;
        RECT 96.170 207.425 96.420 207.885 ;
        RECT 96.590 207.595 96.920 208.055 ;
        RECT 97.090 207.425 97.400 208.245 ;
        RECT 97.720 207.995 97.890 208.785 ;
        RECT 98.065 208.325 98.420 208.695 ;
        RECT 98.700 208.665 98.870 208.875 ;
        RECT 98.700 208.335 98.955 208.665 ;
        RECT 98.700 208.145 98.870 208.335 ;
        RECT 99.125 208.170 99.295 208.900 ;
        RECT 99.470 208.825 99.730 209.975 ;
        RECT 100.825 208.810 101.115 209.975 ;
        RECT 102.210 209.540 107.555 209.975 ;
        RECT 107.730 209.540 113.075 209.975 ;
        RECT 113.250 209.540 118.595 209.975 ;
        RECT 118.770 209.540 124.115 209.975 ;
        RECT 103.800 208.290 104.150 209.540 ;
        RECT 97.570 207.595 97.890 207.995 ;
        RECT 98.155 207.975 98.870 208.145 ;
        RECT 98.155 207.595 98.325 207.975 ;
        RECT 98.540 207.425 98.870 207.805 ;
        RECT 99.040 207.595 99.295 208.170 ;
        RECT 99.470 207.425 99.730 208.265 ;
        RECT 100.825 207.425 101.115 208.150 ;
        RECT 105.630 207.970 105.970 208.800 ;
        RECT 109.320 208.290 109.670 209.540 ;
        RECT 111.150 207.970 111.490 208.800 ;
        RECT 114.840 208.290 115.190 209.540 ;
        RECT 116.670 207.970 117.010 208.800 ;
        RECT 120.360 208.290 120.710 209.540 ;
        RECT 124.475 209.250 124.805 209.975 ;
        RECT 122.190 207.970 122.530 208.800 ;
        RECT 102.210 207.425 107.555 207.970 ;
        RECT 107.730 207.425 113.075 207.970 ;
        RECT 113.250 207.425 118.595 207.970 ;
        RECT 118.770 207.425 124.115 207.970 ;
        RECT 124.285 207.595 124.805 209.080 ;
        RECT 124.975 208.255 125.495 209.805 ;
        RECT 125.665 208.885 126.875 209.975 ;
        RECT 125.665 208.345 126.185 208.885 ;
        RECT 126.355 208.175 126.875 208.715 ;
        RECT 124.975 207.425 125.315 208.085 ;
        RECT 125.665 207.425 126.875 208.175 ;
        RECT 14.260 207.255 126.960 207.425 ;
        RECT 14.345 206.505 15.555 207.255 ;
        RECT 15.775 206.785 16.065 207.255 ;
        RECT 16.235 206.615 16.565 207.085 ;
        RECT 16.735 206.785 16.905 207.255 ;
        RECT 17.075 206.615 17.405 207.085 ;
        RECT 16.235 206.605 17.405 206.615 ;
        RECT 14.345 205.965 14.865 206.505 ;
        RECT 15.805 206.435 17.405 206.605 ;
        RECT 17.575 206.435 17.850 207.255 ;
        RECT 18.115 206.775 18.415 207.255 ;
        RECT 18.585 206.605 18.845 207.060 ;
        RECT 19.015 206.775 19.275 207.255 ;
        RECT 19.455 206.605 19.715 207.060 ;
        RECT 19.885 206.775 20.135 207.255 ;
        RECT 20.315 206.605 20.575 207.060 ;
        RECT 20.745 206.775 20.995 207.255 ;
        RECT 21.175 206.605 21.435 207.060 ;
        RECT 21.605 206.775 21.850 207.255 ;
        RECT 22.020 206.605 22.295 207.060 ;
        RECT 22.465 206.775 22.710 207.255 ;
        RECT 22.880 206.605 23.140 207.060 ;
        RECT 23.310 206.775 23.570 207.255 ;
        RECT 23.740 206.605 24.000 207.060 ;
        RECT 24.170 206.775 24.430 207.255 ;
        RECT 24.600 206.605 24.860 207.060 ;
        RECT 25.030 206.695 25.290 207.255 ;
        RECT 18.115 206.435 24.860 206.605 ;
        RECT 15.035 205.795 15.555 206.335 ;
        RECT 14.345 204.705 15.555 205.795 ;
        RECT 15.805 205.895 16.020 206.435 ;
        RECT 16.190 206.065 16.960 206.265 ;
        RECT 17.130 206.065 17.850 206.265 ;
        RECT 15.805 205.675 16.565 205.895 ;
        RECT 15.765 205.045 16.065 205.505 ;
        RECT 16.235 205.215 16.565 205.675 ;
        RECT 16.735 205.675 17.850 205.885 ;
        RECT 16.735 205.045 16.905 205.675 ;
        RECT 15.765 204.875 16.905 205.045 ;
        RECT 17.075 204.705 17.405 205.505 ;
        RECT 17.575 204.875 17.850 205.675 ;
        RECT 18.115 205.845 19.280 206.435 ;
        RECT 25.460 206.265 25.710 207.075 ;
        RECT 25.890 206.730 26.150 207.255 ;
        RECT 26.320 206.265 26.570 207.075 ;
        RECT 26.750 206.745 27.055 207.255 ;
        RECT 27.315 206.775 27.615 207.255 ;
        RECT 27.785 206.605 28.045 207.060 ;
        RECT 28.215 206.775 28.475 207.255 ;
        RECT 28.655 206.605 28.915 207.060 ;
        RECT 29.085 206.775 29.335 207.255 ;
        RECT 29.515 206.605 29.775 207.060 ;
        RECT 29.945 206.775 30.195 207.255 ;
        RECT 30.375 206.605 30.635 207.060 ;
        RECT 30.805 206.775 31.050 207.255 ;
        RECT 31.220 206.605 31.495 207.060 ;
        RECT 31.665 206.775 31.910 207.255 ;
        RECT 32.080 206.605 32.340 207.060 ;
        RECT 32.510 206.775 32.770 207.255 ;
        RECT 32.940 206.605 33.200 207.060 ;
        RECT 33.370 206.775 33.630 207.255 ;
        RECT 33.800 206.605 34.060 207.060 ;
        RECT 34.230 206.695 34.490 207.255 ;
        RECT 19.450 206.015 26.570 206.265 ;
        RECT 26.740 206.015 27.055 206.575 ;
        RECT 27.315 206.435 34.060 206.605 ;
        RECT 18.115 205.620 24.860 205.845 ;
        RECT 18.115 204.705 18.385 205.450 ;
        RECT 18.555 204.880 18.845 205.620 ;
        RECT 19.455 205.605 24.860 205.620 ;
        RECT 19.015 204.710 19.270 205.435 ;
        RECT 19.455 204.880 19.715 205.605 ;
        RECT 19.885 204.710 20.130 205.435 ;
        RECT 20.315 204.880 20.575 205.605 ;
        RECT 20.745 204.710 20.990 205.435 ;
        RECT 21.175 204.880 21.435 205.605 ;
        RECT 21.605 204.710 21.850 205.435 ;
        RECT 22.020 204.880 22.280 205.605 ;
        RECT 22.450 204.710 22.710 205.435 ;
        RECT 22.880 204.880 23.140 205.605 ;
        RECT 23.310 204.710 23.570 205.435 ;
        RECT 23.740 204.880 24.000 205.605 ;
        RECT 24.170 204.710 24.430 205.435 ;
        RECT 24.600 204.880 24.860 205.605 ;
        RECT 25.030 204.710 25.290 205.505 ;
        RECT 25.460 204.880 25.710 206.015 ;
        RECT 19.015 204.705 25.290 204.710 ;
        RECT 25.890 204.705 26.150 205.515 ;
        RECT 26.325 204.875 26.570 206.015 ;
        RECT 27.315 205.845 28.480 206.435 ;
        RECT 34.660 206.265 34.910 207.075 ;
        RECT 35.090 206.730 35.350 207.255 ;
        RECT 35.520 206.265 35.770 207.075 ;
        RECT 35.950 206.745 36.255 207.255 ;
        RECT 28.650 206.015 35.770 206.265 ;
        RECT 35.940 206.015 36.255 206.575 ;
        RECT 36.425 206.530 36.715 207.255 ;
        RECT 37.345 206.745 37.650 207.255 ;
        RECT 37.345 206.015 37.660 206.575 ;
        RECT 37.830 206.265 38.080 207.075 ;
        RECT 38.250 206.730 38.510 207.255 ;
        RECT 38.690 206.265 38.940 207.075 ;
        RECT 39.110 206.695 39.370 207.255 ;
        RECT 39.540 206.605 39.800 207.060 ;
        RECT 39.970 206.775 40.230 207.255 ;
        RECT 40.400 206.605 40.660 207.060 ;
        RECT 40.830 206.775 41.090 207.255 ;
        RECT 41.260 206.605 41.520 207.060 ;
        RECT 41.690 206.775 41.935 207.255 ;
        RECT 42.105 206.605 42.380 207.060 ;
        RECT 42.550 206.775 42.795 207.255 ;
        RECT 42.965 206.605 43.225 207.060 ;
        RECT 43.405 206.775 43.655 207.255 ;
        RECT 43.825 206.605 44.085 207.060 ;
        RECT 44.265 206.775 44.515 207.255 ;
        RECT 44.685 206.605 44.945 207.060 ;
        RECT 45.125 206.775 45.385 207.255 ;
        RECT 45.555 206.605 45.815 207.060 ;
        RECT 45.985 206.775 46.285 207.255 ;
        RECT 46.590 206.895 46.920 207.255 ;
        RECT 47.090 206.725 47.420 207.085 ;
        RECT 47.590 206.815 47.825 207.255 ;
        RECT 48.415 206.875 48.750 207.255 ;
        RECT 49.710 206.915 50.045 207.085 ;
        RECT 39.540 206.435 46.285 206.605 ;
        RECT 37.830 206.015 44.950 206.265 ;
        RECT 27.315 205.620 34.060 205.845 ;
        RECT 26.750 204.705 27.045 205.515 ;
        RECT 27.315 204.705 27.585 205.450 ;
        RECT 27.755 204.880 28.045 205.620 ;
        RECT 28.655 205.605 34.060 205.620 ;
        RECT 28.215 204.710 28.470 205.435 ;
        RECT 28.655 204.880 28.915 205.605 ;
        RECT 29.085 204.710 29.330 205.435 ;
        RECT 29.515 204.880 29.775 205.605 ;
        RECT 29.945 204.710 30.190 205.435 ;
        RECT 30.375 204.880 30.635 205.605 ;
        RECT 30.805 204.710 31.050 205.435 ;
        RECT 31.220 204.880 31.480 205.605 ;
        RECT 31.650 204.710 31.910 205.435 ;
        RECT 32.080 204.880 32.340 205.605 ;
        RECT 32.510 204.710 32.770 205.435 ;
        RECT 32.940 204.880 33.200 205.605 ;
        RECT 33.370 204.710 33.630 205.435 ;
        RECT 33.800 204.880 34.060 205.605 ;
        RECT 34.230 204.710 34.490 205.505 ;
        RECT 34.660 204.880 34.910 206.015 ;
        RECT 28.215 204.705 34.490 204.710 ;
        RECT 35.090 204.705 35.350 205.515 ;
        RECT 35.525 204.875 35.770 206.015 ;
        RECT 35.950 204.705 36.245 205.515 ;
        RECT 36.425 204.705 36.715 205.870 ;
        RECT 37.355 204.705 37.650 205.515 ;
        RECT 37.830 204.875 38.075 206.015 ;
        RECT 38.250 204.705 38.510 205.515 ;
        RECT 38.690 204.880 38.940 206.015 ;
        RECT 45.120 205.845 46.285 206.435 ;
        RECT 39.540 205.620 46.285 205.845 ;
        RECT 46.600 206.555 47.420 206.725 ;
        RECT 39.540 205.605 44.945 205.620 ;
        RECT 39.110 204.710 39.370 205.505 ;
        RECT 39.540 204.880 39.800 205.605 ;
        RECT 39.970 204.710 40.230 205.435 ;
        RECT 40.400 204.880 40.660 205.605 ;
        RECT 40.830 204.710 41.090 205.435 ;
        RECT 41.260 204.880 41.520 205.605 ;
        RECT 41.690 204.710 41.950 205.435 ;
        RECT 42.120 204.880 42.380 205.605 ;
        RECT 42.550 204.710 42.795 205.435 ;
        RECT 42.965 204.880 43.225 205.605 ;
        RECT 43.410 204.710 43.655 205.435 ;
        RECT 43.825 204.880 44.085 205.605 ;
        RECT 44.270 204.710 44.515 205.435 ;
        RECT 44.685 204.880 44.945 205.605 ;
        RECT 45.130 204.710 45.385 205.435 ;
        RECT 45.555 204.880 45.845 205.620 ;
        RECT 39.110 204.705 45.385 204.710 ;
        RECT 46.015 204.705 46.285 205.450 ;
        RECT 46.600 205.435 46.795 206.555 ;
        RECT 47.990 206.515 49.260 206.705 ;
        RECT 49.430 206.515 50.045 206.915 ;
        RECT 50.685 206.755 50.945 207.085 ;
        RECT 51.115 206.755 51.365 207.255 ;
        RECT 46.965 206.015 47.645 206.345 ;
        RECT 47.815 206.015 48.150 206.345 ;
        RECT 48.320 206.235 48.610 206.345 ;
        RECT 48.320 206.065 48.615 206.235 ;
        RECT 48.320 206.015 48.610 206.065 ;
        RECT 48.900 206.015 49.260 206.345 ;
        RECT 47.475 205.830 47.645 206.015 ;
        RECT 49.430 205.830 49.610 206.515 ;
        RECT 49.780 206.015 50.055 206.345 ;
        RECT 47.475 205.575 50.050 205.830 ;
        RECT 46.600 205.265 47.330 205.435 ;
        RECT 46.640 204.705 46.970 205.085 ;
        RECT 47.140 204.875 47.330 205.265 ;
        RECT 47.510 204.705 47.940 205.405 ;
        RECT 48.445 204.875 49.115 205.575 ;
        RECT 49.285 204.705 49.615 205.405 ;
        RECT 49.785 204.875 50.050 205.575 ;
        RECT 50.685 205.425 50.855 206.755 ;
        RECT 51.025 206.035 51.375 206.575 ;
        RECT 51.545 205.935 51.850 206.915 ;
        RECT 52.025 206.235 52.290 206.920 ;
        RECT 53.020 206.705 53.190 207.085 ;
        RECT 53.460 206.875 53.790 207.255 ;
        RECT 52.795 206.535 53.785 206.705 ;
        RECT 52.025 206.065 52.295 206.235 ;
        RECT 52.455 205.765 52.625 205.940 ;
        RECT 51.445 205.595 52.625 205.765 ;
        RECT 51.445 205.425 51.615 205.595 ;
        RECT 52.795 205.425 52.965 206.535 ;
        RECT 53.135 206.015 53.445 206.345 ;
        RECT 53.615 206.015 53.785 206.535 ;
        RECT 50.685 205.255 51.615 205.425 ;
        RECT 51.785 205.255 52.965 205.425 ;
        RECT 53.275 205.455 53.445 206.015 ;
        RECT 53.960 205.795 54.185 207.085 ;
        RECT 54.355 206.875 54.685 207.255 ;
        RECT 54.855 206.705 55.025 207.085 ;
        RECT 54.530 206.535 55.025 206.705 ;
        RECT 55.285 206.645 55.635 207.085 ;
        RECT 55.805 206.815 55.975 207.255 ;
        RECT 56.145 206.875 57.340 207.085 ;
        RECT 56.145 206.645 56.395 206.875 ;
        RECT 53.880 205.625 54.210 205.795 ;
        RECT 54.530 205.455 54.700 206.535 ;
        RECT 55.285 206.435 56.395 206.645 ;
        RECT 56.565 206.535 56.895 206.705 ;
        RECT 56.565 206.435 56.890 206.535 ;
        RECT 57.065 206.435 57.340 206.875 ;
        RECT 57.575 206.515 57.905 207.255 ;
        RECT 58.075 206.500 58.310 206.830 ;
        RECT 54.870 206.235 55.050 206.345 ;
        RECT 54.870 206.065 55.055 206.235 ;
        RECT 55.285 206.065 56.430 206.265 ;
        RECT 54.870 205.705 55.050 206.065 ;
        RECT 53.275 205.285 55.025 205.455 ;
        RECT 50.685 204.875 50.945 205.255 ;
        RECT 51.115 204.705 51.445 205.085 ;
        RECT 51.785 204.875 51.955 205.255 ;
        RECT 52.125 204.705 52.465 205.085 ;
        RECT 52.635 204.875 52.805 205.255 ;
        RECT 53.040 204.705 53.710 205.085 ;
        RECT 54.355 204.705 54.685 205.085 ;
        RECT 54.855 204.875 55.025 205.285 ;
        RECT 55.285 204.705 55.615 205.845 ;
        RECT 55.785 205.505 56.060 205.845 ;
        RECT 56.240 205.685 56.430 206.065 ;
        RECT 56.610 205.555 56.890 206.435 ;
        RECT 57.060 205.845 57.390 206.265 ;
        RECT 57.620 206.015 57.965 206.345 ;
        RECT 58.140 205.845 58.310 206.500 ;
        RECT 57.060 205.675 58.310 205.845 ;
        RECT 56.610 205.505 56.895 205.555 ;
        RECT 55.785 205.335 57.385 205.505 ;
        RECT 55.785 204.875 56.140 205.335 ;
        RECT 56.310 204.705 56.885 205.165 ;
        RECT 57.055 204.875 57.385 205.335 ;
        RECT 57.585 204.705 57.840 205.505 ;
        RECT 58.010 205.480 58.310 205.675 ;
        RECT 58.965 206.455 59.570 207.085 ;
        RECT 58.965 205.555 59.195 206.455 ;
        RECT 59.365 205.725 59.695 206.265 ;
        RECT 59.905 205.725 60.235 207.085 ;
        RECT 60.630 206.715 60.975 207.085 ;
        RECT 61.165 206.885 61.495 207.255 ;
        RECT 61.665 206.715 61.995 207.085 ;
        RECT 60.630 206.515 61.995 206.715 ;
        RECT 62.185 206.530 62.475 207.255 ;
        RECT 63.565 206.515 64.005 207.075 ;
        RECT 64.175 206.515 64.625 207.255 ;
        RECT 64.795 206.685 64.965 207.085 ;
        RECT 65.135 206.855 65.555 207.255 ;
        RECT 65.725 206.685 65.955 207.085 ;
        RECT 64.795 206.515 65.955 206.685 ;
        RECT 66.125 206.515 66.615 207.085 ;
        RECT 66.845 206.890 67.015 206.915 ;
        RECT 60.405 205.725 60.695 206.345 ;
        RECT 60.865 205.725 61.495 206.345 ;
        RECT 61.665 205.725 61.995 206.335 ;
        RECT 58.965 205.315 60.975 205.555 ;
        RECT 59.170 204.705 59.500 205.145 ;
        RECT 59.670 204.875 59.905 205.315 ;
        RECT 60.090 204.705 60.420 205.085 ;
        RECT 60.630 204.875 60.975 205.315 ;
        RECT 61.150 204.970 61.495 205.725 ;
        RECT 61.665 204.705 61.995 205.545 ;
        RECT 62.185 204.705 62.475 205.870 ;
        RECT 63.565 205.505 63.875 206.515 ;
        RECT 64.045 205.895 64.215 206.345 ;
        RECT 64.385 206.065 64.775 206.345 ;
        RECT 64.960 206.015 65.205 206.345 ;
        RECT 64.045 205.725 64.835 205.895 ;
        RECT 63.565 204.875 64.005 205.505 ;
        RECT 64.180 204.705 64.495 205.555 ;
        RECT 64.665 205.045 64.835 205.725 ;
        RECT 65.005 205.215 65.205 206.015 ;
        RECT 65.405 205.215 65.655 206.345 ;
        RECT 65.870 206.015 66.275 206.345 ;
        RECT 66.445 205.845 66.615 206.515 ;
        RECT 65.845 205.675 66.615 205.845 ;
        RECT 66.785 206.515 67.145 206.890 ;
        RECT 67.410 206.515 67.580 207.255 ;
        RECT 67.860 206.685 68.030 206.890 ;
        RECT 67.860 206.515 68.400 206.685 ;
        RECT 66.785 205.860 67.040 206.515 ;
        RECT 67.210 206.015 67.560 206.345 ;
        RECT 67.730 206.015 68.060 206.345 ;
        RECT 65.845 205.045 66.095 205.675 ;
        RECT 64.665 204.875 66.095 205.045 ;
        RECT 66.275 204.705 66.605 205.505 ;
        RECT 66.785 204.875 67.125 205.860 ;
        RECT 67.295 205.475 67.560 206.015 ;
        RECT 68.230 205.815 68.400 206.515 ;
        RECT 67.775 205.645 68.400 205.815 ;
        RECT 68.570 205.885 68.740 207.085 ;
        RECT 68.970 206.605 69.300 207.085 ;
        RECT 69.470 206.785 69.640 207.255 ;
        RECT 69.810 206.605 70.140 207.070 ;
        RECT 68.970 206.435 70.140 206.605 ;
        RECT 70.470 206.580 70.745 206.925 ;
        RECT 70.935 206.855 71.315 207.255 ;
        RECT 71.485 206.685 71.655 207.035 ;
        RECT 71.825 206.855 72.155 207.255 ;
        RECT 72.325 206.685 72.580 207.035 ;
        RECT 68.910 206.055 69.480 206.265 ;
        RECT 69.650 206.055 70.295 206.265 ;
        RECT 68.570 205.475 69.275 205.885 ;
        RECT 70.470 205.845 70.640 206.580 ;
        RECT 70.915 206.515 72.580 206.685 ;
        RECT 72.765 206.605 73.025 207.085 ;
        RECT 73.195 206.715 73.445 207.255 ;
        RECT 70.915 206.345 71.085 206.515 ;
        RECT 70.810 206.015 71.085 206.345 ;
        RECT 71.255 206.015 72.080 206.345 ;
        RECT 72.250 206.015 72.595 206.345 ;
        RECT 70.915 205.845 71.085 206.015 ;
        RECT 67.295 205.305 69.275 205.475 ;
        RECT 67.295 204.705 67.705 205.135 ;
        RECT 68.450 204.705 68.780 205.125 ;
        RECT 68.950 204.875 69.275 205.305 ;
        RECT 69.750 204.705 70.080 205.805 ;
        RECT 70.470 204.875 70.745 205.845 ;
        RECT 70.915 205.675 71.575 205.845 ;
        RECT 71.885 205.725 72.080 206.015 ;
        RECT 71.405 205.555 71.575 205.675 ;
        RECT 72.250 205.555 72.575 205.845 ;
        RECT 70.955 204.705 71.235 205.505 ;
        RECT 71.405 205.385 72.575 205.555 ;
        RECT 72.765 205.575 72.935 206.605 ;
        RECT 73.615 206.550 73.835 207.035 ;
        RECT 73.105 205.955 73.335 206.350 ;
        RECT 73.505 206.125 73.835 206.550 ;
        RECT 74.005 206.875 74.895 207.045 ;
        RECT 74.005 206.150 74.175 206.875 ;
        RECT 74.345 206.320 74.895 206.705 ;
        RECT 74.005 206.080 74.895 206.150 ;
        RECT 74.000 206.055 74.895 206.080 ;
        RECT 73.990 206.040 74.895 206.055 ;
        RECT 73.985 206.025 74.895 206.040 ;
        RECT 73.975 206.020 74.895 206.025 ;
        RECT 73.970 206.010 74.895 206.020 ;
        RECT 73.965 206.000 74.895 206.010 ;
        RECT 73.955 205.995 74.895 206.000 ;
        RECT 73.945 205.985 74.895 205.995 ;
        RECT 73.935 205.980 74.895 205.985 ;
        RECT 73.935 205.975 74.270 205.980 ;
        RECT 73.920 205.970 74.270 205.975 ;
        RECT 73.905 205.960 74.270 205.970 ;
        RECT 73.880 205.955 74.270 205.960 ;
        RECT 73.105 205.950 74.270 205.955 ;
        RECT 73.105 205.915 74.240 205.950 ;
        RECT 73.105 205.890 74.205 205.915 ;
        RECT 73.105 205.860 74.175 205.890 ;
        RECT 73.105 205.830 74.155 205.860 ;
        RECT 73.105 205.800 74.135 205.830 ;
        RECT 73.105 205.790 74.065 205.800 ;
        RECT 73.105 205.780 74.040 205.790 ;
        RECT 73.105 205.765 74.020 205.780 ;
        RECT 73.105 205.750 74.000 205.765 ;
        RECT 73.210 205.740 73.995 205.750 ;
        RECT 73.210 205.705 73.980 205.740 ;
        RECT 71.405 204.925 72.595 205.215 ;
        RECT 72.765 204.875 73.040 205.575 ;
        RECT 73.210 205.455 73.965 205.705 ;
        RECT 74.135 205.385 74.465 205.630 ;
        RECT 74.635 205.530 74.895 205.980 ;
        RECT 74.280 205.360 74.465 205.385 ;
        RECT 74.280 205.260 74.895 205.360 ;
        RECT 73.210 204.705 73.465 205.250 ;
        RECT 73.635 204.875 74.115 205.215 ;
        RECT 74.290 204.705 74.895 205.260 ;
        RECT 75.065 204.875 75.345 206.975 ;
        RECT 75.575 206.795 75.745 207.255 ;
        RECT 76.015 206.865 77.265 207.045 ;
        RECT 76.400 206.625 76.765 206.695 ;
        RECT 75.515 206.445 76.765 206.625 ;
        RECT 76.935 206.645 77.265 206.865 ;
        RECT 77.435 206.815 77.605 207.255 ;
        RECT 77.775 206.645 78.115 207.060 ;
        RECT 76.935 206.475 78.115 206.645 ;
        RECT 78.285 206.605 78.545 207.085 ;
        RECT 78.715 206.715 78.965 207.255 ;
        RECT 75.515 205.845 75.790 206.445 ;
        RECT 75.960 206.015 76.315 206.265 ;
        RECT 76.510 206.235 76.975 206.265 ;
        RECT 76.505 206.065 76.975 206.235 ;
        RECT 76.510 206.015 76.975 206.065 ;
        RECT 77.145 206.015 77.475 206.265 ;
        RECT 77.650 206.065 78.115 206.265 ;
        RECT 77.295 205.895 77.475 206.015 ;
        RECT 75.515 205.635 77.125 205.845 ;
        RECT 77.295 205.725 77.625 205.895 ;
        RECT 76.715 205.535 77.125 205.635 ;
        RECT 75.535 204.705 76.320 205.465 ;
        RECT 76.715 204.875 77.100 205.535 ;
        RECT 77.425 204.935 77.625 205.725 ;
        RECT 77.795 204.705 78.115 205.885 ;
        RECT 78.285 205.575 78.455 206.605 ;
        RECT 79.135 206.575 79.355 207.035 ;
        RECT 79.105 206.550 79.355 206.575 ;
        RECT 78.625 205.955 78.855 206.350 ;
        RECT 79.025 206.125 79.355 206.550 ;
        RECT 79.525 206.875 80.415 207.045 ;
        RECT 79.525 206.150 79.695 206.875 ;
        RECT 79.865 206.320 80.415 206.705 ;
        RECT 80.645 206.435 80.855 207.255 ;
        RECT 81.025 206.455 81.355 207.085 ;
        RECT 79.525 206.080 80.415 206.150 ;
        RECT 79.520 206.055 80.415 206.080 ;
        RECT 79.510 206.040 80.415 206.055 ;
        RECT 79.505 206.025 80.415 206.040 ;
        RECT 79.495 206.020 80.415 206.025 ;
        RECT 79.490 206.010 80.415 206.020 ;
        RECT 79.485 206.000 80.415 206.010 ;
        RECT 79.475 205.995 80.415 206.000 ;
        RECT 79.465 205.985 80.415 205.995 ;
        RECT 79.455 205.980 80.415 205.985 ;
        RECT 79.455 205.975 79.790 205.980 ;
        RECT 79.440 205.970 79.790 205.975 ;
        RECT 79.425 205.960 79.790 205.970 ;
        RECT 79.400 205.955 79.790 205.960 ;
        RECT 78.625 205.950 79.790 205.955 ;
        RECT 78.625 205.915 79.760 205.950 ;
        RECT 78.625 205.890 79.725 205.915 ;
        RECT 78.625 205.860 79.695 205.890 ;
        RECT 78.625 205.830 79.675 205.860 ;
        RECT 78.625 205.800 79.655 205.830 ;
        RECT 78.625 205.790 79.585 205.800 ;
        RECT 78.625 205.780 79.560 205.790 ;
        RECT 78.625 205.765 79.540 205.780 ;
        RECT 78.625 205.750 79.520 205.765 ;
        RECT 78.730 205.740 79.515 205.750 ;
        RECT 78.730 205.705 79.500 205.740 ;
        RECT 78.285 204.875 78.560 205.575 ;
        RECT 78.730 205.455 79.485 205.705 ;
        RECT 79.655 205.385 79.985 205.630 ;
        RECT 80.155 205.530 80.415 205.980 ;
        RECT 81.025 205.855 81.275 206.455 ;
        RECT 81.525 206.435 81.755 207.255 ;
        RECT 81.445 206.015 81.775 206.265 ;
        RECT 79.800 205.360 79.985 205.385 ;
        RECT 79.800 205.260 80.415 205.360 ;
        RECT 78.730 204.705 78.985 205.250 ;
        RECT 79.155 204.875 79.635 205.215 ;
        RECT 79.810 204.705 80.415 205.260 ;
        RECT 80.645 204.705 80.855 205.845 ;
        RECT 81.025 204.875 81.355 205.855 ;
        RECT 81.525 204.705 81.755 205.845 ;
        RECT 81.975 204.885 82.235 207.075 ;
        RECT 82.495 206.885 83.165 207.255 ;
        RECT 83.345 206.705 83.655 207.075 ;
        RECT 82.425 206.505 83.655 206.705 ;
        RECT 82.425 205.835 82.715 206.505 ;
        RECT 83.835 206.325 84.065 206.965 ;
        RECT 84.245 206.525 84.535 207.255 ;
        RECT 82.895 206.015 83.360 206.325 ;
        RECT 83.540 206.015 84.065 206.325 ;
        RECT 84.245 206.015 84.545 206.345 ;
        RECT 82.425 205.615 83.195 205.835 ;
        RECT 82.405 204.705 82.745 205.435 ;
        RECT 82.925 204.885 83.195 205.615 ;
        RECT 83.375 205.595 84.535 205.835 ;
        RECT 83.375 204.885 83.605 205.595 ;
        RECT 83.775 204.705 84.105 205.415 ;
        RECT 84.275 204.885 84.535 205.595 ;
        RECT 84.725 204.875 85.005 206.975 ;
        RECT 85.235 206.795 85.405 207.255 ;
        RECT 85.675 206.865 86.925 207.045 ;
        RECT 86.060 206.625 86.425 206.695 ;
        RECT 85.175 206.445 86.425 206.625 ;
        RECT 86.595 206.645 86.925 206.865 ;
        RECT 87.095 206.815 87.265 207.255 ;
        RECT 87.435 206.645 87.775 207.060 ;
        RECT 86.595 206.475 87.775 206.645 ;
        RECT 87.945 206.530 88.235 207.255 ;
        RECT 85.175 205.845 85.450 206.445 ;
        RECT 85.620 206.015 85.975 206.265 ;
        RECT 86.170 206.235 86.635 206.265 ;
        RECT 86.165 206.065 86.635 206.235 ;
        RECT 86.170 206.015 86.635 206.065 ;
        RECT 86.805 206.015 87.135 206.265 ;
        RECT 87.310 206.065 87.775 206.265 ;
        RECT 86.955 205.895 87.135 206.015 ;
        RECT 85.175 205.635 86.785 205.845 ;
        RECT 86.955 205.725 87.285 205.895 ;
        RECT 86.375 205.535 86.785 205.635 ;
        RECT 85.195 204.705 85.980 205.465 ;
        RECT 86.375 204.875 86.760 205.535 ;
        RECT 87.085 204.935 87.285 205.725 ;
        RECT 87.455 204.705 87.775 205.885 ;
        RECT 87.945 204.705 88.235 205.870 ;
        RECT 88.405 204.875 88.685 206.975 ;
        RECT 88.915 206.795 89.085 207.255 ;
        RECT 89.355 206.865 90.605 207.045 ;
        RECT 89.740 206.625 90.105 206.695 ;
        RECT 88.855 206.445 90.105 206.625 ;
        RECT 90.275 206.645 90.605 206.865 ;
        RECT 90.775 206.815 90.945 207.255 ;
        RECT 91.115 206.645 91.455 207.060 ;
        RECT 90.275 206.475 91.455 206.645 ;
        RECT 88.855 205.845 89.130 206.445 ;
        RECT 89.300 206.015 89.655 206.265 ;
        RECT 89.850 206.235 90.315 206.265 ;
        RECT 89.845 206.065 90.315 206.235 ;
        RECT 89.850 206.015 90.315 206.065 ;
        RECT 90.485 206.015 90.815 206.265 ;
        RECT 90.990 206.065 91.455 206.265 ;
        RECT 90.635 205.895 90.815 206.015 ;
        RECT 88.855 205.635 90.465 205.845 ;
        RECT 90.635 205.725 90.965 205.895 ;
        RECT 90.055 205.535 90.465 205.635 ;
        RECT 88.875 204.705 89.660 205.465 ;
        RECT 90.055 204.875 90.440 205.535 ;
        RECT 90.765 204.935 90.965 205.725 ;
        RECT 91.135 204.705 91.455 205.885 ;
        RECT 92.555 204.885 92.815 207.075 ;
        RECT 93.075 206.885 93.745 207.255 ;
        RECT 93.925 206.705 94.235 207.075 ;
        RECT 93.005 206.505 94.235 206.705 ;
        RECT 93.005 205.835 93.295 206.505 ;
        RECT 94.415 206.325 94.645 206.965 ;
        RECT 94.825 206.525 95.115 207.255 ;
        RECT 95.330 206.865 95.660 207.255 ;
        RECT 95.830 206.695 96.055 207.075 ;
        RECT 93.475 206.015 93.940 206.325 ;
        RECT 94.120 206.015 94.645 206.325 ;
        RECT 94.825 206.015 95.125 206.345 ;
        RECT 95.315 206.015 95.555 206.665 ;
        RECT 95.725 206.515 96.055 206.695 ;
        RECT 95.725 205.845 95.900 206.515 ;
        RECT 96.255 206.345 96.485 206.965 ;
        RECT 96.665 206.525 96.965 207.255 ;
        RECT 97.150 206.710 102.495 207.255 ;
        RECT 102.670 206.710 108.015 207.255 ;
        RECT 108.190 206.710 113.535 207.255 ;
        RECT 96.070 206.015 96.485 206.345 ;
        RECT 96.665 206.015 96.960 206.345 ;
        RECT 93.005 205.615 93.775 205.835 ;
        RECT 92.985 204.705 93.325 205.435 ;
        RECT 93.505 204.885 93.775 205.615 ;
        RECT 93.955 205.595 95.115 205.835 ;
        RECT 93.955 204.885 94.185 205.595 ;
        RECT 94.355 204.705 94.685 205.415 ;
        RECT 94.855 204.885 95.115 205.595 ;
        RECT 95.315 205.655 95.900 205.845 ;
        RECT 95.315 204.885 95.590 205.655 ;
        RECT 96.070 205.485 96.965 205.815 ;
        RECT 95.760 205.315 96.965 205.485 ;
        RECT 95.760 204.885 96.090 205.315 ;
        RECT 96.260 204.705 96.455 205.145 ;
        RECT 96.635 204.885 96.965 205.315 ;
        RECT 98.740 205.140 99.090 206.390 ;
        RECT 100.570 205.880 100.910 206.710 ;
        RECT 104.260 205.140 104.610 206.390 ;
        RECT 106.090 205.880 106.430 206.710 ;
        RECT 109.780 205.140 110.130 206.390 ;
        RECT 111.610 205.880 111.950 206.710 ;
        RECT 113.705 206.530 113.995 207.255 ;
        RECT 114.630 206.710 119.975 207.255 ;
        RECT 120.150 206.710 125.495 207.255 ;
        RECT 97.150 204.705 102.495 205.140 ;
        RECT 102.670 204.705 108.015 205.140 ;
        RECT 108.190 204.705 113.535 205.140 ;
        RECT 113.705 204.705 113.995 205.870 ;
        RECT 116.220 205.140 116.570 206.390 ;
        RECT 118.050 205.880 118.390 206.710 ;
        RECT 121.740 205.140 122.090 206.390 ;
        RECT 123.570 205.880 123.910 206.710 ;
        RECT 125.665 206.505 126.875 207.255 ;
        RECT 125.665 205.795 126.185 206.335 ;
        RECT 126.355 205.965 126.875 206.505 ;
        RECT 114.630 204.705 119.975 205.140 ;
        RECT 120.150 204.705 125.495 205.140 ;
        RECT 125.665 204.705 126.875 205.795 ;
        RECT 14.260 204.535 126.960 204.705 ;
        RECT 14.345 203.445 15.555 204.535 ;
        RECT 14.345 202.735 14.865 203.275 ;
        RECT 15.035 202.905 15.555 203.445 ;
        RECT 15.785 203.395 15.995 204.535 ;
        RECT 16.165 203.385 16.495 204.365 ;
        RECT 16.665 203.395 16.895 204.535 ;
        RECT 17.180 203.920 17.510 204.295 ;
        RECT 17.735 204.175 18.065 204.535 ;
        RECT 18.235 203.920 18.405 204.365 ;
        RECT 18.575 204.175 18.905 204.535 ;
        RECT 19.075 204.195 20.085 204.365 ;
        RECT 19.075 203.920 19.255 204.195 ;
        RECT 17.180 203.750 19.255 203.920 ;
        RECT 14.345 201.985 15.555 202.735 ;
        RECT 15.785 201.985 15.995 202.805 ;
        RECT 16.165 202.785 16.415 203.385 ;
        RECT 17.180 203.360 17.435 203.750 ;
        RECT 17.605 203.410 18.895 203.580 ;
        RECT 16.585 202.975 16.915 203.225 ;
        RECT 17.605 203.190 17.855 203.410 ;
        RECT 17.440 202.955 17.855 203.190 ;
        RECT 18.720 203.175 18.895 203.410 ;
        RECT 19.075 203.345 19.255 203.750 ;
        RECT 18.025 202.910 18.550 203.175 ;
        RECT 18.720 203.005 19.175 203.175 ;
        RECT 18.720 202.910 19.115 203.005 ;
        RECT 16.165 202.155 16.495 202.785 ;
        RECT 16.665 201.985 16.895 202.805 ;
        RECT 17.315 201.985 17.595 202.785 ;
        RECT 19.495 202.740 19.665 204.025 ;
        RECT 19.915 203.595 20.085 204.195 ;
        RECT 19.835 202.895 20.145 203.425 ;
        RECT 20.375 203.415 20.625 204.535 ;
        RECT 20.805 203.655 21.055 204.085 ;
        RECT 21.235 203.835 21.565 204.535 ;
        RECT 21.745 203.655 21.915 204.085 ;
        RECT 22.095 203.835 22.425 204.535 ;
        RECT 20.805 203.485 22.395 203.655 ;
        RECT 20.335 202.895 21.740 203.225 ;
        RECT 18.175 202.685 19.665 202.740 ;
        RECT 20.335 202.685 20.505 202.895 ;
        RECT 21.910 202.685 22.395 203.485 ;
        RECT 23.545 203.370 23.835 204.535 ;
        RECT 24.100 203.345 24.270 204.535 ;
        RECT 24.440 203.685 24.700 204.365 ;
        RECT 24.870 203.775 25.200 204.535 ;
        RECT 25.370 203.935 25.620 204.365 ;
        RECT 25.790 204.115 26.145 204.535 ;
        RECT 26.335 204.195 27.505 204.365 ;
        RECT 26.335 204.155 26.665 204.195 ;
        RECT 26.775 203.935 27.005 204.025 ;
        RECT 25.370 203.695 27.005 203.935 ;
        RECT 18.175 202.570 20.505 202.685 ;
        RECT 18.175 202.305 18.455 202.570 ;
        RECT 19.495 202.515 20.505 202.570 ;
        RECT 20.805 202.515 22.395 202.685 ;
        RECT 18.955 201.985 19.285 202.345 ;
        RECT 19.495 202.155 19.665 202.515 ;
        RECT 19.855 201.985 20.630 202.345 ;
        RECT 21.235 201.985 21.565 202.345 ;
        RECT 22.095 201.985 22.435 202.345 ;
        RECT 23.545 201.985 23.835 202.710 ;
        RECT 24.100 201.985 24.270 202.885 ;
        RECT 24.440 202.485 24.610 203.685 ;
        RECT 27.175 203.525 27.505 204.195 ;
        RECT 27.775 203.865 27.945 204.365 ;
        RECT 28.155 204.075 28.405 204.535 ;
        RECT 28.775 203.865 28.945 204.365 ;
        RECT 29.155 204.075 29.405 204.535 ;
        RECT 29.615 203.865 29.785 204.365 ;
        RECT 27.775 203.695 29.785 203.865 ;
        RECT 29.955 203.565 30.285 204.325 ;
        RECT 30.475 203.735 30.725 204.535 ;
        RECT 24.785 203.355 27.505 203.525 ;
        RECT 24.785 202.805 24.955 203.355 ;
        RECT 25.185 202.975 25.590 203.175 ;
        RECT 25.760 202.975 26.090 203.185 ;
        RECT 24.785 202.635 25.625 202.805 ;
        RECT 24.440 202.155 24.700 202.485 ;
        RECT 24.915 201.985 25.245 202.465 ;
        RECT 25.455 202.405 25.625 202.635 ;
        RECT 25.880 202.575 26.090 202.975 ;
        RECT 26.360 202.975 26.835 203.185 ;
        RECT 27.025 202.975 27.510 203.175 ;
        RECT 26.360 202.575 26.580 202.975 ;
        RECT 25.455 202.155 26.780 202.405 ;
        RECT 27.055 201.985 27.505 202.750 ;
        RECT 27.735 202.630 27.955 203.525 ;
        RECT 28.190 203.145 28.405 203.525 ;
        RECT 28.650 203.335 29.055 203.525 ;
        RECT 28.190 202.975 28.655 203.145 ;
        RECT 28.190 202.645 28.405 202.975 ;
        RECT 28.885 202.895 29.055 203.335 ;
        RECT 29.405 203.175 29.740 203.525 ;
        RECT 29.955 203.395 30.760 203.565 ;
        RECT 29.405 203.005 29.755 203.175 ;
        RECT 29.405 202.895 29.740 203.005 ;
        RECT 30.010 202.975 30.340 203.195 ;
        RECT 30.590 202.705 30.760 203.395 ;
        RECT 29.195 202.535 30.760 202.705 ;
        RECT 30.955 202.655 31.145 204.365 ;
        RECT 31.315 203.395 31.645 204.535 ;
        RECT 31.915 203.790 32.185 204.535 ;
        RECT 32.815 204.530 39.090 204.535 ;
        RECT 32.355 203.620 32.645 204.360 ;
        RECT 32.815 203.805 33.070 204.530 ;
        RECT 33.255 203.635 33.515 204.360 ;
        RECT 33.685 203.805 33.930 204.530 ;
        RECT 34.115 203.635 34.375 204.360 ;
        RECT 34.545 203.805 34.790 204.530 ;
        RECT 34.975 203.635 35.235 204.360 ;
        RECT 35.405 203.805 35.650 204.530 ;
        RECT 35.820 203.635 36.080 204.360 ;
        RECT 36.250 203.805 36.510 204.530 ;
        RECT 36.680 203.635 36.940 204.360 ;
        RECT 37.110 203.805 37.370 204.530 ;
        RECT 37.540 203.635 37.800 204.360 ;
        RECT 37.970 203.805 38.230 204.530 ;
        RECT 38.400 203.635 38.660 204.360 ;
        RECT 38.830 203.735 39.090 204.530 ;
        RECT 33.255 203.620 38.660 203.635 ;
        RECT 31.915 203.395 38.660 203.620 ;
        RECT 31.915 202.805 33.080 203.395 ;
        RECT 39.260 203.225 39.510 204.360 ;
        RECT 39.690 203.725 39.950 204.535 ;
        RECT 40.125 203.225 40.370 204.365 ;
        RECT 40.550 203.725 40.845 204.535 ;
        RECT 41.025 203.395 41.355 204.535 ;
        RECT 41.525 203.905 41.880 204.365 ;
        RECT 42.050 204.075 42.625 204.535 ;
        RECT 42.795 203.905 43.125 204.365 ;
        RECT 41.525 203.735 43.125 203.905 ;
        RECT 43.325 203.735 43.580 204.535 ;
        RECT 41.525 203.395 41.800 203.735 ;
        RECT 41.980 203.515 42.170 203.555 ;
        RECT 41.545 203.345 41.715 203.395 ;
        RECT 41.980 203.345 42.175 203.515 ;
        RECT 33.250 202.975 40.370 203.225 ;
        RECT 29.195 202.365 29.365 202.535 ;
        RECT 27.695 202.195 29.365 202.365 ;
        RECT 29.535 201.985 29.865 202.365 ;
        RECT 30.035 202.155 30.245 202.535 ;
        RECT 30.475 201.985 30.805 202.365 ;
        RECT 30.975 202.195 31.145 202.655 ;
        RECT 31.315 201.985 31.645 202.705 ;
        RECT 31.915 202.635 38.660 202.805 ;
        RECT 31.915 201.985 32.215 202.465 ;
        RECT 32.385 202.180 32.645 202.635 ;
        RECT 32.815 201.985 33.075 202.465 ;
        RECT 33.255 202.180 33.515 202.635 ;
        RECT 33.685 201.985 33.935 202.465 ;
        RECT 34.115 202.180 34.375 202.635 ;
        RECT 34.545 201.985 34.795 202.465 ;
        RECT 34.975 202.180 35.235 202.635 ;
        RECT 35.405 201.985 35.650 202.465 ;
        RECT 35.820 202.180 36.095 202.635 ;
        RECT 36.265 201.985 36.510 202.465 ;
        RECT 36.680 202.180 36.940 202.635 ;
        RECT 37.110 201.985 37.370 202.465 ;
        RECT 37.540 202.180 37.800 202.635 ;
        RECT 37.970 201.985 38.230 202.465 ;
        RECT 38.400 202.180 38.660 202.635 ;
        RECT 38.830 201.985 39.090 202.545 ;
        RECT 39.260 202.165 39.510 202.975 ;
        RECT 39.690 201.985 39.950 202.510 ;
        RECT 40.120 202.165 40.370 202.975 ;
        RECT 40.540 202.665 40.855 203.225 ;
        RECT 41.980 203.175 42.170 203.345 ;
        RECT 41.025 202.975 42.170 203.175 ;
        RECT 42.350 202.805 42.630 203.735 ;
        RECT 43.750 203.565 44.050 203.760 ;
        RECT 42.800 203.395 44.050 203.565 ;
        RECT 44.370 203.395 44.700 204.535 ;
        RECT 44.900 203.565 45.230 204.365 ;
        RECT 45.400 203.735 45.570 204.535 ;
        RECT 45.740 203.565 46.070 204.365 ;
        RECT 46.240 203.735 46.410 204.535 ;
        RECT 46.580 203.565 46.925 204.365 ;
        RECT 47.095 203.735 47.265 204.535 ;
        RECT 47.435 203.565 47.765 204.365 ;
        RECT 42.800 202.975 43.130 203.395 ;
        RECT 43.360 202.895 43.705 203.225 ;
        RECT 41.025 202.595 42.135 202.805 ;
        RECT 40.550 201.985 40.855 202.495 ;
        RECT 41.025 202.155 41.375 202.595 ;
        RECT 41.545 201.985 41.715 202.425 ;
        RECT 41.885 202.365 42.135 202.595 ;
        RECT 42.305 202.705 42.630 202.805 ;
        RECT 42.305 202.535 42.635 202.705 ;
        RECT 42.805 202.365 43.080 202.805 ;
        RECT 43.880 202.740 44.050 203.395 ;
        RECT 44.900 203.345 47.765 203.565 ;
        RECT 47.935 203.735 48.625 204.535 ;
        RECT 47.935 203.345 48.250 203.735 ;
        RECT 48.795 203.565 49.130 204.365 ;
        RECT 48.440 203.345 49.130 203.565 ;
        RECT 49.305 203.370 49.595 204.535 ;
        RECT 49.765 203.395 50.125 204.535 ;
        RECT 50.795 203.855 51.125 204.365 ;
        RECT 52.295 204.025 52.805 204.535 ;
        RECT 50.295 203.685 52.805 203.855 ;
        RECT 44.280 202.975 46.065 203.175 ;
        RECT 46.580 202.805 46.845 203.345 ;
        RECT 48.440 203.175 48.610 203.345 ;
        RECT 47.015 202.975 48.610 203.175 ;
        RECT 48.780 202.975 49.110 203.175 ;
        RECT 49.765 203.145 50.095 203.225 ;
        RECT 49.765 202.975 50.125 203.145 ;
        RECT 48.440 202.805 48.610 202.975 ;
        RECT 41.885 202.155 43.080 202.365 ;
        RECT 43.315 201.985 43.645 202.725 ;
        RECT 43.815 202.410 44.050 202.740 ;
        RECT 44.370 202.615 46.410 202.805 ;
        RECT 44.370 202.155 44.700 202.615 ;
        RECT 44.910 201.985 45.150 202.445 ;
        RECT 45.320 202.155 45.650 202.615 ;
        RECT 45.820 201.985 45.990 202.445 ;
        RECT 46.160 202.365 46.410 202.615 ;
        RECT 46.580 202.535 47.765 202.805 ;
        RECT 47.935 202.365 48.185 202.805 ;
        RECT 48.440 202.615 49.130 202.805 ;
        RECT 46.160 202.155 48.185 202.365 ;
        RECT 48.430 201.985 48.625 202.445 ;
        RECT 48.795 202.155 49.130 202.615 ;
        RECT 49.305 201.985 49.595 202.710 ;
        RECT 49.765 202.325 50.125 202.805 ;
        RECT 50.295 202.725 50.495 203.685 ;
        RECT 50.665 203.345 50.915 203.515 ;
        RECT 50.665 202.895 50.910 203.345 ;
        RECT 51.185 202.895 51.405 203.515 ;
        RECT 51.660 202.895 51.835 203.515 ;
        RECT 52.105 202.895 52.325 203.515 ;
        RECT 52.495 202.895 52.805 203.685 ;
        RECT 50.295 202.495 50.625 202.725 ;
        RECT 50.795 202.555 52.125 202.725 ;
        RECT 50.795 202.325 51.125 202.555 ;
        RECT 49.765 202.155 51.125 202.325 ;
        RECT 51.295 201.985 51.625 202.385 ;
        RECT 51.795 202.155 52.125 202.555 ;
        RECT 52.395 201.985 52.725 202.725 ;
        RECT 52.975 202.155 53.305 204.365 ;
        RECT 53.475 203.395 53.735 204.535 ;
        RECT 53.995 203.915 54.165 204.345 ;
        RECT 54.335 204.085 54.665 204.535 ;
        RECT 53.995 203.685 54.670 203.915 ;
        RECT 53.475 201.985 53.735 202.785 ;
        RECT 53.965 202.665 54.265 203.515 ;
        RECT 54.435 203.035 54.670 203.685 ;
        RECT 54.840 203.375 55.125 204.320 ;
        RECT 55.305 204.065 55.990 204.535 ;
        RECT 55.300 203.545 55.995 203.855 ;
        RECT 56.170 203.480 56.475 204.265 ;
        RECT 54.840 203.225 55.700 203.375 ;
        RECT 54.840 203.205 56.125 203.225 ;
        RECT 54.435 202.705 54.970 203.035 ;
        RECT 55.140 202.845 56.125 203.205 ;
        RECT 54.435 202.555 54.655 202.705 ;
        RECT 53.910 201.985 54.245 202.490 ;
        RECT 54.415 202.180 54.655 202.555 ;
        RECT 55.140 202.510 55.310 202.845 ;
        RECT 56.300 202.675 56.475 203.480 ;
        RECT 56.665 203.395 56.995 204.535 ;
        RECT 57.165 203.905 57.520 204.365 ;
        RECT 57.690 204.075 58.265 204.535 ;
        RECT 58.435 203.905 58.765 204.365 ;
        RECT 57.165 203.735 58.765 203.905 ;
        RECT 58.965 203.735 59.220 204.535 ;
        RECT 57.165 203.395 57.440 203.735 ;
        RECT 57.620 203.515 57.810 203.555 ;
        RECT 57.620 203.345 57.815 203.515 ;
        RECT 57.620 203.175 57.810 203.345 ;
        RECT 56.665 202.975 57.810 203.175 ;
        RECT 57.990 202.835 58.270 203.735 ;
        RECT 59.390 203.565 59.690 203.760 ;
        RECT 58.440 203.395 59.690 203.565 ;
        RECT 58.440 202.975 58.770 203.395 ;
        RECT 59.000 202.895 59.345 203.225 ;
        RECT 57.990 202.805 58.275 202.835 ;
        RECT 54.935 202.315 55.310 202.510 ;
        RECT 54.935 202.170 55.105 202.315 ;
        RECT 55.670 201.985 56.065 202.480 ;
        RECT 56.235 202.155 56.475 202.675 ;
        RECT 56.665 202.595 57.775 202.805 ;
        RECT 56.665 202.155 57.015 202.595 ;
        RECT 57.185 201.985 57.355 202.425 ;
        RECT 57.525 202.365 57.775 202.595 ;
        RECT 57.945 202.535 58.275 202.805 ;
        RECT 58.445 202.365 58.720 202.805 ;
        RECT 59.520 202.740 59.690 203.395 ;
        RECT 57.525 202.155 58.720 202.365 ;
        RECT 58.955 201.985 59.285 202.725 ;
        RECT 59.455 202.410 59.690 202.740 ;
        RECT 59.905 203.480 60.210 204.265 ;
        RECT 60.390 204.065 61.075 204.535 ;
        RECT 60.385 203.545 61.080 203.855 ;
        RECT 59.905 202.675 60.080 203.480 ;
        RECT 61.255 203.375 61.540 204.320 ;
        RECT 61.715 204.085 62.045 204.535 ;
        RECT 62.215 203.915 62.385 204.345 ;
        RECT 60.680 203.225 61.540 203.375 ;
        RECT 60.255 203.205 61.540 203.225 ;
        RECT 61.710 203.685 62.385 203.915 ;
        RECT 60.255 202.845 61.240 203.205 ;
        RECT 61.710 203.035 61.945 203.685 ;
        RECT 59.905 202.155 60.145 202.675 ;
        RECT 61.070 202.510 61.240 202.845 ;
        RECT 61.410 202.705 61.945 203.035 ;
        RECT 61.725 202.555 61.945 202.705 ;
        RECT 62.115 202.665 62.415 203.515 ;
        RECT 62.645 203.445 63.855 204.535 ;
        RECT 64.065 203.585 64.355 204.355 ;
        RECT 64.925 203.995 65.185 204.355 ;
        RECT 65.355 204.165 65.685 204.535 ;
        RECT 65.855 203.995 66.115 204.355 ;
        RECT 64.925 203.765 66.115 203.995 ;
        RECT 66.305 203.815 66.635 204.535 ;
        RECT 66.805 203.585 67.070 204.355 ;
        RECT 62.645 202.905 63.165 203.445 ;
        RECT 64.065 203.405 66.560 203.585 ;
        RECT 63.335 202.735 63.855 203.275 ;
        RECT 64.035 202.895 64.305 203.225 ;
        RECT 64.485 202.895 64.920 203.225 ;
        RECT 65.100 202.895 65.675 203.225 ;
        RECT 65.855 202.895 66.135 203.225 ;
        RECT 60.315 201.985 60.710 202.480 ;
        RECT 61.070 202.315 61.445 202.510 ;
        RECT 61.275 202.170 61.445 202.315 ;
        RECT 61.725 202.180 61.965 202.555 ;
        RECT 62.135 201.985 62.470 202.490 ;
        RECT 62.645 201.985 63.855 202.735 ;
        RECT 66.335 202.715 66.560 203.405 ;
        RECT 64.075 202.525 66.560 202.715 ;
        RECT 64.075 202.165 64.300 202.525 ;
        RECT 64.480 201.985 64.810 202.355 ;
        RECT 64.990 202.165 65.245 202.525 ;
        RECT 65.810 201.985 66.555 202.355 ;
        RECT 66.735 202.165 67.070 203.585 ;
        RECT 67.255 203.585 67.530 204.355 ;
        RECT 67.700 203.925 68.030 204.355 ;
        RECT 68.200 204.095 68.395 204.535 ;
        RECT 68.575 203.925 68.905 204.355 ;
        RECT 67.700 203.755 68.905 203.925 ;
        RECT 67.255 203.395 67.840 203.585 ;
        RECT 68.010 203.425 68.905 203.755 ;
        RECT 69.085 203.445 70.295 204.535 ;
        RECT 70.465 203.665 70.740 204.365 ;
        RECT 70.910 203.990 71.165 204.535 ;
        RECT 71.335 204.025 71.815 204.365 ;
        RECT 71.990 203.980 72.595 204.535 ;
        RECT 71.980 203.880 72.595 203.980 ;
        RECT 71.980 203.855 72.165 203.880 ;
        RECT 67.255 202.575 67.495 203.225 ;
        RECT 67.665 202.725 67.840 203.395 ;
        RECT 68.010 202.895 68.425 203.225 ;
        RECT 68.605 202.895 68.900 203.225 ;
        RECT 69.085 202.905 69.605 203.445 ;
        RECT 67.665 202.545 67.995 202.725 ;
        RECT 67.270 201.985 67.600 202.375 ;
        RECT 67.770 202.165 67.995 202.545 ;
        RECT 68.195 202.275 68.425 202.895 ;
        RECT 69.775 202.735 70.295 203.275 ;
        RECT 68.605 201.985 68.905 202.715 ;
        RECT 69.085 201.985 70.295 202.735 ;
        RECT 70.465 202.635 70.635 203.665 ;
        RECT 70.910 203.535 71.665 203.785 ;
        RECT 71.835 203.610 72.165 203.855 ;
        RECT 70.910 203.500 71.680 203.535 ;
        RECT 70.910 203.490 71.695 203.500 ;
        RECT 70.805 203.475 71.700 203.490 ;
        RECT 70.805 203.460 71.720 203.475 ;
        RECT 70.805 203.450 71.740 203.460 ;
        RECT 70.805 203.440 71.765 203.450 ;
        RECT 70.805 203.410 71.835 203.440 ;
        RECT 70.805 203.380 71.855 203.410 ;
        RECT 70.805 203.350 71.875 203.380 ;
        RECT 70.805 203.325 71.905 203.350 ;
        RECT 70.805 203.290 71.940 203.325 ;
        RECT 70.805 203.285 71.970 203.290 ;
        RECT 70.805 202.890 71.035 203.285 ;
        RECT 71.580 203.280 71.970 203.285 ;
        RECT 71.605 203.270 71.970 203.280 ;
        RECT 71.620 203.265 71.970 203.270 ;
        RECT 71.635 203.260 71.970 203.265 ;
        RECT 72.335 203.260 72.595 203.710 ;
        RECT 71.635 203.255 72.595 203.260 ;
        RECT 71.645 203.245 72.595 203.255 ;
        RECT 71.655 203.240 72.595 203.245 ;
        RECT 71.665 203.230 72.595 203.240 ;
        RECT 71.670 203.220 72.595 203.230 ;
        RECT 71.675 203.215 72.595 203.220 ;
        RECT 71.685 203.200 72.595 203.215 ;
        RECT 71.690 203.185 72.595 203.200 ;
        RECT 71.700 203.160 72.595 203.185 ;
        RECT 71.205 202.690 71.535 203.115 ;
        RECT 70.465 202.155 70.725 202.635 ;
        RECT 70.895 201.985 71.145 202.525 ;
        RECT 71.315 202.205 71.535 202.690 ;
        RECT 71.705 203.090 72.595 203.160 ;
        RECT 72.765 203.665 73.040 204.365 ;
        RECT 73.210 203.990 73.465 204.535 ;
        RECT 73.635 204.025 74.115 204.365 ;
        RECT 74.290 203.980 74.895 204.535 ;
        RECT 74.280 203.880 74.895 203.980 ;
        RECT 74.280 203.855 74.465 203.880 ;
        RECT 71.705 202.365 71.875 203.090 ;
        RECT 72.045 202.535 72.595 202.920 ;
        RECT 72.765 202.635 72.935 203.665 ;
        RECT 73.210 203.535 73.965 203.785 ;
        RECT 74.135 203.610 74.465 203.855 ;
        RECT 73.210 203.500 73.980 203.535 ;
        RECT 73.210 203.490 73.995 203.500 ;
        RECT 73.105 203.475 74.000 203.490 ;
        RECT 73.105 203.460 74.020 203.475 ;
        RECT 73.105 203.450 74.040 203.460 ;
        RECT 73.105 203.440 74.065 203.450 ;
        RECT 73.105 203.410 74.135 203.440 ;
        RECT 73.105 203.380 74.155 203.410 ;
        RECT 73.105 203.350 74.175 203.380 ;
        RECT 73.105 203.325 74.205 203.350 ;
        RECT 73.105 203.290 74.240 203.325 ;
        RECT 73.105 203.285 74.270 203.290 ;
        RECT 73.105 202.890 73.335 203.285 ;
        RECT 73.880 203.280 74.270 203.285 ;
        RECT 73.905 203.270 74.270 203.280 ;
        RECT 73.920 203.265 74.270 203.270 ;
        RECT 73.935 203.260 74.270 203.265 ;
        RECT 74.635 203.260 74.895 203.710 ;
        RECT 75.065 203.370 75.355 204.535 ;
        RECT 75.525 203.395 75.795 204.365 ;
        RECT 76.005 203.735 76.285 204.535 ;
        RECT 76.455 204.025 78.110 204.315 ;
        RECT 78.290 204.100 83.635 204.535 ;
        RECT 76.520 203.685 78.110 203.855 ;
        RECT 76.520 203.565 76.690 203.685 ;
        RECT 75.965 203.395 76.690 203.565 ;
        RECT 73.935 203.255 74.895 203.260 ;
        RECT 73.945 203.245 74.895 203.255 ;
        RECT 73.955 203.240 74.895 203.245 ;
        RECT 73.965 203.230 74.895 203.240 ;
        RECT 73.970 203.220 74.895 203.230 ;
        RECT 73.975 203.215 74.895 203.220 ;
        RECT 73.985 203.200 74.895 203.215 ;
        RECT 73.990 203.185 74.895 203.200 ;
        RECT 74.000 203.160 74.895 203.185 ;
        RECT 73.505 202.690 73.835 203.115 ;
        RECT 71.705 202.195 72.595 202.365 ;
        RECT 72.765 202.155 73.025 202.635 ;
        RECT 73.195 201.985 73.445 202.525 ;
        RECT 73.615 202.205 73.835 202.690 ;
        RECT 74.005 203.090 74.895 203.160 ;
        RECT 74.005 202.365 74.175 203.090 ;
        RECT 74.345 202.535 74.895 202.920 ;
        RECT 74.005 202.195 74.895 202.365 ;
        RECT 75.065 201.985 75.355 202.710 ;
        RECT 75.525 202.660 75.695 203.395 ;
        RECT 75.965 203.225 76.135 203.395 ;
        RECT 75.865 202.895 76.135 203.225 ;
        RECT 76.305 202.895 76.710 203.225 ;
        RECT 76.880 202.895 77.590 203.515 ;
        RECT 77.790 203.395 78.110 203.685 ;
        RECT 75.965 202.725 76.135 202.895 ;
        RECT 75.525 202.315 75.795 202.660 ;
        RECT 75.965 202.555 77.575 202.725 ;
        RECT 77.760 202.655 78.110 203.225 ;
        RECT 79.880 202.850 80.230 204.100 ;
        RECT 83.805 203.395 84.065 204.535 ;
        RECT 84.235 203.385 84.565 204.365 ;
        RECT 84.735 203.395 85.015 204.535 ;
        RECT 85.195 203.925 85.525 204.355 ;
        RECT 85.705 204.095 85.900 204.535 ;
        RECT 86.070 203.925 86.400 204.355 ;
        RECT 85.195 203.755 86.400 203.925 ;
        RECT 85.195 203.425 86.090 203.755 ;
        RECT 86.570 203.585 86.845 204.355 ;
        RECT 86.260 203.395 86.845 203.585 ;
        RECT 87.210 203.565 87.600 203.740 ;
        RECT 88.085 203.735 88.415 204.535 ;
        RECT 88.585 203.745 89.120 204.365 ;
        RECT 87.210 203.395 88.635 203.565 ;
        RECT 75.985 201.985 76.365 202.385 ;
        RECT 76.535 202.205 76.705 202.555 ;
        RECT 76.875 201.985 77.205 202.385 ;
        RECT 77.405 202.205 77.575 202.555 ;
        RECT 81.710 202.530 82.050 203.360 ;
        RECT 83.825 202.975 84.160 203.225 ;
        RECT 84.330 202.835 84.500 203.385 ;
        RECT 84.670 202.955 85.005 203.225 ;
        RECT 85.200 202.895 85.495 203.225 ;
        RECT 85.675 202.895 86.090 203.225 ;
        RECT 84.325 202.785 84.500 202.835 ;
        RECT 77.775 201.985 78.105 202.485 ;
        RECT 78.290 201.985 83.635 202.530 ;
        RECT 83.805 202.155 84.500 202.785 ;
        RECT 84.705 201.985 85.015 202.785 ;
        RECT 85.195 201.985 85.495 202.715 ;
        RECT 85.675 202.275 85.905 202.895 ;
        RECT 86.260 202.725 86.435 203.395 ;
        RECT 86.105 202.545 86.435 202.725 ;
        RECT 86.605 202.575 86.845 203.225 ;
        RECT 87.085 202.665 87.440 203.225 ;
        RECT 86.105 202.165 86.330 202.545 ;
        RECT 87.610 202.495 87.780 203.395 ;
        RECT 87.950 202.665 88.215 203.225 ;
        RECT 88.465 202.895 88.635 203.395 ;
        RECT 88.805 202.725 89.120 203.745 ;
        RECT 89.415 203.565 89.585 204.365 ;
        RECT 90.345 203.905 90.595 204.365 ;
        RECT 90.795 204.155 91.465 204.535 ;
        RECT 91.655 203.905 91.905 204.365 ;
        RECT 92.080 204.075 92.325 204.535 ;
        RECT 90.345 203.735 91.905 203.905 ;
        RECT 92.495 203.685 92.835 204.325 ;
        RECT 89.415 203.395 92.355 203.565 ;
        RECT 92.185 203.225 92.355 203.395 ;
        RECT 89.385 202.895 89.570 203.225 ;
        RECT 89.825 202.895 90.300 203.225 ;
        RECT 90.610 202.895 90.955 203.225 ;
        RECT 86.500 201.985 86.830 202.375 ;
        RECT 87.190 201.985 87.430 202.495 ;
        RECT 87.610 202.165 87.890 202.495 ;
        RECT 88.120 201.985 88.335 202.495 ;
        RECT 88.505 202.155 89.120 202.725 ;
        RECT 89.415 202.555 90.595 202.725 ;
        RECT 90.765 202.665 90.955 202.895 ;
        RECT 91.215 202.650 91.410 203.225 ;
        RECT 91.680 202.895 92.015 203.225 ;
        RECT 92.185 202.895 92.495 203.225 ;
        RECT 92.185 202.725 92.355 202.895 ;
        RECT 89.415 202.155 89.585 202.555 ;
        RECT 89.825 201.985 90.155 202.385 ;
        RECT 90.425 202.325 90.595 202.555 ;
        RECT 91.660 202.555 92.355 202.725 ;
        RECT 92.665 202.570 92.835 203.685 ;
        RECT 93.465 203.395 93.745 204.535 ;
        RECT 93.915 203.385 94.245 204.365 ;
        RECT 94.415 203.395 94.675 204.535 ;
        RECT 95.310 204.100 100.655 204.535 ;
        RECT 93.980 203.345 94.155 203.385 ;
        RECT 93.475 202.955 93.810 203.225 ;
        RECT 93.980 202.785 94.150 203.345 ;
        RECT 94.320 202.975 94.655 203.225 ;
        RECT 96.900 202.850 97.250 204.100 ;
        RECT 100.825 203.370 101.115 204.535 ;
        RECT 101.745 203.445 103.415 204.535 ;
        RECT 103.585 203.565 103.855 204.335 ;
        RECT 104.025 203.755 104.355 204.535 ;
        RECT 104.560 203.930 104.745 204.335 ;
        RECT 104.915 204.110 105.250 204.535 ;
        RECT 104.560 203.755 105.225 203.930 ;
        RECT 105.625 203.865 105.905 204.535 ;
        RECT 91.660 202.325 91.830 202.555 ;
        RECT 90.425 202.155 91.830 202.325 ;
        RECT 92.000 201.985 92.330 202.365 ;
        RECT 92.525 202.155 92.835 202.570 ;
        RECT 93.465 201.985 93.775 202.785 ;
        RECT 93.980 202.155 94.675 202.785 ;
        RECT 98.730 202.530 99.070 203.360 ;
        RECT 101.745 202.925 102.495 203.445 ;
        RECT 103.585 203.395 104.715 203.565 ;
        RECT 102.665 202.755 103.415 203.275 ;
        RECT 95.310 201.985 100.655 202.530 ;
        RECT 100.825 201.985 101.115 202.710 ;
        RECT 101.745 201.985 103.415 202.755 ;
        RECT 103.585 202.485 103.755 203.395 ;
        RECT 103.925 202.645 104.285 203.225 ;
        RECT 104.465 202.895 104.715 203.395 ;
        RECT 104.885 202.725 105.225 203.755 ;
        RECT 106.075 203.645 106.375 204.195 ;
        RECT 106.575 203.815 106.905 204.535 ;
        RECT 107.095 203.815 107.555 204.365 ;
        RECT 105.440 203.225 105.705 203.585 ;
        RECT 106.075 203.475 107.015 203.645 ;
        RECT 106.845 203.225 107.015 203.475 ;
        RECT 105.440 202.975 106.115 203.225 ;
        RECT 106.335 202.975 106.675 203.225 ;
        RECT 106.845 202.895 107.135 203.225 ;
        RECT 106.845 202.805 107.015 202.895 ;
        RECT 104.540 202.555 105.225 202.725 ;
        RECT 105.625 202.615 107.015 202.805 ;
        RECT 103.585 202.155 103.845 202.485 ;
        RECT 104.055 201.985 104.330 202.465 ;
        RECT 104.540 202.155 104.745 202.555 ;
        RECT 104.915 201.985 105.250 202.385 ;
        RECT 105.625 202.255 105.955 202.615 ;
        RECT 107.305 202.445 107.555 203.815 ;
        RECT 107.725 203.445 110.315 204.535 ;
        RECT 110.485 203.565 110.755 204.335 ;
        RECT 110.925 203.755 111.255 204.535 ;
        RECT 111.460 203.930 111.645 204.335 ;
        RECT 111.815 204.110 112.150 204.535 ;
        RECT 111.460 203.755 112.125 203.930 ;
        RECT 107.725 202.925 108.935 203.445 ;
        RECT 110.485 203.395 111.615 203.565 ;
        RECT 109.105 202.755 110.315 203.275 ;
        RECT 106.575 201.985 106.825 202.445 ;
        RECT 106.995 202.155 107.555 202.445 ;
        RECT 107.725 201.985 110.315 202.755 ;
        RECT 110.485 202.485 110.655 203.395 ;
        RECT 110.825 202.645 111.185 203.225 ;
        RECT 111.365 202.895 111.615 203.395 ;
        RECT 111.785 202.725 112.125 203.755 ;
        RECT 112.785 203.445 114.455 204.535 ;
        RECT 114.630 204.100 119.975 204.535 ;
        RECT 120.150 204.100 125.495 204.535 ;
        RECT 112.785 202.925 113.535 203.445 ;
        RECT 113.705 202.755 114.455 203.275 ;
        RECT 116.220 202.850 116.570 204.100 ;
        RECT 111.440 202.555 112.125 202.725 ;
        RECT 110.485 202.155 110.745 202.485 ;
        RECT 110.955 201.985 111.230 202.465 ;
        RECT 111.440 202.155 111.645 202.555 ;
        RECT 111.815 201.985 112.150 202.385 ;
        RECT 112.785 201.985 114.455 202.755 ;
        RECT 118.050 202.530 118.390 203.360 ;
        RECT 121.740 202.850 122.090 204.100 ;
        RECT 125.665 203.445 126.875 204.535 ;
        RECT 123.570 202.530 123.910 203.360 ;
        RECT 125.665 202.905 126.185 203.445 ;
        RECT 126.355 202.735 126.875 203.275 ;
        RECT 114.630 201.985 119.975 202.530 ;
        RECT 120.150 201.985 125.495 202.530 ;
        RECT 125.665 201.985 126.875 202.735 ;
        RECT 14.260 201.815 126.960 201.985 ;
        RECT 14.345 201.065 15.555 201.815 ;
        RECT 14.345 200.525 14.865 201.065 ;
        RECT 15.730 200.975 15.990 201.815 ;
        RECT 16.165 201.070 16.420 201.645 ;
        RECT 16.590 201.435 16.920 201.815 ;
        RECT 17.135 201.265 17.305 201.645 ;
        RECT 18.025 201.305 18.330 201.815 ;
        RECT 16.590 201.095 17.305 201.265 ;
        RECT 15.035 200.355 15.555 200.895 ;
        RECT 14.345 199.265 15.555 200.355 ;
        RECT 15.730 199.265 15.990 200.415 ;
        RECT 16.165 200.340 16.335 201.070 ;
        RECT 16.590 200.905 16.760 201.095 ;
        RECT 16.505 200.575 16.760 200.905 ;
        RECT 16.590 200.365 16.760 200.575 ;
        RECT 17.040 200.545 17.395 200.915 ;
        RECT 18.025 200.575 18.340 201.135 ;
        RECT 18.510 200.825 18.760 201.635 ;
        RECT 18.930 201.290 19.190 201.815 ;
        RECT 19.370 200.825 19.620 201.635 ;
        RECT 19.790 201.255 20.050 201.815 ;
        RECT 20.220 201.165 20.480 201.620 ;
        RECT 20.650 201.335 20.910 201.815 ;
        RECT 21.080 201.165 21.340 201.620 ;
        RECT 21.510 201.335 21.770 201.815 ;
        RECT 21.940 201.165 22.200 201.620 ;
        RECT 22.370 201.335 22.615 201.815 ;
        RECT 22.785 201.165 23.060 201.620 ;
        RECT 23.230 201.335 23.475 201.815 ;
        RECT 23.645 201.165 23.905 201.620 ;
        RECT 24.085 201.335 24.335 201.815 ;
        RECT 24.505 201.165 24.765 201.620 ;
        RECT 24.945 201.335 25.195 201.815 ;
        RECT 25.365 201.165 25.625 201.620 ;
        RECT 25.805 201.335 26.065 201.815 ;
        RECT 26.235 201.165 26.495 201.620 ;
        RECT 26.665 201.335 26.965 201.815 ;
        RECT 27.315 201.335 27.615 201.815 ;
        RECT 27.785 201.165 28.045 201.620 ;
        RECT 28.215 201.335 28.475 201.815 ;
        RECT 28.655 201.165 28.915 201.620 ;
        RECT 29.085 201.335 29.335 201.815 ;
        RECT 29.515 201.165 29.775 201.620 ;
        RECT 29.945 201.335 30.195 201.815 ;
        RECT 30.375 201.165 30.635 201.620 ;
        RECT 30.805 201.335 31.050 201.815 ;
        RECT 31.220 201.165 31.495 201.620 ;
        RECT 31.665 201.335 31.910 201.815 ;
        RECT 32.080 201.165 32.340 201.620 ;
        RECT 32.510 201.335 32.770 201.815 ;
        RECT 32.940 201.165 33.200 201.620 ;
        RECT 33.370 201.335 33.630 201.815 ;
        RECT 33.800 201.165 34.060 201.620 ;
        RECT 34.230 201.255 34.490 201.815 ;
        RECT 20.220 200.995 26.965 201.165 ;
        RECT 18.510 200.575 25.630 200.825 ;
        RECT 16.165 199.435 16.420 200.340 ;
        RECT 16.590 200.195 17.305 200.365 ;
        RECT 16.590 199.265 16.920 200.025 ;
        RECT 17.135 199.435 17.305 200.195 ;
        RECT 18.035 199.265 18.330 200.075 ;
        RECT 18.510 199.435 18.755 200.575 ;
        RECT 18.930 199.265 19.190 200.075 ;
        RECT 19.370 199.440 19.620 200.575 ;
        RECT 25.800 200.405 26.965 200.995 ;
        RECT 20.220 200.180 26.965 200.405 ;
        RECT 27.315 200.995 34.060 201.165 ;
        RECT 27.315 200.405 28.480 200.995 ;
        RECT 34.660 200.825 34.910 201.635 ;
        RECT 35.090 201.290 35.350 201.815 ;
        RECT 35.520 200.825 35.770 201.635 ;
        RECT 35.950 201.305 36.255 201.815 ;
        RECT 28.650 200.575 35.770 200.825 ;
        RECT 35.940 200.575 36.255 201.135 ;
        RECT 36.425 201.090 36.715 201.815 ;
        RECT 36.885 201.305 37.190 201.815 ;
        RECT 36.885 200.575 37.200 201.135 ;
        RECT 37.370 200.825 37.620 201.635 ;
        RECT 37.790 201.290 38.050 201.815 ;
        RECT 38.230 200.825 38.480 201.635 ;
        RECT 38.650 201.255 38.910 201.815 ;
        RECT 39.080 201.165 39.340 201.620 ;
        RECT 39.510 201.335 39.770 201.815 ;
        RECT 39.940 201.165 40.200 201.620 ;
        RECT 40.370 201.335 40.630 201.815 ;
        RECT 40.800 201.165 41.060 201.620 ;
        RECT 41.230 201.335 41.475 201.815 ;
        RECT 41.645 201.165 41.920 201.620 ;
        RECT 42.090 201.335 42.335 201.815 ;
        RECT 42.505 201.165 42.765 201.620 ;
        RECT 42.945 201.335 43.195 201.815 ;
        RECT 43.365 201.165 43.625 201.620 ;
        RECT 43.805 201.335 44.055 201.815 ;
        RECT 44.225 201.165 44.485 201.620 ;
        RECT 44.665 201.335 44.925 201.815 ;
        RECT 45.095 201.165 45.355 201.620 ;
        RECT 45.525 201.335 45.825 201.815 ;
        RECT 39.080 200.995 45.825 201.165 ;
        RECT 37.370 200.575 44.490 200.825 ;
        RECT 27.315 200.180 34.060 200.405 ;
        RECT 20.220 200.165 25.625 200.180 ;
        RECT 19.790 199.270 20.050 200.065 ;
        RECT 20.220 199.440 20.480 200.165 ;
        RECT 20.650 199.270 20.910 199.995 ;
        RECT 21.080 199.440 21.340 200.165 ;
        RECT 21.510 199.270 21.770 199.995 ;
        RECT 21.940 199.440 22.200 200.165 ;
        RECT 22.370 199.270 22.630 199.995 ;
        RECT 22.800 199.440 23.060 200.165 ;
        RECT 23.230 199.270 23.475 199.995 ;
        RECT 23.645 199.440 23.905 200.165 ;
        RECT 24.090 199.270 24.335 199.995 ;
        RECT 24.505 199.440 24.765 200.165 ;
        RECT 24.950 199.270 25.195 199.995 ;
        RECT 25.365 199.440 25.625 200.165 ;
        RECT 25.810 199.270 26.065 199.995 ;
        RECT 26.235 199.440 26.525 200.180 ;
        RECT 19.790 199.265 26.065 199.270 ;
        RECT 26.695 199.265 26.965 200.010 ;
        RECT 27.315 199.265 27.585 200.010 ;
        RECT 27.755 199.440 28.045 200.180 ;
        RECT 28.655 200.165 34.060 200.180 ;
        RECT 28.215 199.270 28.470 199.995 ;
        RECT 28.655 199.440 28.915 200.165 ;
        RECT 29.085 199.270 29.330 199.995 ;
        RECT 29.515 199.440 29.775 200.165 ;
        RECT 29.945 199.270 30.190 199.995 ;
        RECT 30.375 199.440 30.635 200.165 ;
        RECT 30.805 199.270 31.050 199.995 ;
        RECT 31.220 199.440 31.480 200.165 ;
        RECT 31.650 199.270 31.910 199.995 ;
        RECT 32.080 199.440 32.340 200.165 ;
        RECT 32.510 199.270 32.770 199.995 ;
        RECT 32.940 199.440 33.200 200.165 ;
        RECT 33.370 199.270 33.630 199.995 ;
        RECT 33.800 199.440 34.060 200.165 ;
        RECT 34.230 199.270 34.490 200.065 ;
        RECT 34.660 199.440 34.910 200.575 ;
        RECT 28.215 199.265 34.490 199.270 ;
        RECT 35.090 199.265 35.350 200.075 ;
        RECT 35.525 199.435 35.770 200.575 ;
        RECT 35.950 199.265 36.245 200.075 ;
        RECT 36.425 199.265 36.715 200.430 ;
        RECT 36.895 199.265 37.190 200.075 ;
        RECT 37.370 199.435 37.615 200.575 ;
        RECT 37.790 199.265 38.050 200.075 ;
        RECT 38.230 199.440 38.480 200.575 ;
        RECT 44.660 200.405 45.825 200.995 ;
        RECT 39.080 200.180 45.825 200.405 ;
        RECT 39.080 200.165 44.485 200.180 ;
        RECT 38.650 199.270 38.910 200.065 ;
        RECT 39.080 199.440 39.340 200.165 ;
        RECT 39.510 199.270 39.770 199.995 ;
        RECT 39.940 199.440 40.200 200.165 ;
        RECT 40.370 199.270 40.630 199.995 ;
        RECT 40.800 199.440 41.060 200.165 ;
        RECT 41.230 199.270 41.490 199.995 ;
        RECT 41.660 199.440 41.920 200.165 ;
        RECT 42.090 199.270 42.335 199.995 ;
        RECT 42.505 199.440 42.765 200.165 ;
        RECT 42.950 199.270 43.195 199.995 ;
        RECT 43.365 199.440 43.625 200.165 ;
        RECT 43.810 199.270 44.055 199.995 ;
        RECT 44.225 199.440 44.485 200.165 ;
        RECT 44.670 199.270 44.925 199.995 ;
        RECT 45.095 199.440 45.385 200.180 ;
        RECT 38.650 199.265 44.925 199.270 ;
        RECT 45.555 199.265 45.825 200.010 ;
        RECT 46.100 199.445 46.380 201.635 ;
        RECT 46.580 201.445 47.310 201.815 ;
        RECT 47.890 201.275 48.320 201.635 ;
        RECT 46.580 201.085 48.320 201.275 ;
        RECT 46.580 200.575 46.840 201.085 ;
        RECT 46.570 199.265 46.855 200.405 ;
        RECT 47.050 200.285 47.310 200.905 ;
        RECT 47.505 200.285 47.930 200.905 ;
        RECT 48.100 200.855 48.320 201.085 ;
        RECT 48.490 201.035 48.735 201.815 ;
        RECT 48.100 200.555 48.645 200.855 ;
        RECT 48.935 200.735 49.165 201.635 ;
        RECT 47.120 199.915 48.145 200.115 ;
        RECT 47.120 199.445 47.290 199.915 ;
        RECT 47.465 199.265 47.795 199.745 ;
        RECT 47.965 199.445 48.145 199.915 ;
        RECT 48.315 199.445 48.645 200.555 ;
        RECT 48.825 200.055 49.165 200.735 ;
        RECT 49.345 200.235 49.575 201.575 ;
        RECT 50.225 201.435 50.555 201.815 ;
        RECT 49.780 201.265 50.055 201.405 ;
        RECT 50.725 201.265 50.935 201.435 ;
        RECT 49.780 201.075 50.935 201.265 ;
        RECT 51.105 201.265 51.435 201.645 ;
        RECT 51.625 201.435 51.955 201.815 ;
        RECT 51.105 201.060 51.955 201.265 ;
        RECT 49.775 200.450 50.035 200.905 ;
        RECT 50.290 200.795 50.875 200.875 ;
        RECT 50.285 200.625 50.875 200.795 ;
        RECT 50.290 200.500 50.875 200.625 ;
        RECT 48.825 199.855 49.575 200.055 ;
        RECT 48.815 199.265 49.165 199.675 ;
        RECT 49.335 199.465 49.575 199.855 ;
        RECT 49.780 199.265 50.105 200.250 ;
        RECT 50.290 199.915 50.495 200.500 ;
        RECT 51.045 200.285 51.455 200.890 ;
        RECT 51.625 200.570 51.955 201.060 ;
        RECT 51.625 200.115 51.795 200.570 ;
        RECT 50.675 199.895 51.795 200.115 ;
        RECT 50.675 199.435 50.935 199.895 ;
        RECT 51.105 199.265 51.955 199.715 ;
        RECT 52.125 199.435 52.370 201.645 ;
        RECT 52.555 201.015 52.795 201.815 ;
        RECT 52.985 201.315 53.285 201.645 ;
        RECT 53.455 201.335 53.730 201.815 ;
        RECT 52.985 200.405 53.155 201.315 ;
        RECT 53.910 201.165 54.205 201.555 ;
        RECT 54.375 201.335 54.630 201.815 ;
        RECT 54.805 201.165 55.065 201.555 ;
        RECT 55.235 201.335 55.515 201.815 ;
        RECT 53.325 200.575 53.675 201.145 ;
        RECT 53.910 200.995 55.560 201.165 ;
        RECT 55.750 200.995 56.025 201.815 ;
        RECT 56.195 201.175 56.525 201.645 ;
        RECT 56.695 201.345 56.865 201.815 ;
        RECT 57.035 201.175 57.365 201.645 ;
        RECT 57.535 201.345 57.825 201.815 ;
        RECT 59.010 201.355 59.760 201.645 ;
        RECT 60.270 201.355 60.600 201.815 ;
        RECT 56.195 201.165 57.365 201.175 ;
        RECT 56.195 201.135 57.795 201.165 ;
        RECT 56.195 200.995 57.815 201.135 ;
        RECT 53.845 200.655 54.985 200.825 ;
        RECT 53.845 200.405 54.015 200.655 ;
        RECT 55.155 200.485 55.560 200.995 ;
        RECT 57.580 200.965 57.815 200.995 ;
        RECT 55.750 200.625 56.470 200.825 ;
        RECT 56.640 200.625 57.410 200.825 ;
        RECT 52.555 199.265 52.810 200.265 ;
        RECT 52.985 200.235 54.015 200.405 ;
        RECT 54.805 200.315 55.560 200.485 ;
        RECT 57.580 200.455 57.795 200.965 ;
        RECT 52.985 199.435 53.295 200.235 ;
        RECT 54.805 200.065 55.065 200.315 ;
        RECT 55.750 200.235 56.865 200.445 ;
        RECT 53.465 199.265 53.775 200.065 ;
        RECT 53.945 199.895 55.065 200.065 ;
        RECT 53.945 199.435 54.205 199.895 ;
        RECT 54.375 199.265 54.630 199.725 ;
        RECT 54.805 199.435 55.065 199.895 ;
        RECT 55.235 199.265 55.520 200.135 ;
        RECT 55.750 199.435 56.025 200.235 ;
        RECT 56.195 199.265 56.525 200.065 ;
        RECT 56.695 199.605 56.865 200.235 ;
        RECT 57.035 200.235 57.795 200.455 ;
        RECT 57.035 199.775 57.365 200.235 ;
        RECT 59.010 200.065 59.380 201.355 ;
        RECT 60.820 201.165 61.090 201.375 ;
        RECT 59.755 200.995 61.090 201.165 ;
        RECT 62.185 201.090 62.475 201.815 ;
        RECT 62.645 201.140 62.905 201.645 ;
        RECT 63.085 201.435 63.415 201.815 ;
        RECT 63.595 201.265 63.765 201.645 ;
        RECT 59.755 200.825 59.925 200.995 ;
        RECT 59.550 200.575 59.925 200.825 ;
        RECT 60.095 200.585 60.570 200.825 ;
        RECT 60.740 200.585 61.090 200.825 ;
        RECT 59.755 200.405 59.925 200.575 ;
        RECT 59.755 200.235 61.090 200.405 ;
        RECT 60.810 200.075 61.090 200.235 ;
        RECT 57.535 199.605 57.835 200.065 ;
        RECT 59.010 199.895 60.180 200.065 ;
        RECT 56.695 199.435 57.835 199.605 ;
        RECT 59.465 199.265 59.680 199.725 ;
        RECT 59.850 199.435 60.180 199.895 ;
        RECT 60.350 199.265 60.600 200.065 ;
        RECT 62.185 199.265 62.475 200.430 ;
        RECT 62.645 200.340 62.815 201.140 ;
        RECT 63.100 201.095 63.765 201.265 ;
        RECT 63.100 200.840 63.270 201.095 ;
        RECT 62.985 200.510 63.270 200.840 ;
        RECT 63.505 200.545 63.835 200.915 ;
        RECT 63.100 200.365 63.270 200.510 ;
        RECT 62.645 199.435 62.915 200.340 ;
        RECT 63.100 200.195 63.765 200.365 ;
        RECT 63.085 199.265 63.415 200.025 ;
        RECT 63.595 199.435 63.765 200.195 ;
        RECT 64.025 199.435 64.775 201.645 ;
        RECT 64.970 201.425 65.300 201.815 ;
        RECT 65.470 201.255 65.695 201.635 ;
        RECT 64.955 200.575 65.195 201.225 ;
        RECT 65.365 201.075 65.695 201.255 ;
        RECT 65.365 200.405 65.540 201.075 ;
        RECT 65.895 200.905 66.125 201.525 ;
        RECT 66.305 201.085 66.605 201.815 ;
        RECT 67.265 201.315 67.520 201.645 ;
        RECT 67.735 201.335 68.065 201.815 ;
        RECT 68.235 201.395 69.770 201.645 ;
        RECT 67.265 201.235 67.450 201.315 ;
        RECT 65.710 200.575 66.125 200.905 ;
        RECT 66.305 200.575 66.600 200.905 ;
        RECT 64.955 200.215 65.540 200.405 ;
        RECT 64.955 199.445 65.230 200.215 ;
        RECT 65.710 200.045 66.605 200.375 ;
        RECT 65.400 199.875 66.605 200.045 ;
        RECT 65.400 199.445 65.730 199.875 ;
        RECT 65.900 199.265 66.095 199.705 ;
        RECT 66.275 199.445 66.605 199.875 ;
        RECT 67.265 200.105 67.435 201.235 ;
        RECT 68.235 201.165 68.405 201.395 ;
        RECT 67.605 200.995 68.405 201.165 ;
        RECT 67.605 200.445 67.775 200.995 ;
        RECT 68.585 200.825 68.870 201.225 ;
        RECT 68.005 200.625 68.370 200.825 ;
        RECT 68.540 200.625 68.870 200.825 ;
        RECT 69.140 200.825 69.420 201.225 ;
        RECT 69.600 201.165 69.770 201.395 ;
        RECT 69.995 201.335 70.325 201.815 ;
        RECT 70.495 201.165 70.665 201.645 ;
        RECT 69.600 200.995 70.665 201.165 ;
        RECT 70.965 200.995 71.195 201.815 ;
        RECT 71.365 201.015 71.695 201.645 ;
        RECT 69.140 200.625 69.615 200.825 ;
        RECT 69.785 200.625 70.230 200.825 ;
        RECT 70.400 200.615 70.750 200.825 ;
        RECT 70.945 200.575 71.275 200.825 ;
        RECT 67.605 200.275 70.665 200.445 ;
        RECT 71.445 200.415 71.695 201.015 ;
        RECT 71.865 200.995 72.075 201.815 ;
        RECT 72.305 201.140 72.565 201.645 ;
        RECT 72.745 201.435 73.075 201.815 ;
        RECT 73.255 201.265 73.425 201.645 ;
        RECT 67.265 199.435 67.520 200.105 ;
        RECT 67.690 199.265 68.020 200.025 ;
        RECT 68.190 199.865 69.825 200.105 ;
        RECT 68.190 199.435 68.440 199.865 ;
        RECT 69.595 199.775 69.825 199.865 ;
        RECT 68.610 199.265 68.965 199.685 ;
        RECT 69.155 199.605 69.485 199.645 ;
        RECT 69.995 199.605 70.325 200.105 ;
        RECT 69.155 199.435 70.325 199.605 ;
        RECT 70.495 199.435 70.665 200.275 ;
        RECT 70.965 199.265 71.195 200.405 ;
        RECT 71.365 199.435 71.695 200.415 ;
        RECT 71.865 199.265 72.075 200.405 ;
        RECT 72.305 200.340 72.475 201.140 ;
        RECT 72.760 201.095 73.425 201.265 ;
        RECT 72.760 200.840 72.930 201.095 ;
        RECT 74.615 201.085 74.915 201.815 ;
        RECT 72.645 200.510 72.930 200.840 ;
        RECT 73.165 200.545 73.495 200.915 ;
        RECT 75.095 200.905 75.325 201.525 ;
        RECT 75.525 201.255 75.750 201.635 ;
        RECT 75.920 201.425 76.250 201.815 ;
        RECT 75.525 201.075 75.855 201.255 ;
        RECT 74.620 200.575 74.915 200.905 ;
        RECT 75.095 200.575 75.510 200.905 ;
        RECT 72.760 200.365 72.930 200.510 ;
        RECT 75.680 200.405 75.855 201.075 ;
        RECT 76.025 200.575 76.265 201.225 ;
        RECT 76.465 201.085 76.755 201.815 ;
        RECT 76.455 200.575 76.755 200.905 ;
        RECT 76.935 200.885 77.165 201.525 ;
        RECT 77.345 201.265 77.655 201.635 ;
        RECT 77.835 201.445 78.505 201.815 ;
        RECT 77.345 201.065 78.575 201.265 ;
        RECT 76.935 200.575 77.460 200.885 ;
        RECT 77.640 200.575 78.105 200.885 ;
        RECT 72.305 199.435 72.575 200.340 ;
        RECT 72.760 200.195 73.425 200.365 ;
        RECT 72.745 199.265 73.075 200.025 ;
        RECT 73.255 199.435 73.425 200.195 ;
        RECT 74.615 200.045 75.510 200.375 ;
        RECT 75.680 200.215 76.265 200.405 ;
        RECT 78.285 200.395 78.575 201.065 ;
        RECT 74.615 199.875 75.820 200.045 ;
        RECT 74.615 199.445 74.945 199.875 ;
        RECT 75.125 199.265 75.320 199.705 ;
        RECT 75.490 199.445 75.820 199.875 ;
        RECT 75.990 199.445 76.265 200.215 ;
        RECT 76.465 200.155 77.625 200.395 ;
        RECT 76.465 199.445 76.725 200.155 ;
        RECT 76.895 199.265 77.225 199.975 ;
        RECT 77.395 199.445 77.625 200.155 ;
        RECT 77.805 200.175 78.575 200.395 ;
        RECT 77.805 199.445 78.075 200.175 ;
        RECT 78.255 199.265 78.595 199.995 ;
        RECT 78.765 199.445 79.025 201.635 ;
        RECT 79.205 201.065 80.415 201.815 ;
        RECT 80.590 201.270 85.935 201.815 ;
        RECT 79.205 200.355 79.725 200.895 ;
        RECT 79.895 200.525 80.415 201.065 ;
        RECT 79.205 199.265 80.415 200.355 ;
        RECT 82.180 199.700 82.530 200.950 ;
        RECT 84.010 200.440 84.350 201.270 ;
        RECT 86.195 201.265 86.365 201.645 ;
        RECT 86.580 201.435 86.910 201.815 ;
        RECT 86.195 201.095 86.910 201.265 ;
        RECT 86.105 200.545 86.460 200.915 ;
        RECT 86.740 200.905 86.910 201.095 ;
        RECT 87.080 201.070 87.335 201.645 ;
        RECT 86.740 200.575 86.995 200.905 ;
        RECT 86.740 200.365 86.910 200.575 ;
        RECT 86.195 200.195 86.910 200.365 ;
        RECT 87.165 200.340 87.335 201.070 ;
        RECT 87.510 200.975 87.770 201.815 ;
        RECT 87.945 201.090 88.235 201.815 ;
        RECT 88.865 201.230 89.175 201.645 ;
        RECT 89.370 201.435 89.700 201.815 ;
        RECT 89.870 201.475 91.275 201.645 ;
        RECT 89.870 201.245 90.040 201.475 ;
        RECT 80.590 199.265 85.935 199.700 ;
        RECT 86.195 199.435 86.365 200.195 ;
        RECT 86.580 199.265 86.910 200.025 ;
        RECT 87.080 199.435 87.335 200.340 ;
        RECT 87.510 199.265 87.770 200.415 ;
        RECT 87.945 199.265 88.235 200.430 ;
        RECT 88.865 200.115 89.035 201.230 ;
        RECT 89.345 201.075 90.040 201.245 ;
        RECT 91.105 201.245 91.275 201.475 ;
        RECT 91.545 201.415 91.875 201.815 ;
        RECT 92.115 201.245 92.285 201.645 ;
        RECT 89.345 200.905 89.515 201.075 ;
        RECT 89.205 200.575 89.515 200.905 ;
        RECT 89.685 200.575 90.020 200.905 ;
        RECT 90.290 200.575 90.485 201.150 ;
        RECT 90.745 200.905 90.935 201.135 ;
        RECT 91.105 201.075 92.285 201.245 ;
        RECT 93.050 201.355 93.800 201.645 ;
        RECT 94.310 201.355 94.640 201.815 ;
        RECT 90.745 200.575 91.090 200.905 ;
        RECT 91.400 200.575 91.875 200.905 ;
        RECT 92.130 200.575 92.315 200.905 ;
        RECT 89.345 200.405 89.515 200.575 ;
        RECT 89.345 200.235 92.285 200.405 ;
        RECT 88.865 199.475 89.205 200.115 ;
        RECT 89.795 199.895 91.355 200.065 ;
        RECT 89.375 199.265 89.620 199.725 ;
        RECT 89.795 199.435 90.045 199.895 ;
        RECT 90.235 199.265 90.905 199.645 ;
        RECT 91.105 199.435 91.355 199.895 ;
        RECT 92.115 199.435 92.285 200.235 ;
        RECT 93.050 200.065 93.420 201.355 ;
        RECT 94.860 201.165 95.130 201.375 ;
        RECT 93.795 200.995 95.130 201.165 ;
        RECT 95.325 201.005 95.565 201.815 ;
        RECT 95.735 201.005 96.065 201.645 ;
        RECT 96.235 201.005 96.505 201.815 ;
        RECT 97.145 201.045 99.735 201.815 ;
        RECT 93.795 200.825 93.965 200.995 ;
        RECT 93.590 200.575 93.965 200.825 ;
        RECT 94.135 200.585 94.610 200.825 ;
        RECT 94.780 200.585 95.130 200.825 ;
        RECT 95.305 200.575 95.655 200.825 ;
        RECT 93.795 200.405 93.965 200.575 ;
        RECT 95.825 200.405 95.995 201.005 ;
        RECT 96.165 200.575 96.515 200.825 ;
        RECT 93.795 200.235 95.130 200.405 ;
        RECT 94.850 200.075 95.130 200.235 ;
        RECT 95.315 200.235 95.995 200.405 ;
        RECT 93.050 199.895 94.220 200.065 ;
        RECT 93.505 199.265 93.720 199.725 ;
        RECT 93.890 199.435 94.220 199.895 ;
        RECT 94.390 199.265 94.640 200.065 ;
        RECT 95.315 199.450 95.645 200.235 ;
        RECT 96.175 199.265 96.505 200.405 ;
        RECT 97.145 200.355 98.355 200.875 ;
        RECT 98.525 200.525 99.735 201.045 ;
        RECT 97.145 199.265 99.735 200.355 ;
        RECT 99.910 200.215 100.245 201.635 ;
        RECT 100.425 201.445 101.170 201.815 ;
        RECT 101.735 201.275 101.990 201.635 ;
        RECT 102.170 201.445 102.500 201.815 ;
        RECT 102.680 201.275 102.905 201.635 ;
        RECT 100.420 201.085 102.905 201.275 ;
        RECT 100.420 200.395 100.645 201.085 ;
        RECT 103.585 201.045 106.175 201.815 ;
        RECT 100.845 200.575 101.125 200.905 ;
        RECT 101.305 200.575 101.880 200.905 ;
        RECT 102.060 200.575 102.495 200.905 ;
        RECT 102.675 200.575 102.945 200.905 ;
        RECT 100.420 200.215 102.915 200.395 ;
        RECT 99.910 199.445 100.175 200.215 ;
        RECT 100.345 199.265 100.675 199.985 ;
        RECT 100.865 199.805 102.055 200.035 ;
        RECT 100.865 199.445 101.125 199.805 ;
        RECT 101.295 199.265 101.625 199.635 ;
        RECT 101.795 199.445 102.055 199.805 ;
        RECT 102.625 199.445 102.915 200.215 ;
        RECT 103.585 200.355 104.795 200.875 ;
        RECT 104.965 200.525 106.175 201.045 ;
        RECT 106.365 201.125 106.605 201.645 ;
        RECT 106.775 201.320 107.170 201.815 ;
        RECT 107.735 201.485 107.905 201.630 ;
        RECT 107.530 201.290 107.905 201.485 ;
        RECT 106.365 200.455 106.540 201.125 ;
        RECT 107.530 200.955 107.700 201.290 ;
        RECT 108.185 201.245 108.425 201.620 ;
        RECT 108.595 201.310 108.930 201.815 ;
        RECT 108.185 201.095 108.405 201.245 ;
        RECT 109.105 201.180 109.375 201.815 ;
        RECT 106.715 200.595 107.700 200.955 ;
        RECT 107.870 200.765 108.405 201.095 ;
        RECT 106.715 200.575 108.000 200.595 ;
        RECT 103.585 199.265 106.175 200.355 ;
        RECT 106.365 200.320 106.575 200.455 ;
        RECT 107.140 200.425 108.000 200.575 ;
        RECT 106.365 199.535 106.670 200.320 ;
        RECT 106.845 199.945 107.540 200.255 ;
        RECT 106.850 199.265 107.535 199.735 ;
        RECT 107.715 199.480 108.000 200.425 ;
        RECT 108.170 200.115 108.405 200.765 ;
        RECT 108.575 200.285 108.875 201.135 ;
        RECT 109.560 201.125 109.795 201.645 ;
        RECT 109.965 201.320 110.365 201.815 ;
        RECT 110.955 201.485 111.125 201.630 ;
        RECT 110.725 201.290 111.125 201.485 ;
        RECT 109.560 200.320 109.735 201.125 ;
        RECT 110.725 200.955 110.895 201.290 ;
        RECT 111.405 201.245 111.645 201.620 ;
        RECT 111.815 201.310 112.145 201.815 ;
        RECT 111.405 201.095 111.620 201.245 ;
        RECT 109.905 200.595 110.895 200.955 ;
        RECT 111.065 200.765 111.620 201.095 ;
        RECT 109.905 200.575 111.195 200.595 ;
        RECT 110.335 200.425 111.195 200.575 ;
        RECT 108.170 199.885 108.845 200.115 ;
        RECT 108.175 199.265 108.505 199.715 ;
        RECT 108.675 199.455 108.845 199.885 ;
        RECT 109.105 199.265 109.375 200.220 ;
        RECT 109.560 199.535 109.865 200.320 ;
        RECT 110.040 199.945 110.735 200.255 ;
        RECT 110.045 199.265 110.730 199.735 ;
        RECT 110.910 199.480 111.195 200.425 ;
        RECT 111.385 200.115 111.620 200.765 ;
        RECT 111.790 200.965 112.095 201.135 ;
        RECT 112.325 201.065 113.535 201.815 ;
        RECT 113.705 201.090 113.995 201.815 ;
        RECT 114.630 201.270 119.975 201.815 ;
        RECT 120.150 201.270 125.495 201.815 ;
        RECT 111.790 200.285 112.090 200.965 ;
        RECT 112.325 200.355 112.845 200.895 ;
        RECT 113.015 200.525 113.535 201.065 ;
        RECT 111.385 199.885 112.065 200.115 ;
        RECT 111.395 199.265 111.725 199.715 ;
        RECT 111.895 199.455 112.065 199.885 ;
        RECT 112.325 199.265 113.535 200.355 ;
        RECT 113.705 199.265 113.995 200.430 ;
        RECT 116.220 199.700 116.570 200.950 ;
        RECT 118.050 200.440 118.390 201.270 ;
        RECT 121.740 199.700 122.090 200.950 ;
        RECT 123.570 200.440 123.910 201.270 ;
        RECT 125.665 201.065 126.875 201.815 ;
        RECT 125.665 200.355 126.185 200.895 ;
        RECT 126.355 200.525 126.875 201.065 ;
        RECT 114.630 199.265 119.975 199.700 ;
        RECT 120.150 199.265 125.495 199.700 ;
        RECT 125.665 199.265 126.875 200.355 ;
        RECT 14.260 199.095 126.960 199.265 ;
        RECT 14.345 198.005 15.555 199.095 ;
        RECT 14.345 197.295 14.865 197.835 ;
        RECT 15.035 197.465 15.555 198.005 ;
        RECT 15.725 197.805 15.995 198.905 ;
        RECT 16.165 198.165 16.440 198.670 ;
        RECT 16.610 198.335 16.940 199.095 ;
        RECT 16.165 197.995 16.655 198.165 ;
        RECT 17.110 198.085 17.435 198.925 ;
        RECT 15.725 197.455 16.175 197.805 ;
        RECT 16.360 197.455 16.655 197.995 ;
        RECT 16.825 197.915 17.435 198.085 ;
        RECT 17.910 197.995 18.285 199.095 ;
        RECT 18.555 198.255 18.805 199.095 ;
        RECT 18.975 198.085 19.225 198.925 ;
        RECT 19.395 198.255 19.645 199.095 ;
        RECT 19.815 198.085 20.065 198.925 ;
        RECT 20.290 198.255 20.540 199.095 ;
        RECT 20.825 198.245 21.125 198.835 ;
        RECT 18.495 197.915 20.065 198.085 ;
        RECT 14.345 196.545 15.555 197.295 ;
        RECT 16.360 197.285 16.530 197.455 ;
        RECT 16.825 197.285 16.995 197.915 ;
        RECT 17.165 197.535 17.665 197.745 ;
        RECT 17.835 197.535 18.315 197.745 ;
        RECT 18.495 197.365 18.735 197.915 ;
        RECT 20.270 197.905 20.705 198.075 ;
        RECT 18.905 197.535 20.365 197.705 ;
        RECT 15.725 196.545 16.000 197.285 ;
        RECT 16.220 197.115 16.530 197.285 ;
        RECT 16.220 196.955 16.410 197.115 ;
        RECT 16.755 197.105 16.995 197.285 ;
        RECT 17.210 197.195 18.305 197.365 ;
        RECT 16.755 197.055 16.925 197.105 ;
        RECT 16.705 196.885 16.925 197.055 ;
        RECT 17.210 196.945 17.380 197.195 ;
        RECT 16.755 196.715 16.925 196.885 ;
        RECT 17.130 196.715 17.460 196.945 ;
        RECT 17.635 196.545 17.805 197.015 ;
        RECT 17.975 196.730 18.305 197.195 ;
        RECT 18.495 197.185 20.025 197.365 ;
        RECT 18.595 196.545 18.765 197.015 ;
        RECT 18.935 196.715 19.265 197.185 ;
        RECT 19.435 196.545 19.605 197.015 ;
        RECT 19.775 196.715 20.025 197.185 ;
        RECT 20.195 197.285 20.365 197.535 ;
        RECT 20.535 197.455 20.705 197.905 ;
        RECT 20.935 197.910 21.125 198.245 ;
        RECT 21.305 198.080 21.665 198.835 ;
        RECT 22.095 198.205 22.425 198.910 ;
        RECT 20.935 197.455 21.265 197.910 ;
        RECT 21.495 197.455 21.665 198.080 ;
        RECT 21.835 198.035 22.425 198.205 ;
        RECT 22.675 198.525 22.865 198.915 ;
        RECT 23.095 198.595 23.375 199.095 ;
        RECT 21.835 197.285 22.005 198.035 ;
        RECT 22.675 197.785 22.845 198.525 ;
        RECT 22.245 197.455 22.845 197.785 ;
        RECT 23.015 197.455 23.355 198.415 ;
        RECT 23.545 197.930 23.835 199.095 ;
        RECT 24.010 198.585 25.665 198.875 ;
        RECT 24.010 198.245 25.600 198.415 ;
        RECT 25.835 198.295 26.115 199.095 ;
        RECT 24.010 197.955 24.330 198.245 ;
        RECT 25.430 198.125 25.600 198.245 ;
        RECT 24.525 197.905 25.240 198.075 ;
        RECT 25.430 197.955 26.155 198.125 ;
        RECT 26.325 197.955 26.595 198.925 ;
        RECT 27.015 198.365 27.310 199.095 ;
        RECT 27.480 198.195 27.740 198.920 ;
        RECT 27.910 198.365 28.170 199.095 ;
        RECT 28.340 198.195 28.600 198.920 ;
        RECT 28.770 198.365 29.030 199.095 ;
        RECT 29.200 198.195 29.460 198.920 ;
        RECT 29.630 198.365 29.890 199.095 ;
        RECT 30.060 198.195 30.320 198.920 ;
        RECT 20.195 197.115 22.005 197.285 ;
        RECT 22.675 197.365 22.845 197.455 ;
        RECT 20.205 196.545 20.585 196.945 ;
        RECT 20.805 196.765 20.975 197.115 ;
        RECT 21.145 196.545 21.475 196.945 ;
        RECT 21.675 196.765 21.845 197.115 ;
        RECT 22.175 196.545 22.425 197.045 ;
        RECT 22.675 196.895 22.865 197.365 ;
        RECT 23.115 196.545 23.375 197.285 ;
        RECT 23.545 196.545 23.835 197.270 ;
        RECT 24.010 197.215 24.360 197.785 ;
        RECT 24.530 197.455 25.240 197.905 ;
        RECT 25.985 197.785 26.155 197.955 ;
        RECT 25.410 197.455 25.815 197.785 ;
        RECT 25.985 197.455 26.255 197.785 ;
        RECT 25.985 197.285 26.155 197.455 ;
        RECT 24.545 197.115 26.155 197.285 ;
        RECT 26.425 197.220 26.595 197.955 ;
        RECT 24.015 196.545 24.345 197.045 ;
        RECT 24.545 196.765 24.715 197.115 ;
        RECT 24.915 196.545 25.245 196.945 ;
        RECT 25.415 196.765 25.585 197.115 ;
        RECT 25.755 196.545 26.135 196.945 ;
        RECT 26.325 196.875 26.595 197.220 ;
        RECT 27.010 197.955 30.320 198.195 ;
        RECT 30.490 197.985 30.750 199.095 ;
        RECT 27.010 197.365 27.980 197.955 ;
        RECT 30.920 197.785 31.170 198.920 ;
        RECT 31.350 197.985 31.645 199.095 ;
        RECT 31.915 198.350 32.185 199.095 ;
        RECT 32.815 199.090 39.090 199.095 ;
        RECT 32.355 198.180 32.645 198.920 ;
        RECT 32.815 198.365 33.070 199.090 ;
        RECT 33.255 198.195 33.515 198.920 ;
        RECT 33.685 198.365 33.930 199.090 ;
        RECT 34.115 198.195 34.375 198.920 ;
        RECT 34.545 198.365 34.790 199.090 ;
        RECT 34.975 198.195 35.235 198.920 ;
        RECT 35.405 198.365 35.650 199.090 ;
        RECT 35.820 198.195 36.080 198.920 ;
        RECT 36.250 198.365 36.510 199.090 ;
        RECT 36.680 198.195 36.940 198.920 ;
        RECT 37.110 198.365 37.370 199.090 ;
        RECT 37.540 198.195 37.800 198.920 ;
        RECT 37.970 198.365 38.230 199.090 ;
        RECT 38.400 198.195 38.660 198.920 ;
        RECT 38.830 198.295 39.090 199.090 ;
        RECT 33.255 198.180 38.660 198.195 ;
        RECT 31.915 197.955 38.660 198.180 ;
        RECT 28.150 197.535 31.170 197.785 ;
        RECT 27.010 197.195 30.320 197.365 ;
        RECT 27.010 196.545 27.310 197.025 ;
        RECT 27.480 196.740 27.740 197.195 ;
        RECT 27.910 196.545 28.170 197.025 ;
        RECT 28.340 196.740 28.600 197.195 ;
        RECT 28.770 196.545 29.030 197.025 ;
        RECT 29.200 196.740 29.460 197.195 ;
        RECT 29.630 196.545 29.890 197.025 ;
        RECT 30.060 196.740 30.320 197.195 ;
        RECT 30.490 196.545 30.750 197.070 ;
        RECT 30.920 196.725 31.170 197.535 ;
        RECT 31.340 197.175 31.655 197.785 ;
        RECT 31.915 197.365 33.080 197.955 ;
        RECT 39.260 197.785 39.510 198.920 ;
        RECT 39.690 198.285 39.950 199.095 ;
        RECT 40.125 197.785 40.370 198.925 ;
        RECT 40.550 198.285 40.845 199.095 ;
        RECT 41.025 197.955 41.305 199.095 ;
        RECT 41.475 197.945 41.805 198.925 ;
        RECT 41.975 197.955 42.235 199.095 ;
        RECT 42.405 198.675 42.745 199.095 ;
        RECT 42.915 198.505 43.165 198.925 ;
        RECT 42.405 198.335 43.165 198.505 ;
        RECT 41.540 197.905 41.715 197.945 ;
        RECT 33.250 197.535 40.370 197.785 ;
        RECT 31.915 197.195 38.660 197.365 ;
        RECT 31.350 196.545 31.595 197.005 ;
        RECT 31.915 196.545 32.215 197.025 ;
        RECT 32.385 196.740 32.645 197.195 ;
        RECT 32.815 196.545 33.075 197.025 ;
        RECT 33.255 196.740 33.515 197.195 ;
        RECT 33.685 196.545 33.935 197.025 ;
        RECT 34.115 196.740 34.375 197.195 ;
        RECT 34.545 196.545 34.795 197.025 ;
        RECT 34.975 196.740 35.235 197.195 ;
        RECT 35.405 196.545 35.650 197.025 ;
        RECT 35.820 196.740 36.095 197.195 ;
        RECT 36.265 196.545 36.510 197.025 ;
        RECT 36.680 196.740 36.940 197.195 ;
        RECT 37.110 196.545 37.370 197.025 ;
        RECT 37.540 196.740 37.800 197.195 ;
        RECT 37.970 196.545 38.230 197.025 ;
        RECT 38.400 196.740 38.660 197.195 ;
        RECT 38.830 196.545 39.090 197.105 ;
        RECT 39.260 196.725 39.510 197.535 ;
        RECT 39.690 196.545 39.950 197.070 ;
        RECT 40.120 196.725 40.370 197.535 ;
        RECT 40.540 197.225 40.855 197.785 ;
        RECT 41.035 197.515 41.370 197.785 ;
        RECT 41.540 197.345 41.710 197.905 ;
        RECT 41.880 197.535 42.215 197.785 ;
        RECT 42.405 197.365 42.715 198.335 ;
        RECT 43.335 198.255 43.665 199.095 ;
        RECT 44.155 198.505 44.910 198.925 ;
        RECT 43.835 198.335 45.300 198.505 ;
        RECT 43.835 198.085 44.005 198.335 ;
        RECT 43.045 197.915 44.005 198.085 ;
        RECT 43.045 197.745 43.215 197.915 ;
        RECT 44.175 197.745 44.480 198.165 ;
        RECT 42.885 197.535 43.215 197.745 ;
        RECT 43.385 197.535 43.825 197.745 ;
        RECT 43.995 197.535 44.480 197.745 ;
        RECT 44.670 197.735 44.960 198.165 ;
        RECT 45.130 198.130 45.300 198.335 ;
        RECT 45.470 198.310 45.710 199.095 ;
        RECT 45.880 198.130 46.210 198.925 ;
        RECT 46.545 198.590 47.175 199.095 ;
        RECT 45.130 197.955 46.210 198.130 ;
        RECT 46.560 198.055 46.815 198.420 ;
        RECT 46.985 198.415 47.175 198.590 ;
        RECT 47.355 198.585 47.830 198.925 ;
        RECT 46.985 198.225 47.315 198.415 ;
        RECT 47.540 198.055 47.790 198.350 ;
        RECT 48.015 198.250 48.230 199.095 ;
        RECT 48.430 198.255 48.705 198.925 ;
        RECT 45.130 197.905 45.915 197.955 ;
        RECT 44.670 197.535 45.060 197.735 ;
        RECT 45.230 197.535 45.575 197.735 ;
        RECT 40.550 196.545 40.855 197.055 ;
        RECT 41.025 196.545 41.335 197.345 ;
        RECT 41.540 196.715 42.235 197.345 ;
        RECT 42.405 197.195 43.165 197.365 ;
        RECT 42.495 196.545 42.665 197.025 ;
        RECT 42.835 196.725 43.165 197.195 ;
        RECT 43.335 196.545 43.505 197.365 ;
        RECT 43.675 197.195 45.375 197.365 ;
        RECT 43.675 196.730 44.005 197.195 ;
        RECT 44.990 197.105 45.375 197.195 ;
        RECT 45.745 197.265 45.915 197.905 ;
        RECT 46.560 197.885 48.350 198.055 ;
        RECT 48.535 197.905 48.705 198.255 ;
        RECT 48.875 198.085 49.135 199.095 ;
        RECT 49.305 197.930 49.595 199.095 ;
        RECT 49.855 198.165 50.025 198.925 ;
        RECT 50.205 198.335 50.535 199.095 ;
        RECT 49.855 197.995 50.520 198.165 ;
        RECT 50.705 198.020 50.975 198.925 ;
        RECT 46.115 197.435 46.375 197.785 ;
        RECT 45.745 197.095 46.290 197.265 ;
        RECT 46.545 197.225 46.930 197.705 ;
        RECT 44.175 196.545 44.345 197.015 ;
        RECT 44.605 196.755 45.790 196.925 ;
        RECT 45.960 196.715 46.290 197.095 ;
        RECT 47.100 197.030 47.355 197.885 ;
        RECT 46.565 196.765 47.355 197.030 ;
        RECT 47.525 197.210 47.935 197.705 ;
        RECT 48.120 197.455 48.350 197.885 ;
        RECT 48.520 197.385 49.135 197.905 ;
        RECT 50.350 197.850 50.520 197.995 ;
        RECT 49.785 197.445 50.115 197.815 ;
        RECT 50.350 197.520 50.635 197.850 ;
        RECT 47.525 196.765 47.755 197.210 ;
        RECT 48.520 197.175 48.690 197.385 ;
        RECT 47.935 196.545 48.265 197.040 ;
        RECT 48.440 196.715 48.690 197.175 ;
        RECT 48.860 196.545 49.135 197.205 ;
        RECT 49.305 196.545 49.595 197.270 ;
        RECT 50.350 197.265 50.520 197.520 ;
        RECT 49.855 197.095 50.520 197.265 ;
        RECT 50.805 197.220 50.975 198.020 ;
        RECT 51.150 198.705 51.485 198.925 ;
        RECT 52.490 198.715 52.845 199.095 ;
        RECT 51.150 198.085 51.405 198.705 ;
        RECT 51.655 198.545 51.885 198.585 ;
        RECT 53.015 198.545 53.265 198.925 ;
        RECT 51.655 198.345 53.265 198.545 ;
        RECT 51.655 198.255 51.840 198.345 ;
        RECT 52.430 198.335 53.265 198.345 ;
        RECT 53.515 198.315 53.765 199.095 ;
        RECT 53.935 198.245 54.195 198.925 ;
        RECT 51.995 198.145 52.325 198.175 ;
        RECT 51.995 198.085 53.795 198.145 ;
        RECT 51.150 197.975 53.855 198.085 ;
        RECT 51.150 197.915 52.325 197.975 ;
        RECT 53.655 197.940 53.855 197.975 ;
        RECT 51.145 197.535 51.635 197.735 ;
        RECT 51.825 197.535 52.300 197.745 ;
        RECT 49.855 196.715 50.025 197.095 ;
        RECT 50.205 196.545 50.535 196.925 ;
        RECT 50.715 196.715 50.975 197.220 ;
        RECT 51.150 196.545 51.605 197.310 ;
        RECT 52.080 197.135 52.300 197.535 ;
        RECT 52.545 197.535 52.875 197.745 ;
        RECT 52.545 197.135 52.755 197.535 ;
        RECT 53.045 197.500 53.455 197.805 ;
        RECT 53.685 197.365 53.855 197.940 ;
        RECT 53.585 197.245 53.855 197.365 ;
        RECT 53.010 197.200 53.855 197.245 ;
        RECT 53.010 197.075 53.765 197.200 ;
        RECT 53.010 196.925 53.180 197.075 ;
        RECT 54.025 197.055 54.195 198.245 ;
        RECT 54.405 197.955 54.635 199.095 ;
        RECT 54.805 197.945 55.135 198.925 ;
        RECT 55.305 197.955 55.515 199.095 ;
        RECT 55.750 198.705 56.085 198.925 ;
        RECT 57.090 198.715 57.445 199.095 ;
        RECT 55.750 198.085 56.005 198.705 ;
        RECT 56.255 198.545 56.485 198.585 ;
        RECT 57.615 198.545 57.865 198.925 ;
        RECT 56.255 198.345 57.865 198.545 ;
        RECT 56.255 198.255 56.440 198.345 ;
        RECT 57.030 198.335 57.865 198.345 ;
        RECT 58.115 198.315 58.365 199.095 ;
        RECT 58.535 198.245 58.795 198.925 ;
        RECT 56.595 198.145 56.925 198.175 ;
        RECT 56.595 198.085 58.395 198.145 ;
        RECT 55.750 197.975 58.455 198.085 ;
        RECT 54.385 197.535 54.715 197.785 ;
        RECT 53.965 197.045 54.195 197.055 ;
        RECT 51.880 196.715 53.180 196.925 ;
        RECT 53.435 196.545 53.765 196.905 ;
        RECT 53.935 196.715 54.195 197.045 ;
        RECT 54.405 196.545 54.635 197.365 ;
        RECT 54.885 197.345 55.135 197.945 ;
        RECT 55.750 197.915 56.925 197.975 ;
        RECT 58.255 197.940 58.455 197.975 ;
        RECT 55.745 197.535 56.235 197.735 ;
        RECT 56.425 197.535 56.900 197.745 ;
        RECT 54.805 196.715 55.135 197.345 ;
        RECT 55.305 196.545 55.515 197.365 ;
        RECT 55.750 196.545 56.205 197.310 ;
        RECT 56.680 197.135 56.900 197.535 ;
        RECT 57.145 197.535 57.475 197.745 ;
        RECT 57.145 197.135 57.355 197.535 ;
        RECT 57.645 197.500 58.055 197.805 ;
        RECT 58.285 197.365 58.455 197.940 ;
        RECT 58.185 197.245 58.455 197.365 ;
        RECT 57.610 197.200 58.455 197.245 ;
        RECT 57.610 197.075 58.365 197.200 ;
        RECT 57.610 196.925 57.780 197.075 ;
        RECT 58.625 197.045 58.795 198.245 ;
        RECT 56.480 196.715 57.780 196.925 ;
        RECT 58.035 196.545 58.365 196.905 ;
        RECT 58.535 196.715 58.795 197.045 ;
        RECT 58.965 196.715 59.715 198.925 ;
        RECT 59.975 198.165 60.145 198.925 ;
        RECT 60.360 198.335 60.690 199.095 ;
        RECT 59.975 197.995 60.690 198.165 ;
        RECT 60.860 198.020 61.115 198.925 ;
        RECT 59.885 197.445 60.240 197.815 ;
        RECT 60.520 197.785 60.690 197.995 ;
        RECT 60.520 197.455 60.775 197.785 ;
        RECT 60.520 197.265 60.690 197.455 ;
        RECT 60.945 197.290 61.115 198.020 ;
        RECT 61.290 197.945 61.550 199.095 ;
        RECT 61.725 198.020 61.995 198.925 ;
        RECT 62.165 198.335 62.495 199.095 ;
        RECT 62.675 198.165 62.845 198.925 ;
        RECT 59.975 197.095 60.690 197.265 ;
        RECT 59.975 196.715 60.145 197.095 ;
        RECT 60.360 196.545 60.690 196.925 ;
        RECT 60.860 196.715 61.115 197.290 ;
        RECT 61.290 196.545 61.550 197.385 ;
        RECT 61.725 197.220 61.895 198.020 ;
        RECT 62.180 197.995 62.845 198.165 ;
        RECT 63.105 198.020 63.375 198.925 ;
        RECT 63.545 198.335 63.875 199.095 ;
        RECT 64.055 198.165 64.235 198.925 ;
        RECT 62.180 197.850 62.350 197.995 ;
        RECT 62.065 197.520 62.350 197.850 ;
        RECT 62.180 197.265 62.350 197.520 ;
        RECT 62.585 197.445 62.915 197.815 ;
        RECT 61.725 196.715 61.985 197.220 ;
        RECT 62.180 197.095 62.845 197.265 ;
        RECT 62.165 196.545 62.495 196.925 ;
        RECT 62.675 196.715 62.845 197.095 ;
        RECT 63.105 197.220 63.285 198.020 ;
        RECT 63.560 197.995 64.235 198.165 ;
        RECT 64.485 198.020 64.755 198.925 ;
        RECT 64.925 198.335 65.255 199.095 ;
        RECT 65.435 198.165 65.615 198.925 ;
        RECT 63.560 197.850 63.730 197.995 ;
        RECT 63.455 197.520 63.730 197.850 ;
        RECT 63.560 197.265 63.730 197.520 ;
        RECT 63.955 197.445 64.295 197.815 ;
        RECT 63.105 196.715 63.365 197.220 ;
        RECT 63.560 197.095 64.225 197.265 ;
        RECT 63.545 196.545 63.875 196.925 ;
        RECT 64.055 196.715 64.225 197.095 ;
        RECT 64.485 197.220 64.665 198.020 ;
        RECT 64.940 197.995 65.615 198.165 ;
        RECT 66.325 198.020 66.595 198.925 ;
        RECT 66.765 198.335 67.095 199.095 ;
        RECT 67.275 198.165 67.455 198.925 ;
        RECT 67.710 198.670 68.045 199.095 ;
        RECT 68.215 198.490 68.400 198.895 ;
        RECT 64.940 197.850 65.110 197.995 ;
        RECT 64.835 197.520 65.110 197.850 ;
        RECT 64.940 197.265 65.110 197.520 ;
        RECT 65.335 197.445 65.675 197.815 ;
        RECT 64.485 196.715 64.745 197.220 ;
        RECT 64.940 197.095 65.605 197.265 ;
        RECT 64.925 196.545 65.255 196.925 ;
        RECT 65.435 196.715 65.605 197.095 ;
        RECT 66.325 197.220 66.505 198.020 ;
        RECT 66.780 197.995 67.455 198.165 ;
        RECT 67.735 198.315 68.400 198.490 ;
        RECT 68.605 198.315 68.935 199.095 ;
        RECT 66.780 197.850 66.950 197.995 ;
        RECT 66.675 197.520 66.950 197.850 ;
        RECT 66.780 197.265 66.950 197.520 ;
        RECT 67.175 197.445 67.515 197.815 ;
        RECT 67.735 197.285 68.075 198.315 ;
        RECT 69.105 198.125 69.375 198.895 ;
        RECT 68.245 197.955 69.375 198.125 ;
        RECT 68.245 197.455 68.495 197.955 ;
        RECT 66.325 196.715 66.585 197.220 ;
        RECT 66.780 197.095 67.445 197.265 ;
        RECT 67.735 197.115 68.420 197.285 ;
        RECT 68.675 197.205 69.035 197.785 ;
        RECT 66.765 196.545 67.095 196.925 ;
        RECT 67.275 196.715 67.445 197.095 ;
        RECT 67.710 196.545 68.045 196.945 ;
        RECT 68.215 196.715 68.420 197.115 ;
        RECT 69.205 197.045 69.375 197.955 ;
        RECT 70.675 198.115 71.005 198.925 ;
        RECT 71.175 198.285 71.345 199.095 ;
        RECT 71.515 198.115 71.845 198.925 ;
        RECT 72.015 198.285 72.185 199.095 ;
        RECT 72.355 198.755 74.465 198.925 ;
        RECT 72.355 198.115 72.605 198.755 ;
        RECT 70.675 197.945 72.605 198.115 ;
        RECT 72.820 198.115 73.205 198.585 ;
        RECT 73.375 198.285 73.545 198.755 ;
        RECT 73.715 198.115 74.045 198.585 ;
        RECT 74.215 198.285 74.465 198.755 ;
        RECT 74.635 198.115 74.885 198.925 ;
        RECT 72.820 197.945 74.885 198.115 ;
        RECT 70.480 197.565 71.615 197.735 ;
        RECT 70.480 197.535 71.590 197.565 ;
        RECT 71.880 197.535 72.535 197.735 ;
        RECT 68.630 196.545 68.905 197.025 ;
        RECT 69.115 196.715 69.375 197.045 ;
        RECT 70.605 197.140 71.765 197.310 ;
        RECT 72.820 197.305 73.110 197.945 ;
        RECT 75.065 197.930 75.355 199.095 ;
        RECT 75.530 198.670 75.865 199.095 ;
        RECT 76.035 198.490 76.220 198.895 ;
        RECT 75.555 198.315 76.220 198.490 ;
        RECT 76.425 198.315 76.755 199.095 ;
        RECT 73.280 197.565 73.915 197.735 ;
        RECT 74.200 197.565 74.835 197.735 ;
        RECT 73.280 197.535 73.910 197.565 ;
        RECT 74.200 197.535 74.830 197.565 ;
        RECT 70.605 196.715 70.925 197.140 ;
        RECT 71.095 196.545 71.425 196.970 ;
        RECT 71.595 196.965 71.765 197.140 ;
        RECT 71.935 197.135 73.625 197.305 ;
        RECT 73.795 197.140 74.885 197.310 ;
        RECT 75.555 197.285 75.895 198.315 ;
        RECT 76.925 198.125 77.195 198.895 ;
        RECT 78.290 198.660 83.635 199.095 ;
        RECT 83.810 198.660 89.155 199.095 ;
        RECT 76.065 197.955 77.195 198.125 ;
        RECT 76.065 197.455 76.315 197.955 ;
        RECT 73.795 196.965 73.965 197.140 ;
        RECT 71.595 196.715 72.685 196.965 ;
        RECT 72.875 196.715 73.965 196.965 ;
        RECT 74.135 196.545 74.465 196.970 ;
        RECT 74.635 196.715 74.885 197.140 ;
        RECT 75.065 196.545 75.355 197.270 ;
        RECT 75.555 197.115 76.240 197.285 ;
        RECT 76.495 197.205 76.855 197.785 ;
        RECT 75.530 196.545 75.865 196.945 ;
        RECT 76.035 196.715 76.240 197.115 ;
        RECT 77.025 197.045 77.195 197.955 ;
        RECT 79.880 197.410 80.230 198.660 ;
        RECT 81.710 197.090 82.050 197.920 ;
        RECT 85.400 197.410 85.750 198.660 ;
        RECT 89.335 197.955 89.665 199.095 ;
        RECT 90.195 198.125 90.525 198.910 ;
        RECT 90.795 198.475 90.965 198.905 ;
        RECT 91.135 198.645 91.465 199.095 ;
        RECT 90.795 198.245 91.475 198.475 ;
        RECT 89.845 197.955 90.525 198.125 ;
        RECT 87.230 197.090 87.570 197.920 ;
        RECT 89.325 197.535 89.675 197.785 ;
        RECT 89.845 197.355 90.015 197.955 ;
        RECT 90.185 197.535 90.535 197.785 ;
        RECT 90.770 197.735 91.070 198.075 ;
        RECT 90.765 197.565 91.070 197.735 ;
        RECT 76.450 196.545 76.725 197.025 ;
        RECT 76.935 196.715 77.195 197.045 ;
        RECT 78.290 196.545 83.635 197.090 ;
        RECT 83.810 196.545 89.155 197.090 ;
        RECT 89.335 196.545 89.605 197.355 ;
        RECT 89.775 196.715 90.105 197.355 ;
        RECT 90.275 196.545 90.515 197.355 ;
        RECT 90.770 197.225 91.070 197.565 ;
        RECT 91.240 197.595 91.475 198.245 ;
        RECT 91.665 197.935 91.950 198.880 ;
        RECT 92.130 198.625 92.815 199.095 ;
        RECT 92.125 198.105 92.820 198.415 ;
        RECT 92.995 198.040 93.300 198.825 ;
        RECT 93.485 198.140 93.755 199.095 ;
        RECT 93.930 198.705 94.265 198.925 ;
        RECT 95.270 198.715 95.625 199.095 ;
        RECT 91.665 197.785 92.525 197.935 ;
        RECT 91.665 197.765 92.955 197.785 ;
        RECT 91.240 197.265 91.795 197.595 ;
        RECT 91.965 197.405 92.955 197.765 ;
        RECT 91.240 197.115 91.455 197.265 ;
        RECT 90.715 196.545 91.045 197.050 ;
        RECT 91.215 196.740 91.455 197.115 ;
        RECT 91.965 197.070 92.135 197.405 ;
        RECT 93.125 197.235 93.300 198.040 ;
        RECT 93.930 198.085 94.185 198.705 ;
        RECT 94.435 198.545 94.665 198.585 ;
        RECT 95.795 198.545 96.045 198.925 ;
        RECT 94.435 198.345 96.045 198.545 ;
        RECT 94.435 198.255 94.620 198.345 ;
        RECT 95.210 198.335 96.045 198.345 ;
        RECT 96.295 198.315 96.545 199.095 ;
        RECT 96.715 198.245 96.975 198.925 ;
        RECT 97.235 198.755 98.395 198.925 ;
        RECT 97.235 198.255 97.405 198.755 ;
        RECT 94.775 198.145 95.105 198.175 ;
        RECT 94.775 198.085 96.575 198.145 ;
        RECT 93.930 197.975 96.635 198.085 ;
        RECT 93.930 197.915 95.105 197.975 ;
        RECT 96.435 197.940 96.635 197.975 ;
        RECT 93.925 197.535 94.415 197.735 ;
        RECT 94.605 197.535 95.080 197.745 ;
        RECT 91.735 196.875 92.135 197.070 ;
        RECT 91.735 196.730 91.905 196.875 ;
        RECT 92.495 196.545 92.895 197.040 ;
        RECT 93.065 196.715 93.300 197.235 ;
        RECT 93.485 196.545 93.755 197.180 ;
        RECT 93.930 196.545 94.385 197.310 ;
        RECT 94.860 197.135 95.080 197.535 ;
        RECT 95.325 197.535 95.655 197.745 ;
        RECT 95.325 197.135 95.535 197.535 ;
        RECT 95.825 197.500 96.235 197.805 ;
        RECT 96.465 197.365 96.635 197.940 ;
        RECT 96.365 197.245 96.635 197.365 ;
        RECT 95.790 197.200 96.635 197.245 ;
        RECT 95.790 197.075 96.545 197.200 ;
        RECT 95.790 196.925 95.960 197.075 ;
        RECT 96.805 197.055 96.975 198.245 ;
        RECT 97.665 198.125 97.835 198.585 ;
        RECT 98.065 198.505 98.395 198.755 ;
        RECT 98.620 198.675 98.950 199.095 ;
        RECT 99.205 198.505 99.490 198.925 ;
        RECT 98.065 198.335 99.490 198.505 ;
        RECT 99.735 198.295 100.065 199.095 ;
        RECT 100.315 198.375 100.650 198.885 ;
        RECT 97.210 197.785 97.415 198.075 ;
        RECT 97.665 197.955 100.035 198.125 ;
        RECT 99.865 197.785 100.035 197.955 ;
        RECT 97.210 197.735 97.560 197.785 ;
        RECT 97.205 197.565 97.560 197.735 ;
        RECT 97.210 197.455 97.560 197.565 ;
        RECT 96.745 197.045 96.975 197.055 ;
        RECT 94.660 196.715 95.960 196.925 ;
        RECT 96.215 196.545 96.545 196.905 ;
        RECT 96.715 196.715 96.975 197.045 ;
        RECT 97.155 196.545 97.485 197.265 ;
        RECT 97.870 197.120 98.290 197.785 ;
        RECT 98.460 197.395 98.750 197.785 ;
        RECT 98.940 197.395 99.210 197.785 ;
        RECT 99.420 197.735 99.670 197.785 ;
        RECT 99.420 197.565 99.675 197.735 ;
        RECT 99.420 197.455 99.670 197.565 ;
        RECT 99.865 197.455 100.170 197.785 ;
        RECT 98.460 197.225 98.755 197.395 ;
        RECT 98.940 197.225 99.215 197.395 ;
        RECT 99.865 197.285 100.035 197.455 ;
        RECT 98.460 197.125 98.750 197.225 ;
        RECT 98.940 197.125 99.210 197.225 ;
        RECT 99.475 197.115 100.035 197.285 ;
        RECT 99.475 196.945 99.645 197.115 ;
        RECT 100.395 197.020 100.650 198.375 ;
        RECT 100.825 197.930 101.115 199.095 ;
        RECT 102.205 198.335 102.870 198.925 ;
        RECT 102.205 197.365 102.455 198.335 ;
        RECT 103.040 198.255 103.370 199.095 ;
        RECT 103.880 198.505 104.685 198.925 ;
        RECT 103.540 198.335 105.105 198.505 ;
        RECT 103.540 198.085 103.710 198.335 ;
        RECT 102.790 197.915 103.710 198.085 ;
        RECT 102.790 197.745 102.960 197.915 ;
        RECT 103.880 197.745 104.255 198.165 ;
        RECT 102.625 197.535 102.960 197.745 ;
        RECT 103.130 197.535 103.580 197.745 ;
        RECT 103.770 197.735 104.255 197.745 ;
        RECT 104.445 197.785 104.765 198.165 ;
        RECT 104.935 198.085 105.105 198.335 ;
        RECT 105.275 198.255 105.525 199.095 ;
        RECT 105.720 198.085 106.020 198.925 ;
        RECT 104.935 197.915 106.020 198.085 ;
        RECT 107.270 198.145 107.535 198.915 ;
        RECT 107.705 198.375 108.035 199.095 ;
        RECT 108.225 198.555 108.485 198.915 ;
        RECT 108.655 198.725 108.985 199.095 ;
        RECT 109.155 198.555 109.415 198.915 ;
        RECT 108.225 198.325 109.415 198.555 ;
        RECT 109.985 198.145 110.275 198.915 ;
        RECT 103.770 197.565 104.275 197.735 ;
        RECT 103.770 197.535 104.255 197.565 ;
        RECT 104.445 197.535 104.825 197.785 ;
        RECT 105.005 197.535 105.335 197.745 ;
        RECT 98.030 196.775 99.645 196.945 ;
        RECT 99.815 196.545 100.145 196.945 ;
        RECT 100.315 196.760 100.650 197.020 ;
        RECT 100.825 196.545 101.115 197.270 ;
        RECT 102.205 196.725 102.890 197.365 ;
        RECT 103.060 196.545 103.230 197.365 ;
        RECT 103.400 197.195 105.100 197.365 ;
        RECT 103.400 196.730 103.730 197.195 ;
        RECT 104.715 197.105 105.100 197.195 ;
        RECT 105.505 197.285 105.675 197.915 ;
        RECT 105.845 197.455 106.175 197.745 ;
        RECT 105.505 197.105 106.015 197.285 ;
        RECT 103.900 196.545 104.070 197.015 ;
        RECT 104.330 196.765 105.515 196.935 ;
        RECT 105.685 196.715 106.015 197.105 ;
        RECT 107.270 196.725 107.605 198.145 ;
        RECT 107.780 197.965 110.275 198.145 ;
        RECT 107.780 197.275 108.005 197.965 ;
        RECT 108.205 197.455 108.485 197.785 ;
        RECT 108.665 197.455 109.240 197.785 ;
        RECT 109.420 197.455 109.855 197.785 ;
        RECT 110.035 197.455 110.305 197.785 ;
        RECT 107.780 197.085 110.265 197.275 ;
        RECT 107.785 196.545 108.530 196.915 ;
        RECT 109.095 196.725 109.350 197.085 ;
        RECT 109.530 196.545 109.860 196.915 ;
        RECT 110.040 196.725 110.265 197.085 ;
        RECT 110.495 196.725 110.755 198.915 ;
        RECT 110.925 198.365 111.265 199.095 ;
        RECT 111.445 198.185 111.715 198.915 ;
        RECT 110.945 197.965 111.715 198.185 ;
        RECT 111.895 198.205 112.125 198.915 ;
        RECT 112.295 198.385 112.625 199.095 ;
        RECT 112.795 198.205 113.055 198.915 ;
        RECT 111.895 197.965 113.055 198.205 ;
        RECT 113.245 198.005 114.455 199.095 ;
        RECT 114.625 198.005 118.135 199.095 ;
        RECT 118.310 198.660 123.655 199.095 ;
        RECT 123.830 198.670 124.165 199.095 ;
        RECT 110.945 197.295 111.235 197.965 ;
        RECT 111.415 197.475 111.880 197.785 ;
        RECT 112.060 197.475 112.585 197.785 ;
        RECT 110.945 197.095 112.175 197.295 ;
        RECT 111.015 196.545 111.685 196.915 ;
        RECT 111.865 196.725 112.175 197.095 ;
        RECT 112.355 196.835 112.585 197.475 ;
        RECT 112.765 197.455 113.065 197.785 ;
        RECT 113.245 197.465 113.765 198.005 ;
        RECT 113.935 197.295 114.455 197.835 ;
        RECT 114.625 197.485 116.315 198.005 ;
        RECT 116.485 197.315 118.135 197.835 ;
        RECT 119.900 197.410 120.250 198.660 ;
        RECT 124.335 198.490 124.520 198.895 ;
        RECT 123.855 198.315 124.520 198.490 ;
        RECT 124.725 198.315 125.055 199.095 ;
        RECT 112.765 196.545 113.055 197.275 ;
        RECT 113.245 196.545 114.455 197.295 ;
        RECT 114.625 196.545 118.135 197.315 ;
        RECT 121.730 197.090 122.070 197.920 ;
        RECT 123.855 197.285 124.195 198.315 ;
        RECT 125.225 198.125 125.495 198.895 ;
        RECT 124.365 197.955 125.495 198.125 ;
        RECT 124.365 197.455 124.615 197.955 ;
        RECT 123.855 197.115 124.540 197.285 ;
        RECT 124.795 197.205 125.155 197.785 ;
        RECT 118.310 196.545 123.655 197.090 ;
        RECT 123.830 196.545 124.165 196.945 ;
        RECT 124.335 196.715 124.540 197.115 ;
        RECT 125.325 197.045 125.495 197.955 ;
        RECT 125.665 198.005 126.875 199.095 ;
        RECT 125.665 197.465 126.185 198.005 ;
        RECT 126.355 197.295 126.875 197.835 ;
        RECT 124.750 196.545 125.025 197.025 ;
        RECT 125.235 196.715 125.495 197.045 ;
        RECT 125.665 196.545 126.875 197.295 ;
        RECT 14.260 196.375 126.960 196.545 ;
        RECT 14.345 195.625 15.555 196.375 ;
        RECT 15.815 195.895 16.115 196.375 ;
        RECT 16.285 195.725 16.545 196.180 ;
        RECT 16.715 195.895 16.975 196.375 ;
        RECT 17.155 195.725 17.415 196.180 ;
        RECT 17.585 195.895 17.835 196.375 ;
        RECT 18.015 195.725 18.275 196.180 ;
        RECT 18.445 195.895 18.695 196.375 ;
        RECT 18.875 195.725 19.135 196.180 ;
        RECT 19.305 195.895 19.550 196.375 ;
        RECT 19.720 195.725 19.995 196.180 ;
        RECT 20.165 195.895 20.410 196.375 ;
        RECT 20.580 195.725 20.840 196.180 ;
        RECT 21.010 195.895 21.270 196.375 ;
        RECT 21.440 195.725 21.700 196.180 ;
        RECT 21.870 195.895 22.130 196.375 ;
        RECT 22.300 195.725 22.560 196.180 ;
        RECT 22.730 195.815 22.990 196.375 ;
        RECT 14.345 195.085 14.865 195.625 ;
        RECT 15.815 195.555 22.560 195.725 ;
        RECT 15.035 194.915 15.555 195.455 ;
        RECT 14.345 193.825 15.555 194.915 ;
        RECT 15.815 194.965 16.980 195.555 ;
        RECT 23.160 195.385 23.410 196.195 ;
        RECT 23.590 195.850 23.850 196.375 ;
        RECT 24.020 195.385 24.270 196.195 ;
        RECT 24.450 195.865 24.755 196.375 ;
        RECT 17.150 195.135 24.270 195.385 ;
        RECT 24.440 195.135 24.755 195.695 ;
        RECT 24.965 195.555 25.195 196.375 ;
        RECT 25.365 195.575 25.695 196.205 ;
        RECT 24.945 195.135 25.275 195.385 ;
        RECT 15.815 194.740 22.560 194.965 ;
        RECT 15.815 193.825 16.085 194.570 ;
        RECT 16.255 194.000 16.545 194.740 ;
        RECT 17.155 194.725 22.560 194.740 ;
        RECT 16.715 193.830 16.970 194.555 ;
        RECT 17.155 194.000 17.415 194.725 ;
        RECT 17.585 193.830 17.830 194.555 ;
        RECT 18.015 194.000 18.275 194.725 ;
        RECT 18.445 193.830 18.690 194.555 ;
        RECT 18.875 194.000 19.135 194.725 ;
        RECT 19.305 193.830 19.550 194.555 ;
        RECT 19.720 194.000 19.980 194.725 ;
        RECT 20.150 193.830 20.410 194.555 ;
        RECT 20.580 194.000 20.840 194.725 ;
        RECT 21.010 193.830 21.270 194.555 ;
        RECT 21.440 194.000 21.700 194.725 ;
        RECT 21.870 193.830 22.130 194.555 ;
        RECT 22.300 194.000 22.560 194.725 ;
        RECT 22.730 193.830 22.990 194.625 ;
        RECT 23.160 194.000 23.410 195.135 ;
        RECT 16.715 193.825 22.990 193.830 ;
        RECT 23.590 193.825 23.850 194.635 ;
        RECT 24.025 193.995 24.270 195.135 ;
        RECT 25.445 194.975 25.695 195.575 ;
        RECT 25.865 195.555 26.075 196.375 ;
        RECT 27.315 195.895 27.615 196.375 ;
        RECT 27.785 195.725 28.045 196.180 ;
        RECT 28.215 195.895 28.475 196.375 ;
        RECT 28.655 195.725 28.915 196.180 ;
        RECT 29.085 195.895 29.335 196.375 ;
        RECT 29.515 195.725 29.775 196.180 ;
        RECT 29.945 195.895 30.195 196.375 ;
        RECT 30.375 195.725 30.635 196.180 ;
        RECT 30.805 195.895 31.050 196.375 ;
        RECT 31.220 195.725 31.495 196.180 ;
        RECT 31.665 195.895 31.910 196.375 ;
        RECT 32.080 195.725 32.340 196.180 ;
        RECT 32.510 195.895 32.770 196.375 ;
        RECT 32.940 195.725 33.200 196.180 ;
        RECT 33.370 195.895 33.630 196.375 ;
        RECT 33.800 195.725 34.060 196.180 ;
        RECT 34.230 195.815 34.490 196.375 ;
        RECT 27.315 195.555 34.060 195.725 ;
        RECT 24.450 193.825 24.745 194.635 ;
        RECT 24.965 193.825 25.195 194.965 ;
        RECT 25.365 193.995 25.695 194.975 ;
        RECT 27.315 194.965 28.480 195.555 ;
        RECT 34.660 195.385 34.910 196.195 ;
        RECT 35.090 195.850 35.350 196.375 ;
        RECT 35.520 195.385 35.770 196.195 ;
        RECT 35.950 195.865 36.255 196.375 ;
        RECT 28.650 195.135 35.770 195.385 ;
        RECT 35.940 195.135 36.255 195.695 ;
        RECT 36.425 195.650 36.715 196.375 ;
        RECT 36.945 195.555 37.155 196.375 ;
        RECT 37.325 195.575 37.655 196.205 ;
        RECT 25.865 193.825 26.075 194.965 ;
        RECT 27.315 194.740 34.060 194.965 ;
        RECT 27.315 193.825 27.585 194.570 ;
        RECT 27.755 194.000 28.045 194.740 ;
        RECT 28.655 194.725 34.060 194.740 ;
        RECT 28.215 193.830 28.470 194.555 ;
        RECT 28.655 194.000 28.915 194.725 ;
        RECT 29.085 193.830 29.330 194.555 ;
        RECT 29.515 194.000 29.775 194.725 ;
        RECT 29.945 193.830 30.190 194.555 ;
        RECT 30.375 194.000 30.635 194.725 ;
        RECT 30.805 193.830 31.050 194.555 ;
        RECT 31.220 194.000 31.480 194.725 ;
        RECT 31.650 193.830 31.910 194.555 ;
        RECT 32.080 194.000 32.340 194.725 ;
        RECT 32.510 193.830 32.770 194.555 ;
        RECT 32.940 194.000 33.200 194.725 ;
        RECT 33.370 193.830 33.630 194.555 ;
        RECT 33.800 194.000 34.060 194.725 ;
        RECT 34.230 193.830 34.490 194.625 ;
        RECT 34.660 194.000 34.910 195.135 ;
        RECT 28.215 193.825 34.490 193.830 ;
        RECT 35.090 193.825 35.350 194.635 ;
        RECT 35.525 193.995 35.770 195.135 ;
        RECT 35.950 193.825 36.245 194.635 ;
        RECT 36.425 193.825 36.715 194.990 ;
        RECT 37.325 194.975 37.575 195.575 ;
        RECT 37.825 195.555 38.055 196.375 ;
        RECT 38.795 195.905 38.965 196.375 ;
        RECT 39.135 195.735 39.465 196.185 ;
        RECT 39.635 195.905 39.805 196.375 ;
        RECT 39.975 195.735 40.305 196.185 ;
        RECT 38.630 195.555 40.305 195.735 ;
        RECT 40.475 195.565 40.645 196.375 ;
        RECT 40.815 195.985 41.985 196.155 ;
        RECT 40.815 195.565 41.065 195.985 ;
        RECT 42.155 195.905 42.325 196.375 ;
        RECT 42.595 195.985 43.765 196.205 ;
        RECT 41.235 195.735 41.565 195.815 ;
        RECT 41.235 195.555 42.585 195.735 ;
        RECT 43.015 195.645 43.345 195.815 ;
        RECT 37.745 195.135 38.075 195.385 ;
        RECT 38.630 195.045 38.935 195.555 ;
        RECT 42.395 195.385 42.585 195.555 ;
        RECT 43.095 195.385 43.345 195.645 ;
        RECT 43.515 195.725 43.765 195.985 ;
        RECT 43.935 195.905 44.105 196.375 ;
        RECT 44.275 195.735 44.605 196.205 ;
        RECT 44.775 195.905 44.945 196.375 ;
        RECT 45.115 195.735 45.445 196.205 ;
        RECT 44.275 195.725 45.445 195.735 ;
        RECT 43.515 195.555 45.445 195.725 ;
        RECT 46.750 195.595 47.250 196.205 ;
        RECT 39.105 195.215 40.375 195.385 ;
        RECT 36.945 193.825 37.155 194.965 ;
        RECT 37.325 193.995 37.655 194.975 ;
        RECT 37.825 193.825 38.055 194.965 ;
        RECT 38.630 194.805 39.425 195.045 ;
        RECT 40.085 194.845 40.375 195.215 ;
        RECT 40.575 195.015 40.935 195.385 ;
        RECT 41.105 195.185 41.725 195.385 ;
        RECT 41.895 195.015 42.225 195.385 ;
        RECT 40.575 194.845 42.225 195.015 ;
        RECT 42.395 195.215 42.925 195.385 ;
        RECT 39.175 194.675 39.425 194.805 ;
        RECT 42.395 194.675 42.585 195.215 ;
        RECT 43.095 195.045 43.475 195.385 ;
        RECT 38.755 193.825 39.005 194.635 ;
        RECT 39.175 194.505 40.265 194.675 ;
        RECT 39.175 193.995 39.425 194.505 ;
        RECT 39.595 193.825 39.845 194.295 ;
        RECT 40.015 193.995 40.265 194.505 ;
        RECT 40.435 193.825 40.685 194.665 ;
        RECT 40.855 194.495 42.585 194.675 ;
        RECT 42.925 194.675 43.475 195.045 ;
        RECT 43.645 195.015 43.975 195.385 ;
        RECT 44.195 195.185 44.735 195.385 ;
        RECT 44.965 195.015 45.455 195.385 ;
        RECT 46.545 195.135 46.895 195.385 ;
        RECT 43.645 194.845 45.455 195.015 ;
        RECT 47.080 194.965 47.250 195.595 ;
        RECT 47.880 195.725 48.210 196.205 ;
        RECT 48.380 195.915 48.605 196.375 ;
        RECT 48.775 195.725 49.105 196.205 ;
        RECT 47.880 195.555 49.105 195.725 ;
        RECT 49.295 195.575 49.545 196.375 ;
        RECT 49.715 195.575 50.055 196.205 ;
        RECT 50.250 195.985 50.580 196.375 ;
        RECT 50.750 195.815 50.975 196.195 ;
        RECT 47.420 195.185 47.750 195.385 ;
        RECT 47.920 195.185 48.250 195.385 ;
        RECT 48.420 195.185 48.840 195.385 ;
        RECT 49.015 195.215 49.710 195.385 ;
        RECT 49.015 194.965 49.185 195.215 ;
        RECT 49.880 194.965 50.055 195.575 ;
        RECT 50.235 195.135 50.475 195.785 ;
        RECT 50.645 195.635 50.975 195.815 ;
        RECT 50.645 194.965 50.820 195.635 ;
        RECT 51.175 195.465 51.405 196.085 ;
        RECT 51.585 195.645 51.885 196.375 ;
        RECT 52.565 195.865 52.965 196.375 ;
        RECT 53.540 195.760 53.710 196.205 ;
        RECT 53.880 195.975 54.600 196.375 ;
        RECT 54.770 195.805 54.940 196.205 ;
        RECT 55.175 195.930 55.605 196.375 ;
        RECT 50.990 195.135 51.405 195.465 ;
        RECT 51.585 195.135 51.880 195.465 ;
        RECT 46.750 194.795 49.185 194.965 ;
        RECT 42.925 194.505 44.565 194.675 ;
        RECT 42.925 194.495 43.305 194.505 ;
        RECT 40.855 193.995 41.105 194.495 ;
        RECT 41.695 194.335 41.945 194.495 ;
        RECT 41.275 193.825 41.525 194.325 ;
        RECT 42.115 193.825 42.845 194.325 ;
        RECT 43.015 193.995 43.305 194.495 ;
        RECT 44.315 194.335 44.565 194.505 ;
        RECT 43.475 193.825 43.725 194.335 ;
        RECT 43.895 194.165 44.145 194.335 ;
        RECT 44.735 194.165 44.985 194.675 ;
        RECT 43.895 193.995 44.985 194.165 ;
        RECT 45.195 193.825 45.400 194.665 ;
        RECT 46.750 193.995 47.080 194.795 ;
        RECT 47.250 193.825 47.580 194.625 ;
        RECT 47.880 193.995 48.210 194.795 ;
        RECT 48.855 193.825 49.105 194.625 ;
        RECT 49.375 193.825 49.545 194.965 ;
        RECT 49.715 193.995 50.055 194.965 ;
        RECT 50.235 194.775 50.820 194.965 ;
        RECT 50.235 194.005 50.510 194.775 ;
        RECT 50.990 194.605 51.885 194.935 ;
        RECT 52.580 194.805 52.840 195.695 ;
        RECT 53.040 195.105 53.300 195.695 ;
        RECT 53.540 195.590 53.890 195.760 ;
        RECT 53.040 194.805 53.520 195.105 ;
        RECT 50.680 194.435 51.885 194.605 ;
        RECT 50.680 194.005 51.010 194.435 ;
        RECT 51.180 193.825 51.375 194.265 ;
        RECT 51.555 194.005 51.885 194.435 ;
        RECT 52.605 194.455 53.545 194.625 ;
        RECT 52.605 193.995 52.785 194.455 ;
        RECT 52.955 193.825 53.205 194.285 ;
        RECT 53.375 194.205 53.545 194.455 ;
        RECT 53.720 194.565 53.890 195.590 ;
        RECT 54.060 195.635 54.940 195.805 ;
        RECT 55.775 195.650 56.035 196.205 ;
        RECT 54.060 194.915 54.230 195.635 ;
        RECT 54.420 195.085 54.710 195.465 ;
        RECT 54.060 194.745 54.580 194.915 ;
        RECT 54.880 194.845 55.210 195.465 ;
        RECT 55.435 195.135 55.690 195.465 ;
        RECT 53.720 194.395 54.130 194.565 ;
        RECT 54.410 194.555 54.580 194.745 ;
        RECT 55.435 194.655 55.605 195.135 ;
        RECT 55.860 194.935 56.035 195.650 ;
        RECT 56.210 195.610 56.665 196.375 ;
        RECT 56.940 195.995 58.240 196.205 ;
        RECT 58.495 196.015 58.825 196.375 ;
        RECT 58.070 195.845 58.240 195.995 ;
        RECT 58.995 195.875 59.255 196.205 ;
        RECT 57.140 195.385 57.360 195.785 ;
        RECT 56.205 195.185 56.695 195.385 ;
        RECT 56.885 195.175 57.360 195.385 ;
        RECT 57.605 195.385 57.815 195.785 ;
        RECT 58.070 195.720 58.825 195.845 ;
        RECT 58.070 195.675 58.915 195.720 ;
        RECT 58.645 195.555 58.915 195.675 ;
        RECT 57.605 195.175 57.935 195.385 ;
        RECT 58.105 195.115 58.515 195.420 ;
        RECT 53.875 194.260 54.130 194.395 ;
        RECT 54.845 194.485 55.605 194.655 ;
        RECT 54.845 194.260 55.015 194.485 ;
        RECT 53.375 194.035 53.705 194.205 ;
        RECT 53.875 194.090 55.015 194.260 ;
        RECT 53.875 193.995 54.130 194.090 ;
        RECT 55.275 193.825 55.605 194.225 ;
        RECT 55.775 193.995 56.035 194.935 ;
        RECT 56.210 194.945 57.385 195.005 ;
        RECT 58.745 194.980 58.915 195.555 ;
        RECT 58.715 194.945 58.915 194.980 ;
        RECT 56.210 194.835 58.915 194.945 ;
        RECT 56.210 194.215 56.465 194.835 ;
        RECT 57.055 194.775 58.855 194.835 ;
        RECT 57.055 194.745 57.385 194.775 ;
        RECT 59.085 194.675 59.255 195.875 ;
        RECT 59.435 195.865 59.885 196.375 ;
        RECT 60.160 195.955 61.465 196.205 ;
        RECT 61.645 195.975 61.975 196.375 ;
        RECT 61.285 195.805 61.465 195.955 ;
        RECT 59.465 195.185 59.915 195.695 ;
        RECT 60.330 195.385 60.580 195.785 ;
        RECT 60.105 195.185 60.580 195.385 ;
        RECT 60.830 195.385 61.040 195.785 ;
        RECT 61.285 195.635 62.015 195.805 ;
        RECT 62.185 195.650 62.475 196.375 ;
        RECT 62.645 195.700 62.915 196.045 ;
        RECT 63.105 195.975 63.485 196.375 ;
        RECT 63.655 195.805 63.825 196.155 ;
        RECT 63.995 195.975 64.325 196.375 ;
        RECT 64.525 195.805 64.695 196.155 ;
        RECT 64.895 195.875 65.225 196.375 ;
        RECT 60.830 195.185 61.180 195.385 ;
        RECT 61.350 195.135 61.675 195.465 ;
        RECT 56.715 194.575 56.900 194.665 ;
        RECT 57.490 194.575 58.325 194.585 ;
        RECT 56.715 194.375 58.325 194.575 ;
        RECT 56.715 194.335 56.945 194.375 ;
        RECT 56.210 193.995 56.545 194.215 ;
        RECT 57.550 193.825 57.905 194.205 ;
        RECT 58.075 193.995 58.325 194.375 ;
        RECT 58.575 193.825 58.825 194.605 ;
        RECT 58.995 193.995 59.255 194.675 ;
        RECT 59.435 194.965 61.180 195.015 ;
        RECT 61.845 194.965 62.015 195.635 ;
        RECT 59.435 194.835 62.015 194.965 ;
        RECT 59.435 194.165 59.765 194.835 ;
        RECT 60.955 194.795 62.015 194.835 ;
        RECT 59.935 194.625 60.815 194.665 ;
        RECT 59.935 194.425 61.465 194.625 ;
        RECT 59.935 194.375 60.550 194.425 ;
        RECT 59.935 194.335 60.165 194.375 ;
        RECT 61.295 194.295 61.465 194.425 ;
        RECT 60.275 194.165 60.605 194.205 ;
        RECT 59.435 193.995 60.605 194.165 ;
        RECT 60.775 193.825 61.150 194.205 ;
        RECT 61.700 193.825 61.965 194.605 ;
        RECT 62.185 193.825 62.475 194.990 ;
        RECT 62.645 194.965 62.815 195.700 ;
        RECT 63.085 195.635 64.695 195.805 ;
        RECT 63.085 195.465 63.255 195.635 ;
        RECT 62.985 195.135 63.255 195.465 ;
        RECT 63.425 195.135 63.830 195.465 ;
        RECT 63.085 194.965 63.255 195.135 ;
        RECT 62.645 193.995 62.915 194.965 ;
        RECT 63.085 194.795 63.810 194.965 ;
        RECT 64.000 194.845 64.710 195.465 ;
        RECT 64.880 195.135 65.230 195.705 ;
        RECT 63.640 194.675 63.810 194.795 ;
        RECT 64.910 194.675 65.230 194.965 ;
        RECT 63.125 193.825 63.405 194.625 ;
        RECT 63.640 194.505 65.230 194.675 ;
        RECT 63.575 194.045 65.230 194.335 ;
        RECT 65.865 193.995 66.615 196.205 ;
        RECT 66.810 195.985 67.140 196.375 ;
        RECT 67.310 195.815 67.535 196.195 ;
        RECT 66.795 195.135 67.035 195.785 ;
        RECT 67.205 195.635 67.535 195.815 ;
        RECT 67.205 194.965 67.380 195.635 ;
        RECT 67.735 195.465 67.965 196.085 ;
        RECT 68.145 195.645 68.445 196.375 ;
        RECT 69.095 195.645 69.395 196.375 ;
        RECT 69.575 195.465 69.805 196.085 ;
        RECT 70.005 195.815 70.230 196.195 ;
        RECT 70.400 195.985 70.730 196.375 ;
        RECT 70.005 195.635 70.335 195.815 ;
        RECT 67.550 195.135 67.965 195.465 ;
        RECT 68.145 195.135 68.440 195.465 ;
        RECT 69.100 195.135 69.395 195.465 ;
        RECT 69.575 195.135 69.990 195.465 ;
        RECT 66.795 194.775 67.380 194.965 ;
        RECT 70.160 194.965 70.335 195.635 ;
        RECT 70.505 195.135 70.745 195.785 ;
        RECT 71.845 195.605 75.355 196.375 ;
        RECT 66.795 194.005 67.070 194.775 ;
        RECT 67.550 194.605 68.445 194.935 ;
        RECT 67.240 194.435 68.445 194.605 ;
        RECT 67.240 194.005 67.570 194.435 ;
        RECT 67.740 193.825 67.935 194.265 ;
        RECT 68.115 194.005 68.445 194.435 ;
        RECT 69.095 194.605 69.990 194.935 ;
        RECT 70.160 194.775 70.745 194.965 ;
        RECT 69.095 194.435 70.300 194.605 ;
        RECT 69.095 194.005 69.425 194.435 ;
        RECT 69.605 193.825 69.800 194.265 ;
        RECT 69.970 194.005 70.300 194.435 ;
        RECT 70.470 194.005 70.745 194.775 ;
        RECT 71.845 194.915 73.535 195.435 ;
        RECT 73.705 195.085 75.355 195.605 ;
        RECT 75.560 195.635 76.175 196.205 ;
        RECT 76.345 195.865 76.560 196.375 ;
        RECT 76.790 195.865 77.070 196.195 ;
        RECT 77.250 195.865 77.490 196.375 ;
        RECT 71.845 193.825 75.355 194.915 ;
        RECT 75.560 194.615 75.875 195.635 ;
        RECT 76.045 194.965 76.215 195.465 ;
        RECT 76.465 195.135 76.730 195.695 ;
        RECT 76.900 194.965 77.070 195.865 ;
        RECT 77.240 195.135 77.595 195.695 ;
        RECT 78.265 195.655 78.605 196.375 ;
        RECT 78.795 195.465 78.995 196.045 ;
        RECT 79.255 195.695 79.555 196.115 ;
        RECT 78.210 195.135 78.625 195.445 ;
        RECT 78.795 195.135 79.155 195.465 ;
        RECT 79.365 195.385 79.555 195.695 ;
        RECT 79.795 195.825 80.045 196.165 ;
        RECT 80.535 195.995 80.865 196.375 ;
        RECT 79.795 195.655 80.445 195.825 ;
        RECT 79.365 195.205 79.730 195.385 ;
        RECT 79.935 195.035 80.105 195.465 ;
        RECT 76.045 194.795 77.470 194.965 ;
        RECT 75.560 193.995 76.095 194.615 ;
        RECT 76.265 193.825 76.595 194.625 ;
        RECT 77.080 194.620 77.470 194.795 ;
        RECT 78.265 193.825 78.605 194.965 ;
        RECT 79.705 194.845 80.105 195.035 ;
        RECT 78.775 194.675 78.945 194.715 ;
        RECT 80.275 194.675 80.445 195.655 ;
        RECT 81.250 195.595 81.750 196.205 ;
        RECT 80.615 195.135 80.875 195.465 ;
        RECT 81.045 195.135 81.395 195.385 ;
        RECT 81.580 194.965 81.750 195.595 ;
        RECT 82.380 195.725 82.710 196.205 ;
        RECT 82.880 195.915 83.105 196.375 ;
        RECT 83.275 195.725 83.605 196.205 ;
        RECT 82.380 195.555 83.605 195.725 ;
        RECT 83.795 195.575 84.045 196.375 ;
        RECT 84.215 195.575 84.555 196.205 ;
        RECT 85.185 195.605 87.775 196.375 ;
        RECT 87.945 195.650 88.235 196.375 ;
        RECT 88.405 195.625 89.615 196.375 ;
        RECT 81.920 195.185 82.250 195.385 ;
        RECT 82.420 195.185 82.750 195.385 ;
        RECT 82.920 195.185 83.340 195.385 ;
        RECT 83.515 195.215 84.210 195.385 ;
        RECT 83.515 194.965 83.685 195.215 ;
        RECT 84.380 194.965 84.555 195.575 ;
        RECT 78.775 194.505 79.865 194.675 ;
        RECT 78.775 193.995 78.945 194.505 ;
        RECT 79.155 193.825 79.405 194.325 ;
        RECT 79.615 194.205 79.865 194.505 ;
        RECT 80.095 194.375 80.445 194.675 ;
        RECT 81.250 194.795 83.685 194.965 ;
        RECT 80.615 194.205 80.875 194.625 ;
        RECT 79.615 193.995 80.875 194.205 ;
        RECT 81.250 193.995 81.580 194.795 ;
        RECT 81.750 193.825 82.080 194.625 ;
        RECT 82.380 193.995 82.710 194.795 ;
        RECT 83.355 193.825 83.605 194.625 ;
        RECT 83.875 193.825 84.045 194.965 ;
        RECT 84.215 193.995 84.555 194.965 ;
        RECT 85.185 194.915 86.395 195.435 ;
        RECT 86.565 195.085 87.775 195.605 ;
        RECT 85.185 193.825 87.775 194.915 ;
        RECT 87.945 193.825 88.235 194.990 ;
        RECT 88.405 194.915 88.925 195.455 ;
        RECT 89.095 195.085 89.615 195.625 ;
        RECT 89.785 195.575 90.480 196.205 ;
        RECT 90.685 195.575 90.995 196.375 ;
        RECT 91.625 195.765 91.975 196.205 ;
        RECT 92.145 195.935 92.315 196.375 ;
        RECT 92.485 195.995 93.680 196.205 ;
        RECT 92.485 195.765 92.735 195.995 ;
        RECT 89.805 195.135 90.140 195.385 ;
        RECT 90.310 194.975 90.480 195.575 ;
        RECT 91.625 195.555 92.735 195.765 ;
        RECT 92.905 195.655 93.235 195.825 ;
        RECT 92.905 195.555 93.230 195.655 ;
        RECT 93.405 195.555 93.680 195.995 ;
        RECT 93.915 195.635 94.245 196.375 ;
        RECT 94.415 195.620 94.650 195.950 ;
        RECT 90.650 195.135 90.985 195.405 ;
        RECT 91.625 195.355 92.770 195.385 ;
        RECT 91.625 195.185 92.775 195.355 ;
        RECT 88.405 193.825 89.615 194.915 ;
        RECT 89.785 193.825 90.045 194.965 ;
        RECT 90.215 193.995 90.545 194.975 ;
        RECT 90.715 193.825 90.995 194.965 ;
        RECT 91.625 193.825 91.955 194.965 ;
        RECT 92.125 194.625 92.400 194.965 ;
        RECT 92.580 194.805 92.770 195.185 ;
        RECT 92.950 194.625 93.230 195.555 ;
        RECT 93.400 194.965 93.730 195.385 ;
        RECT 93.960 195.135 94.305 195.465 ;
        RECT 94.480 194.965 94.650 195.620 ;
        RECT 95.305 195.605 96.975 196.375 ;
        RECT 97.150 195.830 102.495 196.375 ;
        RECT 93.400 194.795 94.650 194.965 ;
        RECT 92.125 194.455 93.725 194.625 ;
        RECT 92.125 193.995 92.480 194.455 ;
        RECT 92.650 193.825 93.225 194.285 ;
        RECT 93.395 193.995 93.725 194.455 ;
        RECT 93.925 193.825 94.180 194.625 ;
        RECT 94.350 194.600 94.650 194.795 ;
        RECT 95.305 194.915 96.055 195.435 ;
        RECT 96.225 195.085 96.975 195.605 ;
        RECT 95.305 193.825 96.975 194.915 ;
        RECT 98.740 194.260 99.090 195.510 ;
        RECT 100.570 195.000 100.910 195.830 ;
        RECT 102.700 195.635 103.315 196.205 ;
        RECT 103.485 195.865 103.700 196.375 ;
        RECT 103.930 195.865 104.210 196.195 ;
        RECT 104.390 195.865 104.630 196.375 ;
        RECT 102.700 194.615 103.015 195.635 ;
        RECT 103.185 194.965 103.355 195.465 ;
        RECT 103.605 195.135 103.870 195.695 ;
        RECT 104.040 194.965 104.210 195.865 ;
        RECT 104.380 195.135 104.735 195.695 ;
        RECT 104.970 195.535 105.230 196.375 ;
        RECT 105.405 195.630 105.660 196.205 ;
        RECT 105.830 195.995 106.160 196.375 ;
        RECT 106.375 195.825 106.545 196.205 ;
        RECT 105.830 195.655 106.545 195.825 ;
        RECT 106.805 195.745 107.145 196.205 ;
        RECT 107.315 195.915 107.485 196.375 ;
        RECT 108.115 195.940 108.475 196.205 ;
        RECT 108.120 195.935 108.475 195.940 ;
        RECT 108.125 195.925 108.475 195.935 ;
        RECT 108.130 195.920 108.475 195.925 ;
        RECT 108.135 195.910 108.475 195.920 ;
        RECT 108.715 195.915 108.885 196.375 ;
        RECT 108.140 195.905 108.475 195.910 ;
        RECT 108.150 195.895 108.475 195.905 ;
        RECT 108.160 195.885 108.475 195.895 ;
        RECT 107.655 195.745 107.985 195.825 ;
        RECT 103.185 194.795 104.610 194.965 ;
        RECT 97.150 193.825 102.495 194.260 ;
        RECT 102.700 193.995 103.235 194.615 ;
        RECT 103.405 193.825 103.735 194.625 ;
        RECT 104.220 194.620 104.610 194.795 ;
        RECT 104.970 193.825 105.230 194.975 ;
        RECT 105.405 194.900 105.575 195.630 ;
        RECT 105.830 195.465 106.000 195.655 ;
        RECT 106.805 195.555 107.985 195.745 ;
        RECT 108.175 195.745 108.475 195.885 ;
        RECT 108.175 195.555 108.885 195.745 ;
        RECT 105.745 195.135 106.000 195.465 ;
        RECT 105.830 194.925 106.000 195.135 ;
        RECT 106.280 195.105 106.635 195.475 ;
        RECT 106.805 195.185 107.135 195.385 ;
        RECT 107.445 195.365 107.775 195.385 ;
        RECT 107.325 195.185 107.775 195.365 ;
        RECT 105.405 193.995 105.660 194.900 ;
        RECT 105.830 194.755 106.545 194.925 ;
        RECT 106.805 194.845 107.035 195.185 ;
        RECT 105.830 193.825 106.160 194.585 ;
        RECT 106.375 193.995 106.545 194.755 ;
        RECT 106.815 193.825 107.145 194.545 ;
        RECT 107.325 194.070 107.540 195.185 ;
        RECT 107.945 195.155 108.415 195.385 ;
        RECT 108.600 194.985 108.885 195.555 ;
        RECT 109.055 195.430 109.395 196.205 ;
        RECT 107.735 194.770 108.885 194.985 ;
        RECT 107.735 193.995 108.065 194.770 ;
        RECT 108.235 193.825 108.945 194.600 ;
        RECT 109.115 193.995 109.395 195.430 ;
        RECT 109.565 195.915 110.125 196.205 ;
        RECT 110.295 195.915 110.545 196.375 ;
        RECT 109.565 194.545 109.815 195.915 ;
        RECT 111.165 195.745 111.495 196.105 ;
        RECT 110.105 195.555 111.495 195.745 ;
        RECT 111.865 195.605 113.535 196.375 ;
        RECT 113.705 195.650 113.995 196.375 ;
        RECT 114.165 195.605 115.835 196.375 ;
        RECT 116.010 195.830 121.355 196.375 ;
        RECT 110.105 195.465 110.275 195.555 ;
        RECT 109.985 195.135 110.275 195.465 ;
        RECT 110.445 195.135 110.785 195.385 ;
        RECT 111.005 195.135 111.680 195.385 ;
        RECT 110.105 194.885 110.275 195.135 ;
        RECT 110.105 194.715 111.045 194.885 ;
        RECT 111.415 194.775 111.680 195.135 ;
        RECT 111.865 194.915 112.615 195.435 ;
        RECT 112.785 195.085 113.535 195.605 ;
        RECT 109.565 193.995 110.025 194.545 ;
        RECT 110.215 193.825 110.545 194.545 ;
        RECT 110.745 194.165 111.045 194.715 ;
        RECT 111.215 193.825 111.495 194.495 ;
        RECT 111.865 193.825 113.535 194.915 ;
        RECT 113.705 193.825 113.995 194.990 ;
        RECT 114.165 194.915 114.915 195.435 ;
        RECT 115.085 195.085 115.835 195.605 ;
        RECT 114.165 193.825 115.835 194.915 ;
        RECT 117.600 194.260 117.950 195.510 ;
        RECT 119.430 195.000 119.770 195.830 ;
        RECT 121.615 195.825 121.785 196.205 ;
        RECT 121.965 195.995 122.295 196.375 ;
        RECT 121.615 195.655 122.280 195.825 ;
        RECT 122.475 195.700 122.735 196.205 ;
        RECT 121.545 195.105 121.875 195.475 ;
        RECT 122.110 195.400 122.280 195.655 ;
        RECT 122.110 195.070 122.395 195.400 ;
        RECT 122.110 194.925 122.280 195.070 ;
        RECT 121.615 194.755 122.280 194.925 ;
        RECT 122.565 194.900 122.735 195.700 ;
        RECT 123.915 195.825 124.085 196.205 ;
        RECT 124.300 195.995 124.630 196.375 ;
        RECT 123.915 195.655 124.630 195.825 ;
        RECT 123.825 195.105 124.180 195.475 ;
        RECT 124.460 195.465 124.630 195.655 ;
        RECT 124.800 195.630 125.055 196.205 ;
        RECT 124.460 195.135 124.715 195.465 ;
        RECT 124.460 194.925 124.630 195.135 ;
        RECT 116.010 193.825 121.355 194.260 ;
        RECT 121.615 193.995 121.785 194.755 ;
        RECT 121.965 193.825 122.295 194.585 ;
        RECT 122.465 193.995 122.735 194.900 ;
        RECT 123.915 194.755 124.630 194.925 ;
        RECT 124.885 194.900 125.055 195.630 ;
        RECT 125.230 195.535 125.490 196.375 ;
        RECT 125.665 195.625 126.875 196.375 ;
        RECT 123.915 193.995 124.085 194.755 ;
        RECT 124.300 193.825 124.630 194.585 ;
        RECT 124.800 193.995 125.055 194.900 ;
        RECT 125.230 193.825 125.490 194.975 ;
        RECT 125.665 194.915 126.185 195.455 ;
        RECT 126.355 195.085 126.875 195.625 ;
        RECT 125.665 193.825 126.875 194.915 ;
        RECT 14.260 193.655 126.960 193.825 ;
        RECT 14.345 192.565 15.555 193.655 ;
        RECT 14.345 191.855 14.865 192.395 ;
        RECT 15.035 192.025 15.555 192.565 ;
        RECT 15.730 192.510 16.025 193.655 ;
        RECT 14.345 191.105 15.555 191.855 ;
        RECT 15.730 191.105 16.025 191.925 ;
        RECT 16.195 191.655 16.425 193.355 ;
        RECT 16.640 192.850 16.895 193.655 ;
        RECT 17.095 193.040 17.425 193.485 ;
        RECT 17.595 193.210 17.870 193.655 ;
        RECT 18.105 193.040 18.435 193.485 ;
        RECT 17.095 192.860 18.435 193.040 ;
        RECT 18.895 192.680 19.225 193.345 ;
        RECT 16.640 192.510 19.225 192.680 ;
        RECT 16.640 191.895 16.950 192.510 ;
        RECT 19.505 192.465 19.675 193.655 ;
        RECT 19.845 192.545 20.100 193.485 ;
        RECT 20.270 193.255 20.600 193.655 ;
        RECT 21.820 193.390 21.990 193.485 ;
        RECT 20.860 193.220 21.990 193.390 ;
        RECT 22.195 193.275 22.525 193.445 ;
        RECT 20.860 192.995 21.030 193.220 ;
        RECT 20.270 192.825 21.030 192.995 ;
        RECT 21.760 193.085 21.990 193.220 ;
        RECT 17.120 192.065 17.450 192.295 ;
        RECT 17.620 192.065 18.090 192.295 ;
        RECT 18.260 192.125 18.715 192.295 ;
        RECT 18.260 192.065 18.710 192.125 ;
        RECT 18.900 192.065 19.235 192.295 ;
        RECT 16.640 191.715 19.225 191.895 ;
        RECT 16.195 191.275 16.415 191.655 ;
        RECT 16.585 191.105 17.435 191.465 ;
        RECT 17.915 191.295 18.245 191.715 ;
        RECT 18.450 191.105 18.725 191.545 ;
        RECT 18.895 191.295 19.225 191.715 ;
        RECT 19.505 191.105 19.675 191.950 ;
        RECT 19.845 191.830 20.015 192.545 ;
        RECT 20.270 192.345 20.440 192.825 ;
        RECT 21.295 192.735 21.465 192.925 ;
        RECT 21.760 192.915 22.170 193.085 ;
        RECT 20.185 192.015 20.440 192.345 ;
        RECT 20.665 192.015 20.995 192.635 ;
        RECT 21.295 192.565 21.830 192.735 ;
        RECT 21.165 192.295 21.455 192.395 ;
        RECT 21.165 192.125 21.475 192.295 ;
        RECT 21.165 192.015 21.455 192.125 ;
        RECT 21.660 191.845 21.830 192.565 ;
        RECT 19.845 191.275 20.100 191.830 ;
        RECT 20.935 191.675 21.830 191.845 ;
        RECT 22.000 191.890 22.170 192.915 ;
        RECT 22.355 193.025 22.525 193.275 ;
        RECT 22.695 193.195 22.945 193.655 ;
        RECT 23.115 193.025 23.285 193.485 ;
        RECT 22.355 192.855 23.285 193.025 ;
        RECT 22.370 192.375 22.850 192.675 ;
        RECT 22.590 191.955 22.850 192.375 ;
        RECT 23.050 191.955 23.310 192.675 ;
        RECT 23.545 192.490 23.835 193.655 ;
        RECT 24.930 192.515 25.185 193.655 ;
        RECT 25.355 192.685 25.685 193.485 ;
        RECT 25.855 192.855 26.025 193.655 ;
        RECT 26.195 192.685 26.525 193.485 ;
        RECT 26.695 192.855 26.865 193.655 ;
        RECT 27.035 192.685 27.365 193.485 ;
        RECT 27.535 192.855 27.705 193.655 ;
        RECT 27.875 192.685 28.205 193.485 ;
        RECT 28.375 192.855 28.625 193.655 ;
        RECT 25.355 192.515 28.205 192.685 ;
        RECT 29.135 192.685 29.495 193.485 ;
        RECT 30.040 192.855 30.210 193.655 ;
        RECT 30.420 193.025 30.750 193.485 ;
        RECT 30.920 193.195 31.090 193.655 ;
        RECT 31.260 193.025 31.590 193.485 ;
        RECT 30.420 192.855 31.590 193.025 ;
        RECT 31.760 192.855 31.930 193.655 ;
        RECT 31.260 192.685 31.590 192.855 ;
        RECT 29.135 192.515 30.595 192.685 ;
        RECT 31.260 192.515 32.115 192.685 ;
        RECT 24.950 192.095 26.570 192.345 ;
        RECT 26.750 192.095 27.285 192.515 ;
        RECT 27.455 192.095 28.895 192.345 ;
        RECT 22.000 191.720 22.350 191.890 ;
        RECT 22.590 191.785 22.855 191.955 ;
        RECT 23.050 191.785 23.315 191.955 ;
        RECT 20.270 191.105 20.700 191.550 ;
        RECT 20.935 191.275 21.105 191.675 ;
        RECT 21.275 191.105 22.010 191.505 ;
        RECT 22.180 191.275 22.350 191.720 ;
        RECT 22.925 191.105 23.325 191.615 ;
        RECT 23.545 191.105 23.835 191.830 ;
        RECT 24.930 191.735 26.865 191.925 ;
        RECT 24.930 191.275 25.265 191.735 ;
        RECT 25.435 191.105 25.605 191.565 ;
        RECT 25.775 191.275 26.105 191.735 ;
        RECT 26.275 191.105 26.445 191.565 ;
        RECT 26.615 191.485 26.865 191.735 ;
        RECT 27.035 191.825 27.285 192.095 ;
        RECT 27.035 191.655 28.205 191.825 ;
        RECT 28.375 191.485 28.625 191.905 ;
        RECT 29.070 191.785 29.325 192.345 ;
        RECT 29.495 191.845 29.675 192.515 ;
        RECT 29.845 192.015 30.220 192.345 ;
        RECT 30.390 192.265 30.595 192.515 ;
        RECT 30.390 192.095 31.600 192.265 ;
        RECT 31.770 191.925 32.115 192.515 ;
        RECT 32.745 192.565 35.335 193.655 ;
        RECT 35.515 192.845 35.810 193.655 ;
        RECT 32.745 192.045 33.955 192.565 ;
        RECT 26.615 191.275 28.625 191.485 ;
        RECT 29.085 191.105 29.325 191.615 ;
        RECT 29.495 191.310 29.825 191.845 ;
        RECT 30.040 191.105 30.210 191.845 ;
        RECT 30.420 191.755 32.115 191.925 ;
        RECT 34.125 191.875 35.335 192.395 ;
        RECT 35.990 192.345 36.235 193.485 ;
        RECT 36.410 192.845 36.670 193.655 ;
        RECT 37.270 193.650 43.545 193.655 ;
        RECT 36.850 192.345 37.100 193.480 ;
        RECT 37.270 192.855 37.530 193.650 ;
        RECT 37.700 192.755 37.960 193.480 ;
        RECT 38.130 192.925 38.390 193.650 ;
        RECT 38.560 192.755 38.820 193.480 ;
        RECT 38.990 192.925 39.250 193.650 ;
        RECT 39.420 192.755 39.680 193.480 ;
        RECT 39.850 192.925 40.110 193.650 ;
        RECT 40.280 192.755 40.540 193.480 ;
        RECT 40.710 192.925 40.955 193.650 ;
        RECT 41.125 192.755 41.385 193.480 ;
        RECT 41.570 192.925 41.815 193.650 ;
        RECT 41.985 192.755 42.245 193.480 ;
        RECT 42.430 192.925 42.675 193.650 ;
        RECT 42.845 192.755 43.105 193.480 ;
        RECT 43.290 192.925 43.545 193.650 ;
        RECT 37.700 192.740 43.105 192.755 ;
        RECT 43.715 192.740 44.005 193.480 ;
        RECT 44.175 192.910 44.445 193.655 ;
        RECT 37.700 192.515 44.445 192.740 ;
        RECT 44.710 192.655 44.965 193.655 ;
        RECT 30.420 191.285 30.750 191.755 ;
        RECT 30.920 191.105 31.090 191.585 ;
        RECT 31.260 191.285 31.590 191.755 ;
        RECT 31.760 191.105 31.930 191.585 ;
        RECT 32.745 191.105 35.335 191.875 ;
        RECT 35.505 191.785 35.820 192.345 ;
        RECT 35.990 192.095 43.110 192.345 ;
        RECT 35.505 191.105 35.810 191.615 ;
        RECT 35.990 191.285 36.240 192.095 ;
        RECT 36.410 191.105 36.670 191.630 ;
        RECT 36.850 191.285 37.100 192.095 ;
        RECT 43.280 191.925 44.445 192.515 ;
        RECT 37.700 191.755 44.445 191.925 ;
        RECT 37.270 191.105 37.530 191.665 ;
        RECT 37.700 191.300 37.960 191.755 ;
        RECT 38.130 191.105 38.390 191.585 ;
        RECT 38.560 191.300 38.820 191.755 ;
        RECT 38.990 191.105 39.250 191.585 ;
        RECT 39.420 191.300 39.680 191.755 ;
        RECT 39.850 191.105 40.095 191.585 ;
        RECT 40.265 191.300 40.540 191.755 ;
        RECT 40.710 191.105 40.955 191.585 ;
        RECT 41.125 191.300 41.385 191.755 ;
        RECT 41.565 191.105 41.815 191.585 ;
        RECT 41.985 191.300 42.245 191.755 ;
        RECT 42.425 191.105 42.675 191.585 ;
        RECT 42.845 191.300 43.105 191.755 ;
        RECT 43.285 191.105 43.545 191.585 ;
        RECT 43.715 191.300 43.975 191.755 ;
        RECT 44.145 191.105 44.445 191.585 ;
        RECT 44.725 191.105 44.965 191.905 ;
        RECT 45.150 191.275 45.395 193.485 ;
        RECT 45.565 193.205 46.415 193.655 ;
        RECT 46.585 193.025 46.845 193.485 ;
        RECT 45.725 192.805 46.845 193.025 ;
        RECT 45.725 192.350 45.895 192.805 ;
        RECT 45.565 191.860 45.895 192.350 ;
        RECT 46.065 192.030 46.475 192.635 ;
        RECT 47.025 192.420 47.230 193.005 ;
        RECT 47.415 192.670 47.740 193.655 ;
        RECT 47.965 192.515 48.195 193.655 ;
        RECT 48.365 192.505 48.695 193.485 ;
        RECT 48.865 192.515 49.075 193.655 ;
        RECT 46.645 192.295 47.230 192.420 ;
        RECT 46.645 192.125 47.235 192.295 ;
        RECT 46.645 192.045 47.230 192.125 ;
        RECT 47.485 192.015 47.745 192.470 ;
        RECT 47.945 192.095 48.275 192.345 ;
        RECT 45.565 191.655 46.415 191.860 ;
        RECT 45.565 191.105 45.895 191.485 ;
        RECT 46.085 191.275 46.415 191.655 ;
        RECT 46.585 191.655 47.740 191.845 ;
        RECT 46.585 191.485 46.795 191.655 ;
        RECT 47.465 191.515 47.740 191.655 ;
        RECT 46.965 191.105 47.295 191.485 ;
        RECT 47.965 191.105 48.195 191.925 ;
        RECT 48.445 191.905 48.695 192.505 ;
        RECT 49.305 192.490 49.595 193.655 ;
        RECT 49.775 192.685 50.105 193.470 ;
        RECT 49.775 192.515 50.455 192.685 ;
        RECT 50.635 192.515 50.965 193.655 ;
        RECT 51.145 192.895 51.810 193.485 ;
        RECT 49.765 192.095 50.115 192.345 ;
        RECT 48.365 191.275 48.695 191.905 ;
        RECT 48.865 191.105 49.075 191.925 ;
        RECT 50.285 191.915 50.455 192.515 ;
        RECT 50.625 192.095 50.975 192.345 ;
        RECT 51.145 191.925 51.395 192.895 ;
        RECT 51.980 192.815 52.310 193.655 ;
        RECT 52.820 193.065 53.625 193.485 ;
        RECT 52.480 192.895 54.045 193.065 ;
        RECT 52.480 192.645 52.650 192.895 ;
        RECT 51.730 192.475 52.650 192.645 ;
        RECT 52.820 192.635 53.195 192.725 ;
        RECT 51.730 192.305 51.900 192.475 ;
        RECT 52.820 192.465 53.215 192.635 ;
        RECT 52.820 192.305 53.195 192.465 ;
        RECT 51.565 192.095 51.900 192.305 ;
        RECT 52.070 192.095 52.520 192.305 ;
        RECT 52.710 192.095 53.195 192.305 ;
        RECT 53.385 192.345 53.705 192.725 ;
        RECT 53.875 192.645 54.045 192.895 ;
        RECT 54.215 192.815 54.465 193.655 ;
        RECT 54.660 192.645 54.960 193.485 ;
        RECT 53.875 192.475 54.960 192.645 ;
        RECT 55.755 193.315 56.925 193.485 ;
        RECT 55.755 192.645 56.085 193.315 ;
        RECT 56.595 193.275 56.925 193.315 ;
        RECT 57.095 193.275 57.470 193.655 ;
        RECT 56.255 193.105 56.485 193.145 ;
        RECT 56.255 193.055 56.870 193.105 ;
        RECT 57.615 193.055 57.785 193.185 ;
        RECT 56.255 192.855 57.785 193.055 ;
        RECT 58.020 192.875 58.285 193.655 ;
        RECT 56.255 192.815 57.135 192.855 ;
        RECT 57.275 192.645 58.335 192.685 ;
        RECT 55.755 192.515 58.335 192.645 ;
        RECT 58.505 192.515 58.785 193.655 ;
        RECT 53.385 192.095 53.765 192.345 ;
        RECT 53.945 192.095 54.275 192.305 ;
        RECT 49.305 191.105 49.595 191.830 ;
        RECT 49.785 191.105 50.025 191.915 ;
        RECT 50.195 191.275 50.525 191.915 ;
        RECT 50.695 191.105 50.965 191.915 ;
        RECT 51.145 191.285 51.830 191.925 ;
        RECT 52.000 191.105 52.170 191.925 ;
        RECT 52.340 191.755 54.040 191.925 ;
        RECT 52.340 191.290 52.670 191.755 ;
        RECT 53.655 191.665 54.040 191.755 ;
        RECT 54.445 191.845 54.615 192.475 ;
        RECT 55.755 192.465 57.500 192.515 ;
        RECT 54.785 192.015 55.115 192.305 ;
        RECT 54.445 191.665 54.955 191.845 ;
        RECT 55.785 191.785 56.235 192.295 ;
        RECT 56.425 192.095 56.900 192.295 ;
        RECT 56.650 191.695 56.900 192.095 ;
        RECT 57.150 192.095 57.500 192.295 ;
        RECT 57.150 191.695 57.360 192.095 ;
        RECT 57.670 192.015 57.995 192.345 ;
        RECT 58.165 191.845 58.335 192.515 ;
        RECT 58.955 192.505 59.285 193.485 ;
        RECT 59.455 192.515 59.715 193.655 ;
        RECT 58.515 192.075 58.850 192.345 ;
        RECT 59.020 191.905 59.190 192.505 ;
        RECT 59.360 192.095 59.695 192.345 ;
        RECT 52.840 191.105 53.010 191.575 ;
        RECT 53.270 191.325 54.455 191.495 ;
        RECT 54.625 191.275 54.955 191.665 ;
        RECT 57.605 191.675 58.335 191.845 ;
        RECT 55.755 191.105 56.205 191.615 ;
        RECT 57.605 191.525 57.785 191.675 ;
        RECT 56.480 191.275 57.785 191.525 ;
        RECT 57.965 191.105 58.295 191.505 ;
        RECT 58.505 191.105 58.815 191.905 ;
        RECT 59.020 191.275 59.715 191.905 ;
        RECT 60.360 191.285 60.640 193.475 ;
        RECT 60.830 192.515 61.115 193.655 ;
        RECT 61.380 193.005 61.550 193.475 ;
        RECT 61.725 193.175 62.055 193.655 ;
        RECT 62.225 193.005 62.405 193.475 ;
        RECT 61.380 192.805 62.405 193.005 ;
        RECT 60.840 191.835 61.100 192.345 ;
        RECT 61.310 192.015 61.570 192.635 ;
        RECT 61.765 192.015 62.190 192.635 ;
        RECT 62.575 192.365 62.905 193.475 ;
        RECT 63.075 193.245 63.425 193.655 ;
        RECT 63.595 193.065 63.835 193.455 ;
        RECT 62.360 192.065 62.905 192.365 ;
        RECT 63.085 192.865 63.835 193.065 ;
        RECT 63.085 192.185 63.425 192.865 ;
        RECT 62.360 191.835 62.580 192.065 ;
        RECT 60.840 191.645 62.580 191.835 ;
        RECT 60.840 191.105 61.570 191.475 ;
        RECT 62.150 191.285 62.580 191.645 ;
        RECT 62.750 191.105 62.995 191.885 ;
        RECT 63.195 191.285 63.425 192.185 ;
        RECT 63.605 191.345 63.835 192.685 ;
        RECT 64.040 191.285 64.320 193.475 ;
        RECT 64.510 192.515 64.795 193.655 ;
        RECT 65.060 193.005 65.230 193.475 ;
        RECT 65.405 193.175 65.735 193.655 ;
        RECT 65.905 193.005 66.085 193.475 ;
        RECT 65.060 192.805 66.085 193.005 ;
        RECT 64.520 191.835 64.780 192.345 ;
        RECT 64.990 192.015 65.250 192.635 ;
        RECT 65.445 192.015 65.870 192.635 ;
        RECT 66.255 192.365 66.585 193.475 ;
        RECT 66.755 193.245 67.105 193.655 ;
        RECT 67.275 193.065 67.515 193.455 ;
        RECT 68.720 193.275 69.050 193.655 ;
        RECT 69.220 193.095 69.410 193.485 ;
        RECT 66.040 192.065 66.585 192.365 ;
        RECT 66.765 192.865 67.515 193.065 ;
        RECT 68.680 192.925 69.410 193.095 ;
        RECT 69.590 192.955 70.020 193.655 ;
        RECT 66.765 192.185 67.105 192.865 ;
        RECT 66.040 191.835 66.260 192.065 ;
        RECT 64.520 191.645 66.260 191.835 ;
        RECT 64.520 191.105 65.250 191.475 ;
        RECT 65.830 191.285 66.260 191.645 ;
        RECT 66.430 191.105 66.675 191.885 ;
        RECT 66.875 191.285 67.105 192.185 ;
        RECT 67.285 191.345 67.515 192.685 ;
        RECT 68.680 191.805 68.875 192.925 ;
        RECT 70.525 192.785 71.195 193.485 ;
        RECT 71.365 192.955 71.695 193.655 ;
        RECT 71.865 192.785 72.130 193.485 ;
        RECT 69.555 192.530 72.130 192.785 ;
        RECT 72.315 192.705 72.590 193.475 ;
        RECT 72.760 193.045 73.090 193.475 ;
        RECT 73.260 193.215 73.455 193.655 ;
        RECT 73.635 193.045 73.965 193.475 ;
        RECT 72.760 192.875 73.965 193.045 ;
        RECT 69.555 192.345 69.725 192.530 ;
        RECT 69.045 192.015 69.725 192.345 ;
        RECT 69.895 192.015 70.230 192.345 ;
        RECT 70.400 192.295 70.690 192.345 ;
        RECT 70.400 192.125 70.695 192.295 ;
        RECT 70.400 192.015 70.690 192.125 ;
        RECT 70.980 192.015 71.340 192.345 ;
        RECT 71.510 191.845 71.690 192.530 ;
        RECT 72.315 192.515 72.900 192.705 ;
        RECT 73.070 192.545 73.965 192.875 ;
        RECT 71.860 192.015 72.135 192.345 ;
        RECT 68.680 191.635 69.500 191.805 ;
        RECT 70.070 191.655 71.340 191.845 ;
        RECT 68.670 191.105 69.000 191.465 ;
        RECT 69.170 191.275 69.500 191.635 ;
        RECT 69.670 191.105 69.905 191.545 ;
        RECT 70.495 191.105 70.830 191.485 ;
        RECT 71.510 191.445 72.125 191.845 ;
        RECT 72.315 191.695 72.555 192.345 ;
        RECT 72.725 191.845 72.900 192.515 ;
        RECT 75.065 192.490 75.355 193.655 ;
        RECT 76.745 193.015 77.075 193.445 ;
        RECT 76.620 192.845 77.075 193.015 ;
        RECT 77.255 193.015 77.505 193.435 ;
        RECT 77.735 193.185 78.065 193.655 ;
        RECT 78.295 193.015 78.545 193.435 ;
        RECT 77.255 192.845 78.545 193.015 ;
        RECT 73.070 192.015 73.485 192.345 ;
        RECT 73.665 192.015 73.960 192.345 ;
        RECT 72.725 191.665 73.055 191.845 ;
        RECT 71.790 191.275 72.125 191.445 ;
        RECT 72.330 191.105 72.660 191.495 ;
        RECT 72.830 191.285 73.055 191.665 ;
        RECT 73.255 191.395 73.485 192.015 ;
        RECT 76.620 191.845 76.790 192.845 ;
        RECT 76.960 192.015 77.205 192.675 ;
        RECT 77.420 192.015 77.685 192.675 ;
        RECT 77.880 192.015 78.165 192.675 ;
        RECT 78.340 192.345 78.555 192.675 ;
        RECT 78.735 192.515 78.985 193.655 ;
        RECT 79.155 192.595 79.485 193.445 ;
        RECT 78.340 192.015 78.645 192.345 ;
        RECT 78.815 192.015 79.125 192.345 ;
        RECT 78.815 191.845 78.985 192.015 ;
        RECT 73.665 191.105 73.965 191.835 ;
        RECT 75.065 191.105 75.355 191.830 ;
        RECT 76.620 191.675 78.985 191.845 ;
        RECT 79.295 191.830 79.485 192.595 ;
        RECT 76.775 191.105 77.105 191.505 ;
        RECT 77.275 191.335 77.605 191.675 ;
        RECT 78.655 191.105 78.985 191.505 ;
        RECT 79.155 191.320 79.485 191.830 ;
        RECT 79.665 192.515 79.940 193.485 ;
        RECT 80.150 192.855 80.430 193.655 ;
        RECT 80.600 193.145 82.215 193.475 ;
        RECT 80.600 192.805 81.775 192.975 ;
        RECT 80.600 192.685 80.770 192.805 ;
        RECT 80.110 192.515 80.770 192.685 ;
        RECT 79.665 191.780 79.835 192.515 ;
        RECT 80.110 192.345 80.280 192.515 ;
        RECT 81.030 192.345 81.275 192.635 ;
        RECT 81.445 192.515 81.775 192.805 ;
        RECT 82.035 192.345 82.205 192.905 ;
        RECT 82.455 192.515 82.715 193.655 ;
        RECT 83.345 192.815 83.605 193.485 ;
        RECT 83.775 193.255 84.105 193.655 ;
        RECT 84.975 193.255 85.375 193.655 ;
        RECT 85.665 193.075 85.995 193.310 ;
        RECT 83.915 192.905 85.995 193.075 ;
        RECT 80.005 192.015 80.280 192.345 ;
        RECT 80.450 192.015 81.275 192.345 ;
        RECT 81.490 192.015 82.205 192.345 ;
        RECT 82.375 192.095 82.710 192.345 ;
        RECT 80.110 191.845 80.280 192.015 ;
        RECT 81.955 191.925 82.205 192.015 ;
        RECT 79.665 191.435 79.940 191.780 ;
        RECT 80.110 191.675 81.775 191.845 ;
        RECT 80.130 191.105 80.505 191.505 ;
        RECT 80.675 191.325 80.845 191.675 ;
        RECT 81.015 191.105 81.345 191.505 ;
        RECT 81.515 191.275 81.775 191.675 ;
        RECT 81.955 191.505 82.285 191.925 ;
        RECT 82.455 191.105 82.715 191.925 ;
        RECT 83.345 191.845 83.520 192.815 ;
        RECT 83.915 192.635 84.085 192.905 ;
        RECT 83.690 192.465 84.085 192.635 ;
        RECT 84.255 192.515 85.270 192.735 ;
        RECT 83.690 192.015 83.860 192.465 ;
        RECT 84.995 192.375 85.270 192.515 ;
        RECT 85.440 192.515 85.995 192.905 ;
        RECT 84.030 192.095 84.480 192.295 ;
        RECT 84.650 191.925 84.825 192.120 ;
        RECT 83.345 191.275 83.685 191.845 ;
        RECT 83.880 191.105 84.050 191.770 ;
        RECT 84.330 191.755 84.825 191.925 ;
        RECT 84.330 191.615 84.550 191.755 ;
        RECT 84.325 191.445 84.550 191.615 ;
        RECT 84.995 191.585 85.165 192.375 ;
        RECT 85.440 192.265 85.610 192.515 ;
        RECT 86.165 192.345 86.340 193.445 ;
        RECT 86.510 192.835 86.855 193.655 ;
        RECT 85.415 192.095 85.610 192.265 ;
        RECT 85.780 192.095 86.340 192.345 ;
        RECT 86.510 192.095 86.855 192.665 ;
        RECT 87.025 192.565 89.615 193.655 ;
        RECT 89.790 193.220 95.135 193.655 ;
        RECT 95.310 193.220 100.655 193.655 ;
        RECT 85.415 191.710 85.585 192.095 ;
        RECT 87.025 192.045 88.235 192.565 ;
        RECT 84.330 191.400 84.550 191.445 ;
        RECT 84.720 191.415 85.165 191.585 ;
        RECT 85.335 191.340 85.585 191.710 ;
        RECT 85.755 191.745 86.855 191.925 ;
        RECT 88.405 191.875 89.615 192.395 ;
        RECT 91.380 191.970 91.730 193.220 ;
        RECT 85.755 191.340 86.005 191.745 ;
        RECT 86.175 191.105 86.345 191.575 ;
        RECT 86.515 191.340 86.855 191.745 ;
        RECT 87.025 191.105 89.615 191.875 ;
        RECT 93.210 191.650 93.550 192.480 ;
        RECT 96.900 191.970 97.250 193.220 ;
        RECT 100.825 192.490 101.115 193.655 ;
        RECT 101.745 192.565 105.255 193.655 ;
        RECT 105.425 192.935 105.885 193.485 ;
        RECT 106.075 192.935 106.405 193.655 ;
        RECT 98.730 191.650 99.070 192.480 ;
        RECT 101.745 192.045 103.435 192.565 ;
        RECT 103.605 191.875 105.255 192.395 ;
        RECT 89.790 191.105 95.135 191.650 ;
        RECT 95.310 191.105 100.655 191.650 ;
        RECT 100.825 191.105 101.115 191.830 ;
        RECT 101.745 191.105 105.255 191.875 ;
        RECT 105.425 191.565 105.675 192.935 ;
        RECT 106.605 192.765 106.905 193.315 ;
        RECT 107.075 192.985 107.355 193.655 ;
        RECT 107.725 193.145 107.985 193.655 ;
        RECT 105.965 192.595 106.905 192.765 ;
        RECT 105.965 192.345 106.135 192.595 ;
        RECT 107.275 192.345 107.540 192.705 ;
        RECT 105.845 192.015 106.135 192.345 ;
        RECT 106.305 192.095 106.645 192.345 ;
        RECT 106.865 192.095 107.540 192.345 ;
        RECT 107.725 192.095 108.065 192.975 ;
        RECT 108.235 192.265 108.405 193.485 ;
        RECT 108.645 193.150 109.260 193.655 ;
        RECT 108.645 192.615 108.895 192.980 ;
        RECT 109.065 192.975 109.260 193.150 ;
        RECT 109.430 193.145 109.905 193.485 ;
        RECT 110.075 193.110 110.290 193.655 ;
        RECT 109.065 192.785 109.395 192.975 ;
        RECT 109.615 192.615 110.330 192.910 ;
        RECT 110.500 192.785 110.775 193.485 ;
        RECT 108.645 192.445 110.435 192.615 ;
        RECT 105.965 191.925 106.135 192.015 ;
        RECT 108.235 192.015 109.030 192.265 ;
        RECT 108.235 191.925 108.485 192.015 ;
        RECT 105.965 191.735 107.355 191.925 ;
        RECT 105.425 191.275 105.985 191.565 ;
        RECT 106.155 191.105 106.405 191.565 ;
        RECT 107.025 191.375 107.355 191.735 ;
        RECT 107.725 191.105 107.985 191.925 ;
        RECT 108.155 191.505 108.485 191.925 ;
        RECT 109.200 191.590 109.455 192.445 ;
        RECT 108.665 191.325 109.455 191.590 ;
        RECT 109.625 191.745 110.035 192.265 ;
        RECT 110.205 192.015 110.435 192.445 ;
        RECT 110.605 191.755 110.775 192.785 ;
        RECT 109.625 191.325 109.825 191.745 ;
        RECT 110.015 191.105 110.345 191.565 ;
        RECT 110.515 191.275 110.775 191.755 ;
        RECT 110.945 193.105 111.205 193.485 ;
        RECT 111.375 193.275 111.705 193.655 ;
        RECT 112.045 193.105 112.215 193.485 ;
        RECT 112.385 193.275 112.725 193.655 ;
        RECT 112.895 193.105 113.065 193.485 ;
        RECT 113.300 193.275 113.970 193.655 ;
        RECT 114.615 193.275 114.945 193.655 ;
        RECT 110.945 192.935 111.875 193.105 ;
        RECT 112.045 192.935 113.225 193.105 ;
        RECT 115.115 193.075 115.285 193.485 ;
        RECT 116.010 193.220 121.355 193.655 ;
        RECT 110.945 191.605 111.115 192.935 ;
        RECT 111.705 192.765 111.875 192.935 ;
        RECT 111.705 192.595 112.885 192.765 ;
        RECT 111.285 191.785 111.635 192.325 ;
        RECT 110.945 191.275 111.205 191.605 ;
        RECT 111.375 191.105 111.625 191.605 ;
        RECT 111.805 191.445 112.110 192.425 ;
        RECT 112.715 192.420 112.885 192.595 ;
        RECT 112.285 192.125 112.555 192.295 ;
        RECT 112.285 191.440 112.550 192.125 ;
        RECT 113.055 191.825 113.225 192.935 ;
        RECT 113.535 192.905 115.285 193.075 ;
        RECT 113.535 192.345 113.705 192.905 ;
        RECT 114.140 192.565 114.470 192.735 ;
        RECT 113.395 192.015 113.705 192.345 ;
        RECT 113.875 191.825 114.045 192.345 ;
        RECT 113.055 191.655 114.045 191.825 ;
        RECT 113.280 191.275 113.450 191.655 ;
        RECT 113.720 191.105 114.050 191.485 ;
        RECT 114.220 191.275 114.445 192.565 ;
        RECT 114.790 191.825 114.960 192.905 ;
        RECT 115.130 192.295 115.310 192.655 ;
        RECT 115.130 192.125 115.315 192.295 ;
        RECT 115.130 192.015 115.310 192.125 ;
        RECT 117.600 191.970 117.950 193.220 ;
        RECT 121.615 192.725 121.785 193.485 ;
        RECT 121.965 192.895 122.295 193.655 ;
        RECT 121.615 192.555 122.280 192.725 ;
        RECT 122.465 192.580 122.735 193.485 ;
        RECT 123.830 193.230 124.165 193.655 ;
        RECT 124.335 193.050 124.520 193.455 ;
        RECT 114.790 191.655 115.285 191.825 ;
        RECT 114.615 191.105 114.945 191.485 ;
        RECT 115.115 191.275 115.285 191.655 ;
        RECT 119.430 191.650 119.770 192.480 ;
        RECT 122.110 192.410 122.280 192.555 ;
        RECT 121.545 192.005 121.875 192.375 ;
        RECT 122.110 192.080 122.395 192.410 ;
        RECT 122.110 191.825 122.280 192.080 ;
        RECT 121.615 191.655 122.280 191.825 ;
        RECT 122.565 191.780 122.735 192.580 ;
        RECT 116.010 191.105 121.355 191.650 ;
        RECT 121.615 191.275 121.785 191.655 ;
        RECT 121.965 191.105 122.295 191.485 ;
        RECT 122.475 191.275 122.735 191.780 ;
        RECT 123.855 192.875 124.520 193.050 ;
        RECT 124.725 192.875 125.055 193.655 ;
        RECT 123.855 191.845 124.195 192.875 ;
        RECT 125.225 192.685 125.495 193.455 ;
        RECT 124.365 192.515 125.495 192.685 ;
        RECT 124.365 192.015 124.615 192.515 ;
        RECT 123.855 191.675 124.540 191.845 ;
        RECT 124.795 191.765 125.155 192.345 ;
        RECT 123.830 191.105 124.165 191.505 ;
        RECT 124.335 191.275 124.540 191.675 ;
        RECT 125.325 191.605 125.495 192.515 ;
        RECT 125.665 192.565 126.875 193.655 ;
        RECT 125.665 192.025 126.185 192.565 ;
        RECT 126.355 191.855 126.875 192.395 ;
        RECT 124.750 191.105 125.025 191.585 ;
        RECT 125.235 191.275 125.495 191.605 ;
        RECT 125.665 191.105 126.875 191.855 ;
        RECT 14.260 190.935 126.960 191.105 ;
        RECT 14.345 190.185 15.555 190.935 ;
        RECT 14.345 189.645 14.865 190.185 ;
        RECT 15.730 190.095 15.990 190.935 ;
        RECT 16.165 190.190 16.420 190.765 ;
        RECT 16.590 190.555 16.920 190.935 ;
        RECT 17.135 190.385 17.305 190.765 ;
        RECT 18.115 190.455 18.415 190.935 ;
        RECT 16.590 190.215 17.305 190.385 ;
        RECT 18.585 190.285 18.845 190.740 ;
        RECT 19.015 190.455 19.275 190.935 ;
        RECT 19.455 190.285 19.715 190.740 ;
        RECT 19.885 190.455 20.135 190.935 ;
        RECT 20.315 190.285 20.575 190.740 ;
        RECT 20.745 190.455 20.995 190.935 ;
        RECT 21.175 190.285 21.435 190.740 ;
        RECT 21.605 190.455 21.850 190.935 ;
        RECT 22.020 190.285 22.295 190.740 ;
        RECT 22.465 190.455 22.710 190.935 ;
        RECT 22.880 190.285 23.140 190.740 ;
        RECT 23.310 190.455 23.570 190.935 ;
        RECT 23.740 190.285 24.000 190.740 ;
        RECT 24.170 190.455 24.430 190.935 ;
        RECT 24.600 190.285 24.860 190.740 ;
        RECT 25.030 190.375 25.290 190.935 ;
        RECT 15.035 189.475 15.555 190.015 ;
        RECT 14.345 188.385 15.555 189.475 ;
        RECT 15.730 188.385 15.990 189.535 ;
        RECT 16.165 189.460 16.335 190.190 ;
        RECT 16.590 190.025 16.760 190.215 ;
        RECT 18.115 190.115 24.860 190.285 ;
        RECT 16.505 189.695 16.760 190.025 ;
        RECT 16.590 189.485 16.760 189.695 ;
        RECT 17.040 189.665 17.395 190.035 ;
        RECT 18.115 189.525 19.280 190.115 ;
        RECT 25.460 189.945 25.710 190.755 ;
        RECT 25.890 190.410 26.150 190.935 ;
        RECT 26.320 189.945 26.570 190.755 ;
        RECT 26.750 190.425 27.055 190.935 ;
        RECT 27.315 190.455 27.615 190.935 ;
        RECT 27.785 190.285 28.045 190.740 ;
        RECT 28.215 190.455 28.475 190.935 ;
        RECT 28.655 190.285 28.915 190.740 ;
        RECT 29.085 190.455 29.335 190.935 ;
        RECT 29.515 190.285 29.775 190.740 ;
        RECT 29.945 190.455 30.195 190.935 ;
        RECT 30.375 190.285 30.635 190.740 ;
        RECT 30.805 190.455 31.050 190.935 ;
        RECT 31.220 190.285 31.495 190.740 ;
        RECT 31.665 190.455 31.910 190.935 ;
        RECT 32.080 190.285 32.340 190.740 ;
        RECT 32.510 190.455 32.770 190.935 ;
        RECT 32.940 190.285 33.200 190.740 ;
        RECT 33.370 190.455 33.630 190.935 ;
        RECT 33.800 190.285 34.060 190.740 ;
        RECT 34.230 190.375 34.490 190.935 ;
        RECT 19.450 189.695 26.570 189.945 ;
        RECT 26.740 189.695 27.055 190.255 ;
        RECT 27.315 190.115 34.060 190.285 ;
        RECT 16.165 188.555 16.420 189.460 ;
        RECT 16.590 189.315 17.305 189.485 ;
        RECT 16.590 188.385 16.920 189.145 ;
        RECT 17.135 188.555 17.305 189.315 ;
        RECT 18.115 189.300 24.860 189.525 ;
        RECT 18.115 188.385 18.385 189.130 ;
        RECT 18.555 188.560 18.845 189.300 ;
        RECT 19.455 189.285 24.860 189.300 ;
        RECT 19.015 188.390 19.270 189.115 ;
        RECT 19.455 188.560 19.715 189.285 ;
        RECT 19.885 188.390 20.130 189.115 ;
        RECT 20.315 188.560 20.575 189.285 ;
        RECT 20.745 188.390 20.990 189.115 ;
        RECT 21.175 188.560 21.435 189.285 ;
        RECT 21.605 188.390 21.850 189.115 ;
        RECT 22.020 188.560 22.280 189.285 ;
        RECT 22.450 188.390 22.710 189.115 ;
        RECT 22.880 188.560 23.140 189.285 ;
        RECT 23.310 188.390 23.570 189.115 ;
        RECT 23.740 188.560 24.000 189.285 ;
        RECT 24.170 188.390 24.430 189.115 ;
        RECT 24.600 188.560 24.860 189.285 ;
        RECT 25.030 188.390 25.290 189.185 ;
        RECT 25.460 188.560 25.710 189.695 ;
        RECT 19.015 188.385 25.290 188.390 ;
        RECT 25.890 188.385 26.150 189.195 ;
        RECT 26.325 188.555 26.570 189.695 ;
        RECT 27.315 189.525 28.480 190.115 ;
        RECT 34.660 189.945 34.910 190.755 ;
        RECT 35.090 190.410 35.350 190.935 ;
        RECT 35.520 189.945 35.770 190.755 ;
        RECT 35.950 190.425 36.255 190.935 ;
        RECT 28.650 189.695 35.770 189.945 ;
        RECT 35.940 189.695 36.255 190.255 ;
        RECT 36.425 190.210 36.715 190.935 ;
        RECT 36.885 190.135 37.580 190.765 ;
        RECT 37.785 190.135 38.095 190.935 ;
        RECT 38.265 190.135 38.525 190.935 ;
        RECT 36.905 189.695 37.240 189.945 ;
        RECT 27.315 189.300 34.060 189.525 ;
        RECT 26.750 188.385 27.045 189.195 ;
        RECT 27.315 188.385 27.585 189.130 ;
        RECT 27.755 188.560 28.045 189.300 ;
        RECT 28.655 189.285 34.060 189.300 ;
        RECT 28.215 188.390 28.470 189.115 ;
        RECT 28.655 188.560 28.915 189.285 ;
        RECT 29.085 188.390 29.330 189.115 ;
        RECT 29.515 188.560 29.775 189.285 ;
        RECT 29.945 188.390 30.190 189.115 ;
        RECT 30.375 188.560 30.635 189.285 ;
        RECT 30.805 188.390 31.050 189.115 ;
        RECT 31.220 188.560 31.480 189.285 ;
        RECT 31.650 188.390 31.910 189.115 ;
        RECT 32.080 188.560 32.340 189.285 ;
        RECT 32.510 188.390 32.770 189.115 ;
        RECT 32.940 188.560 33.200 189.285 ;
        RECT 33.370 188.390 33.630 189.115 ;
        RECT 33.800 188.560 34.060 189.285 ;
        RECT 34.230 188.390 34.490 189.185 ;
        RECT 34.660 188.560 34.910 189.695 ;
        RECT 28.215 188.385 34.490 188.390 ;
        RECT 35.090 188.385 35.350 189.195 ;
        RECT 35.525 188.555 35.770 189.695 ;
        RECT 35.950 188.385 36.245 189.195 ;
        RECT 36.425 188.385 36.715 189.550 ;
        RECT 37.410 189.535 37.580 190.135 ;
        RECT 37.750 189.695 38.085 189.965 ;
        RECT 36.885 188.385 37.145 189.525 ;
        RECT 37.315 188.555 37.645 189.535 ;
        RECT 37.815 188.385 38.095 189.525 ;
        RECT 38.265 188.385 38.525 189.525 ;
        RECT 38.695 188.555 39.025 190.765 ;
        RECT 39.275 190.195 39.605 190.935 ;
        RECT 39.875 190.365 40.205 190.765 ;
        RECT 40.375 190.535 40.705 190.935 ;
        RECT 40.875 190.595 42.235 190.765 ;
        RECT 40.875 190.365 41.205 190.595 ;
        RECT 39.875 190.195 41.205 190.365 ;
        RECT 41.375 190.195 41.705 190.425 ;
        RECT 39.195 189.235 39.505 190.025 ;
        RECT 39.675 189.405 39.895 190.025 ;
        RECT 40.165 189.405 40.340 190.025 ;
        RECT 40.595 189.405 40.815 190.025 ;
        RECT 41.090 189.575 41.335 190.025 ;
        RECT 41.085 189.405 41.335 189.575 ;
        RECT 41.505 189.235 41.705 190.195 ;
        RECT 41.875 190.115 42.235 190.595 ;
        RECT 42.405 190.165 45.915 190.935 ;
        RECT 41.875 189.775 42.235 189.945 ;
        RECT 41.905 189.695 42.235 189.775 ;
        RECT 39.195 189.065 41.705 189.235 ;
        RECT 39.195 188.385 39.705 188.895 ;
        RECT 40.875 188.555 41.205 189.065 ;
        RECT 41.875 188.385 42.235 189.525 ;
        RECT 42.405 189.475 44.095 189.995 ;
        RECT 44.265 189.645 45.915 190.165 ;
        RECT 46.105 190.125 46.345 190.935 ;
        RECT 46.515 190.125 46.845 190.765 ;
        RECT 47.015 190.125 47.285 190.935 ;
        RECT 47.465 190.425 47.770 190.935 ;
        RECT 46.085 189.695 46.435 189.945 ;
        RECT 46.605 189.525 46.775 190.125 ;
        RECT 46.945 189.695 47.295 189.945 ;
        RECT 47.465 189.695 47.780 190.255 ;
        RECT 47.950 189.945 48.200 190.755 ;
        RECT 48.370 190.410 48.630 190.935 ;
        RECT 48.810 189.945 49.060 190.755 ;
        RECT 49.230 190.375 49.490 190.935 ;
        RECT 49.660 190.285 49.920 190.740 ;
        RECT 50.090 190.455 50.350 190.935 ;
        RECT 50.520 190.285 50.780 190.740 ;
        RECT 50.950 190.455 51.210 190.935 ;
        RECT 51.380 190.285 51.640 190.740 ;
        RECT 51.810 190.455 52.055 190.935 ;
        RECT 52.225 190.285 52.500 190.740 ;
        RECT 52.670 190.455 52.915 190.935 ;
        RECT 53.085 190.285 53.345 190.740 ;
        RECT 53.525 190.455 53.775 190.935 ;
        RECT 53.945 190.285 54.205 190.740 ;
        RECT 54.385 190.455 54.635 190.935 ;
        RECT 54.805 190.285 55.065 190.740 ;
        RECT 55.245 190.455 55.505 190.935 ;
        RECT 55.675 190.285 55.935 190.740 ;
        RECT 56.105 190.455 56.405 190.935 ;
        RECT 49.660 190.115 56.405 190.285 ;
        RECT 56.670 190.170 57.125 190.935 ;
        RECT 57.400 190.555 58.700 190.765 ;
        RECT 58.955 190.575 59.285 190.935 ;
        RECT 58.530 190.405 58.700 190.555 ;
        RECT 59.455 190.435 59.715 190.765 ;
        RECT 59.485 190.425 59.715 190.435 ;
        RECT 47.950 189.695 55.070 189.945 ;
        RECT 42.405 188.385 45.915 189.475 ;
        RECT 46.095 189.355 46.775 189.525 ;
        RECT 46.095 188.570 46.425 189.355 ;
        RECT 46.955 188.385 47.285 189.525 ;
        RECT 47.475 188.385 47.770 189.195 ;
        RECT 47.950 188.555 48.195 189.695 ;
        RECT 48.370 188.385 48.630 189.195 ;
        RECT 48.810 188.560 49.060 189.695 ;
        RECT 55.240 189.525 56.405 190.115 ;
        RECT 57.600 189.945 57.820 190.345 ;
        RECT 56.665 189.745 57.155 189.945 ;
        RECT 57.345 189.735 57.820 189.945 ;
        RECT 58.065 189.945 58.275 190.345 ;
        RECT 58.530 190.280 59.285 190.405 ;
        RECT 58.530 190.235 59.375 190.280 ;
        RECT 59.105 190.115 59.375 190.235 ;
        RECT 58.065 189.735 58.395 189.945 ;
        RECT 58.565 189.675 58.975 189.980 ;
        RECT 49.660 189.300 56.405 189.525 ;
        RECT 56.670 189.505 57.845 189.565 ;
        RECT 59.205 189.540 59.375 190.115 ;
        RECT 59.175 189.505 59.375 189.540 ;
        RECT 56.670 189.395 59.375 189.505 ;
        RECT 49.660 189.285 55.065 189.300 ;
        RECT 49.230 188.390 49.490 189.185 ;
        RECT 49.660 188.560 49.920 189.285 ;
        RECT 50.090 188.390 50.350 189.115 ;
        RECT 50.520 188.560 50.780 189.285 ;
        RECT 50.950 188.390 51.210 189.115 ;
        RECT 51.380 188.560 51.640 189.285 ;
        RECT 51.810 188.390 52.070 189.115 ;
        RECT 52.240 188.560 52.500 189.285 ;
        RECT 52.670 188.390 52.915 189.115 ;
        RECT 53.085 188.560 53.345 189.285 ;
        RECT 53.530 188.390 53.775 189.115 ;
        RECT 53.945 188.560 54.205 189.285 ;
        RECT 54.390 188.390 54.635 189.115 ;
        RECT 54.805 188.560 55.065 189.285 ;
        RECT 55.250 188.390 55.505 189.115 ;
        RECT 55.675 188.560 55.965 189.300 ;
        RECT 49.230 188.385 55.505 188.390 ;
        RECT 56.135 188.385 56.405 189.130 ;
        RECT 56.670 188.775 56.925 189.395 ;
        RECT 57.515 189.335 59.315 189.395 ;
        RECT 57.515 189.305 57.845 189.335 ;
        RECT 59.545 189.235 59.715 190.425 ;
        RECT 59.905 190.125 60.145 190.935 ;
        RECT 60.315 190.125 60.645 190.765 ;
        RECT 60.815 190.125 61.085 190.935 ;
        RECT 62.185 190.210 62.475 190.935 ;
        RECT 62.645 190.260 62.905 190.765 ;
        RECT 63.085 190.555 63.415 190.935 ;
        RECT 63.595 190.385 63.765 190.765 ;
        RECT 59.885 189.695 60.235 189.945 ;
        RECT 60.405 189.525 60.575 190.125 ;
        RECT 60.745 189.695 61.095 189.945 ;
        RECT 57.175 189.135 57.360 189.225 ;
        RECT 57.950 189.135 58.785 189.145 ;
        RECT 57.175 188.935 58.785 189.135 ;
        RECT 57.175 188.895 57.405 188.935 ;
        RECT 56.670 188.555 57.005 188.775 ;
        RECT 58.010 188.385 58.365 188.765 ;
        RECT 58.535 188.555 58.785 188.935 ;
        RECT 59.035 188.385 59.285 189.165 ;
        RECT 59.455 188.555 59.715 189.235 ;
        RECT 59.895 189.355 60.575 189.525 ;
        RECT 59.895 188.570 60.225 189.355 ;
        RECT 60.755 188.385 61.085 189.525 ;
        RECT 62.185 188.385 62.475 189.550 ;
        RECT 62.645 189.460 62.815 190.260 ;
        RECT 63.100 190.215 63.765 190.385 ;
        RECT 63.100 189.960 63.270 190.215 ;
        RECT 62.985 189.630 63.270 189.960 ;
        RECT 63.505 189.665 63.835 190.035 ;
        RECT 63.100 189.485 63.270 189.630 ;
        RECT 62.645 188.555 62.915 189.460 ;
        RECT 63.100 189.315 63.765 189.485 ;
        RECT 63.085 188.385 63.415 189.145 ;
        RECT 63.595 188.555 63.765 189.315 ;
        RECT 64.025 188.555 64.775 190.765 ;
        RECT 65.875 190.205 66.175 190.935 ;
        RECT 66.355 190.025 66.585 190.645 ;
        RECT 66.785 190.375 67.010 190.755 ;
        RECT 67.180 190.545 67.510 190.935 ;
        RECT 67.790 190.385 68.120 190.765 ;
        RECT 68.290 190.555 69.475 190.725 ;
        RECT 69.735 190.465 69.905 190.935 ;
        RECT 66.785 190.195 67.115 190.375 ;
        RECT 65.880 189.695 66.175 190.025 ;
        RECT 66.355 189.695 66.770 190.025 ;
        RECT 66.940 189.525 67.115 190.195 ;
        RECT 67.285 189.695 67.525 190.345 ;
        RECT 67.790 190.215 68.335 190.385 ;
        RECT 67.705 189.695 67.965 190.045 ;
        RECT 68.165 189.575 68.335 190.215 ;
        RECT 68.705 190.285 69.090 190.375 ;
        RECT 70.075 190.285 70.405 190.750 ;
        RECT 68.705 190.115 70.405 190.285 ;
        RECT 70.575 190.115 70.745 190.935 ;
        RECT 70.915 190.285 71.245 190.755 ;
        RECT 71.415 190.455 71.585 190.935 ;
        RECT 70.915 190.115 71.675 190.285 ;
        RECT 68.505 189.745 68.850 189.945 ;
        RECT 69.020 189.745 69.410 189.945 ;
        RECT 68.165 189.525 68.950 189.575 ;
        RECT 65.875 189.165 66.770 189.495 ;
        RECT 66.940 189.335 67.525 189.525 ;
        RECT 65.875 188.995 67.080 189.165 ;
        RECT 65.875 188.565 66.205 188.995 ;
        RECT 66.385 188.385 66.580 188.825 ;
        RECT 66.750 188.565 67.080 188.995 ;
        RECT 67.250 188.565 67.525 189.335 ;
        RECT 67.870 189.350 68.950 189.525 ;
        RECT 67.870 188.555 68.200 189.350 ;
        RECT 68.370 188.385 68.610 189.170 ;
        RECT 68.780 189.145 68.950 189.350 ;
        RECT 69.120 189.315 69.410 189.745 ;
        RECT 69.600 189.735 70.085 189.945 ;
        RECT 70.255 189.735 70.695 189.945 ;
        RECT 70.865 189.735 71.195 189.945 ;
        RECT 69.600 189.315 69.905 189.735 ;
        RECT 70.865 189.565 71.035 189.735 ;
        RECT 70.075 189.395 71.035 189.565 ;
        RECT 70.075 189.145 70.245 189.395 ;
        RECT 68.780 188.975 70.245 189.145 ;
        RECT 69.170 188.555 69.925 188.975 ;
        RECT 70.415 188.385 70.745 189.225 ;
        RECT 71.365 189.145 71.675 190.115 ;
        RECT 70.915 188.975 71.675 189.145 ;
        RECT 70.915 188.555 71.165 188.975 ;
        RECT 71.335 188.385 71.675 188.805 ;
        RECT 71.845 188.555 72.125 190.655 ;
        RECT 72.355 190.475 72.525 190.935 ;
        RECT 72.795 190.545 74.045 190.725 ;
        RECT 73.180 190.305 73.545 190.375 ;
        RECT 72.295 190.125 73.545 190.305 ;
        RECT 73.715 190.325 74.045 190.545 ;
        RECT 74.215 190.495 74.385 190.935 ;
        RECT 74.555 190.325 74.895 190.740 ;
        RECT 73.715 190.155 74.895 190.325 ;
        RECT 75.065 190.165 76.735 190.935 ;
        RECT 72.295 189.525 72.570 190.125 ;
        RECT 72.740 189.695 73.095 189.945 ;
        RECT 73.290 189.915 73.755 189.945 ;
        RECT 73.285 189.745 73.755 189.915 ;
        RECT 73.290 189.695 73.755 189.745 ;
        RECT 73.925 189.695 74.255 189.945 ;
        RECT 74.430 189.745 74.895 189.945 ;
        RECT 74.075 189.575 74.255 189.695 ;
        RECT 72.295 189.315 73.905 189.525 ;
        RECT 74.075 189.405 74.405 189.575 ;
        RECT 73.495 189.215 73.905 189.315 ;
        RECT 72.315 188.385 73.100 189.145 ;
        RECT 73.495 188.555 73.880 189.215 ;
        RECT 74.205 188.615 74.405 189.405 ;
        RECT 74.575 188.385 74.895 189.565 ;
        RECT 75.065 189.475 75.815 189.995 ;
        RECT 75.985 189.645 76.735 190.165 ;
        RECT 76.905 190.135 77.215 190.935 ;
        RECT 77.420 190.135 78.115 190.765 ;
        RECT 76.915 189.695 77.250 189.965 ;
        RECT 77.420 189.535 77.590 190.135 ;
        RECT 77.760 189.695 78.095 189.945 ;
        RECT 75.065 188.385 76.735 189.475 ;
        RECT 76.905 188.385 77.185 189.525 ;
        RECT 77.355 188.555 77.685 189.535 ;
        RECT 77.855 188.385 78.115 189.525 ;
        RECT 78.295 188.565 78.555 190.755 ;
        RECT 78.815 190.565 79.485 190.935 ;
        RECT 79.665 190.385 79.975 190.755 ;
        RECT 78.745 190.185 79.975 190.385 ;
        RECT 78.745 189.515 79.035 190.185 ;
        RECT 80.155 190.005 80.385 190.645 ;
        RECT 80.565 190.205 80.855 190.935 ;
        RECT 81.045 190.260 81.320 190.605 ;
        RECT 81.510 190.535 81.885 190.935 ;
        RECT 82.055 190.365 82.225 190.715 ;
        RECT 82.395 190.535 82.725 190.935 ;
        RECT 82.895 190.365 83.155 190.765 ;
        RECT 79.215 189.695 79.680 190.005 ;
        RECT 79.860 189.695 80.385 190.005 ;
        RECT 80.565 189.695 80.865 190.025 ;
        RECT 81.045 189.525 81.215 190.260 ;
        RECT 81.490 190.195 83.155 190.365 ;
        RECT 81.490 190.025 81.660 190.195 ;
        RECT 83.335 190.115 83.665 190.535 ;
        RECT 83.835 190.115 84.095 190.935 ;
        RECT 85.205 190.245 85.445 190.765 ;
        RECT 85.615 190.440 86.010 190.935 ;
        RECT 86.575 190.605 86.745 190.750 ;
        RECT 86.370 190.410 86.745 190.605 ;
        RECT 83.335 190.025 83.585 190.115 ;
        RECT 81.385 189.695 81.660 190.025 ;
        RECT 81.830 189.695 82.655 190.025 ;
        RECT 82.870 189.695 83.585 190.025 ;
        RECT 83.755 189.695 84.090 189.945 ;
        RECT 81.490 189.525 81.660 189.695 ;
        RECT 78.745 189.295 79.515 189.515 ;
        RECT 78.725 188.385 79.065 189.115 ;
        RECT 79.245 188.565 79.515 189.295 ;
        RECT 79.695 189.275 80.855 189.515 ;
        RECT 79.695 188.565 79.925 189.275 ;
        RECT 80.095 188.385 80.425 189.095 ;
        RECT 80.595 188.565 80.855 189.275 ;
        RECT 81.045 188.555 81.320 189.525 ;
        RECT 81.490 189.355 82.150 189.525 ;
        RECT 82.410 189.405 82.655 189.695 ;
        RECT 81.980 189.235 82.150 189.355 ;
        RECT 82.825 189.235 83.155 189.525 ;
        RECT 81.530 188.385 81.810 189.185 ;
        RECT 81.980 189.065 83.155 189.235 ;
        RECT 83.415 189.135 83.585 189.695 ;
        RECT 81.980 188.565 83.595 188.895 ;
        RECT 83.835 188.385 84.095 189.525 ;
        RECT 85.205 189.440 85.380 190.245 ;
        RECT 86.370 190.075 86.540 190.410 ;
        RECT 87.025 190.365 87.265 190.740 ;
        RECT 87.435 190.430 87.770 190.935 ;
        RECT 87.025 190.215 87.245 190.365 ;
        RECT 85.555 189.715 86.540 190.075 ;
        RECT 86.710 189.885 87.245 190.215 ;
        RECT 85.555 189.695 86.840 189.715 ;
        RECT 85.980 189.545 86.840 189.695 ;
        RECT 85.205 188.655 85.510 189.440 ;
        RECT 85.685 189.065 86.380 189.375 ;
        RECT 85.690 188.385 86.375 188.855 ;
        RECT 86.555 188.600 86.840 189.545 ;
        RECT 87.010 189.235 87.245 189.885 ;
        RECT 87.415 189.405 87.715 190.255 ;
        RECT 87.945 190.210 88.235 190.935 ;
        RECT 88.865 190.165 92.375 190.935 ;
        RECT 87.010 189.005 87.685 189.235 ;
        RECT 87.015 188.385 87.345 188.835 ;
        RECT 87.515 188.575 87.685 189.005 ;
        RECT 87.945 188.385 88.235 189.550 ;
        RECT 88.865 189.475 90.555 189.995 ;
        RECT 90.725 189.645 92.375 190.165 ;
        RECT 92.605 190.115 92.815 190.935 ;
        RECT 92.985 190.135 93.315 190.765 ;
        RECT 92.985 189.535 93.235 190.135 ;
        RECT 93.485 190.115 93.715 190.935 ;
        RECT 94.390 190.390 99.735 190.935 ;
        RECT 99.930 190.545 100.260 190.935 ;
        RECT 93.405 189.695 93.735 189.945 ;
        RECT 88.865 188.385 92.375 189.475 ;
        RECT 92.605 188.385 92.815 189.525 ;
        RECT 92.985 188.555 93.315 189.535 ;
        RECT 93.485 188.385 93.715 189.525 ;
        RECT 95.980 188.820 96.330 190.070 ;
        RECT 97.810 189.560 98.150 190.390 ;
        RECT 100.430 190.375 100.655 190.755 ;
        RECT 99.915 189.695 100.155 190.345 ;
        RECT 100.325 190.195 100.655 190.375 ;
        RECT 100.325 189.525 100.500 190.195 ;
        RECT 100.855 190.025 101.085 190.645 ;
        RECT 101.265 190.205 101.565 190.935 ;
        RECT 102.665 190.195 103.025 190.570 ;
        RECT 103.290 190.195 103.460 190.935 ;
        RECT 103.740 190.365 103.910 190.570 ;
        RECT 103.740 190.195 104.280 190.365 ;
        RECT 100.670 189.695 101.085 190.025 ;
        RECT 101.265 189.695 101.560 190.025 ;
        RECT 99.915 189.335 100.500 189.525 ;
        RECT 102.665 189.540 102.920 190.195 ;
        RECT 103.090 189.695 103.440 190.025 ;
        RECT 103.610 189.695 103.940 190.025 ;
        RECT 94.390 188.385 99.735 188.820 ;
        RECT 99.915 188.565 100.190 189.335 ;
        RECT 100.670 189.165 101.565 189.495 ;
        RECT 100.360 188.995 101.565 189.165 ;
        RECT 100.360 188.565 100.690 188.995 ;
        RECT 100.860 188.385 101.055 188.825 ;
        RECT 101.235 188.565 101.565 188.995 ;
        RECT 102.665 188.555 103.005 189.540 ;
        RECT 103.175 189.155 103.440 189.695 ;
        RECT 104.110 189.495 104.280 190.195 ;
        RECT 103.655 189.325 104.280 189.495 ;
        RECT 104.450 189.565 104.620 190.765 ;
        RECT 104.850 190.285 105.180 190.765 ;
        RECT 105.350 190.465 105.520 190.935 ;
        RECT 105.690 190.285 106.020 190.750 ;
        RECT 104.850 190.115 106.020 190.285 ;
        RECT 106.345 190.165 109.855 190.935 ;
        RECT 110.030 190.680 110.365 190.725 ;
        RECT 104.790 189.735 105.360 189.945 ;
        RECT 105.530 189.735 106.175 189.945 ;
        RECT 104.450 189.155 105.155 189.565 ;
        RECT 103.175 188.985 105.155 189.155 ;
        RECT 103.175 188.385 103.585 188.815 ;
        RECT 104.330 188.385 104.660 188.805 ;
        RECT 104.830 188.555 105.155 188.985 ;
        RECT 105.630 188.385 105.960 189.485 ;
        RECT 106.345 189.475 108.035 189.995 ;
        RECT 108.205 189.645 109.855 190.165 ;
        RECT 110.025 190.215 110.365 190.680 ;
        RECT 110.535 190.555 110.865 190.935 ;
        RECT 111.325 190.595 111.595 190.600 ;
        RECT 111.325 190.425 111.635 190.595 ;
        RECT 110.025 189.525 110.195 190.215 ;
        RECT 110.365 189.695 110.625 190.025 ;
        RECT 106.345 188.385 109.855 189.475 ;
        RECT 110.025 188.555 110.285 189.525 ;
        RECT 110.455 189.145 110.625 189.695 ;
        RECT 110.795 189.325 111.135 190.355 ;
        RECT 111.325 189.325 111.595 190.425 ;
        RECT 111.820 189.325 112.100 190.600 ;
        RECT 112.300 190.435 112.530 190.765 ;
        RECT 112.775 190.555 113.105 190.935 ;
        RECT 112.300 189.145 112.470 190.435 ;
        RECT 113.275 190.365 113.450 190.765 ;
        RECT 112.820 190.195 113.450 190.365 ;
        RECT 113.705 190.210 113.995 190.935 ;
        RECT 112.820 190.025 112.990 190.195 ;
        RECT 114.165 190.135 114.455 190.935 ;
        RECT 114.625 190.475 115.175 190.765 ;
        RECT 115.345 190.475 115.595 190.935 ;
        RECT 112.640 189.695 112.990 190.025 ;
        RECT 110.455 188.975 112.470 189.145 ;
        RECT 112.820 189.175 112.990 189.695 ;
        RECT 113.170 189.345 113.535 190.025 ;
        RECT 112.820 189.005 113.450 189.175 ;
        RECT 110.480 188.385 110.810 188.795 ;
        RECT 111.010 188.555 111.180 188.975 ;
        RECT 111.395 188.385 112.065 188.795 ;
        RECT 112.300 188.555 112.470 188.975 ;
        RECT 112.775 188.385 113.105 188.825 ;
        RECT 113.275 188.555 113.450 189.005 ;
        RECT 113.705 188.385 113.995 189.550 ;
        RECT 114.165 188.385 114.455 189.525 ;
        RECT 114.625 189.105 114.875 190.475 ;
        RECT 116.225 190.305 116.555 190.665 ;
        RECT 115.165 190.115 116.555 190.305 ;
        RECT 116.945 190.245 117.185 190.765 ;
        RECT 117.355 190.440 117.750 190.935 ;
        RECT 118.315 190.605 118.485 190.750 ;
        RECT 118.110 190.410 118.485 190.605 ;
        RECT 115.165 190.025 115.335 190.115 ;
        RECT 115.045 189.695 115.335 190.025 ;
        RECT 115.505 189.695 115.835 189.945 ;
        RECT 116.065 189.695 116.755 189.945 ;
        RECT 115.165 189.445 115.335 189.695 ;
        RECT 115.165 189.275 116.105 189.445 ;
        RECT 114.625 188.555 115.075 189.105 ;
        RECT 115.265 188.385 115.595 189.105 ;
        RECT 115.805 188.725 116.105 189.275 ;
        RECT 116.440 189.255 116.755 189.695 ;
        RECT 116.945 189.440 117.120 190.245 ;
        RECT 118.110 190.075 118.280 190.410 ;
        RECT 118.765 190.365 119.005 190.740 ;
        RECT 119.175 190.430 119.510 190.935 ;
        RECT 118.765 190.215 118.985 190.365 ;
        RECT 119.685 190.300 119.955 190.935 ;
        RECT 117.295 189.715 118.280 190.075 ;
        RECT 118.450 189.885 118.985 190.215 ;
        RECT 117.295 189.695 118.580 189.715 ;
        RECT 117.720 189.545 118.580 189.695 ;
        RECT 116.275 188.385 116.555 189.055 ;
        RECT 116.945 188.655 117.250 189.440 ;
        RECT 117.425 189.065 118.120 189.375 ;
        RECT 117.430 188.385 118.115 188.855 ;
        RECT 118.295 188.600 118.580 189.545 ;
        RECT 118.750 189.235 118.985 189.885 ;
        RECT 119.155 189.405 119.455 190.255 ;
        RECT 120.140 190.245 120.375 190.765 ;
        RECT 120.545 190.440 120.945 190.935 ;
        RECT 121.535 190.605 121.705 190.750 ;
        RECT 121.305 190.410 121.705 190.605 ;
        RECT 120.140 189.440 120.315 190.245 ;
        RECT 121.305 190.075 121.475 190.410 ;
        RECT 121.985 190.365 122.225 190.740 ;
        RECT 122.395 190.430 122.725 190.935 ;
        RECT 121.985 190.215 122.200 190.365 ;
        RECT 120.485 189.715 121.475 190.075 ;
        RECT 121.645 189.885 122.200 190.215 ;
        RECT 120.485 189.695 121.775 189.715 ;
        RECT 120.915 189.545 121.775 189.695 ;
        RECT 118.750 189.005 119.425 189.235 ;
        RECT 118.755 188.385 119.085 188.835 ;
        RECT 119.255 188.575 119.425 189.005 ;
        RECT 119.685 188.385 119.955 189.340 ;
        RECT 120.140 188.655 120.445 189.440 ;
        RECT 120.620 189.065 121.315 189.375 ;
        RECT 120.625 188.385 121.310 188.855 ;
        RECT 121.490 188.600 121.775 189.545 ;
        RECT 121.965 189.235 122.200 189.885 ;
        RECT 122.370 189.575 122.670 190.255 ;
        RECT 122.965 190.115 123.175 190.935 ;
        RECT 123.345 190.135 123.675 190.765 ;
        RECT 122.370 189.405 122.675 189.575 ;
        RECT 123.345 189.535 123.595 190.135 ;
        RECT 123.845 190.115 124.075 190.935 ;
        RECT 124.285 190.185 125.495 190.935 ;
        RECT 125.665 190.185 126.875 190.935 ;
        RECT 123.765 189.695 124.095 189.945 ;
        RECT 121.965 189.005 122.645 189.235 ;
        RECT 121.975 188.385 122.305 188.835 ;
        RECT 122.475 188.575 122.645 189.005 ;
        RECT 122.965 188.385 123.175 189.525 ;
        RECT 123.345 188.555 123.675 189.535 ;
        RECT 123.845 188.385 124.075 189.525 ;
        RECT 124.285 189.475 124.805 190.015 ;
        RECT 124.975 189.645 125.495 190.185 ;
        RECT 125.665 189.475 126.185 190.015 ;
        RECT 126.355 189.645 126.875 190.185 ;
        RECT 124.285 188.385 125.495 189.475 ;
        RECT 125.665 188.385 126.875 189.475 ;
        RECT 14.260 188.215 126.960 188.385 ;
        RECT 14.345 187.125 15.555 188.215 ;
        RECT 14.345 186.415 14.865 186.955 ;
        RECT 15.035 186.585 15.555 187.125 ;
        RECT 15.725 187.045 16.020 188.215 ;
        RECT 16.190 187.415 16.630 188.045 ;
        RECT 16.190 186.875 16.500 187.415 ;
        RECT 16.805 187.365 17.120 188.215 ;
        RECT 17.290 187.875 18.720 188.045 ;
        RECT 17.290 187.195 17.460 187.875 ;
        RECT 15.725 186.655 16.500 186.875 ;
        RECT 14.345 185.665 15.555 186.415 ;
        RECT 15.725 185.665 16.020 186.485 ;
        RECT 16.190 186.405 16.500 186.655 ;
        RECT 16.670 187.025 17.460 187.195 ;
        RECT 16.670 186.575 16.840 187.025 ;
        RECT 17.630 186.905 17.830 187.705 ;
        RECT 17.010 186.575 17.400 186.855 ;
        RECT 17.585 186.575 17.830 186.905 ;
        RECT 18.030 186.575 18.280 187.705 ;
        RECT 18.470 187.245 18.720 187.875 ;
        RECT 18.895 187.415 19.230 188.215 ;
        RECT 19.495 187.245 19.665 188.045 ;
        RECT 20.435 187.585 20.745 188.045 ;
        RECT 21.005 187.835 21.335 188.215 ;
        RECT 21.620 187.585 21.870 188.045 ;
        RECT 20.435 187.415 21.870 187.585 ;
        RECT 22.080 187.415 22.300 188.215 ;
        RECT 18.470 187.075 19.235 187.245 ;
        RECT 19.495 187.075 22.445 187.245 ;
        RECT 18.495 186.575 18.895 186.905 ;
        RECT 19.065 186.405 19.235 187.075 ;
        RECT 19.455 186.575 19.765 186.905 ;
        RECT 20.225 186.575 20.565 186.905 ;
        RECT 20.785 186.575 21.020 186.905 ;
        RECT 16.190 185.845 16.630 186.405 ;
        RECT 16.800 185.665 17.250 186.405 ;
        RECT 17.420 186.235 18.580 186.405 ;
        RECT 17.420 185.835 17.590 186.235 ;
        RECT 17.760 185.665 18.180 186.065 ;
        RECT 18.350 185.835 18.580 186.235 ;
        RECT 18.750 185.835 19.235 186.405 ;
        RECT 19.495 186.235 20.670 186.405 ;
        RECT 19.495 185.835 19.665 186.235 ;
        RECT 19.910 185.665 20.240 186.065 ;
        RECT 20.500 186.005 20.670 186.235 ;
        RECT 20.840 186.185 21.020 186.575 ;
        RECT 21.295 186.185 21.565 186.905 ;
        RECT 21.750 186.575 21.965 186.905 ;
        RECT 22.275 186.405 22.445 187.075 ;
        RECT 21.765 186.235 22.445 186.405 ;
        RECT 21.765 186.005 21.935 186.235 ;
        RECT 20.500 185.835 21.935 186.005 ;
        RECT 22.115 185.665 22.445 186.045 ;
        RECT 22.615 185.875 22.945 188.005 ;
        RECT 23.115 187.075 23.370 188.215 ;
        RECT 23.545 187.050 23.835 188.215 ;
        RECT 24.060 187.345 24.345 188.215 ;
        RECT 24.515 187.585 24.775 188.045 ;
        RECT 24.950 187.755 25.205 188.215 ;
        RECT 25.375 187.585 25.635 188.045 ;
        RECT 24.515 187.415 25.635 187.585 ;
        RECT 25.805 187.415 26.115 188.215 ;
        RECT 24.515 187.165 24.775 187.415 ;
        RECT 26.285 187.245 26.595 188.045 ;
        RECT 24.020 186.995 24.775 187.165 ;
        RECT 25.565 187.075 26.595 187.245 ;
        RECT 24.020 186.485 24.425 186.995 ;
        RECT 25.565 186.825 25.735 187.075 ;
        RECT 24.595 186.655 25.735 186.825 ;
        RECT 23.115 185.665 23.370 186.465 ;
        RECT 23.545 185.665 23.835 186.390 ;
        RECT 24.020 186.315 25.670 186.485 ;
        RECT 25.905 186.335 26.255 186.905 ;
        RECT 24.065 185.665 24.345 186.145 ;
        RECT 24.515 185.925 24.775 186.315 ;
        RECT 24.950 185.665 25.205 186.145 ;
        RECT 25.375 185.925 25.670 186.315 ;
        RECT 26.425 186.165 26.595 187.075 ;
        RECT 25.850 185.665 26.125 186.145 ;
        RECT 26.295 185.835 26.595 186.165 ;
        RECT 26.765 187.140 27.035 188.045 ;
        RECT 27.205 187.455 27.535 188.215 ;
        RECT 27.715 187.285 27.885 188.045 ;
        RECT 26.765 186.340 26.935 187.140 ;
        RECT 27.220 187.115 27.885 187.285 ;
        RECT 27.220 186.970 27.390 187.115 ;
        RECT 28.145 187.075 28.405 188.215 ;
        RECT 28.575 187.065 28.905 188.045 ;
        RECT 29.075 187.075 29.355 188.215 ;
        RECT 29.985 187.125 33.495 188.215 ;
        RECT 33.675 187.245 34.005 188.030 ;
        RECT 27.105 186.640 27.390 186.970 ;
        RECT 27.220 186.385 27.390 186.640 ;
        RECT 27.625 186.565 27.955 186.935 ;
        RECT 28.165 186.655 28.500 186.905 ;
        RECT 28.670 186.465 28.840 187.065 ;
        RECT 29.010 186.635 29.345 186.905 ;
        RECT 29.985 186.605 31.675 187.125 ;
        RECT 33.675 187.075 34.355 187.245 ;
        RECT 34.535 187.075 34.865 188.215 ;
        RECT 35.135 187.470 35.405 188.215 ;
        RECT 36.035 188.210 42.310 188.215 ;
        RECT 35.575 187.300 35.865 188.040 ;
        RECT 36.035 187.485 36.290 188.210 ;
        RECT 36.475 187.315 36.735 188.040 ;
        RECT 36.905 187.485 37.150 188.210 ;
        RECT 37.335 187.315 37.595 188.040 ;
        RECT 37.765 187.485 38.010 188.210 ;
        RECT 38.195 187.315 38.455 188.040 ;
        RECT 38.625 187.485 38.870 188.210 ;
        RECT 39.040 187.315 39.300 188.040 ;
        RECT 39.470 187.485 39.730 188.210 ;
        RECT 39.900 187.315 40.160 188.040 ;
        RECT 40.330 187.485 40.590 188.210 ;
        RECT 40.760 187.315 41.020 188.040 ;
        RECT 41.190 187.485 41.450 188.210 ;
        RECT 41.620 187.315 41.880 188.040 ;
        RECT 42.050 187.415 42.310 188.210 ;
        RECT 36.475 187.300 41.880 187.315 ;
        RECT 35.135 187.075 41.880 187.300 ;
        RECT 26.765 185.835 27.025 186.340 ;
        RECT 27.220 186.215 27.885 186.385 ;
        RECT 27.205 185.665 27.535 186.045 ;
        RECT 27.715 185.835 27.885 186.215 ;
        RECT 28.145 185.835 28.840 186.465 ;
        RECT 29.045 185.665 29.355 186.465 ;
        RECT 31.845 186.435 33.495 186.955 ;
        RECT 33.665 186.655 34.015 186.905 ;
        RECT 34.185 186.475 34.355 187.075 ;
        RECT 34.525 186.655 34.875 186.905 ;
        RECT 35.135 186.485 36.300 187.075 ;
        RECT 42.480 186.905 42.730 188.040 ;
        RECT 42.910 187.405 43.170 188.215 ;
        RECT 43.345 186.905 43.590 188.045 ;
        RECT 43.770 187.405 44.065 188.215 ;
        RECT 36.470 186.655 43.590 186.905 ;
        RECT 29.985 185.665 33.495 186.435 ;
        RECT 33.685 185.665 33.925 186.475 ;
        RECT 34.095 185.835 34.425 186.475 ;
        RECT 34.595 185.665 34.865 186.475 ;
        RECT 35.135 186.315 41.880 186.485 ;
        RECT 35.135 185.665 35.435 186.145 ;
        RECT 35.605 185.860 35.865 186.315 ;
        RECT 36.035 185.665 36.295 186.145 ;
        RECT 36.475 185.860 36.735 186.315 ;
        RECT 36.905 185.665 37.155 186.145 ;
        RECT 37.335 185.860 37.595 186.315 ;
        RECT 37.765 185.665 38.015 186.145 ;
        RECT 38.195 185.860 38.455 186.315 ;
        RECT 38.625 185.665 38.870 186.145 ;
        RECT 39.040 185.860 39.315 186.315 ;
        RECT 39.485 185.665 39.730 186.145 ;
        RECT 39.900 185.860 40.160 186.315 ;
        RECT 40.330 185.665 40.590 186.145 ;
        RECT 40.760 185.860 41.020 186.315 ;
        RECT 41.190 185.665 41.450 186.145 ;
        RECT 41.620 185.860 41.880 186.315 ;
        RECT 42.050 185.665 42.310 186.225 ;
        RECT 42.480 185.845 42.730 186.655 ;
        RECT 42.910 185.665 43.170 186.190 ;
        RECT 43.340 185.845 43.590 186.655 ;
        RECT 43.760 186.345 44.075 186.905 ;
        RECT 43.770 185.665 44.075 186.175 ;
        RECT 44.245 185.945 44.525 188.045 ;
        RECT 44.715 187.455 45.500 188.215 ;
        RECT 45.895 187.385 46.280 188.045 ;
        RECT 45.895 187.285 46.305 187.385 ;
        RECT 44.695 187.075 46.305 187.285 ;
        RECT 46.605 187.195 46.805 187.985 ;
        RECT 44.695 186.475 44.970 187.075 ;
        RECT 46.475 187.025 46.805 187.195 ;
        RECT 46.975 187.035 47.295 188.215 ;
        RECT 47.465 187.245 47.735 188.015 ;
        RECT 47.905 187.435 48.235 188.215 ;
        RECT 48.440 187.610 48.625 188.015 ;
        RECT 48.795 187.790 49.130 188.215 ;
        RECT 48.440 187.435 49.105 187.610 ;
        RECT 47.465 187.075 48.595 187.245 ;
        RECT 46.475 186.905 46.655 187.025 ;
        RECT 45.140 186.655 45.495 186.905 ;
        RECT 45.690 186.855 46.155 186.905 ;
        RECT 45.685 186.685 46.155 186.855 ;
        RECT 45.690 186.655 46.155 186.685 ;
        RECT 46.325 186.655 46.655 186.905 ;
        RECT 46.830 186.655 47.295 186.855 ;
        RECT 44.695 186.295 45.945 186.475 ;
        RECT 45.580 186.225 45.945 186.295 ;
        RECT 46.115 186.275 47.295 186.445 ;
        RECT 44.755 185.665 44.925 186.125 ;
        RECT 46.115 186.055 46.445 186.275 ;
        RECT 45.195 185.875 46.445 186.055 ;
        RECT 46.615 185.665 46.785 186.105 ;
        RECT 46.955 185.860 47.295 186.275 ;
        RECT 47.465 186.165 47.635 187.075 ;
        RECT 47.805 186.325 48.165 186.905 ;
        RECT 48.345 186.575 48.595 187.075 ;
        RECT 48.765 186.405 49.105 187.435 ;
        RECT 49.305 187.050 49.595 188.215 ;
        RECT 49.805 187.075 50.035 188.215 ;
        RECT 50.205 187.065 50.535 188.045 ;
        RECT 50.705 187.075 50.915 188.215 ;
        RECT 51.225 187.285 51.405 188.045 ;
        RECT 51.585 187.455 51.915 188.215 ;
        RECT 51.225 187.115 51.900 187.285 ;
        RECT 52.085 187.140 52.355 188.045 ;
        RECT 49.785 186.655 50.115 186.905 ;
        RECT 48.420 186.235 49.105 186.405 ;
        RECT 47.465 185.835 47.725 186.165 ;
        RECT 47.935 185.665 48.210 186.145 ;
        RECT 48.420 185.835 48.625 186.235 ;
        RECT 48.795 185.665 49.130 186.065 ;
        RECT 49.305 185.665 49.595 186.390 ;
        RECT 49.805 185.665 50.035 186.485 ;
        RECT 50.285 186.465 50.535 187.065 ;
        RECT 51.730 186.970 51.900 187.115 ;
        RECT 51.165 186.565 51.505 186.935 ;
        RECT 51.730 186.640 52.005 186.970 ;
        RECT 50.205 185.835 50.535 186.465 ;
        RECT 50.705 185.665 50.915 186.485 ;
        RECT 51.730 186.385 51.900 186.640 ;
        RECT 51.235 186.215 51.900 186.385 ;
        RECT 52.175 186.340 52.355 187.140 ;
        RECT 52.710 187.245 53.100 187.420 ;
        RECT 53.585 187.415 53.915 188.215 ;
        RECT 54.085 187.425 54.620 188.045 ;
        RECT 52.710 187.075 54.135 187.245 ;
        RECT 52.585 186.345 52.940 186.905 ;
        RECT 51.235 185.835 51.405 186.215 ;
        RECT 51.585 185.665 51.915 186.045 ;
        RECT 52.095 185.835 52.355 186.340 ;
        RECT 53.110 186.175 53.280 187.075 ;
        RECT 53.450 186.345 53.715 186.905 ;
        RECT 53.965 186.575 54.135 187.075 ;
        RECT 54.305 186.405 54.620 187.425 ;
        RECT 54.830 187.825 55.165 188.045 ;
        RECT 56.170 187.835 56.525 188.215 ;
        RECT 54.830 187.205 55.085 187.825 ;
        RECT 55.335 187.665 55.565 187.705 ;
        RECT 56.695 187.665 56.945 188.045 ;
        RECT 55.335 187.465 56.945 187.665 ;
        RECT 55.335 187.375 55.520 187.465 ;
        RECT 56.110 187.455 56.945 187.465 ;
        RECT 57.195 187.435 57.445 188.215 ;
        RECT 57.615 187.365 57.875 188.045 ;
        RECT 58.055 187.405 58.350 188.215 ;
        RECT 55.675 187.265 56.005 187.295 ;
        RECT 55.675 187.205 57.475 187.265 ;
        RECT 54.830 187.095 57.535 187.205 ;
        RECT 54.830 187.035 56.005 187.095 ;
        RECT 57.335 187.060 57.535 187.095 ;
        RECT 54.825 186.655 55.315 186.855 ;
        RECT 55.505 186.655 55.980 186.865 ;
        RECT 52.690 185.665 52.930 186.175 ;
        RECT 53.110 185.845 53.390 186.175 ;
        RECT 53.620 185.665 53.835 186.175 ;
        RECT 54.005 185.835 54.620 186.405 ;
        RECT 54.830 185.665 55.285 186.430 ;
        RECT 55.760 186.255 55.980 186.655 ;
        RECT 56.225 186.655 56.555 186.865 ;
        RECT 56.225 186.255 56.435 186.655 ;
        RECT 56.725 186.620 57.135 186.925 ;
        RECT 57.365 186.485 57.535 187.060 ;
        RECT 57.265 186.365 57.535 186.485 ;
        RECT 56.690 186.320 57.535 186.365 ;
        RECT 56.690 186.195 57.445 186.320 ;
        RECT 56.690 186.045 56.860 186.195 ;
        RECT 57.705 186.175 57.875 187.365 ;
        RECT 58.530 186.905 58.775 188.045 ;
        RECT 58.950 187.405 59.210 188.215 ;
        RECT 59.810 188.210 66.085 188.215 ;
        RECT 59.390 186.905 59.640 188.040 ;
        RECT 59.810 187.415 60.070 188.210 ;
        RECT 60.240 187.315 60.500 188.040 ;
        RECT 60.670 187.485 60.930 188.210 ;
        RECT 61.100 187.315 61.360 188.040 ;
        RECT 61.530 187.485 61.790 188.210 ;
        RECT 61.960 187.315 62.220 188.040 ;
        RECT 62.390 187.485 62.650 188.210 ;
        RECT 62.820 187.315 63.080 188.040 ;
        RECT 63.250 187.485 63.495 188.210 ;
        RECT 63.665 187.315 63.925 188.040 ;
        RECT 64.110 187.485 64.355 188.210 ;
        RECT 64.525 187.315 64.785 188.040 ;
        RECT 64.970 187.485 65.215 188.210 ;
        RECT 65.385 187.315 65.645 188.040 ;
        RECT 65.830 187.485 66.085 188.210 ;
        RECT 60.240 187.300 65.645 187.315 ;
        RECT 66.255 187.300 66.545 188.040 ;
        RECT 66.715 187.470 66.985 188.215 ;
        RECT 60.240 187.075 66.985 187.300 ;
        RECT 67.250 187.215 67.505 188.215 ;
        RECT 58.045 186.345 58.360 186.905 ;
        RECT 58.530 186.655 65.650 186.905 ;
        RECT 57.645 186.165 57.875 186.175 ;
        RECT 55.560 185.835 56.860 186.045 ;
        RECT 57.115 185.665 57.445 186.025 ;
        RECT 57.615 185.835 57.875 186.165 ;
        RECT 58.045 185.665 58.350 186.175 ;
        RECT 58.530 185.845 58.780 186.655 ;
        RECT 58.950 185.665 59.210 186.190 ;
        RECT 59.390 185.845 59.640 186.655 ;
        RECT 65.820 186.515 66.985 187.075 ;
        RECT 65.820 186.485 67.015 186.515 ;
        RECT 60.240 186.345 67.015 186.485 ;
        RECT 60.240 186.315 66.985 186.345 ;
        RECT 59.810 185.665 60.070 186.225 ;
        RECT 60.240 185.860 60.500 186.315 ;
        RECT 60.670 185.665 60.930 186.145 ;
        RECT 61.100 185.860 61.360 186.315 ;
        RECT 61.530 185.665 61.790 186.145 ;
        RECT 61.960 185.860 62.220 186.315 ;
        RECT 62.390 185.665 62.635 186.145 ;
        RECT 62.805 185.860 63.080 186.315 ;
        RECT 63.250 185.665 63.495 186.145 ;
        RECT 63.665 185.860 63.925 186.315 ;
        RECT 64.105 185.665 64.355 186.145 ;
        RECT 64.525 185.860 64.785 186.315 ;
        RECT 64.965 185.665 65.215 186.145 ;
        RECT 65.385 185.860 65.645 186.315 ;
        RECT 65.825 185.665 66.085 186.145 ;
        RECT 66.255 185.860 66.515 186.315 ;
        RECT 66.685 185.665 66.985 186.145 ;
        RECT 67.265 185.665 67.505 186.465 ;
        RECT 67.690 185.835 67.935 188.045 ;
        RECT 68.105 187.765 68.955 188.215 ;
        RECT 69.125 187.585 69.385 188.045 ;
        RECT 68.265 187.365 69.385 187.585 ;
        RECT 69.565 187.535 69.770 187.565 ;
        RECT 69.565 187.365 69.775 187.535 ;
        RECT 68.265 186.910 68.435 187.365 ;
        RECT 68.105 186.420 68.435 186.910 ;
        RECT 68.605 186.590 69.015 187.195 ;
        RECT 69.565 186.980 69.770 187.365 ;
        RECT 69.955 187.230 70.280 188.215 ;
        RECT 71.385 187.125 74.895 188.215 ;
        RECT 69.185 186.605 69.770 186.980 ;
        RECT 70.025 186.575 70.285 187.030 ;
        RECT 71.385 186.605 73.075 187.125 ;
        RECT 75.065 187.050 75.355 188.215 ;
        RECT 75.985 187.125 77.655 188.215 ;
        RECT 77.830 187.780 83.175 188.215 ;
        RECT 73.245 186.435 74.895 186.955 ;
        RECT 75.985 186.605 76.735 187.125 ;
        RECT 76.905 186.435 77.655 186.955 ;
        RECT 79.420 186.530 79.770 187.780 ;
        RECT 83.425 187.585 83.605 188.045 ;
        RECT 83.775 187.755 84.025 188.215 ;
        RECT 84.195 187.835 84.525 188.005 ;
        RECT 84.695 187.950 84.950 188.045 ;
        RECT 84.195 187.585 84.365 187.835 ;
        RECT 84.695 187.780 85.835 187.950 ;
        RECT 86.095 187.815 86.425 188.215 ;
        RECT 84.695 187.645 84.950 187.780 ;
        RECT 83.425 187.415 84.365 187.585 ;
        RECT 84.540 187.475 84.950 187.645 ;
        RECT 85.665 187.555 85.835 187.780 ;
        RECT 68.105 186.215 68.955 186.420 ;
        RECT 68.105 185.665 68.435 186.045 ;
        RECT 68.625 185.835 68.955 186.215 ;
        RECT 69.125 186.215 70.280 186.405 ;
        RECT 69.125 186.045 69.335 186.215 ;
        RECT 70.005 186.075 70.280 186.215 ;
        RECT 69.505 185.665 69.835 186.045 ;
        RECT 71.385 185.665 74.895 186.435 ;
        RECT 75.065 185.665 75.355 186.390 ;
        RECT 75.985 185.665 77.655 186.435 ;
        RECT 81.250 186.210 81.590 187.040 ;
        RECT 83.400 186.345 83.660 187.235 ;
        RECT 83.860 186.935 84.340 187.235 ;
        RECT 83.860 186.345 84.120 186.935 ;
        RECT 84.540 186.450 84.710 187.475 ;
        RECT 85.230 187.295 85.400 187.485 ;
        RECT 85.665 187.385 86.425 187.555 ;
        RECT 84.360 186.280 84.710 186.450 ;
        RECT 84.880 187.125 85.400 187.295 ;
        RECT 84.880 186.405 85.050 187.125 ;
        RECT 85.240 186.575 85.530 186.955 ;
        RECT 85.700 186.575 86.030 187.195 ;
        RECT 86.255 186.905 86.425 187.385 ;
        RECT 86.595 187.105 86.855 188.045 ;
        RECT 86.255 186.575 86.510 186.905 ;
        RECT 77.830 185.665 83.175 186.210 ;
        RECT 83.385 185.665 83.785 186.175 ;
        RECT 84.360 185.835 84.530 186.280 ;
        RECT 84.880 186.235 85.760 186.405 ;
        RECT 86.680 186.390 86.855 187.105 ;
        RECT 84.700 185.665 85.420 186.065 ;
        RECT 85.590 185.835 85.760 186.235 ;
        RECT 85.995 185.665 86.425 186.110 ;
        RECT 86.595 185.835 86.855 186.390 ;
        RECT 87.045 187.160 87.350 187.945 ;
        RECT 87.530 187.745 88.215 188.215 ;
        RECT 87.525 187.225 88.220 187.535 ;
        RECT 87.045 186.355 87.220 187.160 ;
        RECT 88.395 187.055 88.680 188.000 ;
        RECT 88.855 187.765 89.185 188.215 ;
        RECT 89.355 187.595 89.525 188.025 ;
        RECT 87.820 186.905 88.680 187.055 ;
        RECT 87.395 186.885 88.680 186.905 ;
        RECT 88.850 187.365 89.525 187.595 ;
        RECT 87.395 186.525 88.380 186.885 ;
        RECT 88.850 186.715 89.085 187.365 ;
        RECT 87.045 185.835 87.285 186.355 ;
        RECT 88.210 186.190 88.380 186.525 ;
        RECT 88.550 186.385 89.085 186.715 ;
        RECT 88.865 186.235 89.085 186.385 ;
        RECT 89.255 186.345 89.555 187.195 ;
        RECT 90.245 187.125 91.915 188.215 ;
        RECT 92.090 187.780 97.435 188.215 ;
        RECT 90.245 186.605 90.995 187.125 ;
        RECT 91.165 186.435 91.915 186.955 ;
        RECT 93.680 186.530 94.030 187.780 ;
        RECT 97.615 187.075 97.945 188.215 ;
        RECT 98.475 187.245 98.805 188.030 ;
        RECT 98.125 187.075 98.805 187.245 ;
        RECT 98.995 187.605 99.325 188.035 ;
        RECT 99.505 187.775 99.700 188.215 ;
        RECT 99.870 187.605 100.200 188.035 ;
        RECT 98.995 187.435 100.200 187.605 ;
        RECT 98.995 187.105 99.890 187.435 ;
        RECT 100.370 187.265 100.645 188.035 ;
        RECT 100.060 187.075 100.645 187.265 ;
        RECT 87.455 185.665 87.850 186.160 ;
        RECT 88.210 185.995 88.585 186.190 ;
        RECT 88.415 185.850 88.585 185.995 ;
        RECT 88.865 185.860 89.105 186.235 ;
        RECT 89.275 185.665 89.610 186.170 ;
        RECT 90.245 185.665 91.915 186.435 ;
        RECT 95.510 186.210 95.850 187.040 ;
        RECT 97.605 186.655 97.955 186.905 ;
        RECT 98.125 186.475 98.295 187.075 ;
        RECT 98.465 186.655 98.815 186.905 ;
        RECT 99.000 186.575 99.295 186.905 ;
        RECT 99.475 186.575 99.890 186.905 ;
        RECT 92.090 185.665 97.435 186.210 ;
        RECT 97.615 185.665 97.885 186.475 ;
        RECT 98.055 185.835 98.385 186.475 ;
        RECT 98.555 185.665 98.795 186.475 ;
        RECT 98.995 185.665 99.295 186.395 ;
        RECT 99.475 185.955 99.705 186.575 ;
        RECT 100.060 186.405 100.235 187.075 ;
        RECT 100.825 187.050 101.115 188.215 ;
        RECT 101.335 187.200 101.590 188.040 ;
        RECT 101.765 187.395 102.095 188.215 ;
        RECT 102.335 187.225 102.545 188.040 ;
        RECT 99.905 186.225 100.235 186.405 ;
        RECT 100.405 186.255 100.645 186.905 ;
        RECT 99.905 185.845 100.130 186.225 ;
        RECT 100.300 185.665 100.630 186.055 ;
        RECT 100.825 185.665 101.115 186.390 ;
        RECT 101.335 185.835 101.665 187.200 ;
        RECT 101.895 187.045 102.545 187.225 ;
        RECT 101.895 186.405 102.115 187.045 ;
        RECT 102.715 186.870 102.920 188.045 ;
        RECT 102.490 186.630 102.920 186.870 ;
        RECT 103.090 186.630 103.420 188.045 ;
        RECT 103.600 186.575 103.880 188.045 ;
        RECT 104.060 187.245 104.345 188.040 ;
        RECT 104.525 187.415 104.740 188.215 ;
        RECT 104.920 187.245 105.190 188.040 ;
        RECT 104.060 187.075 105.190 187.245 ;
        RECT 105.435 187.265 105.710 188.035 ;
        RECT 105.880 187.605 106.210 188.035 ;
        RECT 106.380 187.775 106.575 188.215 ;
        RECT 106.755 187.605 107.085 188.035 ;
        RECT 105.880 187.435 107.085 187.605 ;
        RECT 105.435 187.075 106.020 187.265 ;
        RECT 106.190 187.105 107.085 187.435 ;
        RECT 107.265 187.125 109.855 188.215 ;
        RECT 110.035 187.245 110.365 188.030 ;
        RECT 104.105 186.575 104.490 186.905 ;
        RECT 104.710 186.605 105.210 186.870 ;
        RECT 104.185 186.425 104.490 186.575 ;
        RECT 101.895 186.235 104.005 186.405 ;
        RECT 101.895 186.230 103.115 186.235 ;
        RECT 101.835 185.665 102.510 186.050 ;
        RECT 102.785 185.840 103.115 186.230 ;
        RECT 103.285 185.665 103.630 186.065 ;
        RECT 103.800 185.840 104.005 186.235 ;
        RECT 104.185 185.865 104.740 186.425 ;
        RECT 104.915 185.665 105.155 186.340 ;
        RECT 105.435 186.255 105.675 186.905 ;
        RECT 105.845 186.405 106.020 187.075 ;
        RECT 106.190 186.575 106.605 186.905 ;
        RECT 106.785 186.575 107.080 186.905 ;
        RECT 107.265 186.605 108.475 187.125 ;
        RECT 110.035 187.075 110.715 187.245 ;
        RECT 110.895 187.075 111.225 188.215 ;
        RECT 111.405 187.345 111.680 188.045 ;
        RECT 111.890 187.670 112.105 188.215 ;
        RECT 112.275 187.705 112.750 188.045 ;
        RECT 112.920 187.710 113.535 188.215 ;
        RECT 112.920 187.535 113.115 187.710 ;
        RECT 105.845 186.225 106.175 186.405 ;
        RECT 105.450 185.665 105.780 186.055 ;
        RECT 105.950 185.845 106.175 186.225 ;
        RECT 106.375 185.955 106.605 186.575 ;
        RECT 108.645 186.435 109.855 186.955 ;
        RECT 110.025 186.655 110.375 186.905 ;
        RECT 110.545 186.475 110.715 187.075 ;
        RECT 110.885 186.655 111.235 186.905 ;
        RECT 106.785 185.665 107.085 186.395 ;
        RECT 107.265 185.665 109.855 186.435 ;
        RECT 110.045 185.665 110.285 186.475 ;
        RECT 110.455 185.835 110.785 186.475 ;
        RECT 110.955 185.665 111.225 186.475 ;
        RECT 111.405 186.315 111.575 187.345 ;
        RECT 111.850 187.175 112.565 187.470 ;
        RECT 112.785 187.345 113.115 187.535 ;
        RECT 113.285 187.175 113.535 187.540 ;
        RECT 111.745 187.005 113.535 187.175 ;
        RECT 111.745 186.575 111.975 187.005 ;
        RECT 111.405 185.835 111.665 186.315 ;
        RECT 112.145 186.305 112.555 186.825 ;
        RECT 111.835 185.665 112.165 186.125 ;
        RECT 112.355 185.885 112.555 186.305 ;
        RECT 112.725 186.150 112.980 187.005 ;
        RECT 113.775 186.825 113.945 188.045 ;
        RECT 114.195 187.705 114.455 188.215 ;
        RECT 113.150 186.575 113.945 186.825 ;
        RECT 114.115 186.655 114.455 187.535 ;
        RECT 114.625 187.125 118.135 188.215 ;
        RECT 118.310 187.780 123.655 188.215 ;
        RECT 114.625 186.605 116.315 187.125 ;
        RECT 113.695 186.485 113.945 186.575 ;
        RECT 112.725 185.885 113.515 186.150 ;
        RECT 113.695 186.065 114.025 186.485 ;
        RECT 114.195 185.665 114.455 186.485 ;
        RECT 116.485 186.435 118.135 186.955 ;
        RECT 119.900 186.530 120.250 187.780 ;
        RECT 123.915 187.285 124.085 188.045 ;
        RECT 124.300 187.455 124.630 188.215 ;
        RECT 123.915 187.115 124.630 187.285 ;
        RECT 124.800 187.140 125.055 188.045 ;
        RECT 114.625 185.665 118.135 186.435 ;
        RECT 121.730 186.210 122.070 187.040 ;
        RECT 123.825 186.565 124.180 186.935 ;
        RECT 124.460 186.905 124.630 187.115 ;
        RECT 124.460 186.575 124.715 186.905 ;
        RECT 124.460 186.385 124.630 186.575 ;
        RECT 124.885 186.410 125.055 187.140 ;
        RECT 125.230 187.065 125.490 188.215 ;
        RECT 125.665 187.125 126.875 188.215 ;
        RECT 125.665 186.585 126.185 187.125 ;
        RECT 123.915 186.215 124.630 186.385 ;
        RECT 118.310 185.665 123.655 186.210 ;
        RECT 123.915 185.835 124.085 186.215 ;
        RECT 124.300 185.665 124.630 186.045 ;
        RECT 124.800 185.835 125.055 186.410 ;
        RECT 125.230 185.665 125.490 186.505 ;
        RECT 126.355 186.415 126.875 186.955 ;
        RECT 125.665 185.665 126.875 186.415 ;
        RECT 14.260 185.495 126.960 185.665 ;
        RECT 14.345 184.745 15.555 185.495 ;
        RECT 16.275 184.945 16.445 185.325 ;
        RECT 16.625 185.115 16.955 185.495 ;
        RECT 16.275 184.775 16.940 184.945 ;
        RECT 17.135 184.820 17.395 185.325 ;
        RECT 18.115 185.015 18.415 185.495 ;
        RECT 18.585 184.845 18.845 185.300 ;
        RECT 19.015 185.015 19.275 185.495 ;
        RECT 19.455 184.845 19.715 185.300 ;
        RECT 19.885 185.015 20.135 185.495 ;
        RECT 20.315 184.845 20.575 185.300 ;
        RECT 20.745 185.015 20.995 185.495 ;
        RECT 21.175 184.845 21.435 185.300 ;
        RECT 21.605 185.015 21.850 185.495 ;
        RECT 22.020 184.845 22.295 185.300 ;
        RECT 22.465 185.015 22.710 185.495 ;
        RECT 22.880 184.845 23.140 185.300 ;
        RECT 23.310 185.015 23.570 185.495 ;
        RECT 23.740 184.845 24.000 185.300 ;
        RECT 24.170 185.015 24.430 185.495 ;
        RECT 24.600 184.845 24.860 185.300 ;
        RECT 25.030 184.935 25.290 185.495 ;
        RECT 14.345 184.205 14.865 184.745 ;
        RECT 15.035 184.035 15.555 184.575 ;
        RECT 16.205 184.225 16.535 184.595 ;
        RECT 16.770 184.520 16.940 184.775 ;
        RECT 16.770 184.190 17.055 184.520 ;
        RECT 16.770 184.045 16.940 184.190 ;
        RECT 14.345 182.945 15.555 184.035 ;
        RECT 16.275 183.875 16.940 184.045 ;
        RECT 17.225 184.020 17.395 184.820 ;
        RECT 16.275 183.115 16.445 183.875 ;
        RECT 16.625 182.945 16.955 183.705 ;
        RECT 17.125 183.115 17.395 184.020 ;
        RECT 18.115 184.675 24.860 184.845 ;
        RECT 18.115 184.085 19.280 184.675 ;
        RECT 25.460 184.505 25.710 185.315 ;
        RECT 25.890 184.970 26.150 185.495 ;
        RECT 26.320 184.505 26.570 185.315 ;
        RECT 26.750 184.985 27.055 185.495 ;
        RECT 27.225 184.985 27.530 185.495 ;
        RECT 19.450 184.255 26.570 184.505 ;
        RECT 26.740 184.255 27.055 184.815 ;
        RECT 27.225 184.255 27.540 184.815 ;
        RECT 27.710 184.505 27.960 185.315 ;
        RECT 28.130 184.970 28.390 185.495 ;
        RECT 28.570 184.505 28.820 185.315 ;
        RECT 28.990 184.935 29.250 185.495 ;
        RECT 29.420 184.845 29.680 185.300 ;
        RECT 29.850 185.015 30.110 185.495 ;
        RECT 30.280 184.845 30.540 185.300 ;
        RECT 30.710 185.015 30.970 185.495 ;
        RECT 31.140 184.845 31.400 185.300 ;
        RECT 31.570 185.015 31.815 185.495 ;
        RECT 31.985 184.845 32.260 185.300 ;
        RECT 32.430 185.015 32.675 185.495 ;
        RECT 32.845 184.845 33.105 185.300 ;
        RECT 33.285 185.015 33.535 185.495 ;
        RECT 33.705 184.845 33.965 185.300 ;
        RECT 34.145 185.015 34.395 185.495 ;
        RECT 34.565 184.845 34.825 185.300 ;
        RECT 35.005 185.015 35.265 185.495 ;
        RECT 35.435 184.845 35.695 185.300 ;
        RECT 35.865 185.015 36.165 185.495 ;
        RECT 29.420 184.675 36.165 184.845 ;
        RECT 36.425 184.770 36.715 185.495 ;
        RECT 36.895 184.770 37.225 185.495 ;
        RECT 37.415 185.240 37.745 185.285 ;
        RECT 37.410 184.775 37.745 185.240 ;
        RECT 27.710 184.255 34.830 184.505 ;
        RECT 18.115 183.860 24.860 184.085 ;
        RECT 18.115 182.945 18.385 183.690 ;
        RECT 18.555 183.120 18.845 183.860 ;
        RECT 19.455 183.845 24.860 183.860 ;
        RECT 19.015 182.950 19.270 183.675 ;
        RECT 19.455 183.120 19.715 183.845 ;
        RECT 19.885 182.950 20.130 183.675 ;
        RECT 20.315 183.120 20.575 183.845 ;
        RECT 20.745 182.950 20.990 183.675 ;
        RECT 21.175 183.120 21.435 183.845 ;
        RECT 21.605 182.950 21.850 183.675 ;
        RECT 22.020 183.120 22.280 183.845 ;
        RECT 22.450 182.950 22.710 183.675 ;
        RECT 22.880 183.120 23.140 183.845 ;
        RECT 23.310 182.950 23.570 183.675 ;
        RECT 23.740 183.120 24.000 183.845 ;
        RECT 24.170 182.950 24.430 183.675 ;
        RECT 24.600 183.120 24.860 183.845 ;
        RECT 25.030 182.950 25.290 183.745 ;
        RECT 25.460 183.120 25.710 184.255 ;
        RECT 19.015 182.945 25.290 182.950 ;
        RECT 25.890 182.945 26.150 183.755 ;
        RECT 26.325 183.115 26.570 184.255 ;
        RECT 26.750 182.945 27.045 183.755 ;
        RECT 27.235 182.945 27.530 183.755 ;
        RECT 27.710 183.115 27.955 184.255 ;
        RECT 28.130 182.945 28.390 183.755 ;
        RECT 28.570 183.120 28.820 184.255 ;
        RECT 35.000 184.085 36.165 184.675 ;
        RECT 29.420 183.860 36.165 184.085 ;
        RECT 29.420 183.845 34.825 183.860 ;
        RECT 28.990 182.950 29.250 183.745 ;
        RECT 29.420 183.120 29.680 183.845 ;
        RECT 29.850 182.950 30.110 183.675 ;
        RECT 30.280 183.120 30.540 183.845 ;
        RECT 30.710 182.950 30.970 183.675 ;
        RECT 31.140 183.120 31.400 183.845 ;
        RECT 31.570 182.950 31.830 183.675 ;
        RECT 32.000 183.120 32.260 183.845 ;
        RECT 32.430 182.950 32.675 183.675 ;
        RECT 32.845 183.120 33.105 183.845 ;
        RECT 33.290 182.950 33.535 183.675 ;
        RECT 33.705 183.120 33.965 183.845 ;
        RECT 34.150 182.950 34.395 183.675 ;
        RECT 34.565 183.120 34.825 183.845 ;
        RECT 35.010 182.950 35.265 183.675 ;
        RECT 35.435 183.120 35.725 183.860 ;
        RECT 28.990 182.945 35.265 182.950 ;
        RECT 35.895 182.945 36.165 183.690 ;
        RECT 36.425 182.945 36.715 184.110 ;
        RECT 37.410 184.085 37.585 184.775 ;
        RECT 37.915 184.690 38.150 185.495 ;
        RECT 37.755 184.265 38.150 184.505 ;
        RECT 37.925 184.085 38.150 184.265 ;
        RECT 38.320 184.255 38.580 185.165 ;
        RECT 38.760 184.275 39.060 185.165 ;
        RECT 38.890 184.255 39.060 184.275 ;
        RECT 39.235 184.255 39.590 185.160 ;
        RECT 39.810 184.995 40.305 185.325 ;
        RECT 40.565 184.995 40.825 185.325 ;
        RECT 40.995 185.135 41.325 185.495 ;
        RECT 41.580 185.115 42.880 185.325 ;
        RECT 39.810 184.085 39.980 184.995 ;
        RECT 40.565 184.985 40.795 184.995 ;
        RECT 36.905 182.945 37.235 183.745 ;
        RECT 37.410 183.455 37.745 184.085 ;
        RECT 37.925 183.915 39.980 184.085 ;
        RECT 37.405 183.285 37.745 183.455 ;
        RECT 37.410 183.115 37.745 183.285 ;
        RECT 37.915 182.945 38.245 183.745 ;
        RECT 38.645 183.115 38.895 183.915 ;
        RECT 39.080 182.945 39.410 183.665 ;
        RECT 39.630 183.115 39.880 183.915 ;
        RECT 40.150 183.505 40.355 184.825 ;
        RECT 40.565 183.795 40.735 184.985 ;
        RECT 41.580 184.965 41.750 185.115 ;
        RECT 40.995 184.840 41.750 184.965 ;
        RECT 40.905 184.795 41.750 184.840 ;
        RECT 40.905 184.675 41.175 184.795 ;
        RECT 40.905 184.100 41.075 184.675 ;
        RECT 41.305 184.235 41.715 184.540 ;
        RECT 42.005 184.505 42.215 184.905 ;
        RECT 41.885 184.295 42.215 184.505 ;
        RECT 42.460 184.505 42.680 184.905 ;
        RECT 43.155 184.730 43.610 185.495 ;
        RECT 43.785 184.995 44.085 185.325 ;
        RECT 44.255 185.015 44.530 185.495 ;
        RECT 42.460 184.295 42.935 184.505 ;
        RECT 43.125 184.305 43.615 184.505 ;
        RECT 40.905 184.065 41.105 184.100 ;
        RECT 42.435 184.065 43.610 184.125 ;
        RECT 40.905 183.955 43.610 184.065 ;
        RECT 40.965 183.895 42.765 183.955 ;
        RECT 42.435 183.865 42.765 183.895 ;
        RECT 40.055 182.945 40.385 183.325 ;
        RECT 40.565 183.115 40.825 183.795 ;
        RECT 40.995 182.945 41.245 183.725 ;
        RECT 41.495 183.695 42.330 183.705 ;
        RECT 42.920 183.695 43.105 183.785 ;
        RECT 41.495 183.495 43.105 183.695 ;
        RECT 41.495 183.115 41.745 183.495 ;
        RECT 42.875 183.455 43.105 183.495 ;
        RECT 43.355 183.335 43.610 183.955 ;
        RECT 41.915 182.945 42.270 183.325 ;
        RECT 43.275 183.115 43.610 183.335 ;
        RECT 43.785 184.085 43.955 184.995 ;
        RECT 44.710 184.845 45.005 185.235 ;
        RECT 45.175 185.015 45.430 185.495 ;
        RECT 45.605 184.845 45.865 185.235 ;
        RECT 46.035 185.015 46.315 185.495 ;
        RECT 46.555 184.845 46.885 185.310 ;
        RECT 47.055 185.025 47.225 185.495 ;
        RECT 47.400 185.095 47.730 185.325 ;
        RECT 47.935 185.155 48.105 185.325 ;
        RECT 47.480 184.845 47.650 185.095 ;
        RECT 47.935 184.985 48.155 185.155 ;
        RECT 47.935 184.935 48.105 184.985 ;
        RECT 44.125 184.255 44.475 184.825 ;
        RECT 44.710 184.675 46.360 184.845 ;
        RECT 46.555 184.675 47.650 184.845 ;
        RECT 47.865 184.755 48.105 184.935 ;
        RECT 48.450 184.925 48.640 185.085 ;
        RECT 48.330 184.755 48.640 184.925 ;
        RECT 48.860 184.755 49.135 185.495 ;
        RECT 50.425 184.865 50.755 185.225 ;
        RECT 51.375 185.035 51.625 185.495 ;
        RECT 51.795 185.035 52.355 185.325 ;
        RECT 44.645 184.335 45.785 184.505 ;
        RECT 44.645 184.085 44.815 184.335 ;
        RECT 45.955 184.165 46.360 184.675 ;
        RECT 46.545 184.295 47.025 184.505 ;
        RECT 47.195 184.295 47.695 184.505 ;
        RECT 43.785 183.915 44.815 184.085 ;
        RECT 45.605 183.995 46.360 184.165 ;
        RECT 47.865 184.125 48.035 184.755 ;
        RECT 48.330 184.585 48.500 184.755 ;
        RECT 50.425 184.675 51.815 184.865 ;
        RECT 51.645 184.585 51.815 184.675 ;
        RECT 43.785 183.115 44.095 183.915 ;
        RECT 45.605 183.745 45.865 183.995 ;
        RECT 44.265 182.945 44.575 183.745 ;
        RECT 44.745 183.575 45.865 183.745 ;
        RECT 44.745 183.115 45.005 183.575 ;
        RECT 45.175 182.945 45.430 183.405 ;
        RECT 45.605 183.115 45.865 183.575 ;
        RECT 46.035 182.945 46.320 183.815 ;
        RECT 46.575 182.945 46.950 184.045 ;
        RECT 47.425 183.955 48.035 184.125 ;
        RECT 48.205 184.045 48.500 184.585 ;
        RECT 48.685 184.235 49.135 184.585 ;
        RECT 47.425 183.115 47.750 183.955 ;
        RECT 48.205 183.875 48.695 184.045 ;
        RECT 47.920 182.945 48.250 183.705 ;
        RECT 48.420 183.370 48.695 183.875 ;
        RECT 48.865 183.135 49.135 184.235 ;
        RECT 50.240 184.255 50.915 184.505 ;
        RECT 51.135 184.255 51.475 184.505 ;
        RECT 51.645 184.255 51.935 184.585 ;
        RECT 50.240 183.895 50.505 184.255 ;
        RECT 51.645 184.005 51.815 184.255 ;
        RECT 50.875 183.835 51.815 184.005 ;
        RECT 50.425 182.945 50.705 183.615 ;
        RECT 50.875 183.285 51.175 183.835 ;
        RECT 52.105 183.665 52.355 185.035 ;
        RECT 52.525 185.005 52.795 185.495 ;
        RECT 52.585 184.255 52.850 184.835 ;
        RECT 53.020 184.565 53.295 185.275 ;
        RECT 53.495 185.010 54.280 185.275 ;
        RECT 53.020 184.335 53.855 184.565 ;
        RECT 51.375 182.945 51.705 183.665 ;
        RECT 51.895 183.115 52.355 183.665 ;
        RECT 52.525 182.945 52.840 184.005 ;
        RECT 53.020 183.675 53.295 184.335 ;
        RECT 54.025 184.155 54.280 185.010 ;
        RECT 54.450 184.815 54.660 185.275 ;
        RECT 54.850 185.000 55.180 185.495 ;
        RECT 55.355 184.865 55.600 185.325 ;
        RECT 54.450 184.335 54.860 184.815 ;
        RECT 55.430 184.655 55.600 184.865 ;
        RECT 55.770 184.835 56.035 185.495 ;
        RECT 56.205 184.820 56.465 185.325 ;
        RECT 56.645 185.115 56.975 185.495 ;
        RECT 57.155 184.945 57.325 185.325 ;
        RECT 55.030 184.155 55.260 184.585 ;
        RECT 53.490 183.985 55.260 184.155 ;
        RECT 55.430 184.135 56.035 184.655 ;
        RECT 53.490 183.620 53.725 183.985 ;
        RECT 53.895 183.625 54.225 183.815 ;
        RECT 54.450 183.690 54.640 183.985 ;
        RECT 53.895 183.450 54.085 183.625 ;
        RECT 53.470 182.945 54.085 183.450 ;
        RECT 54.255 183.115 54.730 183.455 ;
        RECT 54.900 182.945 55.115 183.790 ;
        RECT 55.430 183.785 55.600 184.135 ;
        RECT 56.205 184.020 56.375 184.820 ;
        RECT 56.660 184.775 57.325 184.945 ;
        RECT 56.660 184.520 56.830 184.775 ;
        RECT 56.545 184.190 56.830 184.520 ;
        RECT 57.065 184.225 57.395 184.595 ;
        RECT 56.660 184.045 56.830 184.190 ;
        RECT 55.315 183.115 55.600 183.785 ;
        RECT 55.770 182.945 56.035 183.955 ;
        RECT 56.205 183.115 56.475 184.020 ;
        RECT 56.660 183.875 57.325 184.045 ;
        RECT 56.645 182.945 56.975 183.705 ;
        RECT 57.155 183.115 57.325 183.875 ;
        RECT 57.585 183.115 58.335 185.325 ;
        RECT 58.515 184.775 58.845 185.495 ;
        RECT 59.390 185.095 61.005 185.265 ;
        RECT 61.175 185.095 61.505 185.495 ;
        RECT 60.835 184.925 61.005 185.095 ;
        RECT 61.675 185.020 62.010 185.280 ;
        RECT 58.570 184.255 58.920 184.585 ;
        RECT 59.230 184.255 59.650 184.920 ;
        RECT 59.820 184.475 60.110 184.915 ;
        RECT 60.300 184.815 60.570 184.915 ;
        RECT 60.300 184.645 60.575 184.815 ;
        RECT 60.835 184.755 61.395 184.925 ;
        RECT 59.820 184.305 60.115 184.475 ;
        RECT 59.820 184.255 60.110 184.305 ;
        RECT 60.300 184.255 60.570 184.645 ;
        RECT 61.225 184.585 61.395 184.755 ;
        RECT 60.780 184.475 61.030 184.585 ;
        RECT 60.780 184.305 61.035 184.475 ;
        RECT 60.780 184.255 61.030 184.305 ;
        RECT 61.225 184.255 61.530 184.585 ;
        RECT 58.570 184.135 58.775 184.255 ;
        RECT 58.565 183.965 58.775 184.135 ;
        RECT 61.225 184.085 61.395 184.255 ;
        RECT 59.025 183.915 61.395 184.085 ;
        RECT 58.595 183.285 58.765 183.785 ;
        RECT 59.025 183.455 59.195 183.915 ;
        RECT 59.425 183.535 60.850 183.705 ;
        RECT 59.425 183.285 59.755 183.535 ;
        RECT 58.595 183.115 59.755 183.285 ;
        RECT 59.980 182.945 60.310 183.365 ;
        RECT 60.565 183.115 60.850 183.535 ;
        RECT 61.095 182.945 61.425 183.745 ;
        RECT 61.755 183.665 62.010 185.020 ;
        RECT 62.185 184.770 62.475 185.495 ;
        RECT 63.565 184.695 63.875 185.495 ;
        RECT 64.080 184.695 64.775 185.325 ;
        RECT 64.945 184.755 65.435 185.325 ;
        RECT 65.605 184.925 65.835 185.325 ;
        RECT 66.005 185.095 66.425 185.495 ;
        RECT 66.595 184.925 66.765 185.325 ;
        RECT 65.605 184.755 66.765 184.925 ;
        RECT 66.935 184.755 67.385 185.495 ;
        RECT 67.555 184.755 67.995 185.315 ;
        RECT 63.575 184.255 63.910 184.525 ;
        RECT 64.080 184.135 64.250 184.695 ;
        RECT 64.420 184.255 64.755 184.505 ;
        RECT 61.675 183.155 62.010 183.665 ;
        RECT 62.185 182.945 62.475 184.110 ;
        RECT 64.080 184.095 64.255 184.135 ;
        RECT 63.565 182.945 63.845 184.085 ;
        RECT 64.015 183.115 64.345 184.095 ;
        RECT 64.945 184.085 65.115 184.755 ;
        RECT 65.285 184.255 65.690 184.585 ;
        RECT 64.515 182.945 64.775 184.085 ;
        RECT 64.945 183.915 65.715 184.085 ;
        RECT 64.955 182.945 65.285 183.745 ;
        RECT 65.465 183.285 65.715 183.915 ;
        RECT 65.905 183.455 66.155 184.585 ;
        RECT 66.355 184.255 66.600 184.585 ;
        RECT 66.785 184.305 67.175 184.585 ;
        RECT 66.355 183.455 66.555 184.255 ;
        RECT 67.345 184.135 67.515 184.585 ;
        RECT 66.725 183.965 67.515 184.135 ;
        RECT 66.725 183.285 66.895 183.965 ;
        RECT 65.465 183.115 66.895 183.285 ;
        RECT 67.065 182.945 67.380 183.795 ;
        RECT 67.685 183.745 67.995 184.755 ;
        RECT 68.165 184.755 68.655 185.325 ;
        RECT 68.825 184.925 69.055 185.325 ;
        RECT 69.225 185.095 69.645 185.495 ;
        RECT 69.815 184.925 69.985 185.325 ;
        RECT 68.825 184.755 69.985 184.925 ;
        RECT 70.155 184.755 70.605 185.495 ;
        RECT 70.775 184.755 71.215 185.315 ;
        RECT 68.165 184.085 68.335 184.755 ;
        RECT 68.505 184.255 68.910 184.585 ;
        RECT 68.165 183.915 68.935 184.085 ;
        RECT 67.555 183.115 67.995 183.745 ;
        RECT 68.175 182.945 68.505 183.745 ;
        RECT 68.685 183.285 68.935 183.915 ;
        RECT 69.125 183.455 69.375 184.585 ;
        RECT 69.575 184.255 69.820 184.585 ;
        RECT 70.005 184.305 70.395 184.585 ;
        RECT 69.575 183.455 69.775 184.255 ;
        RECT 70.565 184.135 70.735 184.585 ;
        RECT 69.945 183.965 70.735 184.135 ;
        RECT 69.945 183.285 70.115 183.965 ;
        RECT 68.685 183.115 70.115 183.285 ;
        RECT 70.285 182.945 70.600 183.795 ;
        RECT 70.905 183.745 71.215 184.755 ;
        RECT 71.475 184.625 71.645 185.190 ;
        RECT 71.835 184.965 72.065 185.270 ;
        RECT 72.235 185.135 72.565 185.495 ;
        RECT 72.760 184.965 73.050 185.315 ;
        RECT 71.835 184.795 73.050 184.965 ;
        RECT 73.225 184.725 74.895 185.495 ;
        RECT 75.070 184.950 80.415 185.495 ;
        RECT 71.475 184.455 71.995 184.625 ;
        RECT 71.390 183.925 71.635 184.285 ;
        RECT 71.825 184.075 71.995 184.455 ;
        RECT 72.165 184.255 72.550 184.585 ;
        RECT 72.730 184.475 72.990 184.585 ;
        RECT 72.730 184.305 72.995 184.475 ;
        RECT 72.730 184.255 72.990 184.305 ;
        RECT 71.825 183.795 72.175 184.075 ;
        RECT 70.775 183.115 71.215 183.745 ;
        RECT 71.390 182.945 71.645 183.745 ;
        RECT 71.845 183.115 72.175 183.795 ;
        RECT 72.355 183.205 72.550 184.255 ;
        RECT 72.730 182.945 73.050 184.085 ;
        RECT 73.225 184.035 73.975 184.555 ;
        RECT 74.145 184.205 74.895 184.725 ;
        RECT 73.225 182.945 74.895 184.035 ;
        RECT 76.660 183.380 77.010 184.630 ;
        RECT 78.490 184.120 78.830 184.950 ;
        RECT 80.675 184.845 80.845 185.325 ;
        RECT 81.015 185.015 81.345 185.495 ;
        RECT 81.570 185.075 83.105 185.325 ;
        RECT 81.570 184.845 81.740 185.075 ;
        RECT 80.675 184.675 81.740 184.845 ;
        RECT 81.920 184.505 82.200 184.905 ;
        RECT 80.590 184.295 80.940 184.505 ;
        RECT 81.110 184.305 81.555 184.505 ;
        RECT 81.725 184.305 82.200 184.505 ;
        RECT 82.470 184.505 82.755 184.905 ;
        RECT 82.935 184.845 83.105 185.075 ;
        RECT 83.275 185.015 83.605 185.495 ;
        RECT 83.820 184.995 84.075 185.325 ;
        RECT 83.865 184.985 84.075 184.995 ;
        RECT 83.890 184.915 84.075 184.985 ;
        RECT 82.935 184.675 83.735 184.845 ;
        RECT 82.470 184.305 82.800 184.505 ;
        RECT 82.970 184.305 83.335 184.505 ;
        RECT 83.565 184.125 83.735 184.675 ;
        RECT 80.675 183.955 83.735 184.125 ;
        RECT 75.070 182.945 80.415 183.380 ;
        RECT 80.675 183.115 80.845 183.955 ;
        RECT 83.905 183.785 84.075 184.915 ;
        RECT 84.275 184.775 84.605 185.495 ;
        RECT 85.150 185.095 86.765 185.265 ;
        RECT 86.935 185.095 87.265 185.495 ;
        RECT 86.595 184.925 86.765 185.095 ;
        RECT 87.435 185.020 87.770 185.280 ;
        RECT 84.330 184.255 84.680 184.585 ;
        RECT 84.990 184.255 85.410 184.920 ;
        RECT 85.580 184.255 85.870 184.915 ;
        RECT 86.060 184.815 86.330 184.915 ;
        RECT 86.060 184.645 86.335 184.815 ;
        RECT 86.595 184.755 87.155 184.925 ;
        RECT 86.060 184.255 86.330 184.645 ;
        RECT 86.985 184.585 87.155 184.755 ;
        RECT 86.540 184.475 86.790 184.585 ;
        RECT 86.540 184.305 86.795 184.475 ;
        RECT 86.540 184.255 86.790 184.305 ;
        RECT 86.985 184.255 87.290 184.585 ;
        RECT 84.330 184.135 84.535 184.255 ;
        RECT 84.325 183.965 84.535 184.135 ;
        RECT 86.985 184.085 87.155 184.255 ;
        RECT 84.785 183.915 87.155 184.085 ;
        RECT 81.015 183.285 81.345 183.785 ;
        RECT 81.515 183.545 83.150 183.785 ;
        RECT 81.515 183.455 81.745 183.545 ;
        RECT 81.855 183.285 82.185 183.325 ;
        RECT 81.015 183.115 82.185 183.285 ;
        RECT 82.375 182.945 82.730 183.365 ;
        RECT 82.900 183.115 83.150 183.545 ;
        RECT 83.320 182.945 83.650 183.705 ;
        RECT 83.820 183.115 84.075 183.785 ;
        RECT 84.355 183.285 84.525 183.785 ;
        RECT 84.785 183.455 84.955 183.915 ;
        RECT 85.185 183.535 86.610 183.705 ;
        RECT 85.185 183.285 85.515 183.535 ;
        RECT 84.355 183.115 85.515 183.285 ;
        RECT 85.740 182.945 86.070 183.365 ;
        RECT 86.325 183.115 86.610 183.535 ;
        RECT 86.855 182.945 87.185 183.745 ;
        RECT 87.515 183.665 87.770 185.020 ;
        RECT 87.945 184.770 88.235 185.495 ;
        RECT 88.430 185.105 88.760 185.495 ;
        RECT 88.930 184.935 89.155 185.315 ;
        RECT 88.415 184.255 88.655 184.905 ;
        RECT 88.825 184.755 89.155 184.935 ;
        RECT 87.435 183.155 87.770 183.665 ;
        RECT 87.945 182.945 88.235 184.110 ;
        RECT 88.825 184.085 89.000 184.755 ;
        RECT 89.355 184.585 89.585 185.205 ;
        RECT 89.765 184.765 90.065 185.495 ;
        RECT 90.265 184.985 90.505 185.495 ;
        RECT 90.675 184.985 90.965 185.325 ;
        RECT 91.195 184.985 91.510 185.495 ;
        RECT 90.305 184.645 90.505 184.815 ;
        RECT 89.170 184.255 89.585 184.585 ;
        RECT 89.765 184.255 90.060 184.585 ;
        RECT 90.310 184.255 90.505 184.645 ;
        RECT 90.675 184.085 90.855 184.985 ;
        RECT 91.680 184.925 91.850 185.195 ;
        RECT 92.020 185.095 92.350 185.495 ;
        RECT 91.025 184.255 91.435 184.815 ;
        RECT 91.680 184.755 92.375 184.925 ;
        RECT 91.605 184.085 91.775 184.585 ;
        RECT 88.415 183.895 89.000 184.085 ;
        RECT 88.415 183.125 88.690 183.895 ;
        RECT 89.170 183.725 90.065 184.055 ;
        RECT 90.315 183.915 91.775 184.085 ;
        RECT 90.315 183.740 90.675 183.915 ;
        RECT 91.945 183.745 92.375 184.755 ;
        RECT 92.635 184.625 92.805 185.190 ;
        RECT 92.995 184.965 93.225 185.270 ;
        RECT 93.395 185.135 93.725 185.495 ;
        RECT 93.920 184.965 94.210 185.315 ;
        RECT 92.995 184.795 94.210 184.965 ;
        RECT 94.585 184.865 94.915 185.225 ;
        RECT 95.535 185.035 95.785 185.495 ;
        RECT 95.955 185.035 96.515 185.325 ;
        RECT 94.585 184.675 95.975 184.865 ;
        RECT 92.635 184.455 93.155 184.625 ;
        RECT 95.805 184.585 95.975 184.675 ;
        RECT 92.550 183.925 92.795 184.285 ;
        RECT 92.985 184.075 93.155 184.455 ;
        RECT 93.325 184.255 93.710 184.585 ;
        RECT 93.890 184.475 94.150 184.585 ;
        RECT 93.890 184.305 94.155 184.475 ;
        RECT 93.890 184.255 94.150 184.305 ;
        RECT 94.400 184.255 95.075 184.505 ;
        RECT 95.295 184.255 95.635 184.505 ;
        RECT 95.805 184.255 96.095 184.585 ;
        RECT 92.985 183.795 93.335 184.075 ;
        RECT 88.860 183.555 90.065 183.725 ;
        RECT 88.860 183.125 89.190 183.555 ;
        RECT 89.360 182.945 89.555 183.385 ;
        RECT 89.735 183.125 90.065 183.555 ;
        RECT 91.260 182.945 91.430 183.745 ;
        RECT 91.600 183.575 92.375 183.745 ;
        RECT 91.600 183.115 91.930 183.575 ;
        RECT 92.100 182.945 92.270 183.405 ;
        RECT 92.550 182.945 92.805 183.745 ;
        RECT 93.005 183.115 93.335 183.795 ;
        RECT 93.515 183.205 93.710 184.255 ;
        RECT 93.890 182.945 94.210 184.085 ;
        RECT 94.400 183.895 94.665 184.255 ;
        RECT 95.805 184.005 95.975 184.255 ;
        RECT 95.035 183.835 95.975 184.005 ;
        RECT 94.585 182.945 94.865 183.615 ;
        RECT 95.035 183.285 95.335 183.835 ;
        RECT 96.265 183.665 96.515 185.035 ;
        RECT 97.145 184.695 97.455 185.495 ;
        RECT 97.660 184.695 98.355 185.325 ;
        RECT 98.525 185.115 99.910 185.325 ;
        RECT 98.525 184.845 98.815 185.115 ;
        RECT 98.985 184.755 99.410 184.945 ;
        RECT 99.580 184.925 99.910 185.115 ;
        RECT 100.145 185.095 100.475 185.495 ;
        RECT 100.650 184.925 100.980 185.325 ;
        RECT 101.185 184.935 101.355 185.495 ;
        RECT 99.580 184.755 100.980 184.925 ;
        RECT 101.525 184.755 102.035 185.325 ;
        RECT 97.155 184.255 97.490 184.525 ;
        RECT 97.660 184.095 97.830 184.695 ;
        RECT 98.000 184.255 98.335 184.505 ;
        RECT 98.525 184.255 98.800 184.585 ;
        RECT 95.535 182.945 95.865 183.665 ;
        RECT 96.055 183.115 96.515 183.665 ;
        RECT 97.145 182.945 97.425 184.085 ;
        RECT 97.595 183.115 97.925 184.095 ;
        RECT 98.095 182.945 98.355 184.085 ;
        RECT 98.525 182.945 98.815 184.085 ;
        RECT 98.985 183.745 99.155 184.755 ;
        RECT 99.325 183.920 99.680 184.585 ;
        RECT 99.865 183.920 100.140 184.585 ;
        RECT 100.310 184.255 100.655 184.585 ;
        RECT 100.945 184.505 101.115 184.585 ;
        RECT 101.485 184.505 101.675 184.585 ;
        RECT 100.865 184.255 101.115 184.505 ;
        RECT 101.310 184.255 101.675 184.505 ;
        RECT 98.985 183.495 99.940 183.745 ;
        RECT 99.610 183.285 99.940 183.495 ;
        RECT 100.310 183.455 100.635 184.255 ;
        RECT 101.310 184.085 101.480 184.255 ;
        RECT 101.860 184.085 102.035 184.755 ;
        RECT 102.210 184.885 102.545 185.300 ;
        RECT 102.715 185.055 102.885 185.495 ;
        RECT 103.070 185.105 104.335 185.285 ;
        RECT 103.070 184.885 103.410 185.105 ;
        RECT 104.595 185.035 104.775 185.495 ;
        RECT 102.210 184.755 103.410 184.885 ;
        RECT 103.585 184.865 103.950 184.935 ;
        RECT 102.210 184.715 103.240 184.755 ;
        RECT 103.585 184.685 104.825 184.865 ;
        RECT 100.805 183.915 101.480 184.085 ;
        RECT 100.805 183.285 100.975 183.915 ;
        RECT 99.610 183.115 100.975 183.285 ;
        RECT 101.145 182.945 101.435 183.745 ;
        RECT 101.650 183.125 102.035 184.085 ;
        RECT 102.210 184.305 102.705 184.505 ;
        RECT 102.210 183.965 102.530 184.305 ;
        RECT 102.875 184.255 103.205 184.505 ;
        RECT 103.375 184.255 103.840 184.505 ;
        RECT 104.010 184.255 104.365 184.505 ;
        RECT 102.875 184.135 103.055 184.255 ;
        RECT 102.700 183.965 103.055 184.135 ;
        RECT 104.545 184.085 104.825 184.685 ;
        RECT 102.210 182.945 102.530 183.785 ;
        RECT 102.700 183.175 102.900 183.965 ;
        RECT 103.225 183.875 104.825 184.085 ;
        RECT 103.225 183.115 103.610 183.875 ;
        RECT 104.005 182.945 104.805 183.705 ;
        RECT 104.995 183.115 105.210 185.215 ;
        RECT 105.445 184.695 105.615 185.495 ;
        RECT 105.885 184.725 108.475 185.495 ;
        RECT 105.435 182.945 105.685 184.135 ;
        RECT 105.885 184.035 107.095 184.555 ;
        RECT 107.265 184.205 108.475 184.725 ;
        RECT 108.705 184.675 108.915 185.495 ;
        RECT 109.085 184.695 109.415 185.325 ;
        RECT 109.085 184.095 109.335 184.695 ;
        RECT 109.585 184.675 109.815 185.495 ;
        RECT 110.115 184.625 110.285 185.190 ;
        RECT 110.475 184.965 110.705 185.270 ;
        RECT 110.875 185.135 111.205 185.495 ;
        RECT 111.400 184.965 111.690 185.315 ;
        RECT 110.475 184.795 111.690 184.965 ;
        RECT 111.870 184.655 112.130 185.495 ;
        RECT 112.305 184.750 112.560 185.325 ;
        RECT 112.730 185.115 113.060 185.495 ;
        RECT 113.275 184.945 113.445 185.325 ;
        RECT 112.730 184.775 113.445 184.945 ;
        RECT 109.505 184.255 109.835 184.505 ;
        RECT 110.115 184.455 110.635 184.625 ;
        RECT 105.885 182.945 108.475 184.035 ;
        RECT 108.705 182.945 108.915 184.085 ;
        RECT 109.085 183.115 109.415 184.095 ;
        RECT 109.585 182.945 109.815 184.085 ;
        RECT 110.030 183.925 110.275 184.285 ;
        RECT 110.465 184.075 110.635 184.455 ;
        RECT 110.805 184.255 111.190 184.585 ;
        RECT 111.370 184.475 111.630 184.585 ;
        RECT 111.370 184.305 111.635 184.475 ;
        RECT 111.370 184.255 111.630 184.305 ;
        RECT 110.465 183.795 110.815 184.075 ;
        RECT 110.030 182.945 110.285 183.745 ;
        RECT 110.485 183.115 110.815 183.795 ;
        RECT 110.995 183.205 111.190 184.255 ;
        RECT 111.370 182.945 111.690 184.085 ;
        RECT 111.870 182.945 112.130 184.095 ;
        RECT 112.305 184.020 112.475 184.750 ;
        RECT 112.730 184.585 112.900 184.775 ;
        RECT 113.705 184.770 113.995 185.495 ;
        RECT 114.255 184.625 114.425 185.190 ;
        RECT 114.615 184.965 114.845 185.270 ;
        RECT 115.015 185.135 115.345 185.495 ;
        RECT 115.540 184.965 115.830 185.315 ;
        RECT 114.615 184.795 115.830 184.965 ;
        RECT 116.005 184.745 117.215 185.495 ;
        RECT 112.645 184.255 112.900 184.585 ;
        RECT 112.730 184.045 112.900 184.255 ;
        RECT 113.180 184.225 113.535 184.595 ;
        RECT 114.255 184.455 114.775 184.625 ;
        RECT 112.305 183.115 112.560 184.020 ;
        RECT 112.730 183.875 113.445 184.045 ;
        RECT 112.730 182.945 113.060 183.705 ;
        RECT 113.275 183.115 113.445 183.875 ;
        RECT 113.705 182.945 113.995 184.110 ;
        RECT 114.170 183.925 114.415 184.285 ;
        RECT 114.605 184.075 114.775 184.455 ;
        RECT 114.945 184.255 115.330 184.585 ;
        RECT 115.510 184.475 115.770 184.585 ;
        RECT 115.510 184.305 115.775 184.475 ;
        RECT 115.510 184.255 115.770 184.305 ;
        RECT 114.605 183.795 114.955 184.075 ;
        RECT 114.170 182.945 114.425 183.745 ;
        RECT 114.625 183.115 114.955 183.795 ;
        RECT 115.135 183.205 115.330 184.255 ;
        RECT 115.510 182.945 115.830 184.085 ;
        RECT 116.005 184.035 116.525 184.575 ;
        RECT 116.695 184.205 117.215 184.745 ;
        RECT 117.385 184.725 120.895 185.495 ;
        RECT 117.385 184.035 119.075 184.555 ;
        RECT 119.245 184.205 120.895 184.725 ;
        RECT 121.065 184.755 121.325 185.325 ;
        RECT 121.495 185.095 121.880 185.495 ;
        RECT 122.050 184.925 122.305 185.325 ;
        RECT 121.495 184.755 122.305 184.925 ;
        RECT 122.495 184.755 122.740 185.325 ;
        RECT 122.910 185.095 123.295 185.495 ;
        RECT 123.465 184.925 123.720 185.325 ;
        RECT 122.910 184.755 123.720 184.925 ;
        RECT 123.910 184.755 124.335 185.325 ;
        RECT 124.505 185.095 124.890 185.495 ;
        RECT 125.060 184.925 125.495 185.325 ;
        RECT 124.505 184.755 125.495 184.925 ;
        RECT 121.065 184.085 121.250 184.755 ;
        RECT 121.495 184.585 121.845 184.755 ;
        RECT 122.495 184.585 122.665 184.755 ;
        RECT 122.910 184.585 123.260 184.755 ;
        RECT 123.910 184.585 124.260 184.755 ;
        RECT 124.505 184.585 124.840 184.755 ;
        RECT 125.665 184.745 126.875 185.495 ;
        RECT 121.420 184.255 121.845 184.585 ;
        RECT 116.005 182.945 117.215 184.035 ;
        RECT 117.385 182.945 120.895 184.035 ;
        RECT 121.065 183.115 121.325 184.085 ;
        RECT 121.495 183.735 121.845 184.255 ;
        RECT 122.015 184.085 122.665 184.585 ;
        RECT 122.835 184.255 123.260 184.585 ;
        RECT 122.015 183.905 122.740 184.085 ;
        RECT 121.495 183.540 122.305 183.735 ;
        RECT 121.495 182.945 121.880 183.370 ;
        RECT 122.050 183.115 122.305 183.540 ;
        RECT 122.495 183.115 122.740 183.905 ;
        RECT 122.910 183.735 123.260 184.255 ;
        RECT 123.430 184.085 124.260 184.585 ;
        RECT 124.430 184.255 124.840 184.585 ;
        RECT 123.430 183.905 124.335 184.085 ;
        RECT 122.910 183.540 123.740 183.735 ;
        RECT 122.910 182.945 123.295 183.370 ;
        RECT 123.465 183.115 123.740 183.540 ;
        RECT 123.910 183.115 124.335 183.905 ;
        RECT 124.505 183.710 124.840 184.255 ;
        RECT 125.010 183.880 125.495 184.585 ;
        RECT 125.665 184.035 126.185 184.575 ;
        RECT 126.355 184.205 126.875 184.745 ;
        RECT 124.505 183.540 125.495 183.710 ;
        RECT 124.505 182.945 124.890 183.370 ;
        RECT 125.060 183.115 125.495 183.540 ;
        RECT 125.665 182.945 126.875 184.035 ;
        RECT 14.260 182.775 126.960 182.945 ;
        RECT 14.345 181.685 15.555 182.775 ;
        RECT 14.345 180.975 14.865 181.515 ;
        RECT 15.035 181.145 15.555 181.685 ;
        RECT 16.275 181.845 16.445 182.605 ;
        RECT 16.625 182.015 16.955 182.775 ;
        RECT 16.275 181.675 16.940 181.845 ;
        RECT 17.125 181.700 17.395 182.605 ;
        RECT 16.770 181.530 16.940 181.675 ;
        RECT 16.205 181.125 16.535 181.495 ;
        RECT 16.770 181.200 17.055 181.530 ;
        RECT 14.345 180.225 15.555 180.975 ;
        RECT 16.770 180.945 16.940 181.200 ;
        RECT 16.275 180.775 16.940 180.945 ;
        RECT 17.225 180.900 17.395 181.700 ;
        RECT 17.780 181.675 18.110 182.775 ;
        RECT 18.585 182.175 18.910 182.605 ;
        RECT 19.080 182.355 19.410 182.775 ;
        RECT 20.155 182.345 20.565 182.775 ;
        RECT 18.585 182.005 20.565 182.175 ;
        RECT 18.585 181.595 19.290 182.005 ;
        RECT 17.565 181.215 18.210 181.425 ;
        RECT 18.380 181.215 18.950 181.425 ;
        RECT 16.275 180.395 16.445 180.775 ;
        RECT 16.625 180.225 16.955 180.605 ;
        RECT 17.135 180.395 17.395 180.900 ;
        RECT 17.720 180.875 18.890 181.045 ;
        RECT 17.720 180.410 18.050 180.875 ;
        RECT 18.220 180.225 18.390 180.695 ;
        RECT 18.560 180.395 18.890 180.875 ;
        RECT 19.120 180.395 19.290 181.595 ;
        RECT 19.460 181.665 20.085 181.835 ;
        RECT 19.460 180.965 19.630 181.665 ;
        RECT 20.300 181.465 20.565 182.005 ;
        RECT 20.735 181.620 21.075 182.605 ;
        RECT 21.285 182.435 22.425 182.605 ;
        RECT 21.285 181.975 21.585 182.435 ;
        RECT 21.755 181.805 22.085 182.265 ;
        RECT 19.800 181.135 20.130 181.465 ;
        RECT 20.300 181.135 20.650 181.465 ;
        RECT 20.820 180.965 21.075 181.620 ;
        RECT 19.460 180.795 20.000 180.965 ;
        RECT 19.830 180.590 20.000 180.795 ;
        RECT 20.280 180.225 20.450 180.965 ;
        RECT 20.715 180.590 21.075 180.965 ;
        RECT 21.325 181.585 22.085 181.805 ;
        RECT 22.255 181.805 22.425 182.435 ;
        RECT 22.595 181.975 22.925 182.775 ;
        RECT 23.095 181.805 23.370 182.605 ;
        RECT 22.255 181.595 23.370 181.805 ;
        RECT 23.545 181.610 23.835 182.775 ;
        RECT 24.545 181.845 24.725 182.605 ;
        RECT 24.905 182.015 25.235 182.775 ;
        RECT 24.545 181.675 25.220 181.845 ;
        RECT 25.405 181.700 25.675 182.605 ;
        RECT 21.325 181.045 21.540 181.585 ;
        RECT 25.050 181.530 25.220 181.675 ;
        RECT 21.710 181.215 22.480 181.415 ;
        RECT 22.650 181.215 23.370 181.415 ;
        RECT 24.485 181.125 24.825 181.495 ;
        RECT 25.050 181.200 25.325 181.530 ;
        RECT 21.325 180.875 22.925 181.045 ;
        RECT 21.755 180.865 22.925 180.875 ;
        RECT 21.295 180.225 21.585 180.695 ;
        RECT 21.755 180.395 22.085 180.865 ;
        RECT 22.255 180.225 22.425 180.695 ;
        RECT 22.595 180.395 22.925 180.865 ;
        RECT 23.095 180.225 23.370 181.045 ;
        RECT 23.545 180.225 23.835 180.950 ;
        RECT 25.050 180.945 25.220 181.200 ;
        RECT 24.555 180.775 25.220 180.945 ;
        RECT 25.495 180.900 25.675 181.700 ;
        RECT 25.985 181.585 26.155 182.775 ;
        RECT 26.325 181.935 26.580 182.605 ;
        RECT 26.750 182.015 27.080 182.775 ;
        RECT 27.250 182.175 27.500 182.605 ;
        RECT 27.670 182.355 28.025 182.775 ;
        RECT 28.215 182.435 29.385 182.605 ;
        RECT 28.215 182.395 28.545 182.435 ;
        RECT 28.655 182.175 28.885 182.265 ;
        RECT 27.250 181.935 28.885 182.175 ;
        RECT 29.055 181.935 29.385 182.435 ;
        RECT 24.555 180.395 24.725 180.775 ;
        RECT 24.905 180.225 25.235 180.605 ;
        RECT 25.415 180.395 25.675 180.900 ;
        RECT 25.985 180.225 26.155 181.120 ;
        RECT 26.325 180.805 26.495 181.935 ;
        RECT 29.555 181.765 29.725 182.605 ;
        RECT 30.035 181.935 30.285 182.775 ;
        RECT 30.455 181.765 30.705 182.605 ;
        RECT 30.875 181.935 31.125 182.775 ;
        RECT 31.295 181.765 31.545 182.605 ;
        RECT 31.770 181.935 32.020 182.775 ;
        RECT 32.305 181.925 32.625 182.515 ;
        RECT 26.665 181.595 29.725 181.765 ;
        RECT 29.985 181.595 31.545 181.765 ;
        RECT 26.665 181.045 26.835 181.595 ;
        RECT 27.065 181.215 27.430 181.415 ;
        RECT 27.600 181.215 27.930 181.415 ;
        RECT 26.665 180.875 27.465 181.045 ;
        RECT 26.325 180.735 26.510 180.805 ;
        RECT 26.325 180.725 26.535 180.735 ;
        RECT 26.325 180.395 26.580 180.725 ;
        RECT 26.795 180.225 27.125 180.705 ;
        RECT 27.295 180.645 27.465 180.875 ;
        RECT 27.645 180.815 27.930 181.215 ;
        RECT 28.200 181.215 28.675 181.415 ;
        RECT 28.845 181.215 29.290 181.415 ;
        RECT 29.460 181.215 29.815 181.425 ;
        RECT 28.200 180.815 28.480 181.215 ;
        RECT 29.985 181.045 30.215 181.595 ;
        RECT 31.750 181.585 32.185 181.755 ;
        RECT 30.385 181.215 31.845 181.385 ;
        RECT 28.660 180.875 29.725 181.045 ;
        RECT 28.660 180.645 28.830 180.875 ;
        RECT 27.295 180.395 28.830 180.645 ;
        RECT 29.055 180.225 29.385 180.705 ;
        RECT 29.555 180.395 29.725 180.875 ;
        RECT 29.985 180.865 31.505 181.045 ;
        RECT 30.075 180.225 30.245 180.695 ;
        RECT 30.415 180.395 30.745 180.865 ;
        RECT 30.915 180.225 31.085 180.695 ;
        RECT 31.255 180.395 31.505 180.865 ;
        RECT 31.675 180.965 31.845 181.215 ;
        RECT 32.015 181.135 32.185 181.585 ;
        RECT 32.415 181.590 32.625 181.925 ;
        RECT 32.975 182.435 34.295 182.605 ;
        RECT 32.415 181.135 32.745 181.590 ;
        RECT 32.975 181.135 33.145 182.435 ;
        RECT 33.315 182.095 33.910 182.265 ;
        RECT 34.125 182.175 34.295 182.435 ;
        RECT 34.575 182.345 34.905 182.775 ;
        RECT 35.075 182.175 35.335 182.595 ;
        RECT 33.315 180.965 33.485 182.095 ;
        RECT 34.125 182.005 35.335 182.175 ;
        RECT 33.825 181.665 34.430 181.835 ;
        RECT 33.825 181.465 34.015 181.665 ;
        RECT 33.725 181.135 34.015 181.465 ;
        RECT 34.185 181.135 34.475 181.465 ;
        RECT 34.645 181.135 34.995 181.835 ;
        RECT 31.675 180.795 33.485 180.965 ;
        RECT 33.825 180.965 34.015 181.135 ;
        RECT 35.165 180.965 35.335 182.005 ;
        RECT 35.530 182.245 35.790 182.605 ;
        RECT 35.960 182.415 36.290 182.775 ;
        RECT 36.470 182.245 36.640 182.605 ;
        RECT 36.895 182.335 37.065 182.775 ;
        RECT 37.235 182.425 38.510 182.605 ;
        RECT 35.530 182.165 36.640 182.245 ;
        RECT 37.235 182.165 37.565 182.425 ;
        RECT 35.530 181.995 37.565 182.165 ;
        RECT 35.565 181.635 37.350 181.815 ;
        RECT 35.565 181.175 36.065 181.635 ;
        RECT 36.235 181.135 36.845 181.465 ;
        RECT 37.025 181.385 37.350 181.635 ;
        RECT 37.025 181.215 37.355 181.385 ;
        RECT 33.825 180.795 34.345 180.965 ;
        RECT 31.685 180.225 32.065 180.625 ;
        RECT 32.285 180.445 32.455 180.795 ;
        RECT 32.625 180.225 32.955 180.625 ;
        RECT 33.155 180.445 33.325 180.795 ;
        RECT 33.575 180.225 33.905 180.620 ;
        RECT 34.175 180.590 34.345 180.795 ;
        RECT 34.595 180.225 34.765 180.965 ;
        RECT 35.020 180.590 35.335 180.965 ;
        RECT 35.520 180.225 35.815 181.005 ;
        RECT 37.735 180.925 38.035 182.255 ;
        RECT 38.205 181.935 38.510 182.425 ;
        RECT 38.775 182.315 39.025 182.775 ;
        RECT 39.235 182.145 39.405 182.605 ;
        RECT 38.730 181.975 39.405 182.145 ;
        RECT 39.575 181.975 39.825 182.775 ;
        RECT 39.995 182.145 40.245 182.565 ;
        RECT 40.455 182.315 40.785 182.775 ;
        RECT 40.975 182.145 41.225 182.565 ;
        RECT 39.995 181.975 41.285 182.145 ;
        RECT 38.220 181.135 38.495 181.765 ;
        RECT 38.730 181.025 38.985 181.975 ;
        RECT 41.515 181.805 41.685 182.605 ;
        RECT 39.195 181.635 41.685 181.805 ;
        RECT 41.945 181.925 42.205 182.605 ;
        RECT 42.375 181.995 42.625 182.775 ;
        RECT 42.875 182.225 43.125 182.605 ;
        RECT 43.295 182.395 43.650 182.775 ;
        RECT 44.655 182.385 44.990 182.605 ;
        RECT 44.255 182.225 44.485 182.265 ;
        RECT 42.875 182.025 44.485 182.225 ;
        RECT 42.875 182.015 43.710 182.025 ;
        RECT 44.300 181.935 44.485 182.025 ;
        RECT 39.195 181.385 39.365 181.635 ;
        RECT 39.195 181.215 39.525 181.385 ;
        RECT 39.705 181.135 40.035 181.465 ;
        RECT 40.265 181.385 40.435 181.400 ;
        RECT 40.265 181.215 40.595 181.385 ;
        RECT 36.375 180.755 38.035 180.925 ;
        RECT 36.375 180.395 36.720 180.755 ;
        RECT 37.180 180.225 37.510 180.585 ;
        RECT 37.715 180.395 38.035 180.755 ;
        RECT 38.215 180.225 38.545 180.965 ;
        RECT 38.730 180.855 39.405 181.025 ;
        RECT 39.705 180.900 39.910 181.135 ;
        RECT 40.265 181.005 40.435 181.215 ;
        RECT 40.825 181.075 40.995 181.465 ;
        RECT 40.715 181.010 40.995 181.075 ;
        RECT 38.730 180.225 38.985 180.685 ;
        RECT 39.235 180.395 39.405 180.855 ;
        RECT 40.170 180.835 40.435 181.005 ;
        RECT 40.605 180.840 40.995 181.010 ;
        RECT 40.170 180.735 40.340 180.835 ;
        RECT 39.655 180.605 39.825 180.685 ;
        RECT 39.595 180.225 39.925 180.605 ;
        RECT 40.165 180.565 40.340 180.735 ;
        RECT 40.170 180.540 40.340 180.565 ;
        RECT 40.605 180.555 40.815 180.840 ;
        RECT 41.175 180.645 41.345 181.635 ;
        RECT 41.535 180.895 41.730 181.465 ;
        RECT 41.945 180.725 42.115 181.925 ;
        RECT 43.815 181.825 44.145 181.855 ;
        RECT 42.345 181.765 44.145 181.825 ;
        RECT 44.735 181.765 44.990 182.385 ;
        RECT 42.285 181.655 44.990 181.765 ;
        RECT 42.285 181.620 42.485 181.655 ;
        RECT 42.285 181.045 42.455 181.620 ;
        RECT 43.815 181.595 44.990 181.655 ;
        RECT 45.165 181.635 45.445 182.775 ;
        RECT 45.615 181.625 45.945 182.605 ;
        RECT 46.115 181.635 46.375 182.775 ;
        RECT 46.545 181.635 46.825 182.775 ;
        RECT 46.995 181.625 47.325 182.605 ;
        RECT 47.495 181.635 47.755 182.775 ;
        RECT 47.925 181.700 48.195 182.605 ;
        RECT 48.365 182.015 48.695 182.775 ;
        RECT 48.875 181.845 49.055 182.605 ;
        RECT 42.685 181.180 43.095 181.485 ;
        RECT 43.265 181.215 43.595 181.425 ;
        RECT 42.285 180.925 42.555 181.045 ;
        RECT 42.285 180.880 43.130 180.925 ;
        RECT 42.375 180.755 43.130 180.880 ;
        RECT 43.385 180.815 43.595 181.215 ;
        RECT 43.840 181.215 44.315 181.425 ;
        RECT 44.505 181.215 44.995 181.415 ;
        RECT 43.840 180.815 44.060 181.215 ;
        RECT 45.175 181.195 45.510 181.465 ;
        RECT 45.680 181.025 45.850 181.625 ;
        RECT 46.020 181.215 46.355 181.465 ;
        RECT 46.555 181.195 46.890 181.465 ;
        RECT 47.060 181.025 47.230 181.625 ;
        RECT 47.400 181.215 47.735 181.465 ;
        RECT 41.015 180.475 41.345 180.645 ;
        RECT 41.100 180.395 41.345 180.475 ;
        RECT 41.515 180.225 41.775 180.705 ;
        RECT 41.945 180.395 42.205 180.725 ;
        RECT 42.960 180.605 43.130 180.755 ;
        RECT 42.375 180.225 42.705 180.585 ;
        RECT 42.960 180.395 44.260 180.605 ;
        RECT 44.535 180.225 44.990 180.990 ;
        RECT 45.165 180.225 45.475 181.025 ;
        RECT 45.680 180.395 46.375 181.025 ;
        RECT 46.545 180.225 46.855 181.025 ;
        RECT 47.060 180.395 47.755 181.025 ;
        RECT 47.925 180.900 48.105 181.700 ;
        RECT 48.380 181.675 49.055 181.845 ;
        RECT 48.380 181.530 48.550 181.675 ;
        RECT 49.305 181.610 49.595 182.775 ;
        RECT 49.775 181.805 50.105 182.590 ;
        RECT 49.775 181.635 50.455 181.805 ;
        RECT 50.635 181.635 50.965 182.775 ;
        RECT 52.065 182.015 52.730 182.605 ;
        RECT 48.275 181.200 48.550 181.530 ;
        RECT 48.380 180.945 48.550 181.200 ;
        RECT 48.775 181.125 49.115 181.495 ;
        RECT 49.765 181.215 50.115 181.465 ;
        RECT 50.285 181.035 50.455 181.635 ;
        RECT 50.625 181.215 50.975 181.465 ;
        RECT 52.065 181.045 52.315 182.015 ;
        RECT 52.900 181.935 53.230 182.775 ;
        RECT 53.740 182.185 54.545 182.605 ;
        RECT 53.400 182.015 54.965 182.185 ;
        RECT 53.400 181.765 53.570 182.015 ;
        RECT 52.650 181.595 53.570 181.765 ;
        RECT 53.740 181.755 54.115 181.845 ;
        RECT 52.650 181.425 52.820 181.595 ;
        RECT 53.740 181.585 54.135 181.755 ;
        RECT 53.740 181.425 54.115 181.585 ;
        RECT 52.485 181.215 52.820 181.425 ;
        RECT 52.990 181.215 53.440 181.425 ;
        RECT 53.630 181.215 54.115 181.425 ;
        RECT 54.305 181.465 54.625 181.845 ;
        RECT 54.795 181.765 54.965 182.015 ;
        RECT 55.135 181.935 55.385 182.775 ;
        RECT 55.580 181.765 55.880 182.605 ;
        RECT 54.795 181.595 55.880 181.765 ;
        RECT 56.205 181.700 56.475 182.605 ;
        RECT 56.645 182.015 56.975 182.775 ;
        RECT 57.155 181.845 57.335 182.605 ;
        RECT 54.305 181.215 54.685 181.465 ;
        RECT 54.865 181.215 55.195 181.425 ;
        RECT 47.925 180.395 48.185 180.900 ;
        RECT 48.380 180.775 49.045 180.945 ;
        RECT 48.365 180.225 48.695 180.605 ;
        RECT 48.875 180.395 49.045 180.775 ;
        RECT 49.305 180.225 49.595 180.950 ;
        RECT 49.785 180.225 50.025 181.035 ;
        RECT 50.195 180.395 50.525 181.035 ;
        RECT 50.695 180.225 50.965 181.035 ;
        RECT 52.065 180.405 52.750 181.045 ;
        RECT 52.920 180.225 53.090 181.045 ;
        RECT 53.260 180.875 54.960 181.045 ;
        RECT 53.260 180.410 53.590 180.875 ;
        RECT 54.575 180.785 54.960 180.875 ;
        RECT 55.365 180.965 55.535 181.595 ;
        RECT 55.705 181.135 56.035 181.425 ;
        RECT 55.365 180.785 55.875 180.965 ;
        RECT 53.760 180.225 53.930 180.695 ;
        RECT 54.190 180.445 55.375 180.615 ;
        RECT 55.545 180.395 55.875 180.785 ;
        RECT 56.205 180.900 56.385 181.700 ;
        RECT 56.660 181.675 57.335 181.845 ;
        RECT 56.660 181.530 56.830 181.675 ;
        RECT 56.555 181.200 56.830 181.530 ;
        RECT 56.660 180.945 56.830 181.200 ;
        RECT 57.055 181.125 57.395 181.495 ;
        RECT 56.205 180.395 56.465 180.900 ;
        RECT 56.660 180.775 57.325 180.945 ;
        RECT 56.645 180.225 56.975 180.605 ;
        RECT 57.155 180.395 57.325 180.775 ;
        RECT 57.585 180.395 58.335 182.605 ;
        RECT 58.595 182.435 59.755 182.605 ;
        RECT 58.595 181.935 58.765 182.435 ;
        RECT 59.025 181.805 59.195 182.265 ;
        RECT 59.425 182.185 59.755 182.435 ;
        RECT 59.980 182.355 60.310 182.775 ;
        RECT 60.565 182.185 60.850 182.605 ;
        RECT 59.425 182.015 60.850 182.185 ;
        RECT 61.095 181.975 61.425 182.775 ;
        RECT 61.675 182.055 62.010 182.565 ;
        RECT 62.650 182.340 67.995 182.775 ;
        RECT 58.570 181.465 58.775 181.755 ;
        RECT 59.025 181.635 61.395 181.805 ;
        RECT 61.225 181.465 61.395 181.635 ;
        RECT 58.570 181.415 58.920 181.465 ;
        RECT 58.565 181.245 58.920 181.415 ;
        RECT 58.570 181.135 58.920 181.245 ;
        RECT 58.515 180.225 58.845 180.945 ;
        RECT 59.230 180.800 59.650 181.465 ;
        RECT 59.820 181.415 60.110 181.465 ;
        RECT 60.300 181.415 60.570 181.465 ;
        RECT 60.780 181.415 61.030 181.465 ;
        RECT 59.820 181.245 60.115 181.415 ;
        RECT 60.300 181.245 60.575 181.415 ;
        RECT 60.780 181.245 61.035 181.415 ;
        RECT 59.820 180.805 60.110 181.245 ;
        RECT 60.300 180.805 60.570 181.245 ;
        RECT 60.780 181.135 61.030 181.245 ;
        RECT 61.225 181.135 61.530 181.465 ;
        RECT 61.225 180.965 61.395 181.135 ;
        RECT 60.835 180.795 61.395 180.965 ;
        RECT 60.835 180.625 61.005 180.795 ;
        RECT 61.755 180.700 62.010 182.055 ;
        RECT 64.240 181.090 64.590 182.340 ;
        RECT 68.165 181.635 68.425 182.775 ;
        RECT 68.595 181.625 68.925 182.605 ;
        RECT 69.095 181.635 69.375 182.775 ;
        RECT 69.545 181.685 71.215 182.775 ;
        RECT 71.390 181.975 71.645 182.775 ;
        RECT 71.845 181.925 72.175 182.605 ;
        RECT 66.070 180.770 66.410 181.600 ;
        RECT 68.185 181.215 68.520 181.465 ;
        RECT 68.690 181.025 68.860 181.625 ;
        RECT 69.030 181.195 69.365 181.465 ;
        RECT 69.545 181.165 70.295 181.685 ;
        RECT 59.390 180.455 61.005 180.625 ;
        RECT 61.175 180.225 61.505 180.625 ;
        RECT 61.675 180.440 62.010 180.700 ;
        RECT 62.650 180.225 67.995 180.770 ;
        RECT 68.165 180.395 68.860 181.025 ;
        RECT 69.065 180.225 69.375 181.025 ;
        RECT 70.465 180.995 71.215 181.515 ;
        RECT 71.390 181.435 71.635 181.795 ;
        RECT 71.825 181.645 72.175 181.925 ;
        RECT 71.825 181.265 71.995 181.645 ;
        RECT 72.355 181.465 72.550 182.515 ;
        RECT 72.730 181.635 73.050 182.775 ;
        RECT 73.685 181.635 73.945 182.775 ;
        RECT 74.115 181.625 74.445 182.605 ;
        RECT 74.615 181.635 74.895 182.775 ;
        RECT 69.545 180.225 71.215 180.995 ;
        RECT 71.475 181.095 71.995 181.265 ;
        RECT 72.165 181.135 72.550 181.465 ;
        RECT 72.730 181.415 72.990 181.465 ;
        RECT 72.730 181.245 72.995 181.415 ;
        RECT 72.730 181.135 72.990 181.245 ;
        RECT 73.705 181.215 74.040 181.465 ;
        RECT 71.475 180.735 71.645 181.095 ;
        RECT 74.210 181.025 74.380 181.625 ;
        RECT 75.065 181.610 75.355 182.775 ;
        RECT 75.525 181.685 76.735 182.775 ;
        RECT 76.910 182.340 82.255 182.775 ;
        RECT 74.550 181.195 74.885 181.465 ;
        RECT 75.525 181.145 76.045 181.685 ;
        RECT 71.445 180.565 71.645 180.735 ;
        RECT 71.475 180.530 71.645 180.565 ;
        RECT 71.835 180.755 73.050 180.925 ;
        RECT 71.835 180.450 72.065 180.755 ;
        RECT 72.235 180.225 72.565 180.585 ;
        RECT 72.760 180.405 73.050 180.755 ;
        RECT 73.685 180.395 74.380 181.025 ;
        RECT 74.585 180.225 74.895 181.025 ;
        RECT 76.215 180.975 76.735 181.515 ;
        RECT 78.500 181.090 78.850 182.340 ;
        RECT 82.425 182.185 83.125 182.605 ;
        RECT 83.325 182.415 83.655 182.775 ;
        RECT 83.825 182.185 84.155 182.585 ;
        RECT 82.425 181.955 84.155 182.185 ;
        RECT 75.065 180.225 75.355 180.950 ;
        RECT 75.525 180.225 76.735 180.975 ;
        RECT 80.330 180.770 80.670 181.600 ;
        RECT 82.425 180.985 82.630 181.955 ;
        RECT 82.800 181.215 83.130 181.755 ;
        RECT 83.305 181.465 83.630 181.755 ;
        RECT 83.825 181.735 84.155 181.955 ;
        RECT 84.325 181.465 84.495 182.435 ;
        RECT 84.675 181.715 85.005 182.775 ;
        RECT 85.185 182.345 85.525 182.605 ;
        RECT 83.305 181.135 83.800 181.465 ;
        RECT 84.120 181.135 84.495 181.465 ;
        RECT 84.705 181.135 85.015 181.465 ;
        RECT 76.910 180.225 82.255 180.770 ;
        RECT 82.425 180.395 83.135 180.985 ;
        RECT 83.645 180.755 85.005 180.965 ;
        RECT 83.645 180.395 83.975 180.755 ;
        RECT 84.175 180.225 84.505 180.585 ;
        RECT 84.675 180.395 85.005 180.755 ;
        RECT 85.185 180.945 85.445 182.345 ;
        RECT 85.695 181.975 86.025 182.775 ;
        RECT 86.490 181.805 86.740 182.605 ;
        RECT 86.925 182.055 87.255 182.775 ;
        RECT 87.475 181.805 87.725 182.605 ;
        RECT 87.895 182.395 88.230 182.775 ;
        RECT 85.635 181.635 87.825 181.805 ;
        RECT 85.635 181.465 85.950 181.635 ;
        RECT 85.620 181.215 85.950 181.465 ;
        RECT 85.185 180.435 85.525 180.945 ;
        RECT 85.695 180.225 85.965 181.025 ;
        RECT 86.145 180.495 86.425 181.465 ;
        RECT 86.605 180.495 86.905 181.465 ;
        RECT 87.085 180.500 87.435 181.465 ;
        RECT 87.655 180.725 87.825 181.635 ;
        RECT 87.995 180.905 88.235 182.215 ;
        RECT 88.405 181.685 89.615 182.775 ;
        RECT 89.785 181.685 93.295 182.775 ;
        RECT 93.470 182.340 98.815 182.775 ;
        RECT 88.405 181.145 88.925 181.685 ;
        RECT 89.095 180.975 89.615 181.515 ;
        RECT 89.785 181.165 91.475 181.685 ;
        RECT 91.645 180.995 93.295 181.515 ;
        RECT 95.060 181.090 95.410 182.340 ;
        RECT 98.985 181.635 99.265 182.775 ;
        RECT 99.435 181.625 99.765 182.605 ;
        RECT 99.935 181.635 100.195 182.775 ;
        RECT 87.655 180.395 88.150 180.725 ;
        RECT 88.405 180.225 89.615 180.975 ;
        RECT 89.785 180.225 93.295 180.995 ;
        RECT 96.890 180.770 97.230 181.600 ;
        RECT 98.995 181.195 99.330 181.465 ;
        RECT 99.500 181.025 99.670 181.625 ;
        RECT 100.825 181.610 101.115 182.775 ;
        RECT 101.805 181.635 102.015 182.775 ;
        RECT 102.185 181.625 102.515 182.605 ;
        RECT 102.685 181.635 102.915 182.775 ;
        RECT 104.045 181.685 107.555 182.775 ;
        RECT 99.840 181.215 100.175 181.465 ;
        RECT 93.470 180.225 98.815 180.770 ;
        RECT 98.985 180.225 99.295 181.025 ;
        RECT 99.500 180.395 100.195 181.025 ;
        RECT 100.825 180.225 101.115 180.950 ;
        RECT 101.805 180.225 102.015 181.045 ;
        RECT 102.185 181.025 102.435 181.625 ;
        RECT 102.605 181.215 102.935 181.465 ;
        RECT 104.045 181.165 105.735 181.685 ;
        RECT 107.765 181.635 107.995 182.775 ;
        RECT 108.165 181.625 108.495 182.605 ;
        RECT 108.665 181.635 108.875 182.775 ;
        RECT 109.600 181.975 109.850 182.775 ;
        RECT 110.020 182.145 110.350 182.605 ;
        RECT 110.520 182.315 110.735 182.775 ;
        RECT 110.020 181.975 111.190 182.145 ;
        RECT 109.110 181.805 109.390 181.965 ;
        RECT 109.110 181.635 110.445 181.805 ;
        RECT 102.185 180.395 102.515 181.025 ;
        RECT 102.685 180.225 102.915 181.045 ;
        RECT 105.905 180.995 107.555 181.515 ;
        RECT 107.745 181.215 108.075 181.465 ;
        RECT 104.045 180.225 107.555 180.995 ;
        RECT 107.765 180.225 107.995 181.045 ;
        RECT 108.245 181.025 108.495 181.625 ;
        RECT 110.275 181.465 110.445 181.635 ;
        RECT 109.110 181.215 109.460 181.455 ;
        RECT 109.630 181.215 110.105 181.455 ;
        RECT 110.275 181.215 110.650 181.465 ;
        RECT 110.275 181.045 110.445 181.215 ;
        RECT 108.165 180.395 108.495 181.025 ;
        RECT 108.665 180.225 108.875 181.045 ;
        RECT 109.110 180.875 110.445 181.045 ;
        RECT 109.110 180.665 109.380 180.875 ;
        RECT 110.820 180.685 111.190 181.975 ;
        RECT 111.405 182.015 111.920 182.425 ;
        RECT 112.155 182.015 112.325 182.775 ;
        RECT 112.495 182.435 114.525 182.605 ;
        RECT 111.405 181.205 111.745 182.015 ;
        RECT 112.495 181.770 112.665 182.435 ;
        RECT 113.060 182.095 114.185 182.265 ;
        RECT 111.915 181.580 112.665 181.770 ;
        RECT 112.835 181.755 113.845 181.925 ;
        RECT 111.405 181.035 112.635 181.205 ;
        RECT 109.600 180.225 109.930 180.685 ;
        RECT 110.440 180.395 111.190 180.685 ;
        RECT 111.680 180.430 111.925 181.035 ;
        RECT 112.145 180.225 112.655 180.760 ;
        RECT 112.835 180.395 113.025 181.755 ;
        RECT 113.195 180.735 113.470 181.555 ;
        RECT 113.675 180.955 113.845 181.755 ;
        RECT 114.015 180.965 114.185 182.095 ;
        RECT 114.355 181.465 114.525 182.435 ;
        RECT 114.695 181.635 114.865 182.775 ;
        RECT 115.035 181.635 115.370 182.605 ;
        RECT 114.355 181.135 114.550 181.465 ;
        RECT 114.775 181.135 115.030 181.465 ;
        RECT 114.775 180.965 114.945 181.135 ;
        RECT 115.200 180.965 115.370 181.635 ;
        RECT 116.465 181.685 119.975 182.775 ;
        RECT 120.150 182.340 125.495 182.775 ;
        RECT 116.465 181.165 118.155 181.685 ;
        RECT 118.325 180.995 119.975 181.515 ;
        RECT 121.740 181.090 122.090 182.340 ;
        RECT 125.665 181.685 126.875 182.775 ;
        RECT 114.015 180.795 114.945 180.965 ;
        RECT 114.015 180.760 114.190 180.795 ;
        RECT 113.195 180.565 113.475 180.735 ;
        RECT 113.195 180.395 113.470 180.565 ;
        RECT 113.660 180.395 114.190 180.760 ;
        RECT 114.615 180.225 114.945 180.625 ;
        RECT 115.115 180.395 115.370 180.965 ;
        RECT 116.465 180.225 119.975 180.995 ;
        RECT 123.570 180.770 123.910 181.600 ;
        RECT 125.665 181.145 126.185 181.685 ;
        RECT 126.355 180.975 126.875 181.515 ;
        RECT 120.150 180.225 125.495 180.770 ;
        RECT 125.665 180.225 126.875 180.975 ;
        RECT 14.260 180.055 126.960 180.225 ;
        RECT 14.345 179.305 15.555 180.055 ;
        RECT 16.185 179.380 16.445 179.885 ;
        RECT 16.625 179.675 16.955 180.055 ;
        RECT 17.135 179.505 17.305 179.885 ;
        RECT 17.625 179.690 17.795 179.715 ;
        RECT 14.345 178.765 14.865 179.305 ;
        RECT 15.035 178.595 15.555 179.135 ;
        RECT 14.345 177.505 15.555 178.595 ;
        RECT 16.185 178.580 16.365 179.380 ;
        RECT 16.640 179.335 17.305 179.505 ;
        RECT 16.640 179.080 16.810 179.335 ;
        RECT 17.565 179.315 17.925 179.690 ;
        RECT 18.190 179.315 18.360 180.055 ;
        RECT 18.640 179.485 18.810 179.690 ;
        RECT 18.640 179.315 19.180 179.485 ;
        RECT 16.535 178.750 16.810 179.080 ;
        RECT 17.035 178.785 17.375 179.155 ;
        RECT 16.640 178.605 16.810 178.750 ;
        RECT 17.565 178.660 17.820 179.315 ;
        RECT 17.990 178.815 18.340 179.145 ;
        RECT 18.510 178.815 18.840 179.145 ;
        RECT 16.185 177.675 16.455 178.580 ;
        RECT 16.640 178.435 17.315 178.605 ;
        RECT 16.625 177.505 16.955 178.265 ;
        RECT 17.135 177.675 17.315 178.435 ;
        RECT 17.565 177.675 17.905 178.660 ;
        RECT 18.075 178.275 18.340 178.815 ;
        RECT 19.010 178.615 19.180 179.315 ;
        RECT 18.555 178.445 19.180 178.615 ;
        RECT 19.350 178.685 19.520 179.885 ;
        RECT 19.750 179.405 20.080 179.885 ;
        RECT 20.250 179.585 20.420 180.055 ;
        RECT 20.590 179.405 20.920 179.870 ;
        RECT 22.165 179.545 22.470 180.055 ;
        RECT 19.750 179.235 20.920 179.405 ;
        RECT 19.690 178.855 20.260 179.065 ;
        RECT 20.430 178.855 21.075 179.065 ;
        RECT 22.165 178.815 22.480 179.375 ;
        RECT 22.650 179.065 22.900 179.875 ;
        RECT 23.070 179.530 23.330 180.055 ;
        RECT 23.510 179.065 23.760 179.875 ;
        RECT 23.930 179.495 24.190 180.055 ;
        RECT 24.360 179.405 24.620 179.860 ;
        RECT 24.790 179.575 25.050 180.055 ;
        RECT 25.220 179.405 25.480 179.860 ;
        RECT 25.650 179.575 25.910 180.055 ;
        RECT 26.080 179.405 26.340 179.860 ;
        RECT 26.510 179.575 26.755 180.055 ;
        RECT 26.925 179.405 27.200 179.860 ;
        RECT 27.370 179.575 27.615 180.055 ;
        RECT 27.785 179.405 28.045 179.860 ;
        RECT 28.225 179.575 28.475 180.055 ;
        RECT 28.645 179.405 28.905 179.860 ;
        RECT 29.085 179.575 29.335 180.055 ;
        RECT 29.505 179.405 29.765 179.860 ;
        RECT 29.945 179.575 30.205 180.055 ;
        RECT 30.375 179.405 30.635 179.860 ;
        RECT 30.805 179.575 31.105 180.055 ;
        RECT 31.455 179.505 31.625 179.885 ;
        RECT 31.805 179.675 32.135 180.055 ;
        RECT 24.360 179.235 31.105 179.405 ;
        RECT 31.455 179.335 32.120 179.505 ;
        RECT 32.315 179.380 32.575 179.885 ;
        RECT 32.790 179.695 33.120 180.055 ;
        RECT 33.290 179.525 33.620 179.885 ;
        RECT 33.790 179.615 34.025 180.055 ;
        RECT 34.615 179.675 34.950 180.055 ;
        RECT 35.910 179.715 36.245 179.885 ;
        RECT 22.650 178.815 29.770 179.065 ;
        RECT 19.350 178.275 20.055 178.685 ;
        RECT 18.075 178.105 20.055 178.275 ;
        RECT 18.075 177.505 18.485 177.935 ;
        RECT 19.230 177.505 19.560 177.925 ;
        RECT 19.730 177.675 20.055 178.105 ;
        RECT 20.530 177.505 20.860 178.605 ;
        RECT 22.175 177.505 22.470 178.315 ;
        RECT 22.650 177.675 22.895 178.815 ;
        RECT 23.070 177.505 23.330 178.315 ;
        RECT 23.510 177.680 23.760 178.815 ;
        RECT 29.940 178.645 31.105 179.235 ;
        RECT 31.385 178.785 31.715 179.155 ;
        RECT 31.950 179.080 32.120 179.335 ;
        RECT 24.360 178.420 31.105 178.645 ;
        RECT 31.950 178.750 32.235 179.080 ;
        RECT 31.950 178.605 32.120 178.750 ;
        RECT 31.455 178.435 32.120 178.605 ;
        RECT 32.405 178.580 32.575 179.380 ;
        RECT 24.360 178.405 29.765 178.420 ;
        RECT 23.930 177.510 24.190 178.305 ;
        RECT 24.360 177.680 24.620 178.405 ;
        RECT 24.790 177.510 25.050 178.235 ;
        RECT 25.220 177.680 25.480 178.405 ;
        RECT 25.650 177.510 25.910 178.235 ;
        RECT 26.080 177.680 26.340 178.405 ;
        RECT 26.510 177.510 26.770 178.235 ;
        RECT 26.940 177.680 27.200 178.405 ;
        RECT 27.370 177.510 27.615 178.235 ;
        RECT 27.785 177.680 28.045 178.405 ;
        RECT 28.230 177.510 28.475 178.235 ;
        RECT 28.645 177.680 28.905 178.405 ;
        RECT 29.090 177.510 29.335 178.235 ;
        RECT 29.505 177.680 29.765 178.405 ;
        RECT 29.950 177.510 30.205 178.235 ;
        RECT 30.375 177.680 30.665 178.420 ;
        RECT 23.930 177.505 30.205 177.510 ;
        RECT 30.835 177.505 31.105 178.250 ;
        RECT 31.455 177.675 31.625 178.435 ;
        RECT 31.805 177.505 32.135 178.265 ;
        RECT 32.305 177.675 32.575 178.580 ;
        RECT 32.800 179.355 33.620 179.525 ;
        RECT 32.800 178.235 32.995 179.355 ;
        RECT 34.190 179.315 35.460 179.505 ;
        RECT 35.630 179.315 36.245 179.715 ;
        RECT 36.425 179.330 36.715 180.055 ;
        RECT 36.895 179.445 37.225 179.865 ;
        RECT 37.395 179.615 37.670 180.055 ;
        RECT 37.875 179.445 38.205 179.865 ;
        RECT 38.685 179.695 39.535 180.055 ;
        RECT 39.705 179.505 39.925 179.885 ;
        RECT 33.165 178.815 33.845 179.145 ;
        RECT 34.015 178.815 34.350 179.145 ;
        RECT 34.520 179.035 34.810 179.145 ;
        RECT 34.520 178.865 34.815 179.035 ;
        RECT 34.520 178.815 34.810 178.865 ;
        RECT 35.100 178.815 35.460 179.145 ;
        RECT 33.675 178.630 33.845 178.815 ;
        RECT 35.630 178.630 35.810 179.315 ;
        RECT 36.895 179.265 39.480 179.445 ;
        RECT 35.980 178.815 36.255 179.145 ;
        RECT 36.885 178.865 37.220 179.095 ;
        RECT 37.410 179.035 37.860 179.095 ;
        RECT 37.405 178.865 37.860 179.035 ;
        RECT 38.030 178.865 38.500 179.095 ;
        RECT 38.670 178.865 39.000 179.095 ;
        RECT 33.675 178.375 36.250 178.630 ;
        RECT 32.800 178.065 33.530 178.235 ;
        RECT 32.840 177.505 33.170 177.885 ;
        RECT 33.340 177.675 33.530 178.065 ;
        RECT 33.710 177.505 34.140 178.205 ;
        RECT 34.645 177.675 35.315 178.375 ;
        RECT 35.485 177.505 35.815 178.205 ;
        RECT 35.985 177.675 36.250 178.375 ;
        RECT 36.425 177.505 36.715 178.670 ;
        RECT 39.170 178.650 39.480 179.265 ;
        RECT 36.895 178.480 39.480 178.650 ;
        RECT 36.895 177.815 37.225 178.480 ;
        RECT 37.685 178.120 39.025 178.300 ;
        RECT 37.685 177.675 38.015 178.120 ;
        RECT 38.250 177.505 38.525 177.950 ;
        RECT 38.695 177.675 39.025 178.120 ;
        RECT 39.225 177.505 39.480 178.310 ;
        RECT 39.695 177.805 39.925 179.505 ;
        RECT 40.095 179.235 40.390 180.055 ;
        RECT 40.600 179.315 41.215 179.885 ;
        RECT 41.385 179.545 41.600 180.055 ;
        RECT 41.830 179.545 42.110 179.875 ;
        RECT 42.290 179.545 42.530 180.055 ;
        RECT 40.095 177.505 40.390 178.650 ;
        RECT 40.600 178.295 40.915 179.315 ;
        RECT 41.085 178.645 41.255 179.145 ;
        RECT 41.505 178.815 41.770 179.375 ;
        RECT 41.940 178.645 42.110 179.545 ;
        RECT 42.955 179.505 43.125 179.885 ;
        RECT 43.305 179.675 43.635 180.055 ;
        RECT 42.280 178.815 42.635 179.375 ;
        RECT 42.955 179.335 43.620 179.505 ;
        RECT 43.815 179.380 44.075 179.885 ;
        RECT 42.885 178.785 43.225 179.155 ;
        RECT 43.450 179.080 43.620 179.335 ;
        RECT 43.450 178.750 43.725 179.080 ;
        RECT 41.085 178.475 42.510 178.645 ;
        RECT 43.450 178.605 43.620 178.750 ;
        RECT 40.600 177.675 41.135 178.295 ;
        RECT 41.305 177.505 41.635 178.305 ;
        RECT 42.120 178.300 42.510 178.475 ;
        RECT 42.945 178.435 43.620 178.605 ;
        RECT 43.895 178.580 44.075 179.380 ;
        RECT 44.335 179.505 44.505 179.885 ;
        RECT 44.685 179.675 45.015 180.055 ;
        RECT 44.335 179.335 45.000 179.505 ;
        RECT 45.195 179.380 45.455 179.885 ;
        RECT 44.265 178.785 44.605 179.155 ;
        RECT 44.830 179.080 45.000 179.335 ;
        RECT 44.830 178.750 45.105 179.080 ;
        RECT 44.830 178.605 45.000 178.750 ;
        RECT 42.945 177.675 43.125 178.435 ;
        RECT 43.305 177.505 43.635 178.265 ;
        RECT 43.805 177.675 44.075 178.580 ;
        RECT 44.325 178.435 45.000 178.605 ;
        RECT 45.275 178.580 45.455 179.380 ;
        RECT 44.325 177.675 44.505 178.435 ;
        RECT 44.685 177.505 45.015 178.265 ;
        RECT 45.185 177.675 45.455 178.580 ;
        RECT 45.625 179.380 45.885 179.885 ;
        RECT 46.065 179.675 46.395 180.055 ;
        RECT 46.575 179.505 46.745 179.885 ;
        RECT 45.625 178.580 45.795 179.380 ;
        RECT 46.080 179.335 46.745 179.505 ;
        RECT 46.080 179.080 46.250 179.335 ;
        RECT 47.045 179.235 47.275 180.055 ;
        RECT 47.445 179.255 47.775 179.885 ;
        RECT 45.965 178.750 46.250 179.080 ;
        RECT 46.485 178.785 46.815 179.155 ;
        RECT 47.025 178.815 47.355 179.065 ;
        RECT 46.080 178.605 46.250 178.750 ;
        RECT 47.525 178.655 47.775 179.255 ;
        RECT 47.945 179.235 48.155 180.055 ;
        RECT 48.425 179.235 48.655 180.055 ;
        RECT 48.825 179.255 49.155 179.885 ;
        RECT 48.405 178.815 48.735 179.065 ;
        RECT 48.905 178.655 49.155 179.255 ;
        RECT 49.325 179.235 49.535 180.055 ;
        RECT 49.785 179.245 50.025 180.055 ;
        RECT 50.195 179.245 50.525 179.885 ;
        RECT 50.695 179.245 50.965 180.055 ;
        RECT 51.145 179.380 51.405 179.885 ;
        RECT 51.585 179.675 51.915 180.055 ;
        RECT 52.095 179.505 52.265 179.885 ;
        RECT 49.765 178.815 50.115 179.065 ;
        RECT 45.625 177.675 45.895 178.580 ;
        RECT 46.080 178.435 46.745 178.605 ;
        RECT 46.065 177.505 46.395 178.265 ;
        RECT 46.575 177.675 46.745 178.435 ;
        RECT 47.045 177.505 47.275 178.645 ;
        RECT 47.445 177.675 47.775 178.655 ;
        RECT 47.945 177.505 48.155 178.645 ;
        RECT 48.425 177.505 48.655 178.645 ;
        RECT 48.825 177.675 49.155 178.655 ;
        RECT 50.285 178.645 50.455 179.245 ;
        RECT 50.625 178.815 50.975 179.065 ;
        RECT 49.325 177.505 49.535 178.645 ;
        RECT 49.775 178.475 50.455 178.645 ;
        RECT 49.775 177.690 50.105 178.475 ;
        RECT 50.635 177.505 50.965 178.645 ;
        RECT 51.145 178.580 51.325 179.380 ;
        RECT 51.600 179.335 52.265 179.505 ;
        RECT 52.525 179.555 52.785 179.885 ;
        RECT 52.955 179.695 53.285 180.055 ;
        RECT 53.540 179.675 54.840 179.885 ;
        RECT 51.600 179.080 51.770 179.335 ;
        RECT 51.495 178.750 51.770 179.080 ;
        RECT 51.995 178.785 52.335 179.155 ;
        RECT 51.600 178.605 51.770 178.750 ;
        RECT 51.145 177.675 51.415 178.580 ;
        RECT 51.600 178.435 52.275 178.605 ;
        RECT 51.585 177.505 51.915 178.265 ;
        RECT 52.095 177.675 52.275 178.435 ;
        RECT 52.525 178.355 52.695 179.555 ;
        RECT 53.540 179.525 53.710 179.675 ;
        RECT 52.955 179.400 53.710 179.525 ;
        RECT 52.865 179.355 53.710 179.400 ;
        RECT 52.865 179.235 53.135 179.355 ;
        RECT 52.865 178.660 53.035 179.235 ;
        RECT 53.265 178.795 53.675 179.100 ;
        RECT 53.965 179.065 54.175 179.465 ;
        RECT 53.845 178.855 54.175 179.065 ;
        RECT 54.420 179.065 54.640 179.465 ;
        RECT 55.115 179.290 55.570 180.055 ;
        RECT 56.665 179.425 57.005 179.885 ;
        RECT 57.175 179.595 57.345 180.055 ;
        RECT 57.975 179.620 58.335 179.885 ;
        RECT 57.980 179.615 58.335 179.620 ;
        RECT 57.985 179.605 58.335 179.615 ;
        RECT 57.990 179.600 58.335 179.605 ;
        RECT 57.995 179.590 58.335 179.600 ;
        RECT 58.575 179.595 58.745 180.055 ;
        RECT 58.000 179.585 58.335 179.590 ;
        RECT 58.010 179.575 58.335 179.585 ;
        RECT 58.020 179.565 58.335 179.575 ;
        RECT 57.515 179.425 57.845 179.505 ;
        RECT 56.665 179.235 57.845 179.425 ;
        RECT 58.035 179.425 58.335 179.565 ;
        RECT 58.035 179.235 58.745 179.425 ;
        RECT 54.420 178.855 54.895 179.065 ;
        RECT 55.085 178.865 55.575 179.065 ;
        RECT 56.665 178.865 56.995 179.065 ;
        RECT 57.305 179.045 57.635 179.065 ;
        RECT 57.185 178.865 57.635 179.045 ;
        RECT 52.865 178.625 53.065 178.660 ;
        RECT 54.395 178.625 55.570 178.685 ;
        RECT 52.865 178.515 55.570 178.625 ;
        RECT 56.665 178.525 56.895 178.865 ;
        RECT 52.925 178.455 54.725 178.515 ;
        RECT 54.395 178.425 54.725 178.455 ;
        RECT 52.525 177.675 52.785 178.355 ;
        RECT 52.955 177.505 53.205 178.285 ;
        RECT 53.455 178.255 54.290 178.265 ;
        RECT 54.880 178.255 55.065 178.345 ;
        RECT 53.455 178.055 55.065 178.255 ;
        RECT 53.455 177.675 53.705 178.055 ;
        RECT 54.835 178.015 55.065 178.055 ;
        RECT 55.315 177.895 55.570 178.515 ;
        RECT 53.875 177.505 54.230 177.885 ;
        RECT 55.235 177.675 55.570 177.895 ;
        RECT 56.675 177.505 57.005 178.225 ;
        RECT 57.185 177.750 57.400 178.865 ;
        RECT 57.805 178.835 58.275 179.065 ;
        RECT 58.460 178.665 58.745 179.235 ;
        RECT 58.915 179.110 59.255 179.885 ;
        RECT 59.425 179.285 62.015 180.055 ;
        RECT 62.185 179.330 62.475 180.055 ;
        RECT 57.595 178.450 58.745 178.665 ;
        RECT 57.595 177.675 57.925 178.450 ;
        RECT 58.095 177.505 58.805 178.280 ;
        RECT 58.975 177.675 59.255 179.110 ;
        RECT 59.425 178.595 60.635 179.115 ;
        RECT 60.805 178.765 62.015 179.285 ;
        RECT 62.920 179.245 63.165 179.850 ;
        RECT 63.385 179.520 63.895 180.055 ;
        RECT 62.645 179.075 63.875 179.245 ;
        RECT 59.425 177.505 62.015 178.595 ;
        RECT 62.185 177.505 62.475 178.670 ;
        RECT 62.645 178.265 62.985 179.075 ;
        RECT 63.155 178.510 63.905 178.700 ;
        RECT 62.645 177.855 63.160 178.265 ;
        RECT 63.395 177.505 63.565 178.265 ;
        RECT 63.735 177.845 63.905 178.510 ;
        RECT 64.075 178.525 64.265 179.885 ;
        RECT 64.435 179.035 64.710 179.885 ;
        RECT 64.900 179.520 65.430 179.885 ;
        RECT 65.855 179.655 66.185 180.055 ;
        RECT 65.255 179.485 65.430 179.520 ;
        RECT 64.435 178.865 64.715 179.035 ;
        RECT 64.435 178.725 64.710 178.865 ;
        RECT 64.915 178.525 65.085 179.325 ;
        RECT 64.075 178.355 65.085 178.525 ;
        RECT 65.255 179.315 66.185 179.485 ;
        RECT 66.355 179.315 66.610 179.885 ;
        RECT 65.255 178.185 65.425 179.315 ;
        RECT 66.015 179.145 66.185 179.315 ;
        RECT 64.300 178.015 65.425 178.185 ;
        RECT 65.595 178.815 65.790 179.145 ;
        RECT 66.015 178.815 66.270 179.145 ;
        RECT 65.595 177.845 65.765 178.815 ;
        RECT 66.440 178.645 66.610 179.315 ;
        RECT 63.735 177.675 65.765 177.845 ;
        RECT 65.935 177.505 66.105 178.645 ;
        RECT 66.275 177.675 66.610 178.645 ;
        RECT 66.790 179.315 67.045 179.885 ;
        RECT 67.215 179.655 67.545 180.055 ;
        RECT 67.970 179.520 68.500 179.885 ;
        RECT 68.690 179.715 68.965 179.885 ;
        RECT 68.685 179.545 68.965 179.715 ;
        RECT 67.970 179.485 68.145 179.520 ;
        RECT 67.215 179.315 68.145 179.485 ;
        RECT 66.790 178.645 66.960 179.315 ;
        RECT 67.215 179.145 67.385 179.315 ;
        RECT 67.130 178.815 67.385 179.145 ;
        RECT 67.610 178.815 67.805 179.145 ;
        RECT 66.790 177.675 67.125 178.645 ;
        RECT 67.295 177.505 67.465 178.645 ;
        RECT 67.635 177.845 67.805 178.815 ;
        RECT 67.975 178.185 68.145 179.315 ;
        RECT 68.315 178.525 68.485 179.325 ;
        RECT 68.690 178.725 68.965 179.545 ;
        RECT 69.135 178.525 69.325 179.885 ;
        RECT 69.505 179.520 70.015 180.055 ;
        RECT 70.235 179.245 70.480 179.850 ;
        RECT 71.845 179.255 72.540 179.885 ;
        RECT 72.745 179.255 73.055 180.055 ;
        RECT 73.225 179.415 73.565 179.820 ;
        RECT 73.735 179.585 73.905 180.055 ;
        RECT 74.075 179.415 74.325 179.820 ;
        RECT 69.525 179.075 70.755 179.245 ;
        RECT 68.315 178.355 69.325 178.525 ;
        RECT 69.495 178.510 70.245 178.700 ;
        RECT 67.975 178.015 69.100 178.185 ;
        RECT 69.495 177.845 69.665 178.510 ;
        RECT 70.415 178.265 70.755 179.075 ;
        RECT 71.865 178.815 72.200 179.065 ;
        RECT 72.370 178.695 72.540 179.255 ;
        RECT 73.225 179.235 74.325 179.415 ;
        RECT 74.495 179.450 74.745 179.820 ;
        RECT 74.915 179.575 75.360 179.745 ;
        RECT 75.530 179.715 75.750 179.760 ;
        RECT 72.710 178.815 73.045 179.085 ;
        RECT 74.495 179.065 74.665 179.450 ;
        RECT 72.365 178.655 72.540 178.695 ;
        RECT 67.635 177.675 69.665 177.845 ;
        RECT 69.835 177.505 70.005 178.265 ;
        RECT 70.240 177.855 70.755 178.265 ;
        RECT 71.845 177.505 72.105 178.645 ;
        RECT 72.275 177.675 72.605 178.655 ;
        RECT 72.775 177.505 73.055 178.645 ;
        RECT 73.225 178.495 73.570 179.065 ;
        RECT 73.740 178.815 74.300 179.065 ;
        RECT 74.470 178.895 74.665 179.065 ;
        RECT 73.225 177.505 73.570 178.325 ;
        RECT 73.740 177.715 73.915 178.815 ;
        RECT 74.470 178.645 74.640 178.895 ;
        RECT 74.915 178.785 75.085 179.575 ;
        RECT 75.530 179.545 75.755 179.715 ;
        RECT 75.530 179.405 75.750 179.545 ;
        RECT 75.255 179.235 75.750 179.405 ;
        RECT 76.030 179.390 76.200 180.055 ;
        RECT 76.395 179.315 76.735 179.885 ;
        RECT 77.455 179.575 77.625 180.055 ;
        RECT 77.795 179.405 78.125 179.875 ;
        RECT 75.255 179.040 75.430 179.235 ;
        RECT 75.600 178.865 76.050 179.065 ;
        RECT 74.085 178.255 74.640 178.645 ;
        RECT 74.810 178.645 75.085 178.785 ;
        RECT 76.220 178.695 76.390 179.145 ;
        RECT 74.810 178.425 75.825 178.645 ;
        RECT 75.995 178.525 76.390 178.695 ;
        RECT 75.995 178.255 76.165 178.525 ;
        RECT 76.560 178.355 76.735 179.315 ;
        RECT 76.505 178.345 76.735 178.355 ;
        RECT 74.085 178.085 76.165 178.255 ;
        RECT 74.085 177.850 74.415 178.085 ;
        RECT 74.705 177.505 75.105 177.905 ;
        RECT 75.975 177.505 76.305 177.905 ;
        RECT 76.475 177.675 76.735 178.345 ;
        RECT 77.365 179.235 78.125 179.405 ;
        RECT 78.295 179.235 78.465 180.055 ;
        RECT 78.635 179.405 78.965 179.870 ;
        RECT 79.135 179.585 79.305 180.055 ;
        RECT 79.565 179.675 80.750 179.845 ;
        RECT 80.920 179.505 81.250 179.885 ;
        RECT 79.950 179.405 80.335 179.495 ;
        RECT 78.635 179.235 80.335 179.405 ;
        RECT 80.705 179.335 81.250 179.505 ;
        RECT 77.365 178.265 77.675 179.235 ;
        RECT 77.845 178.855 78.175 179.065 ;
        RECT 78.345 178.855 78.785 179.065 ;
        RECT 78.955 178.855 79.440 179.065 ;
        RECT 78.005 178.685 78.175 178.855 ;
        RECT 78.005 178.515 78.965 178.685 ;
        RECT 77.365 178.095 78.125 178.265 ;
        RECT 77.365 177.505 77.705 177.925 ;
        RECT 77.875 177.675 78.125 178.095 ;
        RECT 78.295 177.505 78.625 178.345 ;
        RECT 78.795 178.265 78.965 178.515 ;
        RECT 79.135 178.435 79.440 178.855 ;
        RECT 79.630 178.865 80.020 179.065 ;
        RECT 80.190 178.865 80.535 179.065 ;
        RECT 79.630 178.435 79.920 178.865 ;
        RECT 80.705 178.695 80.875 179.335 ;
        RECT 81.965 179.285 84.555 180.055 ;
        RECT 81.075 178.815 81.335 179.165 ;
        RECT 80.090 178.645 80.875 178.695 ;
        RECT 80.090 178.470 81.170 178.645 ;
        RECT 80.090 178.265 80.260 178.470 ;
        RECT 78.795 178.095 80.260 178.265 ;
        RECT 79.115 177.675 79.870 178.095 ;
        RECT 80.430 177.505 80.670 178.290 ;
        RECT 80.840 177.675 81.170 178.470 ;
        RECT 81.965 178.595 83.175 179.115 ;
        RECT 83.345 178.765 84.555 179.285 ;
        RECT 84.735 179.330 85.065 179.840 ;
        RECT 85.235 179.655 85.565 180.055 ;
        RECT 86.615 179.485 86.945 179.825 ;
        RECT 87.115 179.655 87.445 180.055 ;
        RECT 81.965 177.505 84.555 178.595 ;
        RECT 84.735 178.565 84.925 179.330 ;
        RECT 85.235 179.315 87.600 179.485 ;
        RECT 87.945 179.330 88.235 180.055 ;
        RECT 85.235 179.145 85.405 179.315 ;
        RECT 85.095 178.815 85.405 179.145 ;
        RECT 85.575 178.815 85.880 179.145 ;
        RECT 84.735 177.715 85.065 178.565 ;
        RECT 85.235 177.505 85.485 178.645 ;
        RECT 85.665 178.485 85.880 178.815 ;
        RECT 86.055 178.485 86.340 179.145 ;
        RECT 86.535 178.485 86.800 179.145 ;
        RECT 87.015 178.485 87.260 179.145 ;
        RECT 87.430 178.315 87.600 179.315 ;
        RECT 89.325 179.255 89.635 180.055 ;
        RECT 89.840 179.255 90.535 179.885 ;
        RECT 90.705 179.285 92.375 180.055 ;
        RECT 89.335 178.815 89.670 179.085 ;
        RECT 85.675 178.145 86.965 178.315 ;
        RECT 85.675 177.725 85.925 178.145 ;
        RECT 86.155 177.505 86.485 177.975 ;
        RECT 86.715 177.725 86.965 178.145 ;
        RECT 87.145 178.145 87.600 178.315 ;
        RECT 87.145 177.715 87.475 178.145 ;
        RECT 87.945 177.505 88.235 178.670 ;
        RECT 89.840 178.655 90.010 179.255 ;
        RECT 90.180 178.815 90.515 179.065 ;
        RECT 89.325 177.505 89.605 178.645 ;
        RECT 89.775 177.675 90.105 178.655 ;
        RECT 90.275 177.505 90.535 178.645 ;
        RECT 90.705 178.595 91.455 179.115 ;
        RECT 91.625 178.765 92.375 179.285 ;
        RECT 92.820 179.245 93.065 179.850 ;
        RECT 93.285 179.520 93.795 180.055 ;
        RECT 92.545 179.075 93.775 179.245 ;
        RECT 90.705 177.505 92.375 178.595 ;
        RECT 92.545 178.265 92.885 179.075 ;
        RECT 93.055 178.510 93.805 178.700 ;
        RECT 92.545 177.855 93.060 178.265 ;
        RECT 93.295 177.505 93.465 178.265 ;
        RECT 93.635 177.845 93.805 178.510 ;
        RECT 93.975 178.525 94.165 179.885 ;
        RECT 94.335 179.715 94.610 179.885 ;
        RECT 94.335 179.545 94.615 179.715 ;
        RECT 94.335 178.725 94.610 179.545 ;
        RECT 94.800 179.520 95.330 179.885 ;
        RECT 95.755 179.655 96.085 180.055 ;
        RECT 95.155 179.485 95.330 179.520 ;
        RECT 94.815 178.525 94.985 179.325 ;
        RECT 93.975 178.355 94.985 178.525 ;
        RECT 95.155 179.315 96.085 179.485 ;
        RECT 96.255 179.315 96.510 179.885 ;
        RECT 95.155 178.185 95.325 179.315 ;
        RECT 95.915 179.145 96.085 179.315 ;
        RECT 94.200 178.015 95.325 178.185 ;
        RECT 95.495 178.815 95.690 179.145 ;
        RECT 95.915 178.815 96.170 179.145 ;
        RECT 95.495 177.845 95.665 178.815 ;
        RECT 96.340 178.645 96.510 179.315 ;
        RECT 96.685 179.305 97.895 180.055 ;
        RECT 93.635 177.675 95.665 177.845 ;
        RECT 95.835 177.505 96.005 178.645 ;
        RECT 96.175 177.675 96.510 178.645 ;
        RECT 96.685 178.595 97.205 179.135 ;
        RECT 97.375 178.765 97.895 179.305 ;
        RECT 96.685 177.505 97.895 178.595 ;
        RECT 98.075 177.685 98.335 179.875 ;
        RECT 98.595 179.685 99.265 180.055 ;
        RECT 99.445 179.505 99.755 179.875 ;
        RECT 98.525 179.305 99.755 179.505 ;
        RECT 98.525 178.635 98.815 179.305 ;
        RECT 99.935 179.125 100.165 179.765 ;
        RECT 100.345 179.325 100.635 180.055 ;
        RECT 100.850 179.665 101.180 180.055 ;
        RECT 101.350 179.495 101.575 179.875 ;
        RECT 98.995 178.815 99.460 179.125 ;
        RECT 99.640 178.815 100.165 179.125 ;
        RECT 100.345 178.815 100.645 179.145 ;
        RECT 100.835 178.815 101.075 179.465 ;
        RECT 101.245 179.315 101.575 179.495 ;
        RECT 101.245 178.645 101.420 179.315 ;
        RECT 101.775 179.145 102.005 179.765 ;
        RECT 102.185 179.325 102.485 180.055 ;
        RECT 103.585 179.255 103.895 180.055 ;
        RECT 104.100 179.255 104.795 179.885 ;
        RECT 105.425 179.255 106.120 179.885 ;
        RECT 106.325 179.255 106.635 180.055 ;
        RECT 106.805 179.255 107.095 180.055 ;
        RECT 107.265 179.595 107.815 179.885 ;
        RECT 107.985 179.595 108.235 180.055 ;
        RECT 101.590 178.815 102.005 179.145 ;
        RECT 102.185 178.815 102.480 179.145 ;
        RECT 103.595 178.815 103.930 179.085 ;
        RECT 104.100 178.655 104.270 179.255 ;
        RECT 104.440 178.815 104.775 179.065 ;
        RECT 105.445 178.815 105.780 179.065 ;
        RECT 105.950 178.695 106.120 179.255 ;
        RECT 106.290 178.815 106.625 179.085 ;
        RECT 105.945 178.655 106.120 178.695 ;
        RECT 98.525 178.415 99.295 178.635 ;
        RECT 98.505 177.505 98.845 178.235 ;
        RECT 99.025 177.685 99.295 178.415 ;
        RECT 99.475 178.395 100.635 178.635 ;
        RECT 99.475 177.685 99.705 178.395 ;
        RECT 99.875 177.505 100.205 178.215 ;
        RECT 100.375 177.685 100.635 178.395 ;
        RECT 100.835 178.455 101.420 178.645 ;
        RECT 100.835 177.685 101.110 178.455 ;
        RECT 101.590 178.285 102.485 178.615 ;
        RECT 101.280 178.115 102.485 178.285 ;
        RECT 101.280 177.685 101.610 178.115 ;
        RECT 101.780 177.505 101.975 177.945 ;
        RECT 102.155 177.685 102.485 178.115 ;
        RECT 103.585 177.505 103.865 178.645 ;
        RECT 104.035 177.675 104.365 178.655 ;
        RECT 104.535 177.505 104.795 178.645 ;
        RECT 105.425 177.505 105.685 178.645 ;
        RECT 105.855 177.675 106.185 178.655 ;
        RECT 106.355 177.505 106.635 178.645 ;
        RECT 106.805 177.505 107.095 178.645 ;
        RECT 107.265 178.225 107.515 179.595 ;
        RECT 108.865 179.425 109.195 179.785 ;
        RECT 107.805 179.235 109.195 179.425 ;
        RECT 109.840 179.245 110.085 179.850 ;
        RECT 110.305 179.520 110.815 180.055 ;
        RECT 107.805 179.145 107.975 179.235 ;
        RECT 107.685 178.815 107.975 179.145 ;
        RECT 109.565 179.075 110.795 179.245 ;
        RECT 108.145 178.815 108.475 179.065 ;
        RECT 108.705 178.815 109.395 179.065 ;
        RECT 107.805 178.565 107.975 178.815 ;
        RECT 107.805 178.395 108.745 178.565 ;
        RECT 107.265 177.675 107.715 178.225 ;
        RECT 107.905 177.505 108.235 178.225 ;
        RECT 108.445 177.845 108.745 178.395 ;
        RECT 109.080 178.375 109.395 178.815 ;
        RECT 109.565 178.265 109.905 179.075 ;
        RECT 110.075 178.510 110.825 178.700 ;
        RECT 108.915 177.505 109.195 178.175 ;
        RECT 109.565 177.855 110.080 178.265 ;
        RECT 110.315 177.505 110.485 178.265 ;
        RECT 110.655 177.845 110.825 178.510 ;
        RECT 110.995 178.525 111.185 179.885 ;
        RECT 111.355 179.715 111.630 179.885 ;
        RECT 111.355 179.545 111.635 179.715 ;
        RECT 111.355 178.725 111.630 179.545 ;
        RECT 111.820 179.520 112.350 179.885 ;
        RECT 112.775 179.655 113.105 180.055 ;
        RECT 112.175 179.485 112.350 179.520 ;
        RECT 111.835 178.525 112.005 179.325 ;
        RECT 110.995 178.355 112.005 178.525 ;
        RECT 112.175 179.315 113.105 179.485 ;
        RECT 113.275 179.315 113.530 179.885 ;
        RECT 113.705 179.330 113.995 180.055 ;
        RECT 114.165 179.445 114.505 179.860 ;
        RECT 114.675 179.615 114.845 180.055 ;
        RECT 115.015 179.665 116.265 179.845 ;
        RECT 115.015 179.445 115.345 179.665 ;
        RECT 116.535 179.595 116.705 180.055 ;
        RECT 112.175 178.185 112.345 179.315 ;
        RECT 112.935 179.145 113.105 179.315 ;
        RECT 111.220 178.015 112.345 178.185 ;
        RECT 112.515 178.815 112.710 179.145 ;
        RECT 112.935 178.815 113.190 179.145 ;
        RECT 112.515 177.845 112.685 178.815 ;
        RECT 113.360 178.645 113.530 179.315 ;
        RECT 114.165 179.275 115.345 179.445 ;
        RECT 115.515 179.425 115.880 179.495 ;
        RECT 115.515 179.245 116.765 179.425 ;
        RECT 114.165 178.865 114.630 179.065 ;
        RECT 114.805 178.815 115.135 179.065 ;
        RECT 115.305 179.035 115.770 179.065 ;
        RECT 115.305 178.865 115.775 179.035 ;
        RECT 115.305 178.815 115.770 178.865 ;
        RECT 115.965 178.815 116.320 179.065 ;
        RECT 114.805 178.695 114.985 178.815 ;
        RECT 110.655 177.675 112.685 177.845 ;
        RECT 112.855 177.505 113.025 178.645 ;
        RECT 113.195 177.675 113.530 178.645 ;
        RECT 113.705 177.505 113.995 178.670 ;
        RECT 114.165 177.505 114.485 178.685 ;
        RECT 114.655 178.525 114.985 178.695 ;
        RECT 116.490 178.645 116.765 179.245 ;
        RECT 114.655 177.735 114.855 178.525 ;
        RECT 115.155 178.435 116.765 178.645 ;
        RECT 115.155 178.335 115.565 178.435 ;
        RECT 115.180 177.675 115.565 178.335 ;
        RECT 115.960 177.505 116.745 178.265 ;
        RECT 116.935 177.675 117.215 179.775 ;
        RECT 117.385 179.285 119.975 180.055 ;
        RECT 120.150 179.510 125.495 180.055 ;
        RECT 117.385 178.595 118.595 179.115 ;
        RECT 118.765 178.765 119.975 179.285 ;
        RECT 117.385 177.505 119.975 178.595 ;
        RECT 121.740 177.940 122.090 179.190 ;
        RECT 123.570 178.680 123.910 179.510 ;
        RECT 125.665 179.305 126.875 180.055 ;
        RECT 125.665 178.595 126.185 179.135 ;
        RECT 126.355 178.765 126.875 179.305 ;
        RECT 120.150 177.505 125.495 177.940 ;
        RECT 125.665 177.505 126.875 178.595 ;
        RECT 14.260 177.335 126.960 177.505 ;
        RECT 14.345 176.245 15.555 177.335 ;
        RECT 14.345 175.535 14.865 176.075 ;
        RECT 15.035 175.705 15.555 176.245 ;
        RECT 15.730 176.185 15.990 177.335 ;
        RECT 16.165 176.260 16.420 177.165 ;
        RECT 16.590 176.575 16.920 177.335 ;
        RECT 17.135 176.405 17.305 177.165 ;
        RECT 14.345 174.785 15.555 175.535 ;
        RECT 15.730 174.785 15.990 175.625 ;
        RECT 16.165 175.530 16.335 176.260 ;
        RECT 16.590 176.235 17.305 176.405 ;
        RECT 16.590 176.025 16.760 176.235 ;
        RECT 17.565 176.180 17.905 177.165 ;
        RECT 18.075 176.905 18.485 177.335 ;
        RECT 19.230 176.915 19.560 177.335 ;
        RECT 19.730 176.735 20.055 177.165 ;
        RECT 18.075 176.565 20.055 176.735 ;
        RECT 16.505 175.695 16.760 176.025 ;
        RECT 16.165 174.955 16.420 175.530 ;
        RECT 16.590 175.505 16.760 175.695 ;
        RECT 17.040 175.685 17.395 176.055 ;
        RECT 17.565 175.525 17.820 176.180 ;
        RECT 18.075 176.025 18.340 176.565 ;
        RECT 18.555 176.225 19.180 176.395 ;
        RECT 17.990 175.695 18.340 176.025 ;
        RECT 18.510 175.695 18.840 176.025 ;
        RECT 19.010 175.525 19.180 176.225 ;
        RECT 16.590 175.335 17.305 175.505 ;
        RECT 16.590 174.785 16.920 175.165 ;
        RECT 17.135 174.955 17.305 175.335 ;
        RECT 17.565 175.150 17.925 175.525 ;
        RECT 18.190 174.785 18.360 175.525 ;
        RECT 18.640 175.355 19.180 175.525 ;
        RECT 19.350 176.155 20.055 176.565 ;
        RECT 20.530 176.235 20.860 177.335 ;
        RECT 22.245 176.405 22.425 177.165 ;
        RECT 22.605 176.575 22.935 177.335 ;
        RECT 22.245 176.235 22.920 176.405 ;
        RECT 23.105 176.260 23.375 177.165 ;
        RECT 18.640 175.150 18.810 175.355 ;
        RECT 19.350 174.955 19.520 176.155 ;
        RECT 22.750 176.090 22.920 176.235 ;
        RECT 19.690 175.775 20.260 175.985 ;
        RECT 20.430 175.775 21.075 175.985 ;
        RECT 22.185 175.685 22.525 176.055 ;
        RECT 22.750 175.760 23.025 176.090 ;
        RECT 19.750 175.435 20.920 175.605 ;
        RECT 22.750 175.505 22.920 175.760 ;
        RECT 19.750 174.955 20.080 175.435 ;
        RECT 20.250 174.785 20.420 175.255 ;
        RECT 20.590 174.970 20.920 175.435 ;
        RECT 22.255 175.335 22.920 175.505 ;
        RECT 23.195 175.460 23.375 176.260 ;
        RECT 23.545 176.170 23.835 177.335 ;
        RECT 24.925 176.365 25.185 177.335 ;
        RECT 22.255 174.955 22.425 175.335 ;
        RECT 22.605 174.785 22.935 175.165 ;
        RECT 23.115 174.955 23.375 175.460 ;
        RECT 23.545 174.785 23.835 175.510 ;
        RECT 24.925 175.075 25.165 176.025 ;
        RECT 25.355 175.990 25.685 177.165 ;
        RECT 25.855 176.365 26.135 177.335 ;
        RECT 26.755 176.535 26.925 177.335 ;
        RECT 27.095 176.315 27.425 177.165 ;
        RECT 27.595 176.535 27.765 177.335 ;
        RECT 27.935 176.315 28.265 177.165 ;
        RECT 28.435 176.535 28.605 177.335 ;
        RECT 28.775 176.315 29.105 177.165 ;
        RECT 29.275 176.535 29.445 177.335 ;
        RECT 29.615 176.315 29.945 177.165 ;
        RECT 30.115 176.485 30.285 177.335 ;
        RECT 30.455 176.315 30.785 177.165 ;
        RECT 30.955 176.485 31.125 177.335 ;
        RECT 31.295 176.315 31.625 177.165 ;
        RECT 26.305 176.145 29.945 176.315 ;
        RECT 30.115 176.145 31.625 176.315 ;
        RECT 31.815 176.245 32.145 177.165 ;
        RECT 25.355 175.460 26.135 175.990 ;
        RECT 26.305 175.605 26.690 176.145 ;
        RECT 30.115 175.975 30.285 176.145 ;
        RECT 31.815 175.975 31.985 176.245 ;
        RECT 32.315 176.145 32.485 177.335 ;
        RECT 33.215 176.525 33.510 177.335 ;
        RECT 33.690 176.025 33.935 177.165 ;
        RECT 34.110 176.525 34.370 177.335 ;
        RECT 34.970 177.330 41.245 177.335 ;
        RECT 34.550 176.025 34.800 177.160 ;
        RECT 34.970 176.535 35.230 177.330 ;
        RECT 35.400 176.435 35.660 177.160 ;
        RECT 35.830 176.605 36.090 177.330 ;
        RECT 36.260 176.435 36.520 177.160 ;
        RECT 36.690 176.605 36.950 177.330 ;
        RECT 37.120 176.435 37.380 177.160 ;
        RECT 37.550 176.605 37.810 177.330 ;
        RECT 37.980 176.435 38.240 177.160 ;
        RECT 38.410 176.605 38.655 177.330 ;
        RECT 38.825 176.435 39.085 177.160 ;
        RECT 39.270 176.605 39.515 177.330 ;
        RECT 39.685 176.435 39.945 177.160 ;
        RECT 40.130 176.605 40.375 177.330 ;
        RECT 40.545 176.435 40.805 177.160 ;
        RECT 40.990 176.605 41.245 177.330 ;
        RECT 35.400 176.420 40.805 176.435 ;
        RECT 41.415 176.420 41.705 177.160 ;
        RECT 41.875 176.590 42.145 177.335 ;
        RECT 35.400 176.195 42.145 176.420 ;
        RECT 42.415 176.195 42.745 177.335 ;
        RECT 43.275 176.365 43.605 177.150 ;
        RECT 42.925 176.195 43.605 176.365 ;
        RECT 43.790 176.615 44.125 177.125 ;
        RECT 26.900 175.775 30.285 175.975 ;
        RECT 30.455 175.775 31.985 175.975 ;
        RECT 32.155 175.775 32.575 175.975 ;
        RECT 30.115 175.605 30.285 175.775 ;
        RECT 31.815 175.605 31.985 175.775 ;
        RECT 25.355 174.955 25.680 175.460 ;
        RECT 26.305 175.435 29.945 175.605 ;
        RECT 30.115 175.435 31.625 175.605 ;
        RECT 25.850 174.785 26.135 175.290 ;
        RECT 26.755 174.785 26.925 175.265 ;
        RECT 27.095 174.960 27.425 175.435 ;
        RECT 27.595 174.785 27.765 175.265 ;
        RECT 27.935 174.960 28.265 175.435 ;
        RECT 28.435 174.785 28.605 175.265 ;
        RECT 28.775 174.960 29.105 175.435 ;
        RECT 29.275 174.785 29.445 175.265 ;
        RECT 29.615 174.960 29.945 175.435 ;
        RECT 30.115 174.785 30.285 175.265 ;
        RECT 30.455 174.960 30.785 175.435 ;
        RECT 30.955 174.785 31.125 175.265 ;
        RECT 31.295 174.960 31.625 175.435 ;
        RECT 31.815 174.960 32.145 175.605 ;
        RECT 32.315 174.785 32.485 175.605 ;
        RECT 33.205 175.465 33.520 176.025 ;
        RECT 33.690 175.775 40.810 176.025 ;
        RECT 33.205 174.785 33.510 175.295 ;
        RECT 33.690 174.965 33.940 175.775 ;
        RECT 34.110 174.785 34.370 175.310 ;
        RECT 34.550 174.965 34.800 175.775 ;
        RECT 40.980 175.605 42.145 176.195 ;
        RECT 42.405 175.775 42.755 176.025 ;
        RECT 35.400 175.435 42.145 175.605 ;
        RECT 42.925 175.595 43.095 176.195 ;
        RECT 43.265 175.775 43.615 176.025 ;
        RECT 34.970 174.785 35.230 175.345 ;
        RECT 35.400 174.980 35.660 175.435 ;
        RECT 35.830 174.785 36.090 175.265 ;
        RECT 36.260 174.980 36.520 175.435 ;
        RECT 36.690 174.785 36.950 175.265 ;
        RECT 37.120 174.980 37.380 175.435 ;
        RECT 37.550 174.785 37.795 175.265 ;
        RECT 37.965 174.980 38.240 175.435 ;
        RECT 38.410 174.785 38.655 175.265 ;
        RECT 38.825 174.980 39.085 175.435 ;
        RECT 39.265 174.785 39.515 175.265 ;
        RECT 39.685 174.980 39.945 175.435 ;
        RECT 40.125 174.785 40.375 175.265 ;
        RECT 40.545 174.980 40.805 175.435 ;
        RECT 40.985 174.785 41.245 175.265 ;
        RECT 41.415 174.980 41.675 175.435 ;
        RECT 41.845 174.785 42.145 175.265 ;
        RECT 42.415 174.785 42.685 175.595 ;
        RECT 42.855 174.955 43.185 175.595 ;
        RECT 43.355 174.785 43.595 175.595 ;
        RECT 43.790 175.260 44.045 176.615 ;
        RECT 44.375 176.535 44.705 177.335 ;
        RECT 44.950 176.745 45.235 177.165 ;
        RECT 45.490 176.915 45.820 177.335 ;
        RECT 46.045 176.995 47.205 177.165 ;
        RECT 46.045 176.745 46.375 176.995 ;
        RECT 44.950 176.575 46.375 176.745 ;
        RECT 46.605 176.365 46.775 176.825 ;
        RECT 47.035 176.495 47.205 176.995 ;
        RECT 44.405 176.195 46.775 176.365 ;
        RECT 44.405 176.025 44.575 176.195 ;
        RECT 47.025 176.145 47.235 176.315 ;
        RECT 47.985 176.195 48.195 177.335 ;
        RECT 48.365 176.185 48.695 177.165 ;
        RECT 48.865 176.195 49.095 177.335 ;
        RECT 47.025 176.025 47.230 176.145 ;
        RECT 44.270 175.695 44.575 176.025 ;
        RECT 44.770 175.975 45.020 176.025 ;
        RECT 44.765 175.805 45.020 175.975 ;
        RECT 44.770 175.695 45.020 175.805 ;
        RECT 44.405 175.525 44.575 175.695 ;
        RECT 45.230 175.635 45.500 176.025 ;
        RECT 45.690 175.635 45.980 176.025 ;
        RECT 44.405 175.355 44.965 175.525 ;
        RECT 45.225 175.465 45.500 175.635 ;
        RECT 45.685 175.465 45.980 175.635 ;
        RECT 45.230 175.365 45.500 175.465 ;
        RECT 45.690 175.365 45.980 175.465 ;
        RECT 46.150 175.360 46.570 176.025 ;
        RECT 46.880 175.695 47.230 176.025 ;
        RECT 43.790 175.000 44.125 175.260 ;
        RECT 44.795 175.185 44.965 175.355 ;
        RECT 44.295 174.785 44.625 175.185 ;
        RECT 44.795 175.015 46.410 175.185 ;
        RECT 46.955 174.785 47.285 175.505 ;
        RECT 47.985 174.785 48.195 175.605 ;
        RECT 48.365 175.585 48.615 176.185 ;
        RECT 49.305 176.170 49.595 177.335 ;
        RECT 50.695 176.725 51.025 177.155 ;
        RECT 51.205 176.895 51.400 177.335 ;
        RECT 51.570 176.725 51.900 177.155 ;
        RECT 50.695 176.555 51.900 176.725 ;
        RECT 50.695 176.225 51.590 176.555 ;
        RECT 52.070 176.385 52.345 177.155 ;
        RECT 51.760 176.195 52.345 176.385 ;
        RECT 52.530 176.945 52.865 177.165 ;
        RECT 53.870 176.955 54.225 177.335 ;
        RECT 52.530 176.325 52.785 176.945 ;
        RECT 53.035 176.785 53.265 176.825 ;
        RECT 54.395 176.785 54.645 177.165 ;
        RECT 53.035 176.585 54.645 176.785 ;
        RECT 53.035 176.495 53.220 176.585 ;
        RECT 53.810 176.575 54.645 176.585 ;
        RECT 54.895 176.555 55.145 177.335 ;
        RECT 55.315 176.485 55.575 177.165 ;
        RECT 53.375 176.385 53.705 176.415 ;
        RECT 53.375 176.325 55.175 176.385 ;
        RECT 52.530 176.215 55.235 176.325 ;
        RECT 48.785 175.775 49.115 176.025 ;
        RECT 50.700 175.695 50.995 176.025 ;
        RECT 51.175 175.695 51.590 176.025 ;
        RECT 48.365 174.955 48.695 175.585 ;
        RECT 48.865 174.785 49.095 175.605 ;
        RECT 49.305 174.785 49.595 175.510 ;
        RECT 50.695 174.785 50.995 175.515 ;
        RECT 51.175 175.075 51.405 175.695 ;
        RECT 51.760 175.525 51.935 176.195 ;
        RECT 52.530 176.155 53.705 176.215 ;
        RECT 55.035 176.180 55.235 176.215 ;
        RECT 51.605 175.345 51.935 175.525 ;
        RECT 52.105 175.375 52.345 176.025 ;
        RECT 52.525 175.775 53.015 175.975 ;
        RECT 53.205 175.775 53.680 175.985 ;
        RECT 51.605 174.965 51.830 175.345 ;
        RECT 52.000 174.785 52.330 175.175 ;
        RECT 52.530 174.785 52.985 175.550 ;
        RECT 53.460 175.375 53.680 175.775 ;
        RECT 53.925 175.775 54.255 175.985 ;
        RECT 53.925 175.375 54.135 175.775 ;
        RECT 54.425 175.740 54.835 176.045 ;
        RECT 55.065 175.605 55.235 176.180 ;
        RECT 54.965 175.485 55.235 175.605 ;
        RECT 54.390 175.440 55.235 175.485 ;
        RECT 54.390 175.315 55.145 175.440 ;
        RECT 54.390 175.165 54.560 175.315 ;
        RECT 55.405 175.285 55.575 176.485 ;
        RECT 56.675 176.385 56.950 177.155 ;
        RECT 57.120 176.725 57.450 177.155 ;
        RECT 57.620 176.895 57.815 177.335 ;
        RECT 57.995 176.725 58.325 177.155 ;
        RECT 57.120 176.555 58.325 176.725 ;
        RECT 56.675 176.195 57.260 176.385 ;
        RECT 57.430 176.225 58.325 176.555 ;
        RECT 59.445 176.445 59.705 177.155 ;
        RECT 59.875 176.625 60.205 177.335 ;
        RECT 60.375 176.445 60.605 177.155 ;
        RECT 59.445 176.205 60.605 176.445 ;
        RECT 60.785 176.425 61.055 177.155 ;
        RECT 61.235 176.605 61.575 177.335 ;
        RECT 60.785 176.205 61.555 176.425 ;
        RECT 56.675 175.375 56.915 176.025 ;
        RECT 57.085 175.525 57.260 176.195 ;
        RECT 57.430 175.695 57.845 176.025 ;
        RECT 58.025 175.695 58.320 176.025 ;
        RECT 59.435 175.695 59.735 176.025 ;
        RECT 59.915 175.715 60.440 176.025 ;
        RECT 60.620 175.715 61.085 176.025 ;
        RECT 57.085 175.345 57.415 175.525 ;
        RECT 53.260 174.955 54.560 175.165 ;
        RECT 54.815 174.785 55.145 175.145 ;
        RECT 55.315 174.955 55.575 175.285 ;
        RECT 56.690 174.785 57.020 175.175 ;
        RECT 57.190 174.965 57.415 175.345 ;
        RECT 57.615 175.075 57.845 175.695 ;
        RECT 58.025 174.785 58.325 175.515 ;
        RECT 59.445 174.785 59.735 175.515 ;
        RECT 59.915 175.075 60.145 175.715 ;
        RECT 61.265 175.535 61.555 176.205 ;
        RECT 60.325 175.335 61.555 175.535 ;
        RECT 60.325 174.965 60.635 175.335 ;
        RECT 60.815 174.785 61.485 175.155 ;
        RECT 61.745 174.965 62.005 177.155 ;
        RECT 62.185 176.245 63.855 177.335 ;
        RECT 64.025 176.575 64.540 176.985 ;
        RECT 64.775 176.575 64.945 177.335 ;
        RECT 65.115 176.995 67.145 177.165 ;
        RECT 62.185 175.725 62.935 176.245 ;
        RECT 63.105 175.555 63.855 176.075 ;
        RECT 64.025 175.765 64.365 176.575 ;
        RECT 65.115 176.330 65.285 176.995 ;
        RECT 65.680 176.655 66.805 176.825 ;
        RECT 64.535 176.140 65.285 176.330 ;
        RECT 65.455 176.315 66.465 176.485 ;
        RECT 64.025 175.595 65.255 175.765 ;
        RECT 62.185 174.785 63.855 175.555 ;
        RECT 64.300 174.990 64.545 175.595 ;
        RECT 64.765 174.785 65.275 175.320 ;
        RECT 65.455 174.955 65.645 176.315 ;
        RECT 65.815 175.975 66.090 176.115 ;
        RECT 65.815 175.805 66.095 175.975 ;
        RECT 65.815 174.955 66.090 175.805 ;
        RECT 66.295 175.515 66.465 176.315 ;
        RECT 66.635 175.525 66.805 176.655 ;
        RECT 66.975 176.025 67.145 176.995 ;
        RECT 67.315 176.195 67.485 177.335 ;
        RECT 67.655 176.195 67.990 177.165 ;
        RECT 66.975 175.695 67.170 176.025 ;
        RECT 67.395 175.695 67.650 176.025 ;
        RECT 67.395 175.525 67.565 175.695 ;
        RECT 67.820 175.525 67.990 176.195 ;
        RECT 68.165 176.575 68.680 176.985 ;
        RECT 68.915 176.575 69.085 177.335 ;
        RECT 69.255 176.995 71.285 177.165 ;
        RECT 68.165 175.765 68.505 176.575 ;
        RECT 69.255 176.330 69.425 176.995 ;
        RECT 69.820 176.655 70.945 176.825 ;
        RECT 68.675 176.140 69.425 176.330 ;
        RECT 69.595 176.315 70.605 176.485 ;
        RECT 68.165 175.595 69.395 175.765 ;
        RECT 66.635 175.355 67.565 175.525 ;
        RECT 66.635 175.320 66.810 175.355 ;
        RECT 66.280 174.955 66.810 175.320 ;
        RECT 67.235 174.785 67.565 175.185 ;
        RECT 67.735 174.955 67.990 175.525 ;
        RECT 68.440 174.990 68.685 175.595 ;
        RECT 68.905 174.785 69.415 175.320 ;
        RECT 69.595 174.955 69.785 176.315 ;
        RECT 69.955 175.975 70.230 176.115 ;
        RECT 69.955 175.805 70.235 175.975 ;
        RECT 69.955 174.955 70.230 175.805 ;
        RECT 70.435 175.515 70.605 176.315 ;
        RECT 70.775 175.525 70.945 176.655 ;
        RECT 71.115 176.025 71.285 176.995 ;
        RECT 71.455 176.195 71.625 177.335 ;
        RECT 71.795 176.195 72.130 177.165 ;
        RECT 71.115 175.695 71.310 176.025 ;
        RECT 71.535 175.695 71.790 176.025 ;
        RECT 71.535 175.525 71.705 175.695 ;
        RECT 71.960 175.525 72.130 176.195 ;
        RECT 72.305 176.245 74.895 177.335 ;
        RECT 72.305 175.725 73.515 176.245 ;
        RECT 75.065 176.170 75.355 177.335 ;
        RECT 75.525 176.245 78.115 177.335 ;
        RECT 73.685 175.555 74.895 176.075 ;
        RECT 75.525 175.725 76.735 176.245 ;
        RECT 76.905 175.555 78.115 176.075 ;
        RECT 78.285 176.015 78.490 177.055 ;
        RECT 78.660 176.195 78.915 177.335 ;
        RECT 79.140 176.025 79.430 177.070 ;
        RECT 79.605 176.725 79.935 177.165 ;
        RECT 80.145 176.955 80.475 177.335 ;
        RECT 80.660 176.725 80.940 177.165 ;
        RECT 81.145 176.895 81.765 177.335 ;
        RECT 79.605 176.485 81.770 176.725 ;
        RECT 78.285 175.705 78.970 176.015 ;
        RECT 79.140 175.695 79.500 176.025 ;
        RECT 79.700 175.775 80.120 176.315 ;
        RECT 70.775 175.355 71.705 175.525 ;
        RECT 70.775 175.320 70.950 175.355 ;
        RECT 70.420 174.955 70.950 175.320 ;
        RECT 71.375 174.785 71.705 175.185 ;
        RECT 71.875 174.955 72.130 175.525 ;
        RECT 72.305 174.785 74.895 175.555 ;
        RECT 75.065 174.785 75.355 175.510 ;
        RECT 75.525 174.785 78.115 175.555 ;
        RECT 80.410 175.635 80.795 176.315 ;
        RECT 80.965 175.775 81.295 176.315 ;
        RECT 78.585 175.325 79.935 175.525 ;
        RECT 78.585 174.955 78.915 175.325 ;
        RECT 79.085 174.785 79.415 175.155 ;
        RECT 79.605 174.955 79.935 175.325 ;
        RECT 80.410 175.465 80.815 175.635 ;
        RECT 81.495 175.585 81.770 176.485 ;
        RECT 80.410 174.955 80.795 175.465 ;
        RECT 80.995 175.415 81.770 175.585 ;
        RECT 80.995 174.955 81.325 175.415 ;
        RECT 81.515 174.785 81.765 175.245 ;
        RECT 81.945 174.955 82.285 177.165 ;
        RECT 82.455 176.195 82.665 177.335 ;
        RECT 82.455 174.785 82.665 175.585 ;
        RECT 82.895 174.965 83.155 177.155 ;
        RECT 83.325 176.605 83.665 177.335 ;
        RECT 83.845 176.425 84.115 177.155 ;
        RECT 83.345 176.205 84.115 176.425 ;
        RECT 84.295 176.445 84.525 177.155 ;
        RECT 84.695 176.625 85.025 177.335 ;
        RECT 85.195 176.445 85.455 177.155 ;
        RECT 84.295 176.205 85.455 176.445 ;
        RECT 83.345 175.535 83.635 176.205 ;
        RECT 86.565 176.195 86.845 177.335 ;
        RECT 87.015 176.185 87.345 177.165 ;
        RECT 87.515 176.195 87.775 177.335 ;
        RECT 88.405 176.575 88.920 176.985 ;
        RECT 89.155 176.575 89.325 177.335 ;
        RECT 89.495 176.995 91.525 177.165 ;
        RECT 83.815 175.715 84.280 176.025 ;
        RECT 84.460 175.715 84.985 176.025 ;
        RECT 83.345 175.335 84.575 175.535 ;
        RECT 83.415 174.785 84.085 175.155 ;
        RECT 84.265 174.965 84.575 175.335 ;
        RECT 84.755 175.075 84.985 175.715 ;
        RECT 85.165 175.695 85.465 176.025 ;
        RECT 86.575 175.755 86.910 176.025 ;
        RECT 87.080 175.635 87.250 176.185 ;
        RECT 87.420 175.775 87.755 176.025 ;
        RECT 88.405 175.765 88.745 176.575 ;
        RECT 89.495 176.330 89.665 176.995 ;
        RECT 90.060 176.655 91.185 176.825 ;
        RECT 88.915 176.140 89.665 176.330 ;
        RECT 89.835 176.315 90.845 176.485 ;
        RECT 87.080 175.585 87.255 175.635 ;
        RECT 88.405 175.595 89.635 175.765 ;
        RECT 85.165 174.785 85.455 175.515 ;
        RECT 86.565 174.785 86.875 175.585 ;
        RECT 87.080 174.955 87.775 175.585 ;
        RECT 88.680 174.990 88.925 175.595 ;
        RECT 89.145 174.785 89.655 175.320 ;
        RECT 89.835 174.955 90.025 176.315 ;
        RECT 90.195 175.975 90.470 176.115 ;
        RECT 90.195 175.805 90.475 175.975 ;
        RECT 90.195 174.955 90.470 175.805 ;
        RECT 90.675 175.515 90.845 176.315 ;
        RECT 91.015 175.525 91.185 176.655 ;
        RECT 91.355 176.025 91.525 176.995 ;
        RECT 91.695 176.195 91.865 177.335 ;
        RECT 92.035 176.195 92.370 177.165 ;
        RECT 91.355 175.695 91.550 176.025 ;
        RECT 91.775 175.695 92.030 176.025 ;
        RECT 91.775 175.525 91.945 175.695 ;
        RECT 92.200 175.525 92.370 176.195 ;
        RECT 92.545 176.575 93.060 176.985 ;
        RECT 93.295 176.575 93.465 177.335 ;
        RECT 93.635 176.995 95.665 177.165 ;
        RECT 92.545 175.765 92.885 176.575 ;
        RECT 93.635 176.330 93.805 176.995 ;
        RECT 94.200 176.655 95.325 176.825 ;
        RECT 93.055 176.140 93.805 176.330 ;
        RECT 93.975 176.315 94.985 176.485 ;
        RECT 92.545 175.595 93.775 175.765 ;
        RECT 91.015 175.355 91.945 175.525 ;
        RECT 91.015 175.320 91.190 175.355 ;
        RECT 90.660 174.955 91.190 175.320 ;
        RECT 91.615 174.785 91.945 175.185 ;
        RECT 92.115 174.955 92.370 175.525 ;
        RECT 92.820 174.990 93.065 175.595 ;
        RECT 93.285 174.785 93.795 175.320 ;
        RECT 93.975 174.955 94.165 176.315 ;
        RECT 94.335 175.975 94.610 176.115 ;
        RECT 94.335 175.805 94.615 175.975 ;
        RECT 94.335 174.955 94.610 175.805 ;
        RECT 94.815 175.515 94.985 176.315 ;
        RECT 95.155 175.525 95.325 176.655 ;
        RECT 95.495 176.025 95.665 176.995 ;
        RECT 95.835 176.195 96.005 177.335 ;
        RECT 96.175 176.195 96.510 177.165 ;
        RECT 95.495 175.695 95.690 176.025 ;
        RECT 95.915 175.695 96.170 176.025 ;
        RECT 95.915 175.525 96.085 175.695 ;
        RECT 96.340 175.525 96.510 176.195 ;
        RECT 96.685 176.155 97.005 177.335 ;
        RECT 97.175 176.315 97.375 177.105 ;
        RECT 97.700 176.505 98.085 177.165 ;
        RECT 98.480 176.575 99.265 177.335 ;
        RECT 97.675 176.405 98.085 176.505 ;
        RECT 97.175 176.145 97.505 176.315 ;
        RECT 97.675 176.195 99.285 176.405 ;
        RECT 97.325 176.025 97.505 176.145 ;
        RECT 96.685 175.775 97.150 175.975 ;
        RECT 97.325 175.775 97.655 176.025 ;
        RECT 97.825 175.975 98.290 176.025 ;
        RECT 97.825 175.805 98.295 175.975 ;
        RECT 97.825 175.775 98.290 175.805 ;
        RECT 98.485 175.775 98.840 176.025 ;
        RECT 99.010 175.595 99.285 176.195 ;
        RECT 95.155 175.355 96.085 175.525 ;
        RECT 95.155 175.320 95.330 175.355 ;
        RECT 94.800 174.955 95.330 175.320 ;
        RECT 95.755 174.785 96.085 175.185 ;
        RECT 96.255 174.955 96.510 175.525 ;
        RECT 96.685 175.395 97.865 175.565 ;
        RECT 96.685 174.980 97.025 175.395 ;
        RECT 97.195 174.785 97.365 175.225 ;
        RECT 97.535 175.175 97.865 175.395 ;
        RECT 98.035 175.415 99.285 175.595 ;
        RECT 98.035 175.345 98.400 175.415 ;
        RECT 97.535 174.995 98.785 175.175 ;
        RECT 99.055 174.785 99.225 175.245 ;
        RECT 99.455 175.065 99.735 177.165 ;
        RECT 100.825 176.170 101.115 177.335 ;
        RECT 101.320 176.545 101.855 177.165 ;
        RECT 101.320 175.525 101.635 176.545 ;
        RECT 102.025 176.535 102.355 177.335 ;
        RECT 103.620 176.545 104.155 177.165 ;
        RECT 102.840 176.365 103.230 176.540 ;
        RECT 101.805 176.195 103.230 176.365 ;
        RECT 101.805 175.695 101.975 176.195 ;
        RECT 100.825 174.785 101.115 175.510 ;
        RECT 101.320 174.955 101.935 175.525 ;
        RECT 102.225 175.465 102.490 176.025 ;
        RECT 102.660 175.295 102.830 176.195 ;
        RECT 103.000 175.465 103.355 176.025 ;
        RECT 103.620 175.525 103.935 176.545 ;
        RECT 104.325 176.535 104.655 177.335 ;
        RECT 105.140 176.365 105.530 176.540 ;
        RECT 104.105 176.195 105.530 176.365 ;
        RECT 105.885 176.245 108.475 177.335 ;
        RECT 108.645 176.575 109.160 176.985 ;
        RECT 109.395 176.575 109.565 177.335 ;
        RECT 109.735 176.995 111.765 177.165 ;
        RECT 104.105 175.695 104.275 176.195 ;
        RECT 102.105 174.785 102.320 175.295 ;
        RECT 102.550 174.965 102.830 175.295 ;
        RECT 103.010 174.785 103.250 175.295 ;
        RECT 103.620 174.955 104.235 175.525 ;
        RECT 104.525 175.465 104.790 176.025 ;
        RECT 104.960 175.295 105.130 176.195 ;
        RECT 105.300 175.465 105.655 176.025 ;
        RECT 105.885 175.725 107.095 176.245 ;
        RECT 107.265 175.555 108.475 176.075 ;
        RECT 108.645 175.765 108.985 176.575 ;
        RECT 109.735 176.330 109.905 176.995 ;
        RECT 110.300 176.655 111.425 176.825 ;
        RECT 109.155 176.140 109.905 176.330 ;
        RECT 110.075 176.315 111.085 176.485 ;
        RECT 108.645 175.595 109.875 175.765 ;
        RECT 104.405 174.785 104.620 175.295 ;
        RECT 104.850 174.965 105.130 175.295 ;
        RECT 105.310 174.785 105.550 175.295 ;
        RECT 105.885 174.785 108.475 175.555 ;
        RECT 108.920 174.990 109.165 175.595 ;
        RECT 109.385 174.785 109.895 175.320 ;
        RECT 110.075 174.955 110.265 176.315 ;
        RECT 110.435 175.295 110.710 176.115 ;
        RECT 110.915 175.515 111.085 176.315 ;
        RECT 111.255 175.525 111.425 176.655 ;
        RECT 111.595 176.025 111.765 176.995 ;
        RECT 111.935 176.195 112.105 177.335 ;
        RECT 112.275 176.195 112.610 177.165 ;
        RECT 111.595 175.695 111.790 176.025 ;
        RECT 112.015 175.695 112.270 176.025 ;
        RECT 112.015 175.525 112.185 175.695 ;
        RECT 112.440 175.525 112.610 176.195 ;
        RECT 113.245 176.245 115.835 177.335 ;
        RECT 116.010 176.900 121.355 177.335 ;
        RECT 113.245 175.725 114.455 176.245 ;
        RECT 114.625 175.555 115.835 176.075 ;
        RECT 117.600 175.650 117.950 176.900 ;
        RECT 121.615 176.405 121.785 177.165 ;
        RECT 121.965 176.575 122.295 177.335 ;
        RECT 121.615 176.235 122.280 176.405 ;
        RECT 122.465 176.260 122.735 177.165 ;
        RECT 111.255 175.355 112.185 175.525 ;
        RECT 111.255 175.320 111.430 175.355 ;
        RECT 110.435 175.125 110.715 175.295 ;
        RECT 110.435 174.955 110.710 175.125 ;
        RECT 110.900 174.955 111.430 175.320 ;
        RECT 111.855 174.785 112.185 175.185 ;
        RECT 112.355 174.955 112.610 175.525 ;
        RECT 113.245 174.785 115.835 175.555 ;
        RECT 119.430 175.330 119.770 176.160 ;
        RECT 122.110 176.090 122.280 176.235 ;
        RECT 121.545 175.685 121.875 176.055 ;
        RECT 122.110 175.760 122.395 176.090 ;
        RECT 122.110 175.505 122.280 175.760 ;
        RECT 121.615 175.335 122.280 175.505 ;
        RECT 122.565 175.460 122.735 176.260 ;
        RECT 122.905 176.245 125.495 177.335 ;
        RECT 125.665 176.245 126.875 177.335 ;
        RECT 122.905 175.725 124.115 176.245 ;
        RECT 124.285 175.555 125.495 176.075 ;
        RECT 125.665 175.705 126.185 176.245 ;
        RECT 116.010 174.785 121.355 175.330 ;
        RECT 121.615 174.955 121.785 175.335 ;
        RECT 121.965 174.785 122.295 175.165 ;
        RECT 122.475 174.955 122.735 175.460 ;
        RECT 122.905 174.785 125.495 175.555 ;
        RECT 126.355 175.535 126.875 176.075 ;
        RECT 125.665 174.785 126.875 175.535 ;
        RECT 14.260 174.615 126.960 174.785 ;
        RECT 14.345 173.865 15.555 174.615 ;
        RECT 15.735 173.885 16.035 174.615 ;
        RECT 14.345 173.325 14.865 173.865 ;
        RECT 16.215 173.705 16.445 174.325 ;
        RECT 16.645 174.055 16.870 174.435 ;
        RECT 17.040 174.225 17.370 174.615 ;
        RECT 16.645 173.875 16.975 174.055 ;
        RECT 15.035 173.155 15.555 173.695 ;
        RECT 15.740 173.375 16.035 173.705 ;
        RECT 16.215 173.375 16.630 173.705 ;
        RECT 16.800 173.205 16.975 173.875 ;
        RECT 17.145 173.375 17.385 174.025 ;
        RECT 17.720 173.965 18.050 174.430 ;
        RECT 18.220 174.145 18.390 174.615 ;
        RECT 18.560 173.965 18.890 174.445 ;
        RECT 17.720 173.795 18.890 173.965 ;
        RECT 17.565 173.415 18.210 173.625 ;
        RECT 18.380 173.415 18.950 173.625 ;
        RECT 19.120 173.245 19.290 174.445 ;
        RECT 19.830 174.045 20.000 174.250 ;
        RECT 14.345 172.065 15.555 173.155 ;
        RECT 15.735 172.845 16.630 173.175 ;
        RECT 16.800 173.015 17.385 173.205 ;
        RECT 15.735 172.675 16.940 172.845 ;
        RECT 15.735 172.245 16.065 172.675 ;
        RECT 16.245 172.065 16.440 172.505 ;
        RECT 16.610 172.245 16.940 172.675 ;
        RECT 17.110 172.245 17.385 173.015 ;
        RECT 17.780 172.065 18.110 173.165 ;
        RECT 18.585 172.835 19.290 173.245 ;
        RECT 19.460 173.875 20.000 174.045 ;
        RECT 20.280 173.875 20.450 174.615 ;
        RECT 20.845 174.250 21.015 174.275 ;
        RECT 20.715 173.875 21.075 174.250 ;
        RECT 19.460 173.175 19.630 173.875 ;
        RECT 19.800 173.375 20.130 173.705 ;
        RECT 20.300 173.375 20.650 173.705 ;
        RECT 19.460 173.005 20.085 173.175 ;
        RECT 20.300 172.835 20.565 173.375 ;
        RECT 20.820 173.220 21.075 173.875 ;
        RECT 21.250 173.775 21.510 174.615 ;
        RECT 21.685 173.870 21.940 174.445 ;
        RECT 22.110 174.235 22.440 174.615 ;
        RECT 22.655 174.065 22.825 174.445 ;
        RECT 23.635 174.135 23.935 174.615 ;
        RECT 22.110 173.895 22.825 174.065 ;
        RECT 24.105 173.965 24.365 174.420 ;
        RECT 24.535 174.135 24.795 174.615 ;
        RECT 24.975 173.965 25.235 174.420 ;
        RECT 25.405 174.135 25.655 174.615 ;
        RECT 25.835 173.965 26.095 174.420 ;
        RECT 26.265 174.135 26.515 174.615 ;
        RECT 26.695 173.965 26.955 174.420 ;
        RECT 27.125 174.135 27.370 174.615 ;
        RECT 27.540 173.965 27.815 174.420 ;
        RECT 27.985 174.135 28.230 174.615 ;
        RECT 28.400 173.965 28.660 174.420 ;
        RECT 28.830 174.135 29.090 174.615 ;
        RECT 29.260 173.965 29.520 174.420 ;
        RECT 29.690 174.135 29.950 174.615 ;
        RECT 30.120 173.965 30.380 174.420 ;
        RECT 30.550 174.055 30.810 174.615 ;
        RECT 18.585 172.665 20.565 172.835 ;
        RECT 18.585 172.235 18.910 172.665 ;
        RECT 19.080 172.065 19.410 172.485 ;
        RECT 20.155 172.065 20.565 172.495 ;
        RECT 20.735 172.235 21.075 173.220 ;
        RECT 21.250 172.065 21.510 173.215 ;
        RECT 21.685 173.140 21.855 173.870 ;
        RECT 22.110 173.705 22.280 173.895 ;
        RECT 23.635 173.795 30.380 173.965 ;
        RECT 22.025 173.375 22.280 173.705 ;
        RECT 22.110 173.165 22.280 173.375 ;
        RECT 22.560 173.345 22.915 173.715 ;
        RECT 23.635 173.205 24.800 173.795 ;
        RECT 30.980 173.625 31.230 174.435 ;
        RECT 31.410 174.090 31.670 174.615 ;
        RECT 31.840 173.625 32.090 174.435 ;
        RECT 32.270 174.105 32.575 174.615 ;
        RECT 33.865 173.985 34.195 174.345 ;
        RECT 34.825 174.155 35.075 174.615 ;
        RECT 35.245 174.155 35.795 174.445 ;
        RECT 24.970 173.375 32.090 173.625 ;
        RECT 32.260 173.375 32.575 173.935 ;
        RECT 33.865 173.795 35.255 173.985 ;
        RECT 35.085 173.705 35.255 173.795 ;
        RECT 33.665 173.375 34.355 173.625 ;
        RECT 34.585 173.375 34.915 173.625 ;
        RECT 35.085 173.375 35.375 173.705 ;
        RECT 21.685 172.235 21.940 173.140 ;
        RECT 22.110 172.995 22.825 173.165 ;
        RECT 22.110 172.065 22.440 172.825 ;
        RECT 22.655 172.235 22.825 172.995 ;
        RECT 23.635 172.980 30.380 173.205 ;
        RECT 23.635 172.065 23.905 172.810 ;
        RECT 24.075 172.240 24.365 172.980 ;
        RECT 24.975 172.965 30.380 172.980 ;
        RECT 24.535 172.070 24.790 172.795 ;
        RECT 24.975 172.240 25.235 172.965 ;
        RECT 25.405 172.070 25.650 172.795 ;
        RECT 25.835 172.240 26.095 172.965 ;
        RECT 26.265 172.070 26.510 172.795 ;
        RECT 26.695 172.240 26.955 172.965 ;
        RECT 27.125 172.070 27.370 172.795 ;
        RECT 27.540 172.240 27.800 172.965 ;
        RECT 27.970 172.070 28.230 172.795 ;
        RECT 28.400 172.240 28.660 172.965 ;
        RECT 28.830 172.070 29.090 172.795 ;
        RECT 29.260 172.240 29.520 172.965 ;
        RECT 29.690 172.070 29.950 172.795 ;
        RECT 30.120 172.240 30.380 172.965 ;
        RECT 30.550 172.070 30.810 172.865 ;
        RECT 30.980 172.240 31.230 173.375 ;
        RECT 24.535 172.065 30.810 172.070 ;
        RECT 31.410 172.065 31.670 172.875 ;
        RECT 31.845 172.235 32.090 173.375 ;
        RECT 33.665 172.935 33.980 173.375 ;
        RECT 35.085 173.125 35.255 173.375 ;
        RECT 34.315 172.955 35.255 173.125 ;
        RECT 32.270 172.065 32.565 172.875 ;
        RECT 33.865 172.065 34.145 172.735 ;
        RECT 34.315 172.405 34.615 172.955 ;
        RECT 35.545 172.785 35.795 174.155 ;
        RECT 35.965 173.815 36.255 174.615 ;
        RECT 36.425 173.890 36.715 174.615 ;
        RECT 37.435 174.065 37.605 174.445 ;
        RECT 37.785 174.235 38.115 174.615 ;
        RECT 37.435 173.895 38.100 174.065 ;
        RECT 38.295 173.940 38.555 174.445 ;
        RECT 37.365 173.345 37.695 173.715 ;
        RECT 37.930 173.640 38.100 173.895 ;
        RECT 37.930 173.310 38.215 173.640 ;
        RECT 34.825 172.065 35.155 172.785 ;
        RECT 35.345 172.235 35.795 172.785 ;
        RECT 35.965 172.065 36.255 173.205 ;
        RECT 36.425 172.065 36.715 173.230 ;
        RECT 37.930 173.165 38.100 173.310 ;
        RECT 37.435 172.995 38.100 173.165 ;
        RECT 38.385 173.140 38.555 173.940 ;
        RECT 38.925 173.985 39.255 174.345 ;
        RECT 39.875 174.155 40.125 174.615 ;
        RECT 40.295 174.155 40.855 174.445 ;
        RECT 41.135 174.235 42.305 174.445 ;
        RECT 41.135 174.215 41.465 174.235 ;
        RECT 38.925 173.795 40.315 173.985 ;
        RECT 40.145 173.705 40.315 173.795 ;
        RECT 37.435 172.235 37.605 172.995 ;
        RECT 37.785 172.065 38.115 172.825 ;
        RECT 38.285 172.235 38.555 173.140 ;
        RECT 38.740 173.375 39.415 173.625 ;
        RECT 39.635 173.375 39.975 173.625 ;
        RECT 40.145 173.375 40.435 173.705 ;
        RECT 38.740 173.015 39.005 173.375 ;
        RECT 40.145 173.125 40.315 173.375 ;
        RECT 39.375 172.955 40.315 173.125 ;
        RECT 38.925 172.065 39.205 172.735 ;
        RECT 39.375 172.405 39.675 172.955 ;
        RECT 40.605 172.785 40.855 174.155 ;
        RECT 41.025 173.795 41.885 174.045 ;
        RECT 42.055 173.985 42.305 174.235 ;
        RECT 42.475 174.155 42.645 174.615 ;
        RECT 42.815 173.985 43.155 174.445 ;
        RECT 42.055 173.815 43.155 173.985 ;
        RECT 43.415 173.965 43.585 174.445 ;
        RECT 43.755 174.135 44.085 174.615 ;
        RECT 44.255 173.965 44.425 174.440 ;
        RECT 44.595 174.135 44.925 174.615 ;
        RECT 45.095 173.965 45.265 174.445 ;
        RECT 45.435 174.135 45.765 174.615 ;
        RECT 45.935 173.965 46.105 174.445 ;
        RECT 46.275 174.135 46.605 174.615 ;
        RECT 46.775 173.965 46.945 174.445 ;
        RECT 47.115 174.135 47.445 174.615 ;
        RECT 47.615 173.965 47.785 174.445 ;
        RECT 43.415 173.795 44.835 173.965 ;
        RECT 45.095 173.795 47.785 173.965 ;
        RECT 47.955 173.815 48.285 174.615 ;
        RECT 49.765 173.940 50.025 174.445 ;
        RECT 50.205 174.235 50.535 174.615 ;
        RECT 50.715 174.065 50.885 174.445 ;
        RECT 41.025 173.205 41.305 173.795 ;
        RECT 44.660 173.625 44.835 173.795 ;
        RECT 41.475 173.375 42.225 173.625 ;
        RECT 42.395 173.375 43.155 173.625 ;
        RECT 43.380 173.425 44.480 173.625 ;
        RECT 44.660 173.455 47.285 173.625 ;
        RECT 47.530 173.595 47.785 173.795 ;
        RECT 44.660 173.255 44.835 173.455 ;
        RECT 47.525 173.425 47.785 173.595 ;
        RECT 47.530 173.255 47.785 173.425 ;
        RECT 41.025 173.035 42.725 173.205 ;
        RECT 39.875 172.065 40.205 172.785 ;
        RECT 40.395 172.235 40.855 172.785 ;
        RECT 41.130 172.065 41.385 172.865 ;
        RECT 41.555 172.235 41.885 173.035 ;
        RECT 42.055 172.065 42.225 172.865 ;
        RECT 42.395 172.235 42.725 173.035 ;
        RECT 42.895 172.065 43.155 173.205 ;
        RECT 43.335 173.085 44.835 173.255 ;
        RECT 45.095 173.085 47.785 173.255 ;
        RECT 43.335 172.235 43.665 173.085 ;
        RECT 43.835 172.065 44.005 172.865 ;
        RECT 44.175 172.235 44.505 173.085 ;
        RECT 44.675 172.065 44.845 172.865 ;
        RECT 45.095 172.235 45.265 173.085 ;
        RECT 45.435 172.065 45.765 172.865 ;
        RECT 45.935 172.235 46.105 173.085 ;
        RECT 46.275 172.065 46.605 172.865 ;
        RECT 46.775 172.235 46.945 173.085 ;
        RECT 47.115 172.065 47.445 172.865 ;
        RECT 47.615 172.235 47.785 173.085 ;
        RECT 47.955 172.065 48.285 173.215 ;
        RECT 49.765 173.140 49.935 173.940 ;
        RECT 50.220 173.895 50.885 174.065 ;
        RECT 50.220 173.640 50.390 173.895 ;
        RECT 51.165 173.805 51.405 174.615 ;
        RECT 51.575 173.805 51.905 174.445 ;
        RECT 52.075 173.805 52.345 174.615 ;
        RECT 50.105 173.310 50.390 173.640 ;
        RECT 50.625 173.345 50.955 173.715 ;
        RECT 51.145 173.375 51.495 173.625 ;
        RECT 50.220 173.165 50.390 173.310 ;
        RECT 51.665 173.205 51.835 173.805 ;
        RECT 52.585 173.795 52.795 174.615 ;
        RECT 52.965 173.815 53.295 174.445 ;
        RECT 52.005 173.375 52.355 173.625 ;
        RECT 52.965 173.215 53.215 173.815 ;
        RECT 53.465 173.795 53.695 174.615 ;
        RECT 53.905 174.155 54.465 174.445 ;
        RECT 54.635 174.155 54.885 174.615 ;
        RECT 53.385 173.375 53.715 173.625 ;
        RECT 49.765 172.235 50.035 173.140 ;
        RECT 50.220 172.995 50.885 173.165 ;
        RECT 50.205 172.065 50.535 172.825 ;
        RECT 50.715 172.235 50.885 172.995 ;
        RECT 51.155 173.035 51.835 173.205 ;
        RECT 51.155 172.250 51.485 173.035 ;
        RECT 52.015 172.065 52.345 173.205 ;
        RECT 52.585 172.065 52.795 173.205 ;
        RECT 52.965 172.235 53.295 173.215 ;
        RECT 53.465 172.065 53.695 173.205 ;
        RECT 53.905 172.785 54.155 174.155 ;
        RECT 55.505 173.985 55.835 174.345 ;
        RECT 56.830 174.105 57.070 174.615 ;
        RECT 57.250 174.105 57.530 174.435 ;
        RECT 57.760 174.105 57.975 174.615 ;
        RECT 54.445 173.795 55.835 173.985 ;
        RECT 54.445 173.705 54.615 173.795 ;
        RECT 54.325 173.375 54.615 173.705 ;
        RECT 54.785 173.375 55.125 173.625 ;
        RECT 55.345 173.375 56.020 173.625 ;
        RECT 56.725 173.375 57.080 173.935 ;
        RECT 54.445 173.125 54.615 173.375 ;
        RECT 54.445 172.955 55.385 173.125 ;
        RECT 55.755 173.015 56.020 173.375 ;
        RECT 57.250 173.205 57.420 174.105 ;
        RECT 57.590 173.375 57.855 173.935 ;
        RECT 58.145 173.875 58.760 174.445 ;
        RECT 58.105 173.205 58.275 173.705 ;
        RECT 56.850 173.035 58.275 173.205 ;
        RECT 53.905 172.235 54.365 172.785 ;
        RECT 54.555 172.065 54.885 172.785 ;
        RECT 55.085 172.405 55.385 172.955 ;
        RECT 56.850 172.860 57.240 173.035 ;
        RECT 55.555 172.065 55.835 172.735 ;
        RECT 57.725 172.065 58.055 172.865 ;
        RECT 58.445 172.855 58.760 173.875 ;
        RECT 58.225 172.235 58.760 172.855 ;
        RECT 58.965 174.155 59.525 174.445 ;
        RECT 59.695 174.155 59.945 174.615 ;
        RECT 58.965 172.785 59.215 174.155 ;
        RECT 60.565 173.985 60.895 174.345 ;
        RECT 59.505 173.795 60.895 173.985 ;
        RECT 62.185 173.890 62.475 174.615 ;
        RECT 62.645 173.940 62.905 174.445 ;
        RECT 63.085 174.235 63.415 174.615 ;
        RECT 63.595 174.065 63.765 174.445 ;
        RECT 59.505 173.705 59.675 173.795 ;
        RECT 59.385 173.375 59.675 173.705 ;
        RECT 59.845 173.375 60.185 173.625 ;
        RECT 60.405 173.375 61.080 173.625 ;
        RECT 59.505 173.125 59.675 173.375 ;
        RECT 59.505 172.955 60.445 173.125 ;
        RECT 60.815 173.015 61.080 173.375 ;
        RECT 58.965 172.235 59.425 172.785 ;
        RECT 59.615 172.065 59.945 172.785 ;
        RECT 60.145 172.405 60.445 172.955 ;
        RECT 60.615 172.065 60.895 172.735 ;
        RECT 62.185 172.065 62.475 173.230 ;
        RECT 62.645 173.140 62.815 173.940 ;
        RECT 63.100 173.895 63.765 174.065 ;
        RECT 63.100 173.640 63.270 173.895 ;
        RECT 64.085 173.795 64.295 174.615 ;
        RECT 64.465 173.815 64.795 174.445 ;
        RECT 62.985 173.310 63.270 173.640 ;
        RECT 63.505 173.345 63.835 173.715 ;
        RECT 63.100 173.165 63.270 173.310 ;
        RECT 64.465 173.215 64.715 173.815 ;
        RECT 64.965 173.795 65.195 174.615 ;
        RECT 65.865 173.985 66.205 174.445 ;
        RECT 66.375 174.155 66.545 174.615 ;
        RECT 66.715 174.235 67.885 174.445 ;
        RECT 66.715 173.985 66.965 174.235 ;
        RECT 67.555 174.215 67.885 174.235 ;
        RECT 65.865 173.815 66.965 173.985 ;
        RECT 67.135 173.795 67.995 174.045 ;
        RECT 68.165 173.845 70.755 174.615 ;
        RECT 71.090 174.105 71.330 174.615 ;
        RECT 71.510 174.105 71.790 174.435 ;
        RECT 72.020 174.105 72.235 174.615 ;
        RECT 64.885 173.375 65.215 173.625 ;
        RECT 65.865 173.375 66.625 173.625 ;
        RECT 66.795 173.375 67.545 173.625 ;
        RECT 62.645 172.235 62.915 173.140 ;
        RECT 63.100 172.995 63.765 173.165 ;
        RECT 63.085 172.065 63.415 172.825 ;
        RECT 63.595 172.235 63.765 172.995 ;
        RECT 64.085 172.065 64.295 173.205 ;
        RECT 64.465 172.235 64.795 173.215 ;
        RECT 67.715 173.205 67.995 173.795 ;
        RECT 64.965 172.065 65.195 173.205 ;
        RECT 65.865 172.065 66.125 173.205 ;
        RECT 66.295 173.035 67.995 173.205 ;
        RECT 68.165 173.155 69.375 173.675 ;
        RECT 69.545 173.325 70.755 173.845 ;
        RECT 70.985 173.375 71.340 173.935 ;
        RECT 71.510 173.205 71.680 174.105 ;
        RECT 71.850 173.375 72.115 173.935 ;
        RECT 72.405 173.875 73.020 174.445 ;
        RECT 72.365 173.205 72.535 173.705 ;
        RECT 66.295 172.235 66.625 173.035 ;
        RECT 66.795 172.065 66.965 172.865 ;
        RECT 67.135 172.235 67.465 173.035 ;
        RECT 67.635 172.065 67.890 172.865 ;
        RECT 68.165 172.065 70.755 173.155 ;
        RECT 71.110 173.035 72.535 173.205 ;
        RECT 71.110 172.860 71.500 173.035 ;
        RECT 71.985 172.065 72.315 172.865 ;
        RECT 72.705 172.855 73.020 173.875 ;
        RECT 73.225 173.975 73.565 174.380 ;
        RECT 73.735 174.145 73.905 174.615 ;
        RECT 74.075 173.975 74.325 174.380 ;
        RECT 73.225 173.795 74.325 173.975 ;
        RECT 74.495 174.010 74.745 174.380 ;
        RECT 74.915 174.135 75.360 174.305 ;
        RECT 75.530 174.275 75.750 174.320 ;
        RECT 74.495 173.625 74.665 174.010 ;
        RECT 73.225 173.055 73.570 173.625 ;
        RECT 73.740 173.375 74.300 173.625 ;
        RECT 74.470 173.455 74.665 173.625 ;
        RECT 72.485 172.235 73.020 172.855 ;
        RECT 73.225 172.065 73.570 172.885 ;
        RECT 73.740 172.275 73.915 173.375 ;
        RECT 74.470 173.205 74.640 173.455 ;
        RECT 74.915 173.345 75.085 174.135 ;
        RECT 75.530 174.105 75.755 174.275 ;
        RECT 75.530 173.965 75.750 174.105 ;
        RECT 75.255 173.795 75.750 173.965 ;
        RECT 76.030 173.950 76.200 174.615 ;
        RECT 76.395 173.875 76.735 174.445 ;
        RECT 75.255 173.600 75.430 173.795 ;
        RECT 75.600 173.425 76.050 173.625 ;
        RECT 74.085 172.815 74.640 173.205 ;
        RECT 74.810 173.205 75.085 173.345 ;
        RECT 76.220 173.255 76.390 173.705 ;
        RECT 74.810 172.985 75.825 173.205 ;
        RECT 75.995 173.085 76.390 173.255 ;
        RECT 75.995 172.815 76.165 173.085 ;
        RECT 76.560 172.905 76.735 173.875 ;
        RECT 76.905 173.865 78.115 174.615 ;
        RECT 74.085 172.645 76.165 172.815 ;
        RECT 74.085 172.410 74.415 172.645 ;
        RECT 74.705 172.065 75.105 172.465 ;
        RECT 75.975 172.065 76.305 172.465 ;
        RECT 76.475 172.235 76.735 172.905 ;
        RECT 76.905 173.155 77.425 173.695 ;
        RECT 77.595 173.325 78.115 173.865 ;
        RECT 78.305 173.815 78.545 174.615 ;
        RECT 76.905 172.065 78.115 173.155 ;
        RECT 78.290 172.065 78.545 173.065 ;
        RECT 78.730 172.235 78.975 174.445 ;
        RECT 79.145 174.235 79.475 174.615 ;
        RECT 79.665 174.065 79.995 174.445 ;
        RECT 80.545 174.235 80.875 174.615 ;
        RECT 79.145 173.860 79.995 174.065 ;
        RECT 80.165 174.065 80.375 174.235 ;
        RECT 81.045 174.065 81.320 174.205 ;
        RECT 80.165 173.875 81.320 174.065 ;
        RECT 81.595 174.065 81.765 174.445 ;
        RECT 81.945 174.235 82.275 174.615 ;
        RECT 81.595 173.895 82.260 174.065 ;
        RECT 82.455 173.940 82.715 174.445 ;
        RECT 82.910 174.225 83.240 174.615 ;
        RECT 83.410 174.055 83.635 174.435 ;
        RECT 79.145 173.370 79.475 173.860 ;
        RECT 79.305 172.915 79.475 173.370 ;
        RECT 79.645 173.085 80.055 173.690 ;
        RECT 80.225 173.300 80.810 173.675 ;
        RECT 80.605 172.915 80.810 173.300 ;
        RECT 81.065 173.250 81.325 173.705 ;
        RECT 81.525 173.345 81.855 173.715 ;
        RECT 82.090 173.640 82.260 173.895 ;
        RECT 82.090 173.310 82.375 173.640 ;
        RECT 82.090 173.165 82.260 173.310 ;
        RECT 79.305 172.695 80.425 172.915 ;
        RECT 80.605 172.745 80.815 172.915 ;
        RECT 80.605 172.715 80.810 172.745 ;
        RECT 79.145 172.065 79.995 172.515 ;
        RECT 80.165 172.235 80.425 172.695 ;
        RECT 80.995 172.065 81.320 173.050 ;
        RECT 81.595 172.995 82.260 173.165 ;
        RECT 82.545 173.140 82.715 173.940 ;
        RECT 82.895 173.375 83.135 174.025 ;
        RECT 83.305 173.875 83.635 174.055 ;
        RECT 83.305 173.205 83.480 173.875 ;
        RECT 83.835 173.705 84.065 174.325 ;
        RECT 84.245 173.885 84.545 174.615 ;
        RECT 84.815 174.065 84.985 174.445 ;
        RECT 85.200 174.235 85.530 174.615 ;
        RECT 84.815 173.895 85.530 174.065 ;
        RECT 83.650 173.375 84.065 173.705 ;
        RECT 84.245 173.375 84.540 173.705 ;
        RECT 84.725 173.345 85.080 173.715 ;
        RECT 85.360 173.705 85.530 173.895 ;
        RECT 85.700 173.870 85.955 174.445 ;
        RECT 85.360 173.375 85.615 173.705 ;
        RECT 81.595 172.235 81.765 172.995 ;
        RECT 81.945 172.065 82.275 172.825 ;
        RECT 82.445 172.235 82.715 173.140 ;
        RECT 82.895 173.015 83.480 173.205 ;
        RECT 82.895 172.245 83.170 173.015 ;
        RECT 83.650 172.845 84.545 173.175 ;
        RECT 85.360 173.165 85.530 173.375 ;
        RECT 83.340 172.675 84.545 172.845 ;
        RECT 83.340 172.245 83.670 172.675 ;
        RECT 83.840 172.065 84.035 172.505 ;
        RECT 84.215 172.245 84.545 172.675 ;
        RECT 84.815 172.995 85.530 173.165 ;
        RECT 85.785 173.140 85.955 173.870 ;
        RECT 86.130 173.775 86.390 174.615 ;
        RECT 86.565 173.865 87.775 174.615 ;
        RECT 87.945 173.890 88.235 174.615 ;
        RECT 84.815 172.235 84.985 172.995 ;
        RECT 85.200 172.065 85.530 172.825 ;
        RECT 85.700 172.235 85.955 173.140 ;
        RECT 86.130 172.065 86.390 173.215 ;
        RECT 86.565 173.155 87.085 173.695 ;
        RECT 87.255 173.325 87.775 173.865 ;
        RECT 88.865 173.845 90.535 174.615 ;
        RECT 86.565 172.065 87.775 173.155 ;
        RECT 87.945 172.065 88.235 173.230 ;
        RECT 88.865 173.155 89.615 173.675 ;
        RECT 89.785 173.325 90.535 173.845 ;
        RECT 90.705 174.115 90.965 174.445 ;
        RECT 91.175 174.135 91.450 174.615 ;
        RECT 90.705 173.205 90.875 174.115 ;
        RECT 91.660 174.045 91.865 174.445 ;
        RECT 92.035 174.215 92.370 174.615 ;
        RECT 91.045 173.375 91.405 173.955 ;
        RECT 91.660 173.875 92.345 174.045 ;
        RECT 91.585 173.205 91.835 173.705 ;
        RECT 88.865 172.065 90.535 173.155 ;
        RECT 90.705 173.035 91.835 173.205 ;
        RECT 90.705 172.265 90.975 173.035 ;
        RECT 92.005 172.845 92.345 173.875 ;
        RECT 92.820 173.805 93.065 174.410 ;
        RECT 93.285 174.080 93.795 174.615 ;
        RECT 91.145 172.065 91.475 172.845 ;
        RECT 91.680 172.670 92.345 172.845 ;
        RECT 92.545 173.635 93.775 173.805 ;
        RECT 92.545 172.825 92.885 173.635 ;
        RECT 93.055 173.070 93.805 173.260 ;
        RECT 91.680 172.265 91.865 172.670 ;
        RECT 92.035 172.065 92.370 172.490 ;
        RECT 92.545 172.415 93.060 172.825 ;
        RECT 93.295 172.065 93.465 172.825 ;
        RECT 93.635 172.405 93.805 173.070 ;
        RECT 93.975 173.085 94.165 174.445 ;
        RECT 94.335 174.275 94.610 174.445 ;
        RECT 94.335 174.105 94.615 174.275 ;
        RECT 94.335 173.285 94.610 174.105 ;
        RECT 94.800 174.080 95.330 174.445 ;
        RECT 95.755 174.215 96.085 174.615 ;
        RECT 95.155 174.045 95.330 174.080 ;
        RECT 94.815 173.085 94.985 173.885 ;
        RECT 93.975 172.915 94.985 173.085 ;
        RECT 95.155 173.875 96.085 174.045 ;
        RECT 96.255 173.875 96.510 174.445 ;
        RECT 95.155 172.745 95.325 173.875 ;
        RECT 95.915 173.705 96.085 173.875 ;
        RECT 94.200 172.575 95.325 172.745 ;
        RECT 95.495 173.375 95.690 173.705 ;
        RECT 95.915 173.375 96.170 173.705 ;
        RECT 95.495 172.405 95.665 173.375 ;
        RECT 96.340 173.205 96.510 173.875 ;
        RECT 96.685 174.005 97.025 174.420 ;
        RECT 97.195 174.175 97.365 174.615 ;
        RECT 97.535 174.225 98.785 174.405 ;
        RECT 97.535 174.005 97.865 174.225 ;
        RECT 99.055 174.155 99.225 174.615 ;
        RECT 96.685 173.835 97.865 174.005 ;
        RECT 98.035 173.985 98.400 174.055 ;
        RECT 98.035 173.805 99.285 173.985 ;
        RECT 96.685 173.425 97.150 173.625 ;
        RECT 97.325 173.375 97.655 173.625 ;
        RECT 97.825 173.595 98.290 173.625 ;
        RECT 97.825 173.425 98.295 173.595 ;
        RECT 97.825 173.375 98.290 173.425 ;
        RECT 98.485 173.375 98.840 173.625 ;
        RECT 97.325 173.255 97.505 173.375 ;
        RECT 93.635 172.235 95.665 172.405 ;
        RECT 95.835 172.065 96.005 173.205 ;
        RECT 96.175 172.235 96.510 173.205 ;
        RECT 96.685 172.065 97.005 173.245 ;
        RECT 97.175 173.085 97.505 173.255 ;
        RECT 99.010 173.205 99.285 173.805 ;
        RECT 97.175 172.295 97.375 173.085 ;
        RECT 97.675 172.995 99.285 173.205 ;
        RECT 97.675 172.895 98.085 172.995 ;
        RECT 97.700 172.235 98.085 172.895 ;
        RECT 98.480 172.065 99.265 172.825 ;
        RECT 99.455 172.235 99.735 174.335 ;
        RECT 99.915 173.885 100.215 174.615 ;
        RECT 100.395 173.705 100.625 174.325 ;
        RECT 100.825 174.055 101.050 174.435 ;
        RECT 101.220 174.225 101.550 174.615 ;
        RECT 101.770 174.225 102.100 174.615 ;
        RECT 102.270 174.055 102.495 174.435 ;
        RECT 100.825 173.875 101.155 174.055 ;
        RECT 99.920 173.375 100.215 173.705 ;
        RECT 100.395 173.375 100.810 173.705 ;
        RECT 100.980 173.205 101.155 173.875 ;
        RECT 101.325 173.375 101.565 174.025 ;
        RECT 101.755 173.375 101.995 174.025 ;
        RECT 102.165 173.875 102.495 174.055 ;
        RECT 102.165 173.205 102.340 173.875 ;
        RECT 102.695 173.705 102.925 174.325 ;
        RECT 103.105 173.885 103.405 174.615 ;
        RECT 104.045 173.845 105.715 174.615 ;
        RECT 106.050 174.105 106.290 174.615 ;
        RECT 106.470 174.105 106.750 174.435 ;
        RECT 106.980 174.105 107.195 174.615 ;
        RECT 102.510 173.375 102.925 173.705 ;
        RECT 103.105 173.375 103.400 173.705 ;
        RECT 99.915 172.845 100.810 173.175 ;
        RECT 100.980 173.015 101.565 173.205 ;
        RECT 99.915 172.675 101.120 172.845 ;
        RECT 99.915 172.245 100.245 172.675 ;
        RECT 100.425 172.065 100.620 172.505 ;
        RECT 100.790 172.245 101.120 172.675 ;
        RECT 101.290 172.245 101.565 173.015 ;
        RECT 101.755 173.015 102.340 173.205 ;
        RECT 101.755 172.245 102.030 173.015 ;
        RECT 102.510 172.845 103.405 173.175 ;
        RECT 102.200 172.675 103.405 172.845 ;
        RECT 102.200 172.245 102.530 172.675 ;
        RECT 102.700 172.065 102.895 172.505 ;
        RECT 103.075 172.245 103.405 172.675 ;
        RECT 104.045 173.155 104.795 173.675 ;
        RECT 104.965 173.325 105.715 173.845 ;
        RECT 105.945 173.375 106.300 173.935 ;
        RECT 106.470 173.205 106.640 174.105 ;
        RECT 106.810 173.375 107.075 173.935 ;
        RECT 107.365 173.875 107.980 174.445 ;
        RECT 107.325 173.205 107.495 173.705 ;
        RECT 104.045 172.065 105.715 173.155 ;
        RECT 106.070 173.035 107.495 173.205 ;
        RECT 106.070 172.860 106.460 173.035 ;
        RECT 106.945 172.065 107.275 172.865 ;
        RECT 107.665 172.855 107.980 173.875 ;
        RECT 108.460 173.805 108.705 174.410 ;
        RECT 108.925 174.080 109.435 174.615 ;
        RECT 107.445 172.235 107.980 172.855 ;
        RECT 108.185 173.635 109.415 173.805 ;
        RECT 108.185 172.825 108.525 173.635 ;
        RECT 108.695 173.070 109.445 173.260 ;
        RECT 108.185 172.415 108.700 172.825 ;
        RECT 108.935 172.065 109.105 172.825 ;
        RECT 109.275 172.405 109.445 173.070 ;
        RECT 109.615 173.085 109.805 174.445 ;
        RECT 109.975 173.935 110.250 174.445 ;
        RECT 110.440 174.080 110.970 174.445 ;
        RECT 111.395 174.215 111.725 174.615 ;
        RECT 110.795 174.045 110.970 174.080 ;
        RECT 109.975 173.765 110.255 173.935 ;
        RECT 109.975 173.285 110.250 173.765 ;
        RECT 110.455 173.085 110.625 173.885 ;
        RECT 109.615 172.915 110.625 173.085 ;
        RECT 110.795 173.875 111.725 174.045 ;
        RECT 111.895 173.875 112.150 174.445 ;
        RECT 110.795 172.745 110.965 173.875 ;
        RECT 111.555 173.705 111.725 173.875 ;
        RECT 109.840 172.575 110.965 172.745 ;
        RECT 111.135 173.375 111.330 173.705 ;
        RECT 111.555 173.375 111.810 173.705 ;
        RECT 111.135 172.405 111.305 173.375 ;
        RECT 111.980 173.205 112.150 173.875 ;
        RECT 112.325 173.865 113.535 174.615 ;
        RECT 113.705 173.890 113.995 174.615 ;
        RECT 109.275 172.235 111.305 172.405 ;
        RECT 111.475 172.065 111.645 173.205 ;
        RECT 111.815 172.235 112.150 173.205 ;
        RECT 112.325 173.155 112.845 173.695 ;
        RECT 113.015 173.325 113.535 173.865 ;
        RECT 114.165 173.845 115.835 174.615 ;
        RECT 116.010 174.070 121.355 174.615 ;
        RECT 112.325 172.065 113.535 173.155 ;
        RECT 113.705 172.065 113.995 173.230 ;
        RECT 114.165 173.155 114.915 173.675 ;
        RECT 115.085 173.325 115.835 173.845 ;
        RECT 114.165 172.065 115.835 173.155 ;
        RECT 117.600 172.500 117.950 173.750 ;
        RECT 119.430 173.240 119.770 174.070 ;
        RECT 121.615 174.065 121.785 174.445 ;
        RECT 121.965 174.235 122.295 174.615 ;
        RECT 121.615 173.895 122.280 174.065 ;
        RECT 122.475 173.940 122.735 174.445 ;
        RECT 121.545 173.345 121.875 173.715 ;
        RECT 122.110 173.640 122.280 173.895 ;
        RECT 122.110 173.310 122.395 173.640 ;
        RECT 122.110 173.165 122.280 173.310 ;
        RECT 121.615 172.995 122.280 173.165 ;
        RECT 122.565 173.140 122.735 173.940 ;
        RECT 123.915 174.065 124.085 174.445 ;
        RECT 124.300 174.235 124.630 174.615 ;
        RECT 123.915 173.895 124.630 174.065 ;
        RECT 123.825 173.345 124.180 173.715 ;
        RECT 124.460 173.705 124.630 173.895 ;
        RECT 124.800 173.870 125.055 174.445 ;
        RECT 124.460 173.375 124.715 173.705 ;
        RECT 124.460 173.165 124.630 173.375 ;
        RECT 116.010 172.065 121.355 172.500 ;
        RECT 121.615 172.235 121.785 172.995 ;
        RECT 121.965 172.065 122.295 172.825 ;
        RECT 122.465 172.235 122.735 173.140 ;
        RECT 123.915 172.995 124.630 173.165 ;
        RECT 124.885 173.140 125.055 173.870 ;
        RECT 125.230 173.775 125.490 174.615 ;
        RECT 125.665 173.865 126.875 174.615 ;
        RECT 123.915 172.235 124.085 172.995 ;
        RECT 124.300 172.065 124.630 172.825 ;
        RECT 124.800 172.235 125.055 173.140 ;
        RECT 125.230 172.065 125.490 173.215 ;
        RECT 125.665 173.155 126.185 173.695 ;
        RECT 126.355 173.325 126.875 173.865 ;
        RECT 125.665 172.065 126.875 173.155 ;
        RECT 14.260 171.895 126.960 172.065 ;
        RECT 14.345 170.805 15.555 171.895 ;
        RECT 15.725 171.095 15.985 171.895 ;
        RECT 14.345 170.095 14.865 170.635 ;
        RECT 15.035 170.265 15.555 170.805 ;
        RECT 14.345 169.345 15.555 170.095 ;
        RECT 15.725 169.915 15.985 170.925 ;
        RECT 16.245 170.505 16.485 171.710 ;
        RECT 16.655 170.875 16.910 171.710 ;
        RECT 17.515 170.925 17.850 171.710 ;
        RECT 16.655 170.675 17.095 170.875 ;
        RECT 16.245 170.335 16.695 170.505 ;
        RECT 16.865 170.255 17.095 170.675 ;
        RECT 17.265 170.755 17.850 170.925 ;
        RECT 18.025 171.095 18.465 171.725 ;
        RECT 17.265 170.085 17.435 170.755 ;
        RECT 16.235 169.915 17.435 170.085 ;
        RECT 17.605 170.005 17.855 170.585 ;
        RECT 18.025 170.085 18.335 171.095 ;
        RECT 18.640 171.045 18.955 171.895 ;
        RECT 19.125 171.555 20.555 171.725 ;
        RECT 19.125 170.875 19.295 171.555 ;
        RECT 18.505 170.705 19.295 170.875 ;
        RECT 18.505 170.255 18.675 170.705 ;
        RECT 19.465 170.585 19.665 171.385 ;
        RECT 18.845 170.255 19.235 170.535 ;
        RECT 19.420 170.255 19.665 170.585 ;
        RECT 19.865 170.255 20.115 171.385 ;
        RECT 20.305 170.925 20.555 171.555 ;
        RECT 20.735 171.095 21.065 171.895 ;
        RECT 20.305 170.755 21.075 170.925 ;
        RECT 20.330 170.255 20.735 170.585 ;
        RECT 20.905 170.085 21.075 170.755 ;
        RECT 21.710 170.745 21.970 171.895 ;
        RECT 22.145 170.820 22.400 171.725 ;
        RECT 22.570 171.135 22.900 171.895 ;
        RECT 23.115 170.965 23.285 171.725 ;
        RECT 15.735 169.345 16.065 169.745 ;
        RECT 16.235 169.645 16.405 169.915 ;
        RECT 17.080 169.905 17.435 169.915 ;
        RECT 16.575 169.345 16.905 169.745 ;
        RECT 17.080 169.645 17.345 169.905 ;
        RECT 17.595 169.345 17.855 169.835 ;
        RECT 18.025 169.525 18.465 170.085 ;
        RECT 18.635 169.345 19.085 170.085 ;
        RECT 19.255 169.915 20.415 170.085 ;
        RECT 19.255 169.515 19.425 169.915 ;
        RECT 19.595 169.345 20.015 169.745 ;
        RECT 20.185 169.515 20.415 169.915 ;
        RECT 20.585 169.515 21.075 170.085 ;
        RECT 21.710 169.345 21.970 170.185 ;
        RECT 22.145 170.090 22.315 170.820 ;
        RECT 22.570 170.795 23.285 170.965 ;
        RECT 22.570 170.585 22.740 170.795 ;
        RECT 23.545 170.730 23.835 171.895 ;
        RECT 22.485 170.255 22.740 170.585 ;
        RECT 22.145 169.515 22.400 170.090 ;
        RECT 22.570 170.065 22.740 170.255 ;
        RECT 23.020 170.245 23.375 170.615 ;
        RECT 24.005 170.290 24.285 171.725 ;
        RECT 24.455 171.120 25.165 171.895 ;
        RECT 25.335 170.950 25.665 171.725 ;
        RECT 24.515 170.735 25.665 170.950 ;
        RECT 22.570 169.895 23.285 170.065 ;
        RECT 22.570 169.345 22.900 169.725 ;
        RECT 23.115 169.515 23.285 169.895 ;
        RECT 23.545 169.345 23.835 170.070 ;
        RECT 24.005 169.515 24.345 170.290 ;
        RECT 24.515 170.165 24.800 170.735 ;
        RECT 24.985 170.335 25.455 170.565 ;
        RECT 25.860 170.535 26.075 171.650 ;
        RECT 26.255 171.175 26.585 171.895 ;
        RECT 26.845 170.965 27.025 171.725 ;
        RECT 27.205 171.135 27.535 171.895 ;
        RECT 26.365 170.535 26.595 170.875 ;
        RECT 26.845 170.795 27.520 170.965 ;
        RECT 27.705 170.820 27.975 171.725 ;
        RECT 27.350 170.650 27.520 170.795 ;
        RECT 25.625 170.355 26.075 170.535 ;
        RECT 25.625 170.335 25.955 170.355 ;
        RECT 26.265 170.335 26.595 170.535 ;
        RECT 26.785 170.245 27.125 170.615 ;
        RECT 27.350 170.320 27.625 170.650 ;
        RECT 24.515 169.975 25.225 170.165 ;
        RECT 24.925 169.835 25.225 169.975 ;
        RECT 25.415 169.975 26.595 170.165 ;
        RECT 27.350 170.065 27.520 170.320 ;
        RECT 25.415 169.895 25.745 169.975 ;
        RECT 24.925 169.825 25.240 169.835 ;
        RECT 24.925 169.815 25.250 169.825 ;
        RECT 24.925 169.810 25.260 169.815 ;
        RECT 24.515 169.345 24.685 169.805 ;
        RECT 24.925 169.800 25.265 169.810 ;
        RECT 24.925 169.795 25.270 169.800 ;
        RECT 24.925 169.785 25.275 169.795 ;
        RECT 24.925 169.780 25.280 169.785 ;
        RECT 24.925 169.515 25.285 169.780 ;
        RECT 25.915 169.345 26.085 169.805 ;
        RECT 26.255 169.515 26.595 169.975 ;
        RECT 26.855 169.895 27.520 170.065 ;
        RECT 27.795 170.020 27.975 170.820 ;
        RECT 28.235 170.965 28.405 171.725 ;
        RECT 28.585 171.135 28.915 171.895 ;
        RECT 28.235 170.795 28.900 170.965 ;
        RECT 29.085 170.820 29.355 171.725 ;
        RECT 28.730 170.650 28.900 170.795 ;
        RECT 28.165 170.245 28.495 170.615 ;
        RECT 28.730 170.320 29.015 170.650 ;
        RECT 28.730 170.065 28.900 170.320 ;
        RECT 26.855 169.515 27.025 169.895 ;
        RECT 27.205 169.345 27.535 169.725 ;
        RECT 27.715 169.515 27.975 170.020 ;
        RECT 28.235 169.895 28.900 170.065 ;
        RECT 29.185 170.020 29.355 170.820 ;
        RECT 29.565 170.755 29.795 171.895 ;
        RECT 29.965 170.745 30.295 171.725 ;
        RECT 30.465 170.755 30.675 171.895 ;
        RECT 30.905 170.755 31.195 171.895 ;
        RECT 31.365 171.175 31.815 171.725 ;
        RECT 32.005 171.175 32.335 171.895 ;
        RECT 29.545 170.335 29.875 170.585 ;
        RECT 28.235 169.515 28.405 169.895 ;
        RECT 28.585 169.345 28.915 169.725 ;
        RECT 29.095 169.515 29.355 170.020 ;
        RECT 29.565 169.345 29.795 170.165 ;
        RECT 30.045 170.145 30.295 170.745 ;
        RECT 29.965 169.515 30.295 170.145 ;
        RECT 30.465 169.345 30.675 170.165 ;
        RECT 30.905 169.345 31.195 170.145 ;
        RECT 31.365 169.805 31.615 171.175 ;
        RECT 32.545 171.005 32.845 171.555 ;
        RECT 33.015 171.225 33.295 171.895 ;
        RECT 31.905 170.835 32.845 171.005 ;
        RECT 31.905 170.585 32.075 170.835 ;
        RECT 33.180 170.585 33.495 171.025 ;
        RECT 33.755 170.965 33.925 171.725 ;
        RECT 34.140 171.135 34.470 171.895 ;
        RECT 33.755 170.795 34.470 170.965 ;
        RECT 34.640 170.820 34.895 171.725 ;
        RECT 31.785 170.255 32.075 170.585 ;
        RECT 32.245 170.335 32.575 170.585 ;
        RECT 32.805 170.335 33.495 170.585 ;
        RECT 31.905 170.165 32.075 170.255 ;
        RECT 33.665 170.245 34.020 170.615 ;
        RECT 34.300 170.585 34.470 170.795 ;
        RECT 34.300 170.255 34.555 170.585 ;
        RECT 31.905 169.975 33.295 170.165 ;
        RECT 34.300 170.065 34.470 170.255 ;
        RECT 34.725 170.090 34.895 170.820 ;
        RECT 35.070 170.745 35.330 171.895 ;
        RECT 36.425 170.730 36.715 171.895 ;
        RECT 36.885 171.175 37.345 171.725 ;
        RECT 37.535 171.175 37.865 171.895 ;
        RECT 31.365 169.515 31.915 169.805 ;
        RECT 32.085 169.345 32.335 169.805 ;
        RECT 32.965 169.615 33.295 169.975 ;
        RECT 33.755 169.895 34.470 170.065 ;
        RECT 33.755 169.515 33.925 169.895 ;
        RECT 34.140 169.345 34.470 169.725 ;
        RECT 34.640 169.515 34.895 170.090 ;
        RECT 35.070 169.345 35.330 170.185 ;
        RECT 36.425 169.345 36.715 170.070 ;
        RECT 36.885 169.805 37.135 171.175 ;
        RECT 38.065 171.005 38.365 171.555 ;
        RECT 38.535 171.225 38.815 171.895 ;
        RECT 37.425 170.835 38.365 171.005 ;
        RECT 37.425 170.585 37.595 170.835 ;
        RECT 38.735 170.585 39.000 170.945 ;
        RECT 39.370 170.925 39.760 171.100 ;
        RECT 40.245 171.095 40.575 171.895 ;
        RECT 40.745 171.105 41.280 171.725 ;
        RECT 39.370 170.755 40.795 170.925 ;
        RECT 37.305 170.255 37.595 170.585 ;
        RECT 37.765 170.335 38.105 170.585 ;
        RECT 38.325 170.335 39.000 170.585 ;
        RECT 37.425 170.165 37.595 170.255 ;
        RECT 37.425 169.975 38.815 170.165 ;
        RECT 39.245 170.025 39.600 170.585 ;
        RECT 36.885 169.515 37.445 169.805 ;
        RECT 37.615 169.345 37.865 169.805 ;
        RECT 38.485 169.615 38.815 169.975 ;
        RECT 39.770 169.855 39.940 170.755 ;
        RECT 40.110 170.025 40.375 170.585 ;
        RECT 40.625 170.255 40.795 170.755 ;
        RECT 40.965 170.085 41.280 171.105 ;
        RECT 42.035 170.965 42.205 171.725 ;
        RECT 42.385 171.135 42.715 171.895 ;
        RECT 42.035 170.795 42.700 170.965 ;
        RECT 42.885 170.820 43.155 171.725 ;
        RECT 42.530 170.650 42.700 170.795 ;
        RECT 41.965 170.245 42.295 170.615 ;
        RECT 42.530 170.320 42.815 170.650 ;
        RECT 39.350 169.345 39.590 169.855 ;
        RECT 39.770 169.525 40.050 169.855 ;
        RECT 40.280 169.345 40.495 169.855 ;
        RECT 40.665 169.515 41.280 170.085 ;
        RECT 42.530 170.065 42.700 170.320 ;
        RECT 42.035 169.895 42.700 170.065 ;
        RECT 42.985 170.020 43.155 170.820 ;
        RECT 43.415 170.965 43.585 171.725 ;
        RECT 43.800 171.135 44.130 171.895 ;
        RECT 43.415 170.795 44.130 170.965 ;
        RECT 44.300 170.820 44.555 171.725 ;
        RECT 43.325 170.245 43.680 170.615 ;
        RECT 43.960 170.585 44.130 170.795 ;
        RECT 43.960 170.255 44.215 170.585 ;
        RECT 43.960 170.065 44.130 170.255 ;
        RECT 44.385 170.090 44.555 170.820 ;
        RECT 44.730 170.745 44.990 171.895 ;
        RECT 45.245 170.965 45.425 171.725 ;
        RECT 45.605 171.135 45.935 171.895 ;
        RECT 45.245 170.795 45.920 170.965 ;
        RECT 46.105 170.820 46.375 171.725 ;
        RECT 45.750 170.650 45.920 170.795 ;
        RECT 45.185 170.245 45.525 170.615 ;
        RECT 45.750 170.320 46.025 170.650 ;
        RECT 42.035 169.515 42.205 169.895 ;
        RECT 42.385 169.345 42.715 169.725 ;
        RECT 42.895 169.515 43.155 170.020 ;
        RECT 43.415 169.895 44.130 170.065 ;
        RECT 43.415 169.515 43.585 169.895 ;
        RECT 43.800 169.345 44.130 169.725 ;
        RECT 44.300 169.515 44.555 170.090 ;
        RECT 44.730 169.345 44.990 170.185 ;
        RECT 45.750 170.065 45.920 170.320 ;
        RECT 45.255 169.895 45.920 170.065 ;
        RECT 46.195 170.020 46.375 170.820 ;
        RECT 46.635 170.965 46.805 171.725 ;
        RECT 47.020 171.135 47.350 171.895 ;
        RECT 46.635 170.795 47.350 170.965 ;
        RECT 47.520 170.820 47.775 171.725 ;
        RECT 46.545 170.245 46.900 170.615 ;
        RECT 47.180 170.585 47.350 170.795 ;
        RECT 47.180 170.255 47.435 170.585 ;
        RECT 47.180 170.065 47.350 170.255 ;
        RECT 47.605 170.090 47.775 170.820 ;
        RECT 47.950 170.745 48.210 171.895 ;
        RECT 49.305 170.730 49.595 171.895 ;
        RECT 49.855 170.965 50.025 171.725 ;
        RECT 50.240 171.135 50.570 171.895 ;
        RECT 49.855 170.795 50.570 170.965 ;
        RECT 50.740 170.820 50.995 171.725 ;
        RECT 49.765 170.245 50.120 170.615 ;
        RECT 50.400 170.585 50.570 170.795 ;
        RECT 50.400 170.255 50.655 170.585 ;
        RECT 45.255 169.515 45.425 169.895 ;
        RECT 45.605 169.345 45.935 169.725 ;
        RECT 46.115 169.515 46.375 170.020 ;
        RECT 46.635 169.895 47.350 170.065 ;
        RECT 46.635 169.515 46.805 169.895 ;
        RECT 47.020 169.345 47.350 169.725 ;
        RECT 47.520 169.515 47.775 170.090 ;
        RECT 47.950 169.345 48.210 170.185 ;
        RECT 49.305 169.345 49.595 170.070 ;
        RECT 50.400 170.065 50.570 170.255 ;
        RECT 50.825 170.090 50.995 170.820 ;
        RECT 51.170 170.745 51.430 171.895 ;
        RECT 51.605 170.820 51.875 171.725 ;
        RECT 52.045 171.135 52.375 171.895 ;
        RECT 52.555 170.965 52.735 171.725 ;
        RECT 49.855 169.895 50.570 170.065 ;
        RECT 49.855 169.515 50.025 169.895 ;
        RECT 50.240 169.345 50.570 169.725 ;
        RECT 50.740 169.515 50.995 170.090 ;
        RECT 51.170 169.345 51.430 170.185 ;
        RECT 51.605 170.020 51.785 170.820 ;
        RECT 52.060 170.795 52.735 170.965 ;
        RECT 53.525 170.965 53.705 171.725 ;
        RECT 53.885 171.135 54.215 171.895 ;
        RECT 53.525 170.795 54.200 170.965 ;
        RECT 54.385 170.820 54.655 171.725 ;
        RECT 52.060 170.650 52.230 170.795 ;
        RECT 51.955 170.320 52.230 170.650 ;
        RECT 54.030 170.650 54.200 170.795 ;
        RECT 52.060 170.065 52.230 170.320 ;
        RECT 52.455 170.245 52.795 170.615 ;
        RECT 53.465 170.245 53.805 170.615 ;
        RECT 54.030 170.320 54.305 170.650 ;
        RECT 54.030 170.065 54.200 170.320 ;
        RECT 51.605 169.515 51.865 170.020 ;
        RECT 52.060 169.895 52.725 170.065 ;
        RECT 52.045 169.345 52.375 169.725 ;
        RECT 52.555 169.515 52.725 169.895 ;
        RECT 53.535 169.895 54.200 170.065 ;
        RECT 54.475 170.020 54.655 170.820 ;
        RECT 53.535 169.515 53.705 169.895 ;
        RECT 53.885 169.345 54.215 169.725 ;
        RECT 54.395 169.515 54.655 170.020 ;
        RECT 54.825 170.820 55.095 171.725 ;
        RECT 55.265 171.135 55.595 171.895 ;
        RECT 55.775 170.965 55.955 171.725 ;
        RECT 54.825 170.020 55.005 170.820 ;
        RECT 55.280 170.795 55.955 170.965 ;
        RECT 55.280 170.650 55.450 170.795 ;
        RECT 56.210 170.745 56.470 171.895 ;
        RECT 56.645 170.820 56.900 171.725 ;
        RECT 57.070 171.135 57.400 171.895 ;
        RECT 57.615 170.965 57.785 171.725 ;
        RECT 55.175 170.320 55.450 170.650 ;
        RECT 55.280 170.065 55.450 170.320 ;
        RECT 55.675 170.245 56.015 170.615 ;
        RECT 54.825 169.515 55.085 170.020 ;
        RECT 55.280 169.895 55.945 170.065 ;
        RECT 55.265 169.345 55.595 169.725 ;
        RECT 55.775 169.515 55.945 169.895 ;
        RECT 56.210 169.345 56.470 170.185 ;
        RECT 56.645 170.090 56.815 170.820 ;
        RECT 57.070 170.795 57.785 170.965 ;
        RECT 58.045 170.820 58.315 171.725 ;
        RECT 58.485 171.135 58.815 171.895 ;
        RECT 58.995 170.965 59.165 171.725 ;
        RECT 57.070 170.585 57.240 170.795 ;
        RECT 56.985 170.255 57.240 170.585 ;
        RECT 56.645 169.515 56.900 170.090 ;
        RECT 57.070 170.065 57.240 170.255 ;
        RECT 57.520 170.245 57.875 170.615 ;
        RECT 57.070 169.895 57.785 170.065 ;
        RECT 57.070 169.345 57.400 169.725 ;
        RECT 57.615 169.515 57.785 169.895 ;
        RECT 58.045 170.020 58.215 170.820 ;
        RECT 58.500 170.795 59.165 170.965 ;
        RECT 58.500 170.650 58.670 170.795 ;
        RECT 60.350 170.745 60.610 171.895 ;
        RECT 60.785 170.820 61.040 171.725 ;
        RECT 61.210 171.135 61.540 171.895 ;
        RECT 61.755 170.965 61.925 171.725 ;
        RECT 58.385 170.320 58.670 170.650 ;
        RECT 58.500 170.065 58.670 170.320 ;
        RECT 58.905 170.245 59.235 170.615 ;
        RECT 58.045 169.515 58.305 170.020 ;
        RECT 58.500 169.895 59.165 170.065 ;
        RECT 58.485 169.345 58.815 169.725 ;
        RECT 58.995 169.515 59.165 169.895 ;
        RECT 60.350 169.345 60.610 170.185 ;
        RECT 60.785 170.090 60.955 170.820 ;
        RECT 61.210 170.795 61.925 170.965 ;
        RECT 61.210 170.585 61.380 170.795 ;
        RECT 62.185 170.730 62.475 171.895 ;
        RECT 63.105 170.755 63.365 171.725 ;
        RECT 63.535 171.470 63.920 171.895 ;
        RECT 64.090 171.300 64.345 171.725 ;
        RECT 63.535 171.105 64.345 171.300 ;
        RECT 61.125 170.255 61.380 170.585 ;
        RECT 60.785 169.515 61.040 170.090 ;
        RECT 61.210 170.065 61.380 170.255 ;
        RECT 61.660 170.245 62.015 170.615 ;
        RECT 63.105 170.085 63.290 170.755 ;
        RECT 63.535 170.585 63.885 171.105 ;
        RECT 64.535 170.935 64.780 171.725 ;
        RECT 64.950 171.470 65.335 171.895 ;
        RECT 65.505 171.300 65.780 171.725 ;
        RECT 63.460 170.255 63.885 170.585 ;
        RECT 64.055 170.755 64.780 170.935 ;
        RECT 64.950 171.105 65.780 171.300 ;
        RECT 64.055 170.255 64.705 170.755 ;
        RECT 64.950 170.585 65.300 171.105 ;
        RECT 65.950 170.935 66.375 171.725 ;
        RECT 66.545 171.470 66.930 171.895 ;
        RECT 67.100 171.300 67.535 171.725 ;
        RECT 64.875 170.255 65.300 170.585 ;
        RECT 65.470 170.755 66.375 170.935 ;
        RECT 66.545 171.130 67.535 171.300 ;
        RECT 65.470 170.255 66.300 170.755 ;
        RECT 66.545 170.585 66.880 171.130 ;
        RECT 66.470 170.255 66.880 170.585 ;
        RECT 67.050 170.255 67.535 170.960 ;
        RECT 67.705 170.820 67.975 171.725 ;
        RECT 68.145 171.135 68.475 171.895 ;
        RECT 68.655 170.965 68.835 171.725 ;
        RECT 63.535 170.085 63.885 170.255 ;
        RECT 64.535 170.085 64.705 170.255 ;
        RECT 64.950 170.085 65.300 170.255 ;
        RECT 65.950 170.085 66.300 170.255 ;
        RECT 66.545 170.085 66.880 170.255 ;
        RECT 61.210 169.895 61.925 170.065 ;
        RECT 61.210 169.345 61.540 169.725 ;
        RECT 61.755 169.515 61.925 169.895 ;
        RECT 62.185 169.345 62.475 170.070 ;
        RECT 63.105 169.515 63.365 170.085 ;
        RECT 63.535 169.915 64.345 170.085 ;
        RECT 63.535 169.345 63.920 169.745 ;
        RECT 64.090 169.515 64.345 169.915 ;
        RECT 64.535 169.515 64.780 170.085 ;
        RECT 64.950 169.915 65.760 170.085 ;
        RECT 64.950 169.345 65.335 169.745 ;
        RECT 65.505 169.515 65.760 169.915 ;
        RECT 65.950 169.515 66.375 170.085 ;
        RECT 66.545 169.915 67.535 170.085 ;
        RECT 66.545 169.345 66.930 169.745 ;
        RECT 67.100 169.515 67.535 169.915 ;
        RECT 67.705 170.020 67.885 170.820 ;
        RECT 68.160 170.795 68.835 170.965 ;
        RECT 68.160 170.650 68.330 170.795 ;
        RECT 68.055 170.320 68.330 170.650 ;
        RECT 68.160 170.065 68.330 170.320 ;
        RECT 68.555 170.245 68.895 170.615 ;
        RECT 67.705 169.515 67.965 170.020 ;
        RECT 68.160 169.895 68.825 170.065 ;
        RECT 68.145 169.345 68.475 169.725 ;
        RECT 68.655 169.515 68.825 169.895 ;
        RECT 69.085 169.515 69.835 171.725 ;
        RECT 70.005 170.820 70.275 171.725 ;
        RECT 70.445 171.135 70.775 171.895 ;
        RECT 70.955 170.965 71.135 171.725 ;
        RECT 70.005 170.020 70.185 170.820 ;
        RECT 70.460 170.795 71.135 170.965 ;
        RECT 71.385 170.805 72.595 171.895 ;
        RECT 72.845 170.965 73.025 171.725 ;
        RECT 73.205 171.135 73.535 171.895 ;
        RECT 70.460 170.650 70.630 170.795 ;
        RECT 70.355 170.320 70.630 170.650 ;
        RECT 70.460 170.065 70.630 170.320 ;
        RECT 70.855 170.245 71.195 170.615 ;
        RECT 71.385 170.265 71.905 170.805 ;
        RECT 72.845 170.795 73.520 170.965 ;
        RECT 73.705 170.820 73.975 171.725 ;
        RECT 73.350 170.650 73.520 170.795 ;
        RECT 72.075 170.095 72.595 170.635 ;
        RECT 72.785 170.245 73.125 170.615 ;
        RECT 73.350 170.320 73.625 170.650 ;
        RECT 70.005 169.515 70.265 170.020 ;
        RECT 70.460 169.895 71.125 170.065 ;
        RECT 70.445 169.345 70.775 169.725 ;
        RECT 70.955 169.515 71.125 169.895 ;
        RECT 71.385 169.345 72.595 170.095 ;
        RECT 73.350 170.065 73.520 170.320 ;
        RECT 72.855 169.895 73.520 170.065 ;
        RECT 73.795 170.020 73.975 170.820 ;
        RECT 75.065 170.730 75.355 171.895 ;
        RECT 75.985 170.820 76.255 171.725 ;
        RECT 76.425 171.135 76.755 171.895 ;
        RECT 76.935 170.965 77.115 171.725 ;
        RECT 72.855 169.515 73.025 169.895 ;
        RECT 73.205 169.345 73.535 169.725 ;
        RECT 73.715 169.515 73.975 170.020 ;
        RECT 75.065 169.345 75.355 170.070 ;
        RECT 75.985 170.020 76.165 170.820 ;
        RECT 76.440 170.795 77.115 170.965 ;
        RECT 78.285 170.805 81.795 171.895 ;
        RECT 82.055 170.965 82.225 171.725 ;
        RECT 82.440 171.135 82.770 171.895 ;
        RECT 76.440 170.650 76.610 170.795 ;
        RECT 76.335 170.320 76.610 170.650 ;
        RECT 76.440 170.065 76.610 170.320 ;
        RECT 76.835 170.245 77.175 170.615 ;
        RECT 78.285 170.285 79.975 170.805 ;
        RECT 82.055 170.795 82.770 170.965 ;
        RECT 82.940 170.820 83.195 171.725 ;
        RECT 80.145 170.115 81.795 170.635 ;
        RECT 81.965 170.245 82.320 170.615 ;
        RECT 82.600 170.585 82.770 170.795 ;
        RECT 82.600 170.255 82.855 170.585 ;
        RECT 75.985 169.515 76.245 170.020 ;
        RECT 76.440 169.895 77.105 170.065 ;
        RECT 76.425 169.345 76.755 169.725 ;
        RECT 76.935 169.515 77.105 169.895 ;
        RECT 78.285 169.345 81.795 170.115 ;
        RECT 82.600 170.065 82.770 170.255 ;
        RECT 83.025 170.090 83.195 170.820 ;
        RECT 83.370 170.745 83.630 171.895 ;
        RECT 83.805 170.805 85.475 171.895 ;
        RECT 85.645 170.820 85.915 171.725 ;
        RECT 86.085 171.135 86.415 171.895 ;
        RECT 86.595 170.965 86.775 171.725 ;
        RECT 83.805 170.285 84.555 170.805 ;
        RECT 82.055 169.895 82.770 170.065 ;
        RECT 82.055 169.515 82.225 169.895 ;
        RECT 82.440 169.345 82.770 169.725 ;
        RECT 82.940 169.515 83.195 170.090 ;
        RECT 83.370 169.345 83.630 170.185 ;
        RECT 84.725 170.115 85.475 170.635 ;
        RECT 83.805 169.345 85.475 170.115 ;
        RECT 85.645 170.020 85.825 170.820 ;
        RECT 86.100 170.795 86.775 170.965 ;
        RECT 86.100 170.650 86.270 170.795 ;
        RECT 87.945 170.730 88.235 171.895 ;
        RECT 88.405 170.805 89.615 171.895 ;
        RECT 89.790 171.460 95.135 171.895 ;
        RECT 95.310 171.460 100.655 171.895 ;
        RECT 85.995 170.320 86.270 170.650 ;
        RECT 86.100 170.065 86.270 170.320 ;
        RECT 86.495 170.245 86.835 170.615 ;
        RECT 88.405 170.265 88.925 170.805 ;
        RECT 89.095 170.095 89.615 170.635 ;
        RECT 91.380 170.210 91.730 171.460 ;
        RECT 85.645 169.515 85.905 170.020 ;
        RECT 86.100 169.895 86.765 170.065 ;
        RECT 86.085 169.345 86.415 169.725 ;
        RECT 86.595 169.515 86.765 169.895 ;
        RECT 87.945 169.345 88.235 170.070 ;
        RECT 88.405 169.345 89.615 170.095 ;
        RECT 93.210 169.890 93.550 170.720 ;
        RECT 96.900 170.210 97.250 171.460 ;
        RECT 100.825 170.730 101.115 171.895 ;
        RECT 101.745 170.805 104.335 171.895 ;
        RECT 104.510 171.460 109.855 171.895 ;
        RECT 98.730 169.890 99.070 170.720 ;
        RECT 101.745 170.285 102.955 170.805 ;
        RECT 103.125 170.115 104.335 170.635 ;
        RECT 106.100 170.210 106.450 171.460 ;
        RECT 89.790 169.345 95.135 169.890 ;
        RECT 95.310 169.345 100.655 169.890 ;
        RECT 100.825 169.345 101.115 170.070 ;
        RECT 101.745 169.345 104.335 170.115 ;
        RECT 107.930 169.890 108.270 170.720 ;
        RECT 104.510 169.345 109.855 169.890 ;
        RECT 110.025 169.625 110.305 171.725 ;
        RECT 110.495 171.135 111.280 171.895 ;
        RECT 111.675 171.065 112.060 171.725 ;
        RECT 111.675 170.965 112.085 171.065 ;
        RECT 110.475 170.755 112.085 170.965 ;
        RECT 112.385 170.875 112.585 171.665 ;
        RECT 110.475 170.155 110.750 170.755 ;
        RECT 112.255 170.705 112.585 170.875 ;
        RECT 112.755 170.715 113.075 171.895 ;
        RECT 113.705 170.730 113.995 171.895 ;
        RECT 114.165 170.805 116.755 171.895 ;
        RECT 116.930 171.460 122.275 171.895 ;
        RECT 112.255 170.585 112.435 170.705 ;
        RECT 110.920 170.335 111.275 170.585 ;
        RECT 111.470 170.535 111.935 170.585 ;
        RECT 111.465 170.365 111.935 170.535 ;
        RECT 111.470 170.335 111.935 170.365 ;
        RECT 112.105 170.335 112.435 170.585 ;
        RECT 112.610 170.335 113.075 170.535 ;
        RECT 114.165 170.285 115.375 170.805 ;
        RECT 110.475 169.975 111.725 170.155 ;
        RECT 111.360 169.905 111.725 169.975 ;
        RECT 111.895 169.955 113.075 170.125 ;
        RECT 115.545 170.115 116.755 170.635 ;
        RECT 118.520 170.210 118.870 171.460 ;
        RECT 122.635 171.170 122.965 171.895 ;
        RECT 110.535 169.345 110.705 169.805 ;
        RECT 111.895 169.735 112.225 169.955 ;
        RECT 110.975 169.555 112.225 169.735 ;
        RECT 112.395 169.345 112.565 169.785 ;
        RECT 112.735 169.540 113.075 169.955 ;
        RECT 113.705 169.345 113.995 170.070 ;
        RECT 114.165 169.345 116.755 170.115 ;
        RECT 120.350 169.890 120.690 170.720 ;
        RECT 116.930 169.345 122.275 169.890 ;
        RECT 122.445 169.515 122.965 171.000 ;
        RECT 123.135 170.175 123.655 171.725 ;
        RECT 123.915 170.965 124.085 171.725 ;
        RECT 124.300 171.135 124.630 171.895 ;
        RECT 123.915 170.795 124.630 170.965 ;
        RECT 124.800 170.820 125.055 171.725 ;
        RECT 123.825 170.245 124.180 170.615 ;
        RECT 124.460 170.585 124.630 170.795 ;
        RECT 124.460 170.255 124.715 170.585 ;
        RECT 124.460 170.065 124.630 170.255 ;
        RECT 124.885 170.090 125.055 170.820 ;
        RECT 125.230 170.745 125.490 171.895 ;
        RECT 125.665 170.805 126.875 171.895 ;
        RECT 125.665 170.265 126.185 170.805 ;
        RECT 123.135 169.345 123.475 170.005 ;
        RECT 123.915 169.895 124.630 170.065 ;
        RECT 123.915 169.515 124.085 169.895 ;
        RECT 124.300 169.345 124.630 169.725 ;
        RECT 124.800 169.515 125.055 170.090 ;
        RECT 125.230 169.345 125.490 170.185 ;
        RECT 126.355 170.095 126.875 170.635 ;
        RECT 125.665 169.345 126.875 170.095 ;
        RECT 14.260 169.175 126.960 169.345 ;
        RECT 128.405 74.775 134.895 74.945 ;
        RECT 50.705 70.245 110.465 70.695 ;
        RECT 50.705 70.115 110.525 70.245 ;
        RECT 50.485 69.875 110.525 70.115 ;
        RECT 50.485 69.630 52.195 69.875 ;
        RECT 58.775 69.645 60.485 69.875 ;
        RECT 46.190 69.460 50.000 69.630 ;
        RECT 46.190 63.650 46.360 69.460 ;
        RECT 46.840 66.820 47.530 68.980 ;
        RECT 46.840 64.130 47.530 66.290 ;
        RECT 48.010 63.650 48.180 69.460 ;
        RECT 48.660 66.820 49.350 68.980 ;
        RECT 48.660 64.130 49.350 66.290 ;
        RECT 49.830 63.650 50.000 69.460 ;
        RECT 46.190 63.480 50.000 63.650 ;
        RECT 1.470 57.840 13.600 58.010 ;
        RECT 1.470 56.190 1.640 57.840 ;
        RECT 2.120 56.670 4.280 57.360 ;
        RECT 4.810 56.670 6.970 57.360 ;
        RECT 7.450 56.190 7.620 57.840 ;
        RECT 8.100 56.670 10.260 57.360 ;
        RECT 10.790 56.670 12.950 57.360 ;
        RECT 13.430 56.190 13.600 57.840 ;
        RECT 46.190 57.670 46.360 63.480 ;
        RECT 46.840 60.840 47.530 63.000 ;
        RECT 46.840 58.150 47.530 60.310 ;
        RECT 48.010 57.670 48.180 63.480 ;
        RECT 48.660 60.840 49.350 63.000 ;
        RECT 48.660 58.150 49.350 60.310 ;
        RECT 49.830 57.670 50.000 63.480 ;
        RECT 50.480 69.460 52.230 69.630 ;
        RECT 50.480 61.970 50.650 69.460 ;
        RECT 51.190 68.950 51.520 69.120 ;
        RECT 51.050 62.695 51.220 68.735 ;
        RECT 51.490 62.695 51.660 68.735 ;
        RECT 51.190 62.310 51.520 62.480 ;
        RECT 52.060 61.970 52.230 69.460 ;
        RECT 50.480 61.800 52.230 61.970 ;
        RECT 52.655 69.475 58.285 69.645 ;
        RECT 52.655 63.665 52.825 69.475 ;
        RECT 53.305 66.835 53.995 68.995 ;
        RECT 53.305 64.145 53.995 66.305 ;
        RECT 54.475 63.665 54.645 69.475 ;
        RECT 55.125 66.835 55.815 68.995 ;
        RECT 55.125 64.145 55.815 66.305 ;
        RECT 56.295 63.665 56.465 69.475 ;
        RECT 56.945 66.835 57.635 68.995 ;
        RECT 56.945 64.145 57.635 66.305 ;
        RECT 58.115 63.665 58.285 69.475 ;
        RECT 52.655 63.495 58.285 63.665 ;
        RECT 50.460 61.075 52.210 61.245 ;
        RECT 50.460 57.675 50.630 61.075 ;
        RECT 51.170 60.565 51.500 60.735 ;
        RECT 51.030 58.355 51.200 60.395 ;
        RECT 51.470 58.355 51.640 60.395 ;
        RECT 51.170 58.015 51.500 58.185 ;
        RECT 52.040 57.675 52.210 61.075 ;
        RECT 50.460 57.670 52.210 57.675 ;
        RECT 52.655 57.685 52.825 63.495 ;
        RECT 53.305 60.855 53.995 63.015 ;
        RECT 53.305 58.165 53.995 60.325 ;
        RECT 54.475 57.685 54.645 63.495 ;
        RECT 55.125 60.855 55.815 63.015 ;
        RECT 55.125 58.165 55.815 60.325 ;
        RECT 56.295 57.685 56.465 63.495 ;
        RECT 56.945 60.855 57.635 63.015 ;
        RECT 56.945 58.165 57.635 60.325 ;
        RECT 58.115 57.685 58.285 63.495 ;
        RECT 58.775 69.475 60.525 69.645 ;
        RECT 58.775 61.985 58.945 69.475 ;
        RECT 59.485 68.965 59.815 69.135 ;
        RECT 59.345 62.710 59.515 68.750 ;
        RECT 59.785 62.710 59.955 68.750 ;
        RECT 59.485 62.325 59.815 62.495 ;
        RECT 60.355 61.985 60.525 69.475 ;
        RECT 58.775 61.815 60.525 61.985 ;
        RECT 60.985 69.465 66.615 69.635 ;
        RECT 60.985 63.655 61.155 69.465 ;
        RECT 61.635 66.825 62.325 68.985 ;
        RECT 61.635 64.135 62.325 66.295 ;
        RECT 62.805 63.655 62.975 69.465 ;
        RECT 63.455 66.825 64.145 68.985 ;
        RECT 63.455 64.135 64.145 66.295 ;
        RECT 64.625 63.655 64.795 69.465 ;
        RECT 65.275 66.825 65.965 68.985 ;
        RECT 65.275 64.135 65.965 66.295 ;
        RECT 66.445 63.655 66.615 69.465 ;
        RECT 66.915 69.485 69.035 69.875 ;
        RECT 75.425 69.675 77.325 69.875 ;
        RECT 66.915 69.405 69.015 69.485 ;
        RECT 69.280 69.455 74.910 69.625 ;
        RECT 60.985 63.485 66.615 63.655 ;
        RECT 52.655 57.670 58.285 57.685 ;
        RECT 58.765 61.075 60.515 61.245 ;
        RECT 58.765 57.675 58.935 61.075 ;
        RECT 59.475 60.565 59.805 60.735 ;
        RECT 59.335 58.355 59.505 60.395 ;
        RECT 59.775 58.355 59.945 60.395 ;
        RECT 59.475 58.015 59.805 58.185 ;
        RECT 60.345 57.675 60.515 61.075 ;
        RECT 58.765 57.670 60.515 57.675 ;
        RECT 60.985 57.675 61.155 63.485 ;
        RECT 61.635 60.845 62.325 63.005 ;
        RECT 61.635 58.155 62.325 60.315 ;
        RECT 62.805 57.675 62.975 63.485 ;
        RECT 63.455 60.845 64.145 63.005 ;
        RECT 63.455 58.155 64.145 60.315 ;
        RECT 64.625 57.675 64.795 63.485 ;
        RECT 65.275 60.845 65.965 63.005 ;
        RECT 65.275 58.155 65.965 60.315 ;
        RECT 66.445 57.675 66.615 63.485 ;
        RECT 67.090 61.975 67.260 69.405 ;
        RECT 67.800 68.955 68.130 69.125 ;
        RECT 67.660 62.700 67.830 68.740 ;
        RECT 68.100 62.700 68.270 68.740 ;
        RECT 67.800 62.315 68.130 62.485 ;
        RECT 68.670 61.975 68.840 69.405 ;
        RECT 67.090 61.805 68.840 61.975 ;
        RECT 69.280 63.645 69.450 69.455 ;
        RECT 69.930 66.815 70.620 68.975 ;
        RECT 69.930 64.125 70.620 66.285 ;
        RECT 71.100 63.645 71.270 69.455 ;
        RECT 71.750 66.815 72.440 68.975 ;
        RECT 71.750 64.125 72.440 66.285 ;
        RECT 72.920 63.645 73.090 69.455 ;
        RECT 73.570 66.815 74.260 68.975 ;
        RECT 73.570 64.125 74.260 66.285 ;
        RECT 74.740 63.645 74.910 69.455 ;
        RECT 69.280 63.475 74.910 63.645 ;
        RECT 60.985 57.670 66.615 57.675 ;
        RECT 67.025 61.075 68.775 61.245 ;
        RECT 67.025 57.675 67.195 61.075 ;
        RECT 67.735 60.565 68.065 60.735 ;
        RECT 67.595 58.355 67.765 60.395 ;
        RECT 68.035 58.355 68.205 60.395 ;
        RECT 67.735 58.015 68.065 58.185 ;
        RECT 68.605 57.675 68.775 61.075 ;
        RECT 67.025 57.670 68.775 57.675 ;
        RECT 69.280 57.670 69.450 63.475 ;
        RECT 69.930 60.835 70.620 62.995 ;
        RECT 69.930 58.145 70.620 60.305 ;
        RECT 71.100 57.670 71.270 63.475 ;
        RECT 71.750 60.835 72.440 62.995 ;
        RECT 71.750 58.145 72.440 60.305 ;
        RECT 72.920 57.670 73.090 63.475 ;
        RECT 73.570 60.835 74.260 62.995 ;
        RECT 73.570 58.145 74.260 60.305 ;
        RECT 74.740 57.670 74.910 63.475 ;
        RECT 75.470 69.565 77.220 69.675 ;
        RECT 83.865 69.660 85.575 69.875 ;
        RECT 92.195 69.685 93.905 69.875 ;
        RECT 100.485 69.700 102.195 69.875 ;
        RECT 75.470 62.075 75.640 69.565 ;
        RECT 76.180 69.055 76.510 69.225 ;
        RECT 76.040 62.800 76.210 68.840 ;
        RECT 76.480 62.800 76.650 68.840 ;
        RECT 76.180 62.415 76.510 62.585 ;
        RECT 77.050 62.075 77.220 69.565 ;
        RECT 75.470 61.905 77.220 62.075 ;
        RECT 77.725 69.470 83.355 69.640 ;
        RECT 77.725 63.660 77.895 69.470 ;
        RECT 78.375 66.830 79.065 68.990 ;
        RECT 78.375 64.140 79.065 66.300 ;
        RECT 79.545 63.660 79.715 69.470 ;
        RECT 80.195 66.830 80.885 68.990 ;
        RECT 80.195 64.140 80.885 66.300 ;
        RECT 81.365 63.660 81.535 69.470 ;
        RECT 82.015 66.830 82.705 68.990 ;
        RECT 82.015 64.140 82.705 66.300 ;
        RECT 83.185 63.660 83.355 69.470 ;
        RECT 77.725 63.490 83.355 63.660 ;
        RECT 75.445 61.095 77.195 61.265 ;
        RECT 75.445 57.695 75.615 61.095 ;
        RECT 76.155 60.585 76.485 60.755 ;
        RECT 76.015 58.375 76.185 60.415 ;
        RECT 76.455 58.375 76.625 60.415 ;
        RECT 76.155 58.035 76.485 58.205 ;
        RECT 77.025 57.695 77.195 61.095 ;
        RECT 75.445 57.670 77.195 57.695 ;
        RECT 77.725 57.680 77.895 63.490 ;
        RECT 78.375 60.850 79.065 63.010 ;
        RECT 78.375 58.160 79.065 60.320 ;
        RECT 79.545 57.680 79.715 63.490 ;
        RECT 80.195 60.850 80.885 63.010 ;
        RECT 80.195 58.160 80.885 60.320 ;
        RECT 81.365 57.680 81.535 63.490 ;
        RECT 82.015 60.850 82.705 63.010 ;
        RECT 82.015 58.160 82.705 60.320 ;
        RECT 83.185 57.680 83.355 63.490 ;
        RECT 83.860 69.490 85.610 69.660 ;
        RECT 83.860 62.000 84.030 69.490 ;
        RECT 84.570 68.980 84.900 69.150 ;
        RECT 84.430 62.725 84.600 68.765 ;
        RECT 84.870 62.725 85.040 68.765 ;
        RECT 84.570 62.340 84.900 62.510 ;
        RECT 85.440 62.000 85.610 69.490 ;
        RECT 83.860 61.830 85.610 62.000 ;
        RECT 86.055 69.470 91.685 69.640 ;
        RECT 86.055 63.660 86.225 69.470 ;
        RECT 86.705 66.830 87.395 68.990 ;
        RECT 86.705 64.140 87.395 66.300 ;
        RECT 87.875 63.660 88.045 69.470 ;
        RECT 88.525 66.830 89.215 68.990 ;
        RECT 88.525 64.140 89.215 66.300 ;
        RECT 89.695 63.660 89.865 69.470 ;
        RECT 90.345 66.830 91.035 68.990 ;
        RECT 90.345 64.140 91.035 66.300 ;
        RECT 91.515 63.660 91.685 69.470 ;
        RECT 86.055 63.490 91.685 63.660 ;
        RECT 77.725 57.670 83.355 57.680 ;
        RECT 83.795 61.075 85.545 61.245 ;
        RECT 83.795 57.675 83.965 61.075 ;
        RECT 84.505 60.565 84.835 60.735 ;
        RECT 84.365 58.355 84.535 60.395 ;
        RECT 84.805 58.355 84.975 60.395 ;
        RECT 84.505 58.015 84.835 58.185 ;
        RECT 85.375 57.675 85.545 61.075 ;
        RECT 83.795 57.670 85.545 57.675 ;
        RECT 86.055 57.680 86.225 63.490 ;
        RECT 86.705 60.850 87.395 63.010 ;
        RECT 86.705 58.160 87.395 60.320 ;
        RECT 87.875 57.680 88.045 63.490 ;
        RECT 88.525 60.850 89.215 63.010 ;
        RECT 88.525 58.160 89.215 60.320 ;
        RECT 89.695 57.680 89.865 63.490 ;
        RECT 90.345 60.850 91.035 63.010 ;
        RECT 90.345 58.160 91.035 60.320 ;
        RECT 91.515 57.680 91.685 63.490 ;
        RECT 92.190 69.515 93.940 69.685 ;
        RECT 92.190 62.025 92.360 69.515 ;
        RECT 92.900 69.005 93.230 69.175 ;
        RECT 92.760 62.750 92.930 68.790 ;
        RECT 93.200 62.750 93.370 68.790 ;
        RECT 92.900 62.365 93.230 62.535 ;
        RECT 93.770 62.025 93.940 69.515 ;
        RECT 92.190 61.855 93.940 62.025 ;
        RECT 94.385 69.470 100.015 69.640 ;
        RECT 94.385 63.660 94.555 69.470 ;
        RECT 95.035 66.830 95.725 68.990 ;
        RECT 95.035 64.140 95.725 66.300 ;
        RECT 96.205 63.660 96.375 69.470 ;
        RECT 96.855 66.830 97.545 68.990 ;
        RECT 96.855 64.140 97.545 66.300 ;
        RECT 98.025 63.660 98.195 69.470 ;
        RECT 98.675 66.830 99.365 68.990 ;
        RECT 98.675 64.140 99.365 66.300 ;
        RECT 99.845 63.660 100.015 69.470 ;
        RECT 94.385 63.490 100.015 63.660 ;
        RECT 86.055 57.670 91.685 57.680 ;
        RECT 92.180 61.070 93.930 61.240 ;
        RECT 92.180 57.670 92.350 61.070 ;
        RECT 92.890 60.560 93.220 60.730 ;
        RECT 92.750 58.350 92.920 60.390 ;
        RECT 93.190 58.350 93.360 60.390 ;
        RECT 92.890 58.010 93.220 58.180 ;
        RECT 93.760 57.670 93.930 61.070 ;
        RECT 94.385 57.680 94.555 63.490 ;
        RECT 95.035 60.850 95.725 63.010 ;
        RECT 95.035 58.160 95.725 60.320 ;
        RECT 96.205 57.680 96.375 63.490 ;
        RECT 96.855 60.850 97.545 63.010 ;
        RECT 96.855 58.160 97.545 60.320 ;
        RECT 98.025 57.680 98.195 63.490 ;
        RECT 98.675 60.850 99.365 63.010 ;
        RECT 98.675 58.160 99.365 60.320 ;
        RECT 99.845 57.680 100.015 63.490 ;
        RECT 100.485 69.530 102.235 69.700 ;
        RECT 108.815 69.680 110.525 69.875 ;
        RECT 100.485 62.040 100.655 69.530 ;
        RECT 101.195 69.020 101.525 69.190 ;
        RECT 101.055 62.765 101.225 68.805 ;
        RECT 101.495 62.765 101.665 68.805 ;
        RECT 101.195 62.380 101.525 62.550 ;
        RECT 102.065 62.040 102.235 69.530 ;
        RECT 100.485 61.870 102.235 62.040 ;
        RECT 102.690 69.465 108.320 69.635 ;
        RECT 102.690 63.655 102.860 69.465 ;
        RECT 103.340 66.825 104.030 68.985 ;
        RECT 103.340 64.135 104.030 66.295 ;
        RECT 104.510 63.655 104.680 69.465 ;
        RECT 105.160 66.825 105.850 68.985 ;
        RECT 105.160 64.135 105.850 66.295 ;
        RECT 106.330 63.655 106.500 69.465 ;
        RECT 106.980 66.825 107.670 68.985 ;
        RECT 106.980 64.135 107.670 66.295 ;
        RECT 108.150 63.655 108.320 69.465 ;
        RECT 102.690 63.485 108.320 63.655 ;
        RECT 94.385 57.670 100.015 57.680 ;
        RECT 100.420 61.080 102.170 61.250 ;
        RECT 100.420 57.680 100.590 61.080 ;
        RECT 101.130 60.570 101.460 60.740 ;
        RECT 100.990 58.360 101.160 60.400 ;
        RECT 101.430 58.360 101.600 60.400 ;
        RECT 101.130 58.020 101.460 58.190 ;
        RECT 102.000 57.680 102.170 61.080 ;
        RECT 100.420 57.670 102.170 57.680 ;
        RECT 102.690 57.675 102.860 63.485 ;
        RECT 103.340 60.845 104.030 63.005 ;
        RECT 103.340 58.155 104.030 60.315 ;
        RECT 104.510 57.675 104.680 63.485 ;
        RECT 105.160 60.845 105.850 63.005 ;
        RECT 105.160 58.155 105.850 60.315 ;
        RECT 106.330 57.675 106.500 63.485 ;
        RECT 106.980 60.845 107.670 63.005 ;
        RECT 106.980 58.155 107.670 60.315 ;
        RECT 108.150 57.675 108.320 63.485 ;
        RECT 108.785 69.510 110.535 69.680 ;
        RECT 108.785 62.020 108.955 69.510 ;
        RECT 109.495 69.000 109.825 69.170 ;
        RECT 109.355 62.745 109.525 68.785 ;
        RECT 109.795 62.745 109.965 68.785 ;
        RECT 109.495 62.360 109.825 62.530 ;
        RECT 110.365 62.020 110.535 69.510 ;
        RECT 108.785 61.850 110.535 62.020 ;
        RECT 110.990 69.475 114.800 69.645 ;
        RECT 110.990 63.665 111.160 69.475 ;
        RECT 111.640 66.835 112.330 68.995 ;
        RECT 111.640 64.145 112.330 66.305 ;
        RECT 112.810 63.665 112.980 69.475 ;
        RECT 113.460 66.835 114.150 68.995 ;
        RECT 113.460 64.145 114.150 66.305 ;
        RECT 114.630 63.665 114.800 69.475 ;
        RECT 128.405 66.785 128.575 74.775 ;
        RECT 129.115 74.265 129.445 74.435 ;
        RECT 126.540 66.345 128.575 66.785 ;
        RECT 126.350 65.790 128.575 66.345 ;
        RECT 126.350 65.740 126.600 65.790 ;
        RECT 110.990 63.495 114.800 63.665 ;
        RECT 102.690 57.670 108.320 57.675 ;
        RECT 108.785 61.080 110.535 61.250 ;
        RECT 108.785 57.680 108.955 61.080 ;
        RECT 109.495 60.570 109.825 60.740 ;
        RECT 109.355 58.360 109.525 60.400 ;
        RECT 109.795 58.360 109.965 60.400 ;
        RECT 109.495 58.020 109.825 58.190 ;
        RECT 110.365 57.680 110.535 61.080 ;
        RECT 108.785 57.670 110.535 57.680 ;
        RECT 110.990 57.685 111.160 63.495 ;
        RECT 111.640 60.855 112.330 63.015 ;
        RECT 111.640 58.165 112.330 60.325 ;
        RECT 112.810 57.685 112.980 63.495 ;
        RECT 113.460 60.855 114.150 63.015 ;
        RECT 113.460 58.165 114.150 60.325 ;
        RECT 114.630 57.685 114.800 63.495 ;
        RECT 126.370 63.365 126.540 65.740 ;
        RECT 127.080 65.345 127.410 65.515 ;
        RECT 126.940 64.090 127.110 65.130 ;
        RECT 127.380 64.090 127.550 65.130 ;
        RECT 127.080 63.705 127.410 63.875 ;
        RECT 127.950 63.365 128.575 65.790 ;
        RECT 128.975 64.010 129.145 74.050 ;
        RECT 129.415 64.010 129.585 74.050 ;
        RECT 129.115 63.625 129.445 63.795 ;
        RECT 126.370 63.285 128.575 63.365 ;
        RECT 129.985 63.285 130.155 74.775 ;
        RECT 130.695 74.265 131.025 74.435 ;
        RECT 130.555 64.010 130.725 74.050 ;
        RECT 130.995 64.010 131.165 74.050 ;
        RECT 130.695 63.625 131.025 63.795 ;
        RECT 131.565 63.285 131.735 74.775 ;
        RECT 132.275 74.265 132.605 74.435 ;
        RECT 132.135 64.010 132.305 74.050 ;
        RECT 132.575 64.010 132.745 74.050 ;
        RECT 132.275 63.625 132.605 63.795 ;
        RECT 133.145 63.285 133.315 74.775 ;
        RECT 133.855 74.265 134.185 74.435 ;
        RECT 133.715 64.010 133.885 74.050 ;
        RECT 134.155 64.010 134.325 74.050 ;
        RECT 133.855 63.625 134.185 63.795 ;
        RECT 134.725 63.285 134.895 74.775 ;
        RECT 126.370 63.195 134.895 63.285 ;
        RECT 127.980 63.120 134.895 63.195 ;
        RECT 128.405 63.115 134.895 63.120 ;
        RECT 126.370 62.675 128.120 62.715 ;
        RECT 128.405 62.675 134.895 62.720 ;
        RECT 126.370 62.550 134.895 62.675 ;
        RECT 126.370 62.545 128.575 62.550 ;
        RECT 126.370 60.145 126.540 62.545 ;
        RECT 127.080 62.035 127.410 62.205 ;
        RECT 126.940 60.825 127.110 61.865 ;
        RECT 127.380 60.825 127.550 61.865 ;
        RECT 127.080 60.485 127.410 60.655 ;
        RECT 127.950 60.145 128.575 62.545 ;
        RECT 129.115 62.040 129.445 62.210 ;
        RECT 126.370 59.975 128.575 60.145 ;
        RECT 126.415 59.790 128.575 59.975 ;
        RECT 126.490 59.655 128.575 59.790 ;
        RECT 126.550 59.415 128.575 59.655 ;
        RECT 110.990 57.670 114.800 57.685 ;
        RECT 46.190 56.795 114.805 57.670 ;
        RECT 128.405 57.150 128.575 59.415 ;
        RECT 128.975 57.830 129.145 61.870 ;
        RECT 129.415 57.830 129.585 61.870 ;
        RECT 129.115 57.490 129.445 57.660 ;
        RECT 129.985 57.150 130.155 62.550 ;
        RECT 130.695 62.040 131.025 62.210 ;
        RECT 130.555 57.830 130.725 61.870 ;
        RECT 130.995 57.830 131.165 61.870 ;
        RECT 130.695 57.490 131.025 57.660 ;
        RECT 131.565 57.150 131.735 62.550 ;
        RECT 132.275 62.040 132.605 62.210 ;
        RECT 132.135 57.830 132.305 61.870 ;
        RECT 132.575 57.830 132.745 61.870 ;
        RECT 132.275 57.490 132.605 57.660 ;
        RECT 133.145 57.150 133.315 62.550 ;
        RECT 133.855 62.040 134.185 62.210 ;
        RECT 133.715 57.830 133.885 61.870 ;
        RECT 134.155 57.830 134.325 61.870 ;
        RECT 133.855 57.490 134.185 57.660 ;
        RECT 134.725 57.150 134.895 62.550 ;
        RECT 128.405 56.980 134.895 57.150 ;
        RECT 1.470 56.020 13.600 56.190 ;
        RECT 1.470 54.370 1.640 56.020 ;
        RECT 2.120 54.850 4.280 55.540 ;
        RECT 4.810 54.850 6.970 55.540 ;
        RECT 7.450 54.370 7.620 56.020 ;
        RECT 8.100 54.850 10.260 55.540 ;
        RECT 10.790 54.850 12.950 55.540 ;
        RECT 13.430 54.370 13.600 56.020 ;
        RECT 1.470 54.200 13.600 54.370 ;
        RECT 1.470 52.550 1.640 54.200 ;
        RECT 2.120 53.030 4.280 53.720 ;
        RECT 4.810 53.030 6.970 53.720 ;
        RECT 7.450 52.550 7.620 54.200 ;
        RECT 8.100 53.030 10.260 53.720 ;
        RECT 10.790 53.030 12.950 53.720 ;
        RECT 13.430 52.550 13.600 54.200 ;
        RECT 1.470 52.380 31.540 52.550 ;
        RECT 1.470 50.855 1.640 52.380 ;
        RECT 2.120 51.210 4.280 51.900 ;
        RECT 4.810 51.210 6.970 51.900 ;
        RECT 7.450 50.855 7.620 52.380 ;
        RECT 8.100 51.210 10.260 51.900 ;
        RECT 10.790 51.210 12.950 51.900 ;
        RECT 1.470 50.730 9.960 50.855 ;
        RECT 13.430 50.730 13.600 52.380 ;
        RECT 14.080 51.210 16.240 51.900 ;
        RECT 16.770 51.210 18.930 51.900 ;
        RECT 19.410 50.730 19.580 52.380 ;
        RECT 20.060 51.210 22.220 51.900 ;
        RECT 22.750 51.210 24.910 51.900 ;
        RECT 25.390 50.730 25.560 52.380 ;
        RECT 26.040 51.210 28.200 51.900 ;
        RECT 28.730 51.210 30.890 51.900 ;
        RECT 31.370 50.730 31.540 52.380 ;
        RECT 1.470 50.560 31.540 50.730 ;
        RECT 43.490 52.540 61.600 52.550 ;
        RECT 67.490 52.540 85.600 52.550 ;
        RECT 43.490 52.380 85.600 52.540 ;
        RECT 43.490 50.730 43.660 52.380 ;
        RECT 44.140 51.210 46.300 51.900 ;
        RECT 46.830 51.210 48.990 51.900 ;
        RECT 49.470 50.730 49.640 52.380 ;
        RECT 50.120 51.210 52.280 51.900 ;
        RECT 52.810 51.210 54.970 51.900 ;
        RECT 55.450 50.730 55.620 52.380 ;
        RECT 61.430 52.090 67.670 52.380 ;
        RECT 56.100 51.210 58.260 51.900 ;
        RECT 58.790 51.210 60.950 51.900 ;
        RECT 61.430 50.730 61.600 52.090 ;
        RECT 43.490 50.560 61.600 50.730 ;
        RECT 67.490 50.730 67.660 52.090 ;
        RECT 68.140 51.210 70.300 51.900 ;
        RECT 70.830 51.210 72.990 51.900 ;
        RECT 73.470 50.730 73.640 52.380 ;
        RECT 74.120 51.210 76.280 51.900 ;
        RECT 76.810 51.210 78.970 51.900 ;
        RECT 79.450 50.730 79.620 52.380 ;
        RECT 80.100 51.210 82.260 51.900 ;
        RECT 82.790 51.210 84.950 51.900 ;
        RECT 85.430 50.730 85.600 52.380 ;
        RECT 67.490 50.560 85.600 50.730 ;
        RECT 1.585 50.360 9.960 50.560 ;
        RECT 77.790 50.170 80.360 50.560 ;
        RECT 1.450 49.480 27.925 49.960 ;
        RECT 29.450 49.480 55.925 49.960 ;
        RECT 57.450 49.480 83.925 49.960 ;
        RECT 85.450 49.480 111.925 49.960 ;
        RECT 113.450 49.480 139.925 49.960 ;
        RECT 1.435 49.420 27.925 49.480 ;
        RECT 29.435 49.420 55.925 49.480 ;
        RECT 57.435 49.420 83.925 49.480 ;
        RECT 85.435 49.420 111.925 49.480 ;
        RECT 113.435 49.420 139.925 49.480 ;
        RECT 143.470 49.840 149.620 50.010 ;
        RECT 1.435 49.260 27.980 49.420 ;
        RECT 1.435 49.235 14.180 49.260 ;
        RECT 1.435 49.005 5.760 49.235 ;
        RECT 1.470 39.745 1.640 49.005 ;
        RECT 2.365 48.435 4.405 48.605 ;
        RECT 1.980 40.375 2.150 48.375 ;
        RECT 4.620 40.375 4.790 48.375 ;
        RECT 2.365 40.145 4.405 40.315 ;
        RECT 5.130 39.745 5.300 49.005 ;
        RECT 1.470 39.575 5.300 39.745 ;
        RECT 5.590 39.745 5.760 49.005 ;
        RECT 6.390 48.725 8.390 48.895 ;
        RECT 6.160 40.470 6.330 48.510 ;
        RECT 8.450 40.470 8.620 48.510 ;
        RECT 6.390 40.085 8.390 40.255 ;
        RECT 9.020 39.745 9.190 49.235 ;
        RECT 9.820 48.725 11.820 48.895 ;
        RECT 9.590 40.470 9.760 48.510 ;
        RECT 11.880 40.470 12.050 48.510 ;
        RECT 12.450 47.665 14.180 49.235 ;
        RECT 26.230 49.250 27.980 49.260 ;
        RECT 12.450 47.495 20.915 47.665 ;
        RECT 12.450 46.085 14.255 47.495 ;
        RECT 14.595 46.625 14.765 46.955 ;
        RECT 14.980 46.925 20.020 47.095 ;
        RECT 14.980 46.485 20.020 46.655 ;
        RECT 20.235 46.625 20.405 46.955 ;
        RECT 20.745 46.085 20.915 47.495 ;
        RECT 12.450 45.915 20.915 46.085 ;
        RECT 12.450 45.400 14.180 45.915 ;
        RECT 12.450 45.285 23.930 45.400 ;
        RECT 9.820 40.085 11.820 40.255 ;
        RECT 12.450 39.745 12.620 45.285 ;
        RECT 5.590 39.575 12.620 39.745 ;
        RECT 12.900 45.230 23.930 45.285 ;
        RECT 12.900 39.740 13.070 45.230 ;
        RECT 13.700 44.720 17.700 44.890 ;
        RECT 13.470 40.465 13.640 44.505 ;
        RECT 17.760 40.465 17.930 44.505 ;
        RECT 13.700 40.080 17.700 40.250 ;
        RECT 18.330 39.740 18.500 45.230 ;
        RECT 19.130 44.720 23.130 44.890 ;
        RECT 18.900 40.465 19.070 44.505 ;
        RECT 23.190 40.465 23.360 44.505 ;
        RECT 19.130 40.080 23.130 40.250 ;
        RECT 23.760 39.740 23.930 45.230 ;
        RECT 12.900 39.570 23.930 39.740 ;
        RECT 24.205 45.245 25.955 45.415 ;
        RECT 24.205 39.755 24.375 45.245 ;
        RECT 24.915 44.735 25.245 44.905 ;
        RECT 24.775 40.480 24.945 44.520 ;
        RECT 25.215 40.480 25.385 44.520 ;
        RECT 24.915 40.095 25.245 40.265 ;
        RECT 25.785 39.755 25.955 45.245 ;
        RECT 24.205 39.585 25.955 39.755 ;
        RECT 26.230 39.760 26.400 49.250 ;
        RECT 26.940 48.740 27.270 48.910 ;
        RECT 26.800 40.485 26.970 48.525 ;
        RECT 27.240 40.485 27.410 48.525 ;
        RECT 26.940 40.100 27.270 40.270 ;
        RECT 27.810 39.760 27.980 49.250 ;
        RECT 29.435 49.260 55.980 49.420 ;
        RECT 29.435 49.235 42.180 49.260 ;
        RECT 29.435 49.005 33.760 49.235 ;
        RECT 26.230 39.590 27.980 39.760 ;
        RECT 29.470 39.745 29.640 49.005 ;
        RECT 30.365 48.435 32.405 48.605 ;
        RECT 29.980 40.375 30.150 48.375 ;
        RECT 32.620 40.375 32.790 48.375 ;
        RECT 30.365 40.145 32.405 40.315 ;
        RECT 33.130 39.745 33.300 49.005 ;
        RECT 29.470 39.575 33.300 39.745 ;
        RECT 33.590 39.745 33.760 49.005 ;
        RECT 34.390 48.725 36.390 48.895 ;
        RECT 34.160 40.470 34.330 48.510 ;
        RECT 36.450 40.470 36.620 48.510 ;
        RECT 34.390 40.085 36.390 40.255 ;
        RECT 37.020 39.745 37.190 49.235 ;
        RECT 37.820 48.725 39.820 48.895 ;
        RECT 37.590 40.470 37.760 48.510 ;
        RECT 39.880 40.470 40.050 48.510 ;
        RECT 40.450 47.665 42.180 49.235 ;
        RECT 54.230 49.250 55.980 49.260 ;
        RECT 40.450 47.495 48.915 47.665 ;
        RECT 40.450 46.085 42.255 47.495 ;
        RECT 42.595 46.625 42.765 46.955 ;
        RECT 42.980 46.925 48.020 47.095 ;
        RECT 42.980 46.485 48.020 46.655 ;
        RECT 48.235 46.625 48.405 46.955 ;
        RECT 48.745 46.085 48.915 47.495 ;
        RECT 40.450 45.915 48.915 46.085 ;
        RECT 40.450 45.400 42.180 45.915 ;
        RECT 40.450 45.285 51.930 45.400 ;
        RECT 37.820 40.085 39.820 40.255 ;
        RECT 40.450 39.745 40.620 45.285 ;
        RECT 33.590 39.575 40.620 39.745 ;
        RECT 40.900 45.230 51.930 45.285 ;
        RECT 40.900 39.740 41.070 45.230 ;
        RECT 41.700 44.720 45.700 44.890 ;
        RECT 41.470 40.465 41.640 44.505 ;
        RECT 45.760 40.465 45.930 44.505 ;
        RECT 41.700 40.080 45.700 40.250 ;
        RECT 46.330 39.740 46.500 45.230 ;
        RECT 47.130 44.720 51.130 44.890 ;
        RECT 46.900 40.465 47.070 44.505 ;
        RECT 51.190 40.465 51.360 44.505 ;
        RECT 47.130 40.080 51.130 40.250 ;
        RECT 51.760 39.740 51.930 45.230 ;
        RECT 40.900 39.570 51.930 39.740 ;
        RECT 52.205 45.245 53.955 45.415 ;
        RECT 52.205 39.755 52.375 45.245 ;
        RECT 52.915 44.735 53.245 44.905 ;
        RECT 52.775 40.480 52.945 44.520 ;
        RECT 53.215 40.480 53.385 44.520 ;
        RECT 52.915 40.095 53.245 40.265 ;
        RECT 53.785 39.755 53.955 45.245 ;
        RECT 52.205 39.585 53.955 39.755 ;
        RECT 54.230 39.760 54.400 49.250 ;
        RECT 54.940 48.740 55.270 48.910 ;
        RECT 54.800 40.485 54.970 48.525 ;
        RECT 55.240 40.485 55.410 48.525 ;
        RECT 54.940 40.100 55.270 40.270 ;
        RECT 55.810 39.760 55.980 49.250 ;
        RECT 57.435 49.260 83.980 49.420 ;
        RECT 57.435 49.235 70.180 49.260 ;
        RECT 57.435 49.005 61.760 49.235 ;
        RECT 54.230 39.590 55.980 39.760 ;
        RECT 57.470 39.745 57.640 49.005 ;
        RECT 58.365 48.435 60.405 48.605 ;
        RECT 57.980 40.375 58.150 48.375 ;
        RECT 60.620 40.375 60.790 48.375 ;
        RECT 58.365 40.145 60.405 40.315 ;
        RECT 61.130 39.745 61.300 49.005 ;
        RECT 57.470 39.575 61.300 39.745 ;
        RECT 61.590 39.745 61.760 49.005 ;
        RECT 62.390 48.725 64.390 48.895 ;
        RECT 62.160 40.470 62.330 48.510 ;
        RECT 64.450 40.470 64.620 48.510 ;
        RECT 62.390 40.085 64.390 40.255 ;
        RECT 65.020 39.745 65.190 49.235 ;
        RECT 65.820 48.725 67.820 48.895 ;
        RECT 65.590 40.470 65.760 48.510 ;
        RECT 67.880 40.470 68.050 48.510 ;
        RECT 68.450 47.665 70.180 49.235 ;
        RECT 82.230 49.250 83.980 49.260 ;
        RECT 68.450 47.495 76.915 47.665 ;
        RECT 68.450 46.085 70.255 47.495 ;
        RECT 70.595 46.625 70.765 46.955 ;
        RECT 70.980 46.925 76.020 47.095 ;
        RECT 70.980 46.485 76.020 46.655 ;
        RECT 76.235 46.625 76.405 46.955 ;
        RECT 76.745 46.085 76.915 47.495 ;
        RECT 68.450 45.915 76.915 46.085 ;
        RECT 68.450 45.400 70.180 45.915 ;
        RECT 68.450 45.285 79.930 45.400 ;
        RECT 65.820 40.085 67.820 40.255 ;
        RECT 68.450 39.745 68.620 45.285 ;
        RECT 61.590 39.575 68.620 39.745 ;
        RECT 68.900 45.230 79.930 45.285 ;
        RECT 68.900 39.740 69.070 45.230 ;
        RECT 69.700 44.720 73.700 44.890 ;
        RECT 69.470 40.465 69.640 44.505 ;
        RECT 73.760 40.465 73.930 44.505 ;
        RECT 69.700 40.080 73.700 40.250 ;
        RECT 74.330 39.740 74.500 45.230 ;
        RECT 75.130 44.720 79.130 44.890 ;
        RECT 74.900 40.465 75.070 44.505 ;
        RECT 79.190 40.465 79.360 44.505 ;
        RECT 75.130 40.080 79.130 40.250 ;
        RECT 79.760 39.740 79.930 45.230 ;
        RECT 68.900 39.570 79.930 39.740 ;
        RECT 80.205 45.245 81.955 45.415 ;
        RECT 80.205 39.755 80.375 45.245 ;
        RECT 80.915 44.735 81.245 44.905 ;
        RECT 80.775 40.480 80.945 44.520 ;
        RECT 81.215 40.480 81.385 44.520 ;
        RECT 80.915 40.095 81.245 40.265 ;
        RECT 81.785 39.755 81.955 45.245 ;
        RECT 80.205 39.585 81.955 39.755 ;
        RECT 82.230 39.760 82.400 49.250 ;
        RECT 82.940 48.740 83.270 48.910 ;
        RECT 82.800 40.485 82.970 48.525 ;
        RECT 83.240 40.485 83.410 48.525 ;
        RECT 82.940 40.100 83.270 40.270 ;
        RECT 83.810 39.760 83.980 49.250 ;
        RECT 85.435 49.260 111.980 49.420 ;
        RECT 85.435 49.235 98.180 49.260 ;
        RECT 85.435 49.005 89.760 49.235 ;
        RECT 82.230 39.590 83.980 39.760 ;
        RECT 85.470 39.745 85.640 49.005 ;
        RECT 86.365 48.435 88.405 48.605 ;
        RECT 85.980 40.375 86.150 48.375 ;
        RECT 88.620 40.375 88.790 48.375 ;
        RECT 86.365 40.145 88.405 40.315 ;
        RECT 89.130 39.745 89.300 49.005 ;
        RECT 85.470 39.575 89.300 39.745 ;
        RECT 89.590 39.745 89.760 49.005 ;
        RECT 90.390 48.725 92.390 48.895 ;
        RECT 90.160 40.470 90.330 48.510 ;
        RECT 92.450 40.470 92.620 48.510 ;
        RECT 90.390 40.085 92.390 40.255 ;
        RECT 93.020 39.745 93.190 49.235 ;
        RECT 93.820 48.725 95.820 48.895 ;
        RECT 93.590 40.470 93.760 48.510 ;
        RECT 95.880 40.470 96.050 48.510 ;
        RECT 96.450 47.665 98.180 49.235 ;
        RECT 110.230 49.250 111.980 49.260 ;
        RECT 96.450 47.495 104.915 47.665 ;
        RECT 96.450 46.085 98.255 47.495 ;
        RECT 98.595 46.625 98.765 46.955 ;
        RECT 98.980 46.925 104.020 47.095 ;
        RECT 98.980 46.485 104.020 46.655 ;
        RECT 104.235 46.625 104.405 46.955 ;
        RECT 104.745 46.085 104.915 47.495 ;
        RECT 96.450 45.915 104.915 46.085 ;
        RECT 96.450 45.400 98.180 45.915 ;
        RECT 96.450 45.285 107.930 45.400 ;
        RECT 93.820 40.085 95.820 40.255 ;
        RECT 96.450 39.745 96.620 45.285 ;
        RECT 89.590 39.575 96.620 39.745 ;
        RECT 96.900 45.230 107.930 45.285 ;
        RECT 96.900 39.740 97.070 45.230 ;
        RECT 97.700 44.720 101.700 44.890 ;
        RECT 97.470 40.465 97.640 44.505 ;
        RECT 101.760 40.465 101.930 44.505 ;
        RECT 97.700 40.080 101.700 40.250 ;
        RECT 102.330 39.740 102.500 45.230 ;
        RECT 103.130 44.720 107.130 44.890 ;
        RECT 102.900 40.465 103.070 44.505 ;
        RECT 107.190 40.465 107.360 44.505 ;
        RECT 103.130 40.080 107.130 40.250 ;
        RECT 107.760 39.740 107.930 45.230 ;
        RECT 96.900 39.570 107.930 39.740 ;
        RECT 108.205 45.245 109.955 45.415 ;
        RECT 108.205 39.755 108.375 45.245 ;
        RECT 108.915 44.735 109.245 44.905 ;
        RECT 108.775 40.480 108.945 44.520 ;
        RECT 109.215 40.480 109.385 44.520 ;
        RECT 108.915 40.095 109.245 40.265 ;
        RECT 109.785 39.755 109.955 45.245 ;
        RECT 108.205 39.585 109.955 39.755 ;
        RECT 110.230 39.760 110.400 49.250 ;
        RECT 110.940 48.740 111.270 48.910 ;
        RECT 110.800 40.485 110.970 48.525 ;
        RECT 111.240 40.485 111.410 48.525 ;
        RECT 110.940 40.100 111.270 40.270 ;
        RECT 111.810 39.760 111.980 49.250 ;
        RECT 113.435 49.260 139.980 49.420 ;
        RECT 113.435 49.235 126.180 49.260 ;
        RECT 113.435 49.005 117.760 49.235 ;
        RECT 110.230 39.590 111.980 39.760 ;
        RECT 113.470 39.745 113.640 49.005 ;
        RECT 114.365 48.435 116.405 48.605 ;
        RECT 113.980 40.375 114.150 48.375 ;
        RECT 116.620 40.375 116.790 48.375 ;
        RECT 114.365 40.145 116.405 40.315 ;
        RECT 117.130 39.745 117.300 49.005 ;
        RECT 113.470 39.575 117.300 39.745 ;
        RECT 117.590 39.745 117.760 49.005 ;
        RECT 118.390 48.725 120.390 48.895 ;
        RECT 118.160 40.470 118.330 48.510 ;
        RECT 120.450 40.470 120.620 48.510 ;
        RECT 118.390 40.085 120.390 40.255 ;
        RECT 121.020 39.745 121.190 49.235 ;
        RECT 121.820 48.725 123.820 48.895 ;
        RECT 121.590 40.470 121.760 48.510 ;
        RECT 123.880 40.470 124.050 48.510 ;
        RECT 124.450 47.665 126.180 49.235 ;
        RECT 138.230 49.250 139.980 49.260 ;
        RECT 124.450 47.495 132.915 47.665 ;
        RECT 124.450 46.085 126.255 47.495 ;
        RECT 126.595 46.625 126.765 46.955 ;
        RECT 126.980 46.925 132.020 47.095 ;
        RECT 126.980 46.485 132.020 46.655 ;
        RECT 132.235 46.625 132.405 46.955 ;
        RECT 132.745 46.085 132.915 47.495 ;
        RECT 124.450 45.915 132.915 46.085 ;
        RECT 124.450 45.400 126.180 45.915 ;
        RECT 124.450 45.285 135.930 45.400 ;
        RECT 121.820 40.085 123.820 40.255 ;
        RECT 124.450 39.745 124.620 45.285 ;
        RECT 117.590 39.575 124.620 39.745 ;
        RECT 124.900 45.230 135.930 45.285 ;
        RECT 124.900 39.740 125.070 45.230 ;
        RECT 125.700 44.720 129.700 44.890 ;
        RECT 125.470 40.465 125.640 44.505 ;
        RECT 129.760 40.465 129.930 44.505 ;
        RECT 125.700 40.080 129.700 40.250 ;
        RECT 130.330 39.740 130.500 45.230 ;
        RECT 131.130 44.720 135.130 44.890 ;
        RECT 130.900 40.465 131.070 44.505 ;
        RECT 135.190 40.465 135.360 44.505 ;
        RECT 131.130 40.080 135.130 40.250 ;
        RECT 135.760 39.740 135.930 45.230 ;
        RECT 124.900 39.570 135.930 39.740 ;
        RECT 136.205 45.245 137.955 45.415 ;
        RECT 136.205 39.755 136.375 45.245 ;
        RECT 136.915 44.735 137.245 44.905 ;
        RECT 136.775 40.480 136.945 44.520 ;
        RECT 137.215 40.480 137.385 44.520 ;
        RECT 136.915 40.095 137.245 40.265 ;
        RECT 137.785 39.755 137.955 45.245 ;
        RECT 136.205 39.585 137.955 39.755 ;
        RECT 138.230 39.760 138.400 49.250 ;
        RECT 138.940 48.740 139.270 48.910 ;
        RECT 138.800 40.485 138.970 48.525 ;
        RECT 139.240 40.485 139.410 48.525 ;
        RECT 138.940 40.100 139.270 40.270 ;
        RECT 139.810 39.760 139.980 49.250 ;
        RECT 143.470 48.190 143.640 49.840 ;
        RECT 144.120 48.670 146.280 49.360 ;
        RECT 146.810 48.670 148.970 49.360 ;
        RECT 149.450 48.190 149.620 49.840 ;
        RECT 143.470 48.020 149.620 48.190 ;
        RECT 143.470 46.370 143.640 48.020 ;
        RECT 144.120 46.850 146.280 47.540 ;
        RECT 146.810 46.850 148.970 47.540 ;
        RECT 149.450 46.370 149.620 48.020 ;
        RECT 143.470 46.200 149.620 46.370 ;
        RECT 143.470 44.550 143.640 46.200 ;
        RECT 144.120 45.030 146.280 45.720 ;
        RECT 146.810 45.030 148.970 45.720 ;
        RECT 149.450 44.550 149.620 46.200 ;
        RECT 143.470 44.380 155.600 44.550 ;
        RECT 143.470 42.730 143.640 44.380 ;
        RECT 144.120 43.210 146.280 43.900 ;
        RECT 146.810 43.210 148.970 43.900 ;
        RECT 149.450 42.730 149.620 44.380 ;
        RECT 150.100 43.210 152.260 43.900 ;
        RECT 152.790 43.210 154.950 43.900 ;
        RECT 155.430 42.730 155.600 44.380 ;
        RECT 143.470 42.560 155.600 42.730 ;
        RECT 143.470 40.910 143.640 42.560 ;
        RECT 144.120 41.390 146.280 42.080 ;
        RECT 146.810 41.390 148.970 42.080 ;
        RECT 149.450 40.910 149.620 42.560 ;
        RECT 150.100 41.390 152.260 42.080 ;
        RECT 152.790 41.390 154.950 42.080 ;
        RECT 155.430 40.910 155.600 42.560 ;
        RECT 143.470 40.740 155.600 40.910 ;
        RECT 150.780 40.250 154.340 40.740 ;
        RECT 138.230 39.590 139.980 39.760 ;
        RECT 2.130 38.665 24.020 38.835 ;
        RECT 2.130 35.265 2.300 38.665 ;
        RECT 2.930 38.155 6.930 38.325 ;
        RECT 2.700 35.945 2.870 37.985 ;
        RECT 6.990 35.945 7.160 37.985 ;
        RECT 2.930 35.605 6.930 35.775 ;
        RECT 7.560 35.265 7.730 38.665 ;
        RECT 8.360 38.155 12.360 38.325 ;
        RECT 8.130 35.945 8.300 37.985 ;
        RECT 12.420 35.945 12.590 37.985 ;
        RECT 8.360 35.605 12.360 35.775 ;
        RECT 12.990 35.265 13.160 38.665 ;
        RECT 13.790 38.155 17.790 38.325 ;
        RECT 13.560 35.945 13.730 37.985 ;
        RECT 17.850 35.945 18.020 37.985 ;
        RECT 13.790 35.605 17.790 35.775 ;
        RECT 18.420 35.265 18.590 38.665 ;
        RECT 19.220 38.155 23.220 38.325 ;
        RECT 18.990 35.945 19.160 37.985 ;
        RECT 23.280 35.945 23.450 37.985 ;
        RECT 23.850 36.240 24.020 38.665 ;
        RECT 24.290 38.670 26.040 38.840 ;
        RECT 24.290 36.270 24.460 38.670 ;
        RECT 25.000 38.160 25.330 38.330 ;
        RECT 24.860 36.950 25.030 37.990 ;
        RECT 25.300 36.950 25.470 37.990 ;
        RECT 25.000 36.610 25.330 36.780 ;
        RECT 25.870 36.270 26.040 38.670 ;
        RECT 24.290 36.240 26.040 36.270 ;
        RECT 26.315 38.675 28.065 38.845 ;
        RECT 26.315 36.240 26.485 38.675 ;
        RECT 27.025 38.165 27.355 38.335 ;
        RECT 19.220 35.605 23.220 35.775 ;
        RECT 23.850 35.275 26.485 36.240 ;
        RECT 26.885 35.955 27.055 37.995 ;
        RECT 27.325 35.955 27.495 37.995 ;
        RECT 27.025 35.615 27.355 35.785 ;
        RECT 27.895 35.275 28.065 38.675 ;
        RECT 23.850 35.265 28.065 35.275 ;
        RECT 2.130 35.245 28.065 35.265 ;
        RECT 30.130 38.665 52.020 38.835 ;
        RECT 30.130 35.265 30.300 38.665 ;
        RECT 30.930 38.155 34.930 38.325 ;
        RECT 30.700 35.945 30.870 37.985 ;
        RECT 34.990 35.945 35.160 37.985 ;
        RECT 30.930 35.605 34.930 35.775 ;
        RECT 35.560 35.265 35.730 38.665 ;
        RECT 36.360 38.155 40.360 38.325 ;
        RECT 36.130 35.945 36.300 37.985 ;
        RECT 40.420 35.945 40.590 37.985 ;
        RECT 36.360 35.605 40.360 35.775 ;
        RECT 40.990 35.265 41.160 38.665 ;
        RECT 41.790 38.155 45.790 38.325 ;
        RECT 41.560 35.945 41.730 37.985 ;
        RECT 45.850 35.945 46.020 37.985 ;
        RECT 41.790 35.605 45.790 35.775 ;
        RECT 46.420 35.265 46.590 38.665 ;
        RECT 47.220 38.155 51.220 38.325 ;
        RECT 46.990 35.945 47.160 37.985 ;
        RECT 51.280 35.945 51.450 37.985 ;
        RECT 51.850 36.240 52.020 38.665 ;
        RECT 52.290 38.670 54.040 38.840 ;
        RECT 52.290 36.270 52.460 38.670 ;
        RECT 53.000 38.160 53.330 38.330 ;
        RECT 52.860 36.950 53.030 37.990 ;
        RECT 53.300 36.950 53.470 37.990 ;
        RECT 53.000 36.610 53.330 36.780 ;
        RECT 53.870 36.270 54.040 38.670 ;
        RECT 52.290 36.240 54.040 36.270 ;
        RECT 54.315 38.675 56.065 38.845 ;
        RECT 54.315 36.240 54.485 38.675 ;
        RECT 55.025 38.165 55.355 38.335 ;
        RECT 47.220 35.605 51.220 35.775 ;
        RECT 51.850 35.275 54.485 36.240 ;
        RECT 54.885 35.955 55.055 37.995 ;
        RECT 55.325 35.955 55.495 37.995 ;
        RECT 55.025 35.615 55.355 35.785 ;
        RECT 55.895 35.275 56.065 38.675 ;
        RECT 51.850 35.265 56.065 35.275 ;
        RECT 30.130 35.245 56.065 35.265 ;
        RECT 58.130 38.665 80.020 38.835 ;
        RECT 58.130 35.265 58.300 38.665 ;
        RECT 58.930 38.155 62.930 38.325 ;
        RECT 58.700 35.945 58.870 37.985 ;
        RECT 62.990 35.945 63.160 37.985 ;
        RECT 58.930 35.605 62.930 35.775 ;
        RECT 63.560 35.265 63.730 38.665 ;
        RECT 64.360 38.155 68.360 38.325 ;
        RECT 64.130 35.945 64.300 37.985 ;
        RECT 68.420 35.945 68.590 37.985 ;
        RECT 64.360 35.605 68.360 35.775 ;
        RECT 68.990 35.265 69.160 38.665 ;
        RECT 69.790 38.155 73.790 38.325 ;
        RECT 69.560 35.945 69.730 37.985 ;
        RECT 73.850 35.945 74.020 37.985 ;
        RECT 69.790 35.605 73.790 35.775 ;
        RECT 74.420 35.265 74.590 38.665 ;
        RECT 75.220 38.155 79.220 38.325 ;
        RECT 74.990 35.945 75.160 37.985 ;
        RECT 79.280 35.945 79.450 37.985 ;
        RECT 79.850 36.240 80.020 38.665 ;
        RECT 80.290 38.670 82.040 38.840 ;
        RECT 80.290 36.270 80.460 38.670 ;
        RECT 81.000 38.160 81.330 38.330 ;
        RECT 80.860 36.950 81.030 37.990 ;
        RECT 81.300 36.950 81.470 37.990 ;
        RECT 81.000 36.610 81.330 36.780 ;
        RECT 81.870 36.270 82.040 38.670 ;
        RECT 80.290 36.240 82.040 36.270 ;
        RECT 82.315 38.675 84.065 38.845 ;
        RECT 82.315 36.240 82.485 38.675 ;
        RECT 83.025 38.165 83.355 38.335 ;
        RECT 75.220 35.605 79.220 35.775 ;
        RECT 79.850 35.275 82.485 36.240 ;
        RECT 82.885 35.955 83.055 37.995 ;
        RECT 83.325 35.955 83.495 37.995 ;
        RECT 83.025 35.615 83.355 35.785 ;
        RECT 83.895 35.275 84.065 38.675 ;
        RECT 79.850 35.265 84.065 35.275 ;
        RECT 58.130 35.245 84.065 35.265 ;
        RECT 86.130 38.665 108.020 38.835 ;
        RECT 86.130 35.265 86.300 38.665 ;
        RECT 86.930 38.155 90.930 38.325 ;
        RECT 86.700 35.945 86.870 37.985 ;
        RECT 90.990 35.945 91.160 37.985 ;
        RECT 86.930 35.605 90.930 35.775 ;
        RECT 91.560 35.265 91.730 38.665 ;
        RECT 92.360 38.155 96.360 38.325 ;
        RECT 92.130 35.945 92.300 37.985 ;
        RECT 96.420 35.945 96.590 37.985 ;
        RECT 92.360 35.605 96.360 35.775 ;
        RECT 96.990 35.265 97.160 38.665 ;
        RECT 97.790 38.155 101.790 38.325 ;
        RECT 97.560 35.945 97.730 37.985 ;
        RECT 101.850 35.945 102.020 37.985 ;
        RECT 97.790 35.605 101.790 35.775 ;
        RECT 102.420 35.265 102.590 38.665 ;
        RECT 103.220 38.155 107.220 38.325 ;
        RECT 102.990 35.945 103.160 37.985 ;
        RECT 107.280 35.945 107.450 37.985 ;
        RECT 107.850 36.240 108.020 38.665 ;
        RECT 108.290 38.670 110.040 38.840 ;
        RECT 108.290 36.270 108.460 38.670 ;
        RECT 109.000 38.160 109.330 38.330 ;
        RECT 108.860 36.950 109.030 37.990 ;
        RECT 109.300 36.950 109.470 37.990 ;
        RECT 109.000 36.610 109.330 36.780 ;
        RECT 109.870 36.270 110.040 38.670 ;
        RECT 108.290 36.240 110.040 36.270 ;
        RECT 110.315 38.675 112.065 38.845 ;
        RECT 110.315 36.240 110.485 38.675 ;
        RECT 111.025 38.165 111.355 38.335 ;
        RECT 103.220 35.605 107.220 35.775 ;
        RECT 107.850 35.275 110.485 36.240 ;
        RECT 110.885 35.955 111.055 37.995 ;
        RECT 111.325 35.955 111.495 37.995 ;
        RECT 111.025 35.615 111.355 35.785 ;
        RECT 111.895 35.275 112.065 38.675 ;
        RECT 107.850 35.265 112.065 35.275 ;
        RECT 86.130 35.245 112.065 35.265 ;
        RECT 114.130 38.665 136.020 38.835 ;
        RECT 114.130 35.265 114.300 38.665 ;
        RECT 114.930 38.155 118.930 38.325 ;
        RECT 114.700 35.945 114.870 37.985 ;
        RECT 118.990 35.945 119.160 37.985 ;
        RECT 114.930 35.605 118.930 35.775 ;
        RECT 119.560 35.265 119.730 38.665 ;
        RECT 120.360 38.155 124.360 38.325 ;
        RECT 120.130 35.945 120.300 37.985 ;
        RECT 124.420 35.945 124.590 37.985 ;
        RECT 120.360 35.605 124.360 35.775 ;
        RECT 124.990 35.265 125.160 38.665 ;
        RECT 125.790 38.155 129.790 38.325 ;
        RECT 125.560 35.945 125.730 37.985 ;
        RECT 129.850 35.945 130.020 37.985 ;
        RECT 125.790 35.605 129.790 35.775 ;
        RECT 130.420 35.265 130.590 38.665 ;
        RECT 131.220 38.155 135.220 38.325 ;
        RECT 130.990 35.945 131.160 37.985 ;
        RECT 135.280 35.945 135.450 37.985 ;
        RECT 135.850 36.240 136.020 38.665 ;
        RECT 136.290 38.670 138.040 38.840 ;
        RECT 136.290 36.270 136.460 38.670 ;
        RECT 137.000 38.160 137.330 38.330 ;
        RECT 136.860 36.950 137.030 37.990 ;
        RECT 137.300 36.950 137.470 37.990 ;
        RECT 137.000 36.610 137.330 36.780 ;
        RECT 137.870 36.270 138.040 38.670 ;
        RECT 136.290 36.240 138.040 36.270 ;
        RECT 138.315 38.675 140.065 38.845 ;
        RECT 138.315 36.240 138.485 38.675 ;
        RECT 139.025 38.165 139.355 38.335 ;
        RECT 131.220 35.605 135.220 35.775 ;
        RECT 135.850 35.275 138.485 36.240 ;
        RECT 138.885 35.955 139.055 37.995 ;
        RECT 139.325 35.955 139.495 37.995 ;
        RECT 139.025 35.615 139.355 35.785 ;
        RECT 139.895 35.275 140.065 38.675 ;
        RECT 135.850 35.265 140.065 35.275 ;
        RECT 114.130 35.245 140.065 35.265 ;
        RECT 1.475 35.105 28.065 35.245 ;
        RECT 29.475 35.105 56.065 35.245 ;
        RECT 57.475 35.105 84.065 35.245 ;
        RECT 85.475 35.105 112.065 35.245 ;
        RECT 113.475 35.105 140.065 35.245 ;
        RECT 1.475 34.380 28.055 35.105 ;
        RECT 29.475 34.380 56.055 35.105 ;
        RECT 57.475 34.380 84.055 35.105 ;
        RECT 85.475 34.380 112.055 35.105 ;
        RECT 113.475 34.380 140.055 35.105 ;
        RECT 1.450 33.480 27.925 33.960 ;
        RECT 29.450 33.480 55.925 33.960 ;
        RECT 57.450 33.480 83.925 33.960 ;
        RECT 85.450 33.480 111.925 33.960 ;
        RECT 113.450 33.480 139.925 33.960 ;
        RECT 1.435 33.420 27.925 33.480 ;
        RECT 29.435 33.420 55.925 33.480 ;
        RECT 57.435 33.420 83.925 33.480 ;
        RECT 85.435 33.420 111.925 33.480 ;
        RECT 113.435 33.420 139.925 33.480 ;
        RECT 1.435 33.260 27.980 33.420 ;
        RECT 1.435 33.235 14.180 33.260 ;
        RECT 1.435 33.005 5.760 33.235 ;
        RECT 1.470 23.745 1.640 33.005 ;
        RECT 2.365 32.435 4.405 32.605 ;
        RECT 1.980 24.375 2.150 32.375 ;
        RECT 4.620 24.375 4.790 32.375 ;
        RECT 2.365 24.145 4.405 24.315 ;
        RECT 5.130 23.745 5.300 33.005 ;
        RECT 1.470 23.575 5.300 23.745 ;
        RECT 5.590 23.745 5.760 33.005 ;
        RECT 6.390 32.725 8.390 32.895 ;
        RECT 6.160 24.470 6.330 32.510 ;
        RECT 8.450 24.470 8.620 32.510 ;
        RECT 6.390 24.085 8.390 24.255 ;
        RECT 9.020 23.745 9.190 33.235 ;
        RECT 9.820 32.725 11.820 32.895 ;
        RECT 9.590 24.470 9.760 32.510 ;
        RECT 11.880 24.470 12.050 32.510 ;
        RECT 12.450 31.665 14.180 33.235 ;
        RECT 26.230 33.250 27.980 33.260 ;
        RECT 12.450 31.495 20.915 31.665 ;
        RECT 12.450 30.085 14.255 31.495 ;
        RECT 14.595 30.625 14.765 30.955 ;
        RECT 14.980 30.925 20.020 31.095 ;
        RECT 14.980 30.485 20.020 30.655 ;
        RECT 20.235 30.625 20.405 30.955 ;
        RECT 20.745 30.085 20.915 31.495 ;
        RECT 12.450 29.915 20.915 30.085 ;
        RECT 12.450 29.400 14.180 29.915 ;
        RECT 12.450 29.285 23.930 29.400 ;
        RECT 9.820 24.085 11.820 24.255 ;
        RECT 12.450 23.745 12.620 29.285 ;
        RECT 5.590 23.575 12.620 23.745 ;
        RECT 12.900 29.230 23.930 29.285 ;
        RECT 12.900 23.740 13.070 29.230 ;
        RECT 13.700 28.720 17.700 28.890 ;
        RECT 13.470 24.465 13.640 28.505 ;
        RECT 17.760 24.465 17.930 28.505 ;
        RECT 13.700 24.080 17.700 24.250 ;
        RECT 18.330 23.740 18.500 29.230 ;
        RECT 19.130 28.720 23.130 28.890 ;
        RECT 18.900 24.465 19.070 28.505 ;
        RECT 23.190 24.465 23.360 28.505 ;
        RECT 19.130 24.080 23.130 24.250 ;
        RECT 23.760 23.740 23.930 29.230 ;
        RECT 12.900 23.570 23.930 23.740 ;
        RECT 24.205 29.245 25.955 29.415 ;
        RECT 24.205 23.755 24.375 29.245 ;
        RECT 24.915 28.735 25.245 28.905 ;
        RECT 24.775 24.480 24.945 28.520 ;
        RECT 25.215 24.480 25.385 28.520 ;
        RECT 24.915 24.095 25.245 24.265 ;
        RECT 25.785 23.755 25.955 29.245 ;
        RECT 24.205 23.585 25.955 23.755 ;
        RECT 26.230 23.760 26.400 33.250 ;
        RECT 26.940 32.740 27.270 32.910 ;
        RECT 26.800 24.485 26.970 32.525 ;
        RECT 27.240 24.485 27.410 32.525 ;
        RECT 26.940 24.100 27.270 24.270 ;
        RECT 27.810 23.760 27.980 33.250 ;
        RECT 29.435 33.260 55.980 33.420 ;
        RECT 29.435 33.235 42.180 33.260 ;
        RECT 29.435 33.005 33.760 33.235 ;
        RECT 26.230 23.590 27.980 23.760 ;
        RECT 29.470 23.745 29.640 33.005 ;
        RECT 30.365 32.435 32.405 32.605 ;
        RECT 29.980 24.375 30.150 32.375 ;
        RECT 32.620 24.375 32.790 32.375 ;
        RECT 30.365 24.145 32.405 24.315 ;
        RECT 33.130 23.745 33.300 33.005 ;
        RECT 29.470 23.575 33.300 23.745 ;
        RECT 33.590 23.745 33.760 33.005 ;
        RECT 34.390 32.725 36.390 32.895 ;
        RECT 34.160 24.470 34.330 32.510 ;
        RECT 36.450 24.470 36.620 32.510 ;
        RECT 34.390 24.085 36.390 24.255 ;
        RECT 37.020 23.745 37.190 33.235 ;
        RECT 37.820 32.725 39.820 32.895 ;
        RECT 37.590 24.470 37.760 32.510 ;
        RECT 39.880 24.470 40.050 32.510 ;
        RECT 40.450 31.665 42.180 33.235 ;
        RECT 54.230 33.250 55.980 33.260 ;
        RECT 40.450 31.495 48.915 31.665 ;
        RECT 40.450 30.085 42.255 31.495 ;
        RECT 42.595 30.625 42.765 30.955 ;
        RECT 42.980 30.925 48.020 31.095 ;
        RECT 42.980 30.485 48.020 30.655 ;
        RECT 48.235 30.625 48.405 30.955 ;
        RECT 48.745 30.085 48.915 31.495 ;
        RECT 40.450 29.915 48.915 30.085 ;
        RECT 40.450 29.400 42.180 29.915 ;
        RECT 40.450 29.285 51.930 29.400 ;
        RECT 37.820 24.085 39.820 24.255 ;
        RECT 40.450 23.745 40.620 29.285 ;
        RECT 33.590 23.575 40.620 23.745 ;
        RECT 40.900 29.230 51.930 29.285 ;
        RECT 40.900 23.740 41.070 29.230 ;
        RECT 41.700 28.720 45.700 28.890 ;
        RECT 41.470 24.465 41.640 28.505 ;
        RECT 45.760 24.465 45.930 28.505 ;
        RECT 41.700 24.080 45.700 24.250 ;
        RECT 46.330 23.740 46.500 29.230 ;
        RECT 47.130 28.720 51.130 28.890 ;
        RECT 46.900 24.465 47.070 28.505 ;
        RECT 51.190 24.465 51.360 28.505 ;
        RECT 47.130 24.080 51.130 24.250 ;
        RECT 51.760 23.740 51.930 29.230 ;
        RECT 40.900 23.570 51.930 23.740 ;
        RECT 52.205 29.245 53.955 29.415 ;
        RECT 52.205 23.755 52.375 29.245 ;
        RECT 52.915 28.735 53.245 28.905 ;
        RECT 52.775 24.480 52.945 28.520 ;
        RECT 53.215 24.480 53.385 28.520 ;
        RECT 52.915 24.095 53.245 24.265 ;
        RECT 53.785 23.755 53.955 29.245 ;
        RECT 52.205 23.585 53.955 23.755 ;
        RECT 54.230 23.760 54.400 33.250 ;
        RECT 54.940 32.740 55.270 32.910 ;
        RECT 54.800 24.485 54.970 32.525 ;
        RECT 55.240 24.485 55.410 32.525 ;
        RECT 54.940 24.100 55.270 24.270 ;
        RECT 55.810 23.760 55.980 33.250 ;
        RECT 57.435 33.260 83.980 33.420 ;
        RECT 57.435 33.235 70.180 33.260 ;
        RECT 57.435 33.005 61.760 33.235 ;
        RECT 54.230 23.590 55.980 23.760 ;
        RECT 57.470 23.745 57.640 33.005 ;
        RECT 58.365 32.435 60.405 32.605 ;
        RECT 57.980 24.375 58.150 32.375 ;
        RECT 60.620 24.375 60.790 32.375 ;
        RECT 58.365 24.145 60.405 24.315 ;
        RECT 61.130 23.745 61.300 33.005 ;
        RECT 57.470 23.575 61.300 23.745 ;
        RECT 61.590 23.745 61.760 33.005 ;
        RECT 62.390 32.725 64.390 32.895 ;
        RECT 62.160 24.470 62.330 32.510 ;
        RECT 64.450 24.470 64.620 32.510 ;
        RECT 62.390 24.085 64.390 24.255 ;
        RECT 65.020 23.745 65.190 33.235 ;
        RECT 65.820 32.725 67.820 32.895 ;
        RECT 65.590 24.470 65.760 32.510 ;
        RECT 67.880 24.470 68.050 32.510 ;
        RECT 68.450 31.665 70.180 33.235 ;
        RECT 82.230 33.250 83.980 33.260 ;
        RECT 68.450 31.495 76.915 31.665 ;
        RECT 68.450 30.085 70.255 31.495 ;
        RECT 70.595 30.625 70.765 30.955 ;
        RECT 70.980 30.925 76.020 31.095 ;
        RECT 70.980 30.485 76.020 30.655 ;
        RECT 76.235 30.625 76.405 30.955 ;
        RECT 76.745 30.085 76.915 31.495 ;
        RECT 68.450 29.915 76.915 30.085 ;
        RECT 68.450 29.400 70.180 29.915 ;
        RECT 68.450 29.285 79.930 29.400 ;
        RECT 65.820 24.085 67.820 24.255 ;
        RECT 68.450 23.745 68.620 29.285 ;
        RECT 61.590 23.575 68.620 23.745 ;
        RECT 68.900 29.230 79.930 29.285 ;
        RECT 68.900 23.740 69.070 29.230 ;
        RECT 69.700 28.720 73.700 28.890 ;
        RECT 69.470 24.465 69.640 28.505 ;
        RECT 73.760 24.465 73.930 28.505 ;
        RECT 69.700 24.080 73.700 24.250 ;
        RECT 74.330 23.740 74.500 29.230 ;
        RECT 75.130 28.720 79.130 28.890 ;
        RECT 74.900 24.465 75.070 28.505 ;
        RECT 79.190 24.465 79.360 28.505 ;
        RECT 75.130 24.080 79.130 24.250 ;
        RECT 79.760 23.740 79.930 29.230 ;
        RECT 68.900 23.570 79.930 23.740 ;
        RECT 80.205 29.245 81.955 29.415 ;
        RECT 80.205 23.755 80.375 29.245 ;
        RECT 80.915 28.735 81.245 28.905 ;
        RECT 80.775 24.480 80.945 28.520 ;
        RECT 81.215 24.480 81.385 28.520 ;
        RECT 80.915 24.095 81.245 24.265 ;
        RECT 81.785 23.755 81.955 29.245 ;
        RECT 80.205 23.585 81.955 23.755 ;
        RECT 82.230 23.760 82.400 33.250 ;
        RECT 82.940 32.740 83.270 32.910 ;
        RECT 82.800 24.485 82.970 32.525 ;
        RECT 83.240 24.485 83.410 32.525 ;
        RECT 82.940 24.100 83.270 24.270 ;
        RECT 83.810 23.760 83.980 33.250 ;
        RECT 85.435 33.260 111.980 33.420 ;
        RECT 85.435 33.235 98.180 33.260 ;
        RECT 85.435 33.005 89.760 33.235 ;
        RECT 82.230 23.590 83.980 23.760 ;
        RECT 85.470 23.745 85.640 33.005 ;
        RECT 86.365 32.435 88.405 32.605 ;
        RECT 85.980 24.375 86.150 32.375 ;
        RECT 88.620 24.375 88.790 32.375 ;
        RECT 86.365 24.145 88.405 24.315 ;
        RECT 89.130 23.745 89.300 33.005 ;
        RECT 85.470 23.575 89.300 23.745 ;
        RECT 89.590 23.745 89.760 33.005 ;
        RECT 90.390 32.725 92.390 32.895 ;
        RECT 90.160 24.470 90.330 32.510 ;
        RECT 92.450 24.470 92.620 32.510 ;
        RECT 90.390 24.085 92.390 24.255 ;
        RECT 93.020 23.745 93.190 33.235 ;
        RECT 93.820 32.725 95.820 32.895 ;
        RECT 93.590 24.470 93.760 32.510 ;
        RECT 95.880 24.470 96.050 32.510 ;
        RECT 96.450 31.665 98.180 33.235 ;
        RECT 110.230 33.250 111.980 33.260 ;
        RECT 96.450 31.495 104.915 31.665 ;
        RECT 96.450 30.085 98.255 31.495 ;
        RECT 98.595 30.625 98.765 30.955 ;
        RECT 98.980 30.925 104.020 31.095 ;
        RECT 98.980 30.485 104.020 30.655 ;
        RECT 104.235 30.625 104.405 30.955 ;
        RECT 104.745 30.085 104.915 31.495 ;
        RECT 96.450 29.915 104.915 30.085 ;
        RECT 96.450 29.400 98.180 29.915 ;
        RECT 96.450 29.285 107.930 29.400 ;
        RECT 93.820 24.085 95.820 24.255 ;
        RECT 96.450 23.745 96.620 29.285 ;
        RECT 89.590 23.575 96.620 23.745 ;
        RECT 96.900 29.230 107.930 29.285 ;
        RECT 96.900 23.740 97.070 29.230 ;
        RECT 97.700 28.720 101.700 28.890 ;
        RECT 97.470 24.465 97.640 28.505 ;
        RECT 101.760 24.465 101.930 28.505 ;
        RECT 97.700 24.080 101.700 24.250 ;
        RECT 102.330 23.740 102.500 29.230 ;
        RECT 103.130 28.720 107.130 28.890 ;
        RECT 102.900 24.465 103.070 28.505 ;
        RECT 107.190 24.465 107.360 28.505 ;
        RECT 103.130 24.080 107.130 24.250 ;
        RECT 107.760 23.740 107.930 29.230 ;
        RECT 96.900 23.570 107.930 23.740 ;
        RECT 108.205 29.245 109.955 29.415 ;
        RECT 108.205 23.755 108.375 29.245 ;
        RECT 108.915 28.735 109.245 28.905 ;
        RECT 108.775 24.480 108.945 28.520 ;
        RECT 109.215 24.480 109.385 28.520 ;
        RECT 108.915 24.095 109.245 24.265 ;
        RECT 109.785 23.755 109.955 29.245 ;
        RECT 108.205 23.585 109.955 23.755 ;
        RECT 110.230 23.760 110.400 33.250 ;
        RECT 110.940 32.740 111.270 32.910 ;
        RECT 110.800 24.485 110.970 32.525 ;
        RECT 111.240 24.485 111.410 32.525 ;
        RECT 110.940 24.100 111.270 24.270 ;
        RECT 111.810 23.760 111.980 33.250 ;
        RECT 113.435 33.260 139.980 33.420 ;
        RECT 113.435 33.235 126.180 33.260 ;
        RECT 113.435 33.005 117.760 33.235 ;
        RECT 110.230 23.590 111.980 23.760 ;
        RECT 113.470 23.745 113.640 33.005 ;
        RECT 114.365 32.435 116.405 32.605 ;
        RECT 113.980 24.375 114.150 32.375 ;
        RECT 116.620 24.375 116.790 32.375 ;
        RECT 114.365 24.145 116.405 24.315 ;
        RECT 117.130 23.745 117.300 33.005 ;
        RECT 113.470 23.575 117.300 23.745 ;
        RECT 117.590 23.745 117.760 33.005 ;
        RECT 118.390 32.725 120.390 32.895 ;
        RECT 118.160 24.470 118.330 32.510 ;
        RECT 120.450 24.470 120.620 32.510 ;
        RECT 118.390 24.085 120.390 24.255 ;
        RECT 121.020 23.745 121.190 33.235 ;
        RECT 121.820 32.725 123.820 32.895 ;
        RECT 121.590 24.470 121.760 32.510 ;
        RECT 123.880 24.470 124.050 32.510 ;
        RECT 124.450 31.665 126.180 33.235 ;
        RECT 138.230 33.250 139.980 33.260 ;
        RECT 124.450 31.495 132.915 31.665 ;
        RECT 124.450 30.085 126.255 31.495 ;
        RECT 126.595 30.625 126.765 30.955 ;
        RECT 126.980 30.925 132.020 31.095 ;
        RECT 126.980 30.485 132.020 30.655 ;
        RECT 132.235 30.625 132.405 30.955 ;
        RECT 132.745 30.085 132.915 31.495 ;
        RECT 124.450 29.915 132.915 30.085 ;
        RECT 124.450 29.400 126.180 29.915 ;
        RECT 124.450 29.285 135.930 29.400 ;
        RECT 121.820 24.085 123.820 24.255 ;
        RECT 124.450 23.745 124.620 29.285 ;
        RECT 117.590 23.575 124.620 23.745 ;
        RECT 124.900 29.230 135.930 29.285 ;
        RECT 124.900 23.740 125.070 29.230 ;
        RECT 125.700 28.720 129.700 28.890 ;
        RECT 125.470 24.465 125.640 28.505 ;
        RECT 129.760 24.465 129.930 28.505 ;
        RECT 125.700 24.080 129.700 24.250 ;
        RECT 130.330 23.740 130.500 29.230 ;
        RECT 131.130 28.720 135.130 28.890 ;
        RECT 130.900 24.465 131.070 28.505 ;
        RECT 135.190 24.465 135.360 28.505 ;
        RECT 131.130 24.080 135.130 24.250 ;
        RECT 135.760 23.740 135.930 29.230 ;
        RECT 124.900 23.570 135.930 23.740 ;
        RECT 136.205 29.245 137.955 29.415 ;
        RECT 136.205 23.755 136.375 29.245 ;
        RECT 136.915 28.735 137.245 28.905 ;
        RECT 136.775 24.480 136.945 28.520 ;
        RECT 137.215 24.480 137.385 28.520 ;
        RECT 136.915 24.095 137.245 24.265 ;
        RECT 137.785 23.755 137.955 29.245 ;
        RECT 136.205 23.585 137.955 23.755 ;
        RECT 138.230 23.760 138.400 33.250 ;
        RECT 138.940 32.740 139.270 32.910 ;
        RECT 138.800 24.485 138.970 32.525 ;
        RECT 139.240 24.485 139.410 32.525 ;
        RECT 138.940 24.100 139.270 24.270 ;
        RECT 139.810 23.760 139.980 33.250 ;
        RECT 138.230 23.590 139.980 23.760 ;
        RECT 2.130 22.665 24.020 22.835 ;
        RECT 2.130 19.265 2.300 22.665 ;
        RECT 2.930 22.155 6.930 22.325 ;
        RECT 2.700 19.945 2.870 21.985 ;
        RECT 6.990 19.945 7.160 21.985 ;
        RECT 2.930 19.605 6.930 19.775 ;
        RECT 7.560 19.265 7.730 22.665 ;
        RECT 8.360 22.155 12.360 22.325 ;
        RECT 8.130 19.945 8.300 21.985 ;
        RECT 12.420 19.945 12.590 21.985 ;
        RECT 8.360 19.605 12.360 19.775 ;
        RECT 12.990 19.265 13.160 22.665 ;
        RECT 13.790 22.155 17.790 22.325 ;
        RECT 13.560 19.945 13.730 21.985 ;
        RECT 17.850 19.945 18.020 21.985 ;
        RECT 13.790 19.605 17.790 19.775 ;
        RECT 18.420 19.265 18.590 22.665 ;
        RECT 19.220 22.155 23.220 22.325 ;
        RECT 18.990 19.945 19.160 21.985 ;
        RECT 23.280 19.945 23.450 21.985 ;
        RECT 23.850 20.240 24.020 22.665 ;
        RECT 24.290 22.670 26.040 22.840 ;
        RECT 24.290 20.270 24.460 22.670 ;
        RECT 25.000 22.160 25.330 22.330 ;
        RECT 24.860 20.950 25.030 21.990 ;
        RECT 25.300 20.950 25.470 21.990 ;
        RECT 25.000 20.610 25.330 20.780 ;
        RECT 25.870 20.270 26.040 22.670 ;
        RECT 24.290 20.240 26.040 20.270 ;
        RECT 26.315 22.675 28.065 22.845 ;
        RECT 26.315 20.240 26.485 22.675 ;
        RECT 27.025 22.165 27.355 22.335 ;
        RECT 19.220 19.605 23.220 19.775 ;
        RECT 23.850 19.275 26.485 20.240 ;
        RECT 26.885 19.955 27.055 21.995 ;
        RECT 27.325 19.955 27.495 21.995 ;
        RECT 27.025 19.615 27.355 19.785 ;
        RECT 27.895 19.275 28.065 22.675 ;
        RECT 23.850 19.265 28.065 19.275 ;
        RECT 2.130 19.245 28.065 19.265 ;
        RECT 30.130 22.665 52.020 22.835 ;
        RECT 30.130 19.265 30.300 22.665 ;
        RECT 30.930 22.155 34.930 22.325 ;
        RECT 30.700 19.945 30.870 21.985 ;
        RECT 34.990 19.945 35.160 21.985 ;
        RECT 30.930 19.605 34.930 19.775 ;
        RECT 35.560 19.265 35.730 22.665 ;
        RECT 36.360 22.155 40.360 22.325 ;
        RECT 36.130 19.945 36.300 21.985 ;
        RECT 40.420 19.945 40.590 21.985 ;
        RECT 36.360 19.605 40.360 19.775 ;
        RECT 40.990 19.265 41.160 22.665 ;
        RECT 41.790 22.155 45.790 22.325 ;
        RECT 41.560 19.945 41.730 21.985 ;
        RECT 45.850 19.945 46.020 21.985 ;
        RECT 41.790 19.605 45.790 19.775 ;
        RECT 46.420 19.265 46.590 22.665 ;
        RECT 47.220 22.155 51.220 22.325 ;
        RECT 46.990 19.945 47.160 21.985 ;
        RECT 51.280 19.945 51.450 21.985 ;
        RECT 51.850 20.240 52.020 22.665 ;
        RECT 52.290 22.670 54.040 22.840 ;
        RECT 52.290 20.270 52.460 22.670 ;
        RECT 53.000 22.160 53.330 22.330 ;
        RECT 52.860 20.950 53.030 21.990 ;
        RECT 53.300 20.950 53.470 21.990 ;
        RECT 53.000 20.610 53.330 20.780 ;
        RECT 53.870 20.270 54.040 22.670 ;
        RECT 52.290 20.240 54.040 20.270 ;
        RECT 54.315 22.675 56.065 22.845 ;
        RECT 54.315 20.240 54.485 22.675 ;
        RECT 55.025 22.165 55.355 22.335 ;
        RECT 47.220 19.605 51.220 19.775 ;
        RECT 51.850 19.275 54.485 20.240 ;
        RECT 54.885 19.955 55.055 21.995 ;
        RECT 55.325 19.955 55.495 21.995 ;
        RECT 55.025 19.615 55.355 19.785 ;
        RECT 55.895 19.275 56.065 22.675 ;
        RECT 51.850 19.265 56.065 19.275 ;
        RECT 30.130 19.245 56.065 19.265 ;
        RECT 58.130 22.665 80.020 22.835 ;
        RECT 58.130 19.265 58.300 22.665 ;
        RECT 58.930 22.155 62.930 22.325 ;
        RECT 58.700 19.945 58.870 21.985 ;
        RECT 62.990 19.945 63.160 21.985 ;
        RECT 58.930 19.605 62.930 19.775 ;
        RECT 63.560 19.265 63.730 22.665 ;
        RECT 64.360 22.155 68.360 22.325 ;
        RECT 64.130 19.945 64.300 21.985 ;
        RECT 68.420 19.945 68.590 21.985 ;
        RECT 64.360 19.605 68.360 19.775 ;
        RECT 68.990 19.265 69.160 22.665 ;
        RECT 69.790 22.155 73.790 22.325 ;
        RECT 69.560 19.945 69.730 21.985 ;
        RECT 73.850 19.945 74.020 21.985 ;
        RECT 69.790 19.605 73.790 19.775 ;
        RECT 74.420 19.265 74.590 22.665 ;
        RECT 75.220 22.155 79.220 22.325 ;
        RECT 74.990 19.945 75.160 21.985 ;
        RECT 79.280 19.945 79.450 21.985 ;
        RECT 79.850 20.240 80.020 22.665 ;
        RECT 80.290 22.670 82.040 22.840 ;
        RECT 80.290 20.270 80.460 22.670 ;
        RECT 81.000 22.160 81.330 22.330 ;
        RECT 80.860 20.950 81.030 21.990 ;
        RECT 81.300 20.950 81.470 21.990 ;
        RECT 81.000 20.610 81.330 20.780 ;
        RECT 81.870 20.270 82.040 22.670 ;
        RECT 80.290 20.240 82.040 20.270 ;
        RECT 82.315 22.675 84.065 22.845 ;
        RECT 82.315 20.240 82.485 22.675 ;
        RECT 83.025 22.165 83.355 22.335 ;
        RECT 75.220 19.605 79.220 19.775 ;
        RECT 79.850 19.275 82.485 20.240 ;
        RECT 82.885 19.955 83.055 21.995 ;
        RECT 83.325 19.955 83.495 21.995 ;
        RECT 83.025 19.615 83.355 19.785 ;
        RECT 83.895 19.275 84.065 22.675 ;
        RECT 79.850 19.265 84.065 19.275 ;
        RECT 58.130 19.245 84.065 19.265 ;
        RECT 86.130 22.665 108.020 22.835 ;
        RECT 86.130 19.265 86.300 22.665 ;
        RECT 86.930 22.155 90.930 22.325 ;
        RECT 86.700 19.945 86.870 21.985 ;
        RECT 90.990 19.945 91.160 21.985 ;
        RECT 86.930 19.605 90.930 19.775 ;
        RECT 91.560 19.265 91.730 22.665 ;
        RECT 92.360 22.155 96.360 22.325 ;
        RECT 92.130 19.945 92.300 21.985 ;
        RECT 96.420 19.945 96.590 21.985 ;
        RECT 92.360 19.605 96.360 19.775 ;
        RECT 96.990 19.265 97.160 22.665 ;
        RECT 97.790 22.155 101.790 22.325 ;
        RECT 97.560 19.945 97.730 21.985 ;
        RECT 101.850 19.945 102.020 21.985 ;
        RECT 97.790 19.605 101.790 19.775 ;
        RECT 102.420 19.265 102.590 22.665 ;
        RECT 103.220 22.155 107.220 22.325 ;
        RECT 102.990 19.945 103.160 21.985 ;
        RECT 107.280 19.945 107.450 21.985 ;
        RECT 107.850 20.240 108.020 22.665 ;
        RECT 108.290 22.670 110.040 22.840 ;
        RECT 108.290 20.270 108.460 22.670 ;
        RECT 109.000 22.160 109.330 22.330 ;
        RECT 108.860 20.950 109.030 21.990 ;
        RECT 109.300 20.950 109.470 21.990 ;
        RECT 109.000 20.610 109.330 20.780 ;
        RECT 109.870 20.270 110.040 22.670 ;
        RECT 108.290 20.240 110.040 20.270 ;
        RECT 110.315 22.675 112.065 22.845 ;
        RECT 110.315 20.240 110.485 22.675 ;
        RECT 111.025 22.165 111.355 22.335 ;
        RECT 103.220 19.605 107.220 19.775 ;
        RECT 107.850 19.275 110.485 20.240 ;
        RECT 110.885 19.955 111.055 21.995 ;
        RECT 111.325 19.955 111.495 21.995 ;
        RECT 111.025 19.615 111.355 19.785 ;
        RECT 111.895 19.275 112.065 22.675 ;
        RECT 107.850 19.265 112.065 19.275 ;
        RECT 86.130 19.245 112.065 19.265 ;
        RECT 114.130 22.665 136.020 22.835 ;
        RECT 114.130 19.265 114.300 22.665 ;
        RECT 114.930 22.155 118.930 22.325 ;
        RECT 114.700 19.945 114.870 21.985 ;
        RECT 118.990 19.945 119.160 21.985 ;
        RECT 114.930 19.605 118.930 19.775 ;
        RECT 119.560 19.265 119.730 22.665 ;
        RECT 120.360 22.155 124.360 22.325 ;
        RECT 120.130 19.945 120.300 21.985 ;
        RECT 124.420 19.945 124.590 21.985 ;
        RECT 120.360 19.605 124.360 19.775 ;
        RECT 124.990 19.265 125.160 22.665 ;
        RECT 125.790 22.155 129.790 22.325 ;
        RECT 125.560 19.945 125.730 21.985 ;
        RECT 129.850 19.945 130.020 21.985 ;
        RECT 125.790 19.605 129.790 19.775 ;
        RECT 130.420 19.265 130.590 22.665 ;
        RECT 131.220 22.155 135.220 22.325 ;
        RECT 130.990 19.945 131.160 21.985 ;
        RECT 135.280 19.945 135.450 21.985 ;
        RECT 135.850 20.240 136.020 22.665 ;
        RECT 136.290 22.670 138.040 22.840 ;
        RECT 136.290 20.270 136.460 22.670 ;
        RECT 137.000 22.160 137.330 22.330 ;
        RECT 136.860 20.950 137.030 21.990 ;
        RECT 137.300 20.950 137.470 21.990 ;
        RECT 137.000 20.610 137.330 20.780 ;
        RECT 137.870 20.270 138.040 22.670 ;
        RECT 136.290 20.240 138.040 20.270 ;
        RECT 138.315 22.675 140.065 22.845 ;
        RECT 138.315 20.240 138.485 22.675 ;
        RECT 139.025 22.165 139.355 22.335 ;
        RECT 131.220 19.605 135.220 19.775 ;
        RECT 135.850 19.275 138.485 20.240 ;
        RECT 138.885 19.955 139.055 21.995 ;
        RECT 139.325 19.955 139.495 21.995 ;
        RECT 139.025 19.615 139.355 19.785 ;
        RECT 139.895 19.275 140.065 22.675 ;
        RECT 135.850 19.265 140.065 19.275 ;
        RECT 114.130 19.245 140.065 19.265 ;
        RECT 1.475 19.105 28.065 19.245 ;
        RECT 29.475 19.105 56.065 19.245 ;
        RECT 57.475 19.105 84.065 19.245 ;
        RECT 85.475 19.105 112.065 19.245 ;
        RECT 113.475 19.105 140.065 19.245 ;
        RECT 1.475 18.380 28.055 19.105 ;
        RECT 29.475 18.380 56.055 19.105 ;
        RECT 57.475 18.380 84.055 19.105 ;
        RECT 85.475 18.380 112.055 19.105 ;
        RECT 113.475 18.380 140.055 19.105 ;
        RECT 1.450 17.480 27.925 17.960 ;
        RECT 29.450 17.480 55.925 17.960 ;
        RECT 57.450 17.480 83.925 17.960 ;
        RECT 85.450 17.480 111.925 17.960 ;
        RECT 113.450 17.480 139.925 17.960 ;
        RECT 1.435 17.420 27.925 17.480 ;
        RECT 29.435 17.420 55.925 17.480 ;
        RECT 57.435 17.420 83.925 17.480 ;
        RECT 85.435 17.420 111.925 17.480 ;
        RECT 113.435 17.420 139.925 17.480 ;
        RECT 1.435 17.260 27.980 17.420 ;
        RECT 1.435 17.235 14.180 17.260 ;
        RECT 1.435 17.005 5.760 17.235 ;
        RECT 1.470 7.745 1.640 17.005 ;
        RECT 2.365 16.435 4.405 16.605 ;
        RECT 1.980 8.375 2.150 16.375 ;
        RECT 4.620 8.375 4.790 16.375 ;
        RECT 2.365 8.145 4.405 8.315 ;
        RECT 5.130 7.745 5.300 17.005 ;
        RECT 1.470 7.575 5.300 7.745 ;
        RECT 5.590 7.745 5.760 17.005 ;
        RECT 6.390 16.725 8.390 16.895 ;
        RECT 6.160 8.470 6.330 16.510 ;
        RECT 8.450 8.470 8.620 16.510 ;
        RECT 6.390 8.085 8.390 8.255 ;
        RECT 9.020 7.745 9.190 17.235 ;
        RECT 9.820 16.725 11.820 16.895 ;
        RECT 9.590 8.470 9.760 16.510 ;
        RECT 11.880 8.470 12.050 16.510 ;
        RECT 12.450 15.665 14.180 17.235 ;
        RECT 26.230 17.250 27.980 17.260 ;
        RECT 12.450 15.495 20.915 15.665 ;
        RECT 12.450 14.085 14.255 15.495 ;
        RECT 14.595 14.625 14.765 14.955 ;
        RECT 14.980 14.925 20.020 15.095 ;
        RECT 14.980 14.485 20.020 14.655 ;
        RECT 20.235 14.625 20.405 14.955 ;
        RECT 20.745 14.085 20.915 15.495 ;
        RECT 12.450 13.915 20.915 14.085 ;
        RECT 12.450 13.400 14.180 13.915 ;
        RECT 12.450 13.285 23.930 13.400 ;
        RECT 9.820 8.085 11.820 8.255 ;
        RECT 12.450 7.745 12.620 13.285 ;
        RECT 5.590 7.575 12.620 7.745 ;
        RECT 12.900 13.230 23.930 13.285 ;
        RECT 12.900 7.740 13.070 13.230 ;
        RECT 13.700 12.720 17.700 12.890 ;
        RECT 13.470 8.465 13.640 12.505 ;
        RECT 17.760 8.465 17.930 12.505 ;
        RECT 13.700 8.080 17.700 8.250 ;
        RECT 18.330 7.740 18.500 13.230 ;
        RECT 19.130 12.720 23.130 12.890 ;
        RECT 18.900 8.465 19.070 12.505 ;
        RECT 23.190 8.465 23.360 12.505 ;
        RECT 19.130 8.080 23.130 8.250 ;
        RECT 23.760 7.740 23.930 13.230 ;
        RECT 12.900 7.570 23.930 7.740 ;
        RECT 24.205 13.245 25.955 13.415 ;
        RECT 24.205 7.755 24.375 13.245 ;
        RECT 24.915 12.735 25.245 12.905 ;
        RECT 24.775 8.480 24.945 12.520 ;
        RECT 25.215 8.480 25.385 12.520 ;
        RECT 24.915 8.095 25.245 8.265 ;
        RECT 25.785 7.755 25.955 13.245 ;
        RECT 24.205 7.585 25.955 7.755 ;
        RECT 26.230 7.760 26.400 17.250 ;
        RECT 26.940 16.740 27.270 16.910 ;
        RECT 26.800 8.485 26.970 16.525 ;
        RECT 27.240 8.485 27.410 16.525 ;
        RECT 26.940 8.100 27.270 8.270 ;
        RECT 27.810 7.760 27.980 17.250 ;
        RECT 29.435 17.260 55.980 17.420 ;
        RECT 29.435 17.235 42.180 17.260 ;
        RECT 29.435 17.005 33.760 17.235 ;
        RECT 26.230 7.590 27.980 7.760 ;
        RECT 29.470 7.745 29.640 17.005 ;
        RECT 30.365 16.435 32.405 16.605 ;
        RECT 29.980 8.375 30.150 16.375 ;
        RECT 32.620 8.375 32.790 16.375 ;
        RECT 30.365 8.145 32.405 8.315 ;
        RECT 33.130 7.745 33.300 17.005 ;
        RECT 29.470 7.575 33.300 7.745 ;
        RECT 33.590 7.745 33.760 17.005 ;
        RECT 34.390 16.725 36.390 16.895 ;
        RECT 34.160 8.470 34.330 16.510 ;
        RECT 36.450 8.470 36.620 16.510 ;
        RECT 34.390 8.085 36.390 8.255 ;
        RECT 37.020 7.745 37.190 17.235 ;
        RECT 37.820 16.725 39.820 16.895 ;
        RECT 37.590 8.470 37.760 16.510 ;
        RECT 39.880 8.470 40.050 16.510 ;
        RECT 40.450 15.665 42.180 17.235 ;
        RECT 54.230 17.250 55.980 17.260 ;
        RECT 40.450 15.495 48.915 15.665 ;
        RECT 40.450 14.085 42.255 15.495 ;
        RECT 42.595 14.625 42.765 14.955 ;
        RECT 42.980 14.925 48.020 15.095 ;
        RECT 42.980 14.485 48.020 14.655 ;
        RECT 48.235 14.625 48.405 14.955 ;
        RECT 48.745 14.085 48.915 15.495 ;
        RECT 40.450 13.915 48.915 14.085 ;
        RECT 40.450 13.400 42.180 13.915 ;
        RECT 40.450 13.285 51.930 13.400 ;
        RECT 37.820 8.085 39.820 8.255 ;
        RECT 40.450 7.745 40.620 13.285 ;
        RECT 33.590 7.575 40.620 7.745 ;
        RECT 40.900 13.230 51.930 13.285 ;
        RECT 40.900 7.740 41.070 13.230 ;
        RECT 41.700 12.720 45.700 12.890 ;
        RECT 41.470 8.465 41.640 12.505 ;
        RECT 45.760 8.465 45.930 12.505 ;
        RECT 41.700 8.080 45.700 8.250 ;
        RECT 46.330 7.740 46.500 13.230 ;
        RECT 47.130 12.720 51.130 12.890 ;
        RECT 46.900 8.465 47.070 12.505 ;
        RECT 51.190 8.465 51.360 12.505 ;
        RECT 47.130 8.080 51.130 8.250 ;
        RECT 51.760 7.740 51.930 13.230 ;
        RECT 40.900 7.570 51.930 7.740 ;
        RECT 52.205 13.245 53.955 13.415 ;
        RECT 52.205 7.755 52.375 13.245 ;
        RECT 52.915 12.735 53.245 12.905 ;
        RECT 52.775 8.480 52.945 12.520 ;
        RECT 53.215 8.480 53.385 12.520 ;
        RECT 52.915 8.095 53.245 8.265 ;
        RECT 53.785 7.755 53.955 13.245 ;
        RECT 52.205 7.585 53.955 7.755 ;
        RECT 54.230 7.760 54.400 17.250 ;
        RECT 54.940 16.740 55.270 16.910 ;
        RECT 54.800 8.485 54.970 16.525 ;
        RECT 55.240 8.485 55.410 16.525 ;
        RECT 54.940 8.100 55.270 8.270 ;
        RECT 55.810 7.760 55.980 17.250 ;
        RECT 57.435 17.260 83.980 17.420 ;
        RECT 57.435 17.235 70.180 17.260 ;
        RECT 57.435 17.005 61.760 17.235 ;
        RECT 54.230 7.590 55.980 7.760 ;
        RECT 57.470 7.745 57.640 17.005 ;
        RECT 58.365 16.435 60.405 16.605 ;
        RECT 57.980 8.375 58.150 16.375 ;
        RECT 60.620 8.375 60.790 16.375 ;
        RECT 58.365 8.145 60.405 8.315 ;
        RECT 61.130 7.745 61.300 17.005 ;
        RECT 57.470 7.575 61.300 7.745 ;
        RECT 61.590 7.745 61.760 17.005 ;
        RECT 62.390 16.725 64.390 16.895 ;
        RECT 62.160 8.470 62.330 16.510 ;
        RECT 64.450 8.470 64.620 16.510 ;
        RECT 62.390 8.085 64.390 8.255 ;
        RECT 65.020 7.745 65.190 17.235 ;
        RECT 65.820 16.725 67.820 16.895 ;
        RECT 65.590 8.470 65.760 16.510 ;
        RECT 67.880 8.470 68.050 16.510 ;
        RECT 68.450 15.665 70.180 17.235 ;
        RECT 82.230 17.250 83.980 17.260 ;
        RECT 68.450 15.495 76.915 15.665 ;
        RECT 68.450 14.085 70.255 15.495 ;
        RECT 70.595 14.625 70.765 14.955 ;
        RECT 70.980 14.925 76.020 15.095 ;
        RECT 70.980 14.485 76.020 14.655 ;
        RECT 76.235 14.625 76.405 14.955 ;
        RECT 76.745 14.085 76.915 15.495 ;
        RECT 68.450 13.915 76.915 14.085 ;
        RECT 68.450 13.400 70.180 13.915 ;
        RECT 68.450 13.285 79.930 13.400 ;
        RECT 65.820 8.085 67.820 8.255 ;
        RECT 68.450 7.745 68.620 13.285 ;
        RECT 61.590 7.575 68.620 7.745 ;
        RECT 68.900 13.230 79.930 13.285 ;
        RECT 68.900 7.740 69.070 13.230 ;
        RECT 69.700 12.720 73.700 12.890 ;
        RECT 69.470 8.465 69.640 12.505 ;
        RECT 73.760 8.465 73.930 12.505 ;
        RECT 69.700 8.080 73.700 8.250 ;
        RECT 74.330 7.740 74.500 13.230 ;
        RECT 75.130 12.720 79.130 12.890 ;
        RECT 74.900 8.465 75.070 12.505 ;
        RECT 79.190 8.465 79.360 12.505 ;
        RECT 75.130 8.080 79.130 8.250 ;
        RECT 79.760 7.740 79.930 13.230 ;
        RECT 68.900 7.570 79.930 7.740 ;
        RECT 80.205 13.245 81.955 13.415 ;
        RECT 80.205 7.755 80.375 13.245 ;
        RECT 80.915 12.735 81.245 12.905 ;
        RECT 80.775 8.480 80.945 12.520 ;
        RECT 81.215 8.480 81.385 12.520 ;
        RECT 80.915 8.095 81.245 8.265 ;
        RECT 81.785 7.755 81.955 13.245 ;
        RECT 80.205 7.585 81.955 7.755 ;
        RECT 82.230 7.760 82.400 17.250 ;
        RECT 82.940 16.740 83.270 16.910 ;
        RECT 82.800 8.485 82.970 16.525 ;
        RECT 83.240 8.485 83.410 16.525 ;
        RECT 82.940 8.100 83.270 8.270 ;
        RECT 83.810 7.760 83.980 17.250 ;
        RECT 85.435 17.260 111.980 17.420 ;
        RECT 85.435 17.235 98.180 17.260 ;
        RECT 85.435 17.005 89.760 17.235 ;
        RECT 82.230 7.590 83.980 7.760 ;
        RECT 85.470 7.745 85.640 17.005 ;
        RECT 86.365 16.435 88.405 16.605 ;
        RECT 85.980 8.375 86.150 16.375 ;
        RECT 88.620 8.375 88.790 16.375 ;
        RECT 86.365 8.145 88.405 8.315 ;
        RECT 89.130 7.745 89.300 17.005 ;
        RECT 85.470 7.575 89.300 7.745 ;
        RECT 89.590 7.745 89.760 17.005 ;
        RECT 90.390 16.725 92.390 16.895 ;
        RECT 90.160 8.470 90.330 16.510 ;
        RECT 92.450 8.470 92.620 16.510 ;
        RECT 90.390 8.085 92.390 8.255 ;
        RECT 93.020 7.745 93.190 17.235 ;
        RECT 93.820 16.725 95.820 16.895 ;
        RECT 93.590 8.470 93.760 16.510 ;
        RECT 95.880 8.470 96.050 16.510 ;
        RECT 96.450 15.665 98.180 17.235 ;
        RECT 110.230 17.250 111.980 17.260 ;
        RECT 96.450 15.495 104.915 15.665 ;
        RECT 96.450 14.085 98.255 15.495 ;
        RECT 98.595 14.625 98.765 14.955 ;
        RECT 98.980 14.925 104.020 15.095 ;
        RECT 98.980 14.485 104.020 14.655 ;
        RECT 104.235 14.625 104.405 14.955 ;
        RECT 104.745 14.085 104.915 15.495 ;
        RECT 96.450 13.915 104.915 14.085 ;
        RECT 96.450 13.400 98.180 13.915 ;
        RECT 96.450 13.285 107.930 13.400 ;
        RECT 93.820 8.085 95.820 8.255 ;
        RECT 96.450 7.745 96.620 13.285 ;
        RECT 89.590 7.575 96.620 7.745 ;
        RECT 96.900 13.230 107.930 13.285 ;
        RECT 96.900 7.740 97.070 13.230 ;
        RECT 97.700 12.720 101.700 12.890 ;
        RECT 97.470 8.465 97.640 12.505 ;
        RECT 101.760 8.465 101.930 12.505 ;
        RECT 97.700 8.080 101.700 8.250 ;
        RECT 102.330 7.740 102.500 13.230 ;
        RECT 103.130 12.720 107.130 12.890 ;
        RECT 102.900 8.465 103.070 12.505 ;
        RECT 107.190 8.465 107.360 12.505 ;
        RECT 103.130 8.080 107.130 8.250 ;
        RECT 107.760 7.740 107.930 13.230 ;
        RECT 96.900 7.570 107.930 7.740 ;
        RECT 108.205 13.245 109.955 13.415 ;
        RECT 108.205 7.755 108.375 13.245 ;
        RECT 108.915 12.735 109.245 12.905 ;
        RECT 108.775 8.480 108.945 12.520 ;
        RECT 109.215 8.480 109.385 12.520 ;
        RECT 108.915 8.095 109.245 8.265 ;
        RECT 109.785 7.755 109.955 13.245 ;
        RECT 108.205 7.585 109.955 7.755 ;
        RECT 110.230 7.760 110.400 17.250 ;
        RECT 110.940 16.740 111.270 16.910 ;
        RECT 110.800 8.485 110.970 16.525 ;
        RECT 111.240 8.485 111.410 16.525 ;
        RECT 110.940 8.100 111.270 8.270 ;
        RECT 111.810 7.760 111.980 17.250 ;
        RECT 113.435 17.260 139.980 17.420 ;
        RECT 113.435 17.235 126.180 17.260 ;
        RECT 113.435 17.005 117.760 17.235 ;
        RECT 110.230 7.590 111.980 7.760 ;
        RECT 113.470 7.745 113.640 17.005 ;
        RECT 114.365 16.435 116.405 16.605 ;
        RECT 113.980 8.375 114.150 16.375 ;
        RECT 116.620 8.375 116.790 16.375 ;
        RECT 114.365 8.145 116.405 8.315 ;
        RECT 117.130 7.745 117.300 17.005 ;
        RECT 113.470 7.575 117.300 7.745 ;
        RECT 117.590 7.745 117.760 17.005 ;
        RECT 118.390 16.725 120.390 16.895 ;
        RECT 118.160 8.470 118.330 16.510 ;
        RECT 120.450 8.470 120.620 16.510 ;
        RECT 118.390 8.085 120.390 8.255 ;
        RECT 121.020 7.745 121.190 17.235 ;
        RECT 121.820 16.725 123.820 16.895 ;
        RECT 121.590 8.470 121.760 16.510 ;
        RECT 123.880 8.470 124.050 16.510 ;
        RECT 124.450 15.665 126.180 17.235 ;
        RECT 138.230 17.250 139.980 17.260 ;
        RECT 124.450 15.495 132.915 15.665 ;
        RECT 124.450 14.085 126.255 15.495 ;
        RECT 126.595 14.625 126.765 14.955 ;
        RECT 126.980 14.925 132.020 15.095 ;
        RECT 126.980 14.485 132.020 14.655 ;
        RECT 132.235 14.625 132.405 14.955 ;
        RECT 132.745 14.085 132.915 15.495 ;
        RECT 124.450 13.915 132.915 14.085 ;
        RECT 124.450 13.400 126.180 13.915 ;
        RECT 124.450 13.285 135.930 13.400 ;
        RECT 121.820 8.085 123.820 8.255 ;
        RECT 124.450 7.745 124.620 13.285 ;
        RECT 117.590 7.575 124.620 7.745 ;
        RECT 124.900 13.230 135.930 13.285 ;
        RECT 124.900 7.740 125.070 13.230 ;
        RECT 125.700 12.720 129.700 12.890 ;
        RECT 125.470 8.465 125.640 12.505 ;
        RECT 129.760 8.465 129.930 12.505 ;
        RECT 125.700 8.080 129.700 8.250 ;
        RECT 130.330 7.740 130.500 13.230 ;
        RECT 131.130 12.720 135.130 12.890 ;
        RECT 130.900 8.465 131.070 12.505 ;
        RECT 135.190 8.465 135.360 12.505 ;
        RECT 131.130 8.080 135.130 8.250 ;
        RECT 135.760 7.740 135.930 13.230 ;
        RECT 124.900 7.570 135.930 7.740 ;
        RECT 136.205 13.245 137.955 13.415 ;
        RECT 136.205 7.755 136.375 13.245 ;
        RECT 136.915 12.735 137.245 12.905 ;
        RECT 136.775 8.480 136.945 12.520 ;
        RECT 137.215 8.480 137.385 12.520 ;
        RECT 136.915 8.095 137.245 8.265 ;
        RECT 137.785 7.755 137.955 13.245 ;
        RECT 136.205 7.585 137.955 7.755 ;
        RECT 138.230 7.760 138.400 17.250 ;
        RECT 138.940 16.740 139.270 16.910 ;
        RECT 138.800 8.485 138.970 16.525 ;
        RECT 139.240 8.485 139.410 16.525 ;
        RECT 138.940 8.100 139.270 8.270 ;
        RECT 139.810 7.760 139.980 17.250 ;
        RECT 138.230 7.590 139.980 7.760 ;
        RECT 2.130 6.665 24.020 6.835 ;
        RECT 2.130 3.265 2.300 6.665 ;
        RECT 2.930 6.155 6.930 6.325 ;
        RECT 2.700 3.945 2.870 5.985 ;
        RECT 6.990 3.945 7.160 5.985 ;
        RECT 2.930 3.605 6.930 3.775 ;
        RECT 7.560 3.265 7.730 6.665 ;
        RECT 8.360 6.155 12.360 6.325 ;
        RECT 8.130 3.945 8.300 5.985 ;
        RECT 12.420 3.945 12.590 5.985 ;
        RECT 8.360 3.605 12.360 3.775 ;
        RECT 12.990 3.265 13.160 6.665 ;
        RECT 13.790 6.155 17.790 6.325 ;
        RECT 13.560 3.945 13.730 5.985 ;
        RECT 17.850 3.945 18.020 5.985 ;
        RECT 13.790 3.605 17.790 3.775 ;
        RECT 18.420 3.265 18.590 6.665 ;
        RECT 19.220 6.155 23.220 6.325 ;
        RECT 18.990 3.945 19.160 5.985 ;
        RECT 23.280 3.945 23.450 5.985 ;
        RECT 23.850 4.240 24.020 6.665 ;
        RECT 24.290 6.670 26.040 6.840 ;
        RECT 24.290 4.270 24.460 6.670 ;
        RECT 25.000 6.160 25.330 6.330 ;
        RECT 24.860 4.950 25.030 5.990 ;
        RECT 25.300 4.950 25.470 5.990 ;
        RECT 25.000 4.610 25.330 4.780 ;
        RECT 25.870 4.270 26.040 6.670 ;
        RECT 24.290 4.240 26.040 4.270 ;
        RECT 26.315 6.675 28.065 6.845 ;
        RECT 26.315 4.240 26.485 6.675 ;
        RECT 27.025 6.165 27.355 6.335 ;
        RECT 19.220 3.605 23.220 3.775 ;
        RECT 23.850 3.275 26.485 4.240 ;
        RECT 26.885 3.955 27.055 5.995 ;
        RECT 27.325 3.955 27.495 5.995 ;
        RECT 27.025 3.615 27.355 3.785 ;
        RECT 27.895 3.275 28.065 6.675 ;
        RECT 23.850 3.265 28.065 3.275 ;
        RECT 2.130 3.245 28.065 3.265 ;
        RECT 30.130 6.665 52.020 6.835 ;
        RECT 30.130 3.265 30.300 6.665 ;
        RECT 30.930 6.155 34.930 6.325 ;
        RECT 30.700 3.945 30.870 5.985 ;
        RECT 34.990 3.945 35.160 5.985 ;
        RECT 30.930 3.605 34.930 3.775 ;
        RECT 35.560 3.265 35.730 6.665 ;
        RECT 36.360 6.155 40.360 6.325 ;
        RECT 36.130 3.945 36.300 5.985 ;
        RECT 40.420 3.945 40.590 5.985 ;
        RECT 36.360 3.605 40.360 3.775 ;
        RECT 40.990 3.265 41.160 6.665 ;
        RECT 41.790 6.155 45.790 6.325 ;
        RECT 41.560 3.945 41.730 5.985 ;
        RECT 45.850 3.945 46.020 5.985 ;
        RECT 41.790 3.605 45.790 3.775 ;
        RECT 46.420 3.265 46.590 6.665 ;
        RECT 47.220 6.155 51.220 6.325 ;
        RECT 46.990 3.945 47.160 5.985 ;
        RECT 51.280 3.945 51.450 5.985 ;
        RECT 51.850 4.240 52.020 6.665 ;
        RECT 52.290 6.670 54.040 6.840 ;
        RECT 52.290 4.270 52.460 6.670 ;
        RECT 53.000 6.160 53.330 6.330 ;
        RECT 52.860 4.950 53.030 5.990 ;
        RECT 53.300 4.950 53.470 5.990 ;
        RECT 53.000 4.610 53.330 4.780 ;
        RECT 53.870 4.270 54.040 6.670 ;
        RECT 52.290 4.240 54.040 4.270 ;
        RECT 54.315 6.675 56.065 6.845 ;
        RECT 54.315 4.240 54.485 6.675 ;
        RECT 55.025 6.165 55.355 6.335 ;
        RECT 47.220 3.605 51.220 3.775 ;
        RECT 51.850 3.275 54.485 4.240 ;
        RECT 54.885 3.955 55.055 5.995 ;
        RECT 55.325 3.955 55.495 5.995 ;
        RECT 55.025 3.615 55.355 3.785 ;
        RECT 55.895 3.275 56.065 6.675 ;
        RECT 51.850 3.265 56.065 3.275 ;
        RECT 30.130 3.245 56.065 3.265 ;
        RECT 58.130 6.665 80.020 6.835 ;
        RECT 58.130 3.265 58.300 6.665 ;
        RECT 58.930 6.155 62.930 6.325 ;
        RECT 58.700 3.945 58.870 5.985 ;
        RECT 62.990 3.945 63.160 5.985 ;
        RECT 58.930 3.605 62.930 3.775 ;
        RECT 63.560 3.265 63.730 6.665 ;
        RECT 64.360 6.155 68.360 6.325 ;
        RECT 64.130 3.945 64.300 5.985 ;
        RECT 68.420 3.945 68.590 5.985 ;
        RECT 64.360 3.605 68.360 3.775 ;
        RECT 68.990 3.265 69.160 6.665 ;
        RECT 69.790 6.155 73.790 6.325 ;
        RECT 69.560 3.945 69.730 5.985 ;
        RECT 73.850 3.945 74.020 5.985 ;
        RECT 69.790 3.605 73.790 3.775 ;
        RECT 74.420 3.265 74.590 6.665 ;
        RECT 75.220 6.155 79.220 6.325 ;
        RECT 74.990 3.945 75.160 5.985 ;
        RECT 79.280 3.945 79.450 5.985 ;
        RECT 79.850 4.240 80.020 6.665 ;
        RECT 80.290 6.670 82.040 6.840 ;
        RECT 80.290 4.270 80.460 6.670 ;
        RECT 81.000 6.160 81.330 6.330 ;
        RECT 80.860 4.950 81.030 5.990 ;
        RECT 81.300 4.950 81.470 5.990 ;
        RECT 81.000 4.610 81.330 4.780 ;
        RECT 81.870 4.270 82.040 6.670 ;
        RECT 80.290 4.240 82.040 4.270 ;
        RECT 82.315 6.675 84.065 6.845 ;
        RECT 82.315 4.240 82.485 6.675 ;
        RECT 83.025 6.165 83.355 6.335 ;
        RECT 75.220 3.605 79.220 3.775 ;
        RECT 79.850 3.275 82.485 4.240 ;
        RECT 82.885 3.955 83.055 5.995 ;
        RECT 83.325 3.955 83.495 5.995 ;
        RECT 83.025 3.615 83.355 3.785 ;
        RECT 83.895 3.275 84.065 6.675 ;
        RECT 79.850 3.265 84.065 3.275 ;
        RECT 58.130 3.245 84.065 3.265 ;
        RECT 86.130 6.665 108.020 6.835 ;
        RECT 86.130 3.265 86.300 6.665 ;
        RECT 86.930 6.155 90.930 6.325 ;
        RECT 86.700 3.945 86.870 5.985 ;
        RECT 90.990 3.945 91.160 5.985 ;
        RECT 86.930 3.605 90.930 3.775 ;
        RECT 91.560 3.265 91.730 6.665 ;
        RECT 92.360 6.155 96.360 6.325 ;
        RECT 92.130 3.945 92.300 5.985 ;
        RECT 96.420 3.945 96.590 5.985 ;
        RECT 92.360 3.605 96.360 3.775 ;
        RECT 96.990 3.265 97.160 6.665 ;
        RECT 97.790 6.155 101.790 6.325 ;
        RECT 97.560 3.945 97.730 5.985 ;
        RECT 101.850 3.945 102.020 5.985 ;
        RECT 97.790 3.605 101.790 3.775 ;
        RECT 102.420 3.265 102.590 6.665 ;
        RECT 103.220 6.155 107.220 6.325 ;
        RECT 102.990 3.945 103.160 5.985 ;
        RECT 107.280 3.945 107.450 5.985 ;
        RECT 107.850 4.240 108.020 6.665 ;
        RECT 108.290 6.670 110.040 6.840 ;
        RECT 108.290 4.270 108.460 6.670 ;
        RECT 109.000 6.160 109.330 6.330 ;
        RECT 108.860 4.950 109.030 5.990 ;
        RECT 109.300 4.950 109.470 5.990 ;
        RECT 109.000 4.610 109.330 4.780 ;
        RECT 109.870 4.270 110.040 6.670 ;
        RECT 108.290 4.240 110.040 4.270 ;
        RECT 110.315 6.675 112.065 6.845 ;
        RECT 110.315 4.240 110.485 6.675 ;
        RECT 111.025 6.165 111.355 6.335 ;
        RECT 103.220 3.605 107.220 3.775 ;
        RECT 107.850 3.275 110.485 4.240 ;
        RECT 110.885 3.955 111.055 5.995 ;
        RECT 111.325 3.955 111.495 5.995 ;
        RECT 111.025 3.615 111.355 3.785 ;
        RECT 111.895 3.275 112.065 6.675 ;
        RECT 107.850 3.265 112.065 3.275 ;
        RECT 86.130 3.245 112.065 3.265 ;
        RECT 114.130 6.665 136.020 6.835 ;
        RECT 114.130 3.265 114.300 6.665 ;
        RECT 114.930 6.155 118.930 6.325 ;
        RECT 114.700 3.945 114.870 5.985 ;
        RECT 118.990 3.945 119.160 5.985 ;
        RECT 114.930 3.605 118.930 3.775 ;
        RECT 119.560 3.265 119.730 6.665 ;
        RECT 120.360 6.155 124.360 6.325 ;
        RECT 120.130 3.945 120.300 5.985 ;
        RECT 124.420 3.945 124.590 5.985 ;
        RECT 120.360 3.605 124.360 3.775 ;
        RECT 124.990 3.265 125.160 6.665 ;
        RECT 125.790 6.155 129.790 6.325 ;
        RECT 125.560 3.945 125.730 5.985 ;
        RECT 129.850 3.945 130.020 5.985 ;
        RECT 125.790 3.605 129.790 3.775 ;
        RECT 130.420 3.265 130.590 6.665 ;
        RECT 131.220 6.155 135.220 6.325 ;
        RECT 130.990 3.945 131.160 5.985 ;
        RECT 135.280 3.945 135.450 5.985 ;
        RECT 135.850 4.240 136.020 6.665 ;
        RECT 136.290 6.670 138.040 6.840 ;
        RECT 136.290 4.270 136.460 6.670 ;
        RECT 137.000 6.160 137.330 6.330 ;
        RECT 136.860 4.950 137.030 5.990 ;
        RECT 137.300 4.950 137.470 5.990 ;
        RECT 137.000 4.610 137.330 4.780 ;
        RECT 137.870 4.270 138.040 6.670 ;
        RECT 136.290 4.240 138.040 4.270 ;
        RECT 138.315 6.675 140.065 6.845 ;
        RECT 138.315 4.240 138.485 6.675 ;
        RECT 139.025 6.165 139.355 6.335 ;
        RECT 131.220 3.605 135.220 3.775 ;
        RECT 135.850 3.275 138.485 4.240 ;
        RECT 138.885 3.955 139.055 5.995 ;
        RECT 139.325 3.955 139.495 5.995 ;
        RECT 139.025 3.615 139.355 3.785 ;
        RECT 139.895 3.275 140.065 6.675 ;
        RECT 135.850 3.265 140.065 3.275 ;
        RECT 114.130 3.245 140.065 3.265 ;
        RECT 1.475 3.105 28.065 3.245 ;
        RECT 29.475 3.105 56.065 3.245 ;
        RECT 57.475 3.105 84.065 3.245 ;
        RECT 85.475 3.105 112.065 3.245 ;
        RECT 113.475 3.105 140.065 3.245 ;
        RECT 1.475 2.380 28.055 3.105 ;
        RECT 29.475 2.380 56.055 3.105 ;
        RECT 57.475 2.380 84.055 3.105 ;
        RECT 85.475 2.380 112.055 3.105 ;
        RECT 113.475 2.380 140.055 3.105 ;
      LAYER met1 ;
        RECT 35.490 223.220 35.810 223.280 ;
        RECT 79.650 223.220 79.970 223.280 ;
        RECT 35.490 223.080 79.970 223.220 ;
        RECT 35.490 223.020 35.810 223.080 ;
        RECT 79.650 223.020 79.970 223.080 ;
        RECT 22.610 220.500 22.930 220.560 ;
        RECT 82.410 220.500 82.730 220.560 ;
        RECT 22.610 220.360 82.730 220.500 ;
        RECT 22.610 220.300 22.930 220.360 ;
        RECT 82.410 220.300 82.730 220.360 ;
        RECT 54.810 218.800 55.130 218.860 ;
        RECT 67.230 218.800 67.550 218.860 ;
        RECT 54.810 218.660 67.550 218.800 ;
        RECT 54.810 218.600 55.130 218.660 ;
        RECT 67.230 218.600 67.550 218.660 ;
        RECT 48.370 218.460 48.690 218.520 ;
        RECT 75.510 218.460 75.830 218.520 ;
        RECT 48.370 218.320 75.830 218.460 ;
        RECT 48.370 218.260 48.690 218.320 ;
        RECT 75.510 218.260 75.830 218.320 ;
        RECT 41.930 218.120 42.250 218.180 ;
        RECT 81.030 218.120 81.350 218.180 ;
        RECT 41.930 217.980 81.350 218.120 ;
        RECT 41.930 217.920 42.250 217.980 ;
        RECT 81.030 217.920 81.350 217.980 ;
        RECT 51.590 217.780 51.910 217.840 ;
        RECT 71.370 217.780 71.690 217.840 ;
        RECT 51.590 217.640 71.690 217.780 ;
        RECT 51.590 217.580 51.910 217.640 ;
        RECT 71.370 217.580 71.690 217.640 ;
        RECT 45.150 217.440 45.470 217.500 ;
        RECT 76.890 217.440 77.210 217.500 ;
        RECT 45.150 217.300 77.210 217.440 ;
        RECT 45.150 217.240 45.470 217.300 ;
        RECT 76.890 217.240 77.210 217.300 ;
        RECT 38.710 217.100 39.030 217.160 ;
        RECT 75.970 217.100 76.290 217.160 ;
        RECT 38.710 216.960 76.290 217.100 ;
        RECT 38.710 216.900 39.030 216.960 ;
        RECT 75.970 216.900 76.290 216.960 ;
        RECT 54.810 215.740 55.130 215.800 ;
        RECT 61.710 215.740 62.030 215.800 ;
        RECT 54.810 215.600 70.450 215.740 ;
        RECT 54.810 215.540 55.130 215.600 ;
        RECT 61.710 215.540 62.030 215.600 ;
        RECT 58.030 215.400 58.350 215.460 ;
        RECT 68.610 215.400 68.930 215.460 ;
        RECT 58.030 215.260 68.930 215.400 ;
        RECT 70.310 215.400 70.450 215.600 ;
        RECT 92.070 215.400 92.390 215.460 ;
        RECT 70.310 215.260 92.390 215.400 ;
        RECT 58.030 215.200 58.350 215.260 ;
        RECT 68.610 215.200 68.930 215.260 ;
        RECT 92.070 215.200 92.390 215.260 ;
        RECT 34.110 215.060 34.430 215.120 ;
        RECT 66.770 215.060 67.090 215.120 ;
        RECT 34.110 214.920 67.090 215.060 ;
        RECT 34.110 214.860 34.430 214.920 ;
        RECT 66.770 214.860 67.090 214.920 ;
        RECT 48.830 214.720 49.150 214.780 ;
        RECT 84.710 214.720 85.030 214.780 ;
        RECT 48.830 214.580 85.030 214.720 ;
        RECT 48.830 214.520 49.150 214.580 ;
        RECT 84.710 214.520 85.030 214.580 ;
        RECT 57.570 214.380 57.890 214.440 ;
        RECT 81.950 214.380 82.270 214.440 ;
        RECT 57.570 214.240 82.270 214.380 ;
        RECT 57.570 214.180 57.890 214.240 ;
        RECT 81.950 214.180 82.270 214.240 ;
        RECT 33.650 214.040 33.970 214.100 ;
        RECT 77.810 214.040 78.130 214.100 ;
        RECT 33.650 213.900 78.130 214.040 ;
        RECT 33.650 213.840 33.970 213.900 ;
        RECT 77.810 213.840 78.130 213.900 ;
        RECT 58.490 213.700 58.810 213.760 ;
        RECT 73.670 213.700 73.990 213.760 ;
        RECT 58.490 213.560 73.990 213.700 ;
        RECT 58.490 213.500 58.810 213.560 ;
        RECT 73.670 213.500 73.990 213.560 ;
        RECT 48.370 213.360 48.690 213.420 ;
        RECT 76.430 213.360 76.750 213.420 ;
        RECT 48.370 213.220 76.750 213.360 ;
        RECT 48.370 213.160 48.690 213.220 ;
        RECT 76.430 213.160 76.750 213.220 ;
        RECT 14.260 212.540 126.960 213.020 ;
        RECT 20.770 212.340 21.090 212.400 ;
        RECT 34.570 212.340 34.890 212.400 ;
        RECT 35.505 212.340 35.795 212.385 ;
        RECT 20.770 212.200 34.340 212.340 ;
        RECT 20.770 212.140 21.090 212.200 ;
        RECT 23.530 212.000 23.850 212.060 ;
        RECT 16.720 211.860 23.850 212.000 ;
        RECT 16.720 211.705 16.860 211.860 ;
        RECT 23.530 211.800 23.850 211.860 ;
        RECT 23.990 211.800 24.310 212.060 ;
        RECT 33.650 211.800 33.970 212.060 ;
        RECT 34.200 212.000 34.340 212.200 ;
        RECT 34.570 212.200 35.795 212.340 ;
        RECT 34.570 212.140 34.890 212.200 ;
        RECT 35.505 212.155 35.795 212.200 ;
        RECT 48.920 212.200 66.540 212.340 ;
        RECT 35.965 212.000 36.255 212.045 ;
        RECT 46.070 212.000 46.390 212.060 ;
        RECT 34.200 211.860 35.720 212.000 ;
        RECT 16.645 211.475 16.935 211.705 ;
        RECT 18.010 211.460 18.330 211.720 ;
        RECT 30.890 211.660 31.210 211.720 ;
        RECT 34.585 211.660 34.875 211.705 ;
        RECT 30.890 211.520 34.875 211.660 ;
        RECT 35.580 211.660 35.720 211.860 ;
        RECT 35.965 211.860 46.390 212.000 ;
        RECT 35.965 211.815 36.255 211.860 ;
        RECT 46.070 211.800 46.390 211.860 ;
        RECT 46.530 212.000 46.850 212.060 ;
        RECT 48.920 212.045 49.060 212.200 ;
        RECT 48.845 212.000 49.135 212.045 ;
        RECT 46.530 211.860 49.135 212.000 ;
        RECT 46.530 211.800 46.850 211.860 ;
        RECT 48.845 211.815 49.135 211.860 ;
        RECT 53.430 212.000 53.750 212.060 ;
        RECT 60.345 212.000 60.635 212.045 ;
        RECT 53.430 211.860 65.620 212.000 ;
        RECT 53.430 211.800 53.750 211.860 ;
        RECT 60.345 211.815 60.635 211.860 ;
        RECT 35.580 211.520 37.100 211.660 ;
        RECT 30.890 211.460 31.210 211.520 ;
        RECT 34.585 211.475 34.875 211.520 ;
        RECT 17.105 211.320 17.395 211.365 ;
        RECT 19.850 211.320 20.170 211.380 ;
        RECT 17.105 211.180 20.170 211.320 ;
        RECT 17.105 211.135 17.395 211.180 ;
        RECT 19.850 211.120 20.170 211.180 ;
        RECT 20.310 211.320 20.630 211.380 ;
        RECT 21.705 211.320 21.995 211.365 ;
        RECT 20.310 211.180 21.995 211.320 ;
        RECT 20.310 211.120 20.630 211.180 ;
        RECT 21.705 211.135 21.995 211.180 ;
        RECT 23.085 211.320 23.375 211.365 ;
        RECT 32.270 211.320 32.590 211.380 ;
        RECT 23.085 211.180 32.590 211.320 ;
        RECT 23.085 211.135 23.375 211.180 ;
        RECT 32.270 211.120 32.590 211.180 ;
        RECT 32.730 211.320 33.050 211.380 ;
        RECT 35.490 211.320 35.810 211.380 ;
        RECT 32.730 211.180 35.810 211.320 ;
        RECT 36.960 211.320 37.100 211.520 ;
        RECT 37.330 211.460 37.650 211.720 ;
        RECT 39.630 211.460 39.950 211.720 ;
        RECT 40.090 211.460 40.410 211.720 ;
        RECT 42.850 211.660 43.170 211.720 ;
        RECT 49.765 211.660 50.055 211.705 ;
        RECT 42.850 211.520 50.055 211.660 ;
        RECT 42.850 211.460 43.170 211.520 ;
        RECT 49.765 211.475 50.055 211.520 ;
        RECT 59.425 211.660 59.715 211.705 ;
        RECT 60.790 211.660 61.110 211.720 ;
        RECT 59.425 211.520 61.110 211.660 ;
        RECT 59.425 211.475 59.715 211.520 ;
        RECT 60.790 211.460 61.110 211.520 ;
        RECT 61.710 211.460 62.030 211.720 ;
        RECT 63.090 211.460 63.410 211.720 ;
        RECT 65.480 211.705 65.620 211.860 ;
        RECT 66.400 211.705 66.540 212.200 ;
        RECT 68.610 212.140 68.930 212.400 ;
        RECT 69.070 212.340 69.390 212.400 ;
        RECT 70.465 212.340 70.755 212.385 ;
        RECT 69.070 212.200 70.755 212.340 ;
        RECT 69.070 212.140 69.390 212.200 ;
        RECT 70.465 212.155 70.755 212.200 ;
        RECT 71.370 212.140 71.690 212.400 ;
        RECT 75.510 212.140 75.830 212.400 ;
        RECT 76.890 212.140 77.210 212.400 ;
        RECT 81.030 212.140 81.350 212.400 ;
        RECT 82.410 212.140 82.730 212.400 ;
        RECT 83.790 212.140 84.110 212.400 ;
        RECT 89.770 212.140 90.090 212.400 ;
        RECT 97.680 212.200 101.500 212.340 ;
        RECT 66.770 212.000 67.090 212.060 ;
        RECT 66.770 211.860 72.520 212.000 ;
        RECT 66.770 211.800 67.090 211.860 ;
        RECT 65.405 211.475 65.695 211.705 ;
        RECT 66.325 211.475 66.615 211.705 ;
        RECT 67.690 211.460 68.010 211.720 ;
        RECT 70.005 211.660 70.295 211.705 ;
        RECT 70.450 211.660 70.770 211.720 ;
        RECT 70.005 211.520 70.770 211.660 ;
        RECT 70.005 211.475 70.295 211.520 ;
        RECT 70.450 211.460 70.770 211.520 ;
        RECT 70.925 211.660 71.215 211.705 ;
        RECT 71.370 211.660 71.690 211.720 ;
        RECT 72.380 211.705 72.520 211.860 ;
        RECT 79.650 211.800 79.970 212.060 ;
        RECT 70.925 211.520 71.690 211.660 ;
        RECT 70.925 211.475 71.215 211.520 ;
        RECT 71.370 211.460 71.690 211.520 ;
        RECT 72.305 211.475 72.595 211.705 ;
        RECT 73.670 211.460 73.990 211.720 ;
        RECT 76.430 211.460 76.750 211.720 ;
        RECT 77.350 211.660 77.670 211.720 ;
        RECT 77.825 211.660 78.115 211.705 ;
        RECT 77.350 211.520 78.115 211.660 ;
        RECT 77.350 211.460 77.670 211.520 ;
        RECT 77.825 211.475 78.115 211.520 ;
        RECT 78.285 211.475 78.575 211.705 ;
        RECT 78.360 211.320 78.500 211.475 ;
        RECT 81.950 211.460 82.270 211.720 ;
        RECT 84.710 211.460 85.030 211.720 ;
        RECT 86.565 211.475 86.855 211.705 ;
        RECT 89.325 211.660 89.615 211.705 ;
        RECT 89.860 211.660 90.000 212.140 ;
        RECT 92.070 212.000 92.390 212.060 ;
        RECT 93.005 212.000 93.295 212.045 ;
        RECT 92.070 211.860 93.295 212.000 ;
        RECT 92.070 211.800 92.390 211.860 ;
        RECT 93.005 211.815 93.295 211.860 ;
        RECT 93.925 212.000 94.215 212.045 ;
        RECT 96.670 212.000 96.990 212.060 ;
        RECT 93.925 211.860 96.990 212.000 ;
        RECT 93.925 211.815 94.215 211.860 ;
        RECT 96.670 211.800 96.990 211.860 ;
        RECT 89.325 211.520 90.000 211.660 ;
        RECT 92.545 211.660 92.835 211.705 ;
        RECT 93.450 211.660 93.770 211.720 ;
        RECT 92.545 211.520 93.770 211.660 ;
        RECT 89.325 211.475 89.615 211.520 ;
        RECT 92.545 211.475 92.835 211.520 ;
        RECT 36.960 211.180 78.500 211.320 ;
        RECT 82.410 211.320 82.730 211.380 ;
        RECT 86.640 211.320 86.780 211.475 ;
        RECT 93.450 211.460 93.770 211.520 ;
        RECT 95.750 211.460 96.070 211.720 ;
        RECT 97.680 211.705 97.820 212.200 ;
        RECT 101.360 212.000 101.500 212.200 ;
        RECT 104.965 212.155 105.255 212.385 ;
        RECT 105.040 212.000 105.180 212.155 ;
        RECT 101.360 211.860 105.180 212.000 ;
        RECT 97.605 211.475 97.895 211.705 ;
        RECT 102.665 211.660 102.955 211.705 ;
        RECT 103.110 211.660 103.430 211.720 ;
        RECT 102.665 211.520 103.430 211.660 ;
        RECT 102.665 211.475 102.955 211.520 ;
        RECT 92.990 211.320 93.310 211.380 ;
        RECT 97.680 211.320 97.820 211.475 ;
        RECT 103.110 211.460 103.430 211.520 ;
        RECT 105.870 211.460 106.190 211.720 ;
        RECT 109.105 211.660 109.395 211.705 ;
        RECT 109.550 211.660 109.870 211.720 ;
        RECT 109.105 211.520 109.870 211.660 ;
        RECT 109.105 211.475 109.395 211.520 ;
        RECT 109.550 211.460 109.870 211.520 ;
        RECT 112.325 211.660 112.615 211.705 ;
        RECT 112.770 211.660 113.090 211.720 ;
        RECT 112.325 211.520 113.090 211.660 ;
        RECT 112.325 211.475 112.615 211.520 ;
        RECT 112.770 211.460 113.090 211.520 ;
        RECT 82.410 211.180 85.860 211.320 ;
        RECT 86.640 211.180 90.460 211.320 ;
        RECT 32.730 211.120 33.050 211.180 ;
        RECT 35.490 211.120 35.810 211.180 ;
        RECT 82.410 211.120 82.730 211.180 ;
        RECT 17.550 210.780 17.870 211.040 ;
        RECT 35.030 210.980 35.350 211.040 ;
        RECT 42.850 210.980 43.170 211.040 ;
        RECT 35.030 210.840 43.170 210.980 ;
        RECT 35.030 210.780 35.350 210.840 ;
        RECT 42.850 210.780 43.170 210.840 ;
        RECT 66.785 210.795 67.075 211.025 ;
        RECT 67.230 210.980 67.550 211.040 ;
        RECT 72.765 210.980 73.055 211.025 ;
        RECT 67.230 210.840 73.055 210.980 ;
        RECT 15.710 210.440 16.030 210.700 ;
        RECT 35.950 210.640 36.270 210.700 ;
        RECT 37.805 210.640 38.095 210.685 ;
        RECT 35.950 210.500 38.095 210.640 ;
        RECT 35.950 210.440 36.270 210.500 ;
        RECT 37.805 210.455 38.095 210.500 ;
        RECT 46.070 210.640 46.390 210.700 ;
        RECT 49.290 210.640 49.610 210.700 ;
        RECT 46.070 210.500 49.610 210.640 ;
        RECT 46.070 210.440 46.390 210.500 ;
        RECT 49.290 210.440 49.610 210.500 ;
        RECT 49.750 210.640 50.070 210.700 ;
        RECT 56.205 210.640 56.495 210.685 ;
        RECT 63.090 210.640 63.410 210.700 ;
        RECT 49.750 210.500 63.410 210.640 ;
        RECT 66.860 210.640 67.000 210.795 ;
        RECT 67.230 210.780 67.550 210.840 ;
        RECT 72.765 210.795 73.055 210.840 ;
        RECT 73.210 210.980 73.530 211.040 ;
        RECT 85.720 211.025 85.860 211.180 ;
        RECT 90.320 211.040 90.460 211.180 ;
        RECT 92.990 211.180 97.820 211.320 ;
        RECT 92.990 211.120 93.310 211.180 ;
        RECT 98.050 211.120 98.370 211.380 ;
        RECT 73.210 210.840 84.940 210.980 ;
        RECT 73.210 210.780 73.530 210.840 ;
        RECT 77.350 210.640 77.670 210.700 ;
        RECT 66.860 210.500 77.670 210.640 ;
        RECT 84.800 210.640 84.940 210.840 ;
        RECT 85.645 210.795 85.935 211.025 ;
        RECT 88.390 210.780 88.710 211.040 ;
        RECT 90.230 210.980 90.550 211.040 ;
        RECT 108.185 210.980 108.475 211.025 ;
        RECT 90.230 210.840 108.475 210.980 ;
        RECT 90.230 210.780 90.550 210.840 ;
        RECT 108.185 210.795 108.475 210.840 ;
        RECT 91.610 210.640 91.930 210.700 ;
        RECT 84.800 210.500 91.930 210.640 ;
        RECT 49.750 210.440 50.070 210.500 ;
        RECT 56.205 210.455 56.495 210.500 ;
        RECT 63.090 210.440 63.410 210.500 ;
        RECT 77.350 210.440 77.670 210.500 ;
        RECT 91.610 210.440 91.930 210.500 ;
        RECT 94.830 210.440 95.150 210.700 ;
        RECT 95.290 210.640 95.610 210.700 ;
        RECT 95.765 210.640 96.055 210.685 ;
        RECT 95.290 210.500 96.055 210.640 ;
        RECT 95.290 210.440 95.610 210.500 ;
        RECT 95.765 210.455 96.055 210.500 ;
        RECT 101.745 210.640 102.035 210.685 ;
        RECT 104.030 210.640 104.350 210.700 ;
        RECT 101.745 210.500 104.350 210.640 ;
        RECT 101.745 210.455 102.035 210.500 ;
        RECT 104.030 210.440 104.350 210.500 ;
        RECT 109.090 210.640 109.410 210.700 ;
        RECT 111.405 210.640 111.695 210.685 ;
        RECT 109.090 210.500 111.695 210.640 ;
        RECT 109.090 210.440 109.410 210.500 ;
        RECT 111.405 210.455 111.695 210.500 ;
        RECT 14.260 209.820 126.960 210.300 ;
        RECT 33.650 209.420 33.970 209.680 ;
        RECT 34.110 209.620 34.430 209.680 ;
        RECT 34.585 209.620 34.875 209.665 ;
        RECT 45.150 209.620 45.470 209.680 ;
        RECT 34.110 209.480 34.875 209.620 ;
        RECT 34.110 209.420 34.430 209.480 ;
        RECT 34.585 209.435 34.875 209.480 ;
        RECT 35.120 209.480 45.470 209.620 ;
        RECT 35.120 209.280 35.260 209.480 ;
        RECT 45.150 209.420 45.470 209.480 ;
        RECT 49.290 209.620 49.610 209.680 ;
        RECT 59.425 209.620 59.715 209.665 ;
        RECT 61.250 209.620 61.570 209.680 ;
        RECT 63.550 209.620 63.870 209.680 ;
        RECT 67.230 209.620 67.550 209.680 ;
        RECT 49.290 209.480 56.880 209.620 ;
        RECT 49.290 209.420 49.610 209.480 ;
        RECT 17.180 209.140 35.260 209.280 ;
        RECT 35.490 209.280 35.810 209.340 ;
        RECT 56.740 209.280 56.880 209.480 ;
        RECT 59.425 209.480 61.570 209.620 ;
        RECT 59.425 209.435 59.715 209.480 ;
        RECT 61.250 209.420 61.570 209.480 ;
        RECT 63.180 209.480 67.550 209.620 ;
        RECT 60.805 209.280 61.095 209.325 ;
        RECT 35.490 209.140 49.980 209.280 ;
        RECT 56.740 209.140 61.095 209.280 ;
        RECT 17.180 208.645 17.320 209.140 ;
        RECT 35.490 209.080 35.810 209.140 ;
        RECT 21.690 208.940 22.010 209.000 ;
        RECT 23.085 208.940 23.375 208.985 ;
        RECT 39.630 208.940 39.950 209.000 ;
        RECT 21.690 208.800 23.375 208.940 ;
        RECT 21.690 208.740 22.010 208.800 ;
        RECT 23.085 208.755 23.375 208.800 ;
        RECT 34.660 208.800 39.950 208.940 ;
        RECT 17.105 208.415 17.395 208.645 ;
        RECT 18.485 208.415 18.775 208.645 ;
        RECT 19.405 208.415 19.695 208.645 ;
        RECT 15.250 208.260 15.570 208.320 ;
        RECT 18.560 208.260 18.700 208.415 ;
        RECT 15.250 208.120 18.700 208.260 ;
        RECT 19.480 208.260 19.620 208.415 ;
        RECT 20.310 208.400 20.630 208.660 ;
        RECT 22.165 208.600 22.455 208.645 ;
        RECT 29.050 208.600 29.370 208.660 ;
        RECT 22.165 208.460 29.370 208.600 ;
        RECT 22.165 208.415 22.455 208.460 ;
        RECT 29.050 208.400 29.370 208.460 ;
        RECT 23.070 208.260 23.390 208.320 ;
        RECT 19.480 208.120 23.390 208.260 ;
        RECT 15.250 208.060 15.570 208.120 ;
        RECT 23.070 208.060 23.390 208.120 ;
        RECT 24.005 208.075 24.295 208.305 ;
        RECT 32.270 208.260 32.590 208.320 ;
        RECT 34.660 208.305 34.800 208.800 ;
        RECT 39.630 208.740 39.950 208.800 ;
        RECT 46.530 208.740 46.850 209.000 ;
        RECT 35.950 208.400 36.270 208.660 ;
        RECT 46.990 208.400 47.310 208.660 ;
        RECT 49.840 208.645 49.980 209.140 ;
        RECT 60.805 209.095 61.095 209.140 ;
        RECT 61.265 208.940 61.555 208.985 ;
        RECT 63.180 208.940 63.320 209.480 ;
        RECT 63.550 209.420 63.870 209.480 ;
        RECT 67.230 209.420 67.550 209.480 ;
        RECT 67.705 209.620 67.995 209.665 ;
        RECT 69.530 209.620 69.850 209.680 ;
        RECT 67.705 209.480 69.850 209.620 ;
        RECT 67.705 209.435 67.995 209.480 ;
        RECT 69.530 209.420 69.850 209.480 ;
        RECT 71.370 209.620 71.690 209.680 ;
        RECT 75.510 209.620 75.830 209.680 ;
        RECT 71.370 209.480 75.830 209.620 ;
        RECT 71.370 209.420 71.690 209.480 ;
        RECT 75.510 209.420 75.830 209.480 ;
        RECT 75.970 209.620 76.290 209.680 ;
        RECT 76.905 209.620 77.195 209.665 ;
        RECT 75.970 209.480 77.195 209.620 ;
        RECT 75.970 209.420 76.290 209.480 ;
        RECT 76.905 209.435 77.195 209.480 ;
        RECT 77.350 209.620 77.670 209.680 ;
        RECT 78.270 209.620 78.590 209.680 ;
        RECT 86.550 209.620 86.870 209.680 ;
        RECT 77.350 209.480 78.590 209.620 ;
        RECT 77.350 209.420 77.670 209.480 ;
        RECT 78.270 209.420 78.590 209.480 ;
        RECT 78.820 209.480 86.870 209.620 ;
        RECT 78.820 209.280 78.960 209.480 ;
        RECT 86.550 209.420 86.870 209.480 ;
        RECT 87.025 209.435 87.315 209.665 ;
        RECT 87.930 209.620 88.250 209.680 ;
        RECT 91.165 209.620 91.455 209.665 ;
        RECT 95.750 209.620 96.070 209.680 ;
        RECT 87.930 209.480 96.070 209.620 ;
        RECT 87.100 209.280 87.240 209.435 ;
        RECT 87.930 209.420 88.250 209.480 ;
        RECT 91.165 209.435 91.455 209.480 ;
        RECT 95.750 209.420 96.070 209.480 ;
        RECT 125.205 209.620 125.495 209.665 ;
        RECT 128.410 209.620 128.730 209.680 ;
        RECT 125.205 209.480 128.730 209.620 ;
        RECT 125.205 209.435 125.495 209.480 ;
        RECT 128.410 209.420 128.730 209.480 ;
        RECT 97.130 209.280 97.450 209.340 ;
        RECT 72.380 209.140 78.960 209.280 ;
        RECT 83.420 209.140 97.450 209.280 ;
        RECT 61.265 208.800 63.320 208.940 ;
        RECT 63.565 208.940 63.855 208.985 ;
        RECT 71.830 208.940 72.150 209.000 ;
        RECT 63.565 208.800 72.150 208.940 ;
        RECT 61.265 208.755 61.555 208.800 ;
        RECT 63.565 208.755 63.855 208.800 ;
        RECT 71.830 208.740 72.150 208.800 ;
        RECT 48.845 208.600 49.135 208.645 ;
        RECT 48.845 208.460 49.520 208.600 ;
        RECT 48.845 208.415 49.135 208.460 ;
        RECT 32.745 208.260 33.035 208.305 ;
        RECT 32.270 208.120 33.035 208.260 ;
        RECT 16.185 207.920 16.475 207.965 ;
        RECT 17.090 207.920 17.410 207.980 ;
        RECT 16.185 207.780 17.410 207.920 ;
        RECT 16.185 207.735 16.475 207.780 ;
        RECT 17.090 207.720 17.410 207.780 ;
        RECT 18.010 207.920 18.330 207.980 ;
        RECT 20.785 207.920 21.075 207.965 ;
        RECT 18.010 207.780 21.075 207.920 ;
        RECT 18.010 207.720 18.330 207.780 ;
        RECT 20.785 207.735 21.075 207.780 ;
        RECT 22.150 207.920 22.470 207.980 ;
        RECT 24.080 207.920 24.220 208.075 ;
        RECT 32.270 208.060 32.590 208.120 ;
        RECT 32.745 208.075 33.035 208.120 ;
        RECT 34.585 208.075 34.875 208.305 ;
        RECT 35.505 208.260 35.795 208.305 ;
        RECT 37.330 208.260 37.650 208.320 ;
        RECT 35.505 208.120 37.650 208.260 ;
        RECT 49.380 208.260 49.520 208.460 ;
        RECT 49.765 208.415 50.055 208.645 ;
        RECT 60.330 208.400 60.650 208.660 ;
        RECT 62.170 208.400 62.490 208.660 ;
        RECT 63.090 208.400 63.410 208.660 ;
        RECT 64.025 208.415 64.315 208.645 ;
        RECT 54.810 208.260 55.130 208.320 ;
        RECT 64.100 208.260 64.240 208.415 ;
        RECT 64.930 208.400 65.250 208.660 ;
        RECT 66.770 208.400 67.090 208.660 ;
        RECT 67.705 208.600 67.995 208.645 ;
        RECT 68.610 208.600 68.930 208.660 ;
        RECT 67.705 208.460 68.930 208.600 ;
        RECT 67.705 208.415 67.995 208.460 ;
        RECT 49.380 208.120 55.130 208.260 ;
        RECT 35.505 208.075 35.795 208.120 ;
        RECT 37.330 208.060 37.650 208.120 ;
        RECT 54.810 208.060 55.130 208.120 ;
        RECT 56.280 208.120 64.240 208.260 ;
        RECT 64.470 208.260 64.790 208.320 ;
        RECT 67.780 208.260 67.920 208.415 ;
        RECT 68.610 208.400 68.930 208.460 ;
        RECT 69.085 208.600 69.375 208.645 ;
        RECT 69.990 208.600 70.310 208.660 ;
        RECT 69.085 208.460 70.310 208.600 ;
        RECT 69.085 208.415 69.375 208.460 ;
        RECT 69.990 208.400 70.310 208.460 ;
        RECT 70.910 208.600 71.230 208.660 ;
        RECT 72.380 208.645 72.520 209.140 ;
        RECT 72.750 208.940 73.070 209.000 ;
        RECT 75.985 208.940 76.275 208.985 ;
        RECT 72.750 208.800 76.275 208.940 ;
        RECT 72.750 208.740 73.070 208.800 ;
        RECT 75.985 208.755 76.275 208.800 ;
        RECT 77.350 208.940 77.670 209.000 ;
        RECT 78.745 208.940 79.035 208.985 ;
        RECT 77.350 208.800 79.035 208.940 ;
        RECT 77.350 208.740 77.670 208.800 ;
        RECT 78.745 208.755 79.035 208.800 ;
        RECT 79.190 208.940 79.510 209.000 ;
        RECT 83.420 208.940 83.560 209.140 ;
        RECT 97.130 209.080 97.450 209.140 ;
        RECT 89.310 208.940 89.630 209.000 ;
        RECT 91.150 208.940 91.470 209.000 ;
        RECT 79.190 208.800 83.560 208.940 ;
        RECT 79.190 208.740 79.510 208.800 ;
        RECT 72.305 208.600 72.595 208.645 ;
        RECT 70.910 208.460 72.595 208.600 ;
        RECT 70.910 208.400 71.230 208.460 ;
        RECT 72.305 208.415 72.595 208.460 ;
        RECT 73.670 208.400 73.990 208.660 ;
        RECT 74.605 208.415 74.895 208.645 ;
        RECT 75.525 208.415 75.815 208.645 ;
        RECT 76.445 208.600 76.735 208.645 ;
        RECT 76.890 208.600 77.210 208.660 ;
        RECT 76.445 208.460 77.210 208.600 ;
        RECT 76.445 208.415 76.735 208.460 ;
        RECT 74.680 208.260 74.820 208.415 ;
        RECT 64.470 208.120 67.920 208.260 ;
        RECT 71.000 208.120 74.820 208.260 ;
        RECT 75.600 208.260 75.740 208.415 ;
        RECT 76.890 208.400 77.210 208.460 ;
        RECT 77.810 208.400 78.130 208.660 ;
        RECT 78.270 208.400 78.590 208.660 ;
        RECT 80.570 208.400 80.890 208.660 ;
        RECT 81.950 208.400 82.270 208.660 ;
        RECT 82.410 208.400 82.730 208.660 ;
        RECT 83.420 208.645 83.560 208.800 ;
        RECT 84.110 208.800 89.630 208.940 ;
        RECT 83.345 208.415 83.635 208.645 ;
        RECT 75.970 208.260 76.290 208.320 ;
        RECT 82.500 208.260 82.640 208.400 ;
        RECT 84.110 208.260 84.250 208.800 ;
        RECT 89.310 208.740 89.630 208.800 ;
        RECT 89.860 208.800 91.470 208.940 ;
        RECT 87.025 208.600 87.315 208.645 ;
        RECT 87.930 208.600 88.250 208.660 ;
        RECT 87.025 208.460 88.250 208.600 ;
        RECT 87.025 208.415 87.315 208.460 ;
        RECT 87.930 208.400 88.250 208.460 ;
        RECT 88.865 208.600 89.155 208.645 ;
        RECT 89.860 208.600 90.000 208.800 ;
        RECT 91.150 208.740 91.470 208.800 ;
        RECT 91.610 208.940 91.930 209.000 ;
        RECT 91.610 208.800 98.280 208.940 ;
        RECT 91.610 208.740 91.930 208.800 ;
        RECT 88.865 208.460 90.000 208.600 ;
        RECT 88.865 208.415 89.155 208.460 ;
        RECT 90.230 208.400 90.550 208.660 ;
        RECT 92.070 208.400 92.390 208.660 ;
        RECT 95.290 208.400 95.610 208.660 ;
        RECT 95.750 208.600 96.070 208.660 ;
        RECT 96.225 208.600 96.515 208.645 ;
        RECT 95.750 208.460 96.515 208.600 ;
        RECT 95.750 208.400 96.070 208.460 ;
        RECT 96.225 208.415 96.515 208.460 ;
        RECT 97.130 208.400 97.450 208.660 ;
        RECT 98.140 208.645 98.280 208.800 ;
        RECT 98.065 208.415 98.355 208.645 ;
        RECT 75.600 208.120 76.290 208.260 ;
        RECT 22.150 207.780 24.220 207.920 ;
        RECT 35.950 207.920 36.270 207.980 ;
        RECT 40.090 207.920 40.410 207.980 ;
        RECT 42.405 207.920 42.695 207.965 ;
        RECT 35.950 207.780 42.695 207.920 ;
        RECT 22.150 207.720 22.470 207.780 ;
        RECT 35.950 207.720 36.270 207.780 ;
        RECT 40.090 207.720 40.410 207.780 ;
        RECT 42.405 207.735 42.695 207.780 ;
        RECT 48.370 207.720 48.690 207.980 ;
        RECT 55.270 207.920 55.590 207.980 ;
        RECT 56.280 207.965 56.420 208.120 ;
        RECT 64.470 208.060 64.790 208.120 ;
        RECT 71.000 207.980 71.140 208.120 ;
        RECT 75.970 208.060 76.290 208.120 ;
        RECT 77.900 208.120 82.640 208.260 ;
        RECT 83.420 208.120 84.250 208.260 ;
        RECT 77.900 207.980 78.040 208.120 ;
        RECT 56.205 207.920 56.495 207.965 ;
        RECT 55.270 207.780 56.495 207.920 ;
        RECT 55.270 207.720 55.590 207.780 ;
        RECT 56.205 207.735 56.495 207.780 ;
        RECT 59.870 207.920 60.190 207.980 ;
        RECT 61.725 207.920 62.015 207.965 ;
        RECT 59.870 207.780 62.015 207.920 ;
        RECT 59.870 207.720 60.190 207.780 ;
        RECT 61.725 207.735 62.015 207.780 ;
        RECT 65.850 207.720 66.170 207.980 ;
        RECT 68.150 207.920 68.470 207.980 ;
        RECT 68.625 207.920 68.915 207.965 ;
        RECT 68.150 207.780 68.915 207.920 ;
        RECT 68.150 207.720 68.470 207.780 ;
        RECT 68.625 207.735 68.915 207.780 ;
        RECT 69.070 207.920 69.390 207.980 ;
        RECT 69.545 207.920 69.835 207.965 ;
        RECT 69.070 207.780 69.835 207.920 ;
        RECT 69.070 207.720 69.390 207.780 ;
        RECT 69.545 207.735 69.835 207.780 ;
        RECT 70.910 207.720 71.230 207.980 ;
        RECT 71.370 207.720 71.690 207.980 ;
        RECT 77.810 207.720 78.130 207.980 ;
        RECT 78.730 207.920 79.050 207.980 ;
        RECT 79.665 207.920 79.955 207.965 ;
        RECT 78.730 207.780 79.955 207.920 ;
        RECT 78.730 207.720 79.050 207.780 ;
        RECT 79.665 207.735 79.955 207.780 ;
        RECT 81.950 207.920 82.270 207.980 ;
        RECT 83.420 207.920 83.560 208.120 ;
        RECT 85.170 208.060 85.490 208.320 ;
        RECT 93.910 208.060 94.230 208.320 ;
        RECT 81.950 207.780 83.560 207.920 ;
        RECT 83.790 207.920 84.110 207.980 ;
        RECT 86.105 207.920 86.395 207.965 ;
        RECT 83.790 207.780 86.395 207.920 ;
        RECT 81.950 207.720 82.270 207.780 ;
        RECT 83.790 207.720 84.110 207.780 ;
        RECT 86.105 207.735 86.395 207.780 ;
        RECT 93.005 207.920 93.295 207.965 ;
        RECT 94.370 207.920 94.690 207.980 ;
        RECT 95.290 207.920 95.610 207.980 ;
        RECT 93.005 207.780 95.610 207.920 ;
        RECT 93.005 207.735 93.295 207.780 ;
        RECT 94.370 207.720 94.690 207.780 ;
        RECT 95.290 207.720 95.610 207.780 ;
        RECT 97.130 207.920 97.450 207.980 ;
        RECT 98.050 207.920 98.370 207.980 ;
        RECT 98.985 207.920 99.275 207.965 ;
        RECT 97.130 207.780 99.275 207.920 ;
        RECT 97.130 207.720 97.450 207.780 ;
        RECT 98.050 207.720 98.370 207.780 ;
        RECT 98.985 207.735 99.275 207.780 ;
        RECT 14.260 207.100 126.960 207.580 ;
        RECT 17.105 206.900 17.395 206.945 ;
        RECT 28.590 206.900 28.910 206.960 ;
        RECT 17.105 206.760 28.910 206.900 ;
        RECT 17.105 206.715 17.395 206.760 ;
        RECT 28.590 206.700 28.910 206.760 ;
        RECT 29.510 206.900 29.830 206.960 ;
        RECT 34.570 206.900 34.890 206.960 ;
        RECT 29.510 206.760 34.890 206.900 ;
        RECT 29.510 206.700 29.830 206.760 ;
        RECT 34.570 206.700 34.890 206.760 ;
        RECT 37.330 206.900 37.650 206.960 ;
        RECT 44.230 206.900 44.550 206.960 ;
        RECT 51.590 206.900 51.910 206.960 ;
        RECT 37.330 206.760 51.910 206.900 ;
        RECT 37.330 206.700 37.650 206.760 ;
        RECT 44.230 206.700 44.550 206.760 ;
        RECT 51.590 206.700 51.910 206.760 ;
        RECT 53.905 206.900 54.195 206.945 ;
        RECT 58.490 206.900 58.810 206.960 ;
        RECT 53.905 206.760 58.810 206.900 ;
        RECT 53.905 206.715 54.195 206.760 ;
        RECT 58.490 206.700 58.810 206.760 ;
        RECT 59.870 206.700 60.190 206.960 ;
        RECT 60.790 206.900 61.110 206.960 ;
        RECT 62.630 206.900 62.950 206.960 ;
        RECT 60.420 206.760 62.950 206.900 ;
        RECT 26.765 206.560 27.055 206.605 ;
        RECT 32.730 206.560 33.050 206.620 ;
        RECT 26.765 206.420 33.050 206.560 ;
        RECT 26.765 206.375 27.055 206.420 ;
        RECT 32.730 206.360 33.050 206.420 ;
        RECT 46.990 206.560 47.310 206.620 ;
        RECT 51.145 206.560 51.435 206.605 ;
        RECT 60.420 206.560 60.560 206.760 ;
        RECT 60.790 206.700 61.110 206.760 ;
        RECT 62.630 206.700 62.950 206.760 ;
        RECT 63.090 206.900 63.410 206.960 ;
        RECT 66.785 206.900 67.075 206.945 ;
        RECT 63.090 206.760 67.075 206.900 ;
        RECT 63.090 206.700 63.410 206.760 ;
        RECT 66.785 206.715 67.075 206.760 ;
        RECT 67.230 206.900 67.550 206.960 ;
        RECT 68.610 206.900 68.930 206.960 ;
        RECT 67.230 206.760 68.930 206.900 ;
        RECT 67.230 206.700 67.550 206.760 ;
        RECT 68.610 206.700 68.930 206.760 ;
        RECT 70.450 206.900 70.770 206.960 ;
        RECT 74.130 206.900 74.450 206.960 ;
        RECT 70.450 206.760 74.450 206.900 ;
        RECT 70.450 206.700 70.770 206.760 ;
        RECT 74.130 206.700 74.450 206.760 ;
        RECT 76.430 206.900 76.750 206.960 ;
        RECT 81.965 206.900 82.255 206.945 ;
        RECT 76.430 206.760 82.255 206.900 ;
        RECT 76.430 206.700 76.750 206.760 ;
        RECT 81.965 206.715 82.255 206.760 ;
        RECT 83.790 206.700 84.110 206.960 ;
        RECT 93.910 206.900 94.230 206.960 ;
        RECT 89.860 206.760 94.230 206.900 ;
        RECT 71.370 206.560 71.690 206.620 ;
        RECT 46.990 206.420 60.560 206.560 ;
        RECT 61.340 206.420 71.690 206.560 ;
        RECT 46.990 206.360 47.310 206.420 ;
        RECT 51.145 206.375 51.435 206.420 ;
        RECT 16.630 206.020 16.950 206.280 ;
        RECT 17.565 206.220 17.855 206.265 ;
        RECT 25.370 206.220 25.690 206.280 ;
        RECT 35.490 206.220 35.810 206.280 ;
        RECT 35.965 206.220 36.255 206.265 ;
        RECT 17.565 206.080 20.540 206.220 ;
        RECT 17.565 206.035 17.855 206.080 ;
        RECT 20.400 205.585 20.540 206.080 ;
        RECT 25.370 206.080 32.500 206.220 ;
        RECT 25.370 206.020 25.690 206.080 ;
        RECT 26.290 205.880 26.610 205.940 ;
        RECT 31.810 205.880 32.130 205.940 ;
        RECT 26.290 205.740 32.130 205.880 ;
        RECT 32.360 205.880 32.500 206.080 ;
        RECT 35.490 206.080 36.255 206.220 ;
        RECT 35.490 206.020 35.810 206.080 ;
        RECT 35.965 206.035 36.255 206.080 ;
        RECT 37.330 206.020 37.650 206.280 ;
        RECT 47.450 206.220 47.770 206.280 ;
        RECT 47.920 206.220 48.210 206.265 ;
        RECT 47.450 206.080 48.210 206.220 ;
        RECT 47.450 206.020 47.770 206.080 ;
        RECT 47.920 206.035 48.210 206.080 ;
        RECT 48.370 206.020 48.690 206.280 ;
        RECT 48.845 206.035 49.135 206.265 ;
        RECT 43.310 205.880 43.630 205.940 ;
        RECT 32.360 205.740 43.630 205.880 ;
        RECT 26.290 205.680 26.610 205.740 ;
        RECT 31.810 205.680 32.130 205.740 ;
        RECT 43.310 205.680 43.630 205.740 ;
        RECT 45.625 205.880 45.915 205.925 ;
        RECT 48.920 205.880 49.060 206.035 ;
        RECT 49.750 206.020 50.070 206.280 ;
        RECT 50.670 206.220 50.990 206.280 ;
        RECT 52.065 206.220 52.355 206.265 ;
        RECT 50.670 206.080 52.355 206.220 ;
        RECT 50.670 206.020 50.990 206.080 ;
        RECT 52.065 206.035 52.355 206.080 ;
        RECT 54.810 206.020 55.130 206.280 ;
        RECT 55.730 206.020 56.050 206.280 ;
        RECT 56.190 206.220 56.510 206.280 ;
        RECT 57.585 206.220 57.875 206.265 ;
        RECT 56.190 206.080 57.875 206.220 ;
        RECT 56.190 206.020 56.510 206.080 ;
        RECT 57.585 206.035 57.875 206.080 ;
        RECT 58.950 206.220 59.270 206.280 ;
        RECT 61.340 206.265 61.480 206.420 ;
        RECT 71.370 206.360 71.690 206.420 ;
        RECT 73.605 206.560 73.895 206.605 ;
        RECT 73.605 206.420 74.360 206.560 ;
        RECT 73.605 206.375 73.895 206.420 ;
        RECT 60.345 206.220 60.635 206.265 ;
        RECT 58.950 206.080 60.635 206.220 ;
        RECT 58.950 206.020 59.270 206.080 ;
        RECT 60.345 206.035 60.635 206.080 ;
        RECT 61.265 206.035 61.555 206.265 ;
        RECT 61.725 206.220 62.015 206.265 ;
        RECT 64.470 206.220 64.790 206.280 ;
        RECT 61.725 206.080 64.790 206.220 ;
        RECT 61.725 206.035 62.015 206.080 ;
        RECT 57.110 205.880 57.430 205.940 ;
        RECT 45.625 205.740 57.430 205.880 ;
        RECT 45.625 205.695 45.915 205.740 ;
        RECT 57.110 205.680 57.430 205.740 ;
        RECT 59.425 205.695 59.715 205.925 ;
        RECT 20.325 205.540 20.615 205.585 ;
        RECT 46.070 205.540 46.390 205.600 ;
        RECT 20.325 205.400 46.390 205.540 ;
        RECT 20.325 205.355 20.615 205.400 ;
        RECT 46.070 205.340 46.390 205.400 ;
        RECT 46.545 205.540 46.835 205.585 ;
        RECT 49.750 205.540 50.070 205.600 ;
        RECT 46.545 205.400 50.070 205.540 ;
        RECT 46.545 205.355 46.835 205.400 ;
        RECT 49.750 205.340 50.070 205.400 ;
        RECT 54.350 205.540 54.670 205.600 ;
        RECT 56.190 205.540 56.510 205.600 ;
        RECT 54.350 205.400 56.510 205.540 ;
        RECT 54.350 205.340 54.670 205.400 ;
        RECT 56.190 205.340 56.510 205.400 ;
        RECT 56.665 205.540 56.955 205.585 ;
        RECT 58.030 205.540 58.350 205.600 ;
        RECT 56.665 205.400 58.350 205.540 ;
        RECT 56.665 205.355 56.955 205.400 ;
        RECT 58.030 205.340 58.350 205.400 ;
        RECT 58.965 205.355 59.255 205.585 ;
        RECT 23.070 205.200 23.390 205.260 ;
        RECT 27.670 205.200 27.990 205.260 ;
        RECT 23.070 205.060 27.990 205.200 ;
        RECT 23.070 205.000 23.390 205.060 ;
        RECT 27.670 205.000 27.990 205.060 ;
        RECT 29.525 205.200 29.815 205.245 ;
        RECT 31.350 205.200 31.670 205.260 ;
        RECT 29.525 205.060 31.670 205.200 ;
        RECT 29.525 205.015 29.815 205.060 ;
        RECT 31.350 205.000 31.670 205.060 ;
        RECT 31.810 205.200 32.130 205.260 ;
        RECT 59.040 205.200 59.180 205.355 ;
        RECT 31.810 205.060 59.180 205.200 ;
        RECT 59.500 205.200 59.640 205.695 ;
        RECT 60.420 205.540 60.560 206.035 ;
        RECT 64.470 206.020 64.790 206.080 ;
        RECT 65.865 206.220 66.155 206.265 ;
        RECT 67.230 206.220 67.550 206.280 ;
        RECT 65.865 206.080 67.550 206.220 ;
        RECT 65.865 206.035 66.155 206.080 ;
        RECT 67.230 206.020 67.550 206.080 ;
        RECT 67.705 206.035 67.995 206.265 ;
        RECT 69.085 206.035 69.375 206.265 ;
        RECT 69.530 206.220 69.850 206.280 ;
        RECT 70.005 206.220 70.295 206.265 ;
        RECT 70.450 206.220 70.770 206.280 ;
        RECT 69.530 206.080 70.770 206.220 ;
        RECT 64.930 205.680 65.250 205.940 ;
        RECT 65.405 205.880 65.695 205.925 ;
        RECT 66.770 205.880 67.090 205.940 ;
        RECT 65.405 205.740 67.090 205.880 ;
        RECT 65.405 205.695 65.695 205.740 ;
        RECT 66.770 205.680 67.090 205.740 ;
        RECT 67.780 205.540 67.920 206.035 ;
        RECT 69.160 205.880 69.300 206.035 ;
        RECT 69.530 206.020 69.850 206.080 ;
        RECT 70.005 206.035 70.295 206.080 ;
        RECT 70.450 206.020 70.770 206.080 ;
        RECT 70.910 206.220 71.230 206.280 ;
        RECT 71.845 206.220 72.135 206.265 ;
        RECT 70.910 206.080 72.135 206.220 ;
        RECT 70.910 206.020 71.230 206.080 ;
        RECT 71.845 206.035 72.135 206.080 ;
        RECT 72.305 206.220 72.595 206.265 ;
        RECT 72.750 206.220 73.070 206.280 ;
        RECT 72.305 206.080 73.070 206.220 ;
        RECT 74.220 206.220 74.360 206.420 ;
        RECT 74.590 206.360 74.910 206.620 ;
        RECT 79.045 206.560 79.335 206.605 ;
        RECT 76.060 206.420 79.335 206.560 ;
        RECT 76.060 206.280 76.200 206.420 ;
        RECT 79.045 206.375 79.335 206.420 ;
        RECT 80.110 206.360 80.430 206.620 ;
        RECT 83.880 206.560 84.020 206.700 ;
        RECT 89.860 206.560 90.000 206.760 ;
        RECT 93.910 206.700 94.230 206.760 ;
        RECT 94.385 206.900 94.675 206.945 ;
        RECT 94.830 206.900 95.150 206.960 ;
        RECT 96.225 206.900 96.515 206.945 ;
        RECT 94.385 206.760 96.515 206.900 ;
        RECT 94.385 206.715 94.675 206.760 ;
        RECT 94.830 206.700 95.150 206.760 ;
        RECT 96.225 206.715 96.515 206.760 ;
        RECT 82.040 206.420 84.020 206.560 ;
        RECT 85.720 206.420 90.000 206.560 ;
        RECT 75.970 206.220 76.290 206.280 ;
        RECT 74.220 206.080 76.290 206.220 ;
        RECT 72.305 206.035 72.595 206.080 ;
        RECT 72.750 206.020 73.070 206.080 ;
        RECT 75.970 206.020 76.290 206.080 ;
        RECT 76.430 206.020 76.750 206.280 ;
        RECT 76.890 206.220 77.210 206.280 ;
        RECT 77.825 206.220 78.115 206.265 ;
        RECT 81.505 206.220 81.795 206.265 ;
        RECT 82.040 206.220 82.180 206.420 ;
        RECT 76.890 206.080 79.880 206.220 ;
        RECT 76.890 206.020 77.210 206.080 ;
        RECT 77.825 206.035 78.115 206.080 ;
        RECT 69.160 205.740 72.980 205.880 ;
        RECT 69.160 205.540 69.300 205.740 ;
        RECT 72.840 205.585 72.980 205.740 ;
        RECT 73.670 205.680 73.990 205.940 ;
        RECT 74.130 205.880 74.450 205.940 ;
        RECT 77.365 205.880 77.655 205.925 ;
        RECT 74.130 205.740 79.420 205.880 ;
        RECT 74.130 205.680 74.450 205.740 ;
        RECT 77.365 205.695 77.655 205.740 ;
        RECT 60.420 205.400 67.920 205.540 ;
        RECT 68.240 205.400 69.300 205.540 ;
        RECT 66.860 205.260 67.000 205.400 ;
        RECT 63.090 205.200 63.410 205.260 ;
        RECT 59.500 205.060 63.410 205.200 ;
        RECT 31.810 205.000 32.130 205.060 ;
        RECT 63.090 205.000 63.410 205.060 ;
        RECT 63.565 205.200 63.855 205.245 ;
        RECT 64.470 205.200 64.790 205.260 ;
        RECT 63.565 205.060 64.790 205.200 ;
        RECT 63.565 205.015 63.855 205.060 ;
        RECT 64.470 205.000 64.790 205.060 ;
        RECT 66.770 205.000 67.090 205.260 ;
        RECT 67.230 205.200 67.550 205.260 ;
        RECT 68.240 205.200 68.380 205.400 ;
        RECT 72.765 205.355 73.055 205.585 ;
        RECT 73.760 205.540 73.900 205.680 ;
        RECT 78.285 205.540 78.575 205.585 ;
        RECT 73.300 205.400 78.575 205.540 ;
        RECT 67.230 205.060 68.380 205.200 ;
        RECT 69.070 205.200 69.390 205.260 ;
        RECT 70.465 205.200 70.755 205.245 ;
        RECT 69.070 205.060 70.755 205.200 ;
        RECT 67.230 205.000 67.550 205.060 ;
        RECT 69.070 205.000 69.390 205.060 ;
        RECT 70.465 205.015 70.755 205.060 ;
        RECT 72.305 205.200 72.595 205.245 ;
        RECT 73.300 205.200 73.440 205.400 ;
        RECT 78.285 205.355 78.575 205.400 ;
        RECT 72.305 205.060 73.440 205.200 ;
        RECT 73.685 205.200 73.975 205.245 ;
        RECT 74.130 205.200 74.450 205.260 ;
        RECT 73.685 205.060 74.450 205.200 ;
        RECT 72.305 205.015 72.595 205.060 ;
        RECT 73.685 205.015 73.975 205.060 ;
        RECT 74.130 205.000 74.450 205.060 ;
        RECT 75.050 205.000 75.370 205.260 ;
        RECT 76.430 205.200 76.750 205.260 ;
        RECT 77.810 205.200 78.130 205.260 ;
        RECT 79.280 205.245 79.420 205.740 ;
        RECT 79.740 205.540 79.880 206.080 ;
        RECT 81.505 206.080 82.180 206.220 ;
        RECT 81.505 206.035 81.795 206.080 ;
        RECT 82.870 206.020 83.190 206.280 ;
        RECT 84.265 206.220 84.555 206.265 ;
        RECT 85.170 206.220 85.490 206.280 ;
        RECT 85.720 206.265 85.860 206.420 ;
        RECT 84.265 206.080 85.490 206.220 ;
        RECT 84.265 206.035 84.555 206.080 ;
        RECT 85.170 206.020 85.490 206.080 ;
        RECT 85.645 206.035 85.935 206.265 ;
        RECT 86.090 206.020 86.410 206.280 ;
        RECT 87.470 206.220 87.790 206.280 ;
        RECT 88.850 206.220 89.170 206.280 ;
        RECT 89.400 206.265 89.540 206.420 ;
        RECT 87.470 206.080 89.170 206.220 ;
        RECT 87.470 206.020 87.790 206.080 ;
        RECT 88.850 206.020 89.170 206.080 ;
        RECT 89.325 206.035 89.615 206.265 ;
        RECT 89.770 206.020 90.090 206.280 ;
        RECT 91.165 206.035 91.455 206.265 ;
        RECT 91.610 206.220 91.930 206.280 ;
        RECT 93.465 206.220 93.755 206.265 ;
        RECT 91.610 206.080 93.755 206.220 ;
        RECT 94.000 206.220 94.140 206.700 ;
        RECT 95.290 206.360 95.610 206.620 ;
        RECT 94.845 206.220 95.135 206.265 ;
        RECT 96.685 206.220 96.975 206.265 ;
        RECT 94.000 206.080 96.975 206.220 ;
        RECT 80.570 205.880 80.890 205.940 ;
        RECT 84.725 205.880 85.015 205.925 ;
        RECT 80.570 205.740 85.015 205.880 ;
        RECT 85.260 205.880 85.400 206.020 ;
        RECT 87.025 205.880 87.315 205.925 ;
        RECT 90.705 205.880 90.995 205.925 ;
        RECT 85.260 205.740 90.995 205.880 ;
        RECT 91.240 205.880 91.380 206.035 ;
        RECT 91.610 206.020 91.930 206.080 ;
        RECT 93.465 206.035 93.755 206.080 ;
        RECT 94.845 206.035 95.135 206.080 ;
        RECT 96.685 206.035 96.975 206.080 ;
        RECT 93.540 205.880 93.680 206.035 ;
        RECT 95.290 205.880 95.610 205.940 ;
        RECT 91.240 205.740 93.220 205.880 ;
        RECT 93.540 205.740 95.610 205.880 ;
        RECT 80.570 205.680 80.890 205.740 ;
        RECT 84.725 205.695 85.015 205.740 ;
        RECT 87.025 205.695 87.315 205.740 ;
        RECT 90.705 205.695 90.995 205.740 ;
        RECT 92.545 205.540 92.835 205.585 ;
        RECT 79.740 205.400 92.835 205.540 ;
        RECT 93.080 205.540 93.220 205.740 ;
        RECT 95.290 205.680 95.610 205.740 ;
        RECT 96.210 205.540 96.530 205.600 ;
        RECT 93.080 205.400 96.530 205.540 ;
        RECT 92.545 205.355 92.835 205.400 ;
        RECT 96.210 205.340 96.530 205.400 ;
        RECT 76.430 205.060 78.130 205.200 ;
        RECT 76.430 205.000 76.750 205.060 ;
        RECT 77.810 205.000 78.130 205.060 ;
        RECT 79.205 205.015 79.495 205.245 ;
        RECT 81.030 205.000 81.350 205.260 ;
        RECT 81.950 205.200 82.270 205.260 ;
        RECT 88.405 205.200 88.695 205.245 ;
        RECT 81.950 205.060 88.695 205.200 ;
        RECT 81.950 205.000 82.270 205.060 ;
        RECT 88.405 205.015 88.695 205.060 ;
        RECT 92.070 205.200 92.390 205.260 ;
        RECT 95.305 205.200 95.595 205.245 ;
        RECT 92.070 205.060 95.595 205.200 ;
        RECT 92.070 205.000 92.390 205.060 ;
        RECT 95.305 205.015 95.595 205.060 ;
        RECT 14.260 204.380 126.960 204.860 ;
        RECT 25.920 204.040 30.200 204.180 ;
        RECT 20.770 203.640 21.090 203.900 ;
        RECT 24.465 203.840 24.755 203.885 ;
        RECT 22.010 203.700 24.755 203.840 ;
        RECT 16.185 203.500 16.475 203.545 ;
        RECT 21.230 203.500 21.550 203.560 ;
        RECT 16.185 203.360 21.550 203.500 ;
        RECT 16.185 203.315 16.475 203.360 ;
        RECT 21.230 203.300 21.550 203.360 ;
        RECT 16.645 202.975 16.935 203.205 ;
        RECT 16.720 202.820 16.860 202.975 ;
        RECT 18.010 202.960 18.330 203.220 ;
        RECT 18.930 202.960 19.250 203.220 ;
        RECT 19.865 203.160 20.155 203.205 ;
        RECT 22.010 203.160 22.150 203.700 ;
        RECT 24.465 203.655 24.755 203.700 ;
        RECT 25.370 203.205 25.690 203.220 ;
        RECT 25.920 203.205 26.060 204.040 ;
        RECT 29.510 203.840 29.830 203.900 ;
        RECT 27.760 203.700 29.830 203.840 ;
        RECT 27.760 203.500 27.900 203.700 ;
        RECT 29.510 203.640 29.830 203.700 ;
        RECT 27.300 203.360 27.900 203.500 ;
        RECT 25.360 203.160 25.690 203.205 ;
        RECT 19.865 203.020 22.150 203.160 ;
        RECT 25.175 203.020 25.690 203.160 ;
        RECT 19.865 202.975 20.155 203.020 ;
        RECT 25.360 202.975 25.690 203.020 ;
        RECT 25.845 202.975 26.135 203.205 ;
        RECT 25.370 202.960 25.690 202.975 ;
        RECT 26.290 202.960 26.610 203.220 ;
        RECT 27.300 203.205 27.440 203.360 ;
        RECT 28.130 203.300 28.450 203.560 ;
        RECT 28.605 203.500 28.895 203.545 ;
        RECT 29.050 203.500 29.370 203.560 ;
        RECT 28.605 203.360 29.370 203.500 ;
        RECT 30.060 203.500 30.200 204.040 ;
        RECT 30.890 203.980 31.210 204.240 ;
        RECT 51.590 204.180 51.910 204.240 ;
        RECT 52.510 204.180 52.830 204.240 ;
        RECT 58.950 204.180 59.270 204.240 ;
        RECT 51.590 204.040 59.270 204.180 ;
        RECT 51.590 203.980 51.910 204.040 ;
        RECT 52.510 203.980 52.830 204.040 ;
        RECT 34.110 203.640 34.430 203.900 ;
        RECT 55.270 203.840 55.590 203.900 ;
        RECT 42.020 203.700 55.590 203.840 ;
        RECT 39.630 203.500 39.950 203.560 ;
        RECT 30.060 203.360 39.950 203.500 ;
        RECT 28.605 203.315 28.895 203.360 ;
        RECT 29.050 203.300 29.370 203.360 ;
        RECT 39.630 203.300 39.950 203.360 ;
        RECT 40.090 203.500 40.410 203.560 ;
        RECT 42.020 203.545 42.160 203.700 ;
        RECT 55.270 203.640 55.590 203.700 ;
        RECT 55.730 203.640 56.050 203.900 ;
        RECT 41.485 203.500 41.775 203.545 ;
        RECT 40.090 203.360 41.775 203.500 ;
        RECT 40.090 203.300 40.410 203.360 ;
        RECT 41.485 203.315 41.775 203.360 ;
        RECT 41.945 203.315 42.235 203.545 ;
        RECT 45.165 203.500 45.455 203.545 ;
        RECT 42.940 203.360 45.455 203.500 ;
        RECT 27.225 202.975 27.515 203.205 ;
        RECT 27.685 202.975 27.975 203.205 ;
        RECT 28.220 203.160 28.360 203.300 ;
        RECT 29.525 203.160 29.815 203.205 ;
        RECT 28.220 203.020 29.815 203.160 ;
        RECT 29.525 202.975 29.815 203.020 ;
        RECT 29.985 203.160 30.275 203.205 ;
        RECT 36.410 203.160 36.730 203.220 ;
        RECT 29.985 203.020 36.730 203.160 ;
        RECT 29.985 202.975 30.275 203.020 ;
        RECT 20.310 202.820 20.630 202.880 ;
        RECT 16.720 202.680 20.630 202.820 ;
        RECT 20.310 202.620 20.630 202.680 ;
        RECT 20.770 202.820 21.090 202.880 ;
        RECT 27.760 202.820 27.900 202.975 ;
        RECT 36.410 202.960 36.730 203.020 ;
        RECT 40.565 203.160 40.855 203.205 ;
        RECT 42.940 203.160 43.080 203.360 ;
        RECT 45.165 203.315 45.455 203.360 ;
        RECT 46.530 203.500 46.850 203.560 ;
        RECT 50.210 203.500 50.530 203.560 ;
        RECT 50.685 203.500 50.975 203.545 ;
        RECT 46.530 203.360 49.980 203.500 ;
        RECT 46.530 203.300 46.850 203.360 ;
        RECT 40.565 203.020 43.080 203.160 ;
        RECT 43.325 203.160 43.615 203.205 ;
        RECT 45.610 203.160 45.930 203.220 ;
        RECT 43.325 203.020 45.930 203.160 ;
        RECT 40.565 202.975 40.855 203.020 ;
        RECT 43.325 202.975 43.615 203.020 ;
        RECT 45.610 202.960 45.930 203.020 ;
        RECT 46.070 203.160 46.390 203.220 ;
        RECT 48.370 203.160 48.690 203.220 ;
        RECT 49.840 203.205 49.980 203.360 ;
        RECT 50.210 203.360 50.975 203.500 ;
        RECT 50.210 203.300 50.530 203.360 ;
        RECT 50.685 203.315 50.975 203.360 ;
        RECT 51.130 203.300 51.450 203.560 ;
        RECT 52.050 203.300 52.370 203.560 ;
        RECT 53.905 203.500 54.195 203.545 ;
        RECT 54.350 203.500 54.670 203.560 ;
        RECT 53.905 203.360 54.670 203.500 ;
        RECT 53.905 203.315 54.195 203.360 ;
        RECT 54.350 203.300 54.670 203.360 ;
        RECT 54.810 203.500 55.130 203.560 ;
        RECT 55.820 203.500 55.960 203.640 ;
        RECT 57.660 203.545 57.800 204.040 ;
        RECT 58.950 203.980 59.270 204.040 ;
        RECT 59.870 203.980 60.190 204.240 ;
        RECT 66.785 204.180 67.075 204.225 ;
        RECT 69.530 204.180 69.850 204.240 ;
        RECT 66.785 204.040 69.850 204.180 ;
        RECT 66.785 203.995 67.075 204.040 ;
        RECT 69.530 203.980 69.850 204.040 ;
        RECT 70.465 204.180 70.755 204.225 ;
        RECT 70.910 204.180 71.230 204.240 ;
        RECT 70.465 204.040 71.230 204.180 ;
        RECT 70.465 203.995 70.755 204.040 ;
        RECT 70.910 203.980 71.230 204.040 ;
        RECT 71.385 204.180 71.675 204.225 ;
        RECT 72.290 204.180 72.610 204.240 ;
        RECT 73.685 204.180 73.975 204.225 ;
        RECT 75.050 204.180 75.370 204.240 ;
        RECT 71.385 204.040 73.975 204.180 ;
        RECT 71.385 203.995 71.675 204.040 ;
        RECT 72.290 203.980 72.610 204.040 ;
        RECT 73.685 203.995 73.975 204.040 ;
        RECT 74.220 204.040 75.370 204.180 ;
        RECT 60.345 203.840 60.635 203.885 ;
        RECT 66.310 203.840 66.630 203.900 ;
        RECT 58.120 203.700 66.630 203.840 ;
        RECT 54.810 203.360 55.960 203.500 ;
        RECT 54.810 203.300 55.130 203.360 ;
        RECT 57.585 203.315 57.875 203.545 ;
        RECT 48.845 203.160 49.135 203.205 ;
        RECT 46.070 203.020 49.135 203.160 ;
        RECT 46.070 202.960 46.390 203.020 ;
        RECT 48.370 202.960 48.690 203.020 ;
        RECT 48.845 202.975 49.135 203.020 ;
        RECT 49.765 202.975 50.055 203.205 ;
        RECT 51.605 202.975 51.895 203.205 ;
        RECT 20.770 202.680 27.900 202.820 ;
        RECT 20.770 202.620 21.090 202.680 ;
        RECT 28.145 202.635 28.435 202.865 ;
        RECT 33.650 202.820 33.970 202.880 ;
        RECT 51.130 202.820 51.450 202.880 ;
        RECT 33.650 202.680 51.450 202.820 ;
        RECT 51.680 202.820 51.820 202.975 ;
        RECT 52.970 202.960 53.290 203.220 ;
        RECT 54.440 203.160 54.580 203.300 ;
        RECT 58.120 203.160 58.260 203.700 ;
        RECT 60.345 203.655 60.635 203.700 ;
        RECT 66.310 203.640 66.630 203.700 ;
        RECT 67.230 203.640 67.550 203.900 ;
        RECT 69.070 203.840 69.390 203.900 ;
        RECT 67.780 203.700 69.390 203.840 ;
        RECT 67.780 203.500 67.920 203.700 ;
        RECT 69.070 203.640 69.390 203.700 ;
        RECT 72.750 203.640 73.070 203.900 ;
        RECT 74.220 203.840 74.360 204.040 ;
        RECT 75.050 203.980 75.370 204.040 ;
        RECT 75.510 203.980 75.830 204.240 ;
        RECT 77.825 204.180 78.115 204.225 ;
        RECT 80.110 204.180 80.430 204.240 ;
        RECT 87.010 204.180 87.330 204.240 ;
        RECT 77.825 204.040 86.780 204.180 ;
        RECT 77.825 203.995 78.115 204.040 ;
        RECT 80.110 203.980 80.430 204.040 ;
        RECT 73.300 203.700 74.360 203.840 ;
        RECT 74.590 203.840 74.910 203.900 ;
        RECT 85.630 203.840 85.950 203.900 ;
        RECT 86.640 203.885 86.780 204.040 ;
        RECT 87.010 204.040 106.100 204.180 ;
        RECT 87.010 203.980 87.330 204.040 ;
        RECT 74.590 203.700 85.950 203.840 ;
        RECT 70.910 203.500 71.230 203.560 ;
        RECT 73.300 203.500 73.440 203.700 ;
        RECT 74.590 203.640 74.910 203.700 ;
        RECT 75.510 203.500 75.830 203.560 ;
        RECT 65.940 203.360 67.920 203.500 ;
        RECT 68.700 203.360 73.440 203.500 ;
        RECT 73.680 203.360 75.830 203.500 ;
        RECT 54.440 203.020 58.260 203.160 ;
        RECT 58.965 203.160 59.255 203.205 ;
        RECT 59.870 203.160 60.190 203.220 ;
        RECT 61.250 203.160 61.570 203.220 ;
        RECT 58.965 203.020 61.570 203.160 ;
        RECT 58.965 202.975 59.255 203.020 ;
        RECT 59.870 202.960 60.190 203.020 ;
        RECT 61.250 202.960 61.570 203.020 ;
        RECT 62.185 203.160 62.475 203.205 ;
        RECT 63.090 203.160 63.410 203.220 ;
        RECT 62.185 203.020 63.410 203.160 ;
        RECT 62.185 202.975 62.475 203.020 ;
        RECT 63.090 202.960 63.410 203.020 ;
        RECT 64.010 202.960 64.330 203.220 ;
        RECT 64.470 202.960 64.790 203.220 ;
        RECT 64.930 203.160 65.250 203.220 ;
        RECT 65.940 203.205 66.080 203.360 ;
        RECT 68.700 203.205 68.840 203.360 ;
        RECT 70.910 203.300 71.230 203.360 ;
        RECT 65.405 203.160 65.695 203.205 ;
        RECT 64.930 203.020 65.695 203.160 ;
        RECT 64.930 202.960 65.250 203.020 ;
        RECT 65.405 202.975 65.695 203.020 ;
        RECT 65.865 202.975 66.155 203.205 ;
        RECT 68.625 202.975 68.915 203.205 ;
        RECT 73.680 203.160 73.820 203.360 ;
        RECT 75.510 203.300 75.830 203.360 ;
        RECT 76.520 203.205 76.660 203.700 ;
        RECT 85.630 203.640 85.950 203.700 ;
        RECT 86.565 203.655 86.855 203.885 ;
        RECT 89.310 203.840 89.630 203.900 ;
        RECT 90.690 203.840 91.010 203.900 ;
        RECT 92.545 203.840 92.835 203.885 ;
        RECT 89.310 203.700 90.460 203.840 ;
        RECT 86.640 203.500 86.780 203.655 ;
        RECT 89.310 203.640 89.630 203.700 ;
        RECT 83.880 203.360 85.860 203.500 ;
        RECT 86.640 203.360 89.540 203.500 ;
        RECT 83.880 203.220 84.020 203.360 ;
        RECT 69.995 203.020 73.820 203.160 ;
        RECT 53.890 202.820 54.210 202.880 ;
        RECT 58.045 202.820 58.335 202.865 ;
        RECT 67.245 202.820 67.535 202.865 ;
        RECT 51.680 202.680 67.535 202.820 ;
        RECT 25.370 202.480 25.690 202.540 ;
        RECT 28.220 202.480 28.360 202.635 ;
        RECT 33.650 202.620 33.970 202.680 ;
        RECT 51.130 202.620 51.450 202.680 ;
        RECT 53.890 202.620 54.210 202.680 ;
        RECT 58.045 202.635 58.335 202.680 ;
        RECT 67.245 202.635 67.535 202.680 ;
        RECT 25.370 202.340 28.360 202.480 ;
        RECT 46.990 202.480 47.310 202.540 ;
        RECT 55.730 202.480 56.050 202.540 ;
        RECT 56.205 202.480 56.495 202.525 ;
        RECT 46.990 202.340 56.495 202.480 ;
        RECT 25.370 202.280 25.690 202.340 ;
        RECT 46.990 202.280 47.310 202.340 ;
        RECT 55.730 202.280 56.050 202.340 ;
        RECT 56.205 202.295 56.495 202.340 ;
        RECT 57.110 202.480 57.430 202.540 ;
        RECT 61.250 202.480 61.570 202.540 ;
        RECT 57.110 202.340 61.570 202.480 ;
        RECT 57.110 202.280 57.430 202.340 ;
        RECT 61.250 202.280 61.570 202.340 ;
        RECT 65.850 202.480 66.170 202.540 ;
        RECT 68.165 202.480 68.455 202.525 ;
        RECT 69.995 202.480 70.135 203.020 ;
        RECT 76.445 202.975 76.735 203.205 ;
        RECT 76.905 202.975 77.195 203.205 ;
        RECT 72.305 202.820 72.595 202.865 ;
        RECT 74.590 202.820 74.910 202.880 ;
        RECT 72.305 202.680 74.910 202.820 ;
        RECT 72.305 202.635 72.595 202.680 ;
        RECT 74.590 202.620 74.910 202.680 ;
        RECT 75.510 202.820 75.830 202.880 ;
        RECT 76.980 202.820 77.120 202.975 ;
        RECT 83.790 202.960 84.110 203.220 ;
        RECT 84.725 203.160 85.015 203.205 ;
        RECT 85.170 203.160 85.490 203.220 ;
        RECT 85.720 203.205 85.860 203.360 ;
        RECT 84.725 203.020 85.490 203.160 ;
        RECT 84.725 202.975 85.015 203.020 ;
        RECT 85.170 202.960 85.490 203.020 ;
        RECT 85.645 202.975 85.935 203.205 ;
        RECT 86.090 203.160 86.410 203.220 ;
        RECT 86.565 203.160 86.855 203.205 ;
        RECT 88.390 203.160 88.710 203.220 ;
        RECT 89.400 203.205 89.540 203.360 ;
        RECT 86.090 203.020 88.710 203.160 ;
        RECT 86.090 202.960 86.410 203.020 ;
        RECT 86.565 202.975 86.855 203.020 ;
        RECT 88.390 202.960 88.710 203.020 ;
        RECT 89.325 202.975 89.615 203.205 ;
        RECT 89.770 202.960 90.090 203.220 ;
        RECT 90.320 203.160 90.460 203.700 ;
        RECT 90.690 203.700 92.835 203.840 ;
        RECT 90.690 203.640 91.010 203.700 ;
        RECT 92.545 203.655 92.835 203.700 ;
        RECT 93.925 203.500 94.215 203.545 ;
        RECT 91.700 203.360 94.215 203.500 ;
        RECT 90.705 203.160 90.995 203.205 ;
        RECT 90.320 203.020 90.995 203.160 ;
        RECT 90.705 202.975 90.995 203.020 ;
        RECT 91.150 202.960 91.470 203.220 ;
        RECT 91.700 203.205 91.840 203.360 ;
        RECT 93.925 203.315 94.215 203.360 ;
        RECT 105.960 203.220 106.100 204.040 ;
        RECT 91.625 202.975 91.915 203.205 ;
        RECT 75.510 202.680 77.120 202.820 ;
        RECT 75.510 202.620 75.830 202.680 ;
        RECT 77.810 202.620 78.130 202.880 ;
        RECT 84.265 202.820 84.555 202.865 ;
        RECT 87.010 202.820 87.330 202.880 ;
        RECT 84.265 202.680 87.330 202.820 ;
        RECT 84.265 202.635 84.555 202.680 ;
        RECT 87.010 202.620 87.330 202.680 ;
        RECT 87.945 202.820 88.235 202.865 ;
        RECT 91.700 202.820 91.840 202.975 ;
        RECT 93.450 202.960 93.770 203.220 ;
        RECT 94.385 203.160 94.675 203.205 ;
        RECT 94.830 203.160 95.150 203.220 ;
        RECT 94.385 203.020 95.150 203.160 ;
        RECT 94.385 202.975 94.675 203.020 ;
        RECT 94.830 202.960 95.150 203.020 ;
        RECT 105.425 202.975 105.715 203.205 ;
        RECT 105.870 203.160 106.190 203.220 ;
        RECT 106.345 203.160 106.635 203.205 ;
        RECT 111.850 203.160 112.170 203.220 ;
        RECT 105.870 203.020 112.170 203.160 ;
        RECT 87.945 202.680 91.840 202.820 ;
        RECT 87.945 202.635 88.235 202.680 ;
        RECT 104.030 202.620 104.350 202.880 ;
        RECT 105.500 202.820 105.640 202.975 ;
        RECT 105.870 202.960 106.190 203.020 ;
        RECT 106.345 202.975 106.635 203.020 ;
        RECT 111.850 202.960 112.170 203.020 ;
        RECT 108.630 202.820 108.950 202.880 ;
        RECT 104.580 202.680 108.950 202.820 ;
        RECT 65.850 202.340 70.135 202.480 ;
        RECT 71.305 202.480 71.595 202.525 ;
        RECT 71.830 202.480 72.150 202.540 ;
        RECT 71.305 202.340 72.150 202.480 ;
        RECT 65.850 202.280 66.170 202.340 ;
        RECT 68.165 202.295 68.455 202.340 ;
        RECT 71.305 202.295 71.595 202.340 ;
        RECT 71.830 202.280 72.150 202.340 ;
        RECT 73.605 202.480 73.895 202.525 ;
        RECT 77.900 202.480 78.040 202.620 ;
        RECT 73.605 202.340 78.040 202.480 ;
        RECT 88.865 202.480 89.155 202.525 ;
        RECT 90.230 202.480 90.550 202.540 ;
        RECT 93.450 202.480 93.770 202.540 ;
        RECT 88.865 202.340 93.770 202.480 ;
        RECT 73.605 202.295 73.895 202.340 ;
        RECT 88.865 202.295 89.155 202.340 ;
        RECT 90.230 202.280 90.550 202.340 ;
        RECT 93.450 202.280 93.770 202.340 ;
        RECT 99.890 202.480 100.210 202.540 ;
        RECT 104.580 202.525 104.720 202.680 ;
        RECT 108.630 202.620 108.950 202.680 ;
        RECT 109.090 202.820 109.410 202.880 ;
        RECT 110.945 202.820 111.235 202.865 ;
        RECT 109.090 202.680 111.235 202.820 ;
        RECT 109.090 202.620 109.410 202.680 ;
        RECT 110.945 202.635 111.235 202.680 ;
        RECT 104.505 202.480 104.795 202.525 ;
        RECT 99.890 202.340 104.795 202.480 ;
        RECT 99.890 202.280 100.210 202.340 ;
        RECT 104.505 202.295 104.795 202.340 ;
        RECT 107.265 202.480 107.555 202.525 ;
        RECT 108.170 202.480 108.490 202.540 ;
        RECT 107.265 202.340 108.490 202.480 ;
        RECT 107.265 202.295 107.555 202.340 ;
        RECT 108.170 202.280 108.490 202.340 ;
        RECT 14.260 201.660 126.960 202.140 ;
        RECT 16.170 201.260 16.490 201.520 ;
        RECT 44.690 201.460 45.010 201.520 ;
        RECT 46.530 201.460 46.850 201.520 ;
        RECT 49.305 201.460 49.595 201.505 ;
        RECT 50.670 201.460 50.990 201.520 ;
        RECT 58.030 201.460 58.350 201.520 ;
        RECT 44.690 201.320 50.990 201.460 ;
        RECT 44.690 201.260 45.010 201.320 ;
        RECT 46.530 201.260 46.850 201.320 ;
        RECT 49.305 201.275 49.595 201.320 ;
        RECT 50.670 201.260 50.990 201.320 ;
        RECT 55.820 201.320 58.350 201.460 ;
        RECT 35.950 200.920 36.270 201.180 ;
        RECT 48.370 201.120 48.690 201.180 ;
        RECT 53.445 201.120 53.735 201.165 ;
        RECT 48.370 200.980 53.735 201.120 ;
        RECT 48.370 200.920 48.690 200.980 ;
        RECT 53.445 200.935 53.735 200.980 ;
        RECT 16.630 200.780 16.950 200.840 ;
        RECT 17.105 200.780 17.395 200.825 ;
        RECT 16.630 200.640 17.395 200.780 ;
        RECT 16.630 200.580 16.950 200.640 ;
        RECT 17.105 200.595 17.395 200.640 ;
        RECT 18.025 200.780 18.315 200.825 ;
        RECT 19.390 200.780 19.710 200.840 ;
        RECT 18.025 200.640 19.710 200.780 ;
        RECT 18.025 200.595 18.315 200.640 ;
        RECT 17.180 200.440 17.320 200.595 ;
        RECT 19.390 200.580 19.710 200.640 ;
        RECT 29.510 200.780 29.830 200.840 ;
        RECT 36.885 200.780 37.175 200.825 ;
        RECT 29.510 200.640 37.175 200.780 ;
        RECT 29.510 200.580 29.830 200.640 ;
        RECT 36.885 200.595 37.175 200.640 ;
        RECT 46.070 200.580 46.390 200.840 ;
        RECT 46.990 200.580 47.310 200.840 ;
        RECT 47.465 200.780 47.755 200.825 ;
        RECT 49.290 200.780 49.610 200.840 ;
        RECT 47.465 200.640 49.610 200.780 ;
        RECT 47.465 200.595 47.755 200.640 ;
        RECT 49.290 200.580 49.610 200.640 ;
        RECT 49.750 200.580 50.070 200.840 ;
        RECT 50.225 200.780 50.515 200.825 ;
        RECT 50.670 200.780 50.990 200.840 ;
        RECT 50.225 200.640 50.990 200.780 ;
        RECT 50.225 200.595 50.515 200.640 ;
        RECT 50.670 200.580 50.990 200.640 ;
        RECT 51.130 200.580 51.450 200.840 ;
        RECT 52.050 200.780 52.370 200.840 ;
        RECT 55.820 200.825 55.960 201.320 ;
        RECT 58.030 201.260 58.350 201.320 ;
        RECT 61.710 201.460 62.030 201.520 ;
        RECT 62.645 201.460 62.935 201.505 ;
        RECT 61.710 201.320 62.935 201.460 ;
        RECT 61.710 201.260 62.030 201.320 ;
        RECT 62.645 201.275 62.935 201.320 ;
        RECT 65.850 201.260 66.170 201.520 ;
        RECT 67.230 201.460 67.550 201.520 ;
        RECT 67.230 201.320 70.680 201.460 ;
        RECT 67.230 201.260 67.550 201.320 ;
        RECT 57.570 200.920 57.890 201.180 ;
        RECT 58.965 201.120 59.255 201.165 ;
        RECT 64.945 201.120 65.235 201.165 ;
        RECT 68.625 201.120 68.915 201.165 ;
        RECT 58.965 200.980 65.235 201.120 ;
        RECT 58.965 200.935 59.255 200.980 ;
        RECT 64.945 200.935 65.235 200.980 ;
        RECT 65.940 200.980 68.915 201.120 ;
        RECT 55.745 200.780 56.035 200.825 ;
        RECT 52.050 200.640 56.035 200.780 ;
        RECT 52.050 200.580 52.370 200.640 ;
        RECT 55.745 200.595 56.035 200.640 ;
        RECT 57.125 200.595 57.415 200.825 ;
        RECT 20.770 200.440 21.090 200.500 ;
        RECT 54.350 200.440 54.670 200.500 ;
        RECT 57.200 200.440 57.340 200.595 ;
        RECT 17.180 200.300 21.090 200.440 ;
        RECT 20.770 200.240 21.090 200.300 ;
        RECT 29.600 200.300 57.340 200.440 ;
        RECT 29.600 200.145 29.740 200.300 ;
        RECT 54.350 200.240 54.670 200.300 ;
        RECT 29.525 199.915 29.815 200.145 ;
        RECT 39.630 200.100 39.950 200.160 ;
        RECT 44.245 200.100 44.535 200.145 ;
        RECT 50.210 200.100 50.530 200.160 ;
        RECT 39.630 199.960 50.530 200.100 ;
        RECT 39.630 199.900 39.950 199.960 ;
        RECT 44.245 199.915 44.535 199.960 ;
        RECT 50.210 199.900 50.530 199.960 ;
        RECT 51.130 200.100 51.450 200.160 ;
        RECT 58.030 200.100 58.350 200.160 ;
        RECT 51.130 199.960 58.350 200.100 ;
        RECT 51.130 199.900 51.450 199.960 ;
        RECT 58.030 199.900 58.350 199.960 ;
        RECT 25.370 199.560 25.690 199.820 ;
        RECT 28.590 199.760 28.910 199.820 ;
        RECT 47.450 199.760 47.770 199.820 ;
        RECT 28.590 199.620 47.770 199.760 ;
        RECT 28.590 199.560 28.910 199.620 ;
        RECT 47.450 199.560 47.770 199.620 ;
        RECT 49.750 199.760 50.070 199.820 ;
        RECT 52.065 199.760 52.355 199.805 ;
        RECT 49.750 199.620 52.355 199.760 ;
        RECT 49.750 199.560 50.070 199.620 ;
        RECT 52.065 199.575 52.355 199.620 ;
        RECT 52.510 199.760 52.830 199.820 ;
        RECT 59.040 199.760 59.180 200.935 ;
        RECT 65.940 200.840 66.080 200.980 ;
        RECT 68.625 200.935 68.915 200.980 ;
        RECT 69.070 200.920 69.390 201.180 ;
        RECT 59.870 200.825 60.190 200.840 ;
        RECT 59.870 200.595 60.325 200.825 ;
        RECT 60.805 200.780 61.095 200.825 ;
        RECT 62.630 200.780 62.950 200.840 ;
        RECT 60.805 200.640 62.950 200.780 ;
        RECT 60.805 200.595 61.095 200.640 ;
        RECT 59.870 200.580 60.190 200.595 ;
        RECT 62.630 200.580 62.950 200.640 ;
        RECT 63.550 200.780 63.870 200.840 ;
        RECT 64.025 200.780 64.315 200.825 ;
        RECT 63.550 200.640 64.315 200.780 ;
        RECT 63.550 200.580 63.870 200.640 ;
        RECT 64.025 200.595 64.315 200.640 ;
        RECT 65.850 200.580 66.170 200.840 ;
        RECT 66.310 200.580 66.630 200.840 ;
        RECT 68.150 200.825 68.470 200.840 ;
        RECT 68.140 200.595 68.470 200.825 ;
        RECT 69.990 200.780 70.310 200.840 ;
        RECT 70.540 200.825 70.680 201.320 ;
        RECT 71.370 201.260 71.690 201.520 ;
        RECT 72.750 201.460 73.070 201.520 ;
        RECT 75.065 201.460 75.355 201.505 ;
        RECT 76.430 201.460 76.750 201.520 ;
        RECT 76.905 201.460 77.195 201.505 ;
        RECT 72.750 201.320 77.195 201.460 ;
        RECT 72.750 201.260 73.070 201.320 ;
        RECT 75.065 201.275 75.355 201.320 ;
        RECT 76.430 201.260 76.750 201.320 ;
        RECT 76.905 201.275 77.195 201.320 ;
        RECT 77.810 201.460 78.130 201.520 ;
        RECT 78.745 201.460 79.035 201.505 ;
        RECT 77.810 201.320 79.035 201.460 ;
        RECT 77.810 201.260 78.130 201.320 ;
        RECT 78.745 201.275 79.035 201.320 ;
        RECT 92.990 201.260 93.310 201.520 ;
        RECT 71.830 201.120 72.150 201.180 ;
        RECT 75.510 201.120 75.830 201.180 ;
        RECT 71.830 200.980 75.830 201.120 ;
        RECT 71.830 200.920 72.150 200.980 ;
        RECT 75.510 200.920 75.830 200.980 ;
        RECT 75.985 201.120 76.275 201.165 ;
        RECT 90.245 201.120 90.535 201.165 ;
        RECT 91.150 201.120 91.470 201.180 ;
        RECT 93.450 201.120 93.770 201.180 ;
        RECT 75.985 200.980 78.040 201.120 ;
        RECT 75.985 200.935 76.275 200.980 ;
        RECT 69.795 200.640 70.310 200.780 ;
        RECT 68.150 200.580 68.470 200.595 ;
        RECT 69.990 200.580 70.310 200.640 ;
        RECT 70.465 200.595 70.755 200.825 ;
        RECT 70.925 200.595 71.215 200.825 ;
        RECT 73.225 200.595 73.515 200.825 ;
        RECT 61.250 200.440 61.570 200.500 ;
        RECT 71.000 200.440 71.140 200.595 ;
        RECT 61.250 200.300 71.140 200.440 ;
        RECT 61.250 200.240 61.570 200.300 ;
        RECT 64.010 200.100 64.330 200.160 ;
        RECT 64.945 200.100 65.235 200.145 ;
        RECT 72.305 200.100 72.595 200.145 ;
        RECT 64.010 199.960 65.235 200.100 ;
        RECT 64.010 199.900 64.330 199.960 ;
        RECT 64.945 199.915 65.235 199.960 ;
        RECT 65.480 199.960 72.595 200.100 ;
        RECT 52.510 199.620 59.180 199.760 ;
        RECT 60.330 199.760 60.650 199.820 ;
        RECT 65.480 199.760 65.620 199.960 ;
        RECT 72.305 199.915 72.595 199.960 ;
        RECT 60.330 199.620 65.620 199.760 ;
        RECT 67.245 199.760 67.535 199.805 ;
        RECT 68.150 199.760 68.470 199.820 ;
        RECT 67.245 199.620 68.470 199.760 ;
        RECT 52.510 199.560 52.830 199.620 ;
        RECT 60.330 199.560 60.650 199.620 ;
        RECT 67.245 199.575 67.535 199.620 ;
        RECT 68.150 199.560 68.470 199.620 ;
        RECT 68.610 199.760 68.930 199.820 ;
        RECT 73.300 199.760 73.440 200.595 ;
        RECT 74.590 200.580 74.910 200.840 ;
        RECT 76.430 200.580 76.750 200.840 ;
        RECT 77.900 200.825 78.040 200.980 ;
        RECT 90.245 200.980 92.760 201.120 ;
        RECT 90.245 200.935 90.535 200.980 ;
        RECT 91.150 200.920 91.470 200.980 ;
        RECT 77.825 200.780 78.115 200.825 ;
        RECT 83.790 200.780 84.110 200.840 ;
        RECT 77.825 200.640 84.110 200.780 ;
        RECT 77.825 200.595 78.115 200.640 ;
        RECT 83.790 200.580 84.110 200.640 ;
        RECT 86.090 200.580 86.410 200.840 ;
        RECT 87.010 200.780 87.330 200.840 ;
        RECT 89.785 200.780 90.075 200.825 ;
        RECT 87.010 200.640 90.075 200.780 ;
        RECT 87.010 200.580 87.330 200.640 ;
        RECT 89.785 200.595 90.075 200.640 ;
        RECT 90.705 200.595 90.995 200.825 ;
        RECT 91.625 200.595 91.915 200.825 ;
        RECT 75.050 200.440 75.370 200.500 ;
        RECT 76.890 200.440 77.210 200.500 ;
        RECT 75.050 200.300 77.210 200.440 ;
        RECT 75.050 200.240 75.370 200.300 ;
        RECT 76.890 200.240 77.210 200.300 ;
        RECT 89.310 200.440 89.630 200.500 ;
        RECT 90.780 200.440 90.920 200.595 ;
        RECT 89.310 200.300 90.920 200.440 ;
        RECT 91.700 200.440 91.840 200.595 ;
        RECT 92.070 200.580 92.390 200.840 ;
        RECT 92.620 200.780 92.760 200.980 ;
        RECT 93.450 200.980 95.520 201.120 ;
        RECT 93.450 200.920 93.770 200.980 ;
        RECT 93.910 200.825 94.230 200.840 ;
        RECT 93.910 200.780 94.365 200.825 ;
        RECT 92.620 200.640 94.365 200.780 ;
        RECT 93.910 200.595 94.365 200.640 ;
        RECT 93.910 200.580 94.230 200.595 ;
        RECT 94.830 200.580 95.150 200.840 ;
        RECT 95.380 200.825 95.520 200.980 ;
        RECT 108.630 200.920 108.950 201.180 ;
        RECT 111.850 200.920 112.170 201.180 ;
        RECT 95.305 200.595 95.595 200.825 ;
        RECT 96.210 200.580 96.530 200.840 ;
        RECT 96.670 200.780 96.990 200.840 ;
        RECT 100.825 200.780 101.115 200.825 ;
        RECT 96.670 200.640 101.115 200.780 ;
        RECT 96.670 200.580 96.990 200.640 ;
        RECT 100.825 200.595 101.115 200.640 ;
        RECT 101.270 200.580 101.590 200.840 ;
        RECT 102.190 200.580 102.510 200.840 ;
        RECT 102.665 200.595 102.955 200.825 ;
        RECT 95.765 200.440 96.055 200.485 ;
        RECT 91.700 200.300 96.055 200.440 ;
        RECT 89.310 200.240 89.630 200.300 ;
        RECT 75.970 199.900 76.290 200.160 ;
        RECT 90.780 200.100 90.920 200.300 ;
        RECT 95.765 200.255 96.055 200.300 ;
        RECT 100.350 200.440 100.670 200.500 ;
        RECT 102.740 200.440 102.880 200.595 ;
        RECT 100.350 200.300 102.880 200.440 ;
        RECT 100.350 200.240 100.670 200.300 ;
        RECT 106.330 200.240 106.650 200.500 ;
        RECT 92.530 200.100 92.850 200.160 ;
        RECT 94.830 200.100 95.150 200.160 ;
        RECT 102.650 200.100 102.970 200.160 ;
        RECT 90.780 199.960 102.970 200.100 ;
        RECT 92.530 199.900 92.850 199.960 ;
        RECT 94.830 199.900 95.150 199.960 ;
        RECT 102.650 199.900 102.970 199.960 ;
        RECT 105.870 200.100 106.190 200.160 ;
        RECT 106.805 200.100 107.095 200.145 ;
        RECT 107.710 200.100 108.030 200.160 ;
        RECT 105.870 199.960 108.030 200.100 ;
        RECT 105.870 199.900 106.190 199.960 ;
        RECT 106.805 199.915 107.095 199.960 ;
        RECT 107.710 199.900 108.030 199.960 ;
        RECT 108.630 200.100 108.950 200.160 ;
        RECT 110.025 200.100 110.315 200.145 ;
        RECT 108.630 199.960 110.315 200.100 ;
        RECT 108.630 199.900 108.950 199.960 ;
        RECT 110.025 199.915 110.315 199.960 ;
        RECT 68.610 199.620 73.440 199.760 ;
        RECT 74.590 199.760 74.910 199.820 ;
        RECT 78.270 199.760 78.590 199.820 ;
        RECT 74.590 199.620 78.590 199.760 ;
        RECT 68.610 199.560 68.930 199.620 ;
        RECT 74.590 199.560 74.910 199.620 ;
        RECT 78.270 199.560 78.590 199.620 ;
        RECT 87.025 199.760 87.315 199.805 ;
        RECT 88.390 199.760 88.710 199.820 ;
        RECT 87.025 199.620 88.710 199.760 ;
        RECT 87.025 199.575 87.315 199.620 ;
        RECT 88.390 199.560 88.710 199.620 ;
        RECT 88.850 199.560 89.170 199.820 ;
        RECT 91.610 199.760 91.930 199.820 ;
        RECT 93.450 199.760 93.770 199.820 ;
        RECT 91.610 199.620 93.770 199.760 ;
        RECT 91.610 199.560 91.930 199.620 ;
        RECT 93.450 199.560 93.770 199.620 ;
        RECT 98.970 199.760 99.290 199.820 ;
        RECT 99.905 199.760 100.195 199.805 ;
        RECT 98.970 199.620 100.195 199.760 ;
        RECT 98.970 199.560 99.290 199.620 ;
        RECT 99.905 199.575 100.195 199.620 ;
        RECT 104.950 199.760 105.270 199.820 ;
        RECT 109.565 199.760 109.855 199.805 ;
        RECT 104.950 199.620 109.855 199.760 ;
        RECT 104.950 199.560 105.270 199.620 ;
        RECT 109.565 199.575 109.855 199.620 ;
        RECT 14.260 198.940 126.960 199.420 ;
        RECT 18.930 198.540 19.250 198.800 ;
        RECT 20.310 198.740 20.630 198.800 ;
        RECT 21.245 198.740 21.535 198.785 ;
        RECT 20.310 198.600 21.535 198.740 ;
        RECT 20.310 198.540 20.630 198.600 ;
        RECT 21.245 198.555 21.535 198.600 ;
        RECT 22.610 198.740 22.930 198.800 ;
        RECT 24.005 198.740 24.295 198.785 ;
        RECT 22.610 198.600 24.295 198.740 ;
        RECT 22.610 198.540 22.930 198.600 ;
        RECT 24.005 198.555 24.295 198.600 ;
        RECT 34.125 198.740 34.415 198.785 ;
        RECT 35.950 198.740 36.270 198.800 ;
        RECT 37.330 198.740 37.650 198.800 ;
        RECT 43.770 198.740 44.090 198.800 ;
        RECT 34.125 198.600 37.650 198.740 ;
        RECT 34.125 198.555 34.415 198.600 ;
        RECT 35.950 198.540 36.270 198.600 ;
        RECT 37.330 198.540 37.650 198.600 ;
        RECT 43.400 198.600 44.090 198.740 ;
        RECT 20.785 198.400 21.075 198.445 ;
        RECT 22.150 198.400 22.470 198.460 ;
        RECT 26.305 198.400 26.595 198.445 ;
        RECT 43.400 198.400 43.540 198.600 ;
        RECT 43.770 198.540 44.090 198.600 ;
        RECT 46.990 198.740 47.310 198.800 ;
        RECT 47.465 198.740 47.755 198.785 ;
        RECT 46.990 198.600 47.755 198.740 ;
        RECT 46.990 198.540 47.310 198.600 ;
        RECT 47.465 198.555 47.755 198.600 ;
        RECT 48.385 198.740 48.675 198.785 ;
        RECT 48.830 198.740 49.150 198.800 ;
        RECT 48.385 198.600 49.150 198.740 ;
        RECT 48.385 198.555 48.675 198.600 ;
        RECT 48.830 198.540 49.150 198.600 ;
        RECT 50.685 198.740 50.975 198.785 ;
        RECT 55.270 198.740 55.590 198.800 ;
        RECT 50.685 198.600 55.590 198.740 ;
        RECT 50.685 198.555 50.975 198.600 ;
        RECT 55.270 198.540 55.590 198.600 ;
        RECT 56.190 198.740 56.510 198.800 ;
        RECT 58.950 198.740 59.270 198.800 ;
        RECT 56.190 198.600 59.270 198.740 ;
        RECT 56.190 198.540 56.510 198.600 ;
        RECT 58.950 198.540 59.270 198.600 ;
        RECT 59.425 198.740 59.715 198.785 ;
        RECT 62.170 198.740 62.490 198.800 ;
        RECT 59.425 198.600 62.490 198.740 ;
        RECT 59.425 198.555 59.715 198.600 ;
        RECT 62.170 198.540 62.490 198.600 ;
        RECT 63.090 198.540 63.410 198.800 ;
        RECT 64.470 198.540 64.790 198.800 ;
        RECT 66.310 198.540 66.630 198.800 ;
        RECT 66.770 198.740 67.090 198.800 ;
        RECT 68.165 198.740 68.455 198.785 ;
        RECT 99.890 198.740 100.210 198.800 ;
        RECT 66.770 198.600 68.455 198.740 ;
        RECT 66.770 198.540 67.090 198.600 ;
        RECT 68.165 198.555 68.455 198.600 ;
        RECT 70.540 198.600 100.210 198.740 ;
        RECT 58.505 198.400 58.795 198.445 ;
        RECT 60.330 198.400 60.650 198.460 ;
        RECT 20.785 198.260 22.470 198.400 ;
        RECT 20.785 198.215 21.075 198.260 ;
        RECT 22.150 198.200 22.470 198.260 ;
        RECT 23.160 198.260 25.140 198.400 ;
        RECT 20.325 198.060 20.615 198.105 ;
        RECT 23.160 198.060 23.300 198.260 ;
        RECT 20.325 197.920 23.300 198.060 ;
        RECT 23.530 198.060 23.850 198.120 ;
        RECT 24.465 198.060 24.755 198.105 ;
        RECT 23.530 197.920 24.755 198.060 ;
        RECT 25.000 198.060 25.140 198.260 ;
        RECT 26.305 198.260 43.540 198.400 ;
        RECT 43.860 198.260 60.650 198.400 ;
        RECT 26.305 198.215 26.595 198.260 ;
        RECT 28.590 198.060 28.910 198.120 ;
        RECT 25.000 197.920 28.910 198.060 ;
        RECT 20.325 197.875 20.615 197.920 ;
        RECT 23.530 197.860 23.850 197.920 ;
        RECT 24.465 197.875 24.755 197.920 ;
        RECT 28.590 197.860 28.910 197.920 ;
        RECT 41.470 197.860 41.790 198.120 ;
        RECT 43.860 198.060 44.000 198.260 ;
        RECT 58.505 198.215 58.795 198.260 ;
        RECT 60.330 198.200 60.650 198.260 ;
        RECT 60.805 198.215 61.095 198.445 ;
        RECT 61.250 198.400 61.570 198.460 ;
        RECT 61.725 198.400 62.015 198.445 ;
        RECT 61.250 198.260 62.015 198.400 ;
        RECT 42.020 197.920 44.000 198.060 ;
        RECT 44.245 198.060 44.535 198.105 ;
        RECT 53.430 198.060 53.750 198.120 ;
        RECT 44.245 197.920 53.750 198.060 ;
        RECT 15.725 197.720 16.015 197.765 ;
        RECT 16.630 197.720 16.950 197.780 ;
        RECT 15.725 197.580 16.950 197.720 ;
        RECT 15.725 197.535 16.015 197.580 ;
        RECT 16.630 197.520 16.950 197.580 ;
        RECT 17.090 197.520 17.410 197.780 ;
        RECT 17.550 197.720 17.870 197.780 ;
        RECT 18.025 197.720 18.315 197.765 ;
        RECT 17.550 197.580 18.315 197.720 ;
        RECT 17.550 197.520 17.870 197.580 ;
        RECT 18.025 197.535 18.315 197.580 ;
        RECT 23.070 197.520 23.390 197.780 ;
        RECT 23.990 197.520 24.310 197.780 ;
        RECT 25.385 197.720 25.675 197.765 ;
        RECT 25.830 197.720 26.150 197.780 ;
        RECT 25.385 197.580 26.150 197.720 ;
        RECT 25.385 197.535 25.675 197.580 ;
        RECT 25.830 197.520 26.150 197.580 ;
        RECT 26.290 197.720 26.610 197.780 ;
        RECT 37.790 197.720 38.110 197.780 ;
        RECT 26.290 197.580 38.110 197.720 ;
        RECT 26.290 197.520 26.610 197.580 ;
        RECT 37.790 197.520 38.110 197.580 ;
        RECT 40.090 197.720 40.410 197.780 ;
        RECT 42.020 197.765 42.160 197.920 ;
        RECT 44.245 197.875 44.535 197.920 ;
        RECT 40.565 197.720 40.855 197.765 ;
        RECT 40.090 197.580 40.855 197.720 ;
        RECT 40.090 197.520 40.410 197.580 ;
        RECT 40.565 197.535 40.855 197.580 ;
        RECT 41.025 197.535 41.315 197.765 ;
        RECT 41.945 197.535 42.235 197.765 ;
        RECT 43.325 197.535 43.615 197.765 ;
        RECT 23.160 197.380 23.300 197.520 ;
        RECT 28.130 197.380 28.450 197.440 ;
        RECT 23.160 197.240 28.450 197.380 ;
        RECT 28.130 197.180 28.450 197.240 ;
        RECT 31.350 197.180 31.670 197.440 ;
        RECT 41.100 197.380 41.240 197.535 ;
        RECT 42.390 197.380 42.710 197.440 ;
        RECT 41.100 197.240 42.710 197.380 ;
        RECT 42.390 197.180 42.710 197.240 ;
        RECT 16.645 197.040 16.935 197.085 ;
        RECT 17.090 197.040 17.410 197.100 ;
        RECT 16.645 196.900 17.410 197.040 ;
        RECT 16.645 196.855 16.935 196.900 ;
        RECT 17.090 196.840 17.410 196.900 ;
        RECT 19.850 197.040 20.170 197.100 ;
        RECT 23.990 197.040 24.310 197.100 ;
        RECT 19.850 196.900 24.310 197.040 ;
        RECT 19.850 196.840 20.170 196.900 ;
        RECT 23.990 196.840 24.310 196.900 ;
        RECT 26.750 197.040 27.070 197.100 ;
        RECT 42.865 197.040 43.155 197.085 ;
        RECT 26.750 196.900 43.155 197.040 ;
        RECT 43.400 197.040 43.540 197.535 ;
        RECT 44.690 197.520 45.010 197.780 ;
        RECT 45.150 197.720 45.470 197.780 ;
        RECT 45.150 197.580 45.665 197.720 ;
        RECT 45.150 197.520 45.470 197.580 ;
        RECT 46.070 197.520 46.390 197.780 ;
        RECT 51.220 197.765 51.360 197.920 ;
        RECT 53.430 197.860 53.750 197.920 ;
        RECT 53.890 197.860 54.210 198.120 ;
        RECT 56.190 198.060 56.510 198.120 ;
        RECT 55.360 197.920 56.510 198.060 ;
        RECT 49.765 197.535 50.055 197.765 ;
        RECT 51.145 197.535 51.435 197.765 ;
        RECT 44.230 197.380 44.550 197.440 ;
        RECT 46.545 197.380 46.835 197.425 ;
        RECT 48.830 197.380 49.150 197.440 ;
        RECT 44.230 197.240 46.835 197.380 ;
        RECT 44.230 197.180 44.550 197.240 ;
        RECT 46.545 197.195 46.835 197.240 ;
        RECT 47.080 197.240 49.150 197.380 ;
        RECT 49.840 197.380 49.980 197.535 ;
        RECT 52.050 197.520 52.370 197.780 ;
        RECT 52.510 197.520 52.830 197.780 ;
        RECT 52.985 197.720 53.275 197.765 ;
        RECT 53.980 197.720 54.120 197.860 ;
        RECT 52.985 197.580 54.120 197.720 ;
        RECT 52.985 197.535 53.275 197.580 ;
        RECT 54.350 197.520 54.670 197.780 ;
        RECT 55.360 197.380 55.500 197.920 ;
        RECT 56.190 197.860 56.510 197.920 ;
        RECT 57.110 197.860 57.430 198.120 ;
        RECT 60.880 198.060 61.020 198.215 ;
        RECT 61.250 198.200 61.570 198.260 ;
        RECT 61.725 198.215 62.015 198.260 ;
        RECT 62.630 198.400 62.950 198.460 ;
        RECT 70.540 198.400 70.680 198.600 ;
        RECT 99.890 198.540 100.210 198.600 ;
        RECT 100.350 198.540 100.670 198.800 ;
        RECT 102.190 198.540 102.510 198.800 ;
        RECT 102.650 198.740 102.970 198.800 ;
        RECT 102.650 198.600 118.750 198.740 ;
        RECT 102.650 198.540 102.970 198.600 ;
        RECT 62.630 198.260 70.680 198.400 ;
        RECT 70.910 198.400 71.230 198.460 ;
        RECT 92.545 198.400 92.835 198.445 ;
        RECT 93.450 198.400 93.770 198.460 ;
        RECT 99.430 198.400 99.750 198.460 ;
        RECT 108.170 198.400 108.490 198.460 ;
        RECT 118.610 198.400 118.750 198.600 ;
        RECT 123.825 198.400 124.115 198.445 ;
        RECT 70.910 198.260 92.300 198.400 ;
        RECT 62.630 198.200 62.950 198.260 ;
        RECT 70.910 198.200 71.230 198.260 ;
        RECT 73.210 198.060 73.530 198.120 ;
        RECT 76.890 198.060 77.210 198.120 ;
        RECT 58.120 197.920 61.020 198.060 ;
        RECT 64.100 197.920 73.530 198.060 ;
        RECT 55.745 197.720 56.035 197.765 ;
        RECT 57.200 197.720 57.340 197.860 ;
        RECT 58.120 197.780 58.260 197.920 ;
        RECT 55.745 197.580 57.340 197.720 ;
        RECT 57.585 197.720 57.875 197.765 ;
        RECT 58.030 197.720 58.350 197.780 ;
        RECT 57.585 197.580 58.350 197.720 ;
        RECT 55.745 197.535 56.035 197.580 ;
        RECT 57.585 197.535 57.875 197.580 ;
        RECT 58.030 197.520 58.350 197.580 ;
        RECT 58.950 197.720 59.270 197.780 ;
        RECT 59.885 197.720 60.175 197.765 ;
        RECT 58.950 197.580 60.175 197.720 ;
        RECT 58.950 197.520 59.270 197.580 ;
        RECT 59.885 197.535 60.175 197.580 ;
        RECT 62.170 197.720 62.490 197.780 ;
        RECT 64.100 197.765 64.240 197.920 ;
        RECT 73.210 197.860 73.530 197.920 ;
        RECT 73.760 197.920 77.210 198.060 ;
        RECT 62.645 197.720 62.935 197.765 ;
        RECT 62.170 197.580 62.935 197.720 ;
        RECT 62.170 197.520 62.490 197.580 ;
        RECT 62.645 197.535 62.935 197.580 ;
        RECT 64.025 197.535 64.315 197.765 ;
        RECT 65.390 197.520 65.710 197.780 ;
        RECT 67.245 197.535 67.535 197.765 ;
        RECT 49.840 197.240 55.500 197.380 ;
        RECT 47.080 197.040 47.220 197.240 ;
        RECT 48.830 197.180 49.150 197.240 ;
        RECT 56.650 197.180 56.970 197.440 ;
        RECT 57.125 197.195 57.415 197.425 ;
        RECT 61.710 197.380 62.030 197.440 ;
        RECT 67.320 197.380 67.460 197.535 ;
        RECT 71.370 197.520 71.690 197.780 ;
        RECT 72.290 197.520 72.610 197.780 ;
        RECT 73.760 197.765 73.900 197.920 ;
        RECT 76.890 197.860 77.210 197.920 ;
        RECT 78.270 198.060 78.590 198.120 ;
        RECT 92.160 198.060 92.300 198.260 ;
        RECT 92.545 198.260 93.770 198.400 ;
        RECT 92.545 198.215 92.835 198.260 ;
        RECT 93.450 198.200 93.770 198.260 ;
        RECT 94.150 198.260 108.860 198.400 ;
        RECT 118.610 198.260 124.115 198.400 ;
        RECT 94.150 198.060 94.290 198.260 ;
        RECT 99.430 198.200 99.750 198.260 ;
        RECT 108.170 198.200 108.490 198.260 ;
        RECT 78.270 197.920 91.840 198.060 ;
        RECT 92.160 197.920 94.290 198.060 ;
        RECT 101.270 198.060 101.590 198.120 ;
        RECT 101.270 197.920 103.340 198.060 ;
        RECT 78.270 197.860 78.590 197.920 ;
        RECT 72.765 197.720 73.055 197.765 ;
        RECT 72.765 197.580 73.440 197.720 ;
        RECT 72.765 197.535 73.055 197.580 ;
        RECT 61.710 197.240 67.460 197.380 ;
        RECT 68.625 197.380 68.915 197.425 ;
        RECT 69.990 197.380 70.310 197.440 ;
        RECT 68.625 197.240 70.310 197.380 ;
        RECT 73.300 197.380 73.440 197.580 ;
        RECT 73.685 197.535 73.975 197.765 ;
        RECT 74.590 197.520 74.910 197.780 ;
        RECT 75.050 197.720 75.370 197.780 ;
        RECT 76.445 197.720 76.735 197.765 ;
        RECT 75.050 197.580 76.735 197.720 ;
        RECT 75.050 197.520 75.370 197.580 ;
        RECT 76.445 197.535 76.735 197.580 ;
        RECT 87.470 197.720 87.790 197.780 ;
        RECT 89.325 197.720 89.615 197.765 ;
        RECT 89.770 197.720 90.090 197.780 ;
        RECT 87.470 197.580 90.090 197.720 ;
        RECT 87.470 197.520 87.790 197.580 ;
        RECT 89.325 197.535 89.615 197.580 ;
        RECT 89.770 197.520 90.090 197.580 ;
        RECT 90.230 197.520 90.550 197.780 ;
        RECT 90.705 197.720 90.995 197.765 ;
        RECT 91.150 197.720 91.470 197.780 ;
        RECT 90.705 197.580 91.470 197.720 ;
        RECT 91.700 197.720 91.840 197.920 ;
        RECT 101.270 197.860 101.590 197.920 ;
        RECT 92.990 197.720 93.310 197.780 ;
        RECT 93.925 197.720 94.215 197.765 ;
        RECT 91.700 197.580 94.215 197.720 ;
        RECT 90.705 197.535 90.995 197.580 ;
        RECT 91.150 197.520 91.470 197.580 ;
        RECT 92.990 197.520 93.310 197.580 ;
        RECT 93.925 197.535 94.215 197.580 ;
        RECT 94.830 197.520 95.150 197.780 ;
        RECT 95.290 197.520 95.610 197.780 ;
        RECT 95.750 197.520 96.070 197.780 ;
        RECT 97.130 197.520 97.450 197.780 ;
        RECT 99.445 197.730 99.735 197.765 ;
        RECT 99.890 197.730 100.210 197.780 ;
        RECT 103.200 197.765 103.340 197.920 ;
        RECT 99.445 197.590 100.210 197.730 ;
        RECT 99.445 197.535 99.735 197.590 ;
        RECT 99.890 197.520 100.210 197.590 ;
        RECT 103.125 197.720 103.415 197.765 ;
        RECT 103.570 197.720 103.890 197.780 ;
        RECT 103.125 197.580 103.890 197.720 ;
        RECT 103.125 197.535 103.415 197.580 ;
        RECT 103.570 197.520 103.890 197.580 ;
        RECT 104.030 197.520 104.350 197.780 ;
        RECT 104.490 197.520 104.810 197.780 ;
        RECT 104.965 197.535 105.255 197.765 ;
        RECT 105.410 197.720 105.730 197.780 ;
        RECT 108.720 197.765 108.860 198.260 ;
        RECT 123.825 198.215 124.115 198.260 ;
        RECT 105.885 197.720 106.175 197.765 ;
        RECT 105.410 197.580 106.175 197.720 ;
        RECT 74.130 197.380 74.450 197.440 ;
        RECT 73.300 197.240 74.450 197.380 ;
        RECT 43.400 196.900 47.220 197.040 ;
        RECT 47.465 197.040 47.755 197.085 ;
        RECT 50.210 197.040 50.530 197.100 ;
        RECT 53.430 197.040 53.750 197.100 ;
        RECT 47.465 196.900 53.750 197.040 ;
        RECT 26.750 196.840 27.070 196.900 ;
        RECT 42.865 196.855 43.155 196.900 ;
        RECT 47.465 196.855 47.755 196.900 ;
        RECT 50.210 196.840 50.530 196.900 ;
        RECT 53.430 196.840 53.750 196.900 ;
        RECT 53.905 197.040 54.195 197.085 ;
        RECT 54.350 197.040 54.670 197.100 ;
        RECT 53.905 196.900 54.670 197.040 ;
        RECT 53.905 196.855 54.195 196.900 ;
        RECT 54.350 196.840 54.670 196.900 ;
        RECT 55.730 197.040 56.050 197.100 ;
        RECT 57.200 197.040 57.340 197.195 ;
        RECT 61.710 197.180 62.030 197.240 ;
        RECT 68.625 197.195 68.915 197.240 ;
        RECT 69.990 197.180 70.310 197.240 ;
        RECT 74.130 197.180 74.450 197.240 ;
        RECT 75.510 197.380 75.830 197.440 ;
        RECT 98.050 197.425 98.370 197.440 ;
        RECT 75.510 197.240 95.520 197.380 ;
        RECT 75.510 197.180 75.830 197.240 ;
        RECT 64.930 197.040 65.250 197.100 ;
        RECT 55.730 196.900 65.250 197.040 ;
        RECT 55.730 196.840 56.050 196.900 ;
        RECT 64.930 196.840 65.250 196.900 ;
        RECT 75.985 197.040 76.275 197.085 ;
        RECT 76.430 197.040 76.750 197.100 ;
        RECT 75.985 196.900 76.750 197.040 ;
        RECT 75.985 196.855 76.275 196.900 ;
        RECT 76.430 196.840 76.750 196.900 ;
        RECT 89.310 197.040 89.630 197.100 ;
        RECT 89.785 197.040 90.075 197.085 ;
        RECT 89.310 196.900 90.075 197.040 ;
        RECT 89.310 196.840 89.630 196.900 ;
        RECT 89.785 196.855 90.075 196.900 ;
        RECT 92.070 197.040 92.390 197.100 ;
        RECT 93.005 197.040 93.295 197.085 ;
        RECT 94.830 197.040 95.150 197.100 ;
        RECT 92.070 196.900 95.150 197.040 ;
        RECT 95.380 197.040 95.520 197.240 ;
        RECT 97.935 197.195 98.370 197.425 ;
        RECT 98.525 197.195 98.815 197.425 ;
        RECT 98.985 197.195 99.275 197.425 ;
        RECT 99.980 197.380 100.120 197.520 ;
        RECT 105.040 197.380 105.180 197.535 ;
        RECT 105.410 197.520 105.730 197.580 ;
        RECT 105.885 197.535 106.175 197.580 ;
        RECT 108.185 197.535 108.475 197.765 ;
        RECT 108.645 197.535 108.935 197.765 ;
        RECT 109.090 197.720 109.410 197.780 ;
        RECT 109.565 197.720 109.855 197.765 ;
        RECT 109.090 197.580 109.855 197.720 ;
        RECT 108.260 197.380 108.400 197.535 ;
        RECT 109.090 197.520 109.410 197.580 ;
        RECT 109.565 197.535 109.855 197.580 ;
        RECT 110.010 197.520 110.330 197.780 ;
        RECT 111.390 197.520 111.710 197.780 ;
        RECT 112.770 197.720 113.090 197.780 ;
        RECT 111.940 197.580 113.090 197.720 ;
        RECT 110.485 197.380 110.775 197.425 ;
        RECT 99.980 197.240 107.940 197.380 ;
        RECT 108.260 197.240 110.775 197.380 ;
        RECT 98.050 197.180 98.370 197.195 ;
        RECT 96.670 197.040 96.990 197.100 ;
        RECT 95.380 196.900 96.990 197.040 ;
        RECT 92.070 196.840 92.390 196.900 ;
        RECT 93.005 196.855 93.295 196.900 ;
        RECT 94.830 196.840 95.150 196.900 ;
        RECT 96.670 196.840 96.990 196.900 ;
        RECT 97.130 197.040 97.450 197.100 ;
        RECT 98.600 197.040 98.740 197.195 ;
        RECT 97.130 196.900 98.740 197.040 ;
        RECT 99.060 197.040 99.200 197.195 ;
        RECT 99.430 197.040 99.750 197.100 ;
        RECT 99.060 196.900 99.750 197.040 ;
        RECT 97.130 196.840 97.450 196.900 ;
        RECT 99.430 196.840 99.750 196.900 ;
        RECT 101.270 197.040 101.590 197.100 ;
        RECT 107.265 197.040 107.555 197.085 ;
        RECT 101.270 196.900 107.555 197.040 ;
        RECT 107.800 197.040 107.940 197.240 ;
        RECT 110.485 197.195 110.775 197.240 ;
        RECT 111.940 197.040 112.080 197.580 ;
        RECT 112.770 197.520 113.090 197.580 ;
        RECT 124.745 197.720 125.035 197.765 ;
        RECT 129.330 197.720 129.650 197.780 ;
        RECT 124.745 197.580 129.650 197.720 ;
        RECT 124.745 197.535 125.035 197.580 ;
        RECT 129.330 197.520 129.650 197.580 ;
        RECT 107.800 196.900 112.080 197.040 ;
        RECT 101.270 196.840 101.590 196.900 ;
        RECT 107.265 196.855 107.555 196.900 ;
        RECT 112.310 196.840 112.630 197.100 ;
        RECT 14.260 196.220 126.960 196.700 ;
        RECT 49.765 196.020 50.055 196.065 ;
        RECT 51.590 196.020 51.910 196.080 ;
        RECT 60.330 196.020 60.650 196.080 ;
        RECT 65.390 196.020 65.710 196.080 ;
        RECT 65.865 196.020 66.155 196.065 ;
        RECT 73.210 196.020 73.530 196.080 ;
        RECT 49.765 195.880 50.440 196.020 ;
        RECT 49.765 195.835 50.055 195.880 ;
        RECT 35.965 195.680 36.255 195.725 ;
        RECT 41.010 195.680 41.330 195.740 ;
        RECT 46.070 195.680 46.390 195.740 ;
        RECT 50.300 195.725 50.440 195.880 ;
        RECT 51.590 195.880 53.200 196.020 ;
        RECT 51.590 195.820 51.910 195.880 ;
        RECT 53.060 195.725 53.200 195.880 ;
        RECT 60.330 195.880 61.025 196.020 ;
        RECT 60.330 195.820 60.650 195.880 ;
        RECT 35.965 195.540 41.330 195.680 ;
        RECT 35.965 195.495 36.255 195.540 ;
        RECT 41.010 195.480 41.330 195.540 ;
        RECT 41.560 195.540 46.390 195.680 ;
        RECT 16.645 195.340 16.935 195.385 ;
        RECT 16.645 195.200 22.150 195.340 ;
        RECT 16.645 195.155 16.935 195.200 ;
        RECT 22.010 195.000 22.150 195.200 ;
        RECT 24.450 195.140 24.770 195.400 ;
        RECT 24.910 195.140 25.230 195.400 ;
        RECT 37.790 195.140 38.110 195.400 ;
        RECT 41.560 195.385 41.700 195.540 ;
        RECT 46.070 195.480 46.390 195.540 ;
        RECT 47.540 195.540 49.060 195.680 ;
        RECT 41.485 195.155 41.775 195.385 ;
        RECT 41.945 195.340 42.235 195.385 ;
        RECT 42.390 195.340 42.710 195.400 ;
        RECT 41.945 195.200 44.000 195.340 ;
        RECT 41.945 195.155 42.235 195.200 ;
        RECT 42.390 195.140 42.710 195.200 ;
        RECT 25.000 195.000 25.140 195.140 ;
        RECT 22.010 194.860 25.140 195.000 ;
        RECT 29.050 195.000 29.370 195.060 ;
        RECT 37.330 195.000 37.650 195.060 ;
        RECT 29.050 194.860 37.650 195.000 ;
        RECT 29.050 194.800 29.370 194.860 ;
        RECT 37.330 194.800 37.650 194.860 ;
        RECT 40.085 195.000 40.375 195.045 ;
        RECT 42.865 195.000 43.155 195.045 ;
        RECT 40.085 194.860 43.155 195.000 ;
        RECT 40.085 194.815 40.375 194.860 ;
        RECT 42.865 194.815 43.155 194.860 ;
        RECT 16.170 194.660 16.490 194.720 ;
        RECT 23.990 194.660 24.310 194.720 ;
        RECT 16.170 194.520 24.310 194.660 ;
        RECT 16.170 194.460 16.490 194.520 ;
        RECT 23.990 194.460 24.310 194.520 ;
        RECT 25.385 194.660 25.675 194.705 ;
        RECT 39.645 194.660 39.935 194.705 ;
        RECT 41.010 194.660 41.330 194.720 ;
        RECT 25.385 194.520 39.400 194.660 ;
        RECT 25.385 194.475 25.675 194.520 ;
        RECT 29.510 194.120 29.830 194.380 ;
        RECT 34.570 194.320 34.890 194.380 ;
        RECT 37.345 194.320 37.635 194.365 ;
        RECT 34.570 194.180 37.635 194.320 ;
        RECT 39.260 194.320 39.400 194.520 ;
        RECT 39.645 194.520 41.330 194.660 ;
        RECT 43.860 194.660 44.000 195.200 ;
        RECT 44.230 195.140 44.550 195.400 ;
        RECT 46.530 195.140 46.850 195.400 ;
        RECT 47.540 195.385 47.680 195.540 ;
        RECT 47.465 195.155 47.755 195.385 ;
        RECT 47.910 195.140 48.230 195.400 ;
        RECT 48.370 195.140 48.690 195.400 ;
        RECT 48.920 195.340 49.060 195.540 ;
        RECT 50.225 195.495 50.515 195.725 ;
        RECT 50.760 195.540 52.740 195.680 ;
        RECT 50.760 195.340 50.900 195.540 ;
        RECT 52.600 195.400 52.740 195.540 ;
        RECT 52.985 195.495 53.275 195.725 ;
        RECT 55.270 195.480 55.590 195.740 ;
        RECT 56.650 195.680 56.970 195.740 ;
        RECT 60.885 195.725 61.025 195.880 ;
        RECT 65.390 195.880 66.155 196.020 ;
        RECT 65.390 195.820 65.710 195.880 ;
        RECT 65.865 195.835 66.155 195.880 ;
        RECT 69.620 195.880 73.530 196.020 ;
        RECT 56.650 195.540 60.560 195.680 ;
        RECT 56.650 195.480 56.970 195.540 ;
        RECT 48.920 195.200 50.900 195.340 ;
        RECT 51.130 195.140 51.450 195.400 ;
        RECT 51.590 195.140 51.910 195.400 ;
        RECT 52.510 195.140 52.830 195.400 ;
        RECT 54.365 195.340 54.655 195.385 ;
        RECT 55.360 195.340 55.500 195.480 ;
        RECT 54.365 195.200 55.500 195.340 ;
        RECT 55.730 195.340 56.050 195.400 ;
        RECT 56.205 195.340 56.495 195.385 ;
        RECT 55.730 195.200 56.495 195.340 ;
        RECT 54.365 195.155 54.655 195.200 ;
        RECT 55.730 195.140 56.050 195.200 ;
        RECT 56.205 195.155 56.495 195.200 ;
        RECT 57.110 195.140 57.430 195.400 ;
        RECT 57.570 195.140 57.890 195.400 ;
        RECT 58.030 195.140 58.350 195.400 ;
        RECT 59.410 195.140 59.730 195.400 ;
        RECT 60.420 195.385 60.560 195.540 ;
        RECT 60.805 195.495 61.095 195.725 ;
        RECT 62.630 195.680 62.950 195.740 ;
        RECT 62.630 195.540 64.240 195.680 ;
        RECT 62.630 195.480 62.950 195.540 ;
        RECT 60.345 195.155 60.635 195.385 ;
        RECT 62.170 195.340 62.490 195.400 ;
        RECT 64.100 195.385 64.240 195.540 ;
        RECT 64.470 195.480 64.790 195.740 ;
        RECT 64.945 195.680 65.235 195.725 ;
        RECT 67.230 195.680 67.550 195.740 ;
        RECT 64.945 195.540 67.550 195.680 ;
        RECT 64.945 195.495 65.235 195.540 ;
        RECT 67.230 195.480 67.550 195.540 ;
        RECT 67.705 195.680 67.995 195.725 ;
        RECT 69.620 195.680 69.760 195.880 ;
        RECT 73.210 195.820 73.530 195.880 ;
        RECT 76.890 196.020 77.210 196.080 ;
        RECT 79.205 196.020 79.495 196.065 ;
        RECT 83.790 196.020 84.110 196.080 ;
        RECT 98.510 196.020 98.830 196.080 ;
        RECT 102.665 196.020 102.955 196.065 ;
        RECT 76.890 195.880 83.100 196.020 ;
        RECT 76.890 195.820 77.210 195.880 ;
        RECT 79.205 195.835 79.495 195.880 ;
        RECT 67.705 195.540 69.760 195.680 ;
        RECT 69.990 195.680 70.310 195.740 ;
        RECT 70.465 195.680 70.755 195.725 ;
        RECT 75.510 195.680 75.830 195.740 ;
        RECT 69.990 195.540 75.830 195.680 ;
        RECT 67.705 195.495 67.995 195.540 ;
        RECT 69.990 195.480 70.310 195.540 ;
        RECT 70.465 195.495 70.755 195.540 ;
        RECT 75.510 195.480 75.830 195.540 ;
        RECT 75.970 195.680 76.290 195.740 ;
        RECT 76.445 195.680 76.735 195.725 ;
        RECT 79.650 195.680 79.970 195.740 ;
        RECT 81.490 195.680 81.810 195.740 ;
        RECT 82.960 195.680 83.100 195.880 ;
        RECT 83.790 195.880 92.760 196.020 ;
        RECT 83.790 195.820 84.110 195.880 ;
        RECT 92.070 195.680 92.390 195.740 ;
        RECT 75.970 195.540 76.735 195.680 ;
        RECT 75.970 195.480 76.290 195.540 ;
        RECT 76.445 195.495 76.735 195.540 ;
        RECT 76.980 195.540 81.260 195.680 ;
        RECT 63.565 195.340 63.855 195.385 ;
        RECT 61.290 195.240 61.580 195.335 ;
        RECT 60.885 195.105 61.580 195.240 ;
        RECT 62.170 195.200 63.855 195.340 ;
        RECT 62.170 195.140 62.490 195.200 ;
        RECT 63.565 195.155 63.855 195.200 ;
        RECT 64.025 195.155 64.315 195.385 ;
        RECT 60.885 195.100 61.480 195.105 ;
        RECT 45.165 195.000 45.455 195.045 ;
        RECT 52.970 195.000 53.290 195.060 ;
        RECT 45.165 194.860 53.290 195.000 ;
        RECT 45.165 194.815 45.455 194.860 ;
        RECT 52.970 194.800 53.290 194.860 ;
        RECT 54.825 194.815 55.115 195.045 ;
        RECT 60.885 195.000 61.025 195.100 ;
        RECT 58.120 194.860 61.025 195.000 ;
        RECT 48.370 194.660 48.690 194.720 ;
        RECT 49.750 194.660 50.070 194.720 ;
        RECT 43.860 194.520 50.070 194.660 ;
        RECT 54.900 194.660 55.040 194.815 ;
        RECT 55.270 194.660 55.590 194.720 ;
        RECT 54.900 194.520 55.590 194.660 ;
        RECT 39.645 194.475 39.935 194.520 ;
        RECT 41.010 194.460 41.330 194.520 ;
        RECT 48.370 194.460 48.690 194.520 ;
        RECT 49.750 194.460 50.070 194.520 ;
        RECT 55.270 194.460 55.590 194.520 ;
        RECT 40.550 194.320 40.870 194.380 ;
        RECT 39.260 194.180 40.870 194.320 ;
        RECT 34.570 194.120 34.890 194.180 ;
        RECT 37.345 194.135 37.635 194.180 ;
        RECT 40.550 194.120 40.870 194.180 ;
        RECT 45.150 194.320 45.470 194.380 ;
        RECT 47.910 194.320 48.230 194.380 ;
        RECT 45.150 194.180 48.230 194.320 ;
        RECT 45.150 194.120 45.470 194.180 ;
        RECT 47.910 194.120 48.230 194.180 ;
        RECT 50.210 194.120 50.530 194.380 ;
        RECT 55.745 194.320 56.035 194.365 ;
        RECT 56.190 194.320 56.510 194.380 ;
        RECT 58.120 194.320 58.260 194.860 ;
        RECT 58.950 194.460 59.270 194.720 ;
        RECT 64.010 194.660 64.330 194.720 ;
        RECT 60.850 194.520 64.330 194.660 ;
        RECT 55.745 194.180 58.260 194.320 ;
        RECT 59.425 194.320 59.715 194.365 ;
        RECT 60.850 194.320 60.990 194.520 ;
        RECT 64.010 194.460 64.330 194.520 ;
        RECT 59.425 194.180 60.990 194.320 ;
        RECT 62.645 194.320 62.935 194.365 ;
        RECT 63.550 194.320 63.870 194.380 ;
        RECT 64.560 194.365 64.700 195.480 ;
        RECT 66.310 195.340 66.630 195.400 ;
        RECT 66.785 195.340 67.075 195.385 ;
        RECT 66.310 195.200 67.075 195.340 ;
        RECT 66.310 195.140 66.630 195.200 ;
        RECT 66.785 195.155 67.075 195.200 ;
        RECT 68.150 195.140 68.470 195.400 ;
        RECT 69.085 195.155 69.375 195.385 ;
        RECT 69.545 195.340 69.835 195.385 ;
        RECT 76.980 195.340 77.120 195.540 ;
        RECT 79.650 195.480 79.970 195.540 ;
        RECT 69.545 195.200 77.120 195.340 ;
        RECT 69.545 195.155 69.835 195.200 ;
        RECT 77.365 195.155 77.655 195.385 ;
        RECT 65.850 195.000 66.170 195.060 ;
        RECT 69.160 195.000 69.300 195.155 ;
        RECT 65.850 194.860 69.300 195.000 ;
        RECT 71.370 195.000 71.690 195.060 ;
        RECT 75.525 195.000 75.815 195.045 ;
        RECT 71.370 194.860 75.815 195.000 ;
        RECT 65.850 194.800 66.170 194.860 ;
        RECT 71.370 194.800 71.690 194.860 ;
        RECT 75.525 194.815 75.815 194.860 ;
        RECT 66.785 194.660 67.075 194.705 ;
        RECT 74.130 194.660 74.450 194.720 ;
        RECT 66.785 194.520 74.450 194.660 ;
        RECT 66.785 194.475 67.075 194.520 ;
        RECT 74.130 194.460 74.450 194.520 ;
        RECT 62.645 194.180 63.870 194.320 ;
        RECT 55.745 194.135 56.035 194.180 ;
        RECT 56.190 194.120 56.510 194.180 ;
        RECT 59.425 194.135 59.715 194.180 ;
        RECT 62.645 194.135 62.935 194.180 ;
        RECT 63.550 194.120 63.870 194.180 ;
        RECT 64.485 194.320 64.775 194.365 ;
        RECT 64.930 194.320 65.250 194.380 ;
        RECT 64.485 194.180 65.250 194.320 ;
        RECT 64.485 194.135 64.775 194.180 ;
        RECT 64.930 194.120 65.250 194.180 ;
        RECT 70.465 194.320 70.755 194.365 ;
        RECT 72.290 194.320 72.610 194.380 ;
        RECT 70.465 194.180 72.610 194.320 ;
        RECT 75.600 194.320 75.740 194.815 ;
        RECT 77.440 194.660 77.580 195.155 ;
        RECT 78.270 195.140 78.590 195.400 ;
        RECT 78.745 195.155 79.035 195.385 ;
        RECT 80.110 195.340 80.430 195.400 ;
        RECT 81.120 195.385 81.260 195.540 ;
        RECT 81.490 195.540 82.640 195.680 ;
        RECT 82.960 195.540 92.390 195.680 ;
        RECT 92.620 195.680 92.760 195.880 ;
        RECT 98.510 195.880 102.955 196.020 ;
        RECT 98.510 195.820 98.830 195.880 ;
        RECT 102.665 195.835 102.955 195.880 ;
        RECT 109.090 195.820 109.410 196.080 ;
        RECT 109.565 196.020 109.855 196.065 ;
        RECT 110.010 196.020 110.330 196.080 ;
        RECT 109.565 195.880 110.330 196.020 ;
        RECT 109.565 195.835 109.855 195.880 ;
        RECT 110.010 195.820 110.330 195.880 ;
        RECT 124.745 196.020 125.035 196.065 ;
        RECT 128.410 196.020 128.730 196.080 ;
        RECT 124.745 195.880 128.730 196.020 ;
        RECT 124.745 195.835 125.035 195.880 ;
        RECT 128.410 195.820 128.730 195.880 ;
        RECT 111.390 195.680 111.710 195.740 ;
        RECT 92.620 195.540 111.710 195.680 ;
        RECT 81.490 195.480 81.810 195.540 ;
        RECT 80.585 195.340 80.875 195.385 ;
        RECT 80.110 195.200 80.875 195.340 ;
        RECT 77.810 195.000 78.130 195.060 ;
        RECT 78.820 195.000 78.960 195.155 ;
        RECT 80.110 195.140 80.430 195.200 ;
        RECT 80.585 195.155 80.875 195.200 ;
        RECT 81.045 195.155 81.335 195.385 ;
        RECT 81.950 195.140 82.270 195.400 ;
        RECT 82.500 195.385 82.640 195.540 ;
        RECT 92.070 195.480 92.390 195.540 ;
        RECT 82.425 195.155 82.715 195.385 ;
        RECT 82.870 195.140 83.190 195.400 ;
        RECT 83.330 195.340 83.650 195.400 ;
        RECT 89.785 195.340 90.075 195.385 ;
        RECT 83.330 195.200 90.075 195.340 ;
        RECT 83.330 195.140 83.650 195.200 ;
        RECT 89.785 195.155 90.075 195.200 ;
        RECT 90.690 195.140 91.010 195.400 ;
        RECT 92.530 195.140 92.850 195.400 ;
        RECT 93.910 195.140 94.230 195.400 ;
        RECT 103.110 195.340 103.430 195.400 ;
        RECT 103.585 195.340 103.875 195.385 ;
        RECT 103.110 195.200 103.875 195.340 ;
        RECT 103.110 195.140 103.430 195.200 ;
        RECT 103.585 195.155 103.875 195.200 ;
        RECT 104.490 195.140 104.810 195.400 ;
        RECT 105.870 195.340 106.190 195.400 ;
        RECT 106.345 195.340 106.635 195.385 ;
        RECT 105.870 195.200 106.635 195.340 ;
        RECT 105.870 195.140 106.190 195.200 ;
        RECT 106.345 195.155 106.635 195.200 ;
        RECT 107.250 195.140 107.570 195.400 ;
        RECT 108.260 195.385 108.400 195.540 ;
        RECT 111.390 195.480 111.710 195.540 ;
        RECT 108.185 195.155 108.475 195.385 ;
        RECT 109.090 195.340 109.410 195.400 ;
        RECT 110.485 195.340 110.775 195.385 ;
        RECT 109.090 195.200 110.775 195.340 ;
        RECT 109.090 195.140 109.410 195.200 ;
        RECT 110.485 195.155 110.775 195.200 ;
        RECT 112.310 195.340 112.630 195.400 ;
        RECT 121.525 195.340 121.815 195.385 ;
        RECT 123.825 195.340 124.115 195.385 ;
        RECT 112.310 195.200 121.815 195.340 ;
        RECT 112.310 195.140 112.630 195.200 ;
        RECT 121.525 195.155 121.815 195.200 ;
        RECT 122.520 195.200 124.115 195.340 ;
        RECT 77.810 194.860 78.960 195.000 ;
        RECT 79.665 195.000 79.955 195.045 ;
        RECT 83.790 195.000 84.110 195.060 ;
        RECT 79.665 194.860 84.110 195.000 ;
        RECT 77.810 194.800 78.130 194.860 ;
        RECT 79.665 194.815 79.955 194.860 ;
        RECT 83.790 194.800 84.110 194.860 ;
        RECT 87.930 195.000 88.250 195.060 ;
        RECT 94.000 195.000 94.140 195.140 ;
        RECT 87.930 194.860 94.140 195.000 ;
        RECT 104.030 195.000 104.350 195.060 ;
        RECT 106.805 195.000 107.095 195.045 ;
        RECT 104.030 194.860 107.095 195.000 ;
        RECT 107.340 195.000 107.480 195.140 ;
        RECT 111.405 195.000 111.695 195.045 ;
        RECT 107.340 194.860 111.695 195.000 ;
        RECT 87.930 194.800 88.250 194.860 ;
        RECT 104.030 194.800 104.350 194.860 ;
        RECT 106.805 194.815 107.095 194.860 ;
        RECT 111.405 194.815 111.695 194.860 ;
        RECT 80.125 194.660 80.415 194.705 ;
        RECT 81.490 194.660 81.810 194.720 ;
        RECT 104.950 194.660 105.270 194.720 ;
        RECT 107.265 194.660 107.555 194.705 ;
        RECT 108.170 194.660 108.490 194.720 ;
        RECT 77.440 194.520 81.810 194.660 ;
        RECT 80.125 194.475 80.415 194.520 ;
        RECT 81.490 194.460 81.810 194.520 ;
        RECT 82.985 194.520 108.490 194.660 ;
        RECT 111.480 194.660 111.620 194.815 ;
        RECT 112.310 194.660 112.630 194.720 ;
        RECT 122.520 194.705 122.660 195.200 ;
        RECT 123.825 195.155 124.115 195.200 ;
        RECT 111.480 194.520 112.630 194.660 ;
        RECT 78.270 194.320 78.590 194.380 ;
        RECT 75.600 194.180 78.590 194.320 ;
        RECT 70.465 194.135 70.755 194.180 ;
        RECT 72.290 194.120 72.610 194.180 ;
        RECT 78.270 194.120 78.590 194.180 ;
        RECT 80.570 194.320 80.890 194.380 ;
        RECT 82.985 194.320 83.125 194.520 ;
        RECT 104.950 194.460 105.270 194.520 ;
        RECT 107.265 194.475 107.555 194.520 ;
        RECT 108.170 194.460 108.490 194.520 ;
        RECT 112.310 194.460 112.630 194.520 ;
        RECT 122.445 194.475 122.735 194.705 ;
        RECT 80.570 194.180 83.125 194.320 ;
        RECT 80.570 194.120 80.890 194.180 ;
        RECT 84.250 194.120 84.570 194.380 ;
        RECT 87.010 194.320 87.330 194.380 ;
        RECT 90.245 194.320 90.535 194.365 ;
        RECT 87.010 194.180 90.535 194.320 ;
        RECT 87.010 194.120 87.330 194.180 ;
        RECT 90.245 194.135 90.535 194.180 ;
        RECT 90.690 194.320 91.010 194.380 ;
        RECT 92.085 194.320 92.375 194.365 ;
        RECT 90.690 194.180 92.375 194.320 ;
        RECT 90.690 194.120 91.010 194.180 ;
        RECT 92.085 194.135 92.375 194.180 ;
        RECT 104.030 194.320 104.350 194.380 ;
        RECT 105.425 194.320 105.715 194.365 ;
        RECT 104.030 194.180 105.715 194.320 ;
        RECT 104.030 194.120 104.350 194.180 ;
        RECT 105.425 194.135 105.715 194.180 ;
        RECT 14.260 193.500 126.960 193.980 ;
        RECT 16.170 193.100 16.490 193.360 ;
        RECT 19.865 193.300 20.155 193.345 ;
        RECT 21.690 193.300 22.010 193.360 ;
        RECT 19.865 193.160 22.010 193.300 ;
        RECT 19.865 193.115 20.155 193.160 ;
        RECT 21.690 193.100 22.010 193.160 ;
        RECT 23.990 193.300 24.310 193.360 ;
        RECT 38.250 193.300 38.570 193.360 ;
        RECT 23.990 193.160 38.570 193.300 ;
        RECT 23.990 193.100 24.310 193.160 ;
        RECT 38.250 193.100 38.570 193.160 ;
        RECT 41.930 193.100 42.250 193.360 ;
        RECT 44.230 193.300 44.550 193.360 ;
        RECT 49.765 193.300 50.055 193.345 ;
        RECT 44.230 193.160 50.055 193.300 ;
        RECT 44.230 193.100 44.550 193.160 ;
        RECT 49.765 193.115 50.055 193.160 ;
        RECT 51.145 193.300 51.435 193.345 ;
        RECT 51.590 193.300 51.910 193.360 ;
        RECT 51.145 193.160 51.910 193.300 ;
        RECT 51.145 193.115 51.435 193.160 ;
        RECT 51.590 193.100 51.910 193.160 ;
        RECT 52.970 193.300 53.290 193.360 ;
        RECT 55.745 193.300 56.035 193.345 ;
        RECT 60.345 193.300 60.635 193.345 ;
        RECT 65.850 193.300 66.170 193.360 ;
        RECT 72.750 193.300 73.070 193.360 ;
        RECT 79.190 193.300 79.510 193.360 ;
        RECT 52.970 193.160 53.660 193.300 ;
        RECT 52.970 193.100 53.290 193.160 ;
        RECT 18.930 192.960 19.250 193.020 ;
        RECT 52.050 192.960 52.370 193.020 ;
        RECT 17.640 192.820 46.300 192.960 ;
        RECT 17.090 192.080 17.410 192.340 ;
        RECT 17.640 192.325 17.780 192.820 ;
        RECT 18.930 192.760 19.250 192.820 ;
        RECT 20.685 192.620 20.975 192.665 ;
        RECT 22.610 192.620 22.930 192.680 ;
        RECT 23.990 192.620 24.310 192.680 ;
        RECT 20.685 192.480 22.150 192.620 ;
        RECT 20.685 192.435 20.975 192.480 ;
        RECT 17.565 192.095 17.855 192.325 ;
        RECT 18.470 192.080 18.790 192.340 ;
        RECT 18.945 192.095 19.235 192.325 ;
        RECT 19.020 191.600 19.160 192.095 ;
        RECT 21.230 192.080 21.550 192.340 ;
        RECT 22.010 192.280 22.150 192.480 ;
        RECT 22.610 192.480 24.310 192.620 ;
        RECT 22.610 192.420 22.930 192.480 ;
        RECT 23.990 192.420 24.310 192.480 ;
        RECT 24.450 192.620 24.770 192.680 ;
        RECT 36.410 192.620 36.730 192.680 ;
        RECT 46.160 192.665 46.300 192.820 ;
        RECT 52.050 192.820 53.200 192.960 ;
        RECT 52.050 192.760 52.370 192.820 ;
        RECT 45.165 192.620 45.455 192.665 ;
        RECT 24.450 192.480 36.180 192.620 ;
        RECT 24.450 192.420 24.770 192.480 ;
        RECT 22.010 192.140 25.140 192.280 ;
        RECT 22.610 191.740 22.930 192.000 ;
        RECT 23.070 191.740 23.390 192.000 ;
        RECT 25.000 191.940 25.140 192.140 ;
        RECT 25.370 192.080 25.690 192.340 ;
        RECT 26.765 192.280 27.055 192.325 ;
        RECT 27.210 192.280 27.530 192.340 ;
        RECT 28.680 192.325 28.820 192.480 ;
        RECT 26.765 192.140 27.530 192.280 ;
        RECT 26.765 192.095 27.055 192.140 ;
        RECT 27.210 192.080 27.530 192.140 ;
        RECT 28.605 192.095 28.895 192.325 ;
        RECT 29.985 192.280 30.275 192.325 ;
        RECT 34.110 192.280 34.430 192.340 ;
        RECT 35.505 192.280 35.795 192.325 ;
        RECT 29.985 192.140 33.880 192.280 ;
        RECT 29.985 192.095 30.275 192.140 ;
        RECT 29.065 191.940 29.355 191.985 ;
        RECT 31.350 191.940 31.670 192.000 ;
        RECT 25.000 191.800 31.670 191.940 ;
        RECT 29.065 191.755 29.355 191.800 ;
        RECT 31.350 191.740 31.670 191.800 ;
        RECT 31.825 191.940 32.115 191.985 ;
        RECT 32.270 191.940 32.590 192.000 ;
        RECT 31.825 191.800 32.590 191.940 ;
        RECT 33.740 191.940 33.880 192.140 ;
        RECT 34.110 192.140 35.795 192.280 ;
        RECT 36.040 192.280 36.180 192.480 ;
        RECT 36.410 192.480 45.455 192.620 ;
        RECT 36.410 192.420 36.730 192.480 ;
        RECT 45.165 192.435 45.455 192.480 ;
        RECT 46.085 192.435 46.375 192.665 ;
        RECT 48.370 192.620 48.690 192.680 ;
        RECT 53.060 192.665 53.200 192.820 ;
        RECT 53.520 192.665 53.660 193.160 ;
        RECT 55.745 193.160 59.410 193.300 ;
        RECT 55.745 193.115 56.035 193.160 ;
        RECT 54.350 192.960 54.670 193.020 ;
        RECT 56.650 192.960 56.970 193.020 ;
        RECT 54.350 192.820 56.970 192.960 ;
        RECT 59.270 192.960 59.410 193.160 ;
        RECT 60.345 193.160 66.170 193.300 ;
        RECT 60.345 193.115 60.635 193.160 ;
        RECT 65.850 193.100 66.170 193.160 ;
        RECT 69.620 193.160 73.070 193.300 ;
        RECT 68.150 192.960 68.470 193.020 ;
        RECT 59.270 192.820 59.640 192.960 ;
        RECT 54.350 192.760 54.670 192.820 ;
        RECT 56.650 192.760 56.970 192.820 ;
        RECT 47.540 192.480 48.690 192.620 ;
        RECT 41.010 192.280 41.330 192.340 ;
        RECT 36.040 192.140 41.330 192.280 ;
        RECT 34.110 192.080 34.430 192.140 ;
        RECT 35.505 192.095 35.795 192.140 ;
        RECT 41.010 192.080 41.330 192.140 ;
        RECT 43.770 192.280 44.090 192.340 ;
        RECT 46.990 192.280 47.310 192.340 ;
        RECT 47.540 192.325 47.680 192.480 ;
        RECT 48.370 192.420 48.690 192.480 ;
        RECT 50.300 192.480 52.740 192.620 ;
        RECT 43.770 192.140 47.310 192.280 ;
        RECT 43.770 192.080 44.090 192.140 ;
        RECT 46.990 192.080 47.310 192.140 ;
        RECT 47.465 192.095 47.755 192.325 ;
        RECT 47.910 192.080 48.230 192.340 ;
        RECT 49.765 192.280 50.055 192.325 ;
        RECT 50.300 192.280 50.440 192.480 ;
        RECT 49.765 192.140 50.440 192.280 ;
        RECT 50.685 192.280 50.975 192.325 ;
        RECT 51.130 192.280 51.450 192.340 ;
        RECT 50.685 192.140 51.450 192.280 ;
        RECT 49.765 192.095 50.055 192.140 ;
        RECT 50.685 192.095 50.975 192.140 ;
        RECT 51.130 192.080 51.450 192.140 ;
        RECT 52.065 192.095 52.355 192.325 ;
        RECT 52.600 192.280 52.740 192.480 ;
        RECT 52.985 192.435 53.275 192.665 ;
        RECT 53.445 192.435 53.735 192.665 ;
        RECT 55.730 192.420 56.050 192.680 ;
        RECT 56.190 192.620 56.510 192.680 ;
        RECT 59.500 192.620 59.640 192.820 ;
        RECT 63.180 192.820 68.470 192.960 ;
        RECT 61.265 192.620 61.555 192.665 ;
        RECT 56.190 192.480 57.825 192.620 ;
        RECT 56.190 192.420 56.510 192.480 ;
        RECT 53.890 192.280 54.210 192.340 ;
        RECT 52.600 192.140 54.210 192.280 ;
        RECT 50.210 191.940 50.530 192.000 ;
        RECT 33.740 191.800 50.530 191.940 ;
        RECT 52.140 191.940 52.280 192.095 ;
        RECT 53.890 192.080 54.210 192.140 ;
        RECT 54.825 192.280 55.115 192.325 ;
        RECT 55.820 192.280 55.960 192.420 ;
        RECT 54.825 192.140 55.960 192.280 ;
        RECT 54.825 192.095 55.115 192.140 ;
        RECT 56.650 192.080 56.970 192.340 ;
        RECT 57.685 192.325 57.825 192.480 ;
        RECT 58.490 192.325 58.810 192.510 ;
        RECT 59.500 192.480 61.555 192.620 ;
        RECT 61.265 192.435 61.555 192.480 ;
        RECT 61.710 192.420 62.030 192.680 ;
        RECT 57.610 192.095 57.900 192.325 ;
        RECT 58.490 192.280 58.830 192.325 ;
        RECT 59.425 192.280 59.715 192.325 ;
        RECT 58.120 192.140 58.830 192.280 ;
        RECT 55.745 191.940 56.035 191.985 ;
        RECT 56.190 191.940 56.510 192.000 ;
        RECT 52.140 191.800 55.500 191.940 ;
        RECT 31.825 191.755 32.115 191.800 ;
        RECT 32.270 191.740 32.590 191.800 ;
        RECT 50.210 191.740 50.530 191.800 ;
        RECT 55.360 191.660 55.500 191.800 ;
        RECT 55.745 191.800 56.510 191.940 ;
        RECT 55.745 191.755 56.035 191.800 ;
        RECT 56.190 191.740 56.510 191.800 ;
        RECT 57.125 191.940 57.415 191.985 ;
        RECT 58.120 191.940 58.260 192.140 ;
        RECT 58.540 192.095 58.830 192.140 ;
        RECT 59.040 192.140 59.715 192.280 ;
        RECT 57.125 191.800 58.260 191.940 ;
        RECT 57.125 191.755 57.415 191.800 ;
        RECT 50.670 191.600 50.990 191.660 ;
        RECT 19.020 191.460 50.990 191.600 ;
        RECT 50.670 191.400 50.990 191.460 ;
        RECT 55.270 191.400 55.590 191.660 ;
        RECT 56.280 191.600 56.420 191.740 ;
        RECT 59.040 191.600 59.180 192.140 ;
        RECT 59.425 192.095 59.715 192.140 ;
        RECT 63.180 191.940 63.320 192.820 ;
        RECT 64.010 192.620 64.330 192.680 ;
        RECT 65.480 192.665 65.620 192.820 ;
        RECT 68.150 192.760 68.470 192.820 ;
        RECT 64.945 192.620 65.235 192.665 ;
        RECT 64.010 192.480 65.235 192.620 ;
        RECT 64.010 192.420 64.330 192.480 ;
        RECT 64.945 192.435 65.235 192.480 ;
        RECT 65.405 192.435 65.695 192.665 ;
        RECT 69.620 192.620 69.760 193.160 ;
        RECT 72.750 193.100 73.070 193.160 ;
        RECT 77.900 193.160 79.510 193.300 ;
        RECT 69.990 192.960 70.310 193.020 ;
        RECT 72.305 192.960 72.595 193.005 ;
        RECT 69.990 192.820 72.595 192.960 ;
        RECT 69.990 192.760 70.310 192.820 ;
        RECT 72.305 192.775 72.595 192.820 ;
        RECT 75.510 192.620 75.830 192.680 ;
        RECT 76.890 192.620 77.210 192.680 ;
        RECT 77.900 192.665 78.040 193.160 ;
        RECT 79.190 193.100 79.510 193.160 ;
        RECT 79.650 193.100 79.970 193.360 ;
        RECT 80.585 193.115 80.875 193.345 ;
        RECT 84.250 193.300 84.570 193.360 ;
        RECT 86.105 193.300 86.395 193.345 ;
        RECT 84.250 193.160 86.395 193.300 ;
        RECT 78.730 192.960 79.050 193.020 ;
        RECT 80.660 192.960 80.800 193.115 ;
        RECT 84.250 193.100 84.570 193.160 ;
        RECT 86.105 193.115 86.395 193.160 ;
        RECT 104.490 193.300 104.810 193.360 ;
        RECT 105.425 193.300 105.715 193.345 ;
        RECT 104.490 193.160 105.715 193.300 ;
        RECT 104.490 193.100 104.810 193.160 ;
        RECT 105.425 193.115 105.715 193.160 ;
        RECT 108.630 193.300 108.950 193.360 ;
        RECT 109.550 193.300 109.870 193.360 ;
        RECT 108.630 193.160 109.870 193.300 ;
        RECT 108.630 193.100 108.950 193.160 ;
        RECT 109.550 193.100 109.870 193.160 ;
        RECT 78.730 192.820 80.800 192.960 ;
        RECT 81.950 192.960 82.270 193.020 ;
        RECT 92.990 192.960 93.310 193.020 ;
        RECT 81.950 192.820 93.310 192.960 ;
        RECT 78.730 192.760 79.050 192.820 ;
        RECT 81.950 192.760 82.270 192.820 ;
        RECT 92.990 192.760 93.310 192.820 ;
        RECT 104.950 192.960 105.270 193.020 ;
        RECT 107.250 192.960 107.570 193.020 ;
        RECT 104.950 192.820 107.570 192.960 ;
        RECT 104.950 192.760 105.270 192.820 ;
        RECT 107.250 192.760 107.570 192.820 ;
        RECT 107.710 192.760 108.030 193.020 ;
        RECT 109.090 192.960 109.410 193.020 ;
        RECT 110.485 192.960 110.775 193.005 ;
        RECT 114.610 192.960 114.930 193.020 ;
        RECT 109.090 192.820 110.775 192.960 ;
        RECT 109.090 192.760 109.410 192.820 ;
        RECT 110.485 192.775 110.775 192.820 ;
        RECT 111.480 192.820 114.930 192.960 ;
        RECT 67.320 192.480 69.760 192.620 ;
        RECT 70.540 192.480 72.980 192.620 ;
        RECT 67.320 192.325 67.460 192.480 ;
        RECT 63.565 192.280 63.855 192.325 ;
        RECT 67.245 192.280 67.535 192.325 ;
        RECT 63.565 192.140 67.535 192.280 ;
        RECT 63.565 192.095 63.855 192.140 ;
        RECT 67.245 192.095 67.535 192.140 ;
        RECT 69.530 192.280 69.850 192.340 ;
        RECT 70.540 192.325 70.680 192.480 ;
        RECT 70.000 192.280 70.290 192.325 ;
        RECT 69.530 192.140 70.290 192.280 ;
        RECT 69.530 192.080 69.850 192.140 ;
        RECT 70.000 192.095 70.290 192.140 ;
        RECT 70.465 192.095 70.755 192.325 ;
        RECT 70.910 192.080 71.230 192.340 ;
        RECT 71.845 192.095 72.135 192.325 ;
        RECT 59.500 191.800 63.320 191.940 ;
        RECT 59.500 191.645 59.640 191.800 ;
        RECT 68.610 191.740 68.930 192.000 ;
        RECT 56.280 191.460 59.180 191.600 ;
        RECT 59.425 191.415 59.715 191.645 ;
        RECT 64.010 191.400 64.330 191.660 ;
        RECT 67.690 191.600 68.010 191.660 ;
        RECT 71.920 191.600 72.060 192.095 ;
        RECT 72.290 192.080 72.610 192.340 ;
        RECT 72.840 191.940 72.980 192.480 ;
        RECT 75.510 192.480 77.210 192.620 ;
        RECT 75.510 192.420 75.830 192.480 ;
        RECT 76.890 192.420 77.210 192.480 ;
        RECT 77.825 192.435 78.115 192.665 ;
        RECT 78.270 192.420 78.590 192.680 ;
        RECT 81.490 192.620 81.810 192.680 ;
        RECT 103.570 192.620 103.890 192.680 ;
        RECT 111.480 192.620 111.620 192.820 ;
        RECT 114.610 192.760 114.930 192.820 ;
        RECT 81.490 192.480 111.620 192.620 ;
        RECT 111.850 192.620 112.170 192.680 ;
        RECT 114.165 192.620 114.455 192.665 ;
        RECT 111.850 192.480 114.455 192.620 ;
        RECT 81.490 192.420 81.810 192.480 ;
        RECT 103.570 192.420 103.890 192.480 ;
        RECT 73.210 192.080 73.530 192.340 ;
        RECT 73.670 192.080 73.990 192.340 ;
        RECT 77.365 192.280 77.655 192.325 ;
        RECT 80.570 192.280 80.890 192.340 ;
        RECT 77.365 192.140 80.890 192.280 ;
        RECT 77.365 192.095 77.655 192.140 ;
        RECT 80.570 192.080 80.890 192.140 ;
        RECT 81.045 192.280 81.335 192.325 ;
        RECT 81.950 192.280 82.270 192.340 ;
        RECT 81.045 192.140 82.270 192.280 ;
        RECT 81.045 192.095 81.335 192.140 ;
        RECT 81.950 192.080 82.270 192.140 ;
        RECT 82.425 192.280 82.715 192.325 ;
        RECT 82.870 192.280 83.190 192.340 ;
        RECT 82.425 192.140 83.190 192.280 ;
        RECT 82.425 192.095 82.715 192.140 ;
        RECT 82.870 192.080 83.190 192.140 ;
        RECT 83.330 192.280 83.650 192.340 ;
        RECT 84.035 192.280 84.325 192.325 ;
        RECT 83.330 192.140 84.325 192.280 ;
        RECT 83.330 192.080 83.650 192.140 ;
        RECT 84.035 192.095 84.325 192.140 ;
        RECT 84.710 192.280 85.030 192.340 ;
        RECT 86.565 192.280 86.855 192.325 ;
        RECT 90.690 192.280 91.010 192.340 ;
        RECT 84.710 192.140 91.010 192.280 ;
        RECT 84.710 192.080 85.030 192.140 ;
        RECT 86.565 192.095 86.855 192.140 ;
        RECT 90.690 192.080 91.010 192.140 ;
        RECT 104.030 192.280 104.350 192.340 ;
        RECT 106.880 192.325 107.020 192.480 ;
        RECT 111.850 192.420 112.170 192.480 ;
        RECT 114.165 192.435 114.455 192.480 ;
        RECT 106.345 192.280 106.635 192.325 ;
        RECT 104.030 192.140 106.635 192.280 ;
        RECT 104.030 192.080 104.350 192.140 ;
        RECT 106.345 192.095 106.635 192.140 ;
        RECT 106.805 192.095 107.095 192.325 ;
        RECT 107.710 192.280 108.030 192.340 ;
        RECT 110.470 192.280 110.790 192.340 ;
        RECT 107.710 192.140 110.790 192.280 ;
        RECT 107.710 192.080 108.030 192.140 ;
        RECT 110.470 192.080 110.790 192.140 ;
        RECT 110.930 192.280 111.250 192.340 ;
        RECT 111.405 192.280 111.695 192.325 ;
        RECT 110.930 192.140 111.695 192.280 ;
        RECT 110.930 192.080 111.250 192.140 ;
        RECT 111.405 192.095 111.695 192.140 ;
        RECT 112.310 192.080 112.630 192.340 ;
        RECT 115.085 192.280 115.375 192.325 ;
        RECT 115.530 192.280 115.850 192.340 ;
        RECT 115.085 192.140 115.850 192.280 ;
        RECT 115.085 192.095 115.375 192.140 ;
        RECT 99.890 191.940 100.210 192.000 ;
        RECT 72.840 191.800 100.210 191.940 ;
        RECT 99.890 191.740 100.210 191.800 ;
        RECT 109.565 191.940 109.855 191.985 ;
        RECT 115.160 191.940 115.300 192.095 ;
        RECT 115.530 192.080 115.850 192.140 ;
        RECT 121.510 192.080 121.830 192.340 ;
        RECT 124.745 192.280 125.035 192.325 ;
        RECT 128.410 192.280 128.730 192.340 ;
        RECT 124.745 192.140 128.730 192.280 ;
        RECT 124.745 192.095 125.035 192.140 ;
        RECT 128.410 192.080 128.730 192.140 ;
        RECT 109.565 191.800 115.300 191.940 ;
        RECT 109.565 191.755 109.855 191.800 ;
        RECT 67.690 191.460 72.060 191.600 ;
        RECT 67.690 191.400 68.010 191.460 ;
        RECT 79.190 191.400 79.510 191.660 ;
        RECT 80.110 191.600 80.430 191.660 ;
        RECT 83.345 191.600 83.635 191.645 ;
        RECT 80.110 191.460 83.635 191.600 ;
        RECT 80.110 191.400 80.430 191.460 ;
        RECT 83.345 191.415 83.635 191.460 ;
        RECT 84.265 191.600 84.555 191.645 ;
        RECT 88.850 191.600 89.170 191.660 ;
        RECT 84.265 191.460 89.170 191.600 ;
        RECT 84.265 191.415 84.555 191.460 ;
        RECT 88.850 191.400 89.170 191.460 ;
        RECT 95.750 191.600 96.070 191.660 ;
        RECT 108.630 191.600 108.950 191.660 ;
        RECT 95.750 191.460 108.950 191.600 ;
        RECT 95.750 191.400 96.070 191.460 ;
        RECT 108.630 191.400 108.950 191.460 ;
        RECT 111.850 191.400 112.170 191.660 ;
        RECT 122.445 191.600 122.735 191.645 ;
        RECT 123.810 191.600 124.130 191.660 ;
        RECT 122.445 191.460 124.130 191.600 ;
        RECT 122.445 191.415 122.735 191.460 ;
        RECT 123.810 191.400 124.130 191.460 ;
        RECT 124.270 191.400 124.590 191.660 ;
        RECT 14.260 190.780 126.960 191.260 ;
        RECT 16.185 190.580 16.475 190.625 ;
        RECT 23.070 190.580 23.390 190.640 ;
        RECT 28.590 190.580 28.910 190.640 ;
        RECT 16.185 190.440 22.840 190.580 ;
        RECT 16.185 190.395 16.475 190.440 ;
        RECT 18.945 190.240 19.235 190.285 ;
        RECT 19.390 190.240 19.710 190.300 ;
        RECT 21.230 190.240 21.550 190.300 ;
        RECT 18.945 190.100 21.550 190.240 ;
        RECT 22.700 190.240 22.840 190.440 ;
        RECT 23.070 190.440 28.910 190.580 ;
        RECT 23.070 190.380 23.390 190.440 ;
        RECT 28.590 190.380 28.910 190.440 ;
        RECT 29.525 190.580 29.815 190.625 ;
        RECT 36.870 190.580 37.190 190.640 ;
        RECT 42.850 190.580 43.170 190.640 ;
        RECT 29.525 190.440 36.640 190.580 ;
        RECT 29.525 190.395 29.815 190.440 ;
        RECT 26.290 190.240 26.610 190.300 ;
        RECT 22.700 190.100 26.610 190.240 ;
        RECT 18.945 190.055 19.235 190.100 ;
        RECT 19.390 190.040 19.710 190.100 ;
        RECT 21.230 190.040 21.550 190.100 ;
        RECT 26.290 190.040 26.610 190.100 ;
        RECT 35.950 190.040 36.270 190.300 ;
        RECT 36.500 190.240 36.640 190.440 ;
        RECT 36.870 190.440 43.170 190.580 ;
        RECT 36.870 190.380 37.190 190.440 ;
        RECT 42.850 190.380 43.170 190.440 ;
        RECT 44.690 190.580 45.010 190.640 ;
        RECT 46.545 190.580 46.835 190.625 ;
        RECT 47.910 190.580 48.230 190.640 ;
        RECT 44.690 190.440 46.835 190.580 ;
        RECT 44.690 190.380 45.010 190.440 ;
        RECT 46.545 190.395 46.835 190.440 ;
        RECT 47.080 190.440 48.230 190.580 ;
        RECT 47.080 190.240 47.220 190.440 ;
        RECT 47.910 190.380 48.230 190.440 ;
        RECT 48.830 190.580 49.150 190.640 ;
        RECT 51.130 190.580 51.450 190.640 ;
        RECT 48.830 190.440 51.450 190.580 ;
        RECT 48.830 190.380 49.150 190.440 ;
        RECT 51.130 190.380 51.450 190.440 ;
        RECT 53.890 190.380 54.210 190.640 ;
        RECT 54.350 190.580 54.670 190.640 ;
        RECT 55.730 190.580 56.050 190.640 ;
        RECT 54.350 190.440 58.260 190.580 ;
        RECT 54.350 190.380 54.670 190.440 ;
        RECT 55.730 190.380 56.050 190.440 ;
        RECT 36.500 190.100 47.220 190.240 ;
        RECT 47.450 190.040 47.770 190.300 ;
        RECT 49.750 190.240 50.070 190.300 ;
        RECT 57.110 190.240 57.430 190.300 ;
        RECT 58.120 190.285 58.260 190.440 ;
        RECT 59.410 190.380 59.730 190.640 ;
        RECT 60.330 190.380 60.650 190.640 ;
        RECT 62.630 190.380 62.950 190.640 ;
        RECT 63.550 190.580 63.870 190.640 ;
        RECT 64.025 190.580 64.315 190.625 ;
        RECT 63.550 190.440 64.315 190.580 ;
        RECT 63.550 190.380 63.870 190.440 ;
        RECT 64.025 190.395 64.315 190.440 ;
        RECT 65.390 190.580 65.710 190.640 ;
        RECT 70.910 190.580 71.230 190.640 ;
        RECT 71.845 190.580 72.135 190.625 ;
        RECT 79.650 190.580 79.970 190.640 ;
        RECT 80.125 190.580 80.415 190.625 ;
        RECT 65.390 190.440 67.460 190.580 ;
        RECT 65.390 190.380 65.710 190.440 ;
        RECT 49.750 190.100 57.430 190.240 ;
        RECT 49.750 190.040 50.070 190.100 ;
        RECT 57.110 190.040 57.430 190.100 ;
        RECT 58.045 190.240 58.335 190.285 ;
        RECT 58.950 190.240 59.270 190.300 ;
        RECT 64.930 190.240 65.250 190.300 ;
        RECT 67.320 190.285 67.460 190.440 ;
        RECT 70.910 190.440 72.135 190.580 ;
        RECT 70.910 190.380 71.230 190.440 ;
        RECT 71.845 190.395 72.135 190.440 ;
        RECT 74.680 190.440 79.420 190.580 ;
        RECT 58.045 190.100 59.270 190.240 ;
        RECT 58.045 190.055 58.335 190.100 ;
        RECT 58.950 190.040 59.270 190.100 ;
        RECT 59.960 190.100 65.250 190.240 ;
        RECT 17.105 189.715 17.395 189.945 ;
        RECT 17.180 189.560 17.320 189.715 ;
        RECT 26.750 189.700 27.070 189.960 ;
        RECT 36.410 189.900 36.730 189.960 ;
        RECT 27.275 189.760 36.730 189.900 ;
        RECT 27.275 189.560 27.415 189.760 ;
        RECT 36.410 189.700 36.730 189.760 ;
        RECT 36.870 189.700 37.190 189.960 ;
        RECT 37.805 189.900 38.095 189.945 ;
        RECT 38.250 189.900 38.570 189.960 ;
        RECT 37.805 189.760 38.570 189.900 ;
        RECT 37.805 189.715 38.095 189.760 ;
        RECT 38.250 189.700 38.570 189.760 ;
        RECT 39.645 189.900 39.935 189.945 ;
        RECT 39.645 189.760 41.700 189.900 ;
        RECT 39.645 189.715 39.935 189.760 ;
        RECT 41.560 189.620 41.700 189.760 ;
        RECT 41.930 189.700 42.250 189.960 ;
        RECT 43.310 189.900 43.630 189.960 ;
        RECT 45.610 189.900 45.930 189.960 ;
        RECT 43.310 189.760 45.930 189.900 ;
        RECT 43.310 189.700 43.630 189.760 ;
        RECT 45.610 189.700 45.930 189.760 ;
        RECT 46.085 189.715 46.375 189.945 ;
        RECT 47.005 189.900 47.295 189.945 ;
        RECT 49.290 189.900 49.610 189.960 ;
        RECT 47.005 189.760 49.610 189.900 ;
        RECT 47.005 189.715 47.295 189.760 ;
        RECT 17.180 189.420 27.415 189.560 ;
        RECT 35.030 189.560 35.350 189.620 ;
        RECT 38.725 189.560 39.015 189.605 ;
        RECT 35.030 189.420 39.015 189.560 ;
        RECT 35.030 189.360 35.350 189.420 ;
        RECT 38.725 189.375 39.015 189.420 ;
        RECT 40.090 189.360 40.410 189.620 ;
        RECT 40.565 189.375 40.855 189.605 ;
        RECT 10.190 189.220 10.510 189.280 ;
        RECT 10.190 189.080 35.950 189.220 ;
        RECT 10.190 189.020 10.510 189.080 ;
        RECT 21.690 188.880 22.010 188.940 ;
        RECT 34.570 188.880 34.890 188.940 ;
        RECT 21.690 188.740 34.890 188.880 ;
        RECT 35.810 188.880 35.950 189.080 ;
        RECT 37.330 189.020 37.650 189.280 ;
        RECT 40.640 189.220 40.780 189.375 ;
        RECT 41.010 189.360 41.330 189.620 ;
        RECT 41.470 189.560 41.790 189.620 ;
        RECT 45.150 189.560 45.470 189.620 ;
        RECT 41.470 189.420 45.470 189.560 ;
        RECT 46.160 189.560 46.300 189.715 ;
        RECT 49.290 189.700 49.610 189.760 ;
        RECT 55.730 189.900 56.050 189.960 ;
        RECT 56.665 189.900 56.955 189.945 ;
        RECT 55.730 189.760 56.955 189.900 ;
        RECT 55.730 189.700 56.050 189.760 ;
        RECT 56.665 189.715 56.955 189.760 ;
        RECT 57.585 189.715 57.875 189.945 ;
        RECT 52.510 189.560 52.830 189.620 ;
        RECT 46.160 189.420 52.830 189.560 ;
        RECT 41.470 189.360 41.790 189.420 ;
        RECT 45.150 189.360 45.470 189.420 ;
        RECT 52.510 189.360 52.830 189.420 ;
        RECT 57.660 189.560 57.800 189.715 ;
        RECT 58.490 189.700 58.810 189.960 ;
        RECT 59.960 189.945 60.100 190.100 ;
        RECT 64.930 190.040 65.250 190.100 ;
        RECT 67.245 190.055 67.535 190.285 ;
        RECT 69.160 190.100 73.440 190.240 ;
        RECT 69.160 189.960 69.300 190.100 ;
        RECT 59.885 189.715 60.175 189.945 ;
        RECT 60.805 189.900 61.095 189.945 ;
        RECT 61.710 189.900 62.030 189.960 ;
        RECT 60.805 189.760 62.030 189.900 ;
        RECT 60.805 189.715 61.095 189.760 ;
        RECT 61.710 189.700 62.030 189.760 ;
        RECT 63.550 189.700 63.870 189.960 ;
        RECT 64.010 189.900 64.330 189.960 ;
        RECT 65.865 189.900 66.155 189.945 ;
        RECT 64.010 189.760 66.155 189.900 ;
        RECT 64.010 189.700 64.330 189.760 ;
        RECT 65.865 189.715 66.155 189.760 ;
        RECT 66.325 189.715 66.615 189.945 ;
        RECT 60.330 189.560 60.650 189.620 ;
        RECT 57.660 189.420 60.650 189.560 ;
        RECT 66.400 189.560 66.540 189.715 ;
        RECT 67.690 189.700 68.010 189.960 ;
        RECT 68.150 189.900 68.470 189.960 ;
        RECT 68.620 189.900 68.910 189.945 ;
        RECT 68.150 189.760 68.910 189.900 ;
        RECT 68.150 189.700 68.470 189.760 ;
        RECT 68.620 189.715 68.910 189.760 ;
        RECT 69.070 189.700 69.390 189.960 ;
        RECT 69.545 189.900 69.835 189.945 ;
        RECT 69.990 189.900 70.310 189.960 ;
        RECT 69.545 189.760 70.310 189.900 ;
        RECT 69.545 189.715 69.835 189.760 ;
        RECT 69.990 189.700 70.310 189.760 ;
        RECT 70.450 189.900 70.770 189.960 ;
        RECT 72.290 189.900 72.610 189.960 ;
        RECT 73.300 189.945 73.440 190.100 ;
        RECT 74.680 189.960 74.820 190.440 ;
        RECT 75.510 190.240 75.830 190.300 ;
        RECT 78.730 190.240 79.050 190.300 ;
        RECT 75.510 190.100 79.050 190.240 ;
        RECT 75.510 190.040 75.830 190.100 ;
        RECT 72.765 189.900 73.055 189.945 ;
        RECT 70.450 189.760 72.060 189.900 ;
        RECT 70.450 189.700 70.770 189.760 ;
        RECT 70.910 189.560 71.230 189.620 ;
        RECT 66.400 189.420 71.230 189.560 ;
        RECT 41.930 189.220 42.250 189.280 ;
        RECT 40.640 189.080 42.250 189.220 ;
        RECT 41.930 189.020 42.250 189.080 ;
        RECT 42.390 189.220 42.710 189.280 ;
        RECT 43.770 189.220 44.090 189.280 ;
        RECT 52.970 189.220 53.290 189.280 ;
        RECT 55.270 189.220 55.590 189.280 ;
        RECT 42.390 189.080 51.360 189.220 ;
        RECT 42.390 189.020 42.710 189.080 ;
        RECT 43.770 189.020 44.090 189.080 ;
        RECT 50.670 188.880 50.990 188.940 ;
        RECT 35.810 188.740 50.990 188.880 ;
        RECT 51.220 188.880 51.360 189.080 ;
        RECT 52.970 189.080 55.590 189.220 ;
        RECT 52.970 189.020 53.290 189.080 ;
        RECT 55.270 189.020 55.590 189.080 ;
        RECT 56.650 189.220 56.970 189.280 ;
        RECT 57.660 189.220 57.800 189.420 ;
        RECT 60.330 189.360 60.650 189.420 ;
        RECT 70.910 189.360 71.230 189.420 ;
        RECT 71.370 189.360 71.690 189.620 ;
        RECT 71.920 189.560 72.060 189.760 ;
        RECT 72.290 189.760 73.055 189.900 ;
        RECT 72.290 189.700 72.610 189.760 ;
        RECT 72.765 189.715 73.055 189.760 ;
        RECT 73.225 189.715 73.515 189.945 ;
        RECT 74.590 189.900 74.910 189.960 ;
        RECT 73.760 189.760 74.910 189.900 ;
        RECT 73.760 189.560 73.900 189.760 ;
        RECT 74.590 189.700 74.910 189.760 ;
        RECT 75.970 189.900 76.290 189.960 ;
        RECT 77.900 189.945 78.040 190.100 ;
        RECT 78.730 190.040 79.050 190.100 ;
        RECT 79.280 189.945 79.420 190.440 ;
        RECT 79.650 190.440 80.415 190.580 ;
        RECT 79.650 190.380 79.970 190.440 ;
        RECT 80.125 190.395 80.415 190.440 ;
        RECT 80.570 190.580 80.890 190.640 ;
        RECT 81.045 190.580 81.335 190.625 ;
        RECT 80.570 190.440 81.335 190.580 ;
        RECT 80.570 190.380 80.890 190.440 ;
        RECT 81.045 190.395 81.335 190.440 ;
        RECT 83.330 190.580 83.650 190.640 ;
        RECT 92.990 190.580 93.310 190.640 ;
        RECT 102.190 190.580 102.510 190.640 ;
        RECT 83.330 190.440 92.760 190.580 ;
        RECT 83.330 190.380 83.650 190.440 ;
        RECT 87.010 190.240 87.330 190.300 ;
        RECT 80.660 190.100 87.330 190.240 ;
        RECT 92.620 190.240 92.760 190.440 ;
        RECT 92.990 190.440 102.510 190.580 ;
        RECT 92.990 190.380 93.310 190.440 ;
        RECT 102.190 190.380 102.510 190.440 ;
        RECT 103.110 190.580 103.430 190.640 ;
        RECT 110.025 190.580 110.315 190.625 ;
        RECT 103.110 190.440 110.315 190.580 ;
        RECT 103.110 190.380 103.430 190.440 ;
        RECT 110.025 190.395 110.315 190.440 ;
        RECT 110.470 190.580 110.790 190.640 ;
        RECT 111.405 190.580 111.695 190.625 ;
        RECT 112.310 190.580 112.630 190.640 ;
        RECT 110.470 190.440 112.630 190.580 ;
        RECT 110.470 190.380 110.790 190.440 ;
        RECT 111.405 190.395 111.695 190.440 ;
        RECT 112.310 190.380 112.630 190.440 ;
        RECT 114.610 190.380 114.930 190.640 ;
        RECT 116.910 190.380 117.230 190.640 ;
        RECT 120.145 190.580 120.435 190.625 ;
        RECT 118.610 190.440 120.435 190.580 ;
        RECT 100.350 190.240 100.670 190.300 ;
        RECT 100.825 190.240 101.115 190.285 ;
        RECT 106.330 190.240 106.650 190.300 ;
        RECT 109.090 190.240 109.410 190.300 ;
        RECT 92.620 190.100 101.115 190.240 ;
        RECT 80.660 189.945 80.800 190.100 ;
        RECT 87.010 190.040 87.330 190.100 ;
        RECT 100.350 190.040 100.670 190.100 ;
        RECT 100.825 190.055 101.115 190.100 ;
        RECT 105.040 190.100 109.410 190.240 ;
        RECT 76.905 189.900 77.195 189.945 ;
        RECT 75.970 189.760 77.195 189.900 ;
        RECT 75.970 189.700 76.290 189.760 ;
        RECT 76.905 189.715 77.195 189.760 ;
        RECT 77.825 189.715 78.115 189.945 ;
        RECT 79.205 189.715 79.495 189.945 ;
        RECT 80.585 189.715 80.875 189.945 ;
        RECT 82.870 189.900 83.190 189.960 ;
        RECT 83.805 189.900 84.095 189.945 ;
        RECT 82.870 189.760 84.095 189.900 ;
        RECT 82.870 189.700 83.190 189.760 ;
        RECT 83.805 189.715 84.095 189.760 ;
        RECT 84.250 189.900 84.570 189.960 ;
        RECT 87.485 189.900 87.775 189.945 ;
        RECT 87.930 189.900 88.250 189.960 ;
        RECT 84.250 189.760 88.250 189.900 ;
        RECT 71.920 189.420 73.900 189.560 ;
        RECT 74.130 189.360 74.450 189.620 ;
        RECT 78.285 189.560 78.575 189.605 ;
        RECT 78.730 189.560 79.050 189.620 ;
        RECT 81.950 189.560 82.270 189.620 ;
        RECT 82.425 189.560 82.715 189.605 ;
        RECT 78.285 189.420 79.050 189.560 ;
        RECT 78.285 189.375 78.575 189.420 ;
        RECT 78.730 189.360 79.050 189.420 ;
        RECT 79.280 189.420 82.715 189.560 ;
        RECT 83.880 189.560 84.020 189.715 ;
        RECT 84.250 189.700 84.570 189.760 ;
        RECT 87.485 189.715 87.775 189.760 ;
        RECT 87.930 189.700 88.250 189.760 ;
        RECT 92.070 189.900 92.390 189.960 ;
        RECT 93.465 189.900 93.755 189.945 ;
        RECT 92.070 189.760 93.755 189.900 ;
        RECT 92.070 189.700 92.390 189.760 ;
        RECT 93.465 189.715 93.755 189.760 ;
        RECT 99.430 189.900 99.750 189.960 ;
        RECT 99.905 189.900 100.195 189.945 ;
        RECT 99.430 189.760 100.195 189.900 ;
        RECT 99.430 189.700 99.750 189.760 ;
        RECT 99.905 189.715 100.195 189.760 ;
        RECT 101.270 189.700 101.590 189.960 ;
        RECT 103.570 189.700 103.890 189.960 ;
        RECT 105.040 189.945 105.180 190.100 ;
        RECT 106.330 190.040 106.650 190.100 ;
        RECT 109.090 190.040 109.410 190.100 ;
        RECT 109.550 190.240 109.870 190.300 ;
        RECT 111.865 190.240 112.155 190.285 ;
        RECT 118.610 190.240 118.750 190.440 ;
        RECT 120.145 190.395 120.435 190.440 ;
        RECT 121.510 190.580 121.830 190.640 ;
        RECT 123.365 190.580 123.655 190.625 ;
        RECT 121.510 190.440 123.655 190.580 ;
        RECT 121.510 190.380 121.830 190.440 ;
        RECT 123.365 190.395 123.655 190.440 ;
        RECT 109.550 190.100 112.155 190.240 ;
        RECT 109.550 190.040 109.870 190.100 ;
        RECT 111.865 190.055 112.155 190.100 ;
        RECT 112.860 190.100 118.750 190.240 ;
        RECT 104.965 189.715 105.255 189.945 ;
        RECT 105.870 189.700 106.190 189.960 ;
        RECT 108.630 189.900 108.950 189.960 ;
        RECT 112.860 189.900 113.000 190.100 ;
        RECT 108.630 189.760 113.000 189.900 ;
        RECT 113.245 189.900 113.535 189.945 ;
        RECT 115.530 189.900 115.850 189.960 ;
        RECT 113.245 189.760 115.850 189.900 ;
        RECT 108.630 189.700 108.950 189.760 ;
        RECT 113.245 189.715 113.535 189.760 ;
        RECT 115.530 189.700 115.850 189.760 ;
        RECT 116.465 189.900 116.755 189.945 ;
        RECT 119.225 189.900 119.515 189.945 ;
        RECT 123.825 189.900 124.115 189.945 ;
        RECT 124.270 189.900 124.590 189.960 ;
        RECT 116.465 189.760 124.590 189.900 ;
        RECT 116.465 189.715 116.755 189.760 ;
        RECT 119.225 189.715 119.515 189.760 ;
        RECT 102.665 189.560 102.955 189.605 ;
        RECT 83.880 189.420 102.955 189.560 ;
        RECT 79.280 189.220 79.420 189.420 ;
        RECT 81.950 189.360 82.270 189.420 ;
        RECT 82.425 189.375 82.715 189.420 ;
        RECT 102.665 189.375 102.955 189.420 ;
        RECT 110.820 189.560 111.110 189.605 ;
        RECT 111.390 189.560 111.710 189.620 ;
        RECT 116.540 189.560 116.680 189.715 ;
        RECT 110.820 189.420 116.680 189.560 ;
        RECT 110.820 189.375 111.110 189.420 ;
        RECT 111.390 189.360 111.710 189.420 ;
        RECT 56.650 189.080 57.800 189.220 ;
        RECT 65.020 189.080 79.420 189.220 ;
        RECT 80.570 189.220 80.890 189.280 ;
        RECT 85.185 189.220 85.475 189.265 ;
        RECT 80.570 189.080 85.475 189.220 ;
        RECT 56.650 189.020 56.970 189.080 ;
        RECT 65.020 188.880 65.160 189.080 ;
        RECT 80.570 189.020 80.890 189.080 ;
        RECT 85.185 189.035 85.475 189.080 ;
        RECT 86.105 189.220 86.395 189.265 ;
        RECT 92.530 189.220 92.850 189.280 ;
        RECT 86.105 189.080 92.850 189.220 ;
        RECT 86.105 189.035 86.395 189.080 ;
        RECT 92.530 189.020 92.850 189.080 ;
        RECT 99.890 189.020 100.210 189.280 ;
        RECT 101.730 189.220 102.050 189.280 ;
        RECT 105.870 189.220 106.190 189.280 ;
        RECT 101.730 189.080 106.190 189.220 ;
        RECT 101.730 189.020 102.050 189.080 ;
        RECT 105.870 189.020 106.190 189.080 ;
        RECT 115.530 189.220 115.850 189.280 ;
        RECT 121.140 189.265 121.280 189.760 ;
        RECT 123.825 189.715 124.115 189.760 ;
        RECT 124.270 189.700 124.590 189.760 ;
        RECT 122.430 189.360 122.750 189.620 ;
        RECT 117.845 189.220 118.135 189.265 ;
        RECT 115.530 189.080 118.135 189.220 ;
        RECT 115.530 189.020 115.850 189.080 ;
        RECT 117.845 189.035 118.135 189.080 ;
        RECT 121.065 189.035 121.355 189.265 ;
        RECT 51.220 188.740 65.160 188.880 ;
        RECT 65.390 188.880 65.710 188.940 ;
        RECT 67.245 188.880 67.535 188.925 ;
        RECT 65.390 188.740 67.535 188.880 ;
        RECT 21.690 188.680 22.010 188.740 ;
        RECT 34.570 188.680 34.890 188.740 ;
        RECT 50.670 188.680 50.990 188.740 ;
        RECT 65.390 188.680 65.710 188.740 ;
        RECT 67.245 188.695 67.535 188.740 ;
        RECT 77.365 188.880 77.655 188.925 ;
        RECT 81.965 188.880 82.255 188.925 ;
        RECT 82.410 188.880 82.730 188.940 ;
        RECT 77.365 188.740 82.730 188.880 ;
        RECT 77.365 188.695 77.655 188.740 ;
        RECT 81.965 188.695 82.255 188.740 ;
        RECT 82.410 188.680 82.730 188.740 ;
        RECT 82.870 188.880 83.190 188.940 ;
        RECT 93.450 188.880 93.770 188.940 ;
        RECT 82.870 188.740 93.770 188.880 ;
        RECT 82.870 188.680 83.190 188.740 ;
        RECT 93.450 188.680 93.770 188.740 ;
        RECT 95.290 188.880 95.610 188.940 ;
        RECT 103.570 188.880 103.890 188.940 ;
        RECT 110.930 188.880 111.250 188.940 ;
        RECT 95.290 188.740 111.250 188.880 ;
        RECT 117.920 188.880 118.060 189.035 ;
        RECT 122.430 188.880 122.750 188.940 ;
        RECT 117.920 188.740 122.750 188.880 ;
        RECT 95.290 188.680 95.610 188.740 ;
        RECT 103.570 188.680 103.890 188.740 ;
        RECT 110.930 188.680 111.250 188.740 ;
        RECT 122.430 188.680 122.750 188.740 ;
        RECT 14.260 188.060 126.960 188.540 ;
        RECT 20.310 187.860 20.630 187.920 ;
        RECT 26.290 187.860 26.610 187.920 ;
        RECT 26.765 187.860 27.055 187.905 ;
        RECT 20.310 187.720 21.000 187.860 ;
        RECT 20.310 187.660 20.630 187.720 ;
        RECT 15.710 187.520 16.030 187.580 ;
        RECT 18.025 187.520 18.315 187.565 ;
        RECT 15.710 187.380 18.315 187.520 ;
        RECT 15.710 187.320 16.030 187.380 ;
        RECT 18.025 187.335 18.315 187.380 ;
        RECT 16.185 187.180 16.475 187.225 ;
        RECT 20.860 187.180 21.000 187.720 ;
        RECT 26.290 187.720 27.055 187.860 ;
        RECT 26.290 187.660 26.610 187.720 ;
        RECT 26.765 187.675 27.055 187.720 ;
        RECT 28.590 187.660 28.910 187.920 ;
        RECT 29.970 187.860 30.290 187.920 ;
        RECT 35.950 187.860 36.270 187.920 ;
        RECT 36.425 187.860 36.715 187.905 ;
        RECT 29.970 187.720 36.715 187.860 ;
        RECT 29.970 187.660 30.290 187.720 ;
        RECT 35.950 187.660 36.270 187.720 ;
        RECT 36.425 187.675 36.715 187.720 ;
        RECT 41.010 187.860 41.330 187.920 ;
        RECT 46.545 187.860 46.835 187.905 ;
        RECT 46.990 187.860 47.310 187.920 ;
        RECT 41.010 187.720 44.920 187.860 ;
        RECT 41.010 187.660 41.330 187.720 ;
        RECT 24.910 187.520 25.230 187.580 ;
        RECT 39.170 187.520 39.490 187.580 ;
        RECT 24.910 187.380 39.490 187.520 ;
        RECT 24.910 187.320 25.230 187.380 ;
        RECT 39.170 187.320 39.490 187.380 ;
        RECT 34.125 187.180 34.415 187.225 ;
        RECT 16.185 187.040 19.620 187.180 ;
        RECT 20.860 187.040 34.415 187.180 ;
        RECT 44.780 187.180 44.920 187.720 ;
        RECT 46.545 187.720 47.310 187.860 ;
        RECT 46.545 187.675 46.835 187.720 ;
        RECT 46.990 187.660 47.310 187.720 ;
        RECT 50.210 187.660 50.530 187.920 ;
        RECT 51.130 187.860 51.450 187.920 ;
        RECT 52.065 187.860 52.355 187.905 ;
        RECT 86.565 187.860 86.855 187.905 ;
        RECT 87.010 187.860 87.330 187.920 ;
        RECT 100.365 187.860 100.655 187.905 ;
        RECT 51.130 187.720 57.340 187.860 ;
        RECT 51.130 187.660 51.450 187.720 ;
        RECT 52.065 187.675 52.355 187.720 ;
        RECT 45.610 187.520 45.930 187.580 ;
        RECT 49.750 187.520 50.070 187.580 ;
        RECT 56.650 187.520 56.970 187.580 ;
        RECT 45.610 187.380 50.070 187.520 ;
        RECT 45.610 187.320 45.930 187.380 ;
        RECT 49.750 187.320 50.070 187.380 ;
        RECT 52.600 187.380 56.970 187.520 ;
        RECT 57.200 187.520 57.340 187.720 ;
        RECT 86.565 187.720 87.330 187.860 ;
        RECT 86.565 187.675 86.855 187.720 ;
        RECT 87.010 187.660 87.330 187.720 ;
        RECT 87.560 187.720 100.655 187.860 ;
        RECT 61.710 187.520 62.030 187.580 ;
        RECT 57.200 187.380 62.030 187.520 ;
        RECT 48.370 187.180 48.690 187.240 ;
        RECT 44.780 187.040 48.140 187.180 ;
        RECT 16.185 186.995 16.475 187.040 ;
        RECT 17.105 186.655 17.395 186.885 ;
        RECT 17.180 186.500 17.320 186.655 ;
        RECT 17.550 186.640 17.870 186.900 ;
        RECT 18.485 186.840 18.775 186.885 ;
        RECT 18.930 186.840 19.250 186.900 ;
        RECT 19.480 186.885 19.620 187.040 ;
        RECT 34.125 186.995 34.415 187.040 ;
        RECT 18.485 186.700 19.250 186.840 ;
        RECT 18.485 186.655 18.775 186.700 ;
        RECT 18.930 186.640 19.250 186.700 ;
        RECT 19.405 186.655 19.695 186.885 ;
        RECT 20.310 186.640 20.630 186.900 ;
        RECT 21.690 186.640 22.010 186.900 ;
        RECT 24.910 186.840 25.230 186.900 ;
        RECT 27.670 186.840 27.990 186.900 ;
        RECT 24.910 186.700 27.990 186.840 ;
        RECT 24.910 186.640 25.230 186.700 ;
        RECT 27.670 186.640 27.990 186.700 ;
        RECT 28.145 186.840 28.435 186.885 ;
        RECT 28.590 186.840 28.910 186.900 ;
        RECT 33.650 186.885 33.970 186.900 ;
        RECT 28.145 186.700 28.910 186.840 ;
        RECT 28.145 186.655 28.435 186.700 ;
        RECT 28.590 186.640 28.910 186.700 ;
        RECT 29.065 186.655 29.355 186.885 ;
        RECT 33.650 186.655 33.985 186.885 ;
        RECT 34.585 186.840 34.875 186.885 ;
        RECT 44.690 186.840 45.010 186.900 ;
        RECT 34.585 186.700 45.010 186.840 ;
        RECT 34.585 186.655 34.875 186.700 ;
        RECT 18.010 186.500 18.330 186.560 ;
        RECT 17.180 186.360 18.330 186.500 ;
        RECT 18.010 186.300 18.330 186.360 ;
        RECT 20.770 186.300 21.090 186.560 ;
        RECT 21.245 186.500 21.535 186.545 ;
        RECT 25.845 186.500 26.135 186.545 ;
        RECT 26.750 186.500 27.070 186.560 ;
        RECT 21.245 186.360 25.600 186.500 ;
        RECT 21.245 186.315 21.535 186.360 ;
        RECT 22.625 186.160 22.915 186.205 ;
        RECT 24.450 186.160 24.770 186.220 ;
        RECT 22.625 186.020 24.770 186.160 ;
        RECT 25.460 186.160 25.600 186.360 ;
        RECT 25.845 186.360 27.070 186.500 ;
        RECT 29.140 186.500 29.280 186.655 ;
        RECT 33.650 186.640 33.970 186.655 ;
        RECT 44.690 186.640 45.010 186.700 ;
        RECT 45.150 186.640 45.470 186.900 ;
        RECT 45.610 186.640 45.930 186.900 ;
        RECT 46.990 186.640 47.310 186.900 ;
        RECT 48.000 186.885 48.140 187.040 ;
        RECT 48.370 187.040 51.360 187.180 ;
        RECT 48.370 186.980 48.690 187.040 ;
        RECT 47.925 186.655 48.215 186.885 ;
        RECT 49.290 186.840 49.610 186.900 ;
        RECT 51.220 186.885 51.360 187.040 ;
        RECT 49.765 186.840 50.055 186.885 ;
        RECT 49.290 186.700 50.055 186.840 ;
        RECT 49.290 186.640 49.610 186.700 ;
        RECT 49.765 186.655 50.055 186.700 ;
        RECT 51.145 186.655 51.435 186.885 ;
        RECT 41.010 186.500 41.330 186.560 ;
        RECT 29.140 186.360 41.330 186.500 ;
        RECT 25.845 186.315 26.135 186.360 ;
        RECT 26.750 186.300 27.070 186.360 ;
        RECT 41.010 186.300 41.330 186.360 ;
        RECT 43.785 186.500 44.075 186.545 ;
        RECT 46.070 186.500 46.390 186.560 ;
        RECT 52.600 186.545 52.740 187.380 ;
        RECT 56.650 187.320 56.970 187.380 ;
        RECT 61.710 187.320 62.030 187.380 ;
        RECT 69.545 187.520 69.835 187.565 ;
        RECT 87.560 187.520 87.700 187.720 ;
        RECT 100.365 187.675 100.655 187.720 ;
        RECT 101.730 187.860 102.050 187.920 ;
        RECT 102.665 187.860 102.955 187.905 ;
        RECT 101.730 187.720 102.955 187.860 ;
        RECT 101.730 187.660 102.050 187.720 ;
        RECT 102.665 187.675 102.955 187.720 ;
        RECT 108.170 187.860 108.490 187.920 ;
        RECT 110.010 187.860 110.330 187.920 ;
        RECT 108.170 187.720 110.330 187.860 ;
        RECT 108.170 187.660 108.490 187.720 ;
        RECT 110.010 187.660 110.330 187.720 ;
        RECT 110.470 187.860 110.790 187.920 ;
        RECT 112.310 187.860 112.630 187.920 ;
        RECT 110.470 187.720 112.630 187.860 ;
        RECT 110.470 187.660 110.790 187.720 ;
        RECT 112.310 187.660 112.630 187.720 ;
        RECT 124.745 187.860 125.035 187.905 ;
        RECT 131.170 187.860 131.490 187.920 ;
        RECT 124.745 187.720 131.490 187.860 ;
        RECT 124.745 187.675 125.035 187.720 ;
        RECT 131.170 187.660 131.490 187.720 ;
        RECT 69.545 187.380 87.700 187.520 ;
        RECT 87.930 187.520 88.250 187.580 ;
        RECT 90.230 187.520 90.550 187.580 ;
        RECT 87.930 187.380 90.550 187.520 ;
        RECT 69.545 187.335 69.835 187.380 ;
        RECT 87.930 187.320 88.250 187.380 ;
        RECT 90.230 187.320 90.550 187.380 ;
        RECT 98.510 187.520 98.830 187.580 ;
        RECT 103.110 187.520 103.430 187.580 ;
        RECT 98.510 187.380 103.430 187.520 ;
        RECT 98.510 187.320 98.830 187.380 ;
        RECT 103.110 187.320 103.430 187.380 ;
        RECT 105.410 187.320 105.730 187.580 ;
        RECT 105.870 187.520 106.190 187.580 ;
        RECT 111.405 187.520 111.695 187.565 ;
        RECT 105.870 187.380 111.695 187.520 ;
        RECT 105.870 187.320 106.190 187.380 ;
        RECT 111.405 187.335 111.695 187.380 ;
        RECT 55.270 187.180 55.590 187.240 ;
        RECT 55.270 187.040 58.720 187.180 ;
        RECT 55.270 186.980 55.590 187.040 ;
        RECT 53.445 186.840 53.735 186.885 ;
        RECT 54.350 186.840 54.670 186.900 ;
        RECT 54.825 186.840 55.115 186.885 ;
        RECT 53.445 186.700 55.115 186.840 ;
        RECT 53.445 186.655 53.735 186.700 ;
        RECT 54.350 186.640 54.670 186.700 ;
        RECT 54.825 186.655 55.115 186.700 ;
        RECT 55.730 186.640 56.050 186.900 ;
        RECT 56.280 186.885 56.420 187.040 ;
        RECT 58.580 186.900 58.720 187.040 ;
        RECT 67.690 186.980 68.010 187.240 ;
        RECT 68.625 187.180 68.915 187.225 ;
        RECT 71.370 187.180 71.690 187.240 ;
        RECT 79.650 187.180 79.970 187.240 ;
        RECT 68.625 187.040 71.690 187.180 ;
        RECT 68.625 186.995 68.915 187.040 ;
        RECT 71.370 186.980 71.690 187.040 ;
        RECT 71.920 187.040 79.970 187.180 ;
        RECT 56.205 186.655 56.495 186.885 ;
        RECT 56.650 186.640 56.970 186.900 ;
        RECT 58.490 186.840 58.810 186.900 ;
        RECT 69.530 186.840 69.850 186.900 ;
        RECT 70.005 186.840 70.295 186.885 ;
        RECT 71.920 186.840 72.060 187.040 ;
        RECT 79.650 186.980 79.970 187.040 ;
        RECT 83.790 186.980 84.110 187.240 ;
        RECT 86.550 187.180 86.870 187.240 ;
        RECT 84.340 187.040 86.870 187.180 ;
        RECT 58.490 186.700 67.920 186.840 ;
        RECT 58.490 186.640 58.810 186.700 ;
        RECT 52.525 186.500 52.815 186.545 ;
        RECT 43.785 186.360 45.380 186.500 ;
        RECT 43.785 186.315 44.075 186.360 ;
        RECT 45.240 186.220 45.380 186.360 ;
        RECT 46.070 186.360 52.815 186.500 ;
        RECT 46.070 186.300 46.390 186.360 ;
        RECT 52.525 186.315 52.815 186.360 ;
        RECT 53.890 186.500 54.210 186.560 ;
        RECT 58.045 186.500 58.335 186.545 ;
        RECT 53.890 186.360 58.335 186.500 ;
        RECT 53.890 186.300 54.210 186.360 ;
        RECT 58.045 186.315 58.335 186.360 ;
        RECT 66.785 186.500 67.075 186.545 ;
        RECT 67.230 186.500 67.550 186.560 ;
        RECT 66.785 186.360 67.550 186.500 ;
        RECT 67.780 186.500 67.920 186.700 ;
        RECT 69.530 186.700 72.060 186.840 ;
        RECT 73.670 186.840 73.990 186.900 ;
        RECT 80.570 186.840 80.890 186.900 ;
        RECT 73.670 186.700 80.890 186.840 ;
        RECT 69.530 186.640 69.850 186.700 ;
        RECT 70.005 186.655 70.295 186.700 ;
        RECT 73.670 186.640 73.990 186.700 ;
        RECT 80.570 186.640 80.890 186.700 ;
        RECT 83.345 186.840 83.635 186.885 ;
        RECT 84.340 186.840 84.480 187.040 ;
        RECT 86.550 186.980 86.870 187.040 ;
        RECT 89.325 187.180 89.615 187.225 ;
        RECT 91.150 187.180 91.470 187.240 ;
        RECT 92.530 187.180 92.850 187.240 ;
        RECT 101.730 187.180 102.050 187.240 ;
        RECT 112.770 187.180 113.090 187.240 ;
        RECT 89.325 187.040 92.850 187.180 ;
        RECT 89.325 186.995 89.615 187.040 ;
        RECT 91.150 186.980 91.470 187.040 ;
        RECT 92.530 186.980 92.850 187.040 ;
        RECT 97.680 187.040 102.050 187.180 ;
        RECT 83.345 186.700 84.480 186.840 ;
        RECT 83.345 186.655 83.635 186.700 ;
        RECT 85.170 186.640 85.490 186.900 ;
        RECT 85.630 186.640 85.950 186.900 ;
        RECT 97.680 186.885 97.820 187.040 ;
        RECT 101.730 186.980 102.050 187.040 ;
        RECT 105.040 187.040 113.090 187.180 ;
        RECT 97.605 186.655 97.895 186.885 ;
        RECT 98.510 186.640 98.830 186.900 ;
        RECT 98.970 186.640 99.290 186.900 ;
        RECT 99.445 186.840 99.735 186.885 ;
        RECT 99.890 186.840 100.210 186.900 ;
        RECT 105.040 186.885 105.180 187.040 ;
        RECT 106.880 186.885 107.020 187.040 ;
        RECT 112.770 186.980 113.090 187.040 ;
        RECT 99.445 186.700 100.210 186.840 ;
        RECT 99.445 186.655 99.735 186.700 ;
        RECT 99.890 186.640 100.210 186.700 ;
        RECT 103.585 186.655 103.875 186.885 ;
        RECT 104.965 186.655 105.255 186.885 ;
        RECT 106.805 186.655 107.095 186.885 ;
        RECT 110.025 186.840 110.315 186.885 ;
        RECT 110.470 186.840 110.790 186.900 ;
        RECT 110.025 186.700 110.790 186.840 ;
        RECT 110.025 186.655 110.315 186.700 ;
        RECT 71.370 186.500 71.690 186.560 ;
        RECT 100.365 186.500 100.655 186.545 ;
        RECT 100.810 186.500 101.130 186.560 ;
        RECT 67.780 186.360 86.320 186.500 ;
        RECT 66.785 186.315 67.075 186.360 ;
        RECT 67.230 186.300 67.550 186.360 ;
        RECT 71.370 186.300 71.690 186.360 ;
        RECT 86.180 186.220 86.320 186.360 ;
        RECT 100.365 186.360 101.130 186.500 ;
        RECT 103.660 186.500 103.800 186.655 ;
        RECT 110.470 186.640 110.790 186.700 ;
        RECT 110.945 186.840 111.235 186.885 ;
        RECT 114.165 186.840 114.455 186.885 ;
        RECT 110.945 186.700 114.455 186.840 ;
        RECT 110.945 186.655 111.235 186.700 ;
        RECT 114.165 186.655 114.455 186.700 ;
        RECT 105.425 186.500 105.715 186.545 ;
        RECT 105.870 186.500 106.190 186.560 ;
        RECT 103.660 186.360 106.190 186.500 ;
        RECT 100.365 186.315 100.655 186.360 ;
        RECT 100.810 186.300 101.130 186.360 ;
        RECT 105.425 186.315 105.715 186.360 ;
        RECT 105.870 186.300 106.190 186.360 ;
        RECT 106.345 186.500 106.635 186.545 ;
        RECT 109.090 186.500 109.410 186.560 ;
        RECT 111.020 186.500 111.160 186.655 ;
        RECT 123.810 186.640 124.130 186.900 ;
        RECT 106.345 186.360 111.160 186.500 ;
        RECT 111.850 186.500 112.170 186.560 ;
        RECT 112.325 186.500 112.615 186.545 ;
        RECT 111.850 186.360 112.615 186.500 ;
        RECT 106.345 186.315 106.635 186.360 ;
        RECT 28.590 186.160 28.910 186.220 ;
        RECT 25.460 186.020 28.910 186.160 ;
        RECT 22.625 185.975 22.915 186.020 ;
        RECT 24.450 185.960 24.770 186.020 ;
        RECT 28.590 185.960 28.910 186.020 ;
        RECT 33.650 186.160 33.970 186.220 ;
        RECT 41.930 186.160 42.250 186.220 ;
        RECT 44.245 186.160 44.535 186.205 ;
        RECT 33.650 186.020 44.535 186.160 ;
        RECT 33.650 185.960 33.970 186.020 ;
        RECT 41.930 185.960 42.250 186.020 ;
        RECT 44.245 185.975 44.535 186.020 ;
        RECT 45.150 185.960 45.470 186.220 ;
        RECT 54.350 185.960 54.670 186.220 ;
        RECT 56.190 186.160 56.510 186.220 ;
        RECT 57.585 186.160 57.875 186.205 ;
        RECT 56.190 186.020 57.875 186.160 ;
        RECT 56.190 185.960 56.510 186.020 ;
        RECT 57.585 185.975 57.875 186.020 ;
        RECT 60.330 186.160 60.650 186.220 ;
        RECT 82.870 186.160 83.190 186.220 ;
        RECT 60.330 186.020 83.190 186.160 ;
        RECT 60.330 185.960 60.650 186.020 ;
        RECT 82.870 185.960 83.190 186.020 ;
        RECT 86.090 186.160 86.410 186.220 ;
        RECT 87.025 186.160 87.315 186.205 ;
        RECT 86.090 186.020 87.315 186.160 ;
        RECT 86.090 185.960 86.410 186.020 ;
        RECT 87.025 185.975 87.315 186.020 ;
        RECT 98.065 186.160 98.355 186.205 ;
        RECT 98.510 186.160 98.830 186.220 ;
        RECT 98.065 186.020 98.830 186.160 ;
        RECT 98.065 185.975 98.355 186.020 ;
        RECT 98.510 185.960 98.830 186.020 ;
        RECT 101.270 185.960 101.590 186.220 ;
        RECT 104.505 186.160 104.795 186.205 ;
        RECT 106.420 186.160 106.560 186.315 ;
        RECT 109.090 186.300 109.410 186.360 ;
        RECT 111.850 186.300 112.170 186.360 ;
        RECT 112.325 186.315 112.615 186.360 ;
        RECT 104.505 186.020 106.560 186.160 ;
        RECT 108.170 186.160 108.490 186.220 ;
        RECT 110.485 186.160 110.775 186.205 ;
        RECT 108.170 186.020 110.775 186.160 ;
        RECT 104.505 185.975 104.795 186.020 ;
        RECT 108.170 185.960 108.490 186.020 ;
        RECT 110.485 185.975 110.775 186.020 ;
        RECT 14.260 185.340 126.960 185.820 ;
        RECT 18.930 185.140 19.250 185.200 ;
        RECT 20.325 185.140 20.615 185.185 ;
        RECT 26.750 185.140 27.070 185.200 ;
        RECT 18.930 185.000 27.070 185.140 ;
        RECT 18.930 184.940 19.250 185.000 ;
        RECT 20.325 184.955 20.615 185.000 ;
        RECT 26.750 184.940 27.070 185.000 ;
        RECT 39.630 185.140 39.950 185.200 ;
        RECT 40.565 185.140 40.855 185.185 ;
        RECT 39.630 185.000 40.855 185.140 ;
        RECT 39.630 184.940 39.950 185.000 ;
        RECT 40.565 184.955 40.855 185.000 ;
        RECT 41.470 185.140 41.790 185.200 ;
        RECT 46.530 185.140 46.850 185.200 ;
        RECT 47.925 185.140 48.215 185.185 ;
        RECT 41.470 185.000 42.160 185.140 ;
        RECT 41.470 184.940 41.790 185.000 ;
        RECT 27.210 184.600 27.530 184.860 ;
        RECT 35.490 184.600 35.810 184.860 ;
        RECT 42.020 184.845 42.160 185.000 ;
        RECT 46.530 185.000 48.215 185.140 ;
        RECT 46.530 184.940 46.850 185.000 ;
        RECT 47.925 184.955 48.215 185.000 ;
        RECT 50.670 185.140 50.990 185.200 ;
        RECT 53.430 185.140 53.750 185.200 ;
        RECT 54.410 185.140 54.700 185.185 ;
        RECT 50.670 185.000 53.200 185.140 ;
        RECT 50.670 184.940 50.990 185.000 ;
        RECT 39.185 184.800 39.475 184.845 ;
        RECT 37.460 184.660 39.475 184.800 ;
        RECT 16.185 184.275 16.475 184.505 ;
        RECT 26.765 184.460 27.055 184.505 ;
        RECT 29.510 184.460 29.830 184.520 ;
        RECT 37.460 184.460 37.600 184.660 ;
        RECT 39.185 184.615 39.475 184.660 ;
        RECT 41.945 184.615 42.235 184.845 ;
        RECT 45.610 184.800 45.930 184.860 ;
        RECT 51.590 184.800 51.910 184.860 ;
        RECT 42.940 184.660 45.930 184.800 ;
        RECT 26.765 184.320 29.830 184.460 ;
        RECT 26.765 184.275 27.055 184.320 ;
        RECT 16.260 183.780 16.400 184.275 ;
        RECT 29.510 184.260 29.830 184.320 ;
        RECT 35.810 184.320 37.600 184.460 ;
        RECT 28.590 184.120 28.910 184.180 ;
        RECT 35.810 184.120 35.950 184.320 ;
        RECT 38.250 184.260 38.570 184.520 ;
        RECT 38.710 184.260 39.030 184.520 ;
        RECT 39.630 184.460 39.950 184.520 ;
        RECT 41.485 184.460 41.775 184.505 ;
        RECT 39.630 184.320 41.775 184.460 ;
        RECT 39.630 184.260 39.950 184.320 ;
        RECT 41.485 184.275 41.775 184.320 ;
        RECT 28.590 183.980 35.950 184.120 ;
        RECT 36.870 184.120 37.190 184.180 ;
        RECT 40.105 184.120 40.395 184.165 ;
        RECT 36.870 183.980 40.395 184.120 ;
        RECT 41.560 184.120 41.700 184.275 ;
        RECT 42.390 184.260 42.710 184.520 ;
        RECT 42.940 184.120 43.080 184.660 ;
        RECT 45.610 184.600 45.930 184.660 ;
        RECT 50.760 184.660 51.910 184.800 ;
        RECT 43.370 184.505 43.690 184.520 ;
        RECT 43.325 184.275 43.690 184.505 ;
        RECT 44.245 184.275 44.535 184.505 ;
        RECT 44.690 184.460 45.010 184.520 ;
        RECT 46.070 184.460 46.390 184.520 ;
        RECT 44.690 184.320 46.390 184.460 ;
        RECT 43.370 184.260 43.690 184.275 ;
        RECT 44.320 184.120 44.460 184.275 ;
        RECT 44.690 184.260 45.010 184.320 ;
        RECT 46.070 184.260 46.390 184.320 ;
        RECT 46.530 184.260 46.850 184.520 ;
        RECT 47.450 184.260 47.770 184.520 ;
        RECT 47.910 184.460 48.230 184.520 ;
        RECT 48.845 184.460 49.135 184.505 ;
        RECT 49.290 184.460 49.610 184.520 ;
        RECT 50.760 184.505 50.900 184.660 ;
        RECT 51.590 184.600 51.910 184.660 ;
        RECT 52.510 184.600 52.830 184.860 ;
        RECT 53.060 184.800 53.200 185.000 ;
        RECT 53.430 185.000 54.700 185.140 ;
        RECT 53.430 184.940 53.750 185.000 ;
        RECT 54.410 184.955 54.700 185.000 ;
        RECT 67.705 185.140 67.995 185.185 ;
        RECT 68.150 185.140 68.470 185.200 ;
        RECT 67.705 185.000 68.470 185.140 ;
        RECT 67.705 184.955 67.995 185.000 ;
        RECT 68.150 184.940 68.470 185.000 ;
        RECT 70.925 185.140 71.215 185.185 ;
        RECT 71.830 185.140 72.150 185.200 ;
        RECT 70.925 185.000 72.150 185.140 ;
        RECT 70.925 184.955 71.215 185.000 ;
        RECT 71.830 184.940 72.150 185.000 ;
        RECT 72.840 185.000 82.640 185.140 ;
        RECT 57.585 184.800 57.875 184.845 ;
        RECT 53.060 184.660 57.875 184.800 ;
        RECT 47.910 184.320 49.610 184.460 ;
        RECT 47.910 184.260 48.230 184.320 ;
        RECT 48.845 184.275 49.135 184.320 ;
        RECT 49.290 184.260 49.610 184.320 ;
        RECT 50.685 184.275 50.975 184.505 ;
        RECT 51.145 184.460 51.435 184.505 ;
        RECT 54.810 184.460 55.130 184.520 ;
        RECT 57.200 184.505 57.340 184.660 ;
        RECT 57.585 184.615 57.875 184.660 ;
        RECT 60.330 184.600 60.650 184.860 ;
        RECT 69.530 184.800 69.850 184.860 ;
        RECT 72.840 184.800 72.980 185.000 ;
        RECT 82.500 184.860 82.640 185.000 ;
        RECT 83.805 184.955 84.095 185.185 ;
        RECT 84.250 185.140 84.570 185.200 ;
        RECT 112.325 185.140 112.615 185.185 ;
        RECT 112.770 185.140 113.090 185.200 ;
        RECT 84.250 185.000 85.860 185.140 ;
        RECT 63.640 184.660 69.850 184.800 ;
        RECT 58.950 184.505 59.270 184.520 ;
        RECT 57.125 184.460 57.415 184.505 ;
        RECT 51.145 184.320 55.130 184.460 ;
        RECT 57.015 184.320 57.415 184.460 ;
        RECT 51.145 184.275 51.435 184.320 ;
        RECT 54.810 184.260 55.130 184.320 ;
        RECT 57.125 184.275 57.415 184.320 ;
        RECT 58.950 184.275 59.485 184.505 ;
        RECT 58.950 184.260 59.270 184.275 ;
        RECT 59.870 184.260 60.190 184.520 ;
        RECT 60.790 184.260 61.110 184.520 ;
        RECT 63.640 184.505 63.780 184.660 ;
        RECT 61.725 184.460 62.015 184.505 ;
        RECT 63.565 184.460 63.855 184.505 ;
        RECT 61.725 184.320 63.855 184.460 ;
        RECT 61.725 184.275 62.015 184.320 ;
        RECT 63.565 184.275 63.855 184.320 ;
        RECT 64.470 184.260 64.790 184.520 ;
        RECT 65.390 184.260 65.710 184.520 ;
        RECT 66.400 184.505 66.540 184.660 ;
        RECT 69.530 184.600 69.850 184.660 ;
        RECT 72.380 184.660 72.980 184.800 ;
        RECT 72.380 184.520 72.520 184.660 ;
        RECT 81.950 184.600 82.270 184.860 ;
        RECT 82.410 184.600 82.730 184.860 ;
        RECT 66.325 184.275 66.615 184.505 ;
        RECT 66.785 184.460 67.075 184.505 ;
        RECT 68.150 184.460 68.470 184.520 ;
        RECT 66.785 184.320 68.470 184.460 ;
        RECT 66.785 184.275 67.075 184.320 ;
        RECT 68.150 184.260 68.470 184.320 ;
        RECT 68.625 184.275 68.915 184.505 ;
        RECT 69.070 184.460 69.390 184.520 ;
        RECT 70.005 184.460 70.295 184.505 ;
        RECT 69.070 184.320 70.295 184.460 ;
        RECT 41.560 183.980 43.080 184.120 ;
        RECT 43.860 183.980 44.460 184.120 ;
        RECT 45.150 184.120 45.470 184.180 ;
        RECT 53.890 184.120 54.210 184.180 ;
        RECT 45.150 183.980 54.210 184.120 ;
        RECT 28.590 183.920 28.910 183.980 ;
        RECT 36.870 183.920 37.190 183.980 ;
        RECT 40.105 183.935 40.395 183.980 ;
        RECT 29.050 183.780 29.370 183.840 ;
        RECT 16.260 183.640 29.370 183.780 ;
        RECT 29.050 183.580 29.370 183.640 ;
        RECT 34.570 183.780 34.890 183.840 ;
        RECT 35.950 183.780 36.270 183.840 ;
        RECT 34.570 183.640 43.080 183.780 ;
        RECT 34.570 183.580 34.890 183.640 ;
        RECT 35.950 183.580 36.270 183.640 ;
        RECT 17.090 183.240 17.410 183.500 ;
        RECT 20.770 183.440 21.090 183.500 ;
        RECT 36.410 183.440 36.730 183.500 ;
        RECT 20.770 183.300 36.730 183.440 ;
        RECT 20.770 183.240 21.090 183.300 ;
        RECT 36.410 183.240 36.730 183.300 ;
        RECT 36.870 183.440 37.190 183.500 ;
        RECT 37.345 183.440 37.635 183.485 ;
        RECT 36.870 183.300 37.635 183.440 ;
        RECT 36.870 183.240 37.190 183.300 ;
        RECT 37.345 183.255 37.635 183.300 ;
        RECT 38.250 183.440 38.570 183.500 ;
        RECT 39.170 183.440 39.490 183.500 ;
        RECT 42.390 183.440 42.710 183.500 ;
        RECT 38.250 183.300 42.710 183.440 ;
        RECT 42.940 183.440 43.080 183.640 ;
        RECT 43.860 183.440 44.000 183.980 ;
        RECT 45.150 183.920 45.470 183.980 ;
        RECT 53.890 183.920 54.210 183.980 ;
        RECT 54.350 184.120 54.670 184.180 ;
        RECT 55.730 184.120 56.050 184.180 ;
        RECT 58.505 184.120 58.795 184.165 ;
        RECT 54.350 183.980 58.795 184.120 ;
        RECT 54.350 183.920 54.670 183.980 ;
        RECT 55.730 183.920 56.050 183.980 ;
        RECT 58.505 183.935 58.795 183.980 ;
        RECT 64.025 184.120 64.315 184.165 ;
        RECT 68.700 184.120 68.840 184.275 ;
        RECT 69.070 184.260 69.390 184.320 ;
        RECT 70.005 184.275 70.295 184.320 ;
        RECT 72.290 184.260 72.610 184.520 ;
        RECT 72.750 184.260 73.070 184.520 ;
        RECT 80.570 184.505 80.890 184.520 ;
        RECT 82.870 184.505 83.190 184.520 ;
        RECT 80.570 184.460 80.910 184.505 ;
        RECT 80.410 184.320 80.910 184.460 ;
        RECT 80.570 184.275 80.910 184.320 ;
        RECT 81.050 184.275 81.340 184.505 ;
        RECT 82.870 184.460 83.200 184.505 ;
        RECT 83.880 184.460 84.020 184.955 ;
        RECT 84.250 184.940 84.570 185.000 ;
        RECT 85.720 184.845 85.860 185.000 ;
        RECT 91.240 185.000 95.980 185.140 ;
        RECT 91.240 184.860 91.380 185.000 ;
        RECT 85.640 184.615 85.930 184.845 ;
        RECT 86.105 184.800 86.395 184.845 ;
        RECT 87.470 184.800 87.790 184.860 ;
        RECT 86.105 184.660 87.790 184.800 ;
        RECT 86.105 184.615 86.395 184.660 ;
        RECT 87.470 184.600 87.790 184.660 ;
        RECT 90.230 184.600 90.550 184.860 ;
        RECT 91.150 184.600 91.470 184.860 ;
        RECT 94.830 184.800 95.150 184.860 ;
        RECT 91.700 184.660 95.520 184.800 ;
        RECT 84.955 184.460 85.245 184.505 ;
        RECT 82.870 184.320 83.385 184.460 ;
        RECT 83.880 184.320 85.245 184.460 ;
        RECT 82.870 184.275 83.200 184.320 ;
        RECT 84.955 184.275 85.245 184.320 ;
        RECT 80.570 184.260 80.890 184.275 ;
        RECT 64.025 183.980 68.840 184.120 ;
        RECT 71.385 184.120 71.675 184.165 ;
        RECT 73.670 184.120 73.990 184.180 ;
        RECT 71.385 183.980 73.990 184.120 ;
        RECT 64.025 183.935 64.315 183.980 ;
        RECT 71.385 183.935 71.675 183.980 ;
        RECT 73.670 183.920 73.990 183.980 ;
        RECT 79.190 184.120 79.510 184.180 ;
        RECT 81.120 184.120 81.260 184.275 ;
        RECT 82.870 184.260 83.190 184.275 ;
        RECT 86.550 184.260 86.870 184.520 ;
        RECT 88.405 184.275 88.695 184.505 ;
        RECT 79.190 183.980 81.260 184.120 ;
        RECT 84.265 184.120 84.555 184.165 ;
        RECT 86.090 184.120 86.410 184.180 ;
        RECT 88.480 184.120 88.620 184.275 ;
        RECT 89.310 184.260 89.630 184.520 ;
        RECT 89.785 184.275 90.075 184.505 ;
        RECT 90.320 184.460 90.460 184.600 ;
        RECT 91.700 184.460 91.840 184.660 ;
        RECT 94.830 184.600 95.150 184.660 ;
        RECT 90.320 184.320 91.840 184.460 ;
        RECT 92.070 184.460 92.390 184.520 ;
        RECT 93.925 184.460 94.215 184.505 ;
        RECT 94.370 184.460 94.690 184.520 ;
        RECT 95.380 184.505 95.520 184.660 ;
        RECT 92.070 184.320 92.760 184.460 ;
        RECT 84.265 183.980 86.410 184.120 ;
        RECT 79.190 183.920 79.510 183.980 ;
        RECT 84.265 183.935 84.555 183.980 ;
        RECT 86.090 183.920 86.410 183.980 ;
        RECT 86.640 183.980 88.620 184.120 ;
        RECT 52.065 183.780 52.355 183.825 ;
        RECT 60.330 183.780 60.650 183.840 ;
        RECT 52.065 183.640 60.650 183.780 ;
        RECT 52.065 183.595 52.355 183.640 ;
        RECT 42.940 183.300 44.000 183.440 ;
        RECT 44.230 183.440 44.550 183.500 ;
        RECT 46.990 183.440 47.310 183.500 ;
        RECT 54.440 183.485 54.580 183.640 ;
        RECT 60.330 183.580 60.650 183.640 ;
        RECT 65.865 183.780 66.155 183.825 ;
        RECT 66.770 183.780 67.090 183.840 ;
        RECT 65.865 183.640 67.090 183.780 ;
        RECT 65.865 183.595 66.155 183.640 ;
        RECT 66.770 183.580 67.090 183.640 ;
        RECT 69.085 183.595 69.375 183.825 ;
        RECT 44.230 183.300 47.310 183.440 ;
        RECT 38.250 183.240 38.570 183.300 ;
        RECT 39.170 183.240 39.490 183.300 ;
        RECT 42.390 183.240 42.710 183.300 ;
        RECT 44.230 183.240 44.550 183.300 ;
        RECT 46.990 183.240 47.310 183.300 ;
        RECT 54.365 183.255 54.655 183.485 ;
        RECT 55.270 183.240 55.590 183.500 ;
        RECT 56.190 183.240 56.510 183.500 ;
        RECT 66.310 183.440 66.630 183.500 ;
        RECT 69.160 183.440 69.300 183.595 ;
        RECT 69.530 183.580 69.850 183.840 ;
        RECT 80.570 183.780 80.890 183.840 ;
        RECT 86.640 183.780 86.780 183.980 ;
        RECT 80.570 183.640 86.780 183.780 ;
        RECT 87.930 183.780 88.250 183.840 ;
        RECT 88.405 183.780 88.695 183.825 ;
        RECT 87.930 183.640 88.695 183.780 ;
        RECT 80.570 183.580 80.890 183.640 ;
        RECT 87.930 183.580 88.250 183.640 ;
        RECT 88.405 183.595 88.695 183.640 ;
        RECT 66.310 183.300 69.300 183.440 ;
        RECT 66.310 183.240 66.630 183.300 ;
        RECT 71.830 183.240 72.150 183.500 ;
        RECT 81.950 183.440 82.270 183.500 ;
        RECT 84.710 183.440 85.030 183.500 ;
        RECT 81.950 183.300 85.030 183.440 ;
        RECT 81.950 183.240 82.270 183.300 ;
        RECT 84.710 183.240 85.030 183.300 ;
        RECT 87.010 183.440 87.330 183.500 ;
        RECT 87.485 183.440 87.775 183.485 ;
        RECT 87.010 183.300 87.775 183.440 ;
        RECT 89.860 183.440 90.000 184.275 ;
        RECT 92.070 184.260 92.390 184.320 ;
        RECT 92.620 184.165 92.760 184.320 ;
        RECT 93.925 184.320 94.690 184.460 ;
        RECT 93.925 184.275 94.215 184.320 ;
        RECT 94.370 184.260 94.690 184.320 ;
        RECT 95.305 184.275 95.595 184.505 ;
        RECT 95.840 184.460 95.980 185.000 ;
        RECT 112.325 185.000 113.090 185.140 ;
        RECT 112.325 184.955 112.615 185.000 ;
        RECT 112.770 184.940 113.090 185.000 ;
        RECT 96.225 184.800 96.515 184.845 ;
        RECT 98.970 184.800 99.290 184.860 ;
        RECT 101.270 184.800 101.590 184.860 ;
        RECT 108.630 184.800 108.950 184.860 ;
        RECT 96.225 184.660 100.120 184.800 ;
        RECT 96.225 184.615 96.515 184.660 ;
        RECT 98.970 184.600 99.290 184.660 ;
        RECT 97.145 184.460 97.435 184.505 ;
        RECT 95.840 184.320 97.435 184.460 ;
        RECT 97.145 184.275 97.435 184.320 ;
        RECT 98.050 184.260 98.370 184.520 ;
        RECT 98.510 184.260 98.830 184.520 ;
        RECT 99.980 184.505 100.120 184.660 ;
        RECT 100.900 184.660 104.260 184.800 ;
        RECT 100.900 184.505 101.040 184.660 ;
        RECT 101.270 184.600 101.590 184.660 ;
        RECT 99.905 184.275 100.195 184.505 ;
        RECT 100.825 184.275 101.115 184.505 ;
        RECT 101.730 184.460 102.050 184.520 ;
        RECT 104.120 184.505 104.260 184.660 ;
        RECT 108.630 184.660 109.780 184.800 ;
        RECT 108.630 184.600 108.950 184.660 ;
        RECT 103.585 184.460 103.875 184.505 ;
        RECT 101.730 184.320 103.875 184.460 ;
        RECT 101.730 184.260 102.050 184.320 ;
        RECT 103.585 184.275 103.875 184.320 ;
        RECT 104.045 184.275 104.335 184.505 ;
        RECT 109.090 184.260 109.410 184.520 ;
        RECT 109.640 184.505 109.780 184.660 ;
        RECT 111.480 184.660 115.760 184.800 ;
        RECT 111.480 184.520 111.620 184.660 ;
        RECT 109.565 184.275 109.855 184.505 ;
        RECT 111.390 184.260 111.710 184.520 ;
        RECT 113.230 184.260 113.550 184.520 ;
        RECT 115.620 184.505 115.760 184.660 ;
        RECT 115.545 184.275 115.835 184.505 ;
        RECT 122.430 184.460 122.750 184.520 ;
        RECT 123.825 184.460 124.115 184.505 ;
        RECT 122.430 184.320 124.115 184.460 ;
        RECT 122.430 184.260 122.750 184.320 ;
        RECT 123.825 184.275 124.115 184.320 ;
        RECT 125.205 184.460 125.495 184.505 ;
        RECT 130.250 184.460 130.570 184.520 ;
        RECT 125.205 184.320 130.570 184.460 ;
        RECT 125.205 184.275 125.495 184.320 ;
        RECT 130.250 184.260 130.570 184.320 ;
        RECT 92.545 183.935 92.835 184.165 ;
        RECT 99.445 184.120 99.735 184.165 ;
        RECT 102.205 184.120 102.495 184.165 ;
        RECT 93.080 183.980 102.495 184.120 ;
        RECT 93.080 183.825 93.220 183.980 ;
        RECT 99.445 183.935 99.735 183.980 ;
        RECT 102.205 183.935 102.495 183.980 ;
        RECT 102.665 184.120 102.955 184.165 ;
        RECT 105.410 184.120 105.730 184.180 ;
        RECT 102.665 183.980 105.730 184.120 ;
        RECT 102.665 183.935 102.955 183.980 ;
        RECT 105.410 183.920 105.730 183.980 ;
        RECT 110.010 183.920 110.330 184.180 ;
        RECT 114.165 184.120 114.455 184.165 ;
        RECT 110.560 183.980 114.455 184.120 ;
        RECT 93.005 183.595 93.295 183.825 ;
        RECT 97.605 183.780 97.895 183.825 ;
        RECT 99.890 183.780 100.210 183.840 ;
        RECT 100.365 183.780 100.655 183.825 ;
        RECT 97.605 183.640 100.655 183.780 ;
        RECT 97.605 183.595 97.895 183.640 ;
        RECT 99.890 183.580 100.210 183.640 ;
        RECT 100.365 183.595 100.655 183.640 ;
        RECT 104.030 183.780 104.350 183.840 ;
        RECT 110.560 183.780 110.700 183.980 ;
        RECT 114.165 183.935 114.455 183.980 ;
        RECT 104.030 183.640 110.700 183.780 ;
        RECT 110.945 183.780 111.235 183.825 ;
        RECT 115.085 183.780 115.375 183.825 ;
        RECT 115.530 183.780 115.850 183.840 ;
        RECT 110.945 183.640 115.850 183.780 ;
        RECT 104.030 183.580 104.350 183.640 ;
        RECT 110.945 183.595 111.235 183.640 ;
        RECT 115.085 183.595 115.375 183.640 ;
        RECT 115.530 183.580 115.850 183.640 ;
        RECT 93.465 183.440 93.755 183.485 ;
        RECT 96.210 183.440 96.530 183.500 ;
        RECT 98.050 183.440 98.370 183.500 ;
        RECT 89.860 183.300 98.370 183.440 ;
        RECT 87.010 183.240 87.330 183.300 ;
        RECT 87.485 183.255 87.775 183.300 ;
        RECT 93.465 183.255 93.755 183.300 ;
        RECT 96.210 183.240 96.530 183.300 ;
        RECT 98.050 183.240 98.370 183.300 ;
        RECT 101.745 183.440 102.035 183.485 ;
        RECT 103.110 183.440 103.430 183.500 ;
        RECT 101.745 183.300 103.430 183.440 ;
        RECT 101.745 183.255 102.035 183.300 ;
        RECT 103.110 183.240 103.430 183.300 ;
        RECT 104.965 183.440 105.255 183.485 ;
        RECT 105.410 183.440 105.730 183.500 ;
        RECT 104.965 183.300 105.730 183.440 ;
        RECT 104.965 183.255 105.255 183.300 ;
        RECT 105.410 183.240 105.730 183.300 ;
        RECT 109.090 183.440 109.410 183.500 ;
        RECT 110.485 183.440 110.775 183.485 ;
        RECT 109.090 183.300 110.775 183.440 ;
        RECT 109.090 183.240 109.410 183.300 ;
        RECT 110.485 183.255 110.775 183.300 ;
        RECT 113.230 183.440 113.550 183.500 ;
        RECT 114.625 183.440 114.915 183.485 ;
        RECT 113.230 183.300 114.915 183.440 ;
        RECT 113.230 183.240 113.550 183.300 ;
        RECT 114.625 183.255 114.915 183.300 ;
        RECT 14.260 182.620 126.960 183.100 ;
        RECT 41.010 182.420 41.330 182.480 ;
        RECT 41.945 182.420 42.235 182.465 ;
        RECT 41.010 182.280 42.235 182.420 ;
        RECT 41.010 182.220 41.330 182.280 ;
        RECT 41.945 182.235 42.235 182.280 ;
        RECT 42.390 182.420 42.710 182.480 ;
        RECT 47.005 182.420 47.295 182.465 ;
        RECT 42.390 182.280 47.295 182.420 ;
        RECT 42.390 182.220 42.710 182.280 ;
        RECT 47.005 182.235 47.295 182.280 ;
        RECT 47.450 182.420 47.770 182.480 ;
        RECT 48.830 182.420 49.150 182.480 ;
        RECT 63.090 182.420 63.410 182.480 ;
        RECT 47.450 182.280 49.150 182.420 ;
        RECT 47.450 182.220 47.770 182.280 ;
        RECT 48.830 182.220 49.150 182.280 ;
        RECT 53.980 182.280 63.410 182.420 ;
        RECT 21.705 182.080 21.995 182.125 ;
        RECT 39.170 182.080 39.490 182.140 ;
        RECT 21.705 181.940 35.720 182.080 ;
        RECT 21.705 181.895 21.995 181.940 ;
        RECT 31.825 181.740 32.115 181.785 ;
        RECT 33.190 181.740 33.510 181.800 ;
        RECT 35.580 181.785 35.720 181.940 ;
        RECT 37.880 181.940 39.490 182.080 ;
        RECT 29.135 181.600 31.120 181.740 ;
        RECT 11.110 181.400 11.430 181.460 ;
        RECT 16.185 181.400 16.475 181.445 ;
        RECT 11.110 181.260 16.475 181.400 ;
        RECT 11.110 181.200 11.430 181.260 ;
        RECT 16.185 181.215 16.475 181.260 ;
        RECT 17.565 181.215 17.855 181.445 ;
        RECT 18.010 181.400 18.330 181.460 ;
        RECT 18.485 181.400 18.775 181.445 ;
        RECT 18.010 181.260 18.775 181.400 ;
        RECT 17.640 181.060 17.780 181.215 ;
        RECT 18.010 181.200 18.330 181.260 ;
        RECT 18.485 181.215 18.775 181.260 ;
        RECT 19.865 181.215 20.155 181.445 ;
        RECT 19.940 181.060 20.080 181.215 ;
        RECT 20.770 181.200 21.090 181.460 ;
        RECT 22.165 181.400 22.455 181.445 ;
        RECT 22.610 181.400 22.930 181.460 ;
        RECT 22.165 181.260 22.930 181.400 ;
        RECT 22.165 181.215 22.455 181.260 ;
        RECT 22.610 181.200 22.930 181.260 ;
        RECT 23.085 181.400 23.375 181.445 ;
        RECT 23.530 181.400 23.850 181.460 ;
        RECT 23.085 181.260 23.850 181.400 ;
        RECT 23.085 181.215 23.375 181.260 ;
        RECT 23.530 181.200 23.850 181.260 ;
        RECT 24.450 181.200 24.770 181.460 ;
        RECT 27.210 181.445 27.530 181.460 ;
        RECT 29.135 181.445 29.275 181.600 ;
        RECT 27.200 181.400 27.530 181.445 ;
        RECT 27.015 181.260 27.530 181.400 ;
        RECT 27.200 181.215 27.530 181.260 ;
        RECT 29.060 181.215 29.350 181.445 ;
        RECT 29.525 181.400 29.815 181.445 ;
        RECT 30.430 181.400 30.750 181.460 ;
        RECT 29.525 181.260 30.750 181.400 ;
        RECT 29.525 181.215 29.815 181.260 ;
        RECT 27.210 181.200 27.530 181.215 ;
        RECT 30.430 181.200 30.750 181.260 ;
        RECT 23.990 181.060 24.310 181.120 ;
        RECT 25.830 181.060 26.150 181.120 ;
        RECT 17.640 180.920 18.240 181.060 ;
        RECT 19.940 180.920 24.310 181.060 ;
        RECT 16.170 180.720 16.490 180.780 ;
        RECT 17.105 180.720 17.395 180.765 ;
        RECT 16.170 180.580 17.395 180.720 ;
        RECT 18.100 180.720 18.240 180.920 ;
        RECT 23.990 180.860 24.310 180.920 ;
        RECT 25.000 180.920 26.150 181.060 ;
        RECT 25.000 180.720 25.140 180.920 ;
        RECT 25.830 180.860 26.150 180.920 ;
        RECT 27.670 180.860 27.990 181.120 ;
        RECT 28.145 181.060 28.435 181.105 ;
        RECT 29.985 181.060 30.275 181.105 ;
        RECT 28.145 180.920 30.275 181.060 ;
        RECT 28.145 180.875 28.435 180.920 ;
        RECT 29.985 180.875 30.275 180.920 ;
        RECT 18.100 180.580 25.140 180.720 ;
        RECT 16.170 180.520 16.490 180.580 ;
        RECT 17.105 180.535 17.395 180.580 ;
        RECT 25.370 180.520 25.690 180.780 ;
        RECT 26.305 180.720 26.595 180.765 ;
        RECT 26.750 180.720 27.070 180.780 ;
        RECT 26.305 180.580 27.070 180.720 ;
        RECT 30.980 180.720 31.120 181.600 ;
        RECT 31.825 181.600 33.510 181.740 ;
        RECT 31.825 181.555 32.115 181.600 ;
        RECT 33.190 181.540 33.510 181.600 ;
        RECT 35.505 181.555 35.795 181.785 ;
        RECT 37.880 181.740 38.020 181.940 ;
        RECT 39.170 181.880 39.490 181.940 ;
        RECT 39.630 181.880 39.950 182.140 ;
        RECT 41.470 182.080 41.790 182.140 ;
        RECT 44.230 182.080 44.550 182.140 ;
        RECT 41.470 181.940 44.550 182.080 ;
        RECT 41.470 181.880 41.790 181.940 ;
        RECT 44.230 181.880 44.550 181.940 ;
        RECT 45.150 181.880 45.470 182.140 ;
        RECT 47.910 181.880 48.230 182.140 ;
        RECT 36.040 181.600 38.020 181.740 ;
        RECT 38.265 181.740 38.555 181.785 ;
        RECT 38.725 181.740 39.015 181.785 ;
        RECT 38.265 181.600 39.015 181.740 ;
        RECT 39.720 181.740 39.860 181.880 ;
        RECT 45.245 181.740 45.385 181.880 ;
        RECT 49.290 181.740 49.610 181.800 ;
        RECT 53.980 181.785 54.120 182.280 ;
        RECT 63.090 182.220 63.410 182.280 ;
        RECT 65.390 182.420 65.710 182.480 ;
        RECT 68.625 182.420 68.915 182.465 ;
        RECT 65.390 182.280 68.915 182.420 ;
        RECT 65.390 182.220 65.710 182.280 ;
        RECT 68.625 182.235 68.915 182.280 ;
        RECT 72.290 182.220 72.610 182.480 ;
        RECT 72.750 182.420 73.070 182.480 ;
        RECT 72.750 182.280 83.100 182.420 ;
        RECT 72.750 182.220 73.070 182.280 ;
        RECT 55.730 182.080 56.050 182.140 ;
        RECT 82.410 182.080 82.730 182.140 ;
        RECT 55.730 181.940 61.020 182.080 ;
        RECT 55.730 181.880 56.050 181.940 ;
        RECT 39.720 181.600 41.700 181.740 ;
        RECT 45.245 181.600 46.300 181.740 ;
        RECT 31.350 181.400 31.670 181.460 ;
        RECT 32.515 181.400 32.805 181.445 ;
        RECT 31.350 181.260 32.805 181.400 ;
        RECT 31.350 181.200 31.670 181.260 ;
        RECT 32.515 181.215 32.805 181.260 ;
        RECT 33.650 181.400 33.970 181.460 ;
        RECT 34.125 181.400 34.415 181.445 ;
        RECT 33.650 181.260 34.415 181.400 ;
        RECT 33.650 181.200 33.970 181.260 ;
        RECT 34.125 181.215 34.415 181.260 ;
        RECT 34.585 181.400 34.875 181.445 ;
        RECT 36.040 181.400 36.180 181.600 ;
        RECT 38.265 181.555 38.555 181.600 ;
        RECT 38.725 181.555 39.015 181.600 ;
        RECT 34.585 181.260 36.180 181.400 ;
        RECT 36.425 181.400 36.715 181.445 ;
        RECT 39.170 181.400 39.490 181.460 ;
        RECT 41.560 181.445 41.700 181.600 ;
        RECT 39.645 181.400 39.935 181.445 ;
        RECT 36.425 181.260 38.940 181.400 ;
        RECT 34.585 181.215 34.875 181.260 ;
        RECT 36.425 181.215 36.715 181.260 ;
        RECT 34.200 181.060 34.340 181.215 ;
        RECT 37.330 181.060 37.650 181.120 ;
        RECT 34.200 180.920 37.650 181.060 ;
        RECT 37.330 180.860 37.650 180.920 ;
        RECT 38.800 180.780 38.940 181.260 ;
        RECT 39.170 181.260 39.935 181.400 ;
        RECT 39.170 181.200 39.490 181.260 ;
        RECT 39.645 181.215 39.935 181.260 ;
        RECT 41.485 181.215 41.775 181.445 ;
        RECT 42.865 181.215 43.155 181.445 ;
        RECT 40.550 181.105 40.870 181.120 ;
        RECT 40.550 180.875 40.945 181.105 ;
        RECT 42.390 181.060 42.710 181.120 ;
        RECT 42.940 181.060 43.080 181.215 ;
        RECT 43.770 181.200 44.090 181.460 ;
        RECT 44.705 181.215 44.995 181.445 ;
        RECT 45.165 181.400 45.455 181.445 ;
        RECT 45.610 181.400 45.930 181.460 ;
        RECT 46.160 181.445 46.300 181.600 ;
        RECT 49.290 181.600 53.660 181.740 ;
        RECT 49.290 181.540 49.610 181.600 ;
        RECT 45.165 181.260 45.930 181.400 ;
        RECT 45.165 181.215 45.455 181.260 ;
        RECT 42.390 180.920 43.080 181.060 ;
        RECT 43.325 181.060 43.615 181.105 ;
        RECT 44.230 181.060 44.550 181.120 ;
        RECT 43.325 180.920 44.550 181.060 ;
        RECT 44.780 181.060 44.920 181.215 ;
        RECT 45.610 181.200 45.930 181.260 ;
        RECT 46.085 181.215 46.375 181.445 ;
        RECT 46.530 181.200 46.850 181.460 ;
        RECT 47.450 181.200 47.770 181.460 ;
        RECT 48.845 181.215 49.135 181.445 ;
        RECT 47.910 181.060 48.230 181.120 ;
        RECT 44.780 180.920 48.230 181.060 ;
        RECT 40.550 180.860 40.870 180.875 ;
        RECT 42.390 180.860 42.710 180.920 ;
        RECT 43.325 180.875 43.615 180.920 ;
        RECT 44.230 180.860 44.550 180.920 ;
        RECT 47.910 180.860 48.230 180.920 ;
        RECT 36.425 180.720 36.715 180.765 ;
        RECT 30.980 180.580 36.715 180.720 ;
        RECT 26.305 180.535 26.595 180.580 ;
        RECT 26.750 180.520 27.070 180.580 ;
        RECT 36.425 180.535 36.715 180.580 ;
        RECT 38.710 180.720 39.030 180.780 ;
        RECT 40.105 180.720 40.395 180.765 ;
        RECT 45.625 180.720 45.915 180.765 ;
        RECT 38.710 180.580 45.915 180.720 ;
        RECT 38.710 180.520 39.030 180.580 ;
        RECT 40.105 180.535 40.395 180.580 ;
        RECT 45.625 180.535 45.915 180.580 ;
        RECT 46.070 180.720 46.390 180.780 ;
        RECT 48.920 180.720 49.060 181.215 ;
        RECT 49.750 181.200 50.070 181.460 ;
        RECT 50.760 181.445 50.900 181.600 ;
        RECT 50.685 181.215 50.975 181.445 ;
        RECT 52.970 181.200 53.290 181.460 ;
        RECT 50.225 181.060 50.515 181.105 ;
        RECT 50.225 180.920 53.200 181.060 ;
        RECT 50.225 180.875 50.515 180.920 ;
        RECT 53.060 180.780 53.200 180.920 ;
        RECT 46.070 180.580 49.060 180.720 ;
        RECT 46.070 180.520 46.390 180.580 ;
        RECT 52.050 180.520 52.370 180.780 ;
        RECT 52.970 180.520 53.290 180.780 ;
        RECT 53.520 180.720 53.660 181.600 ;
        RECT 53.905 181.555 54.195 181.785 ;
        RECT 57.570 181.740 57.890 181.800 ;
        RECT 57.200 181.600 57.890 181.740 ;
        RECT 54.350 181.200 54.670 181.460 ;
        RECT 54.825 181.215 55.115 181.445 ;
        RECT 53.890 181.060 54.210 181.120 ;
        RECT 54.900 181.060 55.040 181.215 ;
        RECT 55.730 181.200 56.050 181.460 ;
        RECT 57.200 181.445 57.340 181.600 ;
        RECT 57.570 181.540 57.890 181.600 ;
        RECT 59.410 181.740 59.730 181.800 ;
        RECT 59.410 181.600 60.100 181.740 ;
        RECT 59.410 181.540 59.730 181.600 ;
        RECT 59.960 181.445 60.100 181.600 ;
        RECT 57.125 181.215 57.415 181.445 ;
        RECT 58.505 181.215 58.795 181.445 ;
        RECT 59.885 181.215 60.175 181.445 ;
        RECT 53.890 180.920 55.040 181.060 ;
        RECT 53.890 180.860 54.210 180.920 ;
        RECT 56.205 180.720 56.495 180.765 ;
        RECT 53.520 180.580 56.495 180.720 ;
        RECT 58.580 180.720 58.720 181.215 ;
        RECT 60.330 181.200 60.650 181.460 ;
        RECT 60.880 181.445 61.020 181.940 ;
        RECT 72.840 181.940 82.730 182.080 ;
        RECT 82.960 182.080 83.100 182.280 ;
        RECT 84.250 182.220 84.570 182.480 ;
        RECT 89.310 182.420 89.630 182.480 ;
        RECT 84.800 182.280 89.630 182.420 ;
        RECT 84.800 182.080 84.940 182.280 ;
        RECT 89.310 182.220 89.630 182.280 ;
        RECT 93.450 182.420 93.770 182.480 ;
        RECT 104.030 182.420 104.350 182.480 ;
        RECT 104.950 182.420 105.270 182.480 ;
        RECT 107.710 182.420 108.030 182.480 ;
        RECT 93.450 182.280 108.030 182.420 ;
        RECT 93.450 182.220 93.770 182.280 ;
        RECT 104.030 182.220 104.350 182.280 ;
        RECT 104.950 182.220 105.270 182.280 ;
        RECT 107.710 182.220 108.030 182.280 ;
        RECT 82.960 181.940 84.940 182.080 ;
        RECT 71.370 181.540 71.690 181.800 ;
        RECT 60.805 181.215 61.095 181.445 ;
        RECT 65.850 181.400 66.170 181.460 ;
        RECT 68.165 181.400 68.455 181.445 ;
        RECT 65.850 181.260 68.455 181.400 ;
        RECT 65.850 181.200 66.170 181.260 ;
        RECT 68.165 181.215 68.455 181.260 ;
        RECT 69.085 181.400 69.375 181.445 ;
        RECT 69.530 181.400 69.850 181.460 ;
        RECT 72.840 181.445 72.980 181.940 ;
        RECT 82.410 181.880 82.730 181.940 ;
        RECT 85.170 181.880 85.490 182.140 ;
        RECT 87.945 182.080 88.235 182.125 ;
        RECT 91.150 182.080 91.470 182.140 ;
        RECT 87.945 181.940 91.470 182.080 ;
        RECT 87.945 181.895 88.235 181.940 ;
        RECT 91.150 181.880 91.470 181.940 ;
        RECT 99.445 182.080 99.735 182.125 ;
        RECT 101.730 182.080 102.050 182.140 ;
        RECT 99.445 181.940 102.050 182.080 ;
        RECT 99.445 181.895 99.735 181.940 ;
        RECT 101.730 181.880 102.050 181.940 ;
        RECT 102.205 182.080 102.495 182.125 ;
        RECT 102.650 182.080 102.970 182.140 ;
        RECT 102.205 181.940 102.970 182.080 ;
        RECT 102.205 181.895 102.495 181.940 ;
        RECT 76.430 181.740 76.750 181.800 ;
        RECT 73.760 181.600 76.750 181.740 ;
        RECT 73.760 181.445 73.900 181.600 ;
        RECT 76.430 181.540 76.750 181.600 ;
        RECT 83.330 181.540 83.650 181.800 ;
        RECT 85.260 181.740 85.400 181.880 ;
        RECT 87.470 181.740 87.790 181.800 ;
        RECT 102.280 181.740 102.420 181.895 ;
        RECT 102.650 181.880 102.970 181.940 ;
        RECT 85.260 181.600 86.320 181.740 ;
        RECT 69.085 181.260 69.850 181.400 ;
        RECT 69.085 181.215 69.375 181.260 ;
        RECT 69.530 181.200 69.850 181.260 ;
        RECT 72.765 181.215 73.055 181.445 ;
        RECT 73.685 181.215 73.975 181.445 ;
        RECT 74.605 181.400 74.895 181.445 ;
        RECT 75.050 181.400 75.370 181.460 ;
        RECT 82.885 181.400 83.175 181.445 ;
        RECT 84.250 181.400 84.570 181.460 ;
        RECT 86.180 181.445 86.320 181.600 ;
        RECT 86.640 181.600 102.420 181.740 ;
        RECT 105.410 181.740 105.730 181.800 ;
        RECT 111.865 181.740 112.155 181.785 ;
        RECT 105.410 181.600 112.155 181.740 ;
        RECT 86.640 181.445 86.780 181.600 ;
        RECT 87.470 181.540 87.790 181.600 ;
        RECT 105.410 181.540 105.730 181.600 ;
        RECT 111.865 181.555 112.155 181.600 ;
        RECT 74.605 181.260 84.570 181.400 ;
        RECT 74.605 181.215 74.895 181.260 ;
        RECT 75.050 181.200 75.370 181.260 ;
        RECT 82.885 181.215 83.175 181.260 ;
        RECT 84.250 181.200 84.570 181.260 ;
        RECT 84.725 181.400 85.015 181.445 ;
        RECT 85.185 181.400 85.475 181.445 ;
        RECT 84.725 181.260 85.475 181.400 ;
        RECT 84.725 181.215 85.015 181.260 ;
        RECT 85.185 181.215 85.475 181.260 ;
        RECT 86.105 181.215 86.395 181.445 ;
        RECT 86.565 181.215 86.855 181.445 ;
        RECT 98.970 181.200 99.290 181.460 ;
        RECT 99.890 181.200 100.210 181.460 ;
        RECT 102.665 181.400 102.955 181.445 ;
        RECT 104.030 181.400 104.350 181.460 ;
        RECT 107.250 181.400 107.570 181.460 ;
        RECT 102.665 181.260 104.350 181.400 ;
        RECT 102.665 181.215 102.955 181.260 ;
        RECT 104.030 181.200 104.350 181.260 ;
        RECT 104.580 181.260 107.570 181.400 ;
        RECT 58.950 181.105 59.270 181.120 ;
        RECT 58.950 180.875 59.485 181.105 ;
        RECT 70.910 181.060 71.230 181.120 ;
        RECT 79.190 181.060 79.510 181.120 ;
        RECT 83.790 181.060 84.110 181.120 ;
        RECT 87.025 181.060 87.315 181.105 ;
        RECT 87.930 181.060 88.250 181.120 ;
        RECT 97.130 181.060 97.450 181.120 ;
        RECT 104.580 181.060 104.720 181.260 ;
        RECT 107.250 181.200 107.570 181.260 ;
        RECT 107.710 181.200 108.030 181.460 ;
        RECT 108.170 181.400 108.490 181.460 ;
        RECT 109.105 181.400 109.395 181.445 ;
        RECT 108.170 181.260 109.395 181.400 ;
        RECT 108.170 181.200 108.490 181.260 ;
        RECT 109.105 181.215 109.395 181.260 ;
        RECT 109.875 181.400 110.165 181.445 ;
        RECT 112.770 181.400 113.090 181.460 ;
        RECT 109.875 181.260 113.090 181.400 ;
        RECT 109.875 181.215 110.165 181.260 ;
        RECT 70.910 180.920 73.900 181.060 ;
        RECT 58.950 180.860 59.270 180.875 ;
        RECT 70.910 180.860 71.230 180.920 ;
        RECT 59.870 180.720 60.190 180.780 ;
        RECT 58.580 180.580 60.190 180.720 ;
        RECT 56.205 180.535 56.495 180.580 ;
        RECT 59.870 180.520 60.190 180.580 ;
        RECT 61.710 180.520 62.030 180.780 ;
        RECT 64.010 180.720 64.330 180.780 ;
        RECT 69.530 180.720 69.850 180.780 ;
        RECT 73.760 180.765 73.900 180.920 ;
        RECT 79.190 180.920 84.250 181.060 ;
        RECT 79.190 180.860 79.510 180.920 ;
        RECT 83.790 180.860 84.250 180.920 ;
        RECT 87.025 180.920 88.250 181.060 ;
        RECT 87.025 180.875 87.315 180.920 ;
        RECT 87.930 180.860 88.250 180.920 ;
        RECT 93.080 180.920 104.720 181.060 ;
        RECT 104.950 181.060 105.270 181.120 ;
        RECT 109.180 181.060 109.320 181.215 ;
        RECT 112.770 181.200 113.090 181.260 ;
        RECT 111.850 181.060 112.170 181.120 ;
        RECT 104.950 180.920 109.320 181.060 ;
        RECT 110.560 180.920 112.170 181.060 ;
        RECT 71.385 180.720 71.675 180.765 ;
        RECT 64.010 180.580 71.675 180.720 ;
        RECT 64.010 180.520 64.330 180.580 ;
        RECT 69.530 180.520 69.850 180.580 ;
        RECT 71.385 180.535 71.675 180.580 ;
        RECT 73.685 180.535 73.975 180.765 ;
        RECT 82.870 180.520 83.190 180.780 ;
        RECT 84.110 180.720 84.250 180.860 ;
        RECT 93.080 180.720 93.220 180.920 ;
        RECT 97.130 180.860 97.450 180.920 ;
        RECT 104.950 180.860 105.270 180.920 ;
        RECT 84.110 180.580 93.220 180.720 ;
        RECT 93.450 180.720 93.770 180.780 ;
        RECT 105.410 180.720 105.730 180.780 ;
        RECT 93.450 180.580 105.730 180.720 ;
        RECT 93.450 180.520 93.770 180.580 ;
        RECT 105.410 180.520 105.730 180.580 ;
        RECT 108.185 180.720 108.475 180.765 ;
        RECT 110.560 180.720 110.700 180.920 ;
        RECT 111.850 180.860 112.170 180.920 ;
        RECT 108.185 180.580 110.700 180.720 ;
        RECT 110.945 180.720 111.235 180.765 ;
        RECT 111.390 180.720 111.710 180.780 ;
        RECT 112.785 180.720 113.075 180.765 ;
        RECT 110.945 180.580 113.075 180.720 ;
        RECT 108.185 180.535 108.475 180.580 ;
        RECT 110.945 180.535 111.235 180.580 ;
        RECT 111.390 180.520 111.710 180.580 ;
        RECT 112.785 180.535 113.075 180.580 ;
        RECT 113.230 180.520 113.550 180.780 ;
        RECT 115.085 180.720 115.375 180.765 ;
        RECT 115.990 180.720 116.310 180.780 ;
        RECT 115.085 180.580 116.310 180.720 ;
        RECT 115.085 180.535 115.375 180.580 ;
        RECT 115.990 180.520 116.310 180.580 ;
        RECT 14.260 179.900 126.960 180.380 ;
        RECT 17.565 179.700 17.855 179.745 ;
        RECT 18.010 179.700 18.330 179.760 ;
        RECT 17.565 179.560 18.330 179.700 ;
        RECT 17.565 179.515 17.855 179.560 ;
        RECT 18.010 179.500 18.330 179.560 ;
        RECT 25.370 179.700 25.690 179.760 ;
        RECT 30.890 179.700 31.210 179.760 ;
        RECT 35.950 179.700 36.270 179.760 ;
        RECT 25.370 179.560 31.210 179.700 ;
        RECT 25.370 179.500 25.690 179.560 ;
        RECT 30.890 179.500 31.210 179.560 ;
        RECT 31.900 179.560 36.270 179.700 ;
        RECT 21.230 179.360 21.550 179.420 ;
        RECT 22.165 179.360 22.455 179.405 ;
        RECT 21.230 179.220 22.455 179.360 ;
        RECT 21.230 179.160 21.550 179.220 ;
        RECT 22.165 179.175 22.455 179.220 ;
        RECT 17.105 178.835 17.395 179.065 ;
        RECT 17.180 178.680 17.320 178.835 ;
        RECT 18.470 178.820 18.790 179.080 ;
        RECT 19.850 178.820 20.170 179.080 ;
        RECT 20.785 179.020 21.075 179.065 ;
        RECT 21.690 179.020 22.010 179.080 ;
        RECT 20.785 178.880 22.010 179.020 ;
        RECT 20.785 178.835 21.075 178.880 ;
        RECT 21.690 178.820 22.010 178.880 ;
        RECT 22.610 179.020 22.930 179.080 ;
        RECT 31.365 179.020 31.655 179.065 ;
        RECT 31.900 179.020 32.040 179.560 ;
        RECT 35.950 179.500 36.270 179.560 ;
        RECT 37.330 179.700 37.650 179.760 ;
        RECT 40.565 179.700 40.855 179.745 ;
        RECT 37.330 179.560 40.855 179.700 ;
        RECT 37.330 179.500 37.650 179.560 ;
        RECT 40.565 179.515 40.855 179.560 ;
        RECT 42.390 179.700 42.710 179.760 ;
        RECT 45.610 179.700 45.930 179.760 ;
        RECT 42.390 179.560 45.930 179.700 ;
        RECT 42.390 179.500 42.710 179.560 ;
        RECT 45.610 179.500 45.930 179.560 ;
        RECT 47.910 179.700 48.230 179.760 ;
        RECT 47.910 179.560 49.750 179.700 ;
        RECT 47.910 179.500 48.230 179.560 ;
        RECT 32.730 179.160 33.050 179.420 ;
        RECT 33.190 179.360 33.510 179.420 ;
        RECT 49.610 179.360 49.750 179.560 ;
        RECT 58.950 179.500 59.270 179.760 ;
        RECT 64.010 179.500 64.330 179.760 ;
        RECT 66.310 179.500 66.630 179.760 ;
        RECT 66.770 179.500 67.090 179.760 ;
        RECT 68.150 179.700 68.470 179.760 ;
        RECT 68.625 179.700 68.915 179.745 ;
        RECT 68.150 179.560 68.915 179.700 ;
        RECT 68.150 179.500 68.470 179.560 ;
        RECT 68.625 179.515 68.915 179.560 ;
        RECT 69.085 179.700 69.375 179.745 ;
        RECT 70.450 179.700 70.770 179.760 ;
        RECT 71.830 179.700 72.150 179.760 ;
        RECT 69.085 179.560 72.150 179.700 ;
        RECT 69.085 179.515 69.375 179.560 ;
        RECT 70.450 179.500 70.770 179.560 ;
        RECT 71.830 179.500 72.150 179.560 ;
        RECT 72.750 179.700 73.070 179.760 ;
        RECT 75.050 179.700 75.370 179.760 ;
        RECT 72.750 179.560 75.370 179.700 ;
        RECT 72.750 179.500 73.070 179.560 ;
        RECT 75.050 179.500 75.370 179.560 ;
        RECT 75.510 179.500 75.830 179.760 ;
        RECT 76.430 179.700 76.750 179.760 ;
        RECT 86.550 179.700 86.870 179.760 ;
        RECT 76.430 179.560 86.870 179.700 ;
        RECT 76.430 179.500 76.750 179.560 ;
        RECT 86.550 179.500 86.870 179.560 ;
        RECT 88.850 179.700 89.170 179.760 ;
        RECT 94.385 179.700 94.675 179.745 ;
        RECT 88.850 179.560 94.675 179.700 ;
        RECT 88.850 179.500 89.170 179.560 ;
        RECT 94.385 179.515 94.675 179.560 ;
        RECT 99.905 179.700 100.195 179.745 ;
        RECT 99.905 179.560 101.960 179.700 ;
        RECT 99.905 179.515 100.195 179.560 ;
        RECT 65.850 179.360 66.170 179.420 ;
        RECT 33.190 179.220 44.920 179.360 ;
        RECT 49.610 179.220 66.170 179.360 ;
        RECT 33.190 179.160 33.510 179.220 ;
        RECT 34.110 179.020 34.430 179.080 ;
        RECT 22.610 178.880 30.660 179.020 ;
        RECT 22.610 178.820 22.930 178.880 ;
        RECT 20.310 178.680 20.630 178.740 ;
        RECT 17.180 178.540 20.630 178.680 ;
        RECT 30.520 178.680 30.660 178.880 ;
        RECT 31.365 178.880 32.040 179.020 ;
        RECT 33.915 178.880 34.430 179.020 ;
        RECT 31.365 178.835 31.655 178.880 ;
        RECT 34.110 178.820 34.430 178.880 ;
        RECT 34.585 178.835 34.875 179.065 ;
        RECT 34.660 178.680 34.800 178.835 ;
        RECT 35.030 178.820 35.350 179.080 ;
        RECT 35.965 179.020 36.255 179.065 ;
        RECT 36.410 179.020 36.730 179.080 ;
        RECT 35.965 178.880 36.730 179.020 ;
        RECT 35.965 178.835 36.255 178.880 ;
        RECT 36.410 178.820 36.730 178.880 ;
        RECT 36.870 178.820 37.190 179.080 ;
        RECT 37.330 178.820 37.650 179.080 ;
        RECT 38.265 178.835 38.555 179.065 ;
        RECT 38.725 178.835 39.015 179.065 ;
        RECT 41.010 179.020 41.330 179.080 ;
        RECT 41.485 179.020 41.775 179.065 ;
        RECT 41.010 178.880 41.775 179.020 ;
        RECT 30.520 178.540 34.800 178.680 ;
        RECT 20.310 178.480 20.630 178.540 ;
        RECT 38.345 178.400 38.485 178.835 ;
        RECT 27.210 178.340 27.530 178.400 ;
        RECT 27.210 178.200 35.950 178.340 ;
        RECT 27.210 178.140 27.530 178.200 ;
        RECT 12.950 178.000 13.270 178.060 ;
        RECT 16.185 178.000 16.475 178.045 ;
        RECT 12.950 177.860 16.475 178.000 ;
        RECT 12.950 177.800 13.270 177.860 ;
        RECT 16.185 177.815 16.475 177.860 ;
        RECT 28.590 177.800 28.910 178.060 ;
        RECT 32.285 178.000 32.575 178.045 ;
        RECT 33.650 178.000 33.970 178.060 ;
        RECT 32.285 177.860 33.970 178.000 ;
        RECT 35.810 178.000 35.950 178.200 ;
        RECT 38.250 178.140 38.570 178.400 ;
        RECT 38.800 178.000 38.940 178.835 ;
        RECT 41.010 178.820 41.330 178.880 ;
        RECT 41.485 178.835 41.775 178.880 ;
        RECT 41.930 179.020 42.250 179.080 ;
        RECT 42.405 179.020 42.695 179.065 ;
        RECT 41.930 178.880 42.695 179.020 ;
        RECT 41.930 178.820 42.250 178.880 ;
        RECT 42.405 178.835 42.695 178.880 ;
        RECT 42.850 178.820 43.170 179.080 ;
        RECT 44.230 178.820 44.550 179.080 ;
        RECT 44.780 179.020 44.920 179.220 ;
        RECT 65.850 179.160 66.170 179.220 ;
        RECT 67.230 179.360 67.550 179.420 ;
        RECT 92.070 179.360 92.390 179.420 ;
        RECT 100.825 179.360 101.115 179.405 ;
        RECT 101.270 179.360 101.590 179.420 ;
        RECT 67.230 179.220 81.260 179.360 ;
        RECT 67.230 179.160 67.550 179.220 ;
        RECT 81.120 179.080 81.260 179.220 ;
        RECT 85.720 179.220 89.540 179.360 ;
        RECT 46.545 179.020 46.835 179.065 ;
        RECT 44.780 178.880 46.835 179.020 ;
        RECT 46.545 178.835 46.835 178.880 ;
        RECT 46.990 178.820 47.310 179.080 ;
        RECT 48.385 179.040 48.675 179.065 ;
        RECT 48.385 179.020 49.060 179.040 ;
        RECT 49.290 179.020 49.610 179.080 ;
        RECT 48.385 178.900 49.610 179.020 ;
        RECT 48.385 178.835 48.675 178.900 ;
        RECT 48.920 178.880 49.610 178.900 ;
        RECT 49.290 178.820 49.610 178.880 ;
        RECT 49.750 178.820 50.070 179.080 ;
        RECT 50.685 178.835 50.975 179.065 ;
        RECT 51.590 179.020 51.910 179.080 ;
        RECT 53.430 179.065 53.750 179.080 ;
        RECT 52.065 179.020 52.355 179.065 ;
        RECT 51.590 178.880 52.355 179.020 ;
        RECT 44.690 178.680 45.010 178.740 ;
        RECT 47.080 178.680 47.220 178.820 ;
        RECT 44.690 178.540 47.220 178.680 ;
        RECT 47.465 178.680 47.755 178.725 ;
        RECT 48.830 178.680 49.150 178.740 ;
        RECT 50.760 178.680 50.900 178.835 ;
        RECT 51.590 178.820 51.910 178.880 ;
        RECT 52.065 178.835 52.355 178.880 ;
        RECT 53.325 178.835 53.750 179.065 ;
        RECT 53.430 178.820 53.750 178.835 ;
        RECT 53.890 178.820 54.210 179.080 ;
        RECT 54.350 178.820 54.670 179.080 ;
        RECT 55.285 179.020 55.575 179.065 ;
        RECT 56.190 179.020 56.510 179.080 ;
        RECT 55.285 178.880 56.510 179.020 ;
        RECT 55.285 178.835 55.575 178.880 ;
        RECT 56.190 178.820 56.510 178.880 ;
        RECT 56.650 179.020 56.970 179.080 ;
        RECT 57.570 179.020 57.890 179.080 ;
        RECT 56.650 178.880 57.890 179.020 ;
        RECT 56.650 178.820 56.970 178.880 ;
        RECT 57.570 178.820 57.890 178.880 ;
        RECT 58.045 179.020 58.335 179.065 ;
        RECT 59.410 179.020 59.730 179.080 ;
        RECT 58.045 178.880 59.730 179.020 ;
        RECT 58.045 178.835 58.335 178.880 ;
        RECT 59.410 178.820 59.730 178.880 ;
        RECT 64.485 179.020 64.775 179.065 ;
        RECT 70.910 179.020 71.230 179.080 ;
        RECT 64.485 178.880 71.230 179.020 ;
        RECT 64.485 178.835 64.775 178.880 ;
        RECT 70.910 178.820 71.230 178.880 ;
        RECT 71.830 178.820 72.150 179.080 ;
        RECT 72.750 178.820 73.070 179.080 ;
        RECT 75.540 179.020 75.830 179.065 ;
        RECT 77.810 179.020 78.130 179.080 ;
        RECT 73.760 178.880 78.130 179.020 ;
        RECT 47.465 178.540 49.150 178.680 ;
        RECT 44.690 178.480 45.010 178.540 ;
        RECT 47.465 178.495 47.755 178.540 ;
        RECT 48.830 178.480 49.150 178.540 ;
        RECT 49.610 178.540 50.900 178.680 ;
        RECT 63.090 178.680 63.410 178.740 ;
        RECT 69.545 178.680 69.835 178.725 ;
        RECT 72.305 178.680 72.595 178.725 ;
        RECT 63.090 178.540 69.835 178.680 ;
        RECT 40.550 178.340 40.870 178.400 ;
        RECT 43.310 178.340 43.630 178.400 ;
        RECT 40.550 178.200 43.630 178.340 ;
        RECT 40.550 178.140 40.870 178.200 ;
        RECT 43.310 178.140 43.630 178.200 ;
        RECT 45.610 178.140 45.930 178.400 ;
        RECT 46.990 178.340 47.310 178.400 ;
        RECT 49.610 178.340 49.750 178.540 ;
        RECT 63.090 178.480 63.410 178.540 ;
        RECT 69.545 178.495 69.835 178.540 ;
        RECT 69.995 178.540 72.595 178.680 ;
        RECT 46.990 178.200 49.750 178.340 ;
        RECT 46.990 178.140 47.310 178.200 ;
        RECT 51.130 178.140 51.450 178.400 ;
        RECT 52.050 178.340 52.370 178.400 ;
        RECT 56.190 178.340 56.510 178.400 ;
        RECT 52.050 178.200 56.510 178.340 ;
        RECT 52.050 178.140 52.370 178.200 ;
        RECT 56.190 178.140 56.510 178.200 ;
        RECT 68.150 178.340 68.470 178.400 ;
        RECT 69.995 178.340 70.135 178.540 ;
        RECT 72.305 178.495 72.595 178.540 ;
        RECT 73.210 178.480 73.530 178.740 ;
        RECT 73.760 178.340 73.900 178.880 ;
        RECT 75.540 178.835 75.830 178.880 ;
        RECT 77.810 178.820 78.130 178.880 ;
        RECT 78.270 178.820 78.590 179.080 ;
        RECT 79.665 179.020 79.955 179.065 ;
        RECT 78.820 178.880 79.955 179.020 ;
        RECT 74.590 178.680 74.910 178.740 ;
        RECT 78.820 178.680 78.960 178.880 ;
        RECT 79.665 178.835 79.955 178.880 ;
        RECT 80.110 178.820 80.430 179.080 ;
        RECT 81.030 178.820 81.350 179.080 ;
        RECT 85.170 179.020 85.490 179.080 ;
        RECT 85.720 179.065 85.860 179.220 ;
        RECT 85.645 179.020 85.935 179.065 ;
        RECT 85.170 178.880 85.935 179.020 ;
        RECT 85.170 178.820 85.490 178.880 ;
        RECT 85.645 178.835 85.935 178.880 ;
        RECT 86.550 178.820 86.870 179.080 ;
        RECT 87.010 178.820 87.330 179.080 ;
        RECT 89.400 179.065 89.540 179.220 ;
        RECT 90.320 179.220 92.390 179.360 ;
        RECT 90.320 179.065 90.460 179.220 ;
        RECT 92.070 179.160 92.390 179.220 ;
        RECT 99.060 179.220 101.590 179.360 ;
        RECT 89.325 178.835 89.615 179.065 ;
        RECT 90.245 178.835 90.535 179.065 ;
        RECT 90.690 179.020 91.010 179.080 ;
        RECT 99.060 179.065 99.200 179.220 ;
        RECT 100.825 179.175 101.115 179.220 ;
        RECT 101.270 179.160 101.590 179.220 ;
        RECT 101.820 179.080 101.960 179.560 ;
        RECT 104.030 179.500 104.350 179.760 ;
        RECT 107.265 179.700 107.555 179.745 ;
        RECT 108.170 179.700 108.490 179.760 ;
        RECT 107.265 179.560 108.490 179.700 ;
        RECT 107.265 179.515 107.555 179.560 ;
        RECT 108.170 179.500 108.490 179.560 ;
        RECT 111.390 179.500 111.710 179.760 ;
        RECT 110.945 179.360 111.235 179.405 ;
        RECT 113.230 179.360 113.550 179.420 ;
        RECT 105.500 179.220 108.860 179.360 ;
        RECT 98.985 179.020 99.275 179.065 ;
        RECT 90.690 178.880 99.275 179.020 ;
        RECT 74.590 178.540 78.960 178.680 ;
        RECT 74.590 178.480 74.910 178.540 ;
        RECT 79.205 178.495 79.495 178.725 ;
        RECT 84.250 178.680 84.570 178.740 ;
        RECT 86.105 178.680 86.395 178.725 ;
        RECT 87.470 178.680 87.790 178.740 ;
        RECT 90.320 178.680 90.460 178.835 ;
        RECT 90.690 178.820 91.010 178.880 ;
        RECT 98.985 178.835 99.275 178.880 ;
        RECT 100.350 178.820 100.670 179.080 ;
        RECT 101.730 178.820 102.050 179.080 ;
        RECT 102.205 179.020 102.495 179.065 ;
        RECT 102.650 179.020 102.970 179.080 ;
        RECT 102.205 178.880 102.970 179.020 ;
        RECT 102.205 178.835 102.495 178.880 ;
        RECT 102.650 178.820 102.970 178.880 ;
        RECT 103.570 178.820 103.890 179.080 ;
        RECT 104.490 179.020 104.810 179.080 ;
        RECT 105.500 179.065 105.640 179.220 ;
        RECT 105.425 179.020 105.715 179.065 ;
        RECT 104.490 178.880 105.715 179.020 ;
        RECT 104.490 178.820 104.810 178.880 ;
        RECT 105.425 178.835 105.715 178.880 ;
        RECT 106.345 179.020 106.635 179.065 ;
        RECT 107.250 179.020 107.570 179.080 ;
        RECT 108.720 179.065 108.860 179.220 ;
        RECT 110.945 179.220 113.550 179.360 ;
        RECT 110.945 179.175 111.235 179.220 ;
        RECT 113.230 179.160 113.550 179.220 ;
        RECT 108.185 179.020 108.475 179.065 ;
        RECT 106.345 178.880 108.475 179.020 ;
        RECT 106.345 178.835 106.635 178.880 ;
        RECT 107.250 178.820 107.570 178.880 ;
        RECT 108.185 178.835 108.475 178.880 ;
        RECT 108.645 178.835 108.935 179.065 ;
        RECT 114.165 179.020 114.455 179.065 ;
        RECT 109.180 179.010 110.240 179.020 ;
        RECT 110.560 179.010 114.455 179.020 ;
        RECT 109.180 178.880 114.455 179.010 ;
        RECT 84.250 178.540 90.460 178.680 ;
        RECT 68.150 178.200 70.135 178.340 ;
        RECT 70.310 178.200 73.900 178.340 ;
        RECT 76.445 178.340 76.735 178.385 ;
        RECT 79.280 178.340 79.420 178.495 ;
        RECT 84.250 178.480 84.570 178.540 ;
        RECT 86.105 178.495 86.395 178.540 ;
        RECT 87.470 178.480 87.790 178.540 ;
        RECT 93.450 178.480 93.770 178.740 ;
        RECT 93.925 178.495 94.215 178.725 ;
        RECT 95.750 178.680 96.070 178.740 ;
        RECT 104.580 178.680 104.720 178.820 ;
        RECT 95.750 178.540 104.720 178.680 ;
        RECT 105.885 178.680 106.175 178.725 ;
        RECT 106.790 178.680 107.110 178.740 ;
        RECT 109.180 178.680 109.320 178.880 ;
        RECT 110.100 178.870 110.700 178.880 ;
        RECT 114.165 178.835 114.455 178.880 ;
        RECT 115.530 178.820 115.850 179.080 ;
        RECT 115.990 178.820 116.310 179.080 ;
        RECT 105.885 178.540 109.320 178.680 ;
        RECT 76.445 178.200 79.420 178.340 ;
        RECT 85.630 178.340 85.950 178.400 ;
        RECT 87.930 178.340 88.250 178.400 ;
        RECT 94.000 178.340 94.140 178.495 ;
        RECT 95.750 178.480 96.070 178.540 ;
        RECT 105.885 178.495 106.175 178.540 ;
        RECT 106.790 178.480 107.110 178.540 ;
        RECT 110.025 178.495 110.315 178.725 ;
        RECT 85.630 178.200 88.250 178.340 ;
        RECT 68.150 178.140 68.470 178.200 ;
        RECT 35.810 177.860 38.940 178.000 ;
        RECT 32.285 177.815 32.575 177.860 ;
        RECT 33.650 177.800 33.970 177.860 ;
        RECT 39.630 177.800 39.950 178.060 ;
        RECT 43.770 177.800 44.090 178.060 ;
        RECT 45.150 177.800 45.470 178.060 ;
        RECT 48.830 177.800 49.150 178.060 ;
        RECT 49.765 178.000 50.055 178.045 ;
        RECT 50.210 178.000 50.530 178.060 ;
        RECT 49.765 177.860 50.530 178.000 ;
        RECT 49.765 177.815 50.055 177.860 ;
        RECT 50.210 177.800 50.530 177.860 ;
        RECT 50.670 178.000 50.990 178.060 ;
        RECT 52.525 178.000 52.815 178.045 ;
        RECT 50.670 177.860 52.815 178.000 ;
        RECT 50.670 177.800 50.990 177.860 ;
        RECT 52.525 177.815 52.815 177.860 ;
        RECT 54.810 178.000 55.130 178.060 ;
        RECT 56.650 178.000 56.970 178.060 ;
        RECT 54.810 177.860 56.970 178.000 ;
        RECT 54.810 177.800 55.130 177.860 ;
        RECT 56.650 177.800 56.970 177.860 ;
        RECT 57.110 177.800 57.430 178.060 ;
        RECT 64.470 178.000 64.790 178.060 ;
        RECT 70.310 178.000 70.450 178.200 ;
        RECT 76.445 178.155 76.735 178.200 ;
        RECT 85.630 178.140 85.950 178.200 ;
        RECT 87.930 178.140 88.250 178.200 ;
        RECT 89.860 178.200 94.140 178.340 ;
        RECT 89.860 178.060 90.000 178.200 ;
        RECT 100.810 178.140 101.130 178.400 ;
        RECT 105.410 178.340 105.730 178.400 ;
        RECT 110.100 178.340 110.240 178.495 ;
        RECT 105.410 178.200 110.240 178.340 ;
        RECT 113.245 178.340 113.535 178.385 ;
        RECT 114.625 178.340 114.915 178.385 ;
        RECT 113.245 178.200 114.915 178.340 ;
        RECT 105.410 178.140 105.730 178.200 ;
        RECT 113.245 178.155 113.535 178.200 ;
        RECT 114.625 178.155 114.915 178.200 ;
        RECT 64.470 177.860 70.450 178.000 ;
        RECT 64.470 177.800 64.790 177.860 ;
        RECT 73.670 177.800 73.990 178.060 ;
        RECT 77.825 178.000 78.115 178.045 ;
        RECT 79.650 178.000 79.970 178.060 ;
        RECT 77.825 177.860 79.970 178.000 ;
        RECT 77.825 177.815 78.115 177.860 ;
        RECT 79.650 177.800 79.970 177.860 ;
        RECT 84.250 178.000 84.570 178.060 ;
        RECT 84.725 178.000 85.015 178.045 ;
        RECT 84.250 177.860 85.015 178.000 ;
        RECT 84.250 177.800 84.570 177.860 ;
        RECT 84.725 177.815 85.015 177.860 ;
        RECT 89.770 177.800 90.090 178.060 ;
        RECT 96.225 178.000 96.515 178.045 ;
        RECT 97.590 178.000 97.910 178.060 ;
        RECT 96.225 177.860 97.910 178.000 ;
        RECT 96.225 177.815 96.515 177.860 ;
        RECT 97.590 177.800 97.910 177.860 ;
        RECT 98.050 177.800 98.370 178.060 ;
        RECT 102.650 178.000 102.970 178.060 ;
        RECT 116.925 178.000 117.215 178.045 ;
        RECT 102.650 177.860 117.215 178.000 ;
        RECT 102.650 177.800 102.970 177.860 ;
        RECT 116.925 177.815 117.215 177.860 ;
        RECT 14.260 177.180 126.960 177.660 ;
        RECT 16.185 176.980 16.475 177.025 ;
        RECT 18.930 176.980 19.250 177.040 ;
        RECT 23.070 176.980 23.390 177.040 ;
        RECT 16.185 176.840 19.250 176.980 ;
        RECT 16.185 176.795 16.475 176.840 ;
        RECT 18.930 176.780 19.250 176.840 ;
        RECT 22.010 176.840 23.390 176.980 ;
        RECT 15.250 176.640 15.570 176.700 ;
        RECT 17.565 176.640 17.855 176.685 ;
        RECT 20.770 176.640 21.090 176.700 ;
        RECT 15.250 176.500 17.855 176.640 ;
        RECT 15.250 176.440 15.570 176.500 ;
        RECT 17.565 176.455 17.855 176.500 ;
        RECT 19.940 176.500 21.090 176.640 ;
        RECT 17.090 175.760 17.410 176.020 ;
        RECT 18.485 175.960 18.775 176.005 ;
        RECT 19.390 175.960 19.710 176.020 ;
        RECT 19.940 176.005 20.080 176.500 ;
        RECT 20.770 176.440 21.090 176.500 ;
        RECT 22.010 176.300 22.150 176.840 ;
        RECT 23.070 176.780 23.390 176.840 ;
        RECT 23.530 176.980 23.850 177.040 ;
        RECT 39.645 176.980 39.935 177.025 ;
        RECT 40.090 176.980 40.410 177.040 ;
        RECT 23.530 176.840 40.410 176.980 ;
        RECT 23.530 176.780 23.850 176.840 ;
        RECT 39.645 176.795 39.935 176.840 ;
        RECT 40.090 176.780 40.410 176.840 ;
        RECT 42.390 176.980 42.710 177.040 ;
        RECT 43.785 176.980 44.075 177.025 ;
        RECT 42.390 176.840 44.075 176.980 ;
        RECT 42.390 176.780 42.710 176.840 ;
        RECT 43.785 176.795 44.075 176.840 ;
        RECT 45.150 176.980 45.470 177.040 ;
        RECT 49.290 176.980 49.610 177.040 ;
        RECT 45.150 176.840 49.610 176.980 ;
        RECT 45.150 176.780 45.470 176.840 ;
        RECT 49.290 176.780 49.610 176.840 ;
        RECT 52.065 176.980 52.355 177.025 ;
        RECT 56.665 176.980 56.955 177.025 ;
        RECT 63.090 176.980 63.410 177.040 ;
        RECT 52.065 176.840 56.420 176.980 ;
        RECT 52.065 176.795 52.355 176.840 ;
        RECT 43.325 176.640 43.615 176.685 ;
        RECT 44.690 176.640 45.010 176.700 ;
        RECT 48.370 176.640 48.690 176.700 ;
        RECT 55.285 176.640 55.575 176.685 ;
        RECT 56.280 176.640 56.420 176.840 ;
        RECT 56.665 176.840 63.410 176.980 ;
        RECT 56.665 176.795 56.955 176.840 ;
        RECT 63.090 176.780 63.410 176.840 ;
        RECT 71.845 176.980 72.135 177.025 ;
        RECT 73.210 176.980 73.530 177.040 ;
        RECT 71.845 176.840 73.530 176.980 ;
        RECT 71.845 176.795 72.135 176.840 ;
        RECT 73.210 176.780 73.530 176.840 ;
        RECT 81.950 176.780 82.270 177.040 ;
        RECT 82.410 176.980 82.730 177.040 ;
        RECT 95.750 176.980 96.070 177.040 ;
        RECT 82.410 176.840 96.070 176.980 ;
        RECT 82.410 176.780 82.730 176.840 ;
        RECT 95.750 176.780 96.070 176.840 ;
        RECT 96.225 176.980 96.515 177.025 ;
        RECT 97.145 176.980 97.435 177.025 ;
        RECT 96.225 176.840 97.435 176.980 ;
        RECT 96.225 176.795 96.515 176.840 ;
        RECT 97.145 176.795 97.435 176.840 ;
        RECT 99.445 176.980 99.735 177.025 ;
        RECT 100.350 176.980 100.670 177.040 ;
        RECT 99.445 176.840 100.670 176.980 ;
        RECT 99.445 176.795 99.735 176.840 ;
        RECT 100.350 176.780 100.670 176.840 ;
        RECT 101.285 176.980 101.575 177.025 ;
        RECT 101.730 176.980 102.050 177.040 ;
        RECT 101.285 176.840 102.050 176.980 ;
        RECT 101.285 176.795 101.575 176.840 ;
        RECT 101.730 176.780 102.050 176.840 ;
        RECT 107.250 176.980 107.570 177.040 ;
        RECT 111.850 176.980 112.170 177.040 ;
        RECT 107.250 176.840 121.740 176.980 ;
        RECT 107.250 176.780 107.570 176.840 ;
        RECT 111.850 176.780 112.170 176.840 ;
        RECT 61.725 176.640 62.015 176.685 ;
        RECT 62.170 176.640 62.490 176.700 ;
        RECT 43.325 176.500 45.010 176.640 ;
        RECT 43.325 176.455 43.615 176.500 ;
        RECT 44.690 176.440 45.010 176.500 ;
        RECT 46.670 176.500 48.690 176.640 ;
        RECT 20.860 176.160 22.150 176.300 ;
        RECT 25.830 176.300 26.150 176.360 ;
        RECT 41.470 176.300 41.790 176.360 ;
        RECT 25.830 176.160 41.790 176.300 ;
        RECT 20.860 176.005 21.000 176.160 ;
        RECT 25.830 176.100 26.150 176.160 ;
        RECT 41.470 176.100 41.790 176.160 ;
        RECT 41.930 176.100 42.250 176.360 ;
        RECT 46.670 176.300 46.810 176.500 ;
        RECT 48.370 176.440 48.690 176.500 ;
        RECT 51.680 176.500 53.200 176.640 ;
        RECT 44.780 176.160 46.810 176.300 ;
        RECT 18.485 175.820 19.710 175.960 ;
        RECT 18.485 175.775 18.775 175.820 ;
        RECT 19.390 175.760 19.710 175.820 ;
        RECT 19.865 175.775 20.155 176.005 ;
        RECT 20.785 175.775 21.075 176.005 ;
        RECT 22.165 175.775 22.455 176.005 ;
        RECT 24.925 175.960 25.215 176.005 ;
        RECT 28.590 175.960 28.910 176.020 ;
        RECT 24.925 175.820 28.910 175.960 ;
        RECT 24.925 175.775 25.215 175.820 ;
        RECT 9.730 175.620 10.050 175.680 ;
        RECT 22.240 175.620 22.380 175.775 ;
        RECT 28.590 175.760 28.910 175.820 ;
        RECT 31.350 175.960 31.670 176.020 ;
        RECT 32.285 175.960 32.575 176.005 ;
        RECT 31.350 175.820 32.575 175.960 ;
        RECT 31.350 175.760 31.670 175.820 ;
        RECT 32.285 175.775 32.575 175.820 ;
        RECT 33.205 175.960 33.495 176.005 ;
        RECT 35.490 175.960 35.810 176.020 ;
        RECT 33.205 175.820 35.810 175.960 ;
        RECT 33.205 175.775 33.495 175.820 ;
        RECT 35.490 175.760 35.810 175.820 ;
        RECT 38.710 175.960 39.030 176.020 ;
        RECT 42.020 175.960 42.160 176.100 ;
        RECT 38.710 175.820 42.160 175.960 ;
        RECT 38.710 175.760 39.030 175.820 ;
        RECT 42.435 175.775 42.725 176.005 ;
        RECT 43.310 175.960 43.630 176.020 ;
        RECT 44.780 176.005 44.920 176.160 ;
        RECT 46.990 176.100 47.310 176.360 ;
        RECT 51.680 176.300 51.820 176.500 ;
        RECT 51.220 176.160 51.820 176.300 ;
        RECT 53.060 176.300 53.200 176.500 ;
        RECT 55.285 176.500 55.960 176.640 ;
        RECT 56.280 176.500 61.505 176.640 ;
        RECT 55.285 176.455 55.575 176.500 ;
        RECT 55.820 176.300 55.960 176.500 ;
        RECT 61.365 176.300 61.505 176.500 ;
        RECT 61.725 176.500 62.490 176.640 ;
        RECT 61.725 176.455 62.015 176.500 ;
        RECT 62.170 176.440 62.490 176.500 ;
        RECT 67.690 176.640 68.010 176.700 ;
        RECT 75.050 176.640 75.370 176.700 ;
        RECT 98.050 176.640 98.370 176.700 ;
        RECT 103.110 176.640 103.430 176.700 ;
        RECT 67.690 176.500 75.370 176.640 ;
        RECT 67.690 176.440 68.010 176.500 ;
        RECT 75.050 176.440 75.370 176.500 ;
        RECT 84.800 176.500 98.370 176.640 ;
        RECT 64.485 176.300 64.775 176.345 ;
        RECT 68.625 176.300 68.915 176.345 ;
        RECT 53.060 176.160 55.500 176.300 ;
        RECT 55.820 176.160 58.260 176.300 ;
        RECT 61.365 176.160 68.915 176.300 ;
        RECT 43.310 175.820 44.460 175.960 ;
        RECT 9.730 175.480 22.380 175.620 ;
        RECT 41.930 175.620 42.250 175.680 ;
        RECT 42.510 175.620 42.650 175.775 ;
        RECT 43.310 175.760 43.630 175.820 ;
        RECT 41.930 175.480 42.650 175.620 ;
        RECT 44.320 175.620 44.460 175.820 ;
        RECT 44.705 175.775 44.995 176.005 ;
        RECT 46.215 175.970 46.505 176.005 ;
        RECT 46.215 175.960 46.810 175.970 ;
        RECT 47.910 175.960 48.230 176.020 ;
        RECT 46.215 175.830 48.230 175.960 ;
        RECT 46.215 175.820 46.530 175.830 ;
        RECT 46.670 175.820 48.230 175.830 ;
        RECT 46.215 175.775 46.505 175.820 ;
        RECT 47.910 175.760 48.230 175.820 ;
        RECT 48.370 175.760 48.690 176.020 ;
        RECT 48.845 175.960 49.135 176.005 ;
        RECT 48.845 175.820 50.440 175.960 ;
        RECT 48.845 175.775 49.135 175.820 ;
        RECT 45.165 175.620 45.455 175.665 ;
        RECT 44.320 175.480 45.455 175.620 ;
        RECT 9.730 175.420 10.050 175.480 ;
        RECT 41.930 175.420 42.250 175.480 ;
        RECT 45.165 175.435 45.455 175.480 ;
        RECT 45.610 175.620 45.930 175.680 ;
        RECT 50.300 175.620 50.440 175.820 ;
        RECT 50.670 175.760 50.990 176.020 ;
        RECT 51.220 176.005 51.360 176.160 ;
        RECT 51.145 175.775 51.435 176.005 ;
        RECT 52.050 175.760 52.370 176.020 ;
        RECT 52.510 175.760 52.830 176.020 ;
        RECT 53.890 175.960 54.210 176.020 ;
        RECT 53.060 175.820 54.210 175.960 ;
        RECT 53.060 175.620 53.200 175.820 ;
        RECT 53.890 175.760 54.210 175.820 ;
        RECT 54.365 175.960 54.655 176.005 ;
        RECT 54.810 175.960 55.130 176.020 ;
        RECT 54.365 175.820 55.130 175.960 ;
        RECT 55.360 175.960 55.500 176.160 ;
        RECT 58.120 176.005 58.260 176.160 ;
        RECT 64.485 176.115 64.775 176.160 ;
        RECT 68.625 176.115 68.915 176.160 ;
        RECT 69.530 176.100 69.850 176.360 ;
        RECT 70.910 176.300 71.230 176.360 ;
        RECT 70.080 176.160 71.230 176.300 ;
        RECT 58.045 175.960 58.335 176.005 ;
        RECT 59.425 175.960 59.715 176.005 ;
        RECT 55.360 175.820 57.800 175.960 ;
        RECT 54.365 175.775 54.655 175.820 ;
        RECT 54.810 175.760 55.130 175.820 ;
        RECT 45.610 175.480 49.750 175.620 ;
        RECT 50.300 175.480 53.200 175.620 ;
        RECT 45.610 175.420 45.930 175.480 ;
        RECT 48.830 175.280 49.150 175.340 ;
        RECT 13.960 175.140 49.150 175.280 ;
        RECT 49.610 175.280 49.750 175.480 ;
        RECT 53.430 175.420 53.750 175.680 ;
        RECT 56.650 175.420 56.970 175.680 ;
        RECT 57.660 175.665 57.800 175.820 ;
        RECT 58.045 175.820 59.715 175.960 ;
        RECT 58.045 175.775 58.335 175.820 ;
        RECT 59.425 175.775 59.715 175.820 ;
        RECT 59.870 175.760 60.190 176.020 ;
        RECT 60.805 175.960 61.095 176.005 ;
        RECT 61.710 175.960 62.030 176.020 ;
        RECT 60.805 175.820 62.030 175.960 ;
        RECT 60.805 175.775 61.095 175.820 ;
        RECT 61.710 175.760 62.030 175.820 ;
        RECT 65.865 175.960 66.155 176.005 ;
        RECT 68.150 175.960 68.470 176.020 ;
        RECT 70.080 176.005 70.220 176.160 ;
        RECT 70.910 176.100 71.230 176.160 ;
        RECT 78.730 176.300 79.050 176.360 ;
        RECT 79.665 176.300 79.955 176.345 ;
        RECT 78.730 176.160 79.955 176.300 ;
        RECT 78.730 176.100 79.050 176.160 ;
        RECT 79.665 176.115 79.955 176.160 ;
        RECT 81.045 176.300 81.335 176.345 ;
        RECT 82.885 176.300 83.175 176.345 ;
        RECT 81.045 176.160 83.175 176.300 ;
        RECT 81.045 176.115 81.335 176.160 ;
        RECT 82.885 176.115 83.175 176.160 ;
        RECT 65.865 175.820 68.470 175.960 ;
        RECT 65.865 175.775 66.155 175.820 ;
        RECT 68.150 175.760 68.470 175.820 ;
        RECT 70.005 175.775 70.295 176.005 ;
        RECT 78.270 175.960 78.590 176.020 ;
        RECT 71.000 175.820 78.590 175.960 ;
        RECT 57.585 175.620 57.875 175.665 ;
        RECT 59.960 175.620 60.100 175.760 ;
        RECT 57.585 175.480 60.100 175.620 ;
        RECT 65.405 175.620 65.695 175.665 ;
        RECT 70.450 175.620 70.770 175.680 ;
        RECT 65.405 175.480 70.770 175.620 ;
        RECT 57.585 175.435 57.875 175.480 ;
        RECT 65.405 175.435 65.695 175.480 ;
        RECT 70.450 175.420 70.770 175.480 ;
        RECT 66.770 175.280 67.090 175.340 ;
        RECT 49.610 175.140 67.090 175.280 ;
        RECT 13.960 173.580 14.100 175.140 ;
        RECT 48.830 175.080 49.150 175.140 ;
        RECT 66.770 175.080 67.090 175.140 ;
        RECT 67.690 175.080 68.010 175.340 ;
        RECT 68.150 175.280 68.470 175.340 ;
        RECT 69.990 175.280 70.310 175.340 ;
        RECT 71.000 175.280 71.140 175.820 ;
        RECT 78.270 175.760 78.590 175.820 ;
        RECT 79.190 175.760 79.510 176.020 ;
        RECT 80.110 175.960 80.430 176.020 ;
        RECT 84.800 176.005 84.940 176.500 ;
        RECT 98.050 176.440 98.370 176.500 ;
        RECT 98.600 176.500 103.430 176.640 ;
        RECT 89.325 176.300 89.615 176.345 ;
        RECT 93.465 176.300 93.755 176.345 ;
        RECT 98.600 176.300 98.740 176.500 ;
        RECT 103.110 176.440 103.430 176.500 ;
        RECT 108.630 176.640 108.950 176.700 ;
        RECT 112.325 176.640 112.615 176.685 ;
        RECT 108.630 176.500 112.615 176.640 ;
        RECT 108.630 176.440 108.950 176.500 ;
        RECT 112.325 176.455 112.615 176.500 ;
        RECT 104.030 176.300 104.350 176.360 ;
        RECT 109.565 176.300 109.855 176.345 ;
        RECT 89.325 176.160 98.740 176.300 ;
        RECT 102.280 176.160 104.720 176.300 ;
        RECT 89.325 176.115 89.615 176.160 ;
        RECT 93.465 176.115 93.755 176.160 ;
        RECT 83.805 175.960 84.095 176.005 ;
        RECT 80.110 175.820 84.095 175.960 ;
        RECT 80.110 175.760 80.430 175.820 ;
        RECT 83.805 175.775 84.095 175.820 ;
        RECT 84.725 175.775 85.015 176.005 ;
        RECT 85.185 175.775 85.475 176.005 ;
        RECT 86.090 175.960 86.410 176.020 ;
        RECT 86.565 175.960 86.855 176.005 ;
        RECT 86.090 175.820 86.855 175.960 ;
        RECT 80.585 175.620 80.875 175.665 ;
        RECT 81.030 175.620 81.350 175.680 ;
        RECT 80.585 175.480 81.350 175.620 ;
        RECT 80.585 175.435 80.875 175.480 ;
        RECT 81.030 175.420 81.350 175.480 ;
        RECT 82.870 175.620 83.190 175.680 ;
        RECT 85.260 175.620 85.400 175.775 ;
        RECT 86.090 175.760 86.410 175.820 ;
        RECT 86.565 175.775 86.855 175.820 ;
        RECT 87.470 175.760 87.790 176.020 ;
        RECT 88.850 175.960 89.170 176.020 ;
        RECT 90.245 175.960 90.535 176.005 ;
        RECT 88.850 175.820 90.535 175.960 ;
        RECT 88.850 175.760 89.170 175.820 ;
        RECT 90.245 175.775 90.535 175.820 ;
        RECT 90.690 175.960 91.010 176.020 ;
        RECT 97.130 176.005 97.450 176.020 ;
        RECT 94.385 175.960 94.675 176.005 ;
        RECT 90.690 175.820 94.675 175.960 ;
        RECT 90.690 175.760 91.010 175.820 ;
        RECT 94.385 175.775 94.675 175.820 ;
        RECT 96.915 175.960 97.450 176.005 ;
        RECT 96.915 175.820 97.820 175.960 ;
        RECT 96.915 175.775 97.450 175.820 ;
        RECT 97.130 175.760 97.450 175.775 ;
        RECT 82.870 175.480 85.400 175.620 ;
        RECT 87.025 175.620 87.315 175.665 ;
        RECT 93.910 175.620 94.230 175.680 ;
        RECT 87.025 175.480 94.230 175.620 ;
        RECT 97.680 175.620 97.820 175.820 ;
        RECT 98.050 175.760 98.370 176.020 ;
        RECT 98.510 175.760 98.830 176.020 ;
        RECT 102.280 176.005 102.420 176.160 ;
        RECT 104.030 176.100 104.350 176.160 ;
        RECT 102.205 175.775 102.495 176.005 ;
        RECT 103.110 175.760 103.430 176.020 ;
        RECT 104.580 176.005 104.720 176.160 ;
        RECT 105.500 176.160 109.855 176.300 ;
        RECT 105.500 176.020 105.640 176.160 ;
        RECT 109.565 176.115 109.855 176.160 ;
        RECT 104.505 175.775 104.795 176.005 ;
        RECT 105.410 175.760 105.730 176.020 ;
        RECT 109.090 175.960 109.410 176.020 ;
        RECT 121.600 176.005 121.740 176.840 ;
        RECT 110.025 175.960 110.315 176.005 ;
        RECT 109.090 175.820 110.315 175.960 ;
        RECT 109.090 175.760 109.410 175.820 ;
        RECT 110.025 175.775 110.315 175.820 ;
        RECT 121.525 175.775 121.815 176.005 ;
        RECT 106.790 175.620 107.110 175.680 ;
        RECT 97.680 175.480 107.110 175.620 ;
        RECT 82.870 175.420 83.190 175.480 ;
        RECT 87.025 175.435 87.315 175.480 ;
        RECT 93.910 175.420 94.230 175.480 ;
        RECT 106.790 175.420 107.110 175.480 ;
        RECT 68.150 175.140 71.140 175.280 ;
        RECT 71.370 175.280 71.690 175.340 ;
        RECT 74.590 175.280 74.910 175.340 ;
        RECT 71.370 175.140 74.910 175.280 ;
        RECT 68.150 175.080 68.470 175.140 ;
        RECT 69.990 175.080 70.310 175.140 ;
        RECT 71.370 175.080 71.690 175.140 ;
        RECT 74.590 175.080 74.910 175.140 ;
        RECT 89.770 175.080 90.090 175.340 ;
        RECT 92.085 175.280 92.375 175.325 ;
        RECT 97.130 175.280 97.450 175.340 ;
        RECT 92.085 175.140 97.450 175.280 ;
        RECT 92.085 175.095 92.375 175.140 ;
        RECT 97.130 175.080 97.450 175.140 ;
        RECT 98.050 175.280 98.370 175.340 ;
        RECT 102.190 175.280 102.510 175.340 ;
        RECT 98.050 175.140 102.510 175.280 ;
        RECT 98.050 175.080 98.370 175.140 ;
        RECT 102.190 175.080 102.510 175.140 ;
        RECT 103.570 175.080 103.890 175.340 ;
        RECT 109.550 175.280 109.870 175.340 ;
        RECT 110.485 175.280 110.775 175.325 ;
        RECT 109.550 175.140 110.775 175.280 ;
        RECT 109.550 175.080 109.870 175.140 ;
        RECT 110.485 175.095 110.775 175.140 ;
        RECT 122.445 175.280 122.735 175.325 ;
        RECT 123.810 175.280 124.130 175.340 ;
        RECT 122.445 175.140 124.130 175.280 ;
        RECT 122.445 175.095 122.735 175.140 ;
        RECT 123.810 175.080 124.130 175.140 ;
        RECT 14.260 174.460 126.960 174.940 ;
        RECT 16.170 174.060 16.490 174.320 ;
        RECT 19.850 174.260 20.170 174.320 ;
        RECT 20.785 174.260 21.075 174.305 ;
        RECT 19.850 174.120 21.075 174.260 ;
        RECT 19.850 174.060 20.170 174.120 ;
        RECT 20.785 174.075 21.075 174.120 ;
        RECT 25.845 174.260 26.135 174.305 ;
        RECT 31.350 174.260 31.670 174.320 ;
        RECT 51.605 174.260 51.895 174.305 ;
        RECT 53.430 174.260 53.750 174.320 ;
        RECT 25.845 174.120 31.670 174.260 ;
        RECT 25.845 174.075 26.135 174.120 ;
        RECT 31.350 174.060 31.670 174.120 ;
        RECT 31.900 174.120 44.000 174.260 ;
        RECT 17.105 173.920 17.395 173.965 ;
        RECT 25.370 173.920 25.690 173.980 ;
        RECT 17.105 173.780 25.690 173.920 ;
        RECT 17.105 173.735 17.395 173.780 ;
        RECT 25.370 173.720 25.690 173.780 ;
        RECT 26.750 173.920 27.070 173.980 ;
        RECT 31.900 173.920 32.040 174.120 ;
        RECT 26.750 173.780 32.040 173.920 ;
        RECT 26.750 173.720 27.070 173.780 ;
        RECT 32.270 173.720 32.590 173.980 ;
        RECT 40.550 173.720 40.870 173.980 ;
        RECT 41.025 173.735 41.315 173.965 ;
        RECT 15.725 173.580 16.015 173.625 ;
        RECT 13.960 173.440 16.015 173.580 ;
        RECT 15.725 173.395 16.015 173.440 ;
        RECT 16.630 173.580 16.950 173.640 ;
        RECT 17.565 173.580 17.855 173.625 ;
        RECT 16.630 173.440 17.855 173.580 ;
        RECT 16.630 173.380 16.950 173.440 ;
        RECT 17.565 173.395 17.855 173.440 ;
        RECT 18.485 173.395 18.775 173.625 ;
        RECT 18.930 173.580 19.250 173.640 ;
        RECT 19.865 173.580 20.155 173.625 ;
        RECT 18.930 173.440 20.155 173.580 ;
        RECT 18.560 173.240 18.700 173.395 ;
        RECT 18.930 173.380 19.250 173.440 ;
        RECT 19.865 173.395 20.155 173.440 ;
        RECT 22.625 173.580 22.915 173.625 ;
        RECT 26.290 173.580 26.610 173.640 ;
        RECT 22.625 173.440 26.610 173.580 ;
        RECT 22.625 173.395 22.915 173.440 ;
        RECT 26.290 173.380 26.610 173.440 ;
        RECT 34.570 173.380 34.890 173.640 ;
        RECT 36.870 173.580 37.190 173.640 ;
        RECT 35.120 173.440 37.190 173.580 ;
        RECT 17.180 173.100 18.700 173.240 ;
        RECT 29.050 173.240 29.370 173.300 ;
        RECT 33.665 173.240 33.955 173.285 ;
        RECT 35.120 173.240 35.260 173.440 ;
        RECT 36.870 173.380 37.190 173.440 ;
        RECT 37.345 173.395 37.635 173.625 ;
        RECT 38.250 173.580 38.570 173.640 ;
        RECT 38.725 173.580 39.015 173.625 ;
        RECT 38.250 173.440 39.015 173.580 ;
        RECT 29.050 173.100 35.260 173.240 ;
        RECT 35.505 173.240 35.795 173.285 ;
        RECT 36.410 173.240 36.730 173.300 ;
        RECT 35.505 173.100 36.730 173.240 ;
        RECT 37.420 173.240 37.560 173.395 ;
        RECT 38.250 173.380 38.570 173.440 ;
        RECT 38.725 173.395 39.015 173.440 ;
        RECT 39.170 173.580 39.490 173.640 ;
        RECT 39.645 173.580 39.935 173.625 ;
        RECT 39.170 173.440 39.935 173.580 ;
        RECT 41.100 173.580 41.240 173.735 ;
        RECT 41.100 173.440 41.700 173.580 ;
        RECT 39.170 173.380 39.490 173.440 ;
        RECT 39.645 173.395 39.935 173.440 ;
        RECT 41.560 173.300 41.700 173.440 ;
        RECT 41.930 173.380 42.250 173.640 ;
        RECT 42.865 173.580 43.155 173.625 ;
        RECT 43.310 173.580 43.630 173.640 ;
        RECT 43.860 173.625 44.000 174.120 ;
        RECT 51.605 174.120 53.750 174.260 ;
        RECT 51.605 174.075 51.895 174.120 ;
        RECT 53.430 174.060 53.750 174.120 ;
        RECT 53.905 174.260 54.195 174.305 ;
        RECT 54.350 174.260 54.670 174.320 ;
        RECT 53.905 174.120 54.670 174.260 ;
        RECT 53.905 174.075 54.195 174.120 ;
        RECT 54.350 174.060 54.670 174.120 ;
        RECT 58.965 174.260 59.255 174.305 ;
        RECT 59.410 174.260 59.730 174.320 ;
        RECT 58.965 174.120 59.730 174.260 ;
        RECT 58.965 174.075 59.255 174.120 ;
        RECT 59.410 174.060 59.730 174.120 ;
        RECT 60.790 174.060 61.110 174.320 ;
        RECT 72.765 174.260 73.055 174.305 ;
        RECT 73.670 174.260 73.990 174.320 ;
        RECT 72.765 174.120 73.990 174.260 ;
        RECT 72.765 174.075 73.055 174.120 ;
        RECT 52.985 173.920 53.275 173.965 ;
        RECT 58.505 173.920 58.795 173.965 ;
        RECT 60.880 173.920 61.020 174.060 ;
        RECT 68.150 173.920 68.470 173.980 ;
        RECT 51.220 173.780 55.040 173.920 ;
        RECT 42.865 173.440 43.630 173.580 ;
        RECT 42.865 173.395 43.155 173.440 ;
        RECT 43.310 173.380 43.630 173.440 ;
        RECT 43.785 173.395 44.075 173.625 ;
        RECT 47.450 173.380 47.770 173.640 ;
        RECT 51.220 173.625 51.360 173.780 ;
        RECT 52.985 173.735 53.275 173.780 ;
        RECT 54.900 173.625 55.040 173.780 ;
        RECT 55.820 173.780 57.800 173.920 ;
        RECT 55.820 173.625 55.960 173.780 ;
        RECT 50.685 173.580 50.975 173.625 ;
        RECT 51.145 173.580 51.435 173.625 ;
        RECT 50.685 173.440 51.435 173.580 ;
        RECT 50.685 173.395 50.975 173.440 ;
        RECT 51.145 173.395 51.435 173.440 ;
        RECT 52.065 173.395 52.355 173.625 ;
        RECT 53.485 173.530 53.775 173.575 ;
        RECT 41.010 173.240 41.330 173.300 ;
        RECT 37.420 173.100 41.330 173.240 ;
        RECT 17.180 172.945 17.320 173.100 ;
        RECT 29.050 173.040 29.370 173.100 ;
        RECT 33.665 173.055 33.955 173.100 ;
        RECT 35.505 173.055 35.795 173.100 ;
        RECT 36.410 173.040 36.730 173.100 ;
        RECT 41.010 173.040 41.330 173.100 ;
        RECT 41.470 173.040 41.790 173.300 ;
        RECT 42.020 173.240 42.160 173.380 ;
        RECT 43.400 173.240 43.540 173.380 ;
        RECT 42.020 173.100 42.850 173.240 ;
        RECT 43.400 173.100 50.440 173.240 ;
        RECT 17.105 172.715 17.395 172.945 ;
        RECT 42.710 172.900 42.850 173.100 ;
        RECT 45.610 172.900 45.930 172.960 ;
        RECT 42.710 172.760 45.930 172.900 ;
        RECT 45.610 172.700 45.930 172.760 ;
        RECT 21.705 172.560 21.995 172.605 ;
        RECT 22.610 172.560 22.930 172.620 ;
        RECT 21.705 172.420 22.930 172.560 ;
        RECT 21.705 172.375 21.995 172.420 ;
        RECT 22.610 172.360 22.930 172.420 ;
        RECT 24.450 172.560 24.770 172.620 ;
        RECT 37.790 172.560 38.110 172.620 ;
        RECT 24.450 172.420 38.110 172.560 ;
        RECT 24.450 172.360 24.770 172.420 ;
        RECT 37.790 172.360 38.110 172.420 ;
        RECT 38.265 172.560 38.555 172.605 ;
        RECT 43.310 172.560 43.630 172.620 ;
        RECT 38.265 172.420 43.630 172.560 ;
        RECT 38.265 172.375 38.555 172.420 ;
        RECT 43.310 172.360 43.630 172.420 ;
        RECT 49.750 172.360 50.070 172.620 ;
        RECT 50.300 172.560 50.440 173.100 ;
        RECT 52.140 172.900 52.280 173.395 ;
        RECT 53.485 173.390 54.120 173.530 ;
        RECT 54.825 173.395 55.115 173.625 ;
        RECT 55.745 173.395 56.035 173.625 ;
        RECT 56.665 173.580 56.955 173.625 ;
        RECT 57.110 173.580 57.430 173.640 ;
        RECT 57.660 173.625 57.800 173.780 ;
        RECT 58.505 173.780 61.020 173.920 ;
        RECT 63.640 173.780 68.470 173.920 ;
        RECT 58.505 173.735 58.795 173.780 ;
        RECT 63.640 173.640 63.780 173.780 ;
        RECT 68.150 173.720 68.470 173.780 ;
        RECT 69.070 173.920 69.390 173.980 ;
        RECT 70.925 173.920 71.215 173.965 ;
        RECT 69.070 173.780 71.215 173.920 ;
        RECT 69.070 173.720 69.390 173.780 ;
        RECT 70.925 173.735 71.215 173.780 ;
        RECT 56.665 173.440 57.430 173.580 ;
        RECT 56.665 173.395 56.955 173.440 ;
        RECT 53.485 173.345 53.775 173.390 ;
        RECT 53.980 173.240 54.120 173.390 ;
        RECT 55.270 173.240 55.590 173.300 ;
        RECT 56.740 173.240 56.880 173.395 ;
        RECT 57.110 173.380 57.430 173.440 ;
        RECT 57.585 173.395 57.875 173.625 ;
        RECT 58.030 173.580 58.350 173.640 ;
        RECT 59.885 173.580 60.175 173.625 ;
        RECT 58.030 173.440 60.175 173.580 ;
        RECT 53.980 173.100 56.880 173.240 ;
        RECT 57.660 173.240 57.800 173.395 ;
        RECT 58.030 173.380 58.350 173.440 ;
        RECT 59.885 173.395 60.175 173.440 ;
        RECT 60.805 173.580 61.095 173.625 ;
        RECT 61.250 173.580 61.570 173.640 ;
        RECT 60.805 173.440 61.570 173.580 ;
        RECT 60.805 173.395 61.095 173.440 ;
        RECT 60.880 173.240 61.020 173.395 ;
        RECT 61.250 173.380 61.570 173.440 ;
        RECT 63.550 173.380 63.870 173.640 ;
        RECT 64.945 173.580 65.235 173.625 ;
        RECT 66.325 173.580 66.615 173.625 ;
        RECT 64.945 173.440 66.615 173.580 ;
        RECT 64.945 173.395 65.235 173.440 ;
        RECT 66.325 173.395 66.615 173.440 ;
        RECT 57.660 173.100 61.020 173.240 ;
        RECT 66.400 173.240 66.540 173.395 ;
        RECT 66.770 173.380 67.090 173.640 ;
        RECT 67.705 173.580 67.995 173.625 ;
        RECT 71.370 173.580 71.690 173.640 ;
        RECT 67.705 173.440 71.690 173.580 ;
        RECT 67.705 173.395 67.995 173.440 ;
        RECT 71.370 173.380 71.690 173.440 ;
        RECT 71.830 173.380 72.150 173.640 ;
        RECT 73.300 173.625 73.440 174.120 ;
        RECT 73.670 174.060 73.990 174.120 ;
        RECT 75.510 174.060 75.830 174.320 ;
        RECT 76.445 174.260 76.735 174.305 ;
        RECT 79.190 174.260 79.510 174.320 ;
        RECT 76.445 174.120 79.510 174.260 ;
        RECT 76.445 174.075 76.735 174.120 ;
        RECT 79.190 174.060 79.510 174.120 ;
        RECT 83.330 174.260 83.650 174.320 ;
        RECT 83.805 174.260 84.095 174.305 ;
        RECT 85.645 174.260 85.935 174.305 ;
        RECT 83.330 174.120 85.935 174.260 ;
        RECT 83.330 174.060 83.650 174.120 ;
        RECT 83.805 174.075 84.095 174.120 ;
        RECT 85.645 174.075 85.935 174.120 ;
        RECT 93.910 174.060 94.230 174.320 ;
        RECT 94.385 174.260 94.675 174.305 ;
        RECT 94.830 174.260 95.150 174.320 ;
        RECT 94.385 174.120 95.150 174.260 ;
        RECT 94.385 174.075 94.675 174.120 ;
        RECT 75.600 173.920 75.740 174.060 ;
        RECT 73.760 173.780 75.740 173.920 ;
        RECT 73.225 173.395 73.515 173.625 ;
        RECT 69.990 173.240 70.310 173.300 ;
        RECT 66.400 173.100 70.310 173.240 ;
        RECT 71.920 173.240 72.060 173.380 ;
        RECT 73.760 173.240 73.900 173.780 ;
        RECT 78.730 173.720 79.050 173.980 ;
        RECT 92.085 173.920 92.375 173.965 ;
        RECT 94.460 173.920 94.600 174.075 ;
        RECT 94.830 174.060 95.150 174.120 ;
        RECT 96.225 174.260 96.515 174.305 ;
        RECT 98.510 174.260 98.830 174.320 ;
        RECT 96.225 174.120 98.830 174.260 ;
        RECT 96.225 174.075 96.515 174.120 ;
        RECT 98.510 174.060 98.830 174.120 ;
        RECT 100.365 174.260 100.655 174.305 ;
        RECT 102.665 174.260 102.955 174.305 ;
        RECT 103.570 174.260 103.890 174.320 ;
        RECT 100.365 174.120 103.890 174.260 ;
        RECT 100.365 174.075 100.655 174.120 ;
        RECT 102.665 174.075 102.955 174.120 ;
        RECT 103.570 174.060 103.890 174.120 ;
        RECT 107.725 174.260 108.015 174.305 ;
        RECT 109.550 174.260 109.870 174.320 ;
        RECT 107.725 174.120 109.870 174.260 ;
        RECT 107.725 174.075 108.015 174.120 ;
        RECT 109.550 174.060 109.870 174.120 ;
        RECT 124.745 174.260 125.035 174.305 ;
        RECT 130.250 174.260 130.570 174.320 ;
        RECT 124.745 174.120 130.570 174.260 ;
        RECT 124.745 174.075 125.035 174.120 ;
        RECT 130.250 174.060 130.570 174.120 ;
        RECT 79.280 173.780 84.940 173.920 ;
        RECT 75.050 173.580 75.370 173.640 ;
        RECT 75.540 173.580 75.830 173.625 ;
        RECT 79.280 173.580 79.420 173.780 ;
        RECT 75.050 173.440 75.830 173.580 ;
        RECT 75.050 173.380 75.370 173.440 ;
        RECT 75.540 173.395 75.830 173.440 ;
        RECT 76.520 173.440 79.420 173.580 ;
        RECT 71.920 173.100 73.900 173.240 ;
        RECT 74.130 173.240 74.450 173.300 ;
        RECT 76.520 173.240 76.660 173.440 ;
        RECT 79.650 173.380 79.970 173.640 ;
        RECT 80.110 173.580 80.430 173.640 ;
        RECT 81.045 173.580 81.335 173.625 ;
        RECT 80.110 173.440 81.335 173.580 ;
        RECT 80.110 173.380 80.430 173.440 ;
        RECT 81.045 173.395 81.335 173.440 ;
        RECT 81.490 173.380 81.810 173.640 ;
        RECT 82.885 173.580 83.175 173.625 ;
        RECT 82.885 173.440 84.020 173.580 ;
        RECT 82.885 173.395 83.175 173.440 ;
        RECT 74.130 173.100 76.660 173.240 ;
        RECT 55.270 173.040 55.590 173.100 ;
        RECT 57.660 172.900 57.800 173.100 ;
        RECT 69.990 173.040 70.310 173.100 ;
        RECT 74.130 173.040 74.450 173.100 ;
        RECT 52.140 172.760 57.800 172.900 ;
        RECT 58.950 172.900 59.270 172.960 ;
        RECT 64.485 172.900 64.775 172.945 ;
        RECT 58.950 172.760 64.775 172.900 ;
        RECT 58.950 172.700 59.270 172.760 ;
        RECT 64.485 172.715 64.775 172.760 ;
        RECT 67.690 172.900 68.010 172.960 ;
        RECT 73.685 172.900 73.975 172.945 ;
        RECT 67.690 172.760 73.975 172.900 ;
        RECT 67.690 172.700 68.010 172.760 ;
        RECT 73.685 172.715 73.975 172.760 ;
        RECT 80.585 172.900 80.875 172.945 ;
        RECT 82.885 172.900 83.175 172.945 ;
        RECT 80.585 172.760 83.175 172.900 ;
        RECT 83.880 172.900 84.020 173.440 ;
        RECT 84.250 173.380 84.570 173.640 ;
        RECT 84.800 173.625 84.940 173.780 ;
        RECT 92.085 173.780 94.600 173.920 ;
        RECT 97.590 173.920 97.910 173.980 ;
        RECT 101.270 173.920 101.590 173.980 ;
        RECT 101.745 173.920 102.035 173.965 ;
        RECT 97.590 173.780 98.740 173.920 ;
        RECT 92.085 173.735 92.375 173.780 ;
        RECT 97.590 173.720 97.910 173.780 ;
        RECT 84.725 173.395 85.015 173.625 ;
        RECT 85.630 173.580 85.950 173.640 ;
        RECT 91.165 173.580 91.455 173.625 ;
        RECT 85.630 173.440 91.455 173.580 ;
        RECT 85.630 173.380 85.950 173.440 ;
        RECT 91.165 173.395 91.455 173.440 ;
        RECT 96.670 173.380 96.990 173.640 ;
        RECT 98.050 173.380 98.370 173.640 ;
        RECT 98.600 173.625 98.740 173.780 ;
        RECT 101.270 173.780 102.035 173.920 ;
        RECT 101.270 173.720 101.590 173.780 ;
        RECT 101.745 173.735 102.035 173.780 ;
        RECT 106.330 173.920 106.650 173.980 ;
        RECT 106.805 173.920 107.095 173.965 ;
        RECT 106.330 173.780 107.095 173.920 ;
        RECT 106.330 173.720 106.650 173.780 ;
        RECT 106.805 173.735 107.095 173.780 ;
        RECT 109.090 173.920 109.410 173.980 ;
        RECT 110.025 173.920 110.315 173.965 ;
        RECT 109.090 173.780 110.315 173.920 ;
        RECT 109.090 173.720 109.410 173.780 ;
        RECT 110.025 173.735 110.315 173.780 ;
        RECT 98.525 173.395 98.815 173.625 ;
        RECT 99.445 173.580 99.735 173.625 ;
        RECT 99.905 173.580 100.195 173.625 ;
        RECT 99.445 173.440 100.195 173.580 ;
        RECT 99.445 173.395 99.735 173.440 ;
        RECT 99.905 173.395 100.195 173.440 ;
        RECT 103.110 173.380 103.430 173.640 ;
        RECT 104.950 173.580 105.270 173.640 ;
        RECT 105.885 173.580 106.175 173.625 ;
        RECT 104.950 173.440 106.175 173.580 ;
        RECT 104.950 173.380 105.270 173.440 ;
        RECT 105.885 173.395 106.175 173.440 ;
        RECT 115.530 173.580 115.850 173.640 ;
        RECT 121.525 173.580 121.815 173.625 ;
        RECT 115.530 173.440 121.815 173.580 ;
        RECT 115.530 173.380 115.850 173.440 ;
        RECT 121.525 173.395 121.815 173.440 ;
        RECT 123.810 173.380 124.130 173.640 ;
        RECT 93.450 173.040 93.770 173.300 ;
        RECT 97.130 173.040 97.450 173.300 ;
        RECT 105.410 173.240 105.730 173.300 ;
        RECT 108.645 173.240 108.935 173.285 ;
        RECT 105.410 173.100 108.935 173.240 ;
        RECT 105.410 173.040 105.730 173.100 ;
        RECT 108.645 173.055 108.935 173.100 ;
        RECT 101.285 172.900 101.575 172.945 ;
        RECT 83.880 172.760 101.575 172.900 ;
        RECT 80.585 172.715 80.875 172.760 ;
        RECT 82.885 172.715 83.175 172.760 ;
        RECT 101.285 172.715 101.575 172.760 ;
        RECT 59.040 172.560 59.180 172.700 ;
        RECT 50.300 172.420 59.180 172.560 ;
        RECT 62.630 172.360 62.950 172.620 ;
        RECT 69.070 172.560 69.390 172.620 ;
        RECT 71.830 172.560 72.150 172.620 ;
        RECT 69.070 172.420 72.150 172.560 ;
        RECT 69.070 172.360 69.390 172.420 ;
        RECT 71.830 172.360 72.150 172.420 ;
        RECT 82.410 172.360 82.730 172.620 ;
        RECT 99.430 172.560 99.750 172.620 ;
        RECT 101.745 172.560 102.035 172.605 ;
        RECT 99.430 172.420 102.035 172.560 ;
        RECT 99.430 172.360 99.750 172.420 ;
        RECT 101.745 172.375 102.035 172.420 ;
        RECT 111.850 172.360 112.170 172.620 ;
        RECT 122.430 172.360 122.750 172.620 ;
        RECT 14.260 171.740 126.960 172.220 ;
        RECT 17.550 171.340 17.870 171.600 ;
        RECT 18.010 171.340 18.330 171.600 ;
        RECT 21.690 171.540 22.010 171.600 ;
        RECT 19.480 171.400 22.010 171.540 ;
        RECT 16.185 171.200 16.475 171.245 ;
        RECT 18.930 171.200 19.250 171.260 ;
        RECT 16.185 171.060 19.250 171.200 ;
        RECT 16.185 171.015 16.475 171.060 ;
        RECT 18.930 171.000 19.250 171.060 ;
        RECT 16.645 170.860 16.935 170.905 ;
        RECT 19.480 170.860 19.620 171.400 ;
        RECT 21.690 171.340 22.010 171.400 ;
        RECT 22.165 171.540 22.455 171.585 ;
        RECT 24.910 171.540 25.230 171.600 ;
        RECT 22.165 171.400 25.230 171.540 ;
        RECT 22.165 171.355 22.455 171.400 ;
        RECT 24.910 171.340 25.230 171.400 ;
        RECT 25.830 171.340 26.150 171.600 ;
        RECT 29.050 171.340 29.370 171.600 ;
        RECT 29.985 171.540 30.275 171.585 ;
        RECT 35.950 171.540 36.270 171.600 ;
        RECT 36.885 171.540 37.175 171.585 ;
        RECT 29.985 171.400 35.720 171.540 ;
        RECT 29.985 171.355 30.275 171.400 ;
        RECT 20.310 171.200 20.630 171.260 ;
        RECT 31.365 171.200 31.655 171.245 ;
        RECT 34.570 171.200 34.890 171.260 ;
        RECT 20.310 171.060 31.655 171.200 ;
        RECT 20.310 171.000 20.630 171.060 ;
        RECT 31.365 171.015 31.655 171.060 ;
        RECT 32.360 171.060 34.890 171.200 ;
        RECT 35.580 171.200 35.720 171.400 ;
        RECT 35.950 171.400 37.175 171.540 ;
        RECT 35.950 171.340 36.270 171.400 ;
        RECT 36.885 171.355 37.175 171.400 ;
        RECT 37.790 171.540 38.110 171.600 ;
        RECT 37.790 171.400 39.860 171.540 ;
        RECT 37.790 171.340 38.110 171.400 ;
        RECT 39.170 171.200 39.490 171.260 ;
        RECT 35.580 171.060 39.490 171.200 ;
        RECT 39.720 171.200 39.860 171.400 ;
        RECT 41.010 171.340 41.330 171.600 ;
        RECT 46.085 171.540 46.375 171.585 ;
        RECT 48.830 171.540 49.150 171.600 ;
        RECT 41.560 171.400 48.600 171.540 ;
        RECT 41.560 171.200 41.700 171.400 ;
        RECT 46.085 171.355 46.375 171.400 ;
        RECT 39.720 171.060 41.700 171.200 ;
        RECT 42.865 171.200 43.155 171.245 ;
        RECT 46.530 171.200 46.850 171.260 ;
        RECT 42.865 171.060 46.850 171.200 ;
        RECT 48.460 171.200 48.600 171.400 ;
        RECT 48.830 171.400 52.740 171.540 ;
        RECT 48.830 171.340 49.150 171.400 ;
        RECT 49.290 171.200 49.610 171.260 ;
        RECT 48.460 171.060 49.610 171.200 ;
        RECT 16.645 170.720 19.620 170.860 ;
        RECT 19.865 170.860 20.155 170.905 ;
        RECT 24.005 170.860 24.295 170.905 ;
        RECT 19.865 170.720 24.295 170.860 ;
        RECT 16.645 170.675 16.935 170.720 ;
        RECT 19.020 170.565 19.160 170.720 ;
        RECT 19.865 170.675 20.155 170.720 ;
        RECT 24.005 170.675 24.295 170.720 ;
        RECT 26.290 170.660 26.610 170.920 ;
        RECT 18.945 170.335 19.235 170.565 ;
        RECT 19.405 170.335 19.695 170.565 ;
        RECT 15.725 170.180 16.015 170.225 ;
        RECT 16.630 170.180 16.950 170.240 ;
        RECT 15.725 170.040 16.950 170.180 ;
        RECT 15.725 169.995 16.015 170.040 ;
        RECT 16.630 169.980 16.950 170.040 ;
        RECT 17.565 170.180 17.855 170.225 ;
        RECT 18.470 170.180 18.790 170.240 ;
        RECT 19.480 170.180 19.620 170.335 ;
        RECT 20.310 170.320 20.630 170.580 ;
        RECT 23.070 170.320 23.390 170.580 ;
        RECT 24.910 170.320 25.230 170.580 ;
        RECT 26.750 170.320 27.070 170.580 ;
        RECT 28.130 170.320 28.450 170.580 ;
        RECT 32.360 170.565 32.500 171.060 ;
        RECT 34.570 171.000 34.890 171.060 ;
        RECT 39.170 171.000 39.490 171.060 ;
        RECT 42.865 171.015 43.155 171.060 ;
        RECT 46.530 171.000 46.850 171.060 ;
        RECT 49.290 171.000 49.610 171.060 ;
        RECT 50.685 171.200 50.975 171.245 ;
        RECT 52.050 171.200 52.370 171.260 ;
        RECT 50.685 171.060 52.370 171.200 ;
        RECT 52.600 171.200 52.740 171.400 ;
        RECT 54.810 171.340 55.130 171.600 ;
        RECT 67.705 171.540 67.995 171.585 ;
        RECT 55.360 171.400 67.995 171.540 ;
        RECT 55.360 171.200 55.500 171.400 ;
        RECT 67.705 171.355 67.995 171.400 ;
        RECT 68.610 171.540 68.930 171.600 ;
        RECT 69.085 171.540 69.375 171.585 ;
        RECT 68.610 171.400 69.375 171.540 ;
        RECT 68.610 171.340 68.930 171.400 ;
        RECT 69.085 171.355 69.375 171.400 ;
        RECT 69.990 171.340 70.310 171.600 ;
        RECT 74.130 171.540 74.450 171.600 ;
        RECT 75.985 171.540 76.275 171.585 ;
        RECT 74.130 171.400 76.275 171.540 ;
        RECT 74.130 171.340 74.450 171.400 ;
        RECT 75.985 171.355 76.275 171.400 ;
        RECT 85.630 171.340 85.950 171.600 ;
        RECT 103.110 171.540 103.430 171.600 ;
        RECT 110.025 171.540 110.315 171.585 ;
        RECT 103.110 171.400 110.315 171.540 ;
        RECT 103.110 171.340 103.430 171.400 ;
        RECT 110.025 171.355 110.315 171.400 ;
        RECT 111.850 171.540 112.170 171.600 ;
        RECT 112.325 171.540 112.615 171.585 ;
        RECT 111.850 171.400 112.615 171.540 ;
        RECT 111.850 171.340 112.170 171.400 ;
        RECT 112.325 171.355 112.615 171.400 ;
        RECT 124.745 171.540 125.035 171.585 ;
        RECT 130.250 171.540 130.570 171.600 ;
        RECT 124.745 171.400 130.570 171.540 ;
        RECT 124.745 171.355 125.035 171.400 ;
        RECT 130.250 171.340 130.570 171.400 ;
        RECT 52.600 171.060 55.500 171.200 ;
        RECT 50.685 171.015 50.975 171.060 ;
        RECT 52.050 171.000 52.370 171.060 ;
        RECT 58.045 171.015 58.335 171.245 ;
        RECT 71.830 171.200 72.150 171.260 ;
        RECT 104.950 171.200 105.270 171.260 ;
        RECT 71.830 171.060 105.270 171.200 ;
        RECT 33.205 170.860 33.495 170.905 ;
        RECT 33.205 170.720 38.020 170.860 ;
        RECT 33.205 170.675 33.495 170.720 ;
        RECT 29.525 170.335 29.815 170.565 ;
        RECT 32.285 170.335 32.575 170.565 ;
        RECT 19.850 170.180 20.170 170.240 ;
        RECT 17.565 170.040 20.170 170.180 ;
        RECT 17.565 169.995 17.855 170.040 ;
        RECT 18.470 169.980 18.790 170.040 ;
        RECT 19.850 169.980 20.170 170.040 ;
        RECT 29.600 170.180 29.740 170.335 ;
        RECT 33.280 170.180 33.420 170.675 ;
        RECT 33.650 170.320 33.970 170.580 ;
        RECT 37.880 170.565 38.020 170.720 ;
        RECT 37.805 170.335 38.095 170.565 ;
        RECT 38.250 170.320 38.570 170.580 ;
        RECT 39.260 170.565 39.400 171.000 ;
        RECT 39.630 170.860 39.950 170.920 ;
        RECT 39.630 170.720 53.660 170.860 ;
        RECT 39.630 170.660 39.950 170.720 ;
        RECT 39.185 170.520 39.475 170.565 ;
        RECT 41.945 170.520 42.235 170.565 ;
        RECT 39.185 170.380 42.235 170.520 ;
        RECT 39.185 170.335 39.475 170.380 ;
        RECT 41.945 170.335 42.235 170.380 ;
        RECT 43.310 170.320 43.630 170.580 ;
        RECT 43.770 170.520 44.090 170.580 ;
        RECT 45.165 170.520 45.455 170.565 ;
        RECT 43.770 170.380 45.455 170.520 ;
        RECT 43.770 170.320 44.090 170.380 ;
        RECT 45.165 170.335 45.455 170.380 ;
        RECT 46.530 170.320 46.850 170.580 ;
        RECT 49.750 170.320 50.070 170.580 ;
        RECT 53.520 170.565 53.660 170.720 ;
        RECT 52.525 170.335 52.815 170.565 ;
        RECT 53.445 170.335 53.735 170.565 ;
        RECT 55.745 170.520 56.035 170.565 ;
        RECT 57.110 170.520 57.430 170.580 ;
        RECT 55.745 170.380 57.430 170.520 ;
        RECT 55.745 170.335 56.035 170.380 ;
        RECT 29.600 170.040 33.420 170.180 ;
        RECT 38.340 170.180 38.480 170.320 ;
        RECT 40.105 170.180 40.395 170.225 ;
        RECT 38.340 170.040 40.395 170.180 ;
        RECT 27.685 169.840 27.975 169.885 ;
        RECT 29.600 169.840 29.740 170.040 ;
        RECT 40.105 169.995 40.395 170.040 ;
        RECT 42.850 170.180 43.170 170.240 ;
        RECT 52.600 170.180 52.740 170.335 ;
        RECT 57.110 170.320 57.430 170.380 ;
        RECT 57.585 170.520 57.875 170.565 ;
        RECT 58.120 170.520 58.260 171.015 ;
        RECT 71.830 171.000 72.150 171.060 ;
        RECT 104.950 171.000 105.270 171.060 ;
        RECT 65.865 170.860 66.155 170.905 ;
        RECT 66.770 170.860 67.090 170.920 ;
        RECT 65.865 170.720 67.090 170.860 ;
        RECT 65.865 170.675 66.155 170.720 ;
        RECT 66.770 170.660 67.090 170.720 ;
        RECT 108.170 170.860 108.490 170.920 ;
        RECT 123.365 170.860 123.655 170.905 ;
        RECT 125.650 170.860 125.970 170.920 ;
        RECT 108.170 170.720 111.620 170.860 ;
        RECT 108.170 170.660 108.490 170.720 ;
        RECT 57.585 170.380 58.260 170.520 ;
        RECT 57.585 170.335 57.875 170.380 ;
        RECT 58.950 170.320 59.270 170.580 ;
        RECT 61.725 170.520 62.015 170.565 ;
        RECT 62.630 170.520 62.950 170.580 ;
        RECT 61.725 170.380 62.950 170.520 ;
        RECT 61.725 170.335 62.015 170.380 ;
        RECT 62.630 170.320 62.950 170.380 ;
        RECT 67.245 170.520 67.535 170.565 ;
        RECT 67.690 170.520 68.010 170.580 ;
        RECT 67.245 170.380 68.010 170.520 ;
        RECT 67.245 170.335 67.535 170.380 ;
        RECT 67.690 170.320 68.010 170.380 ;
        RECT 68.610 170.320 68.930 170.580 ;
        RECT 70.910 170.320 71.230 170.580 ;
        RECT 72.765 170.335 73.055 170.565 ;
        RECT 76.905 170.520 77.195 170.565 ;
        RECT 77.350 170.520 77.670 170.580 ;
        RECT 76.905 170.380 77.670 170.520 ;
        RECT 76.905 170.335 77.195 170.380 ;
        RECT 42.850 170.040 52.740 170.180 ;
        RECT 56.190 170.180 56.510 170.240 ;
        RECT 72.840 170.180 72.980 170.335 ;
        RECT 77.350 170.320 77.670 170.380 ;
        RECT 81.965 170.520 82.255 170.565 ;
        RECT 82.410 170.520 82.730 170.580 ;
        RECT 81.965 170.380 82.730 170.520 ;
        RECT 81.965 170.335 82.255 170.380 ;
        RECT 82.410 170.320 82.730 170.380 ;
        RECT 86.565 170.520 86.855 170.565 ;
        RECT 87.010 170.520 87.330 170.580 ;
        RECT 86.565 170.380 87.330 170.520 ;
        RECT 86.565 170.335 86.855 170.380 ;
        RECT 87.010 170.320 87.330 170.380 ;
        RECT 108.630 170.520 108.950 170.580 ;
        RECT 111.480 170.565 111.620 170.720 ;
        RECT 123.365 170.720 125.970 170.860 ;
        RECT 123.365 170.675 123.655 170.720 ;
        RECT 125.650 170.660 125.970 170.720 ;
        RECT 110.945 170.520 111.235 170.565 ;
        RECT 108.630 170.380 111.235 170.520 ;
        RECT 108.630 170.320 108.950 170.380 ;
        RECT 110.945 170.335 111.235 170.380 ;
        RECT 111.405 170.335 111.695 170.565 ;
        RECT 112.785 170.520 113.075 170.565 ;
        RECT 115.530 170.520 115.850 170.580 ;
        RECT 112.785 170.380 115.850 170.520 ;
        RECT 112.785 170.335 113.075 170.380 ;
        RECT 115.530 170.320 115.850 170.380 ;
        RECT 122.430 170.520 122.750 170.580 ;
        RECT 123.825 170.520 124.115 170.565 ;
        RECT 122.430 170.380 124.115 170.520 ;
        RECT 122.430 170.320 122.750 170.380 ;
        RECT 123.825 170.335 124.115 170.380 ;
        RECT 56.190 170.040 72.980 170.180 ;
        RECT 42.850 169.980 43.170 170.040 ;
        RECT 56.190 169.980 56.510 170.040 ;
        RECT 27.685 169.700 29.740 169.840 ;
        RECT 34.585 169.840 34.875 169.885 ;
        RECT 35.490 169.840 35.810 169.900 ;
        RECT 34.585 169.700 35.810 169.840 ;
        RECT 27.685 169.655 27.975 169.700 ;
        RECT 34.585 169.655 34.875 169.700 ;
        RECT 35.490 169.640 35.810 169.700 ;
        RECT 44.245 169.840 44.535 169.885 ;
        RECT 45.150 169.840 45.470 169.900 ;
        RECT 44.245 169.700 45.470 169.840 ;
        RECT 44.245 169.655 44.535 169.700 ;
        RECT 45.150 169.640 45.470 169.700 ;
        RECT 47.465 169.840 47.755 169.885 ;
        RECT 48.370 169.840 48.690 169.900 ;
        RECT 47.465 169.700 48.690 169.840 ;
        RECT 47.465 169.655 47.755 169.700 ;
        RECT 48.370 169.640 48.690 169.700 ;
        RECT 51.590 169.640 51.910 169.900 ;
        RECT 54.365 169.840 54.655 169.885 ;
        RECT 54.810 169.840 55.130 169.900 ;
        RECT 54.365 169.700 55.130 169.840 ;
        RECT 54.365 169.655 54.655 169.700 ;
        RECT 54.810 169.640 55.130 169.700 ;
        RECT 56.665 169.840 56.955 169.885 ;
        RECT 58.030 169.840 58.350 169.900 ;
        RECT 56.665 169.700 58.350 169.840 ;
        RECT 56.665 169.655 56.955 169.700 ;
        RECT 58.030 169.640 58.350 169.700 ;
        RECT 60.805 169.840 61.095 169.885 ;
        RECT 64.470 169.840 64.790 169.900 ;
        RECT 60.805 169.700 64.790 169.840 ;
        RECT 60.805 169.655 61.095 169.700 ;
        RECT 64.470 169.640 64.790 169.700 ;
        RECT 73.685 169.840 73.975 169.885 ;
        RECT 74.130 169.840 74.450 169.900 ;
        RECT 73.685 169.700 74.450 169.840 ;
        RECT 73.685 169.655 73.975 169.700 ;
        RECT 74.130 169.640 74.450 169.700 ;
        RECT 82.885 169.840 83.175 169.885 ;
        RECT 83.790 169.840 84.110 169.900 ;
        RECT 82.885 169.700 84.110 169.840 ;
        RECT 82.885 169.655 83.175 169.700 ;
        RECT 83.790 169.640 84.110 169.700 ;
        RECT 14.260 169.020 126.960 169.500 ;
        RECT 18.930 168.820 19.250 168.880 ;
        RECT 24.450 168.820 24.770 168.880 ;
        RECT 18.930 168.680 24.770 168.820 ;
        RECT 18.930 168.620 19.250 168.680 ;
        RECT 24.450 168.620 24.770 168.680 ;
        RECT 24.910 168.820 25.230 168.880 ;
        RECT 50.210 168.820 50.530 168.880 ;
        RECT 24.910 168.680 50.530 168.820 ;
        RECT 24.910 168.620 25.230 168.680 ;
        RECT 50.210 168.620 50.530 168.680 ;
        RECT 57.110 168.820 57.430 168.880 ;
        RECT 61.250 168.820 61.570 168.880 ;
        RECT 57.110 168.680 61.570 168.820 ;
        RECT 57.110 168.620 57.430 168.680 ;
        RECT 61.250 168.620 61.570 168.680 ;
        RECT 29.050 168.480 29.370 168.540 ;
        RECT 47.450 168.480 47.770 168.540 ;
        RECT 29.050 168.340 47.770 168.480 ;
        RECT 29.050 168.280 29.370 168.340 ;
        RECT 47.450 168.280 47.770 168.340 ;
        RECT 16.630 157.260 16.950 157.320 ;
        RECT 51.130 157.260 51.450 157.320 ;
        RECT 16.630 157.120 51.450 157.260 ;
        RECT 16.630 157.060 16.950 157.120 ;
        RECT 51.130 157.060 51.450 157.120 ;
        RECT 129.140 74.465 129.445 74.540 ;
        RECT 130.730 74.505 131.035 74.550 ;
        RECT 129.135 74.280 129.445 74.465 ;
        RECT 130.695 74.290 131.035 74.505 ;
        RECT 132.305 74.465 132.610 74.550 ;
        RECT 132.295 74.290 132.610 74.465 ;
        RECT 129.135 74.235 129.425 74.280 ;
        RECT 130.695 74.245 131.005 74.290 ;
        RECT 130.715 74.235 131.005 74.245 ;
        RECT 132.295 74.235 132.585 74.290 ;
        RECT 133.870 74.280 134.175 74.540 ;
        RECT 133.875 74.235 134.165 74.280 ;
        RECT 128.945 73.980 129.175 74.030 ;
        RECT 77.445 70.840 78.085 70.845 ;
        RECT 50.550 70.835 78.085 70.840 ;
        RECT 81.075 70.840 81.805 70.845 ;
        RECT 81.075 70.835 110.655 70.840 ;
        RECT 50.550 70.300 110.655 70.835 ;
        RECT 50.245 69.600 110.655 70.300 ;
        RECT 50.245 69.435 75.895 69.600 ;
        RECT 76.885 69.435 110.655 69.600 ;
        RECT 46.890 68.900 47.480 68.950 ;
        RECT 48.710 68.900 49.300 68.950 ;
        RECT 46.890 66.945 49.300 68.900 ;
        RECT 50.245 68.670 50.705 69.435 ;
        RECT 51.205 68.920 51.520 69.210 ;
        RECT 51.020 68.670 51.250 68.715 ;
        RECT 50.245 68.000 51.250 68.670 ;
        RECT 46.890 66.845 47.480 66.945 ;
        RECT 48.710 66.845 49.300 66.945 ;
        RECT 46.890 65.940 47.480 66.265 ;
        RECT 48.710 65.960 49.300 66.265 ;
        RECT 46.870 60.920 47.495 65.940 ;
        RECT 48.685 60.940 49.310 65.960 ;
        RECT 50.655 62.795 51.250 68.000 ;
        RECT 51.020 62.715 51.250 62.795 ;
        RECT 51.460 68.655 51.690 68.715 ;
        RECT 53.355 68.670 53.945 68.965 ;
        RECT 51.950 68.655 53.945 68.670 ;
        RECT 51.460 66.885 53.945 68.655 ;
        RECT 51.460 65.275 52.365 66.885 ;
        RECT 53.355 66.860 53.945 66.885 ;
        RECT 55.175 68.870 55.765 68.965 ;
        RECT 56.995 68.870 57.585 68.965 ;
        RECT 55.175 67.085 57.585 68.870 ;
        RECT 58.540 68.670 59.000 69.435 ;
        RECT 59.505 68.945 59.820 69.235 ;
        RECT 59.505 68.935 59.795 68.945 ;
        RECT 61.685 68.755 62.275 68.955 ;
        RECT 59.315 68.670 59.545 68.730 ;
        RECT 58.540 67.840 59.545 68.670 ;
        RECT 55.175 66.860 55.765 67.085 ;
        RECT 56.995 66.860 57.585 67.085 ;
        RECT 53.355 66.100 53.945 66.280 ;
        RECT 55.175 66.100 55.765 66.280 ;
        RECT 51.460 62.820 52.490 65.275 ;
        RECT 53.355 64.315 55.765 66.100 ;
        RECT 56.995 65.950 57.585 66.280 ;
        RECT 53.355 64.175 53.945 64.315 ;
        RECT 55.175 64.175 55.765 64.315 ;
        RECT 56.970 64.175 57.585 65.950 ;
        RECT 56.970 62.985 57.500 64.175 ;
        RECT 51.460 62.715 51.690 62.820 ;
        RECT 51.215 62.510 51.545 62.515 ;
        RECT 51.210 62.280 51.545 62.510 ;
        RECT 51.215 62.255 51.545 62.280 ;
        RECT 51.215 62.085 51.475 62.255 ;
        RECT 50.880 61.085 51.880 62.085 ;
        RECT 46.890 60.865 47.480 60.920 ;
        RECT 48.710 60.865 49.300 60.940 ;
        RECT 51.215 60.765 51.545 61.085 ;
        RECT 51.190 60.550 51.545 60.765 ;
        RECT 51.190 60.535 51.480 60.550 ;
        RECT 51.000 60.315 51.230 60.375 ;
        RECT 46.890 60.195 47.480 60.285 ;
        RECT 46.770 57.670 47.495 60.195 ;
        RECT 48.710 60.185 49.300 60.285 ;
        RECT 48.705 58.090 49.300 60.185 ;
        RECT 50.565 59.530 51.230 60.315 ;
        RECT 50.205 58.445 51.230 59.530 ;
        RECT 48.705 57.670 49.300 57.680 ;
        RECT 50.205 57.670 50.665 58.445 ;
        RECT 51.000 58.375 51.230 58.445 ;
        RECT 51.440 60.305 51.670 60.375 ;
        RECT 52.115 60.305 52.490 62.820 ;
        RECT 53.355 62.805 53.945 62.985 ;
        RECT 55.175 62.805 55.765 62.985 ;
        RECT 53.355 61.020 55.765 62.805 ;
        RECT 53.355 60.880 53.945 61.020 ;
        RECT 55.175 60.880 55.765 61.020 ;
        RECT 56.970 61.005 57.585 62.985 ;
        RECT 58.870 62.795 59.545 67.840 ;
        RECT 59.315 62.730 59.545 62.795 ;
        RECT 59.755 68.675 59.985 68.730 ;
        RECT 60.180 68.675 62.275 68.755 ;
        RECT 59.755 66.970 62.275 68.675 ;
        RECT 59.755 65.390 60.700 66.970 ;
        RECT 61.685 66.850 62.275 66.970 ;
        RECT 63.505 68.705 64.095 68.955 ;
        RECT 65.325 68.705 65.915 68.955 ;
        RECT 63.505 66.920 65.915 68.705 ;
        RECT 66.875 68.650 67.335 69.435 ;
        RECT 67.820 68.920 68.135 69.210 ;
        RECT 67.630 68.650 67.860 68.720 ;
        RECT 66.875 67.850 67.860 68.650 ;
        RECT 63.505 66.850 64.095 66.920 ;
        RECT 65.325 66.850 65.915 66.920 ;
        RECT 61.685 66.015 62.275 66.270 ;
        RECT 63.505 66.015 64.095 66.270 ;
        RECT 59.755 62.840 60.880 65.390 ;
        RECT 61.685 64.230 64.095 66.015 ;
        RECT 65.325 65.940 65.915 66.270 ;
        RECT 61.685 64.165 62.275 64.230 ;
        RECT 63.505 64.165 64.095 64.230 ;
        RECT 59.755 62.730 59.985 62.840 ;
        RECT 59.505 62.495 59.795 62.525 ;
        RECT 59.495 62.080 59.825 62.495 ;
        RECT 59.165 61.080 60.165 62.080 ;
        RECT 56.995 60.880 57.585 61.005 ;
        RECT 59.495 60.530 59.825 61.080 ;
        RECT 51.440 58.485 52.515 60.305 ;
        RECT 51.440 58.375 51.670 58.485 ;
        RECT 51.190 57.930 51.505 58.220 ;
        RECT 53.355 58.195 53.945 60.300 ;
        RECT 55.175 60.085 55.765 60.300 ;
        RECT 55.995 60.085 56.590 60.160 ;
        RECT 56.995 60.085 57.585 60.300 ;
        RECT 59.305 60.285 59.535 60.375 ;
        RECT 59.745 60.295 59.975 60.375 ;
        RECT 60.505 60.295 60.880 62.840 ;
        RECT 61.685 62.845 62.275 62.975 ;
        RECT 63.505 62.845 64.095 62.975 ;
        RECT 61.685 61.060 64.095 62.845 ;
        RECT 61.685 60.870 62.275 61.060 ;
        RECT 63.505 60.870 64.095 61.060 ;
        RECT 65.315 60.920 65.940 65.940 ;
        RECT 67.225 62.775 67.860 67.850 ;
        RECT 67.630 62.720 67.860 62.775 ;
        RECT 68.070 68.700 68.300 68.720 ;
        RECT 68.070 68.680 68.995 68.700 ;
        RECT 69.980 68.680 70.570 68.945 ;
        RECT 68.070 66.865 70.570 68.680 ;
        RECT 68.070 65.265 68.995 66.865 ;
        RECT 69.980 66.840 70.570 66.865 ;
        RECT 71.800 68.760 72.390 68.945 ;
        RECT 73.620 68.760 74.210 68.945 ;
        RECT 71.800 66.945 74.210 68.760 ;
        RECT 75.250 68.790 75.710 69.435 ;
        RECT 76.185 69.045 76.500 69.335 ;
        RECT 76.200 69.025 76.490 69.045 ;
        RECT 76.010 68.790 76.240 68.820 ;
        RECT 75.250 68.230 76.240 68.790 ;
        RECT 71.800 66.840 72.390 66.945 ;
        RECT 73.620 66.840 74.210 66.945 ;
        RECT 69.980 66.120 70.570 66.260 ;
        RECT 71.800 66.120 72.390 66.260 ;
        RECT 68.070 62.865 69.070 65.265 ;
        RECT 69.980 64.305 72.390 66.120 ;
        RECT 69.980 64.155 70.570 64.305 ;
        RECT 71.800 64.155 72.390 64.305 ;
        RECT 73.620 65.980 74.210 66.260 ;
        RECT 68.070 62.720 68.300 62.865 ;
        RECT 67.785 62.285 68.110 62.515 ;
        RECT 67.785 61.965 68.045 62.285 ;
        RECT 67.525 60.965 68.525 61.965 ;
        RECT 65.325 60.870 65.915 60.920 ;
        RECT 67.785 60.765 68.045 60.965 ;
        RECT 67.755 60.535 68.045 60.765 ;
        RECT 55.175 58.300 57.585 60.085 ;
        RECT 58.950 59.680 59.550 60.285 ;
        RECT 55.175 58.195 55.765 58.300 ;
        RECT 56.995 58.195 57.585 58.300 ;
        RECT 58.630 58.415 59.550 59.680 ;
        RECT 59.745 58.605 60.880 60.295 ;
        RECT 59.745 58.475 60.795 58.605 ;
        RECT 58.630 57.670 59.090 58.415 ;
        RECT 59.305 58.375 59.535 58.415 ;
        RECT 59.745 58.375 59.975 58.475 ;
        RECT 59.495 57.940 59.810 58.230 ;
        RECT 61.685 58.185 62.275 60.290 ;
        RECT 63.505 60.025 64.095 60.290 ;
        RECT 64.250 60.025 64.840 60.090 ;
        RECT 65.325 60.025 65.915 60.290 ;
        RECT 67.565 60.275 67.795 60.375 ;
        RECT 63.505 58.240 65.915 60.025 ;
        RECT 67.175 59.690 67.795 60.275 ;
        RECT 63.505 58.185 64.095 58.240 ;
        RECT 65.325 58.185 65.915 58.240 ;
        RECT 66.825 58.405 67.795 59.690 ;
        RECT 61.700 58.160 62.245 58.185 ;
        RECT 66.825 57.670 67.285 58.405 ;
        RECT 67.565 58.375 67.795 58.405 ;
        RECT 68.005 60.280 68.235 60.375 ;
        RECT 68.695 60.280 69.070 62.865 ;
        RECT 69.980 62.815 70.570 62.965 ;
        RECT 71.800 62.815 72.390 62.965 ;
        RECT 69.980 61.000 72.390 62.815 ;
        RECT 69.980 60.860 70.570 61.000 ;
        RECT 71.800 60.860 72.390 61.000 ;
        RECT 73.620 60.960 74.245 65.980 ;
        RECT 75.570 62.915 76.240 68.230 ;
        RECT 76.010 62.820 76.240 62.915 ;
        RECT 76.450 68.750 76.680 68.820 ;
        RECT 76.450 68.700 77.350 68.750 ;
        RECT 78.425 68.700 79.015 68.960 ;
        RECT 76.450 66.885 79.015 68.700 ;
        RECT 76.450 65.315 77.350 66.885 ;
        RECT 78.425 66.855 79.015 66.885 ;
        RECT 80.245 68.820 80.835 68.960 ;
        RECT 82.065 68.820 82.655 68.960 ;
        RECT 80.245 67.005 82.655 68.820 ;
        RECT 83.675 68.700 84.135 69.435 ;
        RECT 84.590 68.960 84.905 69.250 ;
        RECT 84.590 68.950 84.880 68.960 ;
        RECT 86.755 68.760 87.345 68.960 ;
        RECT 84.905 68.745 87.345 68.760 ;
        RECT 84.400 68.700 84.630 68.745 ;
        RECT 83.675 68.210 84.630 68.700 ;
        RECT 80.245 66.855 80.835 67.005 ;
        RECT 82.065 66.855 82.655 67.005 ;
        RECT 78.425 66.020 79.015 66.275 ;
        RECT 80.245 66.020 80.835 66.275 ;
        RECT 82.065 66.205 82.655 66.275 ;
        RECT 76.450 62.915 77.475 65.315 ;
        RECT 78.425 64.205 80.835 66.020 ;
        RECT 78.425 64.170 79.015 64.205 ;
        RECT 80.245 64.170 80.835 64.205 ;
        RECT 76.450 62.820 76.680 62.915 ;
        RECT 76.200 62.385 76.490 62.615 ;
        RECT 76.210 62.125 76.460 62.385 ;
        RECT 75.925 61.125 76.925 62.125 ;
        RECT 73.620 60.860 74.210 60.960 ;
        RECT 76.210 60.785 76.460 61.125 ;
        RECT 76.175 60.555 76.465 60.785 ;
        RECT 75.985 60.315 76.215 60.395 ;
        RECT 68.005 58.460 69.090 60.280 ;
        RECT 69.980 60.130 70.570 60.280 ;
        RECT 68.005 58.375 68.235 58.460 ;
        RECT 67.755 58.195 68.045 58.215 ;
        RECT 67.755 57.985 68.110 58.195 ;
        RECT 69.970 58.175 70.570 60.130 ;
        RECT 71.800 60.035 72.390 60.280 ;
        RECT 73.620 60.035 74.210 60.280 ;
        RECT 71.800 58.220 74.210 60.035 ;
        RECT 75.550 59.830 76.215 60.315 ;
        RECT 75.230 59.780 76.215 59.830 ;
        RECT 71.800 58.175 72.390 58.220 ;
        RECT 73.620 58.175 74.210 58.220 ;
        RECT 75.080 58.445 76.215 59.780 ;
        RECT 69.970 58.140 70.515 58.175 ;
        RECT 67.795 57.905 68.110 57.985 ;
        RECT 75.080 57.710 75.690 58.445 ;
        RECT 75.985 58.395 76.215 58.445 ;
        RECT 76.425 60.305 76.655 60.395 ;
        RECT 77.100 60.305 77.475 62.915 ;
        RECT 78.425 62.715 79.015 62.980 ;
        RECT 80.245 62.715 80.835 62.980 ;
        RECT 78.425 60.900 80.835 62.715 ;
        RECT 78.425 60.875 79.015 60.900 ;
        RECT 80.245 60.875 80.835 60.900 ;
        RECT 82.045 60.885 82.665 66.205 ;
        RECT 84.045 62.825 84.630 68.210 ;
        RECT 84.400 62.745 84.630 62.825 ;
        RECT 84.840 66.945 87.345 68.745 ;
        RECT 84.840 65.250 85.730 66.945 ;
        RECT 86.755 66.855 87.345 66.945 ;
        RECT 88.575 68.800 89.165 68.960 ;
        RECT 90.395 68.800 90.985 68.960 ;
        RECT 88.575 66.985 90.985 68.800 ;
        RECT 92.130 68.750 92.590 69.435 ;
        RECT 92.905 68.995 93.220 69.285 ;
        RECT 92.920 68.975 93.210 68.995 ;
        RECT 92.730 68.750 92.960 68.770 ;
        RECT 92.130 67.930 92.960 68.750 ;
        RECT 88.575 66.855 89.165 66.985 ;
        RECT 90.395 66.855 90.985 66.985 ;
        RECT 86.755 66.060 87.345 66.275 ;
        RECT 88.575 66.060 89.165 66.275 ;
        RECT 84.840 62.815 85.955 65.250 ;
        RECT 86.755 64.245 89.165 66.060 ;
        RECT 90.395 65.980 90.985 66.275 ;
        RECT 86.755 64.170 87.345 64.245 ;
        RECT 88.575 64.170 89.165 64.245 ;
        RECT 84.840 62.745 85.070 62.815 ;
        RECT 84.585 62.540 84.835 62.550 ;
        RECT 84.585 62.310 84.880 62.540 ;
        RECT 84.585 62.085 84.835 62.310 ;
        RECT 84.370 61.085 85.370 62.085 ;
        RECT 82.065 60.875 82.655 60.885 ;
        RECT 84.585 60.765 84.835 61.085 ;
        RECT 84.525 60.565 84.835 60.765 ;
        RECT 84.525 60.535 84.815 60.565 ;
        RECT 76.425 58.485 77.475 60.305 ;
        RECT 84.335 60.295 84.565 60.375 ;
        RECT 76.425 58.395 76.655 58.485 ;
        RECT 76.175 58.220 76.465 58.235 ;
        RECT 76.160 57.930 76.475 58.220 ;
        RECT 78.425 58.175 79.015 60.295 ;
        RECT 80.245 60.055 80.835 60.295 ;
        RECT 82.065 60.055 82.655 60.295 ;
        RECT 80.245 58.240 82.655 60.055 ;
        RECT 83.915 59.840 84.565 60.295 ;
        RECT 80.245 58.190 80.835 58.240 ;
        RECT 82.065 58.190 82.655 58.240 ;
        RECT 83.475 58.395 84.565 59.840 ;
        RECT 74.235 57.670 75.690 57.710 ;
        RECT 83.475 57.670 83.935 58.395 ;
        RECT 84.335 58.375 84.565 58.395 ;
        RECT 84.775 60.255 85.005 60.375 ;
        RECT 85.580 60.255 85.955 62.815 ;
        RECT 86.755 62.795 87.345 62.980 ;
        RECT 88.575 62.795 89.165 62.980 ;
        RECT 86.755 60.980 89.165 62.795 ;
        RECT 86.755 60.875 87.345 60.980 ;
        RECT 88.575 60.875 89.165 60.980 ;
        RECT 90.370 60.960 90.995 65.980 ;
        RECT 92.300 62.875 92.960 67.930 ;
        RECT 92.730 62.770 92.960 62.875 ;
        RECT 93.170 68.685 93.400 68.770 ;
        RECT 93.170 68.680 94.090 68.685 ;
        RECT 95.085 68.680 95.675 68.960 ;
        RECT 93.170 66.865 95.675 68.680 ;
        RECT 93.170 65.275 94.090 66.865 ;
        RECT 95.085 66.855 95.675 66.865 ;
        RECT 96.905 68.780 97.495 68.960 ;
        RECT 98.725 68.780 99.315 68.960 ;
        RECT 96.905 66.965 99.315 68.780 ;
        RECT 100.370 68.710 100.830 69.435 ;
        RECT 101.210 68.970 101.525 69.260 ;
        RECT 101.025 68.710 101.255 68.785 ;
        RECT 100.370 67.980 101.255 68.710 ;
        RECT 96.905 66.855 97.495 66.965 ;
        RECT 98.725 66.855 99.315 66.965 ;
        RECT 95.085 66.020 95.675 66.275 ;
        RECT 96.905 66.020 97.495 66.275 ;
        RECT 98.725 66.020 99.315 66.275 ;
        RECT 93.170 62.850 94.285 65.275 ;
        RECT 95.085 64.205 97.505 66.020 ;
        RECT 95.085 64.170 95.675 64.205 ;
        RECT 96.905 64.170 97.495 64.205 ;
        RECT 93.170 62.770 93.400 62.850 ;
        RECT 92.920 62.335 93.210 62.565 ;
        RECT 92.920 62.070 93.170 62.335 ;
        RECT 92.640 61.070 93.640 62.070 ;
        RECT 90.395 60.875 90.985 60.960 ;
        RECT 92.920 60.760 93.170 61.070 ;
        RECT 92.910 60.530 93.200 60.760 ;
        RECT 92.720 60.315 92.950 60.370 ;
        RECT 84.775 58.465 85.955 60.255 ;
        RECT 86.755 60.280 87.345 60.295 ;
        RECT 84.775 58.435 85.840 58.465 ;
        RECT 84.775 58.375 85.005 58.435 ;
        RECT 86.755 58.260 87.350 60.280 ;
        RECT 88.575 60.075 89.165 60.295 ;
        RECT 90.395 60.075 90.985 60.295 ;
        RECT 88.575 58.260 90.985 60.075 ;
        RECT 92.320 59.850 92.950 60.315 ;
        RECT 84.515 57.940 84.830 58.230 ;
        RECT 86.755 58.190 87.345 58.260 ;
        RECT 88.575 58.190 89.165 58.260 ;
        RECT 89.385 58.175 89.975 58.260 ;
        RECT 90.395 58.190 90.985 58.260 ;
        RECT 91.910 58.415 92.950 59.850 ;
        RECT 91.910 57.670 92.370 58.415 ;
        RECT 92.720 58.370 92.950 58.415 ;
        RECT 93.160 60.245 93.390 60.370 ;
        RECT 93.910 60.245 94.285 62.850 ;
        RECT 95.085 62.775 95.675 62.980 ;
        RECT 96.905 62.775 97.495 62.980 ;
        RECT 95.085 60.960 97.495 62.775 ;
        RECT 98.690 61.000 99.315 66.020 ;
        RECT 100.580 62.835 101.255 67.980 ;
        RECT 101.025 62.785 101.255 62.835 ;
        RECT 101.465 68.680 101.695 68.785 ;
        RECT 103.390 68.680 103.980 68.955 ;
        RECT 101.465 66.865 103.980 68.680 ;
        RECT 101.465 65.375 102.370 66.865 ;
        RECT 103.390 66.850 103.980 66.865 ;
        RECT 105.210 68.780 105.800 68.955 ;
        RECT 107.030 68.780 107.620 68.955 ;
        RECT 105.210 66.965 107.620 68.780 ;
        RECT 108.645 68.710 109.105 69.435 ;
        RECT 109.525 69.200 109.840 69.275 ;
        RECT 109.515 68.985 109.840 69.200 ;
        RECT 109.515 68.970 109.805 68.985 ;
        RECT 111.690 68.780 112.280 68.965 ;
        RECT 113.510 68.780 114.100 68.965 ;
        RECT 109.325 68.710 109.555 68.765 ;
        RECT 108.645 67.750 109.555 68.710 ;
        RECT 105.210 66.850 105.800 66.965 ;
        RECT 107.030 66.850 107.620 66.965 ;
        RECT 103.390 66.020 103.980 66.270 ;
        RECT 105.210 66.020 105.800 66.270 ;
        RECT 101.465 62.825 102.505 65.375 ;
        RECT 103.390 64.205 105.800 66.020 ;
        RECT 103.390 64.165 103.980 64.205 ;
        RECT 105.210 64.165 105.800 64.205 ;
        RECT 107.030 66.000 107.620 66.270 ;
        RECT 107.030 64.165 107.680 66.000 ;
        RECT 107.055 62.975 107.680 64.165 ;
        RECT 101.465 62.785 101.695 62.825 ;
        RECT 101.170 62.100 101.515 62.590 ;
        RECT 100.945 61.100 101.945 62.100 ;
        RECT 95.085 60.875 95.675 60.960 ;
        RECT 96.905 60.875 97.495 60.960 ;
        RECT 98.725 60.875 99.315 61.000 ;
        RECT 101.170 60.770 101.515 61.100 ;
        RECT 101.150 60.555 101.515 60.770 ;
        RECT 101.150 60.540 101.440 60.555 ;
        RECT 100.960 60.305 101.190 60.380 ;
        RECT 93.160 58.490 94.285 60.245 ;
        RECT 95.085 60.200 95.675 60.295 ;
        RECT 93.160 58.425 94.200 58.490 ;
        RECT 93.160 58.370 93.390 58.425 ;
        RECT 92.910 58.195 93.200 58.210 ;
        RECT 92.910 57.980 93.250 58.195 ;
        RECT 95.070 58.190 95.675 60.200 ;
        RECT 96.905 60.075 97.495 60.295 ;
        RECT 98.725 60.075 99.315 60.295 ;
        RECT 96.880 58.260 99.315 60.075 ;
        RECT 100.630 59.810 101.190 60.305 ;
        RECT 96.905 58.190 97.495 58.260 ;
        RECT 98.725 58.190 99.315 58.260 ;
        RECT 100.200 58.405 101.190 59.810 ;
        RECT 95.070 58.170 95.615 58.190 ;
        RECT 92.935 57.905 93.250 57.980 ;
        RECT 100.200 57.670 100.660 58.405 ;
        RECT 100.960 58.380 101.190 58.405 ;
        RECT 101.400 60.280 101.630 60.380 ;
        RECT 102.130 60.280 102.505 62.825 ;
        RECT 103.390 62.775 103.980 62.975 ;
        RECT 105.210 62.775 105.800 62.975 ;
        RECT 103.390 60.960 105.800 62.775 ;
        RECT 103.390 60.870 103.980 60.960 ;
        RECT 105.210 60.870 105.800 60.960 ;
        RECT 107.030 60.980 107.680 62.975 ;
        RECT 108.895 62.835 109.555 67.750 ;
        RECT 109.325 62.765 109.555 62.835 ;
        RECT 109.765 68.745 109.995 68.765 ;
        RECT 109.765 66.160 110.550 68.745 ;
        RECT 111.690 66.965 114.100 68.780 ;
        RECT 111.690 66.860 112.280 66.965 ;
        RECT 113.510 66.860 114.100 66.965 ;
        RECT 127.325 66.785 128.325 66.815 ;
        RECT 111.690 66.160 112.280 66.280 ;
        RECT 109.765 64.345 112.280 66.160 ;
        RECT 113.510 66.040 114.100 66.280 ;
        RECT 126.510 66.255 128.520 66.785 ;
        RECT 109.765 63.580 110.550 64.345 ;
        RECT 111.690 64.175 112.280 64.345 ;
        RECT 113.445 64.175 114.100 66.040 ;
        RECT 126.370 65.770 128.520 66.255 ;
        RECT 126.370 64.985 126.705 65.770 ;
        RECT 127.100 65.525 127.390 65.545 ;
        RECT 127.075 65.260 127.410 65.525 ;
        RECT 126.910 64.985 127.140 65.110 ;
        RECT 126.370 64.580 127.140 64.985 ;
        RECT 109.765 62.845 110.590 63.580 ;
        RECT 109.765 62.765 109.995 62.845 ;
        RECT 109.515 62.505 109.805 62.560 ;
        RECT 109.515 62.495 110.030 62.505 ;
        RECT 109.485 62.060 110.030 62.495 ;
        RECT 110.260 62.265 110.590 62.845 ;
        RECT 111.510 62.695 112.510 63.695 ;
        RECT 113.445 62.985 114.070 64.175 ;
        RECT 126.475 64.125 127.140 64.580 ;
        RECT 126.910 64.110 127.140 64.125 ;
        RECT 127.350 64.970 127.580 65.110 ;
        RECT 127.350 64.130 128.030 64.970 ;
        RECT 127.350 64.110 127.580 64.130 ;
        RECT 127.100 63.815 127.390 63.905 ;
        RECT 127.090 63.675 127.390 63.815 ;
        RECT 127.765 63.830 128.030 64.130 ;
        RECT 128.785 64.095 129.175 73.980 ;
        RECT 128.945 64.030 129.175 64.095 ;
        RECT 129.385 73.995 129.615 74.030 ;
        RECT 129.385 66.020 129.785 73.995 ;
        RECT 130.525 73.980 130.755 74.030 ;
        RECT 129.385 65.915 129.790 66.020 ;
        RECT 129.385 65.270 129.870 65.915 ;
        RECT 129.385 65.005 129.790 65.270 ;
        RECT 129.385 64.110 129.785 65.005 ;
        RECT 129.385 64.030 129.615 64.110 ;
        RECT 130.340 64.095 130.755 73.980 ;
        RECT 130.525 64.030 130.755 64.095 ;
        RECT 130.965 74.000 131.195 74.030 ;
        RECT 130.965 64.070 131.355 74.000 ;
        RECT 132.105 73.990 132.335 74.030 ;
        RECT 131.925 65.870 132.335 73.990 ;
        RECT 131.930 65.255 132.335 65.870 ;
        RECT 131.925 64.105 132.335 65.255 ;
        RECT 130.965 64.030 131.195 64.070 ;
        RECT 132.105 64.030 132.335 64.105 ;
        RECT 132.545 74.025 132.775 74.030 ;
        RECT 132.545 66.130 132.925 74.025 ;
        RECT 133.685 73.955 133.915 74.030 ;
        RECT 132.545 65.910 132.945 66.130 ;
        RECT 132.545 65.265 132.985 65.910 ;
        RECT 133.515 65.870 133.915 73.955 ;
        RECT 132.545 65.115 132.945 65.265 ;
        RECT 133.520 65.255 133.915 65.870 ;
        RECT 132.545 64.140 132.925 65.115 ;
        RECT 132.545 64.030 132.775 64.140 ;
        RECT 133.515 64.070 133.915 65.255 ;
        RECT 133.685 64.030 133.915 64.070 ;
        RECT 134.125 73.990 134.355 74.030 ;
        RECT 134.125 64.555 134.525 73.990 ;
        RECT 134.125 64.030 134.815 64.555 ;
        RECT 127.090 63.430 127.380 63.675 ;
        RECT 127.765 63.570 134.205 63.830 ;
        RECT 127.765 63.535 131.170 63.570 ;
        RECT 132.585 63.550 134.205 63.570 ;
        RECT 132.585 63.535 133.775 63.550 ;
        RECT 109.035 61.060 110.035 62.060 ;
        RECT 110.330 61.265 110.590 62.265 ;
        RECT 107.030 60.870 107.620 60.980 ;
        RECT 109.485 60.595 110.030 61.060 ;
        RECT 110.305 60.970 110.590 61.265 ;
        RECT 111.620 61.010 112.335 62.695 ;
        RECT 113.445 61.020 114.100 62.985 ;
        RECT 126.575 62.430 127.575 63.430 ;
        RECT 127.090 62.235 127.380 62.430 ;
        RECT 127.090 62.005 127.390 62.235 ;
        RECT 126.910 61.750 127.140 61.845 ;
        RECT 126.520 61.245 127.140 61.750 ;
        RECT 109.485 60.585 109.960 60.595 ;
        RECT 109.515 60.570 109.960 60.585 ;
        RECT 109.515 60.540 109.805 60.570 ;
        RECT 109.325 60.335 109.555 60.380 ;
        RECT 101.400 58.590 102.505 60.280 ;
        RECT 103.390 60.180 103.980 60.290 ;
        RECT 101.400 58.460 102.465 58.590 ;
        RECT 101.400 58.380 101.630 58.460 ;
        RECT 101.210 58.220 101.525 58.230 ;
        RECT 101.150 57.990 101.525 58.220 ;
        RECT 103.375 58.185 103.980 60.180 ;
        RECT 105.210 60.135 105.800 60.290 ;
        RECT 107.030 60.135 107.620 60.290 ;
        RECT 105.210 58.320 107.620 60.135 ;
        RECT 108.975 59.900 109.555 60.335 ;
        RECT 105.210 58.185 105.800 58.320 ;
        RECT 103.375 58.160 103.920 58.185 ;
        RECT 106.145 58.170 106.690 58.320 ;
        RECT 107.030 58.185 107.620 58.320 ;
        RECT 108.555 58.435 109.555 59.900 ;
        RECT 101.210 57.940 101.525 57.990 ;
        RECT 108.555 57.670 109.015 58.435 ;
        RECT 109.325 58.380 109.555 58.435 ;
        RECT 109.765 60.320 109.995 60.380 ;
        RECT 110.260 60.320 110.590 60.970 ;
        RECT 111.690 60.975 112.295 61.010 ;
        RECT 111.690 60.880 112.280 60.975 ;
        RECT 113.510 60.880 114.100 61.020 ;
        RECT 126.435 60.895 127.140 61.245 ;
        RECT 109.765 58.825 110.590 60.320 ;
        RECT 111.690 60.115 112.280 60.300 ;
        RECT 113.510 60.115 114.100 60.300 ;
        RECT 109.765 58.440 110.365 58.825 ;
        RECT 109.765 58.380 109.995 58.440 ;
        RECT 111.690 58.300 114.100 60.115 ;
        RECT 126.435 60.075 126.735 60.895 ;
        RECT 126.910 60.845 127.140 60.895 ;
        RECT 127.350 61.735 127.580 61.845 ;
        RECT 127.765 61.735 128.030 63.535 ;
        RECT 134.345 63.410 134.815 64.030 ;
        RECT 131.345 63.385 132.345 63.405 ;
        RECT 128.180 62.705 128.640 63.110 ;
        RECT 128.220 62.275 128.495 62.705 ;
        RECT 131.345 62.405 133.095 63.385 ;
        RECT 133.995 62.410 134.995 63.410 ;
        RECT 128.220 62.265 129.310 62.275 ;
        RECT 128.220 62.015 134.190 62.265 ;
        RECT 128.370 61.995 134.190 62.015 ;
        RECT 129.140 61.990 134.190 61.995 ;
        RECT 134.345 61.850 134.815 62.410 ;
        RECT 128.945 61.740 129.175 61.850 ;
        RECT 127.350 60.895 128.030 61.735 ;
        RECT 127.350 60.845 127.580 60.895 ;
        RECT 127.100 60.670 127.390 60.685 ;
        RECT 127.025 60.455 127.390 60.670 ;
        RECT 127.025 60.405 127.360 60.455 ;
        RECT 127.390 60.075 128.390 60.130 ;
        RECT 126.435 59.385 128.390 60.075 ;
        RECT 126.590 59.365 128.390 59.385 ;
        RECT 127.390 59.130 128.390 59.365 ;
        RECT 109.490 57.930 109.805 58.220 ;
        RECT 111.690 58.195 112.280 58.300 ;
        RECT 113.510 58.195 114.100 58.300 ;
        RECT 128.730 57.870 129.175 61.740 ;
        RECT 128.945 57.850 129.175 57.870 ;
        RECT 129.385 61.765 129.615 61.850 ;
        RECT 129.385 57.895 129.835 61.765 ;
        RECT 130.525 61.740 130.755 61.850 ;
        RECT 129.385 57.850 129.615 57.895 ;
        RECT 130.340 57.870 130.755 61.740 ;
        RECT 130.525 57.850 130.755 57.870 ;
        RECT 130.965 61.740 131.195 61.850 ;
        RECT 132.105 61.755 132.335 61.850 ;
        RECT 130.965 57.870 131.400 61.740 ;
        RECT 131.890 57.885 132.335 61.755 ;
        RECT 130.965 57.850 131.195 57.870 ;
        RECT 132.105 57.850 132.335 57.885 ;
        RECT 132.545 61.740 132.775 61.850 ;
        RECT 132.545 57.870 132.985 61.740 ;
        RECT 133.685 61.710 133.915 61.850 ;
        RECT 132.545 57.850 132.775 57.870 ;
        RECT 133.435 57.850 133.915 61.710 ;
        RECT 134.125 60.935 134.815 61.850 ;
        RECT 134.125 57.870 134.585 60.935 ;
        RECT 134.125 57.850 134.355 57.870 ;
        RECT 133.435 57.840 133.805 57.850 ;
        RECT 10.970 57.310 13.930 57.410 ;
        RECT 2.150 57.280 4.255 57.310 ;
        RECT 2.090 56.720 4.255 57.280 ;
        RECT 4.835 57.280 6.940 57.310 ;
        RECT 8.130 57.280 10.235 57.310 ;
        RECT 4.835 56.720 10.235 57.280 ;
        RECT 10.815 56.720 13.930 57.310 ;
        RECT 46.190 57.190 114.805 57.670 ;
        RECT 129.135 57.640 129.425 57.690 ;
        RECT 130.715 57.640 131.005 57.690 ;
        RECT 132.295 57.640 132.585 57.690 ;
        RECT 133.875 57.655 134.165 57.690 ;
        RECT 129.110 57.375 129.445 57.640 ;
        RECT 130.685 57.375 131.020 57.640 ;
        RECT 132.260 57.375 132.595 57.640 ;
        RECT 133.835 57.390 134.170 57.655 ;
        RECT 2.090 55.490 3.990 56.720 ;
        RECT 4.890 56.680 10.190 56.720 ;
        RECT 10.970 56.630 13.930 56.720 ;
        RECT 46.180 56.610 114.810 57.190 ;
        RECT 2.090 54.900 4.255 55.490 ;
        RECT 4.835 55.480 6.940 55.490 ;
        RECT 8.130 55.480 10.235 55.490 ;
        RECT 4.835 54.900 10.235 55.480 ;
        RECT 10.815 54.900 12.920 55.490 ;
        RECT 2.090 54.880 3.990 54.900 ;
        RECT 4.890 54.880 10.190 54.900 ;
        RECT 2.290 53.670 4.190 53.680 ;
        RECT 4.890 53.670 10.190 53.680 ;
        RECT 10.890 53.670 12.790 54.900 ;
        RECT 2.150 53.080 4.255 53.670 ;
        RECT 4.835 53.080 10.235 53.670 ;
        RECT 10.815 53.080 12.920 53.670 ;
        RECT 2.290 51.850 4.190 53.080 ;
        RECT 61.420 52.540 61.630 52.570 ;
        RECT 61.420 52.090 67.670 52.540 ;
        RECT 61.420 52.060 61.630 52.090 ;
        RECT 10.890 51.875 13.215 51.880 ;
        RECT 10.890 51.850 16.180 51.875 ;
        RECT 25.745 51.850 26.120 51.945 ;
        RECT 41.065 51.875 46.190 51.880 ;
        RECT 28.820 51.850 46.190 51.875 ;
        RECT 46.890 51.850 52.190 51.980 ;
        RECT 52.890 51.850 58.190 51.880 ;
        RECT 58.890 51.850 70.290 51.880 ;
        RECT 70.890 51.850 76.190 51.880 ;
        RECT 76.890 51.850 82.190 51.880 ;
        RECT 2.150 51.260 4.255 51.850 ;
        RECT 4.835 51.780 6.940 51.850 ;
        RECT 8.130 51.780 10.235 51.850 ;
        RECT 4.835 51.260 10.235 51.780 ;
        RECT 10.815 51.260 16.215 51.850 ;
        RECT 16.795 51.260 22.195 51.850 ;
        RECT 22.775 51.810 24.880 51.850 ;
        RECT 25.745 51.810 28.175 51.850 ;
        RECT 22.775 51.260 28.175 51.810 ;
        RECT 28.755 51.270 46.275 51.850 ;
        RECT 28.755 51.260 30.860 51.270 ;
        RECT 41.065 51.260 46.275 51.270 ;
        RECT 46.855 51.280 52.255 51.850 ;
        RECT 46.855 51.260 48.960 51.280 ;
        RECT 50.150 51.260 52.255 51.280 ;
        RECT 52.835 51.260 58.235 51.850 ;
        RECT 58.815 51.260 70.290 51.850 ;
        RECT 70.855 51.260 76.255 51.850 ;
        RECT 76.835 51.280 82.235 51.850 ;
        RECT 76.835 51.260 78.940 51.280 ;
        RECT 80.130 51.260 82.235 51.280 ;
        RECT 82.815 51.260 84.920 51.850 ;
        RECT 4.890 51.180 10.190 51.260 ;
        RECT 10.890 51.180 16.180 51.260 ;
        RECT 16.840 51.255 22.160 51.260 ;
        RECT 12.720 51.170 16.180 51.180 ;
        RECT 1.560 50.360 9.985 50.855 ;
        RECT 10.520 50.500 11.025 50.595 ;
        RECT 17.030 50.500 17.285 51.255 ;
        RECT 22.810 51.215 28.130 51.260 ;
        RECT 28.855 50.575 29.260 51.260 ;
        RECT 41.065 51.180 46.190 51.260 ;
        RECT 47.135 50.630 47.510 51.260 ;
        RECT 52.890 51.180 58.190 51.260 ;
        RECT 58.890 51.180 70.290 51.260 ;
        RECT 70.890 51.180 76.190 51.260 ;
        RECT 59.065 50.680 59.470 51.180 ;
        RECT 10.520 50.245 17.285 50.500 ;
        RECT 10.520 50.150 11.025 50.245 ;
        RECT 26.565 50.170 29.260 50.575 ;
        RECT 38.555 50.255 47.510 50.630 ;
        RECT 54.665 50.275 59.470 50.680 ;
        RECT 71.015 50.655 71.365 51.180 ;
        RECT 81.780 50.735 82.120 51.260 ;
        RECT 82.970 51.160 84.910 51.260 ;
        RECT 83.130 50.755 83.525 51.160 ;
        RECT 66.565 50.305 71.365 50.655 ;
        RECT 77.790 50.170 80.360 50.690 ;
        RECT 81.750 50.395 82.150 50.735 ;
        RECT 82.710 50.360 83.525 50.755 ;
        RECT 84.470 51.100 84.910 51.160 ;
        RECT 144.190 51.100 146.190 51.180 ;
        RECT 84.470 50.660 146.190 51.100 ;
        RECT 27.490 49.960 30.190 49.980 ;
        RECT 55.390 49.960 58.090 49.980 ;
        RECT 83.490 49.960 85.790 49.980 ;
        RECT 111.590 49.960 113.890 49.980 ;
        RECT 1.450 49.280 139.925 49.960 ;
        RECT 144.190 49.310 146.190 50.660 ;
        RECT 1.450 49.260 27.925 49.280 ;
        RECT 29.450 49.260 55.925 49.280 ;
        RECT 57.450 49.260 83.925 49.280 ;
        RECT 85.450 49.260 111.925 49.280 ;
        RECT 113.450 49.260 139.925 49.280 ;
        RECT 2.420 48.635 4.330 49.260 ;
        RECT 6.420 48.925 8.305 48.930 ;
        RECT 9.865 48.925 11.750 48.930 ;
        RECT 6.410 48.695 8.370 48.925 ;
        RECT 9.840 48.695 11.800 48.925 ;
        RECT 2.385 48.405 4.385 48.635 ;
        RECT 6.130 48.410 6.360 48.490 ;
        RECT 1.590 48.355 2.085 48.375 ;
        RECT 1.590 45.060 2.180 48.355 ;
        RECT 4.590 48.275 4.820 48.355 ;
        RECT 4.560 45.060 4.820 48.275 ;
        RECT 1.590 43.245 4.820 45.060 ;
        RECT 1.590 40.395 2.180 43.245 ;
        RECT 3.075 40.640 3.335 40.960 ;
        RECT 4.560 40.645 4.820 43.245 ;
        RECT 5.890 40.990 6.360 48.410 ;
        RECT 6.850 41.775 7.740 48.695 ;
        RECT 8.420 48.390 8.650 48.490 ;
        RECT 8.420 48.380 8.775 48.390 ;
        RECT 9.560 48.380 9.790 48.490 ;
        RECT 3.130 40.480 3.280 40.640 ;
        RECT 1.590 35.255 2.085 40.395 ;
        RECT 3.105 40.345 3.310 40.480 ;
        RECT 4.590 40.395 4.820 40.645 ;
        RECT 5.610 40.550 6.360 40.990 ;
        RECT 6.780 40.775 7.795 41.775 ;
        RECT 2.385 40.115 4.385 40.345 ;
        RECT 5.610 38.355 5.980 40.550 ;
        RECT 6.130 40.490 6.360 40.550 ;
        RECT 6.850 40.285 7.740 40.775 ;
        RECT 8.420 40.580 9.790 48.380 ;
        RECT 10.325 43.635 11.215 48.695 ;
        RECT 11.850 48.410 12.080 48.490 ;
        RECT 10.320 42.015 11.220 43.635 ;
        RECT 10.325 41.605 11.215 42.015 ;
        RECT 10.250 40.605 11.280 41.605 ;
        RECT 11.850 40.625 12.225 48.410 ;
        RECT 12.500 48.025 14.180 49.260 ;
        RECT 15.015 48.025 19.940 48.035 ;
        RECT 12.500 47.545 19.940 48.025 ;
        RECT 12.500 45.285 14.180 47.545 ;
        RECT 15.015 47.125 19.940 47.545 ;
        RECT 14.520 46.935 14.775 46.960 ;
        RECT 14.520 46.920 14.795 46.935 ;
        RECT 14.490 46.645 14.825 46.920 ;
        RECT 15.000 46.895 20.000 47.125 ;
        RECT 20.210 46.935 20.465 46.960 ;
        RECT 14.520 46.630 14.775 46.645 ;
        RECT 15.000 46.455 20.000 46.685 ;
        RECT 20.205 46.645 20.465 46.935 ;
        RECT 20.210 46.630 20.465 46.645 ;
        RECT 15.045 46.445 19.900 46.455 ;
        RECT 15.045 44.920 17.690 44.925 ;
        RECT 13.720 44.720 17.690 44.920 ;
        RECT 13.720 44.690 17.680 44.720 ;
        RECT 12.560 44.335 12.895 44.610 ;
        RECT 13.440 44.440 13.670 44.485 ;
        RECT 8.420 40.560 8.775 40.580 ;
        RECT 8.420 40.490 8.650 40.560 ;
        RECT 9.560 40.490 9.790 40.580 ;
        RECT 10.320 40.465 11.230 40.605 ;
        RECT 11.850 40.490 12.240 40.625 ;
        RECT 10.310 40.285 11.320 40.465 ;
        RECT 6.410 40.055 8.370 40.285 ;
        RECT 9.840 40.055 11.800 40.285 ;
        RECT 7.135 39.065 7.465 40.055 ;
        RECT 9.865 40.050 11.750 40.055 ;
        RECT 12.045 38.355 12.240 40.490 ;
        RECT 12.630 38.830 12.820 44.335 ;
        RECT 13.250 43.105 13.670 44.440 ;
        RECT 14.975 43.105 16.320 44.690 ;
        RECT 13.250 41.720 16.320 43.105 ;
        RECT 13.250 40.990 13.670 41.720 ;
        RECT 13.245 40.485 13.670 40.990 ;
        RECT 12.630 38.640 12.945 38.830 ;
        RECT 2.950 38.125 6.910 38.355 ;
        RECT 8.380 38.125 12.340 38.355 ;
        RECT 12.755 38.130 12.945 38.640 ;
        RECT 2.670 37.515 2.900 37.965 ;
        RECT 4.150 37.515 4.940 38.125 ;
        RECT 2.670 37.210 4.940 37.515 ;
        RECT 2.615 37.195 4.940 37.210 ;
        RECT 2.530 36.350 4.940 37.195 ;
        RECT 2.530 35.975 2.900 36.350 ;
        RECT 2.670 35.965 2.900 35.975 ;
        RECT 4.150 35.805 4.940 36.350 ;
        RECT 6.960 37.880 7.190 37.965 ;
        RECT 8.100 37.880 8.330 37.965 ;
        RECT 6.960 36.055 8.330 37.880 ;
        RECT 6.960 35.965 7.190 36.055 ;
        RECT 2.950 35.575 6.910 35.805 ;
        RECT 2.530 35.255 2.755 35.265 ;
        RECT 7.430 35.255 7.920 36.055 ;
        RECT 8.100 35.965 8.330 36.055 ;
        RECT 9.815 37.745 11.155 38.125 ;
        RECT 12.390 37.745 12.620 37.965 ;
        RECT 9.815 36.150 12.620 37.745 ;
        RECT 9.815 35.805 11.155 36.150 ;
        RECT 12.390 35.965 12.620 36.150 ;
        RECT 8.380 35.575 12.340 35.805 ;
        RECT 12.770 35.785 12.945 38.130 ;
        RECT 13.245 37.965 13.540 40.485 ;
        RECT 14.975 40.280 16.320 41.720 ;
        RECT 17.730 44.390 17.960 44.485 ;
        RECT 18.205 44.390 18.695 46.445 ;
        RECT 19.265 44.920 19.900 44.925 ;
        RECT 19.150 44.690 23.110 44.920 ;
        RECT 18.870 44.390 19.100 44.485 ;
        RECT 17.730 40.565 19.100 44.390 ;
        RECT 17.730 40.485 17.960 40.565 ;
        RECT 18.870 40.485 19.100 40.565 ;
        RECT 20.525 40.280 21.870 44.690 ;
        RECT 23.160 44.420 23.390 44.485 ;
        RECT 24.045 44.425 24.520 49.260 ;
        RECT 25.845 48.455 26.525 49.260 ;
        RECT 26.945 48.735 27.280 48.985 ;
        RECT 26.960 48.710 27.250 48.735 ;
        RECT 30.420 48.635 32.330 49.260 ;
        RECT 34.420 48.925 36.305 48.930 ;
        RECT 37.865 48.925 39.750 48.930 ;
        RECT 34.410 48.695 36.370 48.925 ;
        RECT 37.840 48.695 39.800 48.925 ;
        RECT 26.770 48.455 27.000 48.505 ;
        RECT 25.845 47.955 27.000 48.455 ;
        RECT 24.915 44.735 25.250 44.985 ;
        RECT 24.935 44.705 25.225 44.735 ;
        RECT 24.745 44.425 24.975 44.500 ;
        RECT 23.160 40.485 23.615 44.420 ;
        RECT 24.045 43.680 24.975 44.425 ;
        RECT 24.380 40.565 24.975 43.680 ;
        RECT 24.745 40.500 24.975 40.565 ;
        RECT 25.185 44.475 25.415 44.500 ;
        RECT 25.185 40.920 25.695 44.475 ;
        RECT 25.185 40.550 25.880 40.920 ;
        RECT 26.380 40.600 27.000 47.955 ;
        RECT 25.185 40.500 25.415 40.550 ;
        RECT 13.720 40.250 17.680 40.280 ;
        RECT 19.150 40.250 23.110 40.280 ;
        RECT 13.720 40.090 23.110 40.250 ;
        RECT 13.720 40.050 17.680 40.090 ;
        RECT 19.150 40.050 23.110 40.090 ;
        RECT 23.275 38.660 23.615 40.485 ;
        RECT 24.925 38.660 25.345 40.305 ;
        RECT 23.275 38.505 25.345 38.660 ;
        RECT 23.350 38.390 25.345 38.505 ;
        RECT 13.810 38.125 17.770 38.355 ;
        RECT 19.240 38.125 23.200 38.355 ;
        RECT 13.245 37.205 13.760 37.965 ;
        RECT 13.315 36.025 13.760 37.205 ;
        RECT 13.530 35.965 13.760 36.025 ;
        RECT 15.190 35.805 16.145 38.125 ;
        RECT 17.820 37.900 18.050 37.965 ;
        RECT 18.960 37.900 19.190 37.965 ;
        RECT 17.820 36.030 19.190 37.900 ;
        RECT 17.820 35.965 18.050 36.030 ;
        RECT 12.755 35.255 12.945 35.785 ;
        RECT 13.810 35.575 17.770 35.805 ;
        RECT 18.225 35.255 18.780 36.030 ;
        RECT 18.960 35.965 19.190 36.030 ;
        RECT 20.635 35.805 21.590 38.125 ;
        RECT 23.350 37.970 23.615 38.390 ;
        RECT 24.925 38.115 25.345 38.390 ;
        RECT 25.580 39.355 25.880 40.550 ;
        RECT 26.770 40.505 27.000 40.600 ;
        RECT 27.210 48.430 27.440 48.505 ;
        RECT 27.210 41.110 27.985 48.430 ;
        RECT 30.385 48.405 32.385 48.635 ;
        RECT 34.130 48.410 34.360 48.490 ;
        RECT 29.950 45.060 30.180 48.355 ;
        RECT 32.590 48.275 32.820 48.355 ;
        RECT 32.560 45.060 32.820 48.275 ;
        RECT 29.950 43.245 32.820 45.060 ;
        RECT 27.210 40.580 28.060 41.110 ;
        RECT 29.950 40.825 30.180 43.245 ;
        RECT 27.210 40.505 27.440 40.580 ;
        RECT 26.875 39.825 27.390 40.315 ;
        RECT 27.690 39.825 28.060 40.580 ;
        RECT 29.590 40.395 30.180 40.825 ;
        RECT 31.075 40.640 31.335 40.960 ;
        RECT 32.560 40.645 32.820 43.245 ;
        RECT 33.890 40.990 34.360 48.410 ;
        RECT 34.850 41.775 35.740 48.695 ;
        RECT 36.420 48.390 36.650 48.490 ;
        RECT 36.420 48.380 36.775 48.390 ;
        RECT 37.560 48.380 37.790 48.490 ;
        RECT 31.130 40.480 31.280 40.640 ;
        RECT 26.875 39.360 27.385 39.825 ;
        RECT 26.510 39.355 27.385 39.360 ;
        RECT 25.580 38.950 27.385 39.355 ;
        RECT 25.580 38.110 25.880 38.950 ;
        RECT 26.510 38.935 27.385 38.950 ;
        RECT 26.875 38.825 27.385 38.935 ;
        RECT 26.875 38.125 27.390 38.825 ;
        RECT 27.615 38.795 28.615 39.825 ;
        RECT 23.275 37.965 23.615 37.970 ;
        RECT 23.250 36.020 23.615 37.965 ;
        RECT 24.830 37.900 25.060 37.970 ;
        RECT 24.335 37.230 25.060 37.900 ;
        RECT 24.325 37.040 25.060 37.230 ;
        RECT 24.325 36.240 24.680 37.040 ;
        RECT 24.830 36.970 25.060 37.040 ;
        RECT 25.270 37.925 25.500 37.970 ;
        RECT 25.640 37.925 25.880 38.110 ;
        RECT 25.270 37.595 25.880 37.925 ;
        RECT 26.855 37.870 27.085 37.975 ;
        RECT 25.270 37.040 25.765 37.595 ;
        RECT 25.270 36.970 25.500 37.040 ;
        RECT 25.020 36.785 25.310 36.810 ;
        RECT 25.005 36.535 25.340 36.785 ;
        RECT 26.625 36.765 27.085 37.870 ;
        RECT 26.305 36.240 27.085 36.765 ;
        RECT 23.885 36.060 27.085 36.240 ;
        RECT 23.250 35.965 23.480 36.020 ;
        RECT 19.240 35.575 23.200 35.805 ;
        RECT 23.885 35.620 26.690 36.060 ;
        RECT 26.855 35.975 27.085 36.060 ;
        RECT 27.295 37.910 27.525 37.975 ;
        RECT 27.690 37.910 28.060 38.795 ;
        RECT 27.295 37.585 28.060 37.910 ;
        RECT 27.295 36.045 28.055 37.585 ;
        RECT 27.295 35.975 27.525 36.045 ;
        RECT 27.045 35.795 27.335 35.815 ;
        RECT 23.885 35.255 26.350 35.620 ;
        RECT 27.020 35.545 27.355 35.795 ;
        RECT 29.590 35.280 30.085 40.395 ;
        RECT 31.105 40.345 31.310 40.480 ;
        RECT 32.590 40.395 32.820 40.645 ;
        RECT 33.610 40.550 34.360 40.990 ;
        RECT 34.780 40.775 35.795 41.775 ;
        RECT 30.385 40.115 32.385 40.345 ;
        RECT 33.610 38.355 33.980 40.550 ;
        RECT 34.130 40.490 34.360 40.550 ;
        RECT 34.850 40.285 35.740 40.775 ;
        RECT 36.420 40.580 37.790 48.380 ;
        RECT 38.325 43.635 39.215 48.695 ;
        RECT 39.850 48.410 40.080 48.490 ;
        RECT 38.320 42.015 39.220 43.635 ;
        RECT 38.325 41.605 39.215 42.015 ;
        RECT 38.250 40.605 39.280 41.605 ;
        RECT 39.850 40.625 40.225 48.410 ;
        RECT 40.500 48.025 42.180 49.260 ;
        RECT 43.015 48.025 47.940 48.035 ;
        RECT 40.500 47.545 47.940 48.025 ;
        RECT 40.500 45.285 42.180 47.545 ;
        RECT 43.015 47.125 47.940 47.545 ;
        RECT 42.520 46.935 42.775 46.960 ;
        RECT 42.520 46.920 42.795 46.935 ;
        RECT 42.490 46.645 42.825 46.920 ;
        RECT 43.000 46.895 48.000 47.125 ;
        RECT 48.210 46.935 48.465 46.960 ;
        RECT 42.520 46.630 42.775 46.645 ;
        RECT 43.000 46.455 48.000 46.685 ;
        RECT 48.205 46.645 48.465 46.935 ;
        RECT 48.210 46.630 48.465 46.645 ;
        RECT 43.045 46.445 47.900 46.455 ;
        RECT 43.045 44.920 45.690 44.925 ;
        RECT 41.720 44.720 45.690 44.920 ;
        RECT 41.720 44.690 45.680 44.720 ;
        RECT 40.560 44.335 40.895 44.610 ;
        RECT 41.440 44.440 41.670 44.485 ;
        RECT 36.420 40.560 36.775 40.580 ;
        RECT 36.420 40.490 36.650 40.560 ;
        RECT 37.560 40.490 37.790 40.580 ;
        RECT 38.320 40.465 39.230 40.605 ;
        RECT 39.850 40.490 40.240 40.625 ;
        RECT 38.310 40.285 39.320 40.465 ;
        RECT 34.410 40.055 36.370 40.285 ;
        RECT 37.840 40.055 39.800 40.285 ;
        RECT 35.120 39.340 35.470 40.055 ;
        RECT 37.865 40.050 39.750 40.055 ;
        RECT 40.045 38.355 40.240 40.490 ;
        RECT 40.630 38.830 40.820 44.335 ;
        RECT 41.250 43.105 41.670 44.440 ;
        RECT 42.975 43.105 44.320 44.690 ;
        RECT 41.250 41.720 44.320 43.105 ;
        RECT 41.250 40.990 41.670 41.720 ;
        RECT 41.245 40.485 41.670 40.990 ;
        RECT 40.630 38.640 40.945 38.830 ;
        RECT 30.950 38.125 34.910 38.355 ;
        RECT 36.380 38.125 40.340 38.355 ;
        RECT 40.755 38.130 40.945 38.640 ;
        RECT 30.670 37.515 30.900 37.965 ;
        RECT 32.150 37.515 32.940 38.125 ;
        RECT 30.670 37.210 32.940 37.515 ;
        RECT 30.615 37.195 32.940 37.210 ;
        RECT 30.530 36.350 32.940 37.195 ;
        RECT 30.530 35.975 30.900 36.350 ;
        RECT 30.670 35.965 30.900 35.975 ;
        RECT 32.150 35.805 32.940 36.350 ;
        RECT 34.960 37.880 35.190 37.965 ;
        RECT 36.100 37.880 36.330 37.965 ;
        RECT 34.960 36.055 36.330 37.880 ;
        RECT 34.960 35.965 35.190 36.055 ;
        RECT 30.950 35.575 34.910 35.805 ;
        RECT 27.990 35.255 30.085 35.280 ;
        RECT 30.530 35.255 30.755 35.265 ;
        RECT 35.430 35.255 35.920 36.055 ;
        RECT 36.100 35.965 36.330 36.055 ;
        RECT 37.815 37.745 39.155 38.125 ;
        RECT 40.390 37.745 40.620 37.965 ;
        RECT 37.815 36.150 40.620 37.745 ;
        RECT 37.815 35.805 39.155 36.150 ;
        RECT 40.390 35.965 40.620 36.150 ;
        RECT 36.380 35.575 40.340 35.805 ;
        RECT 40.770 35.785 40.945 38.130 ;
        RECT 41.245 37.965 41.540 40.485 ;
        RECT 42.975 40.280 44.320 41.720 ;
        RECT 45.730 44.390 45.960 44.485 ;
        RECT 46.205 44.390 46.695 46.445 ;
        RECT 47.265 44.920 47.900 44.925 ;
        RECT 47.150 44.690 51.110 44.920 ;
        RECT 46.870 44.390 47.100 44.485 ;
        RECT 45.730 40.565 47.100 44.390 ;
        RECT 45.730 40.485 45.960 40.565 ;
        RECT 46.870 40.485 47.100 40.565 ;
        RECT 48.525 40.280 49.870 44.690 ;
        RECT 51.160 44.420 51.390 44.485 ;
        RECT 52.045 44.425 52.520 49.260 ;
        RECT 53.845 48.455 54.525 49.260 ;
        RECT 54.945 48.735 55.280 48.985 ;
        RECT 54.960 48.710 55.250 48.735 ;
        RECT 58.420 48.635 60.330 49.260 ;
        RECT 62.420 48.925 64.305 48.930 ;
        RECT 65.865 48.925 67.750 48.930 ;
        RECT 62.410 48.695 64.370 48.925 ;
        RECT 65.840 48.695 67.800 48.925 ;
        RECT 54.770 48.455 55.000 48.505 ;
        RECT 53.845 47.955 55.000 48.455 ;
        RECT 52.915 44.735 53.250 44.985 ;
        RECT 52.935 44.705 53.225 44.735 ;
        RECT 52.745 44.425 52.975 44.500 ;
        RECT 51.160 40.485 51.615 44.420 ;
        RECT 52.045 43.680 52.975 44.425 ;
        RECT 52.380 40.565 52.975 43.680 ;
        RECT 52.745 40.500 52.975 40.565 ;
        RECT 53.185 44.475 53.415 44.500 ;
        RECT 53.185 40.920 53.695 44.475 ;
        RECT 53.185 40.550 53.880 40.920 ;
        RECT 54.380 40.600 55.000 47.955 ;
        RECT 53.185 40.500 53.415 40.550 ;
        RECT 41.720 40.250 45.680 40.280 ;
        RECT 47.150 40.250 51.110 40.280 ;
        RECT 41.720 40.090 51.110 40.250 ;
        RECT 41.720 40.050 45.680 40.090 ;
        RECT 47.150 40.050 51.110 40.090 ;
        RECT 51.275 38.660 51.615 40.485 ;
        RECT 52.925 38.660 53.345 40.305 ;
        RECT 51.275 38.505 53.345 38.660 ;
        RECT 51.350 38.390 53.345 38.505 ;
        RECT 41.810 38.125 45.770 38.355 ;
        RECT 47.240 38.125 51.200 38.355 ;
        RECT 41.245 37.205 41.760 37.965 ;
        RECT 41.315 36.025 41.760 37.205 ;
        RECT 41.530 35.965 41.760 36.025 ;
        RECT 43.190 35.805 44.145 38.125 ;
        RECT 45.820 37.900 46.050 37.965 ;
        RECT 46.960 37.900 47.190 37.965 ;
        RECT 45.820 36.030 47.190 37.900 ;
        RECT 45.820 35.965 46.050 36.030 ;
        RECT 40.755 35.255 40.945 35.785 ;
        RECT 41.810 35.575 45.770 35.805 ;
        RECT 46.225 35.255 46.780 36.030 ;
        RECT 46.960 35.965 47.190 36.030 ;
        RECT 48.635 35.805 49.590 38.125 ;
        RECT 51.350 37.970 51.615 38.390 ;
        RECT 52.925 38.115 53.345 38.390 ;
        RECT 53.580 39.355 53.880 40.550 ;
        RECT 54.770 40.505 55.000 40.600 ;
        RECT 55.210 48.430 55.440 48.505 ;
        RECT 55.210 41.110 55.985 48.430 ;
        RECT 58.385 48.405 60.385 48.635 ;
        RECT 62.130 48.410 62.360 48.490 ;
        RECT 57.950 45.060 58.180 48.355 ;
        RECT 60.590 48.275 60.820 48.355 ;
        RECT 60.560 45.060 60.820 48.275 ;
        RECT 57.950 43.245 60.820 45.060 ;
        RECT 55.210 40.580 56.060 41.110 ;
        RECT 57.950 40.825 58.180 43.245 ;
        RECT 55.210 40.505 55.440 40.580 ;
        RECT 54.875 39.825 55.390 40.315 ;
        RECT 54.875 39.360 55.385 39.825 ;
        RECT 55.690 39.795 56.060 40.580 ;
        RECT 57.590 40.395 58.180 40.825 ;
        RECT 59.075 40.640 59.335 40.960 ;
        RECT 60.560 40.645 60.820 43.245 ;
        RECT 61.890 40.990 62.360 48.410 ;
        RECT 62.850 41.775 63.740 48.695 ;
        RECT 64.420 48.390 64.650 48.490 ;
        RECT 64.420 48.380 64.775 48.390 ;
        RECT 65.560 48.380 65.790 48.490 ;
        RECT 59.130 40.480 59.280 40.640 ;
        RECT 54.510 39.355 55.385 39.360 ;
        RECT 53.580 38.950 55.385 39.355 ;
        RECT 53.580 38.110 53.880 38.950 ;
        RECT 54.510 38.935 55.385 38.950 ;
        RECT 54.875 38.825 55.385 38.935 ;
        RECT 54.875 38.125 55.390 38.825 ;
        RECT 55.585 38.795 56.615 39.795 ;
        RECT 51.275 37.965 51.615 37.970 ;
        RECT 51.250 36.020 51.615 37.965 ;
        RECT 52.830 37.900 53.060 37.970 ;
        RECT 52.335 37.230 53.060 37.900 ;
        RECT 52.325 37.040 53.060 37.230 ;
        RECT 52.325 36.240 52.680 37.040 ;
        RECT 52.830 36.970 53.060 37.040 ;
        RECT 53.270 37.925 53.500 37.970 ;
        RECT 53.640 37.925 53.880 38.110 ;
        RECT 53.270 37.595 53.880 37.925 ;
        RECT 54.855 37.870 55.085 37.975 ;
        RECT 53.270 37.040 53.765 37.595 ;
        RECT 53.270 36.970 53.500 37.040 ;
        RECT 53.020 36.785 53.310 36.810 ;
        RECT 53.005 36.535 53.340 36.785 ;
        RECT 54.625 36.765 55.085 37.870 ;
        RECT 54.305 36.240 55.085 36.765 ;
        RECT 51.885 36.060 55.085 36.240 ;
        RECT 51.250 35.965 51.480 36.020 ;
        RECT 47.240 35.575 51.200 35.805 ;
        RECT 51.885 35.620 54.690 36.060 ;
        RECT 54.855 35.975 55.085 36.060 ;
        RECT 55.295 37.910 55.525 37.975 ;
        RECT 55.690 37.910 56.060 38.795 ;
        RECT 55.295 37.585 56.060 37.910 ;
        RECT 55.295 36.045 56.055 37.585 ;
        RECT 55.295 35.975 55.525 36.045 ;
        RECT 55.045 35.795 55.335 35.815 ;
        RECT 51.885 35.255 54.350 35.620 ;
        RECT 55.020 35.545 55.355 35.795 ;
        RECT 57.590 35.280 58.085 40.395 ;
        RECT 59.105 40.345 59.310 40.480 ;
        RECT 60.590 40.395 60.820 40.645 ;
        RECT 61.610 40.550 62.360 40.990 ;
        RECT 62.780 40.775 63.795 41.775 ;
        RECT 58.385 40.115 60.385 40.345 ;
        RECT 61.610 38.355 61.980 40.550 ;
        RECT 62.130 40.490 62.360 40.550 ;
        RECT 62.850 40.285 63.740 40.775 ;
        RECT 64.420 40.580 65.790 48.380 ;
        RECT 66.325 43.635 67.215 48.695 ;
        RECT 67.850 48.410 68.080 48.490 ;
        RECT 66.320 42.015 67.220 43.635 ;
        RECT 66.325 41.605 67.215 42.015 ;
        RECT 66.250 40.605 67.280 41.605 ;
        RECT 67.850 40.625 68.225 48.410 ;
        RECT 68.500 48.025 70.180 49.260 ;
        RECT 71.015 48.025 75.940 48.035 ;
        RECT 68.500 47.545 75.940 48.025 ;
        RECT 68.500 45.285 70.180 47.545 ;
        RECT 71.015 47.125 75.940 47.545 ;
        RECT 70.520 46.935 70.775 46.960 ;
        RECT 70.520 46.920 70.795 46.935 ;
        RECT 70.490 46.645 70.825 46.920 ;
        RECT 71.000 46.895 76.000 47.125 ;
        RECT 76.210 46.935 76.465 46.960 ;
        RECT 70.520 46.630 70.775 46.645 ;
        RECT 71.000 46.455 76.000 46.685 ;
        RECT 76.205 46.645 76.465 46.935 ;
        RECT 76.210 46.630 76.465 46.645 ;
        RECT 71.045 46.445 75.900 46.455 ;
        RECT 71.045 44.920 73.690 44.925 ;
        RECT 69.720 44.720 73.690 44.920 ;
        RECT 69.720 44.690 73.680 44.720 ;
        RECT 68.560 44.335 68.895 44.610 ;
        RECT 69.440 44.440 69.670 44.485 ;
        RECT 64.420 40.560 64.775 40.580 ;
        RECT 64.420 40.490 64.650 40.560 ;
        RECT 65.560 40.490 65.790 40.580 ;
        RECT 66.320 40.465 67.230 40.605 ;
        RECT 67.850 40.490 68.240 40.625 ;
        RECT 66.310 40.285 67.320 40.465 ;
        RECT 62.410 40.055 64.370 40.285 ;
        RECT 65.840 40.055 67.800 40.285 ;
        RECT 63.115 39.230 63.460 40.055 ;
        RECT 65.865 40.050 67.750 40.055 ;
        RECT 68.045 38.355 68.240 40.490 ;
        RECT 68.630 38.830 68.820 44.335 ;
        RECT 69.250 43.105 69.670 44.440 ;
        RECT 70.975 43.105 72.320 44.690 ;
        RECT 69.250 41.720 72.320 43.105 ;
        RECT 69.250 40.990 69.670 41.720 ;
        RECT 69.245 40.485 69.670 40.990 ;
        RECT 68.630 38.640 68.945 38.830 ;
        RECT 58.950 38.125 62.910 38.355 ;
        RECT 64.380 38.125 68.340 38.355 ;
        RECT 68.755 38.130 68.945 38.640 ;
        RECT 58.670 37.515 58.900 37.965 ;
        RECT 60.150 37.515 60.940 38.125 ;
        RECT 58.670 37.210 60.940 37.515 ;
        RECT 58.615 37.195 60.940 37.210 ;
        RECT 58.530 36.350 60.940 37.195 ;
        RECT 58.530 35.975 58.900 36.350 ;
        RECT 58.670 35.965 58.900 35.975 ;
        RECT 60.150 35.805 60.940 36.350 ;
        RECT 62.960 37.880 63.190 37.965 ;
        RECT 64.100 37.880 64.330 37.965 ;
        RECT 62.960 36.055 64.330 37.880 ;
        RECT 62.960 35.965 63.190 36.055 ;
        RECT 58.950 35.575 62.910 35.805 ;
        RECT 55.590 35.255 58.085 35.280 ;
        RECT 58.530 35.255 58.755 35.265 ;
        RECT 63.430 35.255 63.920 36.055 ;
        RECT 64.100 35.965 64.330 36.055 ;
        RECT 65.815 37.745 67.155 38.125 ;
        RECT 68.390 37.745 68.620 37.965 ;
        RECT 65.815 36.150 68.620 37.745 ;
        RECT 65.815 35.805 67.155 36.150 ;
        RECT 68.390 35.965 68.620 36.150 ;
        RECT 64.380 35.575 68.340 35.805 ;
        RECT 68.770 35.785 68.945 38.130 ;
        RECT 69.245 37.965 69.540 40.485 ;
        RECT 70.975 40.280 72.320 41.720 ;
        RECT 73.730 44.390 73.960 44.485 ;
        RECT 74.205 44.390 74.695 46.445 ;
        RECT 75.265 44.920 75.900 44.925 ;
        RECT 75.150 44.690 79.110 44.920 ;
        RECT 74.870 44.390 75.100 44.485 ;
        RECT 73.730 40.565 75.100 44.390 ;
        RECT 73.730 40.485 73.960 40.565 ;
        RECT 74.870 40.485 75.100 40.565 ;
        RECT 76.525 40.280 77.870 44.690 ;
        RECT 79.160 44.420 79.390 44.485 ;
        RECT 80.045 44.425 80.520 49.260 ;
        RECT 81.845 48.455 82.525 49.260 ;
        RECT 82.945 48.735 83.280 48.985 ;
        RECT 82.960 48.710 83.250 48.735 ;
        RECT 86.420 48.635 88.330 49.260 ;
        RECT 90.420 48.925 92.305 48.930 ;
        RECT 93.865 48.925 95.750 48.930 ;
        RECT 90.410 48.695 92.370 48.925 ;
        RECT 93.840 48.695 95.800 48.925 ;
        RECT 82.770 48.455 83.000 48.505 ;
        RECT 81.845 47.955 83.000 48.455 ;
        RECT 80.915 44.735 81.250 44.985 ;
        RECT 80.935 44.705 81.225 44.735 ;
        RECT 80.745 44.425 80.975 44.500 ;
        RECT 79.160 40.485 79.615 44.420 ;
        RECT 80.045 43.680 80.975 44.425 ;
        RECT 80.380 40.565 80.975 43.680 ;
        RECT 80.745 40.500 80.975 40.565 ;
        RECT 81.185 44.475 81.415 44.500 ;
        RECT 81.185 40.920 81.695 44.475 ;
        RECT 81.185 40.550 81.880 40.920 ;
        RECT 82.380 40.600 83.000 47.955 ;
        RECT 81.185 40.500 81.415 40.550 ;
        RECT 69.720 40.250 73.680 40.280 ;
        RECT 75.150 40.250 79.110 40.280 ;
        RECT 69.720 40.090 79.110 40.250 ;
        RECT 69.720 40.050 73.680 40.090 ;
        RECT 75.150 40.050 79.110 40.090 ;
        RECT 79.275 38.660 79.615 40.485 ;
        RECT 80.925 38.660 81.345 40.305 ;
        RECT 79.275 38.505 81.345 38.660 ;
        RECT 79.350 38.390 81.345 38.505 ;
        RECT 69.810 38.125 73.770 38.355 ;
        RECT 75.240 38.125 79.200 38.355 ;
        RECT 69.245 37.205 69.760 37.965 ;
        RECT 69.315 36.025 69.760 37.205 ;
        RECT 69.530 35.965 69.760 36.025 ;
        RECT 71.190 35.805 72.145 38.125 ;
        RECT 73.820 37.900 74.050 37.965 ;
        RECT 74.960 37.900 75.190 37.965 ;
        RECT 73.820 36.030 75.190 37.900 ;
        RECT 73.820 35.965 74.050 36.030 ;
        RECT 68.755 35.255 68.945 35.785 ;
        RECT 69.810 35.575 73.770 35.805 ;
        RECT 74.225 35.255 74.780 36.030 ;
        RECT 74.960 35.965 75.190 36.030 ;
        RECT 76.635 35.805 77.590 38.125 ;
        RECT 79.350 37.970 79.615 38.390 ;
        RECT 80.925 38.115 81.345 38.390 ;
        RECT 81.580 39.355 81.880 40.550 ;
        RECT 82.770 40.505 83.000 40.600 ;
        RECT 83.210 48.430 83.440 48.505 ;
        RECT 83.210 41.110 83.985 48.430 ;
        RECT 86.385 48.405 88.385 48.635 ;
        RECT 90.130 48.410 90.360 48.490 ;
        RECT 85.950 45.060 86.180 48.355 ;
        RECT 88.590 48.275 88.820 48.355 ;
        RECT 88.560 45.060 88.820 48.275 ;
        RECT 85.950 43.245 88.820 45.060 ;
        RECT 83.210 40.580 84.060 41.110 ;
        RECT 85.950 40.825 86.180 43.245 ;
        RECT 83.210 40.505 83.440 40.580 ;
        RECT 82.875 39.825 83.390 40.315 ;
        RECT 82.875 39.360 83.385 39.825 ;
        RECT 83.690 39.795 84.060 40.580 ;
        RECT 85.590 40.395 86.180 40.825 ;
        RECT 87.075 40.640 87.335 40.960 ;
        RECT 88.560 40.645 88.820 43.245 ;
        RECT 89.890 40.990 90.360 48.410 ;
        RECT 90.850 41.775 91.740 48.695 ;
        RECT 92.420 48.390 92.650 48.490 ;
        RECT 92.420 48.380 92.775 48.390 ;
        RECT 93.560 48.380 93.790 48.490 ;
        RECT 87.130 40.480 87.280 40.640 ;
        RECT 82.510 39.355 83.385 39.360 ;
        RECT 81.580 38.950 83.385 39.355 ;
        RECT 81.580 38.110 81.880 38.950 ;
        RECT 82.510 38.935 83.385 38.950 ;
        RECT 82.875 38.825 83.385 38.935 ;
        RECT 82.875 38.125 83.390 38.825 ;
        RECT 83.585 38.795 84.615 39.795 ;
        RECT 79.275 37.965 79.615 37.970 ;
        RECT 79.250 36.020 79.615 37.965 ;
        RECT 80.830 37.900 81.060 37.970 ;
        RECT 80.335 37.230 81.060 37.900 ;
        RECT 80.325 37.040 81.060 37.230 ;
        RECT 80.325 36.240 80.680 37.040 ;
        RECT 80.830 36.970 81.060 37.040 ;
        RECT 81.270 37.925 81.500 37.970 ;
        RECT 81.640 37.925 81.880 38.110 ;
        RECT 81.270 37.595 81.880 37.925 ;
        RECT 82.855 37.870 83.085 37.975 ;
        RECT 81.270 37.040 81.765 37.595 ;
        RECT 81.270 36.970 81.500 37.040 ;
        RECT 81.020 36.785 81.310 36.810 ;
        RECT 81.005 36.535 81.340 36.785 ;
        RECT 82.625 36.765 83.085 37.870 ;
        RECT 82.305 36.240 83.085 36.765 ;
        RECT 79.885 36.060 83.085 36.240 ;
        RECT 79.250 35.965 79.480 36.020 ;
        RECT 79.885 35.960 82.690 36.060 ;
        RECT 82.855 35.975 83.085 36.060 ;
        RECT 83.295 37.910 83.525 37.975 ;
        RECT 83.690 37.910 84.060 38.795 ;
        RECT 83.295 37.585 84.060 37.910 ;
        RECT 83.295 36.045 84.055 37.585 ;
        RECT 83.295 35.975 83.525 36.045 ;
        RECT 75.240 35.575 79.200 35.805 ;
        RECT 79.830 35.785 82.690 35.960 ;
        RECT 83.045 35.795 83.335 35.815 ;
        RECT 79.870 35.620 82.690 35.785 ;
        RECT 79.870 35.255 82.350 35.620 ;
        RECT 83.020 35.545 83.355 35.795 ;
        RECT 85.590 35.280 86.085 40.395 ;
        RECT 87.105 40.345 87.310 40.480 ;
        RECT 88.590 40.395 88.820 40.645 ;
        RECT 89.610 40.550 90.360 40.990 ;
        RECT 90.780 40.775 91.795 41.775 ;
        RECT 86.385 40.115 88.385 40.345 ;
        RECT 89.610 38.355 89.980 40.550 ;
        RECT 90.130 40.490 90.360 40.550 ;
        RECT 90.850 40.285 91.740 40.775 ;
        RECT 92.420 40.580 93.790 48.380 ;
        RECT 94.325 43.635 95.215 48.695 ;
        RECT 95.850 48.410 96.080 48.490 ;
        RECT 94.320 42.015 95.220 43.635 ;
        RECT 94.325 41.605 95.215 42.015 ;
        RECT 94.250 40.605 95.280 41.605 ;
        RECT 95.850 40.625 96.225 48.410 ;
        RECT 96.500 48.025 98.180 49.260 ;
        RECT 99.015 48.025 103.940 48.035 ;
        RECT 96.500 47.545 103.940 48.025 ;
        RECT 96.500 45.285 98.180 47.545 ;
        RECT 99.015 47.125 103.940 47.545 ;
        RECT 98.520 46.935 98.775 46.960 ;
        RECT 98.520 46.920 98.795 46.935 ;
        RECT 98.490 46.645 98.825 46.920 ;
        RECT 99.000 46.895 104.000 47.125 ;
        RECT 104.210 46.935 104.465 46.960 ;
        RECT 98.520 46.630 98.775 46.645 ;
        RECT 99.000 46.455 104.000 46.685 ;
        RECT 104.205 46.645 104.465 46.935 ;
        RECT 104.210 46.630 104.465 46.645 ;
        RECT 99.045 46.445 103.900 46.455 ;
        RECT 99.045 44.920 101.690 44.925 ;
        RECT 97.720 44.720 101.690 44.920 ;
        RECT 97.720 44.690 101.680 44.720 ;
        RECT 96.560 44.335 96.895 44.610 ;
        RECT 97.440 44.440 97.670 44.485 ;
        RECT 92.420 40.560 92.775 40.580 ;
        RECT 92.420 40.490 92.650 40.560 ;
        RECT 93.560 40.490 93.790 40.580 ;
        RECT 94.320 40.465 95.230 40.605 ;
        RECT 95.850 40.490 96.240 40.625 ;
        RECT 94.310 40.285 95.320 40.465 ;
        RECT 90.410 40.055 92.370 40.285 ;
        RECT 93.840 40.055 95.800 40.285 ;
        RECT 91.095 39.170 91.495 40.055 ;
        RECT 93.865 40.050 95.750 40.055 ;
        RECT 96.045 38.355 96.240 40.490 ;
        RECT 96.630 38.830 96.820 44.335 ;
        RECT 97.250 43.105 97.670 44.440 ;
        RECT 98.975 43.105 100.320 44.690 ;
        RECT 97.250 41.720 100.320 43.105 ;
        RECT 97.250 40.990 97.670 41.720 ;
        RECT 97.245 40.485 97.670 40.990 ;
        RECT 96.630 38.640 96.945 38.830 ;
        RECT 86.950 38.125 90.910 38.355 ;
        RECT 92.380 38.125 96.340 38.355 ;
        RECT 96.755 38.130 96.945 38.640 ;
        RECT 86.670 37.515 86.900 37.965 ;
        RECT 88.150 37.515 88.940 38.125 ;
        RECT 86.670 37.210 88.940 37.515 ;
        RECT 86.615 37.195 88.940 37.210 ;
        RECT 86.530 36.350 88.940 37.195 ;
        RECT 86.530 35.975 86.900 36.350 ;
        RECT 86.670 35.965 86.900 35.975 ;
        RECT 88.150 35.805 88.940 36.350 ;
        RECT 90.960 37.880 91.190 37.965 ;
        RECT 92.100 37.880 92.330 37.965 ;
        RECT 90.960 36.055 92.330 37.880 ;
        RECT 90.960 35.965 91.190 36.055 ;
        RECT 86.950 35.575 90.910 35.805 ;
        RECT 83.590 35.255 86.085 35.280 ;
        RECT 86.530 35.255 86.755 35.265 ;
        RECT 91.430 35.255 91.920 36.055 ;
        RECT 92.100 35.965 92.330 36.055 ;
        RECT 93.815 37.745 95.155 38.125 ;
        RECT 96.390 37.745 96.620 37.965 ;
        RECT 93.815 36.150 96.620 37.745 ;
        RECT 93.815 35.805 95.155 36.150 ;
        RECT 96.390 35.965 96.620 36.150 ;
        RECT 92.380 35.575 96.340 35.805 ;
        RECT 96.770 35.785 96.945 38.130 ;
        RECT 97.245 37.965 97.540 40.485 ;
        RECT 98.975 40.280 100.320 41.720 ;
        RECT 101.730 44.390 101.960 44.485 ;
        RECT 102.205 44.390 102.695 46.445 ;
        RECT 103.265 44.920 103.900 44.925 ;
        RECT 103.150 44.690 107.110 44.920 ;
        RECT 102.870 44.390 103.100 44.485 ;
        RECT 101.730 40.565 103.100 44.390 ;
        RECT 101.730 40.485 101.960 40.565 ;
        RECT 102.870 40.485 103.100 40.565 ;
        RECT 104.525 40.280 105.870 44.690 ;
        RECT 107.160 44.420 107.390 44.485 ;
        RECT 108.045 44.425 108.520 49.260 ;
        RECT 109.845 48.455 110.525 49.260 ;
        RECT 110.945 48.735 111.280 48.985 ;
        RECT 110.960 48.710 111.250 48.735 ;
        RECT 114.420 48.635 116.330 49.260 ;
        RECT 118.420 48.925 120.305 48.930 ;
        RECT 121.865 48.925 123.750 48.930 ;
        RECT 118.410 48.695 120.370 48.925 ;
        RECT 121.840 48.695 123.800 48.925 ;
        RECT 110.770 48.455 111.000 48.505 ;
        RECT 109.845 47.955 111.000 48.455 ;
        RECT 108.915 44.735 109.250 44.985 ;
        RECT 108.935 44.705 109.225 44.735 ;
        RECT 108.745 44.425 108.975 44.500 ;
        RECT 107.160 40.485 107.615 44.420 ;
        RECT 108.045 43.680 108.975 44.425 ;
        RECT 108.380 40.565 108.975 43.680 ;
        RECT 108.745 40.500 108.975 40.565 ;
        RECT 109.185 44.475 109.415 44.500 ;
        RECT 109.185 40.920 109.695 44.475 ;
        RECT 109.185 40.550 109.880 40.920 ;
        RECT 110.380 40.600 111.000 47.955 ;
        RECT 109.185 40.500 109.415 40.550 ;
        RECT 97.720 40.250 101.680 40.280 ;
        RECT 103.150 40.250 107.110 40.280 ;
        RECT 97.720 40.090 107.110 40.250 ;
        RECT 97.720 40.050 101.680 40.090 ;
        RECT 103.150 40.050 107.110 40.090 ;
        RECT 107.275 38.660 107.615 40.485 ;
        RECT 108.925 38.660 109.345 40.305 ;
        RECT 107.275 38.505 109.345 38.660 ;
        RECT 107.350 38.390 109.345 38.505 ;
        RECT 97.810 38.125 101.770 38.355 ;
        RECT 103.240 38.125 107.200 38.355 ;
        RECT 97.245 37.205 97.760 37.965 ;
        RECT 97.315 36.025 97.760 37.205 ;
        RECT 97.530 35.965 97.760 36.025 ;
        RECT 99.190 35.805 100.145 38.125 ;
        RECT 101.820 37.900 102.050 37.965 ;
        RECT 102.960 37.900 103.190 37.965 ;
        RECT 101.820 36.030 103.190 37.900 ;
        RECT 101.820 35.965 102.050 36.030 ;
        RECT 96.755 35.255 96.945 35.785 ;
        RECT 97.810 35.575 101.770 35.805 ;
        RECT 102.225 35.255 102.780 36.030 ;
        RECT 102.960 35.965 103.190 36.030 ;
        RECT 104.635 35.805 105.590 38.125 ;
        RECT 107.350 37.970 107.615 38.390 ;
        RECT 108.925 38.115 109.345 38.390 ;
        RECT 109.580 39.355 109.880 40.550 ;
        RECT 110.770 40.505 111.000 40.600 ;
        RECT 111.210 48.430 111.440 48.505 ;
        RECT 111.210 41.110 111.985 48.430 ;
        RECT 114.385 48.405 116.385 48.635 ;
        RECT 118.130 48.410 118.360 48.490 ;
        RECT 113.950 45.060 114.180 48.355 ;
        RECT 116.590 48.275 116.820 48.355 ;
        RECT 116.560 45.060 116.820 48.275 ;
        RECT 113.950 43.245 116.820 45.060 ;
        RECT 111.210 40.580 112.060 41.110 ;
        RECT 113.950 40.825 114.180 43.245 ;
        RECT 111.210 40.505 111.440 40.580 ;
        RECT 110.875 39.825 111.390 40.315 ;
        RECT 110.875 39.360 111.385 39.825 ;
        RECT 111.690 39.795 112.060 40.580 ;
        RECT 113.590 40.395 114.180 40.825 ;
        RECT 115.075 40.640 115.335 40.960 ;
        RECT 116.560 40.645 116.820 43.245 ;
        RECT 117.890 40.990 118.360 48.410 ;
        RECT 118.850 41.775 119.740 48.695 ;
        RECT 120.420 48.390 120.650 48.490 ;
        RECT 120.420 48.380 120.775 48.390 ;
        RECT 121.560 48.380 121.790 48.490 ;
        RECT 115.130 40.480 115.280 40.640 ;
        RECT 110.510 39.355 111.385 39.360 ;
        RECT 109.580 38.950 111.385 39.355 ;
        RECT 109.580 38.110 109.880 38.950 ;
        RECT 110.510 38.935 111.385 38.950 ;
        RECT 110.875 38.825 111.385 38.935 ;
        RECT 110.875 38.125 111.390 38.825 ;
        RECT 111.585 38.795 112.615 39.795 ;
        RECT 107.275 37.965 107.615 37.970 ;
        RECT 107.250 36.020 107.615 37.965 ;
        RECT 108.830 37.900 109.060 37.970 ;
        RECT 108.335 37.230 109.060 37.900 ;
        RECT 108.325 37.040 109.060 37.230 ;
        RECT 108.325 36.240 108.680 37.040 ;
        RECT 108.830 36.970 109.060 37.040 ;
        RECT 109.270 37.925 109.500 37.970 ;
        RECT 109.640 37.925 109.880 38.110 ;
        RECT 109.270 37.595 109.880 37.925 ;
        RECT 110.855 37.870 111.085 37.975 ;
        RECT 109.270 37.040 109.765 37.595 ;
        RECT 109.270 36.970 109.500 37.040 ;
        RECT 109.020 36.785 109.310 36.810 ;
        RECT 109.005 36.535 109.340 36.785 ;
        RECT 110.625 36.765 111.085 37.870 ;
        RECT 110.305 36.240 111.085 36.765 ;
        RECT 107.885 36.060 111.085 36.240 ;
        RECT 107.250 35.965 107.480 36.020 ;
        RECT 103.240 35.575 107.200 35.805 ;
        RECT 107.885 35.620 110.690 36.060 ;
        RECT 110.855 35.975 111.085 36.060 ;
        RECT 111.295 37.910 111.525 37.975 ;
        RECT 111.690 37.910 112.060 38.795 ;
        RECT 111.295 37.585 112.060 37.910 ;
        RECT 111.295 36.045 112.055 37.585 ;
        RECT 111.295 35.975 111.525 36.045 ;
        RECT 111.045 35.795 111.335 35.815 ;
        RECT 107.885 35.255 110.350 35.620 ;
        RECT 111.020 35.545 111.355 35.795 ;
        RECT 113.590 35.280 114.085 40.395 ;
        RECT 115.105 40.345 115.310 40.480 ;
        RECT 116.590 40.395 116.820 40.645 ;
        RECT 117.610 40.550 118.360 40.990 ;
        RECT 118.780 40.775 119.795 41.775 ;
        RECT 114.385 40.115 116.385 40.345 ;
        RECT 117.610 38.355 117.980 40.550 ;
        RECT 118.130 40.490 118.360 40.550 ;
        RECT 118.850 40.285 119.740 40.775 ;
        RECT 120.420 40.580 121.790 48.380 ;
        RECT 122.325 43.635 123.215 48.695 ;
        RECT 123.850 48.410 124.080 48.490 ;
        RECT 122.320 42.015 123.220 43.635 ;
        RECT 122.325 41.605 123.215 42.015 ;
        RECT 122.250 40.605 123.280 41.605 ;
        RECT 123.850 40.625 124.225 48.410 ;
        RECT 124.500 48.025 126.180 49.260 ;
        RECT 127.015 48.025 131.940 48.035 ;
        RECT 124.500 47.545 131.940 48.025 ;
        RECT 124.500 45.285 126.180 47.545 ;
        RECT 127.015 47.125 131.940 47.545 ;
        RECT 126.520 46.935 126.775 46.960 ;
        RECT 126.520 46.920 126.795 46.935 ;
        RECT 126.490 46.645 126.825 46.920 ;
        RECT 127.000 46.895 132.000 47.125 ;
        RECT 132.210 46.935 132.465 46.960 ;
        RECT 126.520 46.630 126.775 46.645 ;
        RECT 127.000 46.455 132.000 46.685 ;
        RECT 132.205 46.645 132.465 46.935 ;
        RECT 132.210 46.630 132.465 46.645 ;
        RECT 127.045 46.445 131.900 46.455 ;
        RECT 127.045 44.920 129.690 44.925 ;
        RECT 125.720 44.720 129.690 44.920 ;
        RECT 125.720 44.690 129.680 44.720 ;
        RECT 124.560 44.335 124.895 44.610 ;
        RECT 125.440 44.440 125.670 44.485 ;
        RECT 120.420 40.560 120.775 40.580 ;
        RECT 120.420 40.490 120.650 40.560 ;
        RECT 121.560 40.490 121.790 40.580 ;
        RECT 122.320 40.465 123.230 40.605 ;
        RECT 123.850 40.490 124.240 40.625 ;
        RECT 122.310 40.285 123.320 40.465 ;
        RECT 118.410 40.055 120.370 40.285 ;
        RECT 121.840 40.055 123.800 40.285 ;
        RECT 119.145 39.135 119.430 40.055 ;
        RECT 121.865 40.050 123.750 40.055 ;
        RECT 124.045 38.355 124.240 40.490 ;
        RECT 124.630 38.830 124.820 44.335 ;
        RECT 125.250 43.105 125.670 44.440 ;
        RECT 126.975 43.105 128.320 44.690 ;
        RECT 125.250 41.720 128.320 43.105 ;
        RECT 125.250 40.990 125.670 41.720 ;
        RECT 125.245 40.485 125.670 40.990 ;
        RECT 124.630 38.640 124.945 38.830 ;
        RECT 114.950 38.125 118.910 38.355 ;
        RECT 120.380 38.125 124.340 38.355 ;
        RECT 124.755 38.130 124.945 38.640 ;
        RECT 114.670 37.515 114.900 37.965 ;
        RECT 116.150 37.515 116.940 38.125 ;
        RECT 114.670 37.210 116.940 37.515 ;
        RECT 114.615 37.195 116.940 37.210 ;
        RECT 114.530 36.350 116.940 37.195 ;
        RECT 114.530 35.975 114.900 36.350 ;
        RECT 114.670 35.965 114.900 35.975 ;
        RECT 116.150 35.805 116.940 36.350 ;
        RECT 118.960 37.880 119.190 37.965 ;
        RECT 120.100 37.880 120.330 37.965 ;
        RECT 118.960 36.055 120.330 37.880 ;
        RECT 118.960 35.965 119.190 36.055 ;
        RECT 114.950 35.575 118.910 35.805 ;
        RECT 111.490 35.255 114.190 35.280 ;
        RECT 114.530 35.255 114.755 35.265 ;
        RECT 119.430 35.255 119.920 36.055 ;
        RECT 120.100 35.965 120.330 36.055 ;
        RECT 121.815 37.745 123.155 38.125 ;
        RECT 124.390 37.745 124.620 37.965 ;
        RECT 121.815 36.150 124.620 37.745 ;
        RECT 121.815 35.805 123.155 36.150 ;
        RECT 124.390 35.965 124.620 36.150 ;
        RECT 120.380 35.575 124.340 35.805 ;
        RECT 124.770 35.785 124.945 38.130 ;
        RECT 125.245 37.965 125.540 40.485 ;
        RECT 126.975 40.280 128.320 41.720 ;
        RECT 129.730 44.390 129.960 44.485 ;
        RECT 130.205 44.390 130.695 46.445 ;
        RECT 131.265 44.920 131.900 44.925 ;
        RECT 131.150 44.690 135.110 44.920 ;
        RECT 130.870 44.390 131.100 44.485 ;
        RECT 129.730 40.565 131.100 44.390 ;
        RECT 129.730 40.485 129.960 40.565 ;
        RECT 130.870 40.485 131.100 40.565 ;
        RECT 132.525 40.280 133.870 44.690 ;
        RECT 135.160 44.420 135.390 44.485 ;
        RECT 136.045 44.425 136.520 49.260 ;
        RECT 137.845 48.455 138.525 49.260 ;
        RECT 138.945 48.735 139.280 48.985 ;
        RECT 138.960 48.710 139.250 48.735 ;
        RECT 144.150 48.720 146.255 49.310 ;
        RECT 146.835 48.720 148.940 49.310 ;
        RECT 138.770 48.455 139.000 48.505 ;
        RECT 137.845 47.955 139.000 48.455 ;
        RECT 136.915 44.735 137.250 44.985 ;
        RECT 136.935 44.705 137.225 44.735 ;
        RECT 136.745 44.425 136.975 44.500 ;
        RECT 135.160 40.485 135.615 44.420 ;
        RECT 136.045 43.680 136.975 44.425 ;
        RECT 136.380 40.565 136.975 43.680 ;
        RECT 136.745 40.500 136.975 40.565 ;
        RECT 137.185 44.475 137.415 44.500 ;
        RECT 137.185 40.920 137.695 44.475 ;
        RECT 137.185 40.550 137.880 40.920 ;
        RECT 138.380 40.600 139.000 47.955 ;
        RECT 137.185 40.500 137.415 40.550 ;
        RECT 125.720 40.250 129.680 40.280 ;
        RECT 131.150 40.250 135.110 40.280 ;
        RECT 125.720 40.090 135.110 40.250 ;
        RECT 125.720 40.050 129.680 40.090 ;
        RECT 131.150 40.050 135.110 40.090 ;
        RECT 135.275 38.660 135.615 40.485 ;
        RECT 136.925 38.660 137.345 40.305 ;
        RECT 135.275 38.505 137.345 38.660 ;
        RECT 135.350 38.390 137.345 38.505 ;
        RECT 125.810 38.125 129.770 38.355 ;
        RECT 131.240 38.125 135.200 38.355 ;
        RECT 125.245 37.205 125.760 37.965 ;
        RECT 125.315 36.025 125.760 37.205 ;
        RECT 125.530 35.965 125.760 36.025 ;
        RECT 127.190 35.805 128.145 38.125 ;
        RECT 129.820 37.900 130.050 37.965 ;
        RECT 130.960 37.900 131.190 37.965 ;
        RECT 129.820 36.030 131.190 37.900 ;
        RECT 129.820 35.965 130.050 36.030 ;
        RECT 124.755 35.255 124.945 35.785 ;
        RECT 125.810 35.575 129.770 35.805 ;
        RECT 130.225 35.255 130.780 36.030 ;
        RECT 130.960 35.965 131.190 36.030 ;
        RECT 132.635 35.805 133.590 38.125 ;
        RECT 135.350 37.970 135.615 38.390 ;
        RECT 136.925 38.115 137.345 38.390 ;
        RECT 137.580 39.355 137.880 40.550 ;
        RECT 138.770 40.505 139.000 40.600 ;
        RECT 139.210 48.430 139.440 48.505 ;
        RECT 139.210 41.110 139.985 48.430 ;
        RECT 146.860 47.490 148.890 48.720 ;
        RECT 144.150 46.900 146.255 47.490 ;
        RECT 146.835 46.900 148.940 47.490 ;
        RECT 144.160 45.670 146.190 46.900 ;
        RECT 146.890 46.880 148.890 46.900 ;
        RECT 146.890 45.670 154.890 45.680 ;
        RECT 144.150 45.080 146.255 45.670 ;
        RECT 146.835 45.180 154.890 45.670 ;
        RECT 146.835 45.080 148.940 45.180 ;
        RECT 144.190 43.850 146.190 43.880 ;
        RECT 144.150 43.260 146.255 43.850 ;
        RECT 146.835 43.780 148.940 43.850 ;
        RECT 149.425 43.780 149.925 44.125 ;
        RECT 152.890 43.850 154.890 45.180 ;
        RECT 150.130 43.780 152.235 43.850 ;
        RECT 146.835 43.280 152.235 43.780 ;
        RECT 146.835 43.260 148.940 43.280 ;
        RECT 150.130 43.260 152.235 43.280 ;
        RECT 152.815 43.260 154.920 43.850 ;
        RECT 144.190 42.945 146.190 43.260 ;
        RECT 141.790 42.505 146.190 42.945 ;
        RECT 144.190 42.030 146.190 42.505 ;
        RECT 144.150 41.440 146.255 42.030 ;
        RECT 146.835 41.980 148.940 42.030 ;
        RECT 150.130 41.980 152.235 42.030 ;
        RECT 146.835 41.480 152.235 41.980 ;
        RECT 146.835 41.440 148.940 41.480 ;
        RECT 149.530 41.440 152.235 41.480 ;
        RECT 152.815 41.440 154.920 42.030 ;
        RECT 149.530 41.240 150.310 41.440 ;
        RECT 139.210 40.580 140.060 41.110 ;
        RECT 149.530 41.035 150.030 41.240 ;
        RECT 139.210 40.505 139.440 40.580 ;
        RECT 138.875 39.825 139.390 40.315 ;
        RECT 138.875 39.360 139.385 39.825 ;
        RECT 139.690 39.795 140.060 40.580 ;
        RECT 142.350 40.535 150.030 41.035 ;
        RECT 153.565 40.995 154.355 41.440 ;
        RECT 150.785 40.205 154.355 40.995 ;
        RECT 150.785 40.055 151.575 40.205 ;
        RECT 138.510 39.355 139.385 39.360 ;
        RECT 137.580 38.950 139.385 39.355 ;
        RECT 137.580 38.110 137.880 38.950 ;
        RECT 138.510 38.935 139.385 38.950 ;
        RECT 138.875 38.825 139.385 38.935 ;
        RECT 138.875 38.125 139.390 38.825 ;
        RECT 139.585 38.795 140.615 39.795 ;
        RECT 141.105 39.265 151.575 40.055 ;
        RECT 135.275 37.965 135.615 37.970 ;
        RECT 135.250 36.020 135.615 37.965 ;
        RECT 136.830 37.900 137.060 37.970 ;
        RECT 136.335 37.230 137.060 37.900 ;
        RECT 136.325 37.040 137.060 37.230 ;
        RECT 136.325 36.240 136.680 37.040 ;
        RECT 136.830 36.970 137.060 37.040 ;
        RECT 137.270 37.925 137.500 37.970 ;
        RECT 137.640 37.925 137.880 38.110 ;
        RECT 137.270 37.595 137.880 37.925 ;
        RECT 138.855 37.870 139.085 37.975 ;
        RECT 137.270 37.040 137.765 37.595 ;
        RECT 137.270 36.970 137.500 37.040 ;
        RECT 137.020 36.785 137.310 36.810 ;
        RECT 137.005 36.535 137.340 36.785 ;
        RECT 138.625 36.765 139.085 37.870 ;
        RECT 138.305 36.240 139.085 36.765 ;
        RECT 135.885 36.060 139.085 36.240 ;
        RECT 135.250 35.965 135.480 36.020 ;
        RECT 131.240 35.575 135.200 35.805 ;
        RECT 135.885 35.620 138.690 36.060 ;
        RECT 138.855 35.975 139.085 36.060 ;
        RECT 139.295 37.910 139.525 37.975 ;
        RECT 139.690 37.910 140.060 38.795 ;
        RECT 139.295 37.585 140.060 37.910 ;
        RECT 139.295 36.045 140.055 37.585 ;
        RECT 139.295 35.975 139.525 36.045 ;
        RECT 139.045 35.795 139.335 35.815 ;
        RECT 135.885 35.335 138.350 35.620 ;
        RECT 139.020 35.545 139.355 35.795 ;
        RECT 141.105 35.335 141.895 39.265 ;
        RECT 135.885 35.255 141.895 35.335 ;
        RECT 1.475 34.545 141.895 35.255 ;
        RECT 1.475 34.380 140.080 34.545 ;
        RECT 27.790 33.960 30.490 33.980 ;
        RECT 55.390 33.960 57.990 33.980 ;
        RECT 83.390 33.960 86.290 33.980 ;
        RECT 111.190 33.960 114.190 33.980 ;
        RECT 1.450 33.280 139.925 33.960 ;
        RECT 1.450 33.260 27.925 33.280 ;
        RECT 29.450 33.260 83.925 33.280 ;
        RECT 85.450 33.260 111.925 33.280 ;
        RECT 113.450 33.260 139.925 33.280 ;
        RECT 2.420 32.635 4.330 33.260 ;
        RECT 6.420 32.925 8.305 32.930 ;
        RECT 9.865 32.925 11.750 32.930 ;
        RECT 6.410 32.695 8.370 32.925 ;
        RECT 9.840 32.695 11.800 32.925 ;
        RECT 2.385 32.405 4.385 32.635 ;
        RECT 6.130 32.410 6.360 32.490 ;
        RECT 1.950 29.060 2.180 32.355 ;
        RECT 4.590 32.275 4.820 32.355 ;
        RECT 4.560 29.060 4.820 32.275 ;
        RECT 1.950 27.245 4.820 29.060 ;
        RECT 1.950 24.825 2.180 27.245 ;
        RECT 1.590 24.395 2.180 24.825 ;
        RECT 3.075 24.640 3.335 24.960 ;
        RECT 4.560 24.645 4.820 27.245 ;
        RECT 5.890 24.990 6.360 32.410 ;
        RECT 6.850 25.775 7.740 32.695 ;
        RECT 8.420 32.390 8.650 32.490 ;
        RECT 8.420 32.380 8.775 32.390 ;
        RECT 9.560 32.380 9.790 32.490 ;
        RECT 3.130 24.480 3.280 24.640 ;
        RECT 1.590 19.255 2.085 24.395 ;
        RECT 3.105 24.345 3.310 24.480 ;
        RECT 4.590 24.395 4.820 24.645 ;
        RECT 5.610 24.550 6.360 24.990 ;
        RECT 6.780 24.775 7.795 25.775 ;
        RECT 2.385 24.115 4.385 24.345 ;
        RECT 5.610 22.355 5.980 24.550 ;
        RECT 6.130 24.490 6.360 24.550 ;
        RECT 6.850 24.285 7.740 24.775 ;
        RECT 8.420 24.580 9.790 32.380 ;
        RECT 10.325 27.635 11.215 32.695 ;
        RECT 11.850 32.410 12.080 32.490 ;
        RECT 10.320 26.015 11.220 27.635 ;
        RECT 10.325 25.605 11.215 26.015 ;
        RECT 10.250 24.605 11.280 25.605 ;
        RECT 11.850 24.625 12.225 32.410 ;
        RECT 12.500 32.025 14.180 33.260 ;
        RECT 15.015 32.025 19.940 32.035 ;
        RECT 12.500 31.545 19.940 32.025 ;
        RECT 12.500 29.285 14.180 31.545 ;
        RECT 15.015 31.125 19.940 31.545 ;
        RECT 14.520 30.935 14.775 30.960 ;
        RECT 14.520 30.920 14.795 30.935 ;
        RECT 14.490 30.645 14.825 30.920 ;
        RECT 15.000 30.895 20.000 31.125 ;
        RECT 20.210 30.935 20.465 30.960 ;
        RECT 14.520 30.630 14.775 30.645 ;
        RECT 15.000 30.455 20.000 30.685 ;
        RECT 20.205 30.645 20.465 30.935 ;
        RECT 20.210 30.630 20.465 30.645 ;
        RECT 15.045 30.445 19.900 30.455 ;
        RECT 15.045 28.920 17.690 28.925 ;
        RECT 13.720 28.720 17.690 28.920 ;
        RECT 13.720 28.690 17.680 28.720 ;
        RECT 12.560 28.335 12.895 28.610 ;
        RECT 13.440 28.440 13.670 28.485 ;
        RECT 8.420 24.560 8.775 24.580 ;
        RECT 8.420 24.490 8.650 24.560 ;
        RECT 9.560 24.490 9.790 24.580 ;
        RECT 10.320 24.465 11.230 24.605 ;
        RECT 11.850 24.490 12.240 24.625 ;
        RECT 10.310 24.285 11.320 24.465 ;
        RECT 6.410 24.055 8.370 24.285 ;
        RECT 9.840 24.055 11.800 24.285 ;
        RECT 7.165 23.035 7.495 24.055 ;
        RECT 9.865 24.050 11.750 24.055 ;
        RECT 12.045 22.355 12.240 24.490 ;
        RECT 12.630 22.830 12.820 28.335 ;
        RECT 13.250 27.105 13.670 28.440 ;
        RECT 14.975 27.105 16.320 28.690 ;
        RECT 13.250 25.720 16.320 27.105 ;
        RECT 13.250 24.990 13.670 25.720 ;
        RECT 13.245 24.485 13.670 24.990 ;
        RECT 12.630 22.640 12.945 22.830 ;
        RECT 2.950 22.125 6.910 22.355 ;
        RECT 8.380 22.125 12.340 22.355 ;
        RECT 12.755 22.130 12.945 22.640 ;
        RECT 2.670 21.515 2.900 21.965 ;
        RECT 4.150 21.515 4.940 22.125 ;
        RECT 2.670 21.210 4.940 21.515 ;
        RECT 2.615 21.195 4.940 21.210 ;
        RECT 2.530 20.350 4.940 21.195 ;
        RECT 2.530 19.975 2.900 20.350 ;
        RECT 2.670 19.965 2.900 19.975 ;
        RECT 4.150 19.805 4.940 20.350 ;
        RECT 6.960 21.880 7.190 21.965 ;
        RECT 8.100 21.880 8.330 21.965 ;
        RECT 6.960 20.055 8.330 21.880 ;
        RECT 6.960 19.965 7.190 20.055 ;
        RECT 2.950 19.575 6.910 19.805 ;
        RECT 2.530 19.255 2.755 19.265 ;
        RECT 7.430 19.255 7.920 20.055 ;
        RECT 8.100 19.965 8.330 20.055 ;
        RECT 9.815 21.745 11.155 22.125 ;
        RECT 12.390 21.745 12.620 21.965 ;
        RECT 9.815 20.150 12.620 21.745 ;
        RECT 9.815 19.805 11.155 20.150 ;
        RECT 12.390 19.965 12.620 20.150 ;
        RECT 8.380 19.575 12.340 19.805 ;
        RECT 12.770 19.785 12.945 22.130 ;
        RECT 13.245 21.965 13.540 24.485 ;
        RECT 14.975 24.280 16.320 25.720 ;
        RECT 17.730 28.390 17.960 28.485 ;
        RECT 18.205 28.390 18.695 30.445 ;
        RECT 19.265 28.920 19.900 28.925 ;
        RECT 19.150 28.690 23.110 28.920 ;
        RECT 18.870 28.390 19.100 28.485 ;
        RECT 17.730 24.565 19.100 28.390 ;
        RECT 17.730 24.485 17.960 24.565 ;
        RECT 18.870 24.485 19.100 24.565 ;
        RECT 20.525 24.280 21.870 28.690 ;
        RECT 23.160 28.420 23.390 28.485 ;
        RECT 24.045 28.425 24.520 33.260 ;
        RECT 25.845 32.455 26.525 33.260 ;
        RECT 26.945 32.735 27.280 32.985 ;
        RECT 26.960 32.710 27.250 32.735 ;
        RECT 30.420 32.635 32.330 33.260 ;
        RECT 34.420 32.925 36.305 32.930 ;
        RECT 37.865 32.925 39.750 32.930 ;
        RECT 34.410 32.695 36.370 32.925 ;
        RECT 37.840 32.695 39.800 32.925 ;
        RECT 26.770 32.455 27.000 32.505 ;
        RECT 25.845 31.955 27.000 32.455 ;
        RECT 24.915 28.735 25.250 28.985 ;
        RECT 24.935 28.705 25.225 28.735 ;
        RECT 24.745 28.425 24.975 28.500 ;
        RECT 23.160 24.485 23.615 28.420 ;
        RECT 24.045 27.680 24.975 28.425 ;
        RECT 24.380 24.565 24.975 27.680 ;
        RECT 24.745 24.500 24.975 24.565 ;
        RECT 25.185 28.475 25.415 28.500 ;
        RECT 25.185 24.920 25.695 28.475 ;
        RECT 25.185 24.550 25.880 24.920 ;
        RECT 26.380 24.600 27.000 31.955 ;
        RECT 25.185 24.500 25.415 24.550 ;
        RECT 13.720 24.250 17.680 24.280 ;
        RECT 19.150 24.250 23.110 24.280 ;
        RECT 13.720 24.090 23.110 24.250 ;
        RECT 13.720 24.050 17.680 24.090 ;
        RECT 19.150 24.050 23.110 24.090 ;
        RECT 23.275 22.660 23.615 24.485 ;
        RECT 24.925 22.660 25.345 24.305 ;
        RECT 23.275 22.505 25.345 22.660 ;
        RECT 23.350 22.390 25.345 22.505 ;
        RECT 13.810 22.125 17.770 22.355 ;
        RECT 19.240 22.125 23.200 22.355 ;
        RECT 13.245 21.205 13.760 21.965 ;
        RECT 13.315 20.025 13.760 21.205 ;
        RECT 13.530 19.965 13.760 20.025 ;
        RECT 15.190 19.805 16.145 22.125 ;
        RECT 17.820 21.900 18.050 21.965 ;
        RECT 18.960 21.900 19.190 21.965 ;
        RECT 17.820 20.030 19.190 21.900 ;
        RECT 17.820 19.965 18.050 20.030 ;
        RECT 12.755 19.255 12.945 19.785 ;
        RECT 13.810 19.575 17.770 19.805 ;
        RECT 18.225 19.255 18.780 20.030 ;
        RECT 18.960 19.965 19.190 20.030 ;
        RECT 20.635 19.805 21.590 22.125 ;
        RECT 23.350 21.970 23.615 22.390 ;
        RECT 24.925 22.115 25.345 22.390 ;
        RECT 25.580 23.355 25.880 24.550 ;
        RECT 26.770 24.505 27.000 24.600 ;
        RECT 27.210 32.430 27.440 32.505 ;
        RECT 27.210 25.110 27.985 32.430 ;
        RECT 30.385 32.405 32.385 32.635 ;
        RECT 34.130 32.410 34.360 32.490 ;
        RECT 29.950 29.060 30.180 32.355 ;
        RECT 32.590 32.275 32.820 32.355 ;
        RECT 32.560 29.060 32.820 32.275 ;
        RECT 29.950 27.245 32.820 29.060 ;
        RECT 27.210 24.580 28.060 25.110 ;
        RECT 29.950 24.825 30.180 27.245 ;
        RECT 27.210 24.505 27.440 24.580 ;
        RECT 26.875 23.825 27.390 24.315 ;
        RECT 27.690 23.825 28.060 24.580 ;
        RECT 29.590 24.395 30.180 24.825 ;
        RECT 31.075 24.640 31.335 24.960 ;
        RECT 32.560 24.645 32.820 27.245 ;
        RECT 33.890 24.990 34.360 32.410 ;
        RECT 34.850 25.775 35.740 32.695 ;
        RECT 36.420 32.390 36.650 32.490 ;
        RECT 36.420 32.380 36.775 32.390 ;
        RECT 37.560 32.380 37.790 32.490 ;
        RECT 31.130 24.480 31.280 24.640 ;
        RECT 26.875 23.360 27.385 23.825 ;
        RECT 26.510 23.355 27.385 23.360 ;
        RECT 25.580 22.950 27.385 23.355 ;
        RECT 25.580 22.110 25.880 22.950 ;
        RECT 26.510 22.935 27.385 22.950 ;
        RECT 26.875 22.825 27.385 22.935 ;
        RECT 26.875 22.125 27.390 22.825 ;
        RECT 27.615 22.795 28.615 23.825 ;
        RECT 23.275 21.965 23.615 21.970 ;
        RECT 23.250 20.020 23.615 21.965 ;
        RECT 24.830 21.900 25.060 21.970 ;
        RECT 24.335 21.230 25.060 21.900 ;
        RECT 24.325 21.040 25.060 21.230 ;
        RECT 24.325 20.240 24.680 21.040 ;
        RECT 24.830 20.970 25.060 21.040 ;
        RECT 25.270 21.925 25.500 21.970 ;
        RECT 25.640 21.925 25.880 22.110 ;
        RECT 25.270 21.595 25.880 21.925 ;
        RECT 26.855 21.870 27.085 21.975 ;
        RECT 25.270 21.040 25.765 21.595 ;
        RECT 25.270 20.970 25.500 21.040 ;
        RECT 25.020 20.785 25.310 20.810 ;
        RECT 25.005 20.535 25.340 20.785 ;
        RECT 26.625 20.765 27.085 21.870 ;
        RECT 26.305 20.240 27.085 20.765 ;
        RECT 23.885 20.060 27.085 20.240 ;
        RECT 23.250 19.965 23.480 20.020 ;
        RECT 19.240 19.575 23.200 19.805 ;
        RECT 23.885 19.620 26.690 20.060 ;
        RECT 26.855 19.975 27.085 20.060 ;
        RECT 27.295 21.910 27.525 21.975 ;
        RECT 27.690 21.910 28.060 22.795 ;
        RECT 27.295 21.585 28.060 21.910 ;
        RECT 27.295 20.045 28.055 21.585 ;
        RECT 27.295 19.975 27.525 20.045 ;
        RECT 27.045 19.795 27.335 19.815 ;
        RECT 23.885 19.255 26.350 19.620 ;
        RECT 27.020 19.545 27.355 19.795 ;
        RECT 29.590 19.280 30.085 24.395 ;
        RECT 31.105 24.345 31.310 24.480 ;
        RECT 32.590 24.395 32.820 24.645 ;
        RECT 33.610 24.550 34.360 24.990 ;
        RECT 34.780 24.775 35.795 25.775 ;
        RECT 30.385 24.115 32.385 24.345 ;
        RECT 33.610 22.355 33.980 24.550 ;
        RECT 34.130 24.490 34.360 24.550 ;
        RECT 34.850 24.285 35.740 24.775 ;
        RECT 36.420 24.580 37.790 32.380 ;
        RECT 38.325 27.635 39.215 32.695 ;
        RECT 39.850 32.410 40.080 32.490 ;
        RECT 38.320 26.015 39.220 27.635 ;
        RECT 38.325 25.605 39.215 26.015 ;
        RECT 38.250 24.605 39.280 25.605 ;
        RECT 39.850 24.625 40.225 32.410 ;
        RECT 40.500 32.025 42.180 33.260 ;
        RECT 43.015 32.025 47.940 32.035 ;
        RECT 40.500 31.545 47.940 32.025 ;
        RECT 40.500 29.285 42.180 31.545 ;
        RECT 43.015 31.125 47.940 31.545 ;
        RECT 42.520 30.935 42.775 30.960 ;
        RECT 42.520 30.920 42.795 30.935 ;
        RECT 42.490 30.645 42.825 30.920 ;
        RECT 43.000 30.895 48.000 31.125 ;
        RECT 48.210 30.935 48.465 30.960 ;
        RECT 42.520 30.630 42.775 30.645 ;
        RECT 43.000 30.455 48.000 30.685 ;
        RECT 48.205 30.645 48.465 30.935 ;
        RECT 48.210 30.630 48.465 30.645 ;
        RECT 43.045 30.445 47.900 30.455 ;
        RECT 43.045 28.920 45.690 28.925 ;
        RECT 41.720 28.720 45.690 28.920 ;
        RECT 41.720 28.690 45.680 28.720 ;
        RECT 40.560 28.335 40.895 28.610 ;
        RECT 41.440 28.440 41.670 28.485 ;
        RECT 36.420 24.560 36.775 24.580 ;
        RECT 36.420 24.490 36.650 24.560 ;
        RECT 37.560 24.490 37.790 24.580 ;
        RECT 38.320 24.465 39.230 24.605 ;
        RECT 39.850 24.490 40.240 24.625 ;
        RECT 38.310 24.285 39.320 24.465 ;
        RECT 34.410 24.055 36.370 24.285 ;
        RECT 37.840 24.055 39.800 24.285 ;
        RECT 35.115 23.005 35.465 24.055 ;
        RECT 37.865 24.050 39.750 24.055 ;
        RECT 40.045 22.355 40.240 24.490 ;
        RECT 40.630 22.830 40.820 28.335 ;
        RECT 41.250 27.105 41.670 28.440 ;
        RECT 42.975 27.105 44.320 28.690 ;
        RECT 41.250 25.720 44.320 27.105 ;
        RECT 41.250 24.990 41.670 25.720 ;
        RECT 41.245 24.485 41.670 24.990 ;
        RECT 40.630 22.640 40.945 22.830 ;
        RECT 30.950 22.125 34.910 22.355 ;
        RECT 36.380 22.125 40.340 22.355 ;
        RECT 40.755 22.130 40.945 22.640 ;
        RECT 30.670 21.515 30.900 21.965 ;
        RECT 32.150 21.515 32.940 22.125 ;
        RECT 30.670 21.210 32.940 21.515 ;
        RECT 30.615 21.195 32.940 21.210 ;
        RECT 30.530 20.350 32.940 21.195 ;
        RECT 30.530 19.975 30.900 20.350 ;
        RECT 30.670 19.965 30.900 19.975 ;
        RECT 32.150 19.805 32.940 20.350 ;
        RECT 34.960 21.880 35.190 21.965 ;
        RECT 36.100 21.880 36.330 21.965 ;
        RECT 34.960 20.055 36.330 21.880 ;
        RECT 34.960 19.965 35.190 20.055 ;
        RECT 30.950 19.575 34.910 19.805 ;
        RECT 27.890 19.255 30.085 19.280 ;
        RECT 30.530 19.255 30.755 19.265 ;
        RECT 35.430 19.255 35.920 20.055 ;
        RECT 36.100 19.965 36.330 20.055 ;
        RECT 37.815 21.745 39.155 22.125 ;
        RECT 40.390 21.745 40.620 21.965 ;
        RECT 37.815 20.150 40.620 21.745 ;
        RECT 37.815 19.805 39.155 20.150 ;
        RECT 40.390 19.965 40.620 20.150 ;
        RECT 36.380 19.575 40.340 19.805 ;
        RECT 40.770 19.785 40.945 22.130 ;
        RECT 41.245 21.965 41.540 24.485 ;
        RECT 42.975 24.280 44.320 25.720 ;
        RECT 45.730 28.390 45.960 28.485 ;
        RECT 46.205 28.390 46.695 30.445 ;
        RECT 47.265 28.920 47.900 28.925 ;
        RECT 47.150 28.690 51.110 28.920 ;
        RECT 46.870 28.390 47.100 28.485 ;
        RECT 45.730 24.565 47.100 28.390 ;
        RECT 45.730 24.485 45.960 24.565 ;
        RECT 46.870 24.485 47.100 24.565 ;
        RECT 48.525 24.280 49.870 28.690 ;
        RECT 51.160 28.420 51.390 28.485 ;
        RECT 52.045 28.425 52.520 33.260 ;
        RECT 53.845 32.455 54.525 33.260 ;
        RECT 55.390 33.180 57.990 33.260 ;
        RECT 54.945 32.735 55.280 32.985 ;
        RECT 54.960 32.710 55.250 32.735 ;
        RECT 58.420 32.635 60.330 33.260 ;
        RECT 62.420 32.925 64.305 32.930 ;
        RECT 65.865 32.925 67.750 32.930 ;
        RECT 62.410 32.695 64.370 32.925 ;
        RECT 65.840 32.695 67.800 32.925 ;
        RECT 54.770 32.455 55.000 32.505 ;
        RECT 53.845 31.955 55.000 32.455 ;
        RECT 52.915 28.735 53.250 28.985 ;
        RECT 52.935 28.705 53.225 28.735 ;
        RECT 52.745 28.425 52.975 28.500 ;
        RECT 51.160 24.485 51.615 28.420 ;
        RECT 52.045 27.680 52.975 28.425 ;
        RECT 52.380 24.565 52.975 27.680 ;
        RECT 52.745 24.500 52.975 24.565 ;
        RECT 53.185 28.475 53.415 28.500 ;
        RECT 53.185 24.920 53.695 28.475 ;
        RECT 53.185 24.550 53.880 24.920 ;
        RECT 54.380 24.600 55.000 31.955 ;
        RECT 53.185 24.500 53.415 24.550 ;
        RECT 41.720 24.250 45.680 24.280 ;
        RECT 47.150 24.250 51.110 24.280 ;
        RECT 41.720 24.090 51.110 24.250 ;
        RECT 41.720 24.050 45.680 24.090 ;
        RECT 47.150 24.050 51.110 24.090 ;
        RECT 51.275 22.660 51.615 24.485 ;
        RECT 52.925 22.660 53.345 24.305 ;
        RECT 51.275 22.505 53.345 22.660 ;
        RECT 51.350 22.390 53.345 22.505 ;
        RECT 41.810 22.125 45.770 22.355 ;
        RECT 47.240 22.125 51.200 22.355 ;
        RECT 41.245 21.205 41.760 21.965 ;
        RECT 41.315 20.025 41.760 21.205 ;
        RECT 41.530 19.965 41.760 20.025 ;
        RECT 43.190 19.805 44.145 22.125 ;
        RECT 45.820 21.900 46.050 21.965 ;
        RECT 46.960 21.900 47.190 21.965 ;
        RECT 45.820 20.030 47.190 21.900 ;
        RECT 45.820 19.965 46.050 20.030 ;
        RECT 40.755 19.255 40.945 19.785 ;
        RECT 41.810 19.575 45.770 19.805 ;
        RECT 46.225 19.255 46.780 20.030 ;
        RECT 46.960 19.965 47.190 20.030 ;
        RECT 48.635 19.805 49.590 22.125 ;
        RECT 51.350 21.970 51.615 22.390 ;
        RECT 52.925 22.115 53.345 22.390 ;
        RECT 53.580 23.355 53.880 24.550 ;
        RECT 54.770 24.505 55.000 24.600 ;
        RECT 55.210 32.430 55.440 32.505 ;
        RECT 55.210 25.110 55.985 32.430 ;
        RECT 58.385 32.405 60.385 32.635 ;
        RECT 62.130 32.410 62.360 32.490 ;
        RECT 57.950 29.060 58.180 32.355 ;
        RECT 60.590 32.275 60.820 32.355 ;
        RECT 60.560 29.060 60.820 32.275 ;
        RECT 57.950 27.245 60.820 29.060 ;
        RECT 55.210 24.580 56.060 25.110 ;
        RECT 57.950 24.825 58.180 27.245 ;
        RECT 55.210 24.505 55.440 24.580 ;
        RECT 54.875 23.825 55.390 24.315 ;
        RECT 54.875 23.360 55.385 23.825 ;
        RECT 55.690 23.795 56.060 24.580 ;
        RECT 57.590 24.395 58.180 24.825 ;
        RECT 59.075 24.640 59.335 24.960 ;
        RECT 60.560 24.645 60.820 27.245 ;
        RECT 61.890 24.990 62.360 32.410 ;
        RECT 62.850 25.775 63.740 32.695 ;
        RECT 64.420 32.390 64.650 32.490 ;
        RECT 64.420 32.380 64.775 32.390 ;
        RECT 65.560 32.380 65.790 32.490 ;
        RECT 59.130 24.480 59.280 24.640 ;
        RECT 54.510 23.355 55.385 23.360 ;
        RECT 53.580 22.950 55.385 23.355 ;
        RECT 53.580 22.110 53.880 22.950 ;
        RECT 54.510 22.935 55.385 22.950 ;
        RECT 54.875 22.825 55.385 22.935 ;
        RECT 54.875 22.125 55.390 22.825 ;
        RECT 55.585 22.795 56.615 23.795 ;
        RECT 51.275 21.965 51.615 21.970 ;
        RECT 51.250 20.020 51.615 21.965 ;
        RECT 52.830 21.900 53.060 21.970 ;
        RECT 52.335 21.230 53.060 21.900 ;
        RECT 52.325 21.040 53.060 21.230 ;
        RECT 52.325 20.240 52.680 21.040 ;
        RECT 52.830 20.970 53.060 21.040 ;
        RECT 53.270 21.925 53.500 21.970 ;
        RECT 53.640 21.925 53.880 22.110 ;
        RECT 53.270 21.595 53.880 21.925 ;
        RECT 54.855 21.870 55.085 21.975 ;
        RECT 53.270 21.040 53.765 21.595 ;
        RECT 53.270 20.970 53.500 21.040 ;
        RECT 53.020 20.785 53.310 20.810 ;
        RECT 53.005 20.535 53.340 20.785 ;
        RECT 54.625 20.765 55.085 21.870 ;
        RECT 54.305 20.240 55.085 20.765 ;
        RECT 51.885 20.060 55.085 20.240 ;
        RECT 51.250 19.965 51.480 20.020 ;
        RECT 47.240 19.575 51.200 19.805 ;
        RECT 51.885 19.620 54.690 20.060 ;
        RECT 54.855 19.975 55.085 20.060 ;
        RECT 55.295 21.910 55.525 21.975 ;
        RECT 55.690 21.910 56.060 22.795 ;
        RECT 55.295 21.585 56.060 21.910 ;
        RECT 55.295 20.045 56.055 21.585 ;
        RECT 55.295 19.975 55.525 20.045 ;
        RECT 55.045 19.795 55.335 19.815 ;
        RECT 51.885 19.255 54.350 19.620 ;
        RECT 55.020 19.545 55.355 19.795 ;
        RECT 57.590 19.280 58.085 24.395 ;
        RECT 59.105 24.345 59.310 24.480 ;
        RECT 60.590 24.395 60.820 24.645 ;
        RECT 61.610 24.550 62.360 24.990 ;
        RECT 62.780 24.775 63.795 25.775 ;
        RECT 58.385 24.115 60.385 24.345 ;
        RECT 61.610 22.355 61.980 24.550 ;
        RECT 62.130 24.490 62.360 24.550 ;
        RECT 62.850 24.285 63.740 24.775 ;
        RECT 64.420 24.580 65.790 32.380 ;
        RECT 66.325 27.635 67.215 32.695 ;
        RECT 67.850 32.410 68.080 32.490 ;
        RECT 66.320 26.015 67.220 27.635 ;
        RECT 66.325 25.605 67.215 26.015 ;
        RECT 66.250 24.605 67.280 25.605 ;
        RECT 67.850 24.625 68.225 32.410 ;
        RECT 68.500 32.025 70.180 33.260 ;
        RECT 71.015 32.025 75.940 32.035 ;
        RECT 68.500 31.545 75.940 32.025 ;
        RECT 68.500 29.285 70.180 31.545 ;
        RECT 71.015 31.125 75.940 31.545 ;
        RECT 70.520 30.935 70.775 30.960 ;
        RECT 70.520 30.920 70.795 30.935 ;
        RECT 70.490 30.645 70.825 30.920 ;
        RECT 71.000 30.895 76.000 31.125 ;
        RECT 76.210 30.935 76.465 30.960 ;
        RECT 70.520 30.630 70.775 30.645 ;
        RECT 71.000 30.455 76.000 30.685 ;
        RECT 76.205 30.645 76.465 30.935 ;
        RECT 76.210 30.630 76.465 30.645 ;
        RECT 71.045 30.445 75.900 30.455 ;
        RECT 71.045 28.920 73.690 28.925 ;
        RECT 69.720 28.720 73.690 28.920 ;
        RECT 69.720 28.690 73.680 28.720 ;
        RECT 68.560 28.335 68.895 28.610 ;
        RECT 69.440 28.440 69.670 28.485 ;
        RECT 64.420 24.560 64.775 24.580 ;
        RECT 64.420 24.490 64.650 24.560 ;
        RECT 65.560 24.490 65.790 24.580 ;
        RECT 66.320 24.465 67.230 24.605 ;
        RECT 67.850 24.490 68.240 24.625 ;
        RECT 66.310 24.285 67.320 24.465 ;
        RECT 62.410 24.055 64.370 24.285 ;
        RECT 65.840 24.055 67.800 24.285 ;
        RECT 63.165 23.050 63.510 24.055 ;
        RECT 65.865 24.050 67.750 24.055 ;
        RECT 68.045 22.355 68.240 24.490 ;
        RECT 68.630 22.830 68.820 28.335 ;
        RECT 69.250 27.105 69.670 28.440 ;
        RECT 70.975 27.105 72.320 28.690 ;
        RECT 69.250 25.720 72.320 27.105 ;
        RECT 69.250 24.990 69.670 25.720 ;
        RECT 69.245 24.485 69.670 24.990 ;
        RECT 68.630 22.640 68.945 22.830 ;
        RECT 58.950 22.125 62.910 22.355 ;
        RECT 64.380 22.125 68.340 22.355 ;
        RECT 68.755 22.130 68.945 22.640 ;
        RECT 58.670 21.515 58.900 21.965 ;
        RECT 60.150 21.515 60.940 22.125 ;
        RECT 58.670 21.210 60.940 21.515 ;
        RECT 58.615 21.195 60.940 21.210 ;
        RECT 58.530 20.350 60.940 21.195 ;
        RECT 58.530 19.975 58.900 20.350 ;
        RECT 58.670 19.965 58.900 19.975 ;
        RECT 60.150 19.805 60.940 20.350 ;
        RECT 62.960 21.880 63.190 21.965 ;
        RECT 64.100 21.880 64.330 21.965 ;
        RECT 62.960 20.055 64.330 21.880 ;
        RECT 62.960 19.965 63.190 20.055 ;
        RECT 58.950 19.575 62.910 19.805 ;
        RECT 55.490 19.255 58.085 19.280 ;
        RECT 58.530 19.255 58.755 19.265 ;
        RECT 63.430 19.255 63.920 20.055 ;
        RECT 64.100 19.965 64.330 20.055 ;
        RECT 65.815 21.745 67.155 22.125 ;
        RECT 68.390 21.745 68.620 21.965 ;
        RECT 65.815 20.150 68.620 21.745 ;
        RECT 65.815 19.805 67.155 20.150 ;
        RECT 68.390 19.965 68.620 20.150 ;
        RECT 64.380 19.575 68.340 19.805 ;
        RECT 68.770 19.785 68.945 22.130 ;
        RECT 69.245 21.965 69.540 24.485 ;
        RECT 70.975 24.280 72.320 25.720 ;
        RECT 73.730 28.390 73.960 28.485 ;
        RECT 74.205 28.390 74.695 30.445 ;
        RECT 75.265 28.920 75.900 28.925 ;
        RECT 75.150 28.690 79.110 28.920 ;
        RECT 74.870 28.390 75.100 28.485 ;
        RECT 73.730 24.565 75.100 28.390 ;
        RECT 73.730 24.485 73.960 24.565 ;
        RECT 74.870 24.485 75.100 24.565 ;
        RECT 76.525 24.280 77.870 28.690 ;
        RECT 79.160 28.420 79.390 28.485 ;
        RECT 80.045 28.425 80.520 33.260 ;
        RECT 81.845 32.455 82.525 33.260 ;
        RECT 82.945 32.735 83.280 32.985 ;
        RECT 82.960 32.710 83.250 32.735 ;
        RECT 86.420 32.635 88.330 33.260 ;
        RECT 90.420 32.925 92.305 32.930 ;
        RECT 93.865 32.925 95.750 32.930 ;
        RECT 90.410 32.695 92.370 32.925 ;
        RECT 93.840 32.695 95.800 32.925 ;
        RECT 82.770 32.455 83.000 32.505 ;
        RECT 81.845 31.955 83.000 32.455 ;
        RECT 80.915 28.735 81.250 28.985 ;
        RECT 80.935 28.705 81.225 28.735 ;
        RECT 80.745 28.425 80.975 28.500 ;
        RECT 79.160 24.485 79.615 28.420 ;
        RECT 80.045 27.680 80.975 28.425 ;
        RECT 80.380 24.565 80.975 27.680 ;
        RECT 80.745 24.500 80.975 24.565 ;
        RECT 81.185 28.475 81.415 28.500 ;
        RECT 81.185 24.920 81.695 28.475 ;
        RECT 81.185 24.550 81.880 24.920 ;
        RECT 82.380 24.600 83.000 31.955 ;
        RECT 81.185 24.500 81.415 24.550 ;
        RECT 69.720 24.250 73.680 24.280 ;
        RECT 75.150 24.250 79.110 24.280 ;
        RECT 69.720 24.090 79.110 24.250 ;
        RECT 69.720 24.050 73.680 24.090 ;
        RECT 75.150 24.050 79.110 24.090 ;
        RECT 79.275 22.660 79.615 24.485 ;
        RECT 80.925 22.660 81.345 24.305 ;
        RECT 79.275 22.505 81.345 22.660 ;
        RECT 79.350 22.390 81.345 22.505 ;
        RECT 69.810 22.125 73.770 22.355 ;
        RECT 75.240 22.125 79.200 22.355 ;
        RECT 69.245 21.205 69.760 21.965 ;
        RECT 69.315 20.025 69.760 21.205 ;
        RECT 69.530 19.965 69.760 20.025 ;
        RECT 71.190 19.805 72.145 22.125 ;
        RECT 73.820 21.900 74.050 21.965 ;
        RECT 74.960 21.900 75.190 21.965 ;
        RECT 73.820 20.030 75.190 21.900 ;
        RECT 73.820 19.965 74.050 20.030 ;
        RECT 68.755 19.255 68.945 19.785 ;
        RECT 69.810 19.575 73.770 19.805 ;
        RECT 74.225 19.255 74.780 20.030 ;
        RECT 74.960 19.965 75.190 20.030 ;
        RECT 76.635 19.805 77.590 22.125 ;
        RECT 79.350 21.970 79.615 22.390 ;
        RECT 80.925 22.115 81.345 22.390 ;
        RECT 81.580 23.355 81.880 24.550 ;
        RECT 82.770 24.505 83.000 24.600 ;
        RECT 83.210 32.430 83.440 32.505 ;
        RECT 83.210 25.110 83.985 32.430 ;
        RECT 86.385 32.405 88.385 32.635 ;
        RECT 90.130 32.410 90.360 32.490 ;
        RECT 85.950 29.060 86.180 32.355 ;
        RECT 88.590 32.275 88.820 32.355 ;
        RECT 88.560 29.060 88.820 32.275 ;
        RECT 85.950 27.245 88.820 29.060 ;
        RECT 83.210 24.580 84.060 25.110 ;
        RECT 85.950 24.825 86.180 27.245 ;
        RECT 83.210 24.505 83.440 24.580 ;
        RECT 82.875 23.825 83.390 24.315 ;
        RECT 82.875 23.360 83.385 23.825 ;
        RECT 83.690 23.795 84.060 24.580 ;
        RECT 85.590 24.395 86.180 24.825 ;
        RECT 87.075 24.640 87.335 24.960 ;
        RECT 88.560 24.645 88.820 27.245 ;
        RECT 89.890 24.990 90.360 32.410 ;
        RECT 90.850 25.775 91.740 32.695 ;
        RECT 92.420 32.390 92.650 32.490 ;
        RECT 92.420 32.380 92.775 32.390 ;
        RECT 93.560 32.380 93.790 32.490 ;
        RECT 87.130 24.480 87.280 24.640 ;
        RECT 82.510 23.355 83.385 23.360 ;
        RECT 81.580 22.950 83.385 23.355 ;
        RECT 81.580 22.110 81.880 22.950 ;
        RECT 82.510 22.935 83.385 22.950 ;
        RECT 82.875 22.825 83.385 22.935 ;
        RECT 82.875 22.125 83.390 22.825 ;
        RECT 83.615 22.795 84.645 23.795 ;
        RECT 79.275 21.965 79.615 21.970 ;
        RECT 79.250 20.020 79.615 21.965 ;
        RECT 80.830 21.900 81.060 21.970 ;
        RECT 80.335 21.230 81.060 21.900 ;
        RECT 80.325 21.040 81.060 21.230 ;
        RECT 80.325 20.240 80.680 21.040 ;
        RECT 80.830 20.970 81.060 21.040 ;
        RECT 81.270 21.925 81.500 21.970 ;
        RECT 81.640 21.925 81.880 22.110 ;
        RECT 81.270 21.595 81.880 21.925 ;
        RECT 82.855 21.870 83.085 21.975 ;
        RECT 81.270 21.040 81.765 21.595 ;
        RECT 81.270 20.970 81.500 21.040 ;
        RECT 81.020 20.785 81.310 20.810 ;
        RECT 81.005 20.535 81.340 20.785 ;
        RECT 82.625 20.765 83.085 21.870 ;
        RECT 82.305 20.240 83.085 20.765 ;
        RECT 79.885 20.060 83.085 20.240 ;
        RECT 79.250 19.965 79.480 20.020 ;
        RECT 75.240 19.575 79.200 19.805 ;
        RECT 79.885 19.620 82.690 20.060 ;
        RECT 82.855 19.975 83.085 20.060 ;
        RECT 83.295 21.910 83.525 21.975 ;
        RECT 83.690 21.910 84.060 22.795 ;
        RECT 83.295 21.585 84.060 21.910 ;
        RECT 83.295 20.045 84.055 21.585 ;
        RECT 83.295 19.975 83.525 20.045 ;
        RECT 83.045 19.795 83.335 19.815 ;
        RECT 79.885 19.255 82.350 19.620 ;
        RECT 83.020 19.545 83.355 19.795 ;
        RECT 85.590 19.280 86.085 24.395 ;
        RECT 87.105 24.345 87.310 24.480 ;
        RECT 88.590 24.395 88.820 24.645 ;
        RECT 89.610 24.550 90.360 24.990 ;
        RECT 90.780 24.775 91.795 25.775 ;
        RECT 86.385 24.115 88.385 24.345 ;
        RECT 89.610 22.355 89.980 24.550 ;
        RECT 90.130 24.490 90.360 24.550 ;
        RECT 90.850 24.285 91.740 24.775 ;
        RECT 92.420 24.580 93.790 32.380 ;
        RECT 94.325 27.635 95.215 32.695 ;
        RECT 95.850 32.410 96.080 32.490 ;
        RECT 94.320 26.015 95.220 27.635 ;
        RECT 94.325 25.605 95.215 26.015 ;
        RECT 94.250 24.605 95.280 25.605 ;
        RECT 95.850 24.625 96.225 32.410 ;
        RECT 96.500 32.025 98.180 33.260 ;
        RECT 99.015 32.025 103.940 32.035 ;
        RECT 96.500 31.545 103.940 32.025 ;
        RECT 96.500 29.285 98.180 31.545 ;
        RECT 99.015 31.125 103.940 31.545 ;
        RECT 98.520 30.935 98.775 30.960 ;
        RECT 98.520 30.920 98.795 30.935 ;
        RECT 98.490 30.645 98.825 30.920 ;
        RECT 99.000 30.895 104.000 31.125 ;
        RECT 104.210 30.935 104.465 30.960 ;
        RECT 98.520 30.630 98.775 30.645 ;
        RECT 99.000 30.455 104.000 30.685 ;
        RECT 104.205 30.645 104.465 30.935 ;
        RECT 104.210 30.630 104.465 30.645 ;
        RECT 99.045 30.445 103.900 30.455 ;
        RECT 99.045 28.920 101.690 28.925 ;
        RECT 97.720 28.720 101.690 28.920 ;
        RECT 97.720 28.690 101.680 28.720 ;
        RECT 96.560 28.335 96.895 28.610 ;
        RECT 97.440 28.440 97.670 28.485 ;
        RECT 92.420 24.560 92.775 24.580 ;
        RECT 92.420 24.490 92.650 24.560 ;
        RECT 93.560 24.490 93.790 24.580 ;
        RECT 94.320 24.465 95.230 24.605 ;
        RECT 95.850 24.490 96.240 24.625 ;
        RECT 94.310 24.285 95.320 24.465 ;
        RECT 90.410 24.055 92.370 24.285 ;
        RECT 93.840 24.055 95.800 24.285 ;
        RECT 91.125 22.980 91.525 24.055 ;
        RECT 93.865 24.050 95.750 24.055 ;
        RECT 96.045 22.355 96.240 24.490 ;
        RECT 96.630 22.830 96.820 28.335 ;
        RECT 97.250 27.105 97.670 28.440 ;
        RECT 98.975 27.105 100.320 28.690 ;
        RECT 97.250 25.720 100.320 27.105 ;
        RECT 97.250 24.990 97.670 25.720 ;
        RECT 97.245 24.485 97.670 24.990 ;
        RECT 96.630 22.640 96.945 22.830 ;
        RECT 86.950 22.125 90.910 22.355 ;
        RECT 92.380 22.125 96.340 22.355 ;
        RECT 96.755 22.130 96.945 22.640 ;
        RECT 86.670 21.515 86.900 21.965 ;
        RECT 88.150 21.515 88.940 22.125 ;
        RECT 86.670 21.210 88.940 21.515 ;
        RECT 86.615 21.195 88.940 21.210 ;
        RECT 86.530 20.350 88.940 21.195 ;
        RECT 86.530 19.975 86.900 20.350 ;
        RECT 86.670 19.965 86.900 19.975 ;
        RECT 88.150 19.805 88.940 20.350 ;
        RECT 90.960 21.880 91.190 21.965 ;
        RECT 92.100 21.880 92.330 21.965 ;
        RECT 90.960 20.055 92.330 21.880 ;
        RECT 90.960 19.965 91.190 20.055 ;
        RECT 86.950 19.575 90.910 19.805 ;
        RECT 83.790 19.255 86.085 19.280 ;
        RECT 86.530 19.255 86.755 19.265 ;
        RECT 91.430 19.255 91.920 20.055 ;
        RECT 92.100 19.965 92.330 20.055 ;
        RECT 93.815 21.745 95.155 22.125 ;
        RECT 96.390 21.745 96.620 21.965 ;
        RECT 93.815 20.150 96.620 21.745 ;
        RECT 93.815 19.805 95.155 20.150 ;
        RECT 96.390 19.965 96.620 20.150 ;
        RECT 92.380 19.575 96.340 19.805 ;
        RECT 96.770 19.785 96.945 22.130 ;
        RECT 97.245 21.965 97.540 24.485 ;
        RECT 98.975 24.280 100.320 25.720 ;
        RECT 101.730 28.390 101.960 28.485 ;
        RECT 102.205 28.390 102.695 30.445 ;
        RECT 103.265 28.920 103.900 28.925 ;
        RECT 103.150 28.690 107.110 28.920 ;
        RECT 102.870 28.390 103.100 28.485 ;
        RECT 101.730 24.565 103.100 28.390 ;
        RECT 101.730 24.485 101.960 24.565 ;
        RECT 102.870 24.485 103.100 24.565 ;
        RECT 104.525 24.280 105.870 28.690 ;
        RECT 107.160 28.420 107.390 28.485 ;
        RECT 108.045 28.425 108.520 33.260 ;
        RECT 109.845 32.455 110.525 33.260 ;
        RECT 110.945 32.735 111.280 32.985 ;
        RECT 110.960 32.710 111.250 32.735 ;
        RECT 114.420 32.635 116.330 33.260 ;
        RECT 118.420 32.925 120.305 32.930 ;
        RECT 121.865 32.925 123.750 32.930 ;
        RECT 118.410 32.695 120.370 32.925 ;
        RECT 121.840 32.695 123.800 32.925 ;
        RECT 110.770 32.455 111.000 32.505 ;
        RECT 109.845 31.955 111.000 32.455 ;
        RECT 108.915 28.735 109.250 28.985 ;
        RECT 108.935 28.705 109.225 28.735 ;
        RECT 108.745 28.425 108.975 28.500 ;
        RECT 107.160 24.485 107.615 28.420 ;
        RECT 108.045 27.680 108.975 28.425 ;
        RECT 108.380 24.565 108.975 27.680 ;
        RECT 108.745 24.500 108.975 24.565 ;
        RECT 109.185 28.475 109.415 28.500 ;
        RECT 109.185 24.920 109.695 28.475 ;
        RECT 109.185 24.550 109.880 24.920 ;
        RECT 110.380 24.600 111.000 31.955 ;
        RECT 109.185 24.500 109.415 24.550 ;
        RECT 97.720 24.250 101.680 24.280 ;
        RECT 103.150 24.250 107.110 24.280 ;
        RECT 97.720 24.090 107.110 24.250 ;
        RECT 97.720 24.050 101.680 24.090 ;
        RECT 103.150 24.050 107.110 24.090 ;
        RECT 107.275 22.660 107.615 24.485 ;
        RECT 108.925 22.660 109.345 24.305 ;
        RECT 107.275 22.505 109.345 22.660 ;
        RECT 107.350 22.390 109.345 22.505 ;
        RECT 97.810 22.125 101.770 22.355 ;
        RECT 103.240 22.125 107.200 22.355 ;
        RECT 97.245 21.205 97.760 21.965 ;
        RECT 97.315 20.025 97.760 21.205 ;
        RECT 97.530 19.965 97.760 20.025 ;
        RECT 99.190 19.805 100.145 22.125 ;
        RECT 101.820 21.900 102.050 21.965 ;
        RECT 102.960 21.900 103.190 21.965 ;
        RECT 101.820 20.030 103.190 21.900 ;
        RECT 101.820 19.965 102.050 20.030 ;
        RECT 96.755 19.255 96.945 19.785 ;
        RECT 97.810 19.575 101.770 19.805 ;
        RECT 102.225 19.255 102.780 20.030 ;
        RECT 102.960 19.965 103.190 20.030 ;
        RECT 104.635 19.805 105.590 22.125 ;
        RECT 107.350 21.970 107.615 22.390 ;
        RECT 108.925 22.115 109.345 22.390 ;
        RECT 109.580 23.355 109.880 24.550 ;
        RECT 110.770 24.505 111.000 24.600 ;
        RECT 111.210 32.430 111.440 32.505 ;
        RECT 111.210 25.110 111.985 32.430 ;
        RECT 114.385 32.405 116.385 32.635 ;
        RECT 118.130 32.410 118.360 32.490 ;
        RECT 113.950 29.060 114.180 32.355 ;
        RECT 116.590 32.275 116.820 32.355 ;
        RECT 116.560 29.060 116.820 32.275 ;
        RECT 113.950 27.245 116.820 29.060 ;
        RECT 111.210 24.580 112.060 25.110 ;
        RECT 113.950 24.825 114.180 27.245 ;
        RECT 111.210 24.505 111.440 24.580 ;
        RECT 110.875 23.825 111.390 24.315 ;
        RECT 110.875 23.360 111.385 23.825 ;
        RECT 111.690 23.795 112.060 24.580 ;
        RECT 113.590 24.395 114.180 24.825 ;
        RECT 115.075 24.640 115.335 24.960 ;
        RECT 116.560 24.645 116.820 27.245 ;
        RECT 117.890 24.990 118.360 32.410 ;
        RECT 118.850 25.775 119.740 32.695 ;
        RECT 120.420 32.390 120.650 32.490 ;
        RECT 120.420 32.380 120.775 32.390 ;
        RECT 121.560 32.380 121.790 32.490 ;
        RECT 115.130 24.480 115.280 24.640 ;
        RECT 110.510 23.355 111.385 23.360 ;
        RECT 109.580 22.950 111.385 23.355 ;
        RECT 109.580 22.110 109.880 22.950 ;
        RECT 110.510 22.935 111.385 22.950 ;
        RECT 110.875 22.825 111.385 22.935 ;
        RECT 110.875 22.125 111.390 22.825 ;
        RECT 111.585 22.795 112.615 23.795 ;
        RECT 107.275 21.965 107.615 21.970 ;
        RECT 107.250 20.020 107.615 21.965 ;
        RECT 108.830 21.900 109.060 21.970 ;
        RECT 108.335 21.230 109.060 21.900 ;
        RECT 108.325 21.040 109.060 21.230 ;
        RECT 108.325 20.240 108.680 21.040 ;
        RECT 108.830 20.970 109.060 21.040 ;
        RECT 109.270 21.925 109.500 21.970 ;
        RECT 109.640 21.925 109.880 22.110 ;
        RECT 109.270 21.595 109.880 21.925 ;
        RECT 110.855 21.870 111.085 21.975 ;
        RECT 109.270 21.040 109.765 21.595 ;
        RECT 109.270 20.970 109.500 21.040 ;
        RECT 109.020 20.785 109.310 20.810 ;
        RECT 109.005 20.535 109.340 20.785 ;
        RECT 110.625 20.765 111.085 21.870 ;
        RECT 110.305 20.240 111.085 20.765 ;
        RECT 107.885 20.060 111.085 20.240 ;
        RECT 107.250 19.965 107.480 20.020 ;
        RECT 103.240 19.575 107.200 19.805 ;
        RECT 107.885 19.620 110.690 20.060 ;
        RECT 110.855 19.975 111.085 20.060 ;
        RECT 111.295 21.910 111.525 21.975 ;
        RECT 111.690 21.910 112.060 22.795 ;
        RECT 111.295 21.585 112.060 21.910 ;
        RECT 111.295 20.045 112.055 21.585 ;
        RECT 111.295 19.975 111.525 20.045 ;
        RECT 111.045 19.795 111.335 19.815 ;
        RECT 107.885 19.255 110.350 19.620 ;
        RECT 111.020 19.545 111.355 19.795 ;
        RECT 113.590 19.255 114.085 24.395 ;
        RECT 115.105 24.345 115.310 24.480 ;
        RECT 116.590 24.395 116.820 24.645 ;
        RECT 117.610 24.550 118.360 24.990 ;
        RECT 118.780 24.775 119.795 25.775 ;
        RECT 114.385 24.115 116.385 24.345 ;
        RECT 117.610 22.355 117.980 24.550 ;
        RECT 118.130 24.490 118.360 24.550 ;
        RECT 118.850 24.285 119.740 24.775 ;
        RECT 120.420 24.580 121.790 32.380 ;
        RECT 122.325 27.635 123.215 32.695 ;
        RECT 123.850 32.410 124.080 32.490 ;
        RECT 122.320 26.015 123.220 27.635 ;
        RECT 122.325 25.605 123.215 26.015 ;
        RECT 122.250 24.605 123.280 25.605 ;
        RECT 123.850 24.625 124.225 32.410 ;
        RECT 124.500 32.025 126.180 33.260 ;
        RECT 127.015 32.025 131.940 32.035 ;
        RECT 124.500 31.545 131.940 32.025 ;
        RECT 124.500 29.285 126.180 31.545 ;
        RECT 127.015 31.125 131.940 31.545 ;
        RECT 126.520 30.935 126.775 30.960 ;
        RECT 126.520 30.920 126.795 30.935 ;
        RECT 126.490 30.645 126.825 30.920 ;
        RECT 127.000 30.895 132.000 31.125 ;
        RECT 132.210 30.935 132.465 30.960 ;
        RECT 126.520 30.630 126.775 30.645 ;
        RECT 127.000 30.455 132.000 30.685 ;
        RECT 132.205 30.645 132.465 30.935 ;
        RECT 132.210 30.630 132.465 30.645 ;
        RECT 127.045 30.445 131.900 30.455 ;
        RECT 127.045 28.920 129.690 28.925 ;
        RECT 125.720 28.720 129.690 28.920 ;
        RECT 125.720 28.690 129.680 28.720 ;
        RECT 124.560 28.335 124.895 28.610 ;
        RECT 125.440 28.440 125.670 28.485 ;
        RECT 120.420 24.560 120.775 24.580 ;
        RECT 120.420 24.490 120.650 24.560 ;
        RECT 121.560 24.490 121.790 24.580 ;
        RECT 122.320 24.465 123.230 24.605 ;
        RECT 123.850 24.490 124.240 24.625 ;
        RECT 122.310 24.285 123.320 24.465 ;
        RECT 118.410 24.055 120.370 24.285 ;
        RECT 121.840 24.055 123.800 24.285 ;
        RECT 119.160 23.115 119.445 24.055 ;
        RECT 121.865 24.050 123.750 24.055 ;
        RECT 124.045 22.355 124.240 24.490 ;
        RECT 124.630 22.830 124.820 28.335 ;
        RECT 125.250 27.105 125.670 28.440 ;
        RECT 126.975 27.105 128.320 28.690 ;
        RECT 125.250 25.720 128.320 27.105 ;
        RECT 125.250 24.990 125.670 25.720 ;
        RECT 125.245 24.485 125.670 24.990 ;
        RECT 124.630 22.640 124.945 22.830 ;
        RECT 114.950 22.125 118.910 22.355 ;
        RECT 120.380 22.125 124.340 22.355 ;
        RECT 124.755 22.130 124.945 22.640 ;
        RECT 114.670 21.515 114.900 21.965 ;
        RECT 116.150 21.515 116.940 22.125 ;
        RECT 114.670 21.210 116.940 21.515 ;
        RECT 114.615 21.195 116.940 21.210 ;
        RECT 114.530 20.350 116.940 21.195 ;
        RECT 114.530 19.975 114.900 20.350 ;
        RECT 114.670 19.965 114.900 19.975 ;
        RECT 116.150 19.805 116.940 20.350 ;
        RECT 118.960 21.880 119.190 21.965 ;
        RECT 120.100 21.880 120.330 21.965 ;
        RECT 118.960 20.055 120.330 21.880 ;
        RECT 118.960 19.965 119.190 20.055 ;
        RECT 114.950 19.575 118.910 19.805 ;
        RECT 114.530 19.255 114.755 19.265 ;
        RECT 119.430 19.255 119.920 20.055 ;
        RECT 120.100 19.965 120.330 20.055 ;
        RECT 121.815 21.745 123.155 22.125 ;
        RECT 124.390 21.745 124.620 21.965 ;
        RECT 121.815 20.150 124.620 21.745 ;
        RECT 121.815 19.805 123.155 20.150 ;
        RECT 124.390 19.965 124.620 20.150 ;
        RECT 120.380 19.575 124.340 19.805 ;
        RECT 124.770 19.785 124.945 22.130 ;
        RECT 125.245 21.965 125.540 24.485 ;
        RECT 126.975 24.280 128.320 25.720 ;
        RECT 129.730 28.390 129.960 28.485 ;
        RECT 130.205 28.390 130.695 30.445 ;
        RECT 131.265 28.920 131.900 28.925 ;
        RECT 131.150 28.690 135.110 28.920 ;
        RECT 130.870 28.390 131.100 28.485 ;
        RECT 129.730 24.565 131.100 28.390 ;
        RECT 129.730 24.485 129.960 24.565 ;
        RECT 130.870 24.485 131.100 24.565 ;
        RECT 132.525 24.280 133.870 28.690 ;
        RECT 135.160 28.420 135.390 28.485 ;
        RECT 136.045 28.425 136.520 33.260 ;
        RECT 137.845 32.455 138.525 33.260 ;
        RECT 138.945 32.735 139.280 32.985 ;
        RECT 138.960 32.710 139.250 32.735 ;
        RECT 138.770 32.455 139.000 32.505 ;
        RECT 137.845 31.955 139.000 32.455 ;
        RECT 136.915 28.735 137.250 28.985 ;
        RECT 136.935 28.705 137.225 28.735 ;
        RECT 136.745 28.425 136.975 28.500 ;
        RECT 135.160 24.485 135.615 28.420 ;
        RECT 136.045 27.680 136.975 28.425 ;
        RECT 136.380 24.565 136.975 27.680 ;
        RECT 136.745 24.500 136.975 24.565 ;
        RECT 137.185 28.475 137.415 28.500 ;
        RECT 137.185 24.920 137.695 28.475 ;
        RECT 137.185 24.550 137.880 24.920 ;
        RECT 138.380 24.600 139.000 31.955 ;
        RECT 137.185 24.500 137.415 24.550 ;
        RECT 125.720 24.250 129.680 24.280 ;
        RECT 131.150 24.250 135.110 24.280 ;
        RECT 125.720 24.090 135.110 24.250 ;
        RECT 125.720 24.050 129.680 24.090 ;
        RECT 131.150 24.050 135.110 24.090 ;
        RECT 135.275 22.660 135.615 24.485 ;
        RECT 136.925 22.660 137.345 24.305 ;
        RECT 135.275 22.505 137.345 22.660 ;
        RECT 135.350 22.390 137.345 22.505 ;
        RECT 125.810 22.125 129.770 22.355 ;
        RECT 131.240 22.125 135.200 22.355 ;
        RECT 125.245 21.205 125.760 21.965 ;
        RECT 125.315 20.025 125.760 21.205 ;
        RECT 125.530 19.965 125.760 20.025 ;
        RECT 127.190 19.805 128.145 22.125 ;
        RECT 129.820 21.900 130.050 21.965 ;
        RECT 130.960 21.900 131.190 21.965 ;
        RECT 129.820 20.030 131.190 21.900 ;
        RECT 129.820 19.965 130.050 20.030 ;
        RECT 124.755 19.255 124.945 19.785 ;
        RECT 125.810 19.575 129.770 19.805 ;
        RECT 130.225 19.255 130.780 20.030 ;
        RECT 130.960 19.965 131.190 20.030 ;
        RECT 132.635 19.805 133.590 22.125 ;
        RECT 135.350 21.970 135.615 22.390 ;
        RECT 136.925 22.115 137.345 22.390 ;
        RECT 137.580 23.355 137.880 24.550 ;
        RECT 138.770 24.505 139.000 24.600 ;
        RECT 139.210 32.430 139.440 32.505 ;
        RECT 139.210 25.110 139.985 32.430 ;
        RECT 139.210 24.580 140.060 25.110 ;
        RECT 139.210 24.505 139.440 24.580 ;
        RECT 138.875 23.825 139.390 24.315 ;
        RECT 138.875 23.360 139.385 23.825 ;
        RECT 139.690 23.795 140.060 24.580 ;
        RECT 138.510 23.355 139.385 23.360 ;
        RECT 137.580 22.950 139.385 23.355 ;
        RECT 137.580 22.110 137.880 22.950 ;
        RECT 138.510 22.935 139.385 22.950 ;
        RECT 138.875 22.825 139.385 22.935 ;
        RECT 138.875 22.125 139.390 22.825 ;
        RECT 139.615 22.795 140.645 23.795 ;
        RECT 135.275 21.965 135.615 21.970 ;
        RECT 135.250 20.020 135.615 21.965 ;
        RECT 136.830 21.900 137.060 21.970 ;
        RECT 136.335 21.230 137.060 21.900 ;
        RECT 136.325 21.040 137.060 21.230 ;
        RECT 136.325 20.240 136.680 21.040 ;
        RECT 136.830 20.970 137.060 21.040 ;
        RECT 137.270 21.925 137.500 21.970 ;
        RECT 137.640 21.925 137.880 22.110 ;
        RECT 137.270 21.595 137.880 21.925 ;
        RECT 138.855 21.870 139.085 21.975 ;
        RECT 137.270 21.040 137.765 21.595 ;
        RECT 137.270 20.970 137.500 21.040 ;
        RECT 137.020 20.785 137.310 20.810 ;
        RECT 137.005 20.535 137.340 20.785 ;
        RECT 138.625 20.765 139.085 21.870 ;
        RECT 138.305 20.240 139.085 20.765 ;
        RECT 135.885 20.060 139.085 20.240 ;
        RECT 135.250 19.965 135.480 20.020 ;
        RECT 131.240 19.575 135.200 19.805 ;
        RECT 135.885 19.620 138.690 20.060 ;
        RECT 138.855 19.975 139.085 20.060 ;
        RECT 139.295 21.910 139.525 21.975 ;
        RECT 139.690 21.910 140.060 22.795 ;
        RECT 139.295 21.585 140.060 21.910 ;
        RECT 139.295 20.045 140.055 21.585 ;
        RECT 139.295 19.975 139.525 20.045 ;
        RECT 139.045 19.795 139.335 19.815 ;
        RECT 135.885 19.255 138.350 19.620 ;
        RECT 139.020 19.545 139.355 19.795 ;
        RECT 1.475 18.380 112.080 19.255 ;
        RECT 113.475 18.380 140.080 19.255 ;
        RECT 27.790 17.960 30.690 17.980 ;
        RECT 55.390 17.960 57.890 17.980 ;
        RECT 68.845 17.960 69.785 17.985 ;
        RECT 83.690 17.960 86.190 17.980 ;
        RECT 1.450 17.280 111.925 17.960 ;
        RECT 1.450 17.260 27.925 17.280 ;
        RECT 29.450 17.260 55.925 17.280 ;
        RECT 57.450 17.260 83.925 17.280 ;
        RECT 85.450 17.260 111.925 17.280 ;
        RECT 113.450 17.260 139.925 17.960 ;
        RECT 2.420 16.635 4.330 17.260 ;
        RECT 6.420 16.925 8.305 16.930 ;
        RECT 9.865 16.925 11.750 16.930 ;
        RECT 6.410 16.695 8.370 16.925 ;
        RECT 9.840 16.695 11.800 16.925 ;
        RECT 2.385 16.405 4.385 16.635 ;
        RECT 6.130 16.410 6.360 16.490 ;
        RECT 1.950 13.060 2.180 16.355 ;
        RECT 4.590 16.275 4.820 16.355 ;
        RECT 4.560 13.060 4.820 16.275 ;
        RECT 1.950 11.245 4.820 13.060 ;
        RECT 1.950 8.825 2.180 11.245 ;
        RECT 1.590 8.395 2.180 8.825 ;
        RECT 3.075 8.640 3.335 8.960 ;
        RECT 4.560 8.645 4.820 11.245 ;
        RECT 5.890 8.990 6.360 16.410 ;
        RECT 6.850 9.775 7.740 16.695 ;
        RECT 8.420 16.390 8.650 16.490 ;
        RECT 8.420 16.380 8.775 16.390 ;
        RECT 9.560 16.380 9.790 16.490 ;
        RECT 3.130 8.480 3.280 8.640 ;
        RECT 1.590 3.255 2.085 8.395 ;
        RECT 3.105 8.345 3.310 8.480 ;
        RECT 4.590 8.395 4.820 8.645 ;
        RECT 5.610 8.550 6.360 8.990 ;
        RECT 6.780 8.775 7.795 9.775 ;
        RECT 2.385 8.115 4.385 8.345 ;
        RECT 5.610 6.355 5.980 8.550 ;
        RECT 6.130 8.490 6.360 8.550 ;
        RECT 6.850 8.285 7.740 8.775 ;
        RECT 8.420 8.580 9.790 16.380 ;
        RECT 10.325 11.635 11.215 16.695 ;
        RECT 11.850 16.410 12.080 16.490 ;
        RECT 10.320 10.015 11.220 11.635 ;
        RECT 10.325 9.605 11.215 10.015 ;
        RECT 10.250 8.605 11.280 9.605 ;
        RECT 11.850 8.625 12.225 16.410 ;
        RECT 12.500 16.025 14.180 17.260 ;
        RECT 15.015 16.025 19.940 16.035 ;
        RECT 12.500 15.545 19.940 16.025 ;
        RECT 12.500 13.285 14.180 15.545 ;
        RECT 15.015 15.125 19.940 15.545 ;
        RECT 14.520 14.935 14.775 14.960 ;
        RECT 14.520 14.920 14.795 14.935 ;
        RECT 14.490 14.645 14.825 14.920 ;
        RECT 15.000 14.895 20.000 15.125 ;
        RECT 20.210 14.935 20.465 14.960 ;
        RECT 14.520 14.630 14.775 14.645 ;
        RECT 15.000 14.455 20.000 14.685 ;
        RECT 20.205 14.645 20.465 14.935 ;
        RECT 20.210 14.630 20.465 14.645 ;
        RECT 15.045 14.445 19.900 14.455 ;
        RECT 15.045 12.920 17.690 12.925 ;
        RECT 13.720 12.720 17.690 12.920 ;
        RECT 13.720 12.690 17.680 12.720 ;
        RECT 12.560 12.335 12.895 12.610 ;
        RECT 13.440 12.440 13.670 12.485 ;
        RECT 8.420 8.560 8.775 8.580 ;
        RECT 8.420 8.490 8.650 8.560 ;
        RECT 9.560 8.490 9.790 8.580 ;
        RECT 10.320 8.465 11.230 8.605 ;
        RECT 11.850 8.490 12.240 8.625 ;
        RECT 10.310 8.285 11.320 8.465 ;
        RECT 6.410 8.055 8.370 8.285 ;
        RECT 9.840 8.055 11.800 8.285 ;
        RECT 7.130 7.085 7.460 8.055 ;
        RECT 9.865 8.050 11.750 8.055 ;
        RECT 12.045 6.355 12.240 8.490 ;
        RECT 12.630 6.830 12.820 12.335 ;
        RECT 13.250 11.105 13.670 12.440 ;
        RECT 14.975 11.105 16.320 12.690 ;
        RECT 13.250 9.720 16.320 11.105 ;
        RECT 13.250 8.990 13.670 9.720 ;
        RECT 13.245 8.485 13.670 8.990 ;
        RECT 12.630 6.640 12.945 6.830 ;
        RECT 2.950 6.125 6.910 6.355 ;
        RECT 8.380 6.125 12.340 6.355 ;
        RECT 12.755 6.130 12.945 6.640 ;
        RECT 2.670 5.515 2.900 5.965 ;
        RECT 4.150 5.515 4.940 6.125 ;
        RECT 2.670 5.210 4.940 5.515 ;
        RECT 2.615 5.195 4.940 5.210 ;
        RECT 2.530 4.350 4.940 5.195 ;
        RECT 2.530 3.975 2.900 4.350 ;
        RECT 2.670 3.965 2.900 3.975 ;
        RECT 4.150 3.805 4.940 4.350 ;
        RECT 6.960 5.880 7.190 5.965 ;
        RECT 8.100 5.880 8.330 5.965 ;
        RECT 6.960 4.055 8.330 5.880 ;
        RECT 6.960 3.965 7.190 4.055 ;
        RECT 2.950 3.575 6.910 3.805 ;
        RECT 2.530 3.255 2.755 3.265 ;
        RECT 7.430 3.255 7.920 4.055 ;
        RECT 8.100 3.965 8.330 4.055 ;
        RECT 9.815 5.745 11.155 6.125 ;
        RECT 12.390 5.745 12.620 5.965 ;
        RECT 9.815 4.150 12.620 5.745 ;
        RECT 9.815 3.805 11.155 4.150 ;
        RECT 12.390 3.965 12.620 4.150 ;
        RECT 8.380 3.575 12.340 3.805 ;
        RECT 12.770 3.785 12.945 6.130 ;
        RECT 13.245 5.965 13.540 8.485 ;
        RECT 14.975 8.280 16.320 9.720 ;
        RECT 17.730 12.390 17.960 12.485 ;
        RECT 18.205 12.390 18.695 14.445 ;
        RECT 19.265 12.920 19.900 12.925 ;
        RECT 19.150 12.690 23.110 12.920 ;
        RECT 18.870 12.390 19.100 12.485 ;
        RECT 17.730 8.565 19.100 12.390 ;
        RECT 17.730 8.485 17.960 8.565 ;
        RECT 18.870 8.485 19.100 8.565 ;
        RECT 20.525 8.280 21.870 12.690 ;
        RECT 23.160 12.420 23.390 12.485 ;
        RECT 24.045 12.425 24.520 17.260 ;
        RECT 25.845 16.455 26.525 17.260 ;
        RECT 26.945 16.735 27.280 16.985 ;
        RECT 26.960 16.710 27.250 16.735 ;
        RECT 30.420 16.635 32.330 17.260 ;
        RECT 34.420 16.925 36.305 16.930 ;
        RECT 37.865 16.925 39.750 16.930 ;
        RECT 34.410 16.695 36.370 16.925 ;
        RECT 37.840 16.695 39.800 16.925 ;
        RECT 26.770 16.455 27.000 16.505 ;
        RECT 25.845 15.955 27.000 16.455 ;
        RECT 24.915 12.735 25.250 12.985 ;
        RECT 24.935 12.705 25.225 12.735 ;
        RECT 24.745 12.425 24.975 12.500 ;
        RECT 23.160 8.485 23.615 12.420 ;
        RECT 24.045 11.680 24.975 12.425 ;
        RECT 24.380 8.565 24.975 11.680 ;
        RECT 24.745 8.500 24.975 8.565 ;
        RECT 25.185 12.475 25.415 12.500 ;
        RECT 25.185 8.920 25.695 12.475 ;
        RECT 25.185 8.550 25.880 8.920 ;
        RECT 26.380 8.600 27.000 15.955 ;
        RECT 25.185 8.500 25.415 8.550 ;
        RECT 13.720 8.250 17.680 8.280 ;
        RECT 19.150 8.250 23.110 8.280 ;
        RECT 13.720 8.090 23.110 8.250 ;
        RECT 13.720 8.050 17.680 8.090 ;
        RECT 19.150 8.050 23.110 8.090 ;
        RECT 23.275 6.660 23.615 8.485 ;
        RECT 24.925 6.660 25.345 8.305 ;
        RECT 23.275 6.505 25.345 6.660 ;
        RECT 23.350 6.390 25.345 6.505 ;
        RECT 13.810 6.125 17.770 6.355 ;
        RECT 19.240 6.125 23.200 6.355 ;
        RECT 13.245 5.205 13.760 5.965 ;
        RECT 13.315 4.025 13.760 5.205 ;
        RECT 13.530 3.965 13.760 4.025 ;
        RECT 15.190 3.805 16.145 6.125 ;
        RECT 17.820 5.900 18.050 5.965 ;
        RECT 18.960 5.900 19.190 5.965 ;
        RECT 17.820 4.030 19.190 5.900 ;
        RECT 17.820 3.965 18.050 4.030 ;
        RECT 12.755 3.255 12.945 3.785 ;
        RECT 13.810 3.575 17.770 3.805 ;
        RECT 18.225 3.255 18.780 4.030 ;
        RECT 18.960 3.965 19.190 4.030 ;
        RECT 20.635 3.805 21.590 6.125 ;
        RECT 23.350 5.970 23.615 6.390 ;
        RECT 24.925 6.115 25.345 6.390 ;
        RECT 25.580 7.355 25.880 8.550 ;
        RECT 26.770 8.505 27.000 8.600 ;
        RECT 27.210 16.430 27.440 16.505 ;
        RECT 27.210 9.110 27.985 16.430 ;
        RECT 30.385 16.405 32.385 16.635 ;
        RECT 34.130 16.410 34.360 16.490 ;
        RECT 29.950 13.060 30.180 16.355 ;
        RECT 32.590 16.275 32.820 16.355 ;
        RECT 32.560 13.060 32.820 16.275 ;
        RECT 29.950 11.245 32.820 13.060 ;
        RECT 27.210 8.580 28.060 9.110 ;
        RECT 29.950 8.825 30.180 11.245 ;
        RECT 27.210 8.505 27.440 8.580 ;
        RECT 26.875 7.825 27.390 8.315 ;
        RECT 27.690 7.825 28.060 8.580 ;
        RECT 29.590 8.395 30.180 8.825 ;
        RECT 31.075 8.640 31.335 8.960 ;
        RECT 32.560 8.645 32.820 11.245 ;
        RECT 33.890 8.990 34.360 16.410 ;
        RECT 34.850 9.775 35.740 16.695 ;
        RECT 36.420 16.390 36.650 16.490 ;
        RECT 36.420 16.380 36.775 16.390 ;
        RECT 37.560 16.380 37.790 16.490 ;
        RECT 31.130 8.480 31.280 8.640 ;
        RECT 26.875 7.360 27.385 7.825 ;
        RECT 26.510 7.355 27.385 7.360 ;
        RECT 25.580 6.950 27.385 7.355 ;
        RECT 25.580 6.110 25.880 6.950 ;
        RECT 26.510 6.935 27.385 6.950 ;
        RECT 26.875 6.825 27.385 6.935 ;
        RECT 26.875 6.125 27.390 6.825 ;
        RECT 27.615 6.795 28.615 7.825 ;
        RECT 23.275 5.965 23.615 5.970 ;
        RECT 23.250 4.020 23.615 5.965 ;
        RECT 24.830 5.900 25.060 5.970 ;
        RECT 24.335 5.230 25.060 5.900 ;
        RECT 24.325 5.040 25.060 5.230 ;
        RECT 24.325 4.240 24.680 5.040 ;
        RECT 24.830 4.970 25.060 5.040 ;
        RECT 25.270 5.925 25.500 5.970 ;
        RECT 25.640 5.925 25.880 6.110 ;
        RECT 25.270 5.595 25.880 5.925 ;
        RECT 26.855 5.870 27.085 5.975 ;
        RECT 25.270 5.040 25.765 5.595 ;
        RECT 25.270 4.970 25.500 5.040 ;
        RECT 25.020 4.785 25.310 4.810 ;
        RECT 25.005 4.535 25.340 4.785 ;
        RECT 26.625 4.765 27.085 5.870 ;
        RECT 26.305 4.240 27.085 4.765 ;
        RECT 23.885 4.060 27.085 4.240 ;
        RECT 23.250 3.965 23.480 4.020 ;
        RECT 19.240 3.575 23.200 3.805 ;
        RECT 23.885 3.620 26.690 4.060 ;
        RECT 26.855 3.975 27.085 4.060 ;
        RECT 27.295 5.910 27.525 5.975 ;
        RECT 27.690 5.910 28.060 6.795 ;
        RECT 27.295 5.585 28.060 5.910 ;
        RECT 27.295 4.045 28.055 5.585 ;
        RECT 27.295 3.975 27.525 4.045 ;
        RECT 27.045 3.795 27.335 3.815 ;
        RECT 23.885 3.255 26.350 3.620 ;
        RECT 27.020 3.545 27.355 3.795 ;
        RECT 29.590 3.280 30.085 8.395 ;
        RECT 31.105 8.345 31.310 8.480 ;
        RECT 32.590 8.395 32.820 8.645 ;
        RECT 33.610 8.550 34.360 8.990 ;
        RECT 34.780 8.775 35.795 9.775 ;
        RECT 30.385 8.115 32.385 8.345 ;
        RECT 33.610 6.355 33.980 8.550 ;
        RECT 34.130 8.490 34.360 8.550 ;
        RECT 34.850 8.285 35.740 8.775 ;
        RECT 36.420 8.580 37.790 16.380 ;
        RECT 38.325 11.635 39.215 16.695 ;
        RECT 39.850 16.410 40.080 16.490 ;
        RECT 38.320 10.015 39.220 11.635 ;
        RECT 38.325 9.605 39.215 10.015 ;
        RECT 38.250 8.605 39.280 9.605 ;
        RECT 39.850 8.625 40.225 16.410 ;
        RECT 40.500 16.025 42.180 17.260 ;
        RECT 43.015 16.025 47.940 16.035 ;
        RECT 40.500 15.545 47.940 16.025 ;
        RECT 40.500 13.285 42.180 15.545 ;
        RECT 43.015 15.125 47.940 15.545 ;
        RECT 42.520 14.935 42.775 14.960 ;
        RECT 42.520 14.920 42.795 14.935 ;
        RECT 42.490 14.645 42.825 14.920 ;
        RECT 43.000 14.895 48.000 15.125 ;
        RECT 48.210 14.935 48.465 14.960 ;
        RECT 42.520 14.630 42.775 14.645 ;
        RECT 43.000 14.455 48.000 14.685 ;
        RECT 48.205 14.645 48.465 14.935 ;
        RECT 48.210 14.630 48.465 14.645 ;
        RECT 43.045 14.445 47.900 14.455 ;
        RECT 43.045 12.920 45.690 12.925 ;
        RECT 41.720 12.720 45.690 12.920 ;
        RECT 41.720 12.690 45.680 12.720 ;
        RECT 40.560 12.335 40.895 12.610 ;
        RECT 41.440 12.440 41.670 12.485 ;
        RECT 36.420 8.560 36.775 8.580 ;
        RECT 36.420 8.490 36.650 8.560 ;
        RECT 37.560 8.490 37.790 8.580 ;
        RECT 38.320 8.465 39.230 8.605 ;
        RECT 39.850 8.490 40.240 8.625 ;
        RECT 38.310 8.285 39.320 8.465 ;
        RECT 34.410 8.055 36.370 8.285 ;
        RECT 37.840 8.055 39.800 8.285 ;
        RECT 35.210 7.040 35.560 8.055 ;
        RECT 37.865 8.050 39.750 8.055 ;
        RECT 40.045 6.355 40.240 8.490 ;
        RECT 40.630 6.830 40.820 12.335 ;
        RECT 41.250 11.105 41.670 12.440 ;
        RECT 42.975 11.105 44.320 12.690 ;
        RECT 41.250 9.720 44.320 11.105 ;
        RECT 41.250 8.990 41.670 9.720 ;
        RECT 41.245 8.485 41.670 8.990 ;
        RECT 40.630 6.640 40.945 6.830 ;
        RECT 30.950 6.125 34.910 6.355 ;
        RECT 36.380 6.125 40.340 6.355 ;
        RECT 40.755 6.130 40.945 6.640 ;
        RECT 30.670 5.515 30.900 5.965 ;
        RECT 32.150 5.515 32.940 6.125 ;
        RECT 30.670 5.210 32.940 5.515 ;
        RECT 30.615 5.195 32.940 5.210 ;
        RECT 30.530 4.350 32.940 5.195 ;
        RECT 30.530 3.975 30.900 4.350 ;
        RECT 30.670 3.965 30.900 3.975 ;
        RECT 32.150 3.805 32.940 4.350 ;
        RECT 34.960 5.880 35.190 5.965 ;
        RECT 36.100 5.880 36.330 5.965 ;
        RECT 34.960 4.055 36.330 5.880 ;
        RECT 34.960 3.965 35.190 4.055 ;
        RECT 30.950 3.575 34.910 3.805 ;
        RECT 27.990 3.255 30.090 3.280 ;
        RECT 30.530 3.255 30.755 3.265 ;
        RECT 35.430 3.255 35.920 4.055 ;
        RECT 36.100 3.965 36.330 4.055 ;
        RECT 37.815 5.745 39.155 6.125 ;
        RECT 40.390 5.745 40.620 5.965 ;
        RECT 37.815 4.150 40.620 5.745 ;
        RECT 37.815 3.805 39.155 4.150 ;
        RECT 40.390 3.965 40.620 4.150 ;
        RECT 36.380 3.575 40.340 3.805 ;
        RECT 40.770 3.785 40.945 6.130 ;
        RECT 41.245 5.965 41.540 8.485 ;
        RECT 42.975 8.280 44.320 9.720 ;
        RECT 45.730 12.390 45.960 12.485 ;
        RECT 46.205 12.390 46.695 14.445 ;
        RECT 47.265 12.920 47.900 12.925 ;
        RECT 47.150 12.690 51.110 12.920 ;
        RECT 46.870 12.390 47.100 12.485 ;
        RECT 45.730 8.565 47.100 12.390 ;
        RECT 45.730 8.485 45.960 8.565 ;
        RECT 46.870 8.485 47.100 8.565 ;
        RECT 48.525 8.280 49.870 12.690 ;
        RECT 51.160 12.420 51.390 12.485 ;
        RECT 52.045 12.425 52.520 17.260 ;
        RECT 53.845 16.455 54.525 17.260 ;
        RECT 54.945 16.735 55.280 16.985 ;
        RECT 54.960 16.710 55.250 16.735 ;
        RECT 58.420 16.635 60.330 17.260 ;
        RECT 62.420 16.925 64.305 16.930 ;
        RECT 65.865 16.925 67.750 16.930 ;
        RECT 62.410 16.695 64.370 16.925 ;
        RECT 65.840 16.695 67.800 16.925 ;
        RECT 54.770 16.455 55.000 16.505 ;
        RECT 53.845 15.955 55.000 16.455 ;
        RECT 52.915 12.735 53.250 12.985 ;
        RECT 52.935 12.705 53.225 12.735 ;
        RECT 52.745 12.425 52.975 12.500 ;
        RECT 51.160 8.485 51.615 12.420 ;
        RECT 52.045 11.680 52.975 12.425 ;
        RECT 52.380 8.565 52.975 11.680 ;
        RECT 52.745 8.500 52.975 8.565 ;
        RECT 53.185 12.475 53.415 12.500 ;
        RECT 53.185 8.920 53.695 12.475 ;
        RECT 53.185 8.550 53.880 8.920 ;
        RECT 54.380 8.600 55.000 15.955 ;
        RECT 53.185 8.500 53.415 8.550 ;
        RECT 41.720 8.250 45.680 8.280 ;
        RECT 47.150 8.250 51.110 8.280 ;
        RECT 41.720 8.090 51.110 8.250 ;
        RECT 41.720 8.050 45.680 8.090 ;
        RECT 47.150 8.050 51.110 8.090 ;
        RECT 51.275 6.660 51.615 8.485 ;
        RECT 52.925 6.660 53.345 8.305 ;
        RECT 51.275 6.505 53.345 6.660 ;
        RECT 51.350 6.390 53.345 6.505 ;
        RECT 41.810 6.125 45.770 6.355 ;
        RECT 47.240 6.125 51.200 6.355 ;
        RECT 41.245 5.205 41.760 5.965 ;
        RECT 41.315 4.025 41.760 5.205 ;
        RECT 41.530 3.965 41.760 4.025 ;
        RECT 43.190 3.805 44.145 6.125 ;
        RECT 45.820 5.900 46.050 5.965 ;
        RECT 46.960 5.900 47.190 5.965 ;
        RECT 45.820 4.030 47.190 5.900 ;
        RECT 45.820 3.965 46.050 4.030 ;
        RECT 40.755 3.255 40.945 3.785 ;
        RECT 41.810 3.575 45.770 3.805 ;
        RECT 46.225 3.255 46.780 4.030 ;
        RECT 46.960 3.965 47.190 4.030 ;
        RECT 48.635 3.805 49.590 6.125 ;
        RECT 51.350 5.970 51.615 6.390 ;
        RECT 52.925 6.115 53.345 6.390 ;
        RECT 53.580 7.355 53.880 8.550 ;
        RECT 54.770 8.505 55.000 8.600 ;
        RECT 55.210 16.430 55.440 16.505 ;
        RECT 55.210 9.110 55.985 16.430 ;
        RECT 58.385 16.405 60.385 16.635 ;
        RECT 62.130 16.410 62.360 16.490 ;
        RECT 57.950 13.060 58.180 16.355 ;
        RECT 60.590 16.275 60.820 16.355 ;
        RECT 60.560 13.060 60.820 16.275 ;
        RECT 57.950 11.245 60.820 13.060 ;
        RECT 55.210 8.580 56.060 9.110 ;
        RECT 57.950 8.825 58.180 11.245 ;
        RECT 55.210 8.505 55.440 8.580 ;
        RECT 54.875 7.825 55.390 8.315 ;
        RECT 54.875 7.360 55.385 7.825 ;
        RECT 55.690 7.795 56.060 8.580 ;
        RECT 57.590 8.395 58.180 8.825 ;
        RECT 59.075 8.640 59.335 8.960 ;
        RECT 60.560 8.645 60.820 11.245 ;
        RECT 61.890 8.990 62.360 16.410 ;
        RECT 62.850 9.775 63.740 16.695 ;
        RECT 64.420 16.390 64.650 16.490 ;
        RECT 64.420 16.380 64.775 16.390 ;
        RECT 65.560 16.380 65.790 16.490 ;
        RECT 59.130 8.480 59.280 8.640 ;
        RECT 54.510 7.355 55.385 7.360 ;
        RECT 53.580 6.950 55.385 7.355 ;
        RECT 53.580 6.110 53.880 6.950 ;
        RECT 54.510 6.935 55.385 6.950 ;
        RECT 54.875 6.825 55.385 6.935 ;
        RECT 54.875 6.125 55.390 6.825 ;
        RECT 55.615 6.795 56.645 7.795 ;
        RECT 51.275 5.965 51.615 5.970 ;
        RECT 51.250 4.020 51.615 5.965 ;
        RECT 52.830 5.900 53.060 5.970 ;
        RECT 52.335 5.230 53.060 5.900 ;
        RECT 52.325 5.040 53.060 5.230 ;
        RECT 52.325 4.240 52.680 5.040 ;
        RECT 52.830 4.970 53.060 5.040 ;
        RECT 53.270 5.925 53.500 5.970 ;
        RECT 53.640 5.925 53.880 6.110 ;
        RECT 53.270 5.595 53.880 5.925 ;
        RECT 54.855 5.870 55.085 5.975 ;
        RECT 53.270 5.040 53.765 5.595 ;
        RECT 53.270 4.970 53.500 5.040 ;
        RECT 53.020 4.785 53.310 4.810 ;
        RECT 53.005 4.535 53.340 4.785 ;
        RECT 54.625 4.765 55.085 5.870 ;
        RECT 54.305 4.240 55.085 4.765 ;
        RECT 51.885 4.060 55.085 4.240 ;
        RECT 51.250 3.965 51.480 4.020 ;
        RECT 47.240 3.575 51.200 3.805 ;
        RECT 51.885 3.620 54.690 4.060 ;
        RECT 54.855 3.975 55.085 4.060 ;
        RECT 55.295 5.910 55.525 5.975 ;
        RECT 55.690 5.910 56.060 6.795 ;
        RECT 55.295 5.585 56.060 5.910 ;
        RECT 55.295 4.045 56.055 5.585 ;
        RECT 55.295 3.975 55.525 4.045 ;
        RECT 55.045 3.795 55.335 3.815 ;
        RECT 51.885 3.255 54.350 3.620 ;
        RECT 55.020 3.545 55.355 3.795 ;
        RECT 57.590 3.280 58.085 8.395 ;
        RECT 59.105 8.345 59.310 8.480 ;
        RECT 60.590 8.395 60.820 8.645 ;
        RECT 61.610 8.550 62.360 8.990 ;
        RECT 62.780 8.775 63.795 9.775 ;
        RECT 58.385 8.115 60.385 8.345 ;
        RECT 61.610 6.355 61.980 8.550 ;
        RECT 62.130 8.490 62.360 8.550 ;
        RECT 62.850 8.285 63.740 8.775 ;
        RECT 64.420 8.580 65.790 16.380 ;
        RECT 66.325 11.635 67.215 16.695 ;
        RECT 67.850 16.410 68.080 16.490 ;
        RECT 66.320 10.015 67.220 11.635 ;
        RECT 66.325 9.605 67.215 10.015 ;
        RECT 66.250 8.605 67.280 9.605 ;
        RECT 67.850 8.625 68.225 16.410 ;
        RECT 68.500 16.025 70.180 17.260 ;
        RECT 71.015 16.025 75.940 16.035 ;
        RECT 68.500 15.545 75.940 16.025 ;
        RECT 68.500 13.285 70.180 15.545 ;
        RECT 71.015 15.125 75.940 15.545 ;
        RECT 70.520 14.935 70.775 14.960 ;
        RECT 70.520 14.920 70.795 14.935 ;
        RECT 70.490 14.645 70.825 14.920 ;
        RECT 71.000 14.895 76.000 15.125 ;
        RECT 76.210 14.935 76.465 14.960 ;
        RECT 70.520 14.630 70.775 14.645 ;
        RECT 71.000 14.455 76.000 14.685 ;
        RECT 76.205 14.645 76.465 14.935 ;
        RECT 76.210 14.630 76.465 14.645 ;
        RECT 71.045 14.445 75.900 14.455 ;
        RECT 71.045 12.920 73.690 12.925 ;
        RECT 69.720 12.720 73.690 12.920 ;
        RECT 69.720 12.690 73.680 12.720 ;
        RECT 68.560 12.335 68.895 12.610 ;
        RECT 69.440 12.440 69.670 12.485 ;
        RECT 64.420 8.560 64.775 8.580 ;
        RECT 64.420 8.490 64.650 8.560 ;
        RECT 65.560 8.490 65.790 8.580 ;
        RECT 66.320 8.465 67.230 8.605 ;
        RECT 67.850 8.490 68.240 8.625 ;
        RECT 66.310 8.285 67.320 8.465 ;
        RECT 62.410 8.055 64.370 8.285 ;
        RECT 65.840 8.055 67.800 8.285 ;
        RECT 63.125 7.090 63.470 8.055 ;
        RECT 65.865 8.050 67.750 8.055 ;
        RECT 68.045 6.355 68.240 8.490 ;
        RECT 68.630 6.830 68.820 12.335 ;
        RECT 69.250 11.105 69.670 12.440 ;
        RECT 70.975 11.105 72.320 12.690 ;
        RECT 69.250 9.720 72.320 11.105 ;
        RECT 69.250 8.990 69.670 9.720 ;
        RECT 69.245 8.485 69.670 8.990 ;
        RECT 68.630 6.640 68.945 6.830 ;
        RECT 58.950 6.125 62.910 6.355 ;
        RECT 64.380 6.125 68.340 6.355 ;
        RECT 68.755 6.130 68.945 6.640 ;
        RECT 58.670 5.515 58.900 5.965 ;
        RECT 60.150 5.515 60.940 6.125 ;
        RECT 58.670 5.210 60.940 5.515 ;
        RECT 58.615 5.195 60.940 5.210 ;
        RECT 58.530 4.350 60.940 5.195 ;
        RECT 58.530 3.975 58.900 4.350 ;
        RECT 58.670 3.965 58.900 3.975 ;
        RECT 60.150 3.805 60.940 4.350 ;
        RECT 62.960 5.880 63.190 5.965 ;
        RECT 64.100 5.880 64.330 5.965 ;
        RECT 62.960 4.055 64.330 5.880 ;
        RECT 62.960 3.965 63.190 4.055 ;
        RECT 58.950 3.575 62.910 3.805 ;
        RECT 55.790 3.255 58.085 3.280 ;
        RECT 58.530 3.255 58.755 3.265 ;
        RECT 63.430 3.255 63.920 4.055 ;
        RECT 64.100 3.965 64.330 4.055 ;
        RECT 65.815 5.745 67.155 6.125 ;
        RECT 68.390 5.745 68.620 5.965 ;
        RECT 65.815 4.150 68.620 5.745 ;
        RECT 65.815 3.805 67.155 4.150 ;
        RECT 68.390 3.965 68.620 4.150 ;
        RECT 64.380 3.575 68.340 3.805 ;
        RECT 68.770 3.785 68.945 6.130 ;
        RECT 69.245 5.965 69.540 8.485 ;
        RECT 70.975 8.280 72.320 9.720 ;
        RECT 73.730 12.390 73.960 12.485 ;
        RECT 74.205 12.390 74.695 14.445 ;
        RECT 75.265 12.920 75.900 12.925 ;
        RECT 75.150 12.690 79.110 12.920 ;
        RECT 74.870 12.390 75.100 12.485 ;
        RECT 73.730 8.565 75.100 12.390 ;
        RECT 73.730 8.485 73.960 8.565 ;
        RECT 74.870 8.485 75.100 8.565 ;
        RECT 76.525 8.280 77.870 12.690 ;
        RECT 79.160 12.420 79.390 12.485 ;
        RECT 80.045 12.425 80.520 17.260 ;
        RECT 81.845 16.455 82.525 17.260 ;
        RECT 82.945 16.735 83.280 16.985 ;
        RECT 82.960 16.710 83.250 16.735 ;
        RECT 86.420 16.635 88.330 17.260 ;
        RECT 90.420 16.925 92.305 16.930 ;
        RECT 93.865 16.925 95.750 16.930 ;
        RECT 90.410 16.695 92.370 16.925 ;
        RECT 93.840 16.695 95.800 16.925 ;
        RECT 82.770 16.455 83.000 16.505 ;
        RECT 81.845 15.955 83.000 16.455 ;
        RECT 80.915 12.735 81.250 12.985 ;
        RECT 80.935 12.705 81.225 12.735 ;
        RECT 80.745 12.425 80.975 12.500 ;
        RECT 79.160 8.485 79.615 12.420 ;
        RECT 80.045 11.680 80.975 12.425 ;
        RECT 80.380 8.565 80.975 11.680 ;
        RECT 80.745 8.500 80.975 8.565 ;
        RECT 81.185 12.475 81.415 12.500 ;
        RECT 81.185 8.920 81.695 12.475 ;
        RECT 81.185 8.550 81.880 8.920 ;
        RECT 82.380 8.600 83.000 15.955 ;
        RECT 81.185 8.500 81.415 8.550 ;
        RECT 69.720 8.250 73.680 8.280 ;
        RECT 75.150 8.250 79.110 8.280 ;
        RECT 69.720 8.090 79.110 8.250 ;
        RECT 69.720 8.050 73.680 8.090 ;
        RECT 75.150 8.050 79.110 8.090 ;
        RECT 79.275 6.660 79.615 8.485 ;
        RECT 80.925 6.660 81.345 8.305 ;
        RECT 79.275 6.505 81.345 6.660 ;
        RECT 79.350 6.390 81.345 6.505 ;
        RECT 69.810 6.125 73.770 6.355 ;
        RECT 75.240 6.125 79.200 6.355 ;
        RECT 69.245 5.205 69.760 5.965 ;
        RECT 69.315 4.025 69.760 5.205 ;
        RECT 69.530 3.965 69.760 4.025 ;
        RECT 71.190 3.805 72.145 6.125 ;
        RECT 73.820 5.900 74.050 5.965 ;
        RECT 74.960 5.900 75.190 5.965 ;
        RECT 73.820 4.030 75.190 5.900 ;
        RECT 73.820 3.965 74.050 4.030 ;
        RECT 68.755 3.255 68.945 3.785 ;
        RECT 69.810 3.575 73.770 3.805 ;
        RECT 74.225 3.255 74.780 4.030 ;
        RECT 74.960 3.965 75.190 4.030 ;
        RECT 76.635 3.805 77.590 6.125 ;
        RECT 79.350 5.970 79.615 6.390 ;
        RECT 80.925 6.115 81.345 6.390 ;
        RECT 81.580 7.355 81.880 8.550 ;
        RECT 82.770 8.505 83.000 8.600 ;
        RECT 83.210 16.430 83.440 16.505 ;
        RECT 83.210 9.110 83.985 16.430 ;
        RECT 86.385 16.405 88.385 16.635 ;
        RECT 90.130 16.410 90.360 16.490 ;
        RECT 85.950 13.060 86.180 16.355 ;
        RECT 88.590 16.275 88.820 16.355 ;
        RECT 88.560 13.060 88.820 16.275 ;
        RECT 85.950 11.245 88.820 13.060 ;
        RECT 83.210 8.580 84.060 9.110 ;
        RECT 85.950 8.825 86.180 11.245 ;
        RECT 83.210 8.505 83.440 8.580 ;
        RECT 82.875 7.825 83.390 8.315 ;
        RECT 82.875 7.360 83.385 7.825 ;
        RECT 83.690 7.795 84.060 8.580 ;
        RECT 85.590 8.395 86.180 8.825 ;
        RECT 87.075 8.640 87.335 8.960 ;
        RECT 88.560 8.645 88.820 11.245 ;
        RECT 89.890 8.990 90.360 16.410 ;
        RECT 90.850 9.775 91.740 16.695 ;
        RECT 92.420 16.390 92.650 16.490 ;
        RECT 92.420 16.380 92.775 16.390 ;
        RECT 93.560 16.380 93.790 16.490 ;
        RECT 87.130 8.480 87.280 8.640 ;
        RECT 82.510 7.355 83.385 7.360 ;
        RECT 81.580 6.950 83.385 7.355 ;
        RECT 81.580 6.110 81.880 6.950 ;
        RECT 82.510 6.935 83.385 6.950 ;
        RECT 82.875 6.825 83.385 6.935 ;
        RECT 82.875 6.125 83.390 6.825 ;
        RECT 83.615 6.795 84.645 7.795 ;
        RECT 79.275 5.965 79.615 5.970 ;
        RECT 79.250 4.020 79.615 5.965 ;
        RECT 80.830 5.900 81.060 5.970 ;
        RECT 80.335 5.230 81.060 5.900 ;
        RECT 80.325 5.040 81.060 5.230 ;
        RECT 80.325 4.240 80.680 5.040 ;
        RECT 80.830 4.970 81.060 5.040 ;
        RECT 81.270 5.925 81.500 5.970 ;
        RECT 81.640 5.925 81.880 6.110 ;
        RECT 81.270 5.595 81.880 5.925 ;
        RECT 82.855 5.870 83.085 5.975 ;
        RECT 81.270 5.040 81.765 5.595 ;
        RECT 81.270 4.970 81.500 5.040 ;
        RECT 81.020 4.785 81.310 4.810 ;
        RECT 81.005 4.535 81.340 4.785 ;
        RECT 82.625 4.765 83.085 5.870 ;
        RECT 82.305 4.240 83.085 4.765 ;
        RECT 79.885 4.060 83.085 4.240 ;
        RECT 79.250 3.965 79.480 4.020 ;
        RECT 75.240 3.575 79.200 3.805 ;
        RECT 79.885 3.620 82.690 4.060 ;
        RECT 82.855 3.975 83.085 4.060 ;
        RECT 83.295 5.910 83.525 5.975 ;
        RECT 83.690 5.910 84.060 6.795 ;
        RECT 83.295 5.585 84.060 5.910 ;
        RECT 83.295 4.045 84.055 5.585 ;
        RECT 83.295 3.975 83.525 4.045 ;
        RECT 83.045 3.795 83.335 3.815 ;
        RECT 79.885 3.255 82.350 3.620 ;
        RECT 83.020 3.545 83.355 3.795 ;
        RECT 85.590 3.280 86.085 8.395 ;
        RECT 87.105 8.345 87.310 8.480 ;
        RECT 88.590 8.395 88.820 8.645 ;
        RECT 89.610 8.550 90.360 8.990 ;
        RECT 90.780 8.775 91.795 9.775 ;
        RECT 86.385 8.115 88.385 8.345 ;
        RECT 89.610 6.355 89.980 8.550 ;
        RECT 90.130 8.490 90.360 8.550 ;
        RECT 90.850 8.285 91.740 8.775 ;
        RECT 92.420 8.580 93.790 16.380 ;
        RECT 94.325 11.635 95.215 16.695 ;
        RECT 95.850 16.410 96.080 16.490 ;
        RECT 94.320 10.015 95.220 11.635 ;
        RECT 94.325 9.605 95.215 10.015 ;
        RECT 94.250 8.605 95.280 9.605 ;
        RECT 95.850 8.625 96.225 16.410 ;
        RECT 96.500 16.025 98.180 17.260 ;
        RECT 99.015 16.025 103.940 16.035 ;
        RECT 96.500 15.545 103.940 16.025 ;
        RECT 96.500 13.285 98.180 15.545 ;
        RECT 99.015 15.125 103.940 15.545 ;
        RECT 98.520 14.935 98.775 14.960 ;
        RECT 98.520 14.920 98.795 14.935 ;
        RECT 98.490 14.645 98.825 14.920 ;
        RECT 99.000 14.895 104.000 15.125 ;
        RECT 104.210 14.935 104.465 14.960 ;
        RECT 98.520 14.630 98.775 14.645 ;
        RECT 99.000 14.455 104.000 14.685 ;
        RECT 104.205 14.645 104.465 14.935 ;
        RECT 104.210 14.630 104.465 14.645 ;
        RECT 99.045 14.445 103.900 14.455 ;
        RECT 99.045 12.920 101.690 12.925 ;
        RECT 97.720 12.720 101.690 12.920 ;
        RECT 97.720 12.690 101.680 12.720 ;
        RECT 96.560 12.335 96.895 12.610 ;
        RECT 97.440 12.440 97.670 12.485 ;
        RECT 92.420 8.560 92.775 8.580 ;
        RECT 92.420 8.490 92.650 8.560 ;
        RECT 93.560 8.490 93.790 8.580 ;
        RECT 94.320 8.465 95.230 8.605 ;
        RECT 95.850 8.490 96.240 8.625 ;
        RECT 94.310 8.285 95.320 8.465 ;
        RECT 90.410 8.055 92.370 8.285 ;
        RECT 93.840 8.055 95.800 8.285 ;
        RECT 91.095 6.975 91.495 8.055 ;
        RECT 93.865 8.050 95.750 8.055 ;
        RECT 96.045 6.355 96.240 8.490 ;
        RECT 96.630 6.830 96.820 12.335 ;
        RECT 97.250 11.105 97.670 12.440 ;
        RECT 98.975 11.105 100.320 12.690 ;
        RECT 97.250 9.720 100.320 11.105 ;
        RECT 97.250 8.990 97.670 9.720 ;
        RECT 97.245 8.485 97.670 8.990 ;
        RECT 96.630 6.640 96.945 6.830 ;
        RECT 86.950 6.125 90.910 6.355 ;
        RECT 92.380 6.125 96.340 6.355 ;
        RECT 96.755 6.130 96.945 6.640 ;
        RECT 86.670 5.515 86.900 5.965 ;
        RECT 88.150 5.515 88.940 6.125 ;
        RECT 86.670 5.210 88.940 5.515 ;
        RECT 86.615 5.195 88.940 5.210 ;
        RECT 86.530 4.350 88.940 5.195 ;
        RECT 86.530 3.975 86.900 4.350 ;
        RECT 86.670 3.965 86.900 3.975 ;
        RECT 88.150 3.805 88.940 4.350 ;
        RECT 90.960 5.880 91.190 5.965 ;
        RECT 92.100 5.880 92.330 5.965 ;
        RECT 90.960 4.055 92.330 5.880 ;
        RECT 90.960 3.965 91.190 4.055 ;
        RECT 86.950 3.575 90.910 3.805 ;
        RECT 83.890 3.255 86.085 3.280 ;
        RECT 86.530 3.255 86.755 3.265 ;
        RECT 91.430 3.255 91.920 4.055 ;
        RECT 92.100 3.965 92.330 4.055 ;
        RECT 93.815 5.745 95.155 6.125 ;
        RECT 96.390 5.745 96.620 5.965 ;
        RECT 93.815 4.150 96.620 5.745 ;
        RECT 93.815 3.805 95.155 4.150 ;
        RECT 96.390 3.965 96.620 4.150 ;
        RECT 92.380 3.575 96.340 3.805 ;
        RECT 96.770 3.785 96.945 6.130 ;
        RECT 97.245 5.965 97.540 8.485 ;
        RECT 98.975 8.280 100.320 9.720 ;
        RECT 101.730 12.390 101.960 12.485 ;
        RECT 102.205 12.390 102.695 14.445 ;
        RECT 103.265 12.920 103.900 12.925 ;
        RECT 103.150 12.690 107.110 12.920 ;
        RECT 102.870 12.390 103.100 12.485 ;
        RECT 101.730 8.565 103.100 12.390 ;
        RECT 101.730 8.485 101.960 8.565 ;
        RECT 102.870 8.485 103.100 8.565 ;
        RECT 104.525 8.280 105.870 12.690 ;
        RECT 107.160 12.420 107.390 12.485 ;
        RECT 108.045 12.425 108.520 17.260 ;
        RECT 109.845 16.455 110.525 17.260 ;
        RECT 110.945 16.735 111.280 16.985 ;
        RECT 110.960 16.710 111.250 16.735 ;
        RECT 114.420 16.635 116.330 17.260 ;
        RECT 118.420 16.925 120.305 16.930 ;
        RECT 121.865 16.925 123.750 16.930 ;
        RECT 118.410 16.695 120.370 16.925 ;
        RECT 121.840 16.695 123.800 16.925 ;
        RECT 110.770 16.455 111.000 16.505 ;
        RECT 109.845 15.955 111.000 16.455 ;
        RECT 108.915 12.735 109.250 12.985 ;
        RECT 108.935 12.705 109.225 12.735 ;
        RECT 108.745 12.425 108.975 12.500 ;
        RECT 107.160 8.485 107.615 12.420 ;
        RECT 108.045 11.680 108.975 12.425 ;
        RECT 108.380 8.565 108.975 11.680 ;
        RECT 108.745 8.500 108.975 8.565 ;
        RECT 109.185 12.475 109.415 12.500 ;
        RECT 109.185 8.920 109.695 12.475 ;
        RECT 109.185 8.550 109.880 8.920 ;
        RECT 110.380 8.600 111.000 15.955 ;
        RECT 109.185 8.500 109.415 8.550 ;
        RECT 97.720 8.250 101.680 8.280 ;
        RECT 103.150 8.250 107.110 8.280 ;
        RECT 97.720 8.090 107.110 8.250 ;
        RECT 97.720 8.050 101.680 8.090 ;
        RECT 103.150 8.050 107.110 8.090 ;
        RECT 107.275 6.660 107.615 8.485 ;
        RECT 108.925 6.660 109.345 8.305 ;
        RECT 107.275 6.505 109.345 6.660 ;
        RECT 107.350 6.390 109.345 6.505 ;
        RECT 97.810 6.125 101.770 6.355 ;
        RECT 103.240 6.125 107.200 6.355 ;
        RECT 97.245 5.205 97.760 5.965 ;
        RECT 97.315 4.025 97.760 5.205 ;
        RECT 97.530 3.965 97.760 4.025 ;
        RECT 99.190 3.805 100.145 6.125 ;
        RECT 101.820 5.900 102.050 5.965 ;
        RECT 102.960 5.900 103.190 5.965 ;
        RECT 101.820 4.030 103.190 5.900 ;
        RECT 101.820 3.965 102.050 4.030 ;
        RECT 96.755 3.255 96.945 3.785 ;
        RECT 97.810 3.575 101.770 3.805 ;
        RECT 102.225 3.255 102.780 4.030 ;
        RECT 102.960 3.965 103.190 4.030 ;
        RECT 104.635 3.805 105.590 6.125 ;
        RECT 107.350 5.970 107.615 6.390 ;
        RECT 108.925 6.115 109.345 6.390 ;
        RECT 109.580 7.355 109.880 8.550 ;
        RECT 110.770 8.505 111.000 8.600 ;
        RECT 111.210 16.430 111.440 16.505 ;
        RECT 111.210 9.110 111.985 16.430 ;
        RECT 114.385 16.405 116.385 16.635 ;
        RECT 118.130 16.410 118.360 16.490 ;
        RECT 113.950 13.060 114.180 16.355 ;
        RECT 116.590 16.275 116.820 16.355 ;
        RECT 116.560 13.060 116.820 16.275 ;
        RECT 113.950 11.245 116.820 13.060 ;
        RECT 111.210 8.580 112.060 9.110 ;
        RECT 113.950 8.825 114.180 11.245 ;
        RECT 111.210 8.505 111.440 8.580 ;
        RECT 110.875 7.825 111.390 8.315 ;
        RECT 110.875 7.360 111.385 7.825 ;
        RECT 111.690 7.795 112.060 8.580 ;
        RECT 113.590 8.395 114.180 8.825 ;
        RECT 115.075 8.640 115.335 8.960 ;
        RECT 116.560 8.645 116.820 11.245 ;
        RECT 117.890 8.990 118.360 16.410 ;
        RECT 118.850 9.775 119.740 16.695 ;
        RECT 120.420 16.390 120.650 16.490 ;
        RECT 120.420 16.380 120.775 16.390 ;
        RECT 121.560 16.380 121.790 16.490 ;
        RECT 115.130 8.480 115.280 8.640 ;
        RECT 110.510 7.355 111.385 7.360 ;
        RECT 109.580 6.950 111.385 7.355 ;
        RECT 109.580 6.110 109.880 6.950 ;
        RECT 110.510 6.935 111.385 6.950 ;
        RECT 110.875 6.825 111.385 6.935 ;
        RECT 110.875 6.125 111.390 6.825 ;
        RECT 111.615 6.795 112.645 7.795 ;
        RECT 107.275 5.965 107.615 5.970 ;
        RECT 107.250 4.020 107.615 5.965 ;
        RECT 108.830 5.900 109.060 5.970 ;
        RECT 108.335 5.230 109.060 5.900 ;
        RECT 108.325 5.040 109.060 5.230 ;
        RECT 108.325 4.240 108.680 5.040 ;
        RECT 108.830 4.970 109.060 5.040 ;
        RECT 109.270 5.925 109.500 5.970 ;
        RECT 109.640 5.925 109.880 6.110 ;
        RECT 109.270 5.595 109.880 5.925 ;
        RECT 110.855 5.870 111.085 5.975 ;
        RECT 109.270 5.040 109.765 5.595 ;
        RECT 109.270 4.970 109.500 5.040 ;
        RECT 109.020 4.785 109.310 4.810 ;
        RECT 109.005 4.535 109.340 4.785 ;
        RECT 110.625 4.765 111.085 5.870 ;
        RECT 110.305 4.240 111.085 4.765 ;
        RECT 107.885 4.060 111.085 4.240 ;
        RECT 107.250 3.965 107.480 4.020 ;
        RECT 103.240 3.575 107.200 3.805 ;
        RECT 107.885 3.620 110.690 4.060 ;
        RECT 110.855 3.975 111.085 4.060 ;
        RECT 111.295 5.910 111.525 5.975 ;
        RECT 111.690 5.910 112.060 6.795 ;
        RECT 111.295 5.585 112.060 5.910 ;
        RECT 111.295 4.045 112.055 5.585 ;
        RECT 111.295 3.975 111.525 4.045 ;
        RECT 111.045 3.795 111.335 3.815 ;
        RECT 107.885 3.255 110.350 3.620 ;
        RECT 111.020 3.545 111.355 3.795 ;
        RECT 113.590 3.280 114.085 8.395 ;
        RECT 115.105 8.345 115.310 8.480 ;
        RECT 116.590 8.395 116.820 8.645 ;
        RECT 117.610 8.550 118.360 8.990 ;
        RECT 118.780 8.775 119.795 9.775 ;
        RECT 114.385 8.115 116.385 8.345 ;
        RECT 117.610 6.355 117.980 8.550 ;
        RECT 118.130 8.490 118.360 8.550 ;
        RECT 118.850 8.285 119.740 8.775 ;
        RECT 120.420 8.580 121.790 16.380 ;
        RECT 122.325 11.635 123.215 16.695 ;
        RECT 123.850 16.410 124.080 16.490 ;
        RECT 122.320 10.015 123.220 11.635 ;
        RECT 122.325 9.605 123.215 10.015 ;
        RECT 122.250 8.605 123.280 9.605 ;
        RECT 123.850 8.625 124.225 16.410 ;
        RECT 124.500 16.025 126.180 17.260 ;
        RECT 127.015 16.025 131.940 16.035 ;
        RECT 124.500 15.545 131.940 16.025 ;
        RECT 124.500 13.285 126.180 15.545 ;
        RECT 127.015 15.125 131.940 15.545 ;
        RECT 126.520 14.935 126.775 14.960 ;
        RECT 126.520 14.920 126.795 14.935 ;
        RECT 126.490 14.645 126.825 14.920 ;
        RECT 127.000 14.895 132.000 15.125 ;
        RECT 132.210 14.935 132.465 14.960 ;
        RECT 126.520 14.630 126.775 14.645 ;
        RECT 127.000 14.455 132.000 14.685 ;
        RECT 132.205 14.645 132.465 14.935 ;
        RECT 132.210 14.630 132.465 14.645 ;
        RECT 127.045 14.445 131.900 14.455 ;
        RECT 127.045 12.920 129.690 12.925 ;
        RECT 125.720 12.720 129.690 12.920 ;
        RECT 125.720 12.690 129.680 12.720 ;
        RECT 124.560 12.335 124.895 12.610 ;
        RECT 125.440 12.440 125.670 12.485 ;
        RECT 120.420 8.560 120.775 8.580 ;
        RECT 120.420 8.490 120.650 8.560 ;
        RECT 121.560 8.490 121.790 8.580 ;
        RECT 122.320 8.465 123.230 8.605 ;
        RECT 123.850 8.490 124.240 8.625 ;
        RECT 122.310 8.285 123.320 8.465 ;
        RECT 118.410 8.055 120.370 8.285 ;
        RECT 121.840 8.055 123.800 8.285 ;
        RECT 119.150 7.155 119.435 8.055 ;
        RECT 121.865 8.050 123.750 8.055 ;
        RECT 124.045 6.355 124.240 8.490 ;
        RECT 124.630 6.830 124.820 12.335 ;
        RECT 125.250 11.105 125.670 12.440 ;
        RECT 126.975 11.105 128.320 12.690 ;
        RECT 125.250 9.720 128.320 11.105 ;
        RECT 125.250 8.990 125.670 9.720 ;
        RECT 125.245 8.485 125.670 8.990 ;
        RECT 124.630 6.640 124.945 6.830 ;
        RECT 114.950 6.125 118.910 6.355 ;
        RECT 120.380 6.125 124.340 6.355 ;
        RECT 124.755 6.130 124.945 6.640 ;
        RECT 114.670 5.515 114.900 5.965 ;
        RECT 116.150 5.515 116.940 6.125 ;
        RECT 114.670 5.210 116.940 5.515 ;
        RECT 114.615 5.195 116.940 5.210 ;
        RECT 114.530 4.350 116.940 5.195 ;
        RECT 114.530 3.975 114.900 4.350 ;
        RECT 114.670 3.965 114.900 3.975 ;
        RECT 116.150 3.805 116.940 4.350 ;
        RECT 118.960 5.880 119.190 5.965 ;
        RECT 120.100 5.880 120.330 5.965 ;
        RECT 118.960 4.055 120.330 5.880 ;
        RECT 118.960 3.965 119.190 4.055 ;
        RECT 114.950 3.575 118.910 3.805 ;
        RECT 111.590 3.255 114.085 3.280 ;
        RECT 114.530 3.255 114.755 3.265 ;
        RECT 119.430 3.255 119.920 4.055 ;
        RECT 120.100 3.965 120.330 4.055 ;
        RECT 121.815 5.745 123.155 6.125 ;
        RECT 124.390 5.745 124.620 5.965 ;
        RECT 121.815 4.150 124.620 5.745 ;
        RECT 121.815 3.805 123.155 4.150 ;
        RECT 124.390 3.965 124.620 4.150 ;
        RECT 120.380 3.575 124.340 3.805 ;
        RECT 124.770 3.785 124.945 6.130 ;
        RECT 125.245 5.965 125.540 8.485 ;
        RECT 126.975 8.280 128.320 9.720 ;
        RECT 129.730 12.390 129.960 12.485 ;
        RECT 130.205 12.390 130.695 14.445 ;
        RECT 131.265 12.920 131.900 12.925 ;
        RECT 131.150 12.690 135.110 12.920 ;
        RECT 130.870 12.390 131.100 12.485 ;
        RECT 129.730 8.565 131.100 12.390 ;
        RECT 129.730 8.485 129.960 8.565 ;
        RECT 130.870 8.485 131.100 8.565 ;
        RECT 132.525 8.280 133.870 12.690 ;
        RECT 135.160 12.420 135.390 12.485 ;
        RECT 136.045 12.425 136.520 17.260 ;
        RECT 137.845 16.455 138.525 17.260 ;
        RECT 138.945 16.735 139.280 16.985 ;
        RECT 138.960 16.710 139.250 16.735 ;
        RECT 138.770 16.455 139.000 16.505 ;
        RECT 137.845 15.955 139.000 16.455 ;
        RECT 136.915 12.735 137.250 12.985 ;
        RECT 136.935 12.705 137.225 12.735 ;
        RECT 136.745 12.425 136.975 12.500 ;
        RECT 135.160 8.485 135.615 12.420 ;
        RECT 136.045 11.680 136.975 12.425 ;
        RECT 136.380 8.565 136.975 11.680 ;
        RECT 136.745 8.500 136.975 8.565 ;
        RECT 137.185 12.475 137.415 12.500 ;
        RECT 137.185 8.920 137.695 12.475 ;
        RECT 137.185 8.550 137.880 8.920 ;
        RECT 138.380 8.600 139.000 15.955 ;
        RECT 137.185 8.500 137.415 8.550 ;
        RECT 125.720 8.250 129.680 8.280 ;
        RECT 131.150 8.250 135.110 8.280 ;
        RECT 125.720 8.090 135.110 8.250 ;
        RECT 125.720 8.050 129.680 8.090 ;
        RECT 131.150 8.050 135.110 8.090 ;
        RECT 135.275 6.660 135.615 8.485 ;
        RECT 136.925 6.660 137.345 8.305 ;
        RECT 135.275 6.505 137.345 6.660 ;
        RECT 135.350 6.390 137.345 6.505 ;
        RECT 125.810 6.125 129.770 6.355 ;
        RECT 131.240 6.125 135.200 6.355 ;
        RECT 125.245 5.205 125.760 5.965 ;
        RECT 125.315 4.025 125.760 5.205 ;
        RECT 125.530 3.965 125.760 4.025 ;
        RECT 127.190 3.805 128.145 6.125 ;
        RECT 129.820 5.900 130.050 5.965 ;
        RECT 130.960 5.900 131.190 5.965 ;
        RECT 129.820 4.030 131.190 5.900 ;
        RECT 129.820 3.965 130.050 4.030 ;
        RECT 124.755 3.255 124.945 3.785 ;
        RECT 125.810 3.575 129.770 3.805 ;
        RECT 130.225 3.255 130.780 4.030 ;
        RECT 130.960 3.965 131.190 4.030 ;
        RECT 132.635 3.805 133.590 6.125 ;
        RECT 135.350 5.970 135.615 6.390 ;
        RECT 136.925 6.115 137.345 6.390 ;
        RECT 137.580 7.355 137.880 8.550 ;
        RECT 138.770 8.505 139.000 8.600 ;
        RECT 139.210 16.430 139.440 16.505 ;
        RECT 139.210 9.110 139.985 16.430 ;
        RECT 139.210 8.580 140.060 9.110 ;
        RECT 139.210 8.505 139.440 8.580 ;
        RECT 138.875 7.825 139.390 8.315 ;
        RECT 138.875 7.360 139.385 7.825 ;
        RECT 139.690 7.795 140.060 8.580 ;
        RECT 138.510 7.355 139.385 7.360 ;
        RECT 137.580 6.950 139.385 7.355 ;
        RECT 137.580 6.110 137.880 6.950 ;
        RECT 138.510 6.935 139.385 6.950 ;
        RECT 138.875 6.825 139.385 6.935 ;
        RECT 138.875 6.125 139.390 6.825 ;
        RECT 139.615 6.795 140.645 7.795 ;
        RECT 135.275 5.965 135.615 5.970 ;
        RECT 135.250 4.020 135.615 5.965 ;
        RECT 136.830 5.900 137.060 5.970 ;
        RECT 136.335 5.230 137.060 5.900 ;
        RECT 136.325 5.040 137.060 5.230 ;
        RECT 136.325 4.240 136.680 5.040 ;
        RECT 136.830 4.970 137.060 5.040 ;
        RECT 137.270 5.925 137.500 5.970 ;
        RECT 137.640 5.925 137.880 6.110 ;
        RECT 137.270 5.595 137.880 5.925 ;
        RECT 138.855 5.870 139.085 5.975 ;
        RECT 137.270 5.040 137.765 5.595 ;
        RECT 137.270 4.970 137.500 5.040 ;
        RECT 137.020 4.785 137.310 4.810 ;
        RECT 137.005 4.535 137.340 4.785 ;
        RECT 138.625 4.765 139.085 5.870 ;
        RECT 138.305 4.240 139.085 4.765 ;
        RECT 135.885 4.060 139.085 4.240 ;
        RECT 135.250 3.965 135.480 4.020 ;
        RECT 131.240 3.575 135.200 3.805 ;
        RECT 135.885 3.620 138.690 4.060 ;
        RECT 138.855 3.975 139.085 4.060 ;
        RECT 139.295 5.910 139.525 5.975 ;
        RECT 139.690 5.910 140.060 6.795 ;
        RECT 139.295 5.585 140.060 5.910 ;
        RECT 139.295 4.045 140.055 5.585 ;
        RECT 139.295 3.975 139.525 4.045 ;
        RECT 139.045 3.795 139.335 3.815 ;
        RECT 135.885 3.255 138.350 3.620 ;
        RECT 139.020 3.545 139.355 3.795 ;
        RECT 1.475 2.380 140.080 3.255 ;
      LAYER met2 ;
        RECT 22.630 223.160 22.910 223.660 ;
        RECT 32.290 223.160 32.570 223.660 ;
        RECT 35.510 223.160 35.790 223.660 ;
        RECT 38.730 223.160 39.010 223.660 ;
        RECT 41.950 223.160 42.230 223.660 ;
        RECT 45.170 223.160 45.450 223.660 ;
        RECT 48.390 223.160 48.670 223.660 ;
        RECT 51.610 223.160 51.890 223.660 ;
        RECT 54.830 223.160 55.110 223.660 ;
        RECT 58.050 223.160 58.330 223.660 ;
        RECT 61.270 223.160 61.550 223.660 ;
        RECT 22.700 220.590 22.840 223.160 ;
        RECT 22.640 220.270 22.900 220.590 ;
        RECT 16.190 219.735 16.470 220.105 ;
        RECT 15.740 210.410 16.000 210.730 ;
        RECT 15.280 208.030 15.540 208.350 ;
        RECT 10.220 188.990 10.480 189.310 ;
        RECT 10.280 182.705 10.420 188.990 ;
        RECT 10.210 182.335 10.490 182.705 ;
        RECT 11.140 181.170 11.400 181.490 ;
        RECT 9.760 175.390 10.020 175.710 ;
        RECT 9.820 157.310 9.960 175.390 ;
        RECT 11.200 158.905 11.340 181.170 ;
        RECT 12.980 177.770 13.240 178.090 ;
        RECT 11.130 158.535 11.410 158.905 ;
        RECT 13.040 157.310 13.180 177.770 ;
        RECT 15.340 176.730 15.480 208.030 ;
        RECT 15.800 187.610 15.940 210.410 ;
        RECT 16.260 201.550 16.400 219.735 ;
        RECT 24.010 212.935 24.290 213.305 ;
        RECT 20.800 212.110 21.060 212.430 ;
        RECT 18.040 211.430 18.300 211.750 ;
        RECT 17.570 210.895 17.850 211.265 ;
        RECT 17.580 210.750 17.840 210.895 ;
        RECT 18.100 210.585 18.240 211.430 ;
        RECT 19.880 211.090 20.140 211.410 ;
        RECT 20.340 211.090 20.600 211.410 ;
        RECT 18.030 210.215 18.310 210.585 ;
        RECT 17.120 207.690 17.380 208.010 ;
        RECT 18.040 207.690 18.300 208.010 ;
        RECT 16.660 205.990 16.920 206.310 ;
        RECT 16.200 201.230 16.460 201.550 ;
        RECT 16.720 200.870 16.860 205.990 ;
        RECT 16.660 200.550 16.920 200.870 ;
        RECT 17.180 197.810 17.320 207.690 ;
        RECT 18.100 203.250 18.240 207.690 ;
        RECT 18.040 202.930 18.300 203.250 ;
        RECT 18.960 202.930 19.220 203.250 ;
        RECT 19.020 198.830 19.160 202.930 ;
        RECT 19.420 200.550 19.680 200.870 ;
        RECT 18.960 198.510 19.220 198.830 ;
        RECT 16.660 197.490 16.920 197.810 ;
        RECT 17.120 197.490 17.380 197.810 ;
        RECT 17.580 197.490 17.840 197.810 ;
        RECT 16.200 194.430 16.460 194.750 ;
        RECT 16.260 193.390 16.400 194.430 ;
        RECT 16.200 193.070 16.460 193.390 ;
        RECT 16.720 191.430 16.860 197.490 ;
        RECT 17.120 196.810 17.380 197.130 ;
        RECT 17.180 192.370 17.320 196.810 ;
        RECT 17.640 194.945 17.780 197.490 ;
        RECT 17.570 194.575 17.850 194.945 ;
        RECT 17.120 192.050 17.380 192.370 ;
        RECT 17.110 191.430 17.390 191.545 ;
        RECT 16.720 191.290 17.390 191.430 ;
        RECT 17.110 191.175 17.390 191.290 ;
        RECT 17.180 189.230 17.320 191.175 ;
        RECT 17.640 189.900 17.780 194.575 ;
        RECT 18.960 192.730 19.220 193.050 ;
        RECT 18.500 192.225 18.760 192.370 ;
        RECT 18.490 191.855 18.770 192.225 ;
        RECT 17.640 189.760 18.240 189.900 ;
        RECT 17.180 189.090 17.780 189.230 ;
        RECT 15.740 187.290 16.000 187.610 ;
        RECT 17.640 186.930 17.780 189.090 ;
        RECT 17.580 186.610 17.840 186.930 ;
        RECT 18.100 186.590 18.240 189.760 ;
        RECT 19.020 186.930 19.160 192.730 ;
        RECT 19.480 190.330 19.620 200.550 ;
        RECT 19.940 197.130 20.080 211.090 ;
        RECT 20.400 208.690 20.540 211.090 ;
        RECT 20.340 208.370 20.600 208.690 ;
        RECT 20.400 207.865 20.540 208.370 ;
        RECT 20.330 207.495 20.610 207.865 ;
        RECT 20.860 203.930 21.000 212.110 ;
        RECT 24.080 212.090 24.220 212.935 ;
        RECT 23.560 211.770 23.820 212.090 ;
        RECT 24.020 211.770 24.280 212.090 ;
        RECT 21.720 208.710 21.980 209.030 ;
        RECT 20.800 203.610 21.060 203.930 ;
        RECT 21.260 203.270 21.520 203.590 ;
        RECT 20.340 202.590 20.600 202.910 ;
        RECT 20.800 202.590 21.060 202.910 ;
        RECT 20.400 198.830 20.540 202.590 ;
        RECT 20.860 200.530 21.000 202.590 ;
        RECT 20.800 200.210 21.060 200.530 ;
        RECT 20.340 198.510 20.600 198.830 ;
        RECT 19.880 196.810 20.140 197.130 ;
        RECT 19.420 190.010 19.680 190.330 ;
        RECT 19.940 189.230 20.080 196.810 ;
        RECT 19.480 189.090 20.080 189.230 ;
        RECT 18.960 186.610 19.220 186.930 ;
        RECT 18.040 186.270 18.300 186.590 ;
        RECT 19.020 185.230 19.160 186.610 ;
        RECT 18.960 184.910 19.220 185.230 ;
        RECT 17.120 183.210 17.380 183.530 ;
        RECT 16.200 180.490 16.460 180.810 ;
        RECT 15.280 176.410 15.540 176.730 ;
        RECT 16.260 174.350 16.400 180.490 ;
        RECT 16.650 177.575 16.930 177.945 ;
        RECT 16.200 174.030 16.460 174.350 ;
        RECT 16.720 173.670 16.860 177.575 ;
        RECT 17.180 176.050 17.320 183.210 ;
        RECT 17.570 181.655 17.850 182.025 ;
        RECT 17.120 175.730 17.380 176.050 ;
        RECT 16.660 173.350 16.920 173.670 ;
        RECT 16.720 170.270 16.860 173.350 ;
        RECT 17.640 171.630 17.780 181.655 ;
        RECT 18.040 181.170 18.300 181.490 ;
        RECT 18.100 179.790 18.240 181.170 ;
        RECT 18.040 179.470 18.300 179.790 ;
        RECT 18.500 178.790 18.760 179.110 ;
        RECT 18.030 174.855 18.310 175.225 ;
        RECT 18.100 171.630 18.240 174.855 ;
        RECT 17.580 171.310 17.840 171.630 ;
        RECT 18.040 171.310 18.300 171.630 ;
        RECT 18.560 170.270 18.700 178.790 ;
        RECT 18.960 176.750 19.220 177.070 ;
        RECT 19.020 175.430 19.160 176.750 ;
        RECT 19.480 176.050 19.620 189.090 ;
        RECT 20.400 187.950 20.540 198.510 ;
        RECT 20.340 187.630 20.600 187.950 ;
        RECT 20.330 187.095 20.610 187.465 ;
        RECT 20.400 186.930 20.540 187.095 ;
        RECT 20.340 186.610 20.600 186.930 ;
        RECT 20.860 186.590 21.000 200.210 ;
        RECT 21.320 192.370 21.460 203.270 ;
        RECT 21.780 193.390 21.920 208.710 ;
        RECT 23.100 208.030 23.360 208.350 ;
        RECT 22.180 207.690 22.440 208.010 ;
        RECT 22.240 198.490 22.380 207.690 ;
        RECT 23.160 205.290 23.300 208.030 ;
        RECT 23.100 204.970 23.360 205.290 ;
        RECT 22.640 198.510 22.900 198.830 ;
        RECT 22.180 198.170 22.440 198.490 ;
        RECT 21.720 193.070 21.980 193.390 ;
        RECT 21.260 192.050 21.520 192.370 ;
        RECT 21.260 190.010 21.520 190.330 ;
        RECT 20.800 186.270 21.060 186.590 ;
        RECT 20.860 183.530 21.000 186.270 ;
        RECT 20.800 183.210 21.060 183.530 ;
        RECT 20.800 181.170 21.060 181.490 ;
        RECT 19.880 178.790 20.140 179.110 ;
        RECT 19.420 175.730 19.680 176.050 ;
        RECT 19.020 175.290 19.620 175.430 ;
        RECT 18.960 173.350 19.220 173.670 ;
        RECT 19.020 171.290 19.160 173.350 ;
        RECT 18.960 170.970 19.220 171.290 ;
        RECT 16.660 169.950 16.920 170.270 ;
        RECT 18.500 169.950 18.760 170.270 ;
        RECT 19.020 168.910 19.160 170.970 ;
        RECT 18.960 168.590 19.220 168.910 ;
        RECT 16.260 157.350 16.860 157.430 ;
        RECT 16.260 157.310 16.920 157.350 ;
        RECT 19.480 157.310 19.620 175.290 ;
        RECT 19.940 174.350 20.080 178.790 ;
        RECT 20.340 178.450 20.600 178.770 ;
        RECT 19.880 174.030 20.140 174.350 ;
        RECT 20.400 171.290 20.540 178.450 ;
        RECT 20.860 176.730 21.000 181.170 ;
        RECT 21.320 179.450 21.460 190.010 ;
        RECT 21.720 188.650 21.980 188.970 ;
        RECT 21.780 186.930 21.920 188.650 ;
        RECT 21.720 186.610 21.980 186.930 ;
        RECT 21.260 179.130 21.520 179.450 ;
        RECT 21.710 178.935 21.990 179.305 ;
        RECT 22.240 179.020 22.380 198.170 ;
        RECT 22.700 192.710 22.840 198.510 ;
        RECT 23.620 198.150 23.760 211.770 ;
        RECT 30.920 211.430 31.180 211.750 ;
        RECT 29.080 208.370 29.340 208.690 ;
        RECT 28.620 206.670 28.880 206.990 ;
        RECT 25.400 205.990 25.660 206.310 ;
        RECT 25.460 203.250 25.600 205.990 ;
        RECT 26.320 205.650 26.580 205.970 ;
        RECT 26.380 203.250 26.520 205.650 ;
        RECT 27.700 204.970 27.960 205.290 ;
        RECT 25.400 202.930 25.660 203.250 ;
        RECT 26.320 202.930 26.580 203.250 ;
        RECT 25.400 202.250 25.660 202.570 ;
        RECT 25.460 199.850 25.600 202.250 ;
        RECT 25.400 199.530 25.660 199.850 ;
        RECT 23.560 197.830 23.820 198.150 ;
        RECT 23.100 197.490 23.360 197.810 ;
        RECT 22.640 192.390 22.900 192.710 ;
        RECT 23.160 192.030 23.300 197.490 ;
        RECT 22.640 191.710 22.900 192.030 ;
        RECT 23.100 191.710 23.360 192.030 ;
        RECT 22.700 188.825 22.840 191.710 ;
        RECT 23.160 190.670 23.300 191.710 ;
        RECT 23.100 190.350 23.360 190.670 ;
        RECT 23.620 190.070 23.760 197.830 ;
        RECT 24.020 197.665 24.280 197.810 ;
        RECT 24.010 197.295 24.290 197.665 ;
        RECT 24.080 197.130 24.220 197.295 ;
        RECT 24.020 196.810 24.280 197.130 ;
        RECT 24.480 195.110 24.740 195.430 ;
        RECT 24.940 195.110 25.200 195.430 ;
        RECT 24.020 194.430 24.280 194.750 ;
        RECT 24.080 193.390 24.220 194.430 ;
        RECT 24.020 193.070 24.280 193.390 ;
        RECT 24.540 192.710 24.680 195.110 ;
        RECT 24.020 192.390 24.280 192.710 ;
        RECT 24.480 192.390 24.740 192.710 ;
        RECT 23.160 189.930 23.760 190.070 ;
        RECT 22.630 188.455 22.910 188.825 ;
        RECT 22.640 181.345 22.900 181.490 ;
        RECT 22.630 180.975 22.910 181.345 ;
        RECT 22.640 179.020 22.900 179.110 ;
        RECT 21.720 178.790 21.980 178.935 ;
        RECT 22.240 178.880 22.900 179.020 ;
        RECT 22.640 178.790 22.900 178.880 ;
        RECT 20.800 176.410 21.060 176.730 ;
        RECT 21.780 171.630 21.920 178.790 ;
        RECT 23.160 177.070 23.300 189.930 ;
        RECT 24.080 183.385 24.220 192.390 ;
        RECT 25.000 187.610 25.140 195.110 ;
        RECT 25.460 192.370 25.600 199.530 ;
        RECT 25.860 197.490 26.120 197.810 ;
        RECT 26.320 197.490 26.580 197.810 ;
        RECT 25.400 192.050 25.660 192.370 ;
        RECT 24.940 187.290 25.200 187.610 ;
        RECT 24.940 186.610 25.200 186.930 ;
        RECT 24.480 185.930 24.740 186.250 ;
        RECT 24.010 183.015 24.290 183.385 ;
        RECT 23.560 181.170 23.820 181.490 ;
        RECT 23.620 177.070 23.760 181.170 ;
        RECT 24.080 181.150 24.220 183.015 ;
        RECT 24.540 181.490 24.680 185.930 ;
        RECT 24.480 181.170 24.740 181.490 ;
        RECT 24.020 180.830 24.280 181.150 ;
        RECT 23.100 176.750 23.360 177.070 ;
        RECT 23.560 176.750 23.820 177.070 ;
        RECT 22.640 172.330 22.900 172.650 ;
        RECT 24.480 172.330 24.740 172.650 ;
        RECT 21.720 171.310 21.980 171.630 ;
        RECT 20.340 170.970 20.600 171.290 ;
        RECT 20.340 170.465 20.600 170.610 ;
        RECT 19.880 169.950 20.140 170.270 ;
        RECT 20.330 170.095 20.610 170.465 ;
        RECT 19.940 169.785 20.080 169.950 ;
        RECT 19.870 169.415 20.150 169.785 ;
        RECT 22.700 157.310 22.840 172.330 ;
        RECT 23.090 171.455 23.370 171.825 ;
        RECT 23.160 170.610 23.300 171.455 ;
        RECT 23.100 170.290 23.360 170.610 ;
        RECT 24.540 168.910 24.680 172.330 ;
        RECT 25.000 171.630 25.140 186.610 ;
        RECT 25.920 182.025 26.060 197.490 ;
        RECT 26.380 190.330 26.520 197.490 ;
        RECT 26.780 196.810 27.040 197.130 ;
        RECT 26.320 190.010 26.580 190.330 ;
        RECT 26.840 189.990 26.980 196.810 ;
        RECT 27.240 192.050 27.500 192.370 ;
        RECT 26.780 189.670 27.040 189.990 ;
        RECT 26.320 187.630 26.580 187.950 ;
        RECT 25.850 181.655 26.130 182.025 ;
        RECT 25.920 181.150 26.060 181.655 ;
        RECT 25.860 180.830 26.120 181.150 ;
        RECT 25.400 180.490 25.660 180.810 ;
        RECT 25.460 179.790 25.600 180.490 ;
        RECT 25.400 179.470 25.660 179.790 ;
        RECT 25.860 176.070 26.120 176.390 ;
        RECT 25.400 173.920 25.660 174.010 ;
        RECT 25.920 173.920 26.060 176.070 ;
        RECT 25.400 173.780 26.060 173.920 ;
        RECT 25.400 173.690 25.660 173.780 ;
        RECT 25.920 171.630 26.060 173.780 ;
        RECT 26.380 173.670 26.520 187.630 ;
        RECT 26.780 186.270 27.040 186.590 ;
        RECT 26.840 185.230 26.980 186.270 ;
        RECT 26.780 184.910 27.040 185.230 ;
        RECT 26.840 184.120 26.980 184.910 ;
        RECT 27.300 184.890 27.440 192.050 ;
        RECT 27.760 190.185 27.900 204.970 ;
        RECT 28.160 203.270 28.420 203.590 ;
        RECT 28.220 197.470 28.360 203.270 ;
        RECT 28.680 199.850 28.820 206.670 ;
        RECT 29.140 203.590 29.280 208.370 ;
        RECT 29.540 206.670 29.800 206.990 ;
        RECT 29.600 203.930 29.740 206.670 ;
        RECT 30.980 204.270 31.120 211.430 ;
        RECT 32.360 211.410 32.500 223.160 ;
        RECT 35.520 222.990 35.780 223.160 ;
        RECT 38.800 217.190 38.940 223.160 ;
        RECT 42.020 218.210 42.160 223.160 ;
        RECT 41.960 217.890 42.220 218.210 ;
        RECT 45.240 217.530 45.380 223.160 ;
        RECT 48.460 218.550 48.600 223.160 ;
        RECT 48.400 218.230 48.660 218.550 ;
        RECT 51.680 217.870 51.820 223.160 ;
        RECT 54.900 218.890 55.040 223.160 ;
        RECT 54.840 218.570 55.100 218.890 ;
        RECT 51.620 217.550 51.880 217.870 ;
        RECT 45.180 217.210 45.440 217.530 ;
        RECT 38.740 216.870 39.000 217.190 ;
        RECT 54.840 215.510 55.100 215.830 ;
        RECT 34.140 214.830 34.400 215.150 ;
        RECT 33.680 213.810 33.940 214.130 ;
        RECT 33.740 212.090 33.880 213.810 ;
        RECT 33.680 211.770 33.940 212.090 ;
        RECT 32.300 211.090 32.560 211.410 ;
        RECT 32.760 211.090 33.020 211.410 ;
        RECT 34.200 211.320 34.340 214.830 ;
        RECT 48.860 214.490 49.120 214.810 ;
        RECT 48.400 213.130 48.660 213.450 ;
        RECT 34.600 212.110 34.860 212.430 ;
        RECT 33.740 211.180 34.340 211.320 ;
        RECT 32.300 208.030 32.560 208.350 ;
        RECT 31.840 205.650 32.100 205.970 ;
        RECT 31.900 205.290 32.040 205.650 ;
        RECT 31.380 204.970 31.640 205.290 ;
        RECT 31.840 204.970 32.100 205.290 ;
        RECT 30.920 203.950 31.180 204.270 ;
        RECT 29.540 203.840 29.800 203.930 ;
        RECT 29.540 203.700 30.200 203.840 ;
        RECT 29.540 203.610 29.800 203.700 ;
        RECT 29.080 203.270 29.340 203.590 ;
        RECT 28.620 199.530 28.880 199.850 ;
        RECT 28.620 197.830 28.880 198.150 ;
        RECT 28.160 197.150 28.420 197.470 ;
        RECT 28.680 196.870 28.820 197.830 ;
        RECT 28.220 196.730 28.820 196.870 ;
        RECT 28.220 190.865 28.360 196.730 ;
        RECT 29.140 195.090 29.280 203.270 ;
        RECT 29.540 200.550 29.800 200.870 ;
        RECT 29.080 194.770 29.340 195.090 ;
        RECT 29.600 194.410 29.740 200.550 ;
        RECT 29.540 194.090 29.800 194.410 ;
        RECT 28.150 190.495 28.430 190.865 ;
        RECT 27.690 189.815 27.970 190.185 ;
        RECT 27.700 186.840 27.960 186.930 ;
        RECT 28.220 186.840 28.360 190.495 ;
        RECT 28.620 190.350 28.880 190.670 ;
        RECT 28.680 187.950 28.820 190.350 ;
        RECT 28.620 187.630 28.880 187.950 ;
        RECT 27.700 186.700 28.360 186.840 ;
        RECT 28.620 186.840 28.880 186.930 ;
        RECT 28.620 186.700 29.280 186.840 ;
        RECT 27.700 186.610 27.960 186.700 ;
        RECT 28.620 186.610 28.880 186.700 ;
        RECT 28.620 185.930 28.880 186.250 ;
        RECT 27.240 184.570 27.500 184.890 ;
        RECT 28.680 184.210 28.820 185.930 ;
        RECT 29.140 184.745 29.280 186.700 ;
        RECT 29.070 184.375 29.350 184.745 ;
        RECT 29.600 184.550 29.740 194.090 ;
        RECT 30.060 187.950 30.200 203.700 ;
        RECT 31.440 197.470 31.580 204.970 ;
        RECT 31.380 197.150 31.640 197.470 ;
        RECT 31.440 192.030 31.580 197.150 ;
        RECT 32.360 192.030 32.500 208.030 ;
        RECT 32.820 206.650 32.960 211.090 ;
        RECT 33.740 209.710 33.880 211.180 ;
        RECT 33.680 209.390 33.940 209.710 ;
        RECT 34.140 209.390 34.400 209.710 ;
        RECT 32.760 206.330 33.020 206.650 ;
        RECT 34.200 204.350 34.340 209.390 ;
        RECT 34.660 206.990 34.800 212.110 ;
        RECT 46.100 211.770 46.360 212.090 ;
        RECT 46.560 211.770 46.820 212.090 ;
        RECT 37.360 211.430 37.620 211.750 ;
        RECT 39.660 211.430 39.920 211.750 ;
        RECT 40.120 211.430 40.380 211.750 ;
        RECT 42.880 211.430 43.140 211.750 ;
        RECT 35.520 211.090 35.780 211.410 ;
        RECT 35.060 210.750 35.320 211.070 ;
        RECT 34.600 206.670 34.860 206.990 ;
        RECT 33.740 204.210 34.340 204.350 ;
        RECT 33.740 202.910 33.880 204.210 ;
        RECT 34.140 203.840 34.400 203.930 ;
        RECT 35.120 203.840 35.260 210.750 ;
        RECT 35.580 209.370 35.720 211.090 ;
        RECT 35.980 210.410 36.240 210.730 ;
        RECT 35.520 209.050 35.780 209.370 ;
        RECT 36.040 208.690 36.180 210.410 ;
        RECT 35.980 208.370 36.240 208.690 ;
        RECT 37.420 208.350 37.560 211.430 ;
        RECT 39.720 209.030 39.860 211.430 ;
        RECT 39.660 208.710 39.920 209.030 ;
        RECT 37.360 208.030 37.620 208.350 ;
        RECT 35.980 207.690 36.240 208.010 ;
        RECT 35.520 205.990 35.780 206.310 ;
        RECT 34.140 203.700 35.260 203.840 ;
        RECT 34.140 203.610 34.400 203.700 ;
        RECT 33.680 202.590 33.940 202.910 ;
        RECT 34.200 192.370 34.340 203.610 ;
        RECT 34.600 194.090 34.860 194.410 ;
        RECT 31.380 191.710 31.640 192.030 ;
        RECT 32.300 191.710 32.560 192.030 ;
        RECT 32.750 191.855 33.030 192.225 ;
        RECT 34.140 192.050 34.400 192.370 ;
        RECT 30.000 187.630 30.260 187.950 ;
        RECT 26.840 183.980 27.440 184.120 ;
        RECT 27.300 181.490 27.440 183.980 ;
        RECT 28.620 183.890 28.880 184.210 ;
        RECT 27.240 181.170 27.500 181.490 ;
        RECT 26.780 180.490 27.040 180.810 ;
        RECT 26.840 174.010 26.980 180.490 ;
        RECT 27.300 178.430 27.440 181.170 ;
        RECT 27.700 180.830 27.960 181.150 ;
        RECT 27.760 180.665 27.900 180.830 ;
        RECT 27.690 180.295 27.970 180.665 ;
        RECT 27.240 178.110 27.500 178.430 ;
        RECT 28.680 178.090 28.820 183.890 ;
        RECT 29.140 183.870 29.280 184.375 ;
        RECT 29.540 184.230 29.800 184.550 ;
        RECT 29.080 183.550 29.340 183.870 ;
        RECT 30.460 181.170 30.720 181.490 ;
        RECT 31.380 181.170 31.640 181.490 ;
        RECT 28.620 177.770 28.880 178.090 ;
        RECT 28.680 176.050 28.820 177.770 ;
        RECT 28.620 175.730 28.880 176.050 ;
        RECT 26.780 173.690 27.040 174.010 ;
        RECT 30.520 173.865 30.660 181.170 ;
        RECT 30.920 179.470 31.180 179.790 ;
        RECT 26.320 173.350 26.580 173.670 ;
        RECT 30.450 173.495 30.730 173.865 ;
        RECT 29.080 173.010 29.340 173.330 ;
        RECT 29.140 171.630 29.280 173.010 ;
        RECT 24.940 171.310 25.200 171.630 ;
        RECT 25.860 171.310 26.120 171.630 ;
        RECT 29.080 171.310 29.340 171.630 ;
        RECT 26.310 170.775 26.590 171.145 ;
        RECT 26.320 170.630 26.580 170.775 ;
        RECT 24.940 170.290 25.200 170.610 ;
        RECT 26.780 170.290 27.040 170.610 ;
        RECT 28.160 170.290 28.420 170.610 ;
        RECT 25.000 168.910 25.140 170.290 ;
        RECT 24.480 168.590 24.740 168.910 ;
        RECT 24.940 168.590 25.200 168.910 ;
        RECT 25.850 168.055 26.130 168.425 ;
        RECT 25.920 157.310 26.060 168.055 ;
        RECT 26.840 163.665 26.980 170.290 ;
        RECT 28.220 164.345 28.360 170.290 ;
        RECT 29.080 168.250 29.340 168.570 ;
        RECT 28.150 163.975 28.430 164.345 ;
        RECT 26.770 163.295 27.050 163.665 ;
        RECT 29.140 157.310 29.280 168.250 ;
        RECT 9.750 156.810 10.030 157.310 ;
        RECT 12.970 156.810 13.250 157.310 ;
        RECT 16.190 157.290 16.920 157.310 ;
        RECT 16.190 156.810 16.470 157.290 ;
        RECT 16.660 157.030 16.920 157.290 ;
        RECT 19.410 156.810 19.690 157.310 ;
        RECT 22.630 156.810 22.910 157.310 ;
        RECT 25.850 156.810 26.130 157.310 ;
        RECT 29.070 156.810 29.350 157.310 ;
        RECT 30.980 157.130 31.120 179.470 ;
        RECT 31.440 176.050 31.580 181.170 ;
        RECT 31.380 175.730 31.640 176.050 ;
        RECT 31.440 174.350 31.580 175.730 ;
        RECT 31.380 174.030 31.640 174.350 ;
        RECT 32.360 174.010 32.500 191.710 ;
        RECT 32.820 179.450 32.960 191.855 ;
        RECT 34.660 188.970 34.800 194.090 ;
        RECT 35.060 189.330 35.320 189.650 ;
        RECT 34.600 188.650 34.860 188.970 ;
        RECT 33.680 186.610 33.940 186.930 ;
        RECT 33.740 186.250 33.880 186.610 ;
        RECT 33.680 185.930 33.940 186.250 ;
        RECT 34.130 185.055 34.410 185.425 ;
        RECT 33.210 184.375 33.490 184.745 ;
        RECT 33.280 181.830 33.420 184.375 ;
        RECT 33.220 181.510 33.480 181.830 ;
        RECT 33.680 181.345 33.940 181.490 ;
        RECT 33.670 180.975 33.950 181.345 ;
        RECT 32.760 179.130 33.020 179.450 ;
        RECT 33.220 179.130 33.480 179.450 ;
        RECT 32.300 173.690 32.560 174.010 ;
        RECT 33.280 172.505 33.420 179.130 ;
        RECT 34.200 179.110 34.340 185.055 ;
        RECT 34.600 183.550 34.860 183.870 ;
        RECT 34.140 178.790 34.400 179.110 ;
        RECT 33.680 177.770 33.940 178.090 ;
        RECT 33.210 172.135 33.490 172.505 ;
        RECT 33.740 170.610 33.880 177.770 ;
        RECT 34.660 173.670 34.800 183.550 ;
        RECT 35.120 179.110 35.260 189.330 ;
        RECT 35.580 184.890 35.720 205.990 ;
        RECT 36.040 201.210 36.180 207.690 ;
        RECT 37.420 206.990 37.560 208.030 ;
        RECT 37.360 206.670 37.620 206.990 ;
        RECT 37.360 205.990 37.620 206.310 ;
        RECT 36.890 204.095 37.170 204.465 ;
        RECT 36.440 202.930 36.700 203.250 ;
        RECT 35.980 200.890 36.240 201.210 ;
        RECT 35.980 198.510 36.240 198.830 ;
        RECT 36.040 190.330 36.180 198.510 ;
        RECT 36.500 192.710 36.640 202.930 ;
        RECT 36.440 192.390 36.700 192.710 ;
        RECT 36.960 190.670 37.100 204.095 ;
        RECT 37.420 198.830 37.560 205.990 ;
        RECT 39.720 203.590 39.860 208.710 ;
        RECT 40.180 208.010 40.320 211.430 ;
        RECT 42.940 211.070 43.080 211.430 ;
        RECT 42.880 210.750 43.140 211.070 ;
        RECT 46.160 210.730 46.300 211.770 ;
        RECT 46.100 210.410 46.360 210.730 ;
        RECT 45.180 209.390 45.440 209.710 ;
        RECT 40.120 207.690 40.380 208.010 ;
        RECT 41.030 207.495 41.310 207.865 ;
        RECT 39.660 203.270 39.920 203.590 ;
        RECT 40.120 203.270 40.380 203.590 ;
        RECT 39.720 200.190 39.860 203.270 ;
        RECT 39.660 199.870 39.920 200.190 ;
        RECT 37.360 198.510 37.620 198.830 ;
        RECT 37.810 198.655 38.090 199.025 ;
        RECT 37.880 197.810 38.020 198.655 ;
        RECT 40.180 197.810 40.320 203.270 ;
        RECT 37.820 197.490 38.080 197.810 ;
        RECT 40.120 197.490 40.380 197.810 ;
        RECT 41.100 195.770 41.240 207.495 ;
        RECT 44.260 206.670 44.520 206.990 ;
        RECT 43.340 205.650 43.600 205.970 ;
        RECT 41.950 203.415 42.230 203.785 ;
        RECT 41.500 197.830 41.760 198.150 ;
        RECT 41.560 196.985 41.700 197.830 ;
        RECT 41.490 196.615 41.770 196.985 ;
        RECT 41.040 195.450 41.300 195.770 ;
        RECT 37.820 195.110 38.080 195.430 ;
        RECT 37.360 194.770 37.620 195.090 ;
        RECT 36.900 190.580 37.160 190.670 ;
        RECT 36.500 190.440 37.160 190.580 ;
        RECT 35.980 190.010 36.240 190.330 ;
        RECT 36.500 189.990 36.640 190.440 ;
        RECT 36.900 190.350 37.160 190.440 ;
        RECT 36.440 189.670 36.700 189.990 ;
        RECT 36.900 189.670 37.160 189.990 ;
        RECT 35.980 187.630 36.240 187.950 ;
        RECT 36.960 187.860 37.100 189.670 ;
        RECT 37.420 189.310 37.560 194.770 ;
        RECT 37.880 192.225 38.020 195.110 ;
        RECT 41.040 194.430 41.300 194.750 ;
        RECT 40.580 194.090 40.840 194.410 ;
        RECT 38.270 193.215 38.550 193.585 ;
        RECT 39.190 193.215 39.470 193.585 ;
        RECT 38.280 193.070 38.540 193.215 ;
        RECT 37.810 191.855 38.090 192.225 ;
        RECT 38.280 189.670 38.540 189.990 ;
        RECT 37.360 188.990 37.620 189.310 ;
        RECT 36.960 187.720 38.020 187.860 ;
        RECT 35.520 184.570 35.780 184.890 ;
        RECT 35.060 178.790 35.320 179.110 ;
        RECT 35.580 176.050 35.720 184.570 ;
        RECT 36.040 183.870 36.180 187.630 ;
        RECT 36.890 186.415 37.170 186.785 ;
        RECT 36.960 184.210 37.100 186.415 ;
        RECT 36.900 184.120 37.160 184.210 ;
        RECT 36.500 183.980 37.160 184.120 ;
        RECT 35.980 183.550 36.240 183.870 ;
        RECT 36.500 183.530 36.640 183.980 ;
        RECT 36.900 183.890 37.160 183.980 ;
        RECT 36.440 183.210 36.700 183.530 ;
        RECT 36.900 183.210 37.160 183.530 ;
        RECT 35.980 179.470 36.240 179.790 ;
        RECT 35.520 175.730 35.780 176.050 ;
        RECT 34.600 173.350 34.860 173.670 ;
        RECT 34.660 171.290 34.800 173.350 ;
        RECT 36.040 171.630 36.180 179.470 ;
        RECT 36.500 179.110 36.640 183.210 ;
        RECT 36.960 179.110 37.100 183.210 ;
        RECT 37.360 180.830 37.620 181.150 ;
        RECT 37.420 179.790 37.560 180.830 ;
        RECT 37.880 179.985 38.020 187.720 ;
        RECT 38.340 185.140 38.480 189.670 ;
        RECT 39.260 187.610 39.400 193.215 ;
        RECT 39.650 191.855 39.930 192.225 ;
        RECT 39.200 187.290 39.460 187.610 ;
        RECT 39.720 185.230 39.860 191.855 ;
        RECT 40.120 189.330 40.380 189.650 ;
        RECT 38.340 185.000 39.400 185.140 ;
        RECT 38.280 184.230 38.540 184.550 ;
        RECT 38.740 184.230 39.000 184.550 ;
        RECT 39.260 184.460 39.400 185.000 ;
        RECT 39.660 184.910 39.920 185.230 ;
        RECT 39.660 184.460 39.920 184.550 ;
        RECT 39.260 184.320 39.920 184.460 ;
        RECT 39.660 184.230 39.920 184.320 ;
        RECT 38.340 183.530 38.480 184.230 ;
        RECT 38.280 183.210 38.540 183.530 ;
        RECT 38.800 180.810 38.940 184.230 ;
        RECT 39.650 183.695 39.930 184.065 ;
        RECT 39.200 183.210 39.460 183.530 ;
        RECT 39.260 182.170 39.400 183.210 ;
        RECT 39.720 182.170 39.860 183.695 ;
        RECT 39.200 181.850 39.460 182.170 ;
        RECT 39.660 181.850 39.920 182.170 ;
        RECT 39.260 181.490 39.400 181.850 ;
        RECT 39.200 181.170 39.460 181.490 ;
        RECT 39.650 180.975 39.930 181.345 ;
        RECT 38.740 180.490 39.000 180.810 ;
        RECT 37.360 179.470 37.620 179.790 ;
        RECT 37.810 179.615 38.090 179.985 ;
        RECT 36.440 178.790 36.700 179.110 ;
        RECT 36.900 178.790 37.160 179.110 ;
        RECT 37.360 178.790 37.620 179.110 ;
        RECT 37.420 178.625 37.560 178.790 ;
        RECT 37.350 178.255 37.630 178.625 ;
        RECT 39.720 178.510 39.860 180.975 ;
        RECT 38.280 178.340 38.540 178.430 ;
        RECT 38.800 178.370 39.860 178.510 ;
        RECT 38.800 178.340 38.940 178.370 ;
        RECT 38.280 178.200 38.940 178.340 ;
        RECT 38.280 178.110 38.540 178.200 ;
        RECT 39.660 177.770 39.920 178.090 ;
        RECT 38.740 175.730 39.000 176.050 ;
        RECT 36.430 174.175 36.710 174.545 ;
        RECT 36.500 173.330 36.640 174.175 ;
        RECT 36.900 173.580 37.160 173.670 ;
        RECT 38.280 173.580 38.540 173.670 ;
        RECT 36.900 173.440 38.540 173.580 ;
        RECT 36.900 173.350 37.160 173.440 ;
        RECT 38.280 173.350 38.540 173.440 ;
        RECT 36.440 173.010 36.700 173.330 ;
        RECT 37.820 172.330 38.080 172.650 ;
        RECT 37.880 171.630 38.020 172.330 ;
        RECT 35.980 171.310 36.240 171.630 ;
        RECT 37.820 171.310 38.080 171.630 ;
        RECT 34.600 170.970 34.860 171.290 ;
        RECT 38.340 170.610 38.480 173.350 ;
        RECT 33.680 170.290 33.940 170.610 ;
        RECT 38.280 170.290 38.540 170.610 ;
        RECT 35.520 169.610 35.780 169.930 ;
        RECT 31.900 157.310 32.500 157.430 ;
        RECT 35.580 157.310 35.720 169.610 ;
        RECT 38.800 165.705 38.940 175.730 ;
        RECT 39.200 173.350 39.460 173.670 ;
        RECT 39.260 171.290 39.400 173.350 ;
        RECT 39.200 170.970 39.460 171.290 ;
        RECT 39.720 170.950 39.860 177.770 ;
        RECT 40.180 177.070 40.320 189.330 ;
        RECT 40.640 181.150 40.780 194.090 ;
        RECT 41.100 192.370 41.240 194.430 ;
        RECT 42.020 193.390 42.160 203.415 ;
        RECT 42.410 200.695 42.690 201.065 ;
        RECT 42.480 197.470 42.620 200.695 ;
        RECT 42.420 197.150 42.680 197.470 ;
        RECT 42.410 195.255 42.690 195.625 ;
        RECT 42.420 195.110 42.680 195.255 ;
        RECT 41.960 193.070 42.220 193.390 ;
        RECT 41.040 192.050 41.300 192.370 ;
        RECT 41.100 189.650 41.240 192.050 ;
        RECT 41.950 191.855 42.230 192.225 ;
        RECT 42.020 189.990 42.160 191.855 ;
        RECT 42.880 190.350 43.140 190.670 ;
        RECT 41.960 189.670 42.220 189.990 ;
        RECT 41.040 189.330 41.300 189.650 ;
        RECT 41.500 189.330 41.760 189.650 ;
        RECT 41.100 187.950 41.240 189.330 ;
        RECT 41.040 187.630 41.300 187.950 ;
        RECT 41.040 186.270 41.300 186.590 ;
        RECT 41.100 184.065 41.240 186.270 ;
        RECT 41.560 185.230 41.700 189.330 ;
        RECT 41.960 188.990 42.220 189.310 ;
        RECT 42.420 188.990 42.680 189.310 ;
        RECT 42.020 186.250 42.160 188.990 ;
        RECT 41.960 185.930 42.220 186.250 ;
        RECT 41.500 184.910 41.760 185.230 ;
        RECT 41.030 183.695 41.310 184.065 ;
        RECT 41.100 182.510 41.240 183.695 ;
        RECT 41.040 182.190 41.300 182.510 ;
        RECT 41.500 181.850 41.760 182.170 ;
        RECT 40.580 180.830 40.840 181.150 ;
        RECT 41.030 179.615 41.310 179.985 ;
        RECT 41.100 179.110 41.240 179.615 ;
        RECT 41.040 178.790 41.300 179.110 ;
        RECT 40.580 178.110 40.840 178.430 ;
        RECT 41.560 178.340 41.700 181.850 ;
        RECT 42.020 179.110 42.160 185.930 ;
        RECT 42.480 185.425 42.620 188.990 ;
        RECT 42.410 185.055 42.690 185.425 ;
        RECT 42.420 184.230 42.680 184.550 ;
        RECT 42.480 184.065 42.620 184.230 ;
        RECT 42.410 183.695 42.690 184.065 ;
        RECT 42.420 183.210 42.680 183.530 ;
        RECT 42.480 182.510 42.620 183.210 ;
        RECT 42.420 182.190 42.680 182.510 ;
        RECT 42.420 181.060 42.680 181.150 ;
        RECT 42.940 181.060 43.080 190.350 ;
        RECT 43.400 189.990 43.540 205.650 ;
        RECT 43.800 198.510 44.060 198.830 ;
        RECT 43.860 192.370 44.000 198.510 ;
        RECT 44.320 197.470 44.460 206.670 ;
        RECT 45.240 201.745 45.380 209.390 ;
        RECT 46.620 209.030 46.760 211.770 ;
        RECT 46.560 208.710 46.820 209.030 ;
        RECT 47.020 208.370 47.280 208.690 ;
        RECT 47.080 206.650 47.220 208.370 ;
        RECT 48.460 208.010 48.600 213.130 ;
        RECT 48.400 207.690 48.660 208.010 ;
        RECT 47.020 206.330 47.280 206.650 ;
        RECT 47.480 205.990 47.740 206.310 ;
        RECT 48.400 206.220 48.660 206.310 ;
        RECT 48.000 206.080 48.660 206.220 ;
        RECT 46.100 205.310 46.360 205.630 ;
        RECT 46.160 203.250 46.300 205.310 ;
        RECT 47.540 205.145 47.680 205.990 ;
        RECT 47.470 204.775 47.750 205.145 ;
        RECT 46.560 203.270 46.820 203.590 ;
        RECT 45.640 202.930 45.900 203.250 ;
        RECT 46.100 202.930 46.360 203.250 ;
        RECT 44.720 201.230 44.980 201.550 ;
        RECT 45.170 201.375 45.450 201.745 ;
        RECT 44.780 197.810 44.920 201.230 ;
        RECT 45.700 200.385 45.840 202.930 ;
        RECT 46.620 201.550 46.760 203.270 ;
        RECT 47.020 202.250 47.280 202.570 ;
        RECT 46.560 201.230 46.820 201.550 ;
        RECT 47.080 200.870 47.220 202.250 ;
        RECT 46.100 200.550 46.360 200.870 ;
        RECT 47.020 200.780 47.280 200.870 ;
        RECT 46.620 200.640 47.280 200.780 ;
        RECT 45.630 200.015 45.910 200.385 ;
        RECT 46.160 197.810 46.300 200.550 ;
        RECT 44.720 197.490 44.980 197.810 ;
        RECT 45.180 197.490 45.440 197.810 ;
        RECT 46.100 197.490 46.360 197.810 ;
        RECT 44.260 197.150 44.520 197.470 ;
        RECT 44.260 195.110 44.520 195.430 ;
        RECT 44.320 193.390 44.460 195.110 ;
        RECT 44.260 193.070 44.520 193.390 ;
        RECT 43.800 192.050 44.060 192.370 ;
        RECT 44.780 190.670 44.920 197.490 ;
        RECT 45.240 194.410 45.380 197.490 ;
        RECT 46.100 195.625 46.360 195.770 ;
        RECT 46.090 195.255 46.370 195.625 ;
        RECT 46.620 195.430 46.760 200.640 ;
        RECT 47.020 200.550 47.280 200.640 ;
        RECT 47.480 199.530 47.740 199.850 ;
        RECT 47.010 198.655 47.290 199.025 ;
        RECT 47.020 198.510 47.280 198.655 ;
        RECT 47.010 197.975 47.290 198.345 ;
        RECT 46.560 195.110 46.820 195.430 ;
        RECT 47.080 194.830 47.220 197.975 ;
        RECT 46.620 194.690 47.220 194.830 ;
        RECT 45.180 194.090 45.440 194.410 ;
        RECT 44.720 190.350 44.980 190.670 ;
        RECT 43.340 189.670 43.600 189.990 ;
        RECT 45.640 189.900 45.900 189.990 ;
        RECT 45.640 189.760 46.300 189.900 ;
        RECT 45.640 189.670 45.900 189.760 ;
        RECT 45.180 189.330 45.440 189.650 ;
        RECT 43.800 188.990 44.060 189.310 ;
        RECT 43.400 184.460 43.660 184.550 ;
        RECT 43.860 184.460 44.000 188.990 ;
        RECT 45.240 188.710 45.380 189.330 ;
        RECT 46.160 188.880 46.300 189.760 ;
        RECT 46.620 189.230 46.760 194.690 ;
        RECT 47.020 192.050 47.280 192.370 ;
        RECT 47.080 189.560 47.220 192.050 ;
        RECT 47.540 190.330 47.680 199.530 ;
        RECT 48.000 198.345 48.140 206.080 ;
        RECT 48.400 205.990 48.660 206.080 ;
        RECT 48.400 202.930 48.660 203.250 ;
        RECT 48.460 201.210 48.600 202.930 ;
        RECT 48.400 200.890 48.660 201.210 ;
        RECT 48.920 198.830 49.060 214.490 ;
        RECT 53.460 211.770 53.720 212.090 ;
        RECT 49.320 210.410 49.580 210.730 ;
        RECT 49.780 210.410 50.040 210.730 ;
        RECT 49.380 209.710 49.520 210.410 ;
        RECT 49.320 209.390 49.580 209.710 ;
        RECT 49.840 206.310 49.980 210.410 ;
        RECT 51.620 206.670 51.880 206.990 ;
        RECT 49.780 205.990 50.040 206.310 ;
        RECT 50.700 205.990 50.960 206.310 ;
        RECT 49.780 205.310 50.040 205.630 ;
        RECT 49.840 200.870 49.980 205.310 ;
        RECT 50.230 203.415 50.510 203.785 ;
        RECT 50.240 203.270 50.500 203.415 ;
        RECT 50.760 202.990 50.900 205.990 ;
        RECT 51.680 204.270 51.820 206.670 ;
        RECT 52.070 204.775 52.350 205.145 ;
        RECT 51.620 203.950 51.880 204.270 ;
        RECT 51.150 203.415 51.430 203.785 ;
        RECT 52.140 203.590 52.280 204.775 ;
        RECT 52.540 203.950 52.800 204.270 ;
        RECT 52.080 203.500 52.340 203.590 ;
        RECT 51.160 203.270 51.420 203.415 ;
        RECT 51.680 203.360 52.340 203.500 ;
        RECT 50.300 202.850 50.900 202.990 ;
        RECT 49.320 200.550 49.580 200.870 ;
        RECT 49.780 200.550 50.040 200.870 ;
        RECT 48.860 198.510 49.120 198.830 ;
        RECT 47.930 197.975 48.210 198.345 ;
        RECT 49.380 198.230 49.520 200.550 ;
        RECT 50.300 200.190 50.440 202.850 ;
        RECT 51.160 202.590 51.420 202.910 ;
        RECT 50.700 201.230 50.960 201.550 ;
        RECT 50.760 200.870 50.900 201.230 ;
        RECT 51.220 200.870 51.360 202.590 ;
        RECT 50.700 200.550 50.960 200.870 ;
        RECT 51.160 200.550 51.420 200.870 ;
        RECT 51.220 200.190 51.360 200.550 ;
        RECT 50.240 199.870 50.500 200.190 ;
        RECT 51.160 199.870 51.420 200.190 ;
        RECT 49.780 199.530 50.040 199.850 ;
        RECT 48.460 198.090 49.520 198.230 ;
        RECT 47.930 197.295 48.210 197.665 ;
        RECT 48.000 195.430 48.140 197.295 ;
        RECT 48.460 195.430 48.600 198.090 ;
        RECT 48.860 197.150 49.120 197.470 ;
        RECT 49.310 197.295 49.590 197.665 ;
        RECT 47.940 195.110 48.200 195.430 ;
        RECT 48.400 195.110 48.660 195.430 ;
        RECT 48.460 194.750 48.600 195.110 ;
        RECT 48.400 194.430 48.660 194.750 ;
        RECT 47.940 194.090 48.200 194.410 ;
        RECT 48.000 192.370 48.140 194.090 ;
        RECT 48.400 192.390 48.660 192.710 ;
        RECT 47.940 192.050 48.200 192.370 ;
        RECT 48.000 190.670 48.140 192.050 ;
        RECT 47.940 190.350 48.200 190.670 ;
        RECT 47.480 190.010 47.740 190.330 ;
        RECT 48.460 190.070 48.600 192.390 ;
        RECT 48.920 190.670 49.060 197.150 ;
        RECT 48.860 190.350 49.120 190.670 ;
        RECT 48.000 189.930 48.600 190.070 ;
        RECT 47.080 189.420 47.680 189.560 ;
        RECT 46.620 189.090 47.220 189.230 ;
        RECT 46.160 188.740 46.760 188.880 ;
        RECT 45.240 188.570 45.840 188.710 ;
        RECT 45.170 187.775 45.450 188.145 ;
        RECT 45.240 187.520 45.380 187.775 ;
        RECT 45.700 187.610 45.840 188.570 ;
        RECT 45.240 187.380 45.385 187.520 ;
        RECT 45.245 186.930 45.385 187.380 ;
        RECT 45.640 187.290 45.900 187.610 ;
        RECT 44.720 186.610 44.980 186.930 ;
        RECT 45.180 186.610 45.440 186.930 ;
        RECT 45.640 186.610 45.900 186.930 ;
        RECT 44.250 185.055 44.530 185.425 ;
        RECT 43.400 184.320 44.000 184.460 ;
        RECT 43.400 184.230 43.660 184.320 ;
        RECT 44.320 183.950 44.460 185.055 ;
        RECT 44.780 184.550 44.920 186.610 ;
        RECT 45.180 185.930 45.440 186.250 ;
        RECT 44.720 184.230 44.980 184.550 ;
        RECT 42.420 180.920 43.080 181.060 ;
        RECT 43.400 183.810 44.460 183.950 ;
        RECT 43.400 181.400 43.540 183.810 ;
        RECT 44.260 183.210 44.520 183.530 ;
        RECT 44.320 182.170 44.460 183.210 ;
        RECT 44.260 181.850 44.520 182.170 ;
        RECT 44.780 182.080 44.920 184.230 ;
        RECT 45.240 184.210 45.380 185.930 ;
        RECT 45.700 185.425 45.840 186.610 ;
        RECT 46.100 186.270 46.360 186.590 ;
        RECT 45.630 185.055 45.910 185.425 ;
        RECT 45.640 184.570 45.900 184.890 ;
        RECT 45.180 183.890 45.440 184.210 ;
        RECT 45.180 182.080 45.440 182.170 ;
        RECT 44.780 181.940 45.440 182.080 ;
        RECT 45.180 181.850 45.440 181.940 ;
        RECT 43.800 181.400 44.060 181.490 ;
        RECT 43.400 181.260 44.060 181.400 ;
        RECT 42.420 180.830 42.680 180.920 ;
        RECT 42.420 179.470 42.680 179.790 ;
        RECT 41.960 178.790 42.220 179.110 ;
        RECT 41.100 178.200 41.700 178.340 ;
        RECT 40.120 176.750 40.380 177.070 ;
        RECT 40.640 174.010 40.780 178.110 ;
        RECT 40.580 173.690 40.840 174.010 ;
        RECT 41.100 173.330 41.240 178.200 ;
        RECT 42.480 177.070 42.620 179.470 ;
        RECT 42.880 178.790 43.140 179.110 ;
        RECT 42.420 176.750 42.680 177.070 ;
        RECT 41.490 176.215 41.770 176.585 ;
        RECT 41.960 176.300 42.220 176.390 ;
        RECT 42.940 176.300 43.080 178.790 ;
        RECT 43.400 178.430 43.540 181.260 ;
        RECT 43.800 181.170 44.060 181.260 ;
        RECT 44.320 181.150 44.460 181.850 ;
        RECT 45.700 181.490 45.840 184.570 ;
        RECT 46.160 184.550 46.300 186.270 ;
        RECT 46.620 185.230 46.760 188.740 ;
        RECT 47.080 187.950 47.220 189.090 ;
        RECT 47.020 187.630 47.280 187.950 ;
        RECT 47.020 186.610 47.280 186.930 ;
        RECT 46.560 184.910 46.820 185.230 ;
        RECT 46.100 184.230 46.360 184.550 ;
        RECT 46.560 184.230 46.820 184.550 ;
        RECT 46.090 183.695 46.370 184.065 ;
        RECT 45.640 181.170 45.900 181.490 ;
        RECT 46.160 181.400 46.300 183.695 ;
        RECT 46.620 182.705 46.760 184.230 ;
        RECT 47.080 183.530 47.220 186.610 ;
        RECT 47.540 184.550 47.680 189.420 ;
        RECT 48.000 184.550 48.140 189.930 ;
        RECT 48.390 189.135 48.670 189.505 ;
        RECT 48.460 187.270 48.600 189.135 ;
        RECT 48.400 186.950 48.660 187.270 ;
        RECT 47.480 184.230 47.740 184.550 ;
        RECT 47.940 184.230 48.200 184.550 ;
        RECT 48.390 183.695 48.670 184.065 ;
        RECT 47.020 183.210 47.280 183.530 ;
        RECT 46.550 182.335 46.830 182.705 ;
        RECT 47.480 182.420 47.740 182.510 ;
        RECT 47.080 182.280 47.740 182.420 ;
        RECT 47.930 182.335 48.210 182.705 ;
        RECT 46.560 181.400 46.820 181.490 ;
        RECT 46.160 181.260 46.820 181.400 ;
        RECT 46.560 181.170 46.820 181.260 ;
        RECT 44.260 180.830 44.520 181.150 ;
        RECT 45.700 179.790 45.840 181.170 ;
        RECT 46.100 180.490 46.360 180.810 ;
        RECT 47.080 180.720 47.220 182.280 ;
        RECT 47.480 182.190 47.740 182.280 ;
        RECT 48.000 182.170 48.140 182.335 ;
        RECT 47.940 181.850 48.200 182.170 ;
        RECT 47.480 181.170 47.740 181.490 ;
        RECT 46.620 180.580 47.220 180.720 ;
        RECT 45.640 179.470 45.900 179.790 ;
        RECT 44.260 178.790 44.520 179.110 ;
        RECT 43.340 178.110 43.600 178.430 ;
        RECT 43.800 177.945 44.060 178.090 ;
        RECT 43.790 177.575 44.070 177.945 ;
        RECT 41.500 176.070 41.760 176.215 ;
        RECT 41.960 176.160 43.080 176.300 ;
        RECT 41.960 176.070 42.220 176.160 ;
        RECT 42.480 175.820 43.080 175.960 ;
        RECT 41.960 175.390 42.220 175.710 ;
        RECT 41.490 174.855 41.770 175.225 ;
        RECT 41.560 173.330 41.700 174.855 ;
        RECT 42.020 173.670 42.160 175.390 ;
        RECT 41.960 173.350 42.220 173.670 ;
        RECT 41.040 173.010 41.300 173.330 ;
        RECT 41.500 173.010 41.760 173.330 ;
        RECT 42.480 173.185 42.620 175.820 ;
        RECT 41.100 171.630 41.240 173.010 ;
        RECT 42.410 172.815 42.690 173.185 ;
        RECT 41.040 171.310 41.300 171.630 ;
        RECT 39.660 170.630 39.920 170.950 ;
        RECT 42.940 170.270 43.080 175.820 ;
        RECT 43.340 175.730 43.600 176.050 ;
        RECT 43.860 175.905 44.000 177.575 ;
        RECT 44.320 175.960 44.460 178.790 ;
        RECT 44.720 178.450 44.980 178.770 ;
        RECT 44.780 176.730 44.920 178.450 ;
        RECT 45.640 178.110 45.900 178.430 ;
        RECT 45.180 177.770 45.440 178.090 ;
        RECT 45.700 177.945 45.840 178.110 ;
        RECT 45.240 177.070 45.380 177.770 ;
        RECT 45.630 177.575 45.910 177.945 ;
        RECT 46.160 177.265 46.300 180.490 ;
        RECT 46.620 179.020 46.760 180.580 ;
        RECT 47.020 179.020 47.280 179.110 ;
        RECT 46.620 178.880 47.280 179.020 ;
        RECT 47.540 179.020 47.680 181.170 ;
        RECT 47.940 180.830 48.200 181.150 ;
        RECT 48.000 179.790 48.140 180.830 ;
        RECT 47.940 179.470 48.200 179.790 ;
        RECT 47.540 178.880 48.140 179.020 ;
        RECT 47.020 178.790 47.280 178.880 ;
        RECT 47.020 178.110 47.280 178.430 ;
        RECT 48.000 178.340 48.140 178.880 ;
        RECT 47.540 178.200 48.140 178.340 ;
        RECT 47.080 177.265 47.220 178.110 ;
        RECT 45.180 176.750 45.440 177.070 ;
        RECT 46.090 176.895 46.370 177.265 ;
        RECT 47.010 176.895 47.290 177.265 ;
        RECT 44.720 176.410 44.980 176.730 ;
        RECT 43.400 173.670 43.540 175.730 ;
        RECT 43.790 175.535 44.070 175.905 ;
        RECT 44.320 175.820 44.920 175.960 ;
        RECT 43.340 173.350 43.600 173.670 ;
        RECT 43.340 172.330 43.600 172.650 ;
        RECT 43.400 170.610 43.540 172.330 ;
        RECT 43.340 170.290 43.600 170.610 ;
        RECT 43.800 170.290 44.060 170.610 ;
        RECT 42.880 169.950 43.140 170.270 ;
        RECT 38.730 165.335 39.010 165.705 ;
        RECT 41.950 163.975 42.230 164.345 ;
        RECT 38.730 163.295 39.010 163.665 ;
        RECT 38.800 157.310 38.940 163.295 ;
        RECT 42.020 157.310 42.160 163.975 ;
        RECT 43.860 162.305 44.000 170.290 ;
        RECT 44.780 169.105 44.920 175.820 ;
        RECT 45.240 171.145 45.380 176.750 ;
        RECT 47.020 176.070 47.280 176.390 ;
        RECT 47.080 175.905 47.220 176.070 ;
        RECT 45.640 175.390 45.900 175.710 ;
        RECT 47.010 175.535 47.290 175.905 ;
        RECT 47.540 175.430 47.680 178.200 ;
        RECT 48.460 176.730 48.600 183.695 ;
        RECT 48.920 182.510 49.060 190.350 ;
        RECT 49.380 189.990 49.520 197.295 ;
        RECT 49.840 195.625 49.980 199.530 ;
        RECT 50.300 197.130 50.440 199.870 ;
        RECT 50.240 196.810 50.500 197.130 ;
        RECT 51.680 196.110 51.820 203.360 ;
        RECT 52.080 203.270 52.340 203.360 ;
        RECT 52.600 202.425 52.740 203.950 ;
        RECT 53.000 202.930 53.260 203.250 ;
        RECT 52.530 202.055 52.810 202.425 ;
        RECT 52.080 200.550 52.340 200.870 ;
        RECT 52.140 197.810 52.280 200.550 ;
        RECT 52.540 199.530 52.800 199.850 ;
        RECT 52.600 197.810 52.740 199.530 ;
        RECT 52.080 197.490 52.340 197.810 ;
        RECT 52.540 197.665 52.800 197.810 ;
        RECT 51.620 195.790 51.880 196.110 ;
        RECT 49.770 195.255 50.050 195.625 ;
        RECT 51.160 195.110 51.420 195.430 ;
        RECT 51.620 195.110 51.880 195.430 ;
        RECT 49.780 194.430 50.040 194.750 ;
        RECT 49.840 190.330 49.980 194.430 ;
        RECT 50.240 194.090 50.500 194.410 ;
        RECT 50.300 192.030 50.440 194.090 ;
        RECT 51.220 192.370 51.360 195.110 ;
        RECT 51.680 193.390 51.820 195.110 ;
        RECT 51.620 193.070 51.880 193.390 ;
        RECT 52.140 193.050 52.280 197.490 ;
        RECT 52.530 197.295 52.810 197.665 ;
        RECT 52.540 195.110 52.800 195.430 ;
        RECT 52.600 193.585 52.740 195.110 ;
        RECT 53.060 195.090 53.200 202.930 ;
        RECT 53.520 198.150 53.660 211.770 ;
        RECT 54.900 208.350 55.040 215.510 ;
        RECT 58.120 215.490 58.260 223.160 ;
        RECT 58.060 215.170 58.320 215.490 ;
        RECT 57.600 214.150 57.860 214.470 ;
        RECT 55.750 210.895 56.030 211.265 ;
        RECT 54.840 208.030 55.100 208.350 ;
        RECT 54.900 206.310 55.040 208.030 ;
        RECT 55.300 207.690 55.560 208.010 ;
        RECT 54.840 205.990 55.100 206.310 ;
        RECT 54.900 205.825 55.040 205.990 ;
        RECT 54.380 205.310 54.640 205.630 ;
        RECT 54.830 205.455 55.110 205.825 ;
        RECT 54.440 203.590 54.580 205.310 ;
        RECT 55.360 203.930 55.500 207.690 ;
        RECT 55.820 206.310 55.960 210.895 ;
        RECT 56.670 206.815 56.950 207.185 ;
        RECT 55.760 205.990 56.020 206.310 ;
        RECT 56.220 205.990 56.480 206.310 ;
        RECT 55.820 203.930 55.960 205.990 ;
        RECT 56.280 205.630 56.420 205.990 ;
        RECT 56.220 205.310 56.480 205.630 ;
        RECT 55.300 203.610 55.560 203.930 ;
        RECT 55.760 203.610 56.020 203.930 ;
        RECT 54.380 203.270 54.640 203.590 ;
        RECT 54.840 203.270 55.100 203.590 ;
        RECT 53.920 202.590 54.180 202.910 ;
        RECT 53.980 198.345 54.120 202.590 ;
        RECT 54.440 202.425 54.580 203.270 ;
        RECT 54.370 202.055 54.650 202.425 ;
        RECT 54.380 200.210 54.640 200.530 ;
        RECT 53.460 197.830 53.720 198.150 ;
        RECT 53.910 197.975 54.190 198.345 ;
        RECT 53.920 197.830 54.180 197.975 ;
        RECT 53.520 197.550 53.660 197.830 ;
        RECT 54.440 197.810 54.580 200.210 ;
        RECT 53.520 197.410 54.120 197.550 ;
        RECT 54.380 197.490 54.640 197.810 ;
        RECT 53.460 196.810 53.720 197.130 ;
        RECT 53.000 194.770 53.260 195.090 ;
        RECT 52.530 193.215 52.810 193.585 ;
        RECT 52.080 192.730 52.340 193.050 ;
        RECT 51.160 192.050 51.420 192.370 ;
        RECT 50.240 191.710 50.500 192.030 ;
        RECT 50.700 191.370 50.960 191.690 ;
        RECT 49.780 190.010 50.040 190.330 ;
        RECT 49.320 189.670 49.580 189.990 ;
        RECT 50.760 189.505 50.900 191.370 ;
        RECT 51.220 190.670 51.360 192.050 ;
        RECT 51.610 191.855 51.890 192.225 ;
        RECT 51.160 190.350 51.420 190.670 ;
        RECT 51.150 189.815 51.430 190.185 ;
        RECT 49.310 189.135 49.590 189.505 ;
        RECT 50.690 189.135 50.970 189.505 ;
        RECT 49.380 186.930 49.520 189.135 ;
        RECT 50.230 188.455 50.510 188.825 ;
        RECT 50.700 188.650 50.960 188.970 ;
        RECT 50.300 187.950 50.440 188.455 ;
        RECT 50.240 187.630 50.500 187.950 ;
        RECT 49.780 187.350 50.040 187.610 ;
        RECT 49.780 187.290 50.440 187.350 ;
        RECT 49.840 187.210 50.440 187.290 ;
        RECT 49.320 186.610 49.580 186.930 ;
        RECT 49.320 184.230 49.580 184.550 ;
        RECT 49.380 182.705 49.520 184.230 ;
        RECT 49.770 183.015 50.050 183.385 ;
        RECT 48.860 182.190 49.120 182.510 ;
        RECT 49.310 182.335 49.590 182.705 ;
        RECT 49.310 181.655 49.590 182.025 ;
        RECT 49.320 181.510 49.580 181.655 ;
        RECT 49.840 181.490 49.980 183.015 ;
        RECT 49.780 181.170 50.040 181.490 ;
        RECT 50.300 179.305 50.440 187.210 ;
        RECT 50.760 185.230 50.900 188.650 ;
        RECT 51.220 187.950 51.360 189.815 ;
        RECT 51.160 187.630 51.420 187.950 ;
        RECT 50.700 184.910 50.960 185.230 ;
        RECT 51.680 184.890 51.820 191.855 ;
        RECT 52.140 188.145 52.280 192.730 ;
        RECT 52.600 189.650 52.740 193.215 ;
        RECT 53.000 193.070 53.260 193.390 ;
        RECT 52.540 189.330 52.800 189.650 ;
        RECT 53.060 189.310 53.200 193.070 ;
        RECT 53.000 188.990 53.260 189.310 ;
        RECT 52.990 188.455 53.270 188.825 ;
        RECT 52.070 187.775 52.350 188.145 ;
        RECT 52.530 185.055 52.810 185.425 ;
        RECT 52.600 184.890 52.740 185.055 ;
        RECT 51.620 184.570 51.880 184.890 ;
        RECT 52.540 184.570 52.800 184.890 ;
        RECT 53.060 181.490 53.200 188.455 ;
        RECT 53.520 185.230 53.660 196.810 ;
        RECT 53.980 192.370 54.120 197.410 ;
        RECT 54.380 196.810 54.640 197.130 ;
        RECT 54.440 193.050 54.580 196.810 ;
        RECT 54.380 192.730 54.640 193.050 ;
        RECT 53.920 192.050 54.180 192.370 ;
        RECT 53.920 190.350 54.180 190.670 ;
        RECT 54.380 190.350 54.640 190.670 ;
        RECT 53.980 186.590 54.120 190.350 ;
        RECT 54.440 186.930 54.580 190.350 ;
        RECT 54.380 186.610 54.640 186.930 ;
        RECT 53.920 186.270 54.180 186.590 ;
        RECT 53.460 184.910 53.720 185.230 ;
        RECT 53.980 184.210 54.120 186.270 ;
        RECT 54.380 185.930 54.640 186.250 ;
        RECT 54.440 184.210 54.580 185.930 ;
        RECT 54.900 184.550 55.040 203.270 ;
        RECT 56.740 203.160 56.880 206.815 ;
        RECT 57.140 205.650 57.400 205.970 ;
        RECT 55.360 203.020 56.880 203.160 ;
        RECT 55.360 198.830 55.500 203.020 ;
        RECT 57.200 202.570 57.340 205.650 ;
        RECT 55.760 202.250 56.020 202.570 ;
        RECT 57.140 202.250 57.400 202.570 ;
        RECT 55.300 198.510 55.560 198.830 ;
        RECT 55.820 198.345 55.960 202.250 ;
        RECT 57.660 201.210 57.800 214.150 ;
        RECT 58.520 213.470 58.780 213.790 ;
        RECT 58.580 206.990 58.720 213.470 ;
        RECT 60.820 211.430 61.080 211.750 ;
        RECT 60.360 208.370 60.620 208.690 ;
        RECT 59.900 207.690 60.160 208.010 ;
        RECT 59.960 206.990 60.100 207.690 ;
        RECT 58.520 206.670 58.780 206.990 ;
        RECT 59.900 206.900 60.160 206.990 ;
        RECT 59.500 206.760 60.160 206.900 ;
        RECT 58.980 205.990 59.240 206.310 ;
        RECT 58.060 205.310 58.320 205.630 ;
        RECT 58.120 201.550 58.260 205.310 ;
        RECT 59.040 204.270 59.180 205.990 ;
        RECT 58.980 203.950 59.240 204.270 ;
        RECT 58.060 201.230 58.320 201.550 ;
        RECT 57.600 200.890 57.860 201.210 ;
        RECT 58.510 200.695 58.790 201.065 ;
        RECT 58.060 199.870 58.320 200.190 ;
        RECT 56.220 198.510 56.480 198.830 ;
        RECT 56.670 198.655 56.950 199.025 ;
        RECT 55.750 197.975 56.030 198.345 ;
        RECT 56.280 198.150 56.420 198.510 ;
        RECT 56.220 197.830 56.480 198.150 ;
        RECT 55.290 197.295 55.570 197.665 ;
        RECT 56.740 197.470 56.880 198.655 ;
        RECT 57.140 198.060 57.400 198.150 ;
        RECT 57.140 197.920 57.800 198.060 ;
        RECT 57.140 197.830 57.400 197.920 ;
        RECT 56.680 197.380 56.940 197.470 ;
        RECT 55.360 195.770 55.500 197.295 ;
        RECT 56.680 197.240 57.340 197.380 ;
        RECT 56.680 197.150 56.940 197.240 ;
        RECT 55.760 196.810 56.020 197.130 ;
        RECT 55.300 195.450 55.560 195.770 ;
        RECT 55.820 195.430 55.960 196.810 ;
        RECT 56.680 195.450 56.940 195.770 ;
        RECT 55.760 195.110 56.020 195.430 ;
        RECT 55.300 194.430 55.560 194.750 ;
        RECT 55.360 192.110 55.500 194.430 ;
        RECT 55.820 192.710 55.960 195.110 ;
        RECT 56.220 194.090 56.480 194.410 ;
        RECT 56.280 192.710 56.420 194.090 ;
        RECT 56.740 193.050 56.880 195.450 ;
        RECT 57.200 195.430 57.340 197.240 ;
        RECT 57.660 195.430 57.800 197.920 ;
        RECT 58.120 197.810 58.260 199.870 ;
        RECT 58.060 197.490 58.320 197.810 ;
        RECT 58.120 195.430 58.260 197.490 ;
        RECT 57.140 195.110 57.400 195.430 ;
        RECT 57.600 195.110 57.860 195.430 ;
        RECT 58.060 195.110 58.320 195.430 ;
        RECT 58.580 195.340 58.720 200.695 ;
        RECT 58.980 198.740 59.240 198.830 ;
        RECT 59.500 198.740 59.640 206.760 ;
        RECT 59.900 206.670 60.160 206.760 ;
        RECT 59.890 204.095 60.170 204.465 ;
        RECT 59.900 203.950 60.160 204.095 ;
        RECT 59.900 202.930 60.160 203.250 ;
        RECT 59.960 200.870 60.100 202.930 ;
        RECT 59.900 200.550 60.160 200.870 ;
        RECT 60.420 199.850 60.560 208.370 ;
        RECT 60.880 206.990 61.020 211.430 ;
        RECT 61.340 209.710 61.480 223.160 ;
        RECT 79.680 222.990 79.940 223.310 ;
        RECT 83.810 223.135 84.090 223.505 ;
        RECT 93.470 223.160 93.750 223.660 ;
        RECT 96.690 223.160 96.970 223.660 ;
        RECT 103.130 223.160 103.410 223.660 ;
        RECT 106.350 223.160 106.630 223.660 ;
        RECT 109.570 223.160 109.850 223.660 ;
        RECT 112.790 223.160 113.070 223.660 ;
        RECT 67.260 218.570 67.520 218.890 ;
        RECT 61.740 215.510 62.000 215.830 ;
        RECT 61.800 211.750 61.940 215.510 ;
        RECT 66.800 214.830 67.060 215.150 ;
        RECT 66.860 212.090 67.000 214.830 ;
        RECT 66.800 211.770 67.060 212.090 ;
        RECT 61.740 211.430 62.000 211.750 ;
        RECT 63.120 211.430 63.380 211.750 ;
        RECT 63.180 210.730 63.320 211.430 ;
        RECT 67.320 211.070 67.460 218.570 ;
        RECT 75.540 218.230 75.800 218.550 ;
        RECT 71.400 217.550 71.660 217.870 ;
        RECT 68.640 215.170 68.900 215.490 ;
        RECT 68.700 212.430 68.840 215.170 ;
        RECT 71.460 212.430 71.600 217.550 ;
        RECT 73.700 213.470 73.960 213.790 ;
        RECT 68.640 212.110 68.900 212.430 ;
        RECT 69.100 212.110 69.360 212.430 ;
        RECT 71.400 212.110 71.660 212.430 ;
        RECT 67.720 211.430 67.980 211.750 ;
        RECT 67.260 210.750 67.520 211.070 ;
        RECT 63.120 210.410 63.380 210.730 ;
        RECT 61.280 209.390 61.540 209.710 ;
        RECT 63.580 209.390 63.840 209.710 ;
        RECT 67.260 209.390 67.520 209.710 ;
        RECT 61.270 208.175 61.550 208.545 ;
        RECT 62.200 208.370 62.460 208.690 ;
        RECT 63.120 208.370 63.380 208.690 ;
        RECT 60.820 206.670 61.080 206.990 ;
        RECT 60.810 206.135 61.090 206.505 ;
        RECT 60.360 199.530 60.620 199.850 ;
        RECT 60.880 199.760 61.020 206.135 ;
        RECT 61.340 203.250 61.480 208.175 ;
        RECT 62.260 206.505 62.400 208.370 ;
        RECT 63.180 206.990 63.320 208.370 ;
        RECT 62.660 206.670 62.920 206.990 ;
        RECT 63.120 206.670 63.380 206.990 ;
        RECT 62.190 206.135 62.470 206.505 ;
        RECT 61.280 202.930 61.540 203.250 ;
        RECT 62.720 203.160 62.860 206.670 ;
        RECT 63.120 205.030 63.380 205.290 ;
        RECT 63.640 205.030 63.780 209.390 ;
        RECT 64.950 208.855 65.230 209.225 ;
        RECT 65.020 208.690 65.160 208.855 ;
        RECT 64.960 208.370 65.220 208.690 ;
        RECT 66.800 208.370 67.060 208.690 ;
        RECT 64.500 208.030 64.760 208.350 ;
        RECT 64.560 206.310 64.700 208.030 ;
        RECT 65.880 207.865 66.140 208.010 ;
        RECT 65.870 207.495 66.150 207.865 ;
        RECT 64.500 205.990 64.760 206.310 ;
        RECT 66.860 205.970 67.000 208.370 ;
        RECT 67.320 206.990 67.460 209.390 ;
        RECT 67.780 207.185 67.920 211.430 ;
        RECT 68.640 208.600 68.900 208.690 ;
        RECT 69.160 208.600 69.300 212.110 ;
        RECT 73.760 211.750 73.900 213.470 ;
        RECT 75.600 212.430 75.740 218.230 ;
        RECT 76.920 217.210 77.180 217.530 ;
        RECT 76.000 216.870 76.260 217.190 ;
        RECT 75.540 212.110 75.800 212.430 ;
        RECT 70.480 211.430 70.740 211.750 ;
        RECT 71.400 211.430 71.660 211.750 ;
        RECT 73.700 211.430 73.960 211.750 ;
        RECT 69.560 209.390 69.820 209.710 ;
        RECT 68.640 208.460 69.300 208.600 ;
        RECT 68.640 208.370 68.900 208.460 ;
        RECT 68.180 207.690 68.440 208.010 ;
        RECT 69.100 207.920 69.360 208.010 ;
        RECT 68.700 207.780 69.360 207.920 ;
        RECT 67.260 206.670 67.520 206.990 ;
        RECT 67.710 206.815 67.990 207.185 ;
        RECT 67.260 206.220 67.520 206.310 ;
        RECT 67.260 206.080 67.920 206.220 ;
        RECT 67.260 205.990 67.520 206.080 ;
        RECT 64.960 205.650 65.220 205.970 ;
        RECT 63.120 204.970 63.780 205.030 ;
        RECT 64.500 204.970 64.760 205.290 ;
        RECT 63.180 204.890 63.780 204.970 ;
        RECT 64.560 203.250 64.700 204.970 ;
        RECT 65.020 204.465 65.160 205.650 ;
        RECT 66.330 205.455 66.610 205.825 ;
        RECT 66.800 205.710 67.060 205.970 ;
        RECT 66.800 205.650 67.460 205.710 ;
        RECT 66.860 205.570 67.460 205.650 ;
        RECT 64.950 204.095 65.230 204.465 ;
        RECT 66.400 203.930 66.540 205.455 ;
        RECT 67.320 205.290 67.460 205.570 ;
        RECT 66.800 204.970 67.060 205.290 ;
        RECT 67.260 204.970 67.520 205.290 ;
        RECT 66.340 203.610 66.600 203.930 ;
        RECT 63.120 203.160 63.380 203.250 ;
        RECT 62.720 203.020 63.380 203.160 ;
        RECT 63.120 202.930 63.380 203.020 ;
        RECT 64.040 202.930 64.300 203.250 ;
        RECT 64.500 202.930 64.760 203.250 ;
        RECT 64.960 202.930 65.220 203.250 ;
        RECT 61.280 202.250 61.540 202.570 ;
        RECT 61.340 200.530 61.480 202.250 ;
        RECT 61.740 201.230 62.000 201.550 ;
        RECT 61.800 201.065 61.940 201.230 ;
        RECT 61.730 200.695 62.010 201.065 ;
        RECT 62.660 200.550 62.920 200.870 ;
        RECT 61.280 200.210 61.540 200.530 ;
        RECT 60.880 199.620 61.940 199.760 ;
        RECT 58.980 198.600 60.100 198.740 ;
        RECT 58.980 198.510 59.240 198.600 ;
        RECT 58.970 197.975 59.250 198.345 ;
        RECT 59.040 197.810 59.180 197.975 ;
        RECT 58.980 197.490 59.240 197.810 ;
        RECT 59.440 195.340 59.700 195.430 ;
        RECT 58.580 195.200 59.700 195.340 ;
        RECT 59.440 195.110 59.700 195.200 ;
        RECT 56.680 192.730 56.940 193.050 ;
        RECT 55.760 192.390 56.020 192.710 ;
        RECT 56.220 192.390 56.480 192.710 ;
        RECT 56.740 192.370 56.880 192.730 ;
        RECT 55.360 191.970 55.960 192.110 ;
        RECT 56.680 192.050 56.940 192.370 ;
        RECT 55.300 191.370 55.560 191.690 ;
        RECT 55.360 189.900 55.500 191.370 ;
        RECT 55.820 190.670 55.960 191.970 ;
        RECT 56.220 191.710 56.480 192.030 ;
        RECT 55.760 190.350 56.020 190.670 ;
        RECT 55.760 189.900 56.020 189.990 ;
        RECT 55.360 189.760 56.020 189.900 ;
        RECT 55.760 189.670 56.020 189.760 ;
        RECT 55.300 188.990 55.560 189.310 ;
        RECT 55.360 187.270 55.500 188.990 ;
        RECT 55.820 188.825 55.960 189.670 ;
        RECT 55.750 188.455 56.030 188.825 ;
        RECT 55.300 186.950 55.560 187.270 ;
        RECT 55.820 186.930 55.960 188.455 ;
        RECT 55.760 186.610 56.020 186.930 ;
        RECT 56.280 186.250 56.420 191.710 ;
        RECT 57.200 191.600 57.340 195.110 ;
        RECT 57.660 192.225 57.800 195.110 ;
        RECT 57.590 191.855 57.870 192.225 ;
        RECT 57.200 191.460 57.800 191.600 ;
        RECT 57.140 190.010 57.400 190.330 ;
        RECT 56.680 188.990 56.940 189.310 ;
        RECT 56.740 187.610 56.880 188.990 ;
        RECT 57.200 188.145 57.340 190.010 ;
        RECT 57.130 187.775 57.410 188.145 ;
        RECT 56.680 187.290 56.940 187.610 ;
        RECT 56.740 186.930 56.880 187.290 ;
        RECT 56.680 186.610 56.940 186.930 ;
        RECT 57.660 186.500 57.800 191.460 ;
        RECT 57.200 186.360 57.800 186.500 ;
        RECT 56.220 185.930 56.480 186.250 ;
        RECT 54.840 184.230 55.100 184.550 ;
        RECT 53.920 183.890 54.180 184.210 ;
        RECT 54.380 183.890 54.640 184.210 ;
        RECT 55.760 183.890 56.020 184.210 ;
        RECT 55.300 183.210 55.560 183.530 ;
        RECT 53.000 181.170 53.260 181.490 ;
        RECT 54.380 181.170 54.640 181.490 ;
        RECT 53.920 180.830 54.180 181.150 ;
        RECT 52.080 180.490 52.340 180.810 ;
        RECT 53.000 180.490 53.260 180.810 ;
        RECT 48.850 178.935 49.130 179.305 ;
        RECT 48.920 178.770 49.060 178.935 ;
        RECT 49.320 178.790 49.580 179.110 ;
        RECT 49.780 178.790 50.040 179.110 ;
        RECT 50.230 178.935 50.510 179.305 ;
        RECT 51.620 178.790 51.880 179.110 ;
        RECT 48.860 178.450 49.120 178.770 ;
        RECT 48.860 177.770 49.120 178.090 ;
        RECT 47.930 176.215 48.210 176.585 ;
        RECT 48.400 176.410 48.660 176.730 ;
        RECT 48.000 176.050 48.140 176.215 ;
        RECT 47.940 175.730 48.200 176.050 ;
        RECT 48.400 175.730 48.660 176.050 ;
        RECT 48.460 175.430 48.600 175.730 ;
        RECT 45.700 172.990 45.840 175.390 ;
        RECT 47.540 175.290 48.600 175.430 ;
        RECT 48.920 175.370 49.060 177.770 ;
        RECT 49.380 177.070 49.520 178.790 ;
        RECT 49.320 176.750 49.580 177.070 ;
        RECT 47.480 173.350 47.740 173.670 ;
        RECT 45.640 172.670 45.900 172.990 ;
        RECT 45.170 170.775 45.450 171.145 ;
        RECT 46.560 170.970 46.820 171.290 ;
        RECT 46.620 170.610 46.760 170.970 ;
        RECT 46.560 170.290 46.820 170.610 ;
        RECT 45.180 169.610 45.440 169.930 ;
        RECT 44.710 168.735 44.990 169.105 ;
        RECT 43.790 161.935 44.070 162.305 ;
        RECT 45.240 157.310 45.380 169.610 ;
        RECT 47.540 168.570 47.680 173.350 ;
        RECT 48.460 171.825 48.600 175.290 ;
        RECT 48.860 175.050 49.120 175.370 ;
        RECT 49.840 173.070 49.980 178.790 ;
        RECT 51.160 178.110 51.420 178.430 ;
        RECT 50.240 177.770 50.500 178.090 ;
        RECT 50.700 177.770 50.960 178.090 ;
        RECT 49.380 172.930 49.980 173.070 ;
        RECT 48.390 171.455 48.670 171.825 ;
        RECT 48.860 171.310 49.120 171.630 ;
        RECT 48.400 169.610 48.660 169.930 ;
        RECT 48.920 169.785 49.060 171.310 ;
        RECT 49.380 171.290 49.520 172.930 ;
        RECT 49.780 172.330 50.040 172.650 ;
        RECT 49.320 170.970 49.580 171.290 ;
        RECT 49.840 170.610 49.980 172.330 ;
        RECT 49.780 170.290 50.040 170.610 ;
        RECT 47.480 168.250 47.740 168.570 ;
        RECT 48.460 157.310 48.600 169.610 ;
        RECT 48.850 169.415 49.130 169.785 ;
        RECT 50.300 168.910 50.440 177.770 ;
        RECT 50.760 176.050 50.900 177.770 ;
        RECT 50.700 175.730 50.960 176.050 ;
        RECT 50.240 168.590 50.500 168.910 ;
        RECT 51.220 157.350 51.360 178.110 ;
        RECT 51.680 174.545 51.820 178.790 ;
        RECT 52.140 178.430 52.280 180.490 ;
        RECT 52.530 179.615 52.810 179.985 ;
        RECT 52.080 178.110 52.340 178.430 ;
        RECT 52.140 176.050 52.280 178.110 ;
        RECT 52.600 176.050 52.740 179.615 ;
        RECT 52.080 175.730 52.340 176.050 ;
        RECT 52.540 175.730 52.800 176.050 ;
        RECT 51.610 174.175 51.890 174.545 ;
        RECT 52.080 170.970 52.340 171.290 ;
        RECT 51.620 169.610 51.880 169.930 ;
        RECT 51.680 168.425 51.820 169.610 ;
        RECT 51.610 168.055 51.890 168.425 ;
        RECT 52.140 167.630 52.280 170.970 ;
        RECT 53.060 170.465 53.200 180.490 ;
        RECT 53.980 179.110 54.120 180.830 ;
        RECT 54.440 179.985 54.580 181.170 ;
        RECT 54.370 179.615 54.650 179.985 ;
        RECT 54.440 179.110 54.580 179.615 ;
        RECT 53.460 178.790 53.720 179.110 ;
        RECT 53.920 178.790 54.180 179.110 ;
        RECT 54.380 178.790 54.640 179.110 ;
        RECT 53.520 177.945 53.660 178.790 ;
        RECT 53.450 177.575 53.730 177.945 ;
        RECT 53.520 176.585 53.660 177.575 ;
        RECT 53.450 176.215 53.730 176.585 ;
        RECT 53.520 175.710 53.660 176.215 ;
        RECT 53.980 176.050 54.120 178.790 ;
        RECT 53.920 175.730 54.180 176.050 ;
        RECT 53.460 175.390 53.720 175.710 ;
        RECT 53.460 174.260 53.720 174.350 ;
        RECT 53.980 174.260 54.120 175.730 ;
        RECT 54.440 174.350 54.580 178.790 ;
        RECT 54.840 177.770 55.100 178.090 ;
        RECT 54.900 176.050 55.040 177.770 ;
        RECT 54.840 175.730 55.100 176.050 ;
        RECT 55.360 175.430 55.500 183.210 ;
        RECT 55.820 182.170 55.960 183.890 ;
        RECT 56.220 183.385 56.480 183.530 ;
        RECT 56.210 183.015 56.490 183.385 ;
        RECT 55.760 181.850 56.020 182.170 ;
        RECT 55.820 181.490 55.960 181.850 ;
        RECT 56.210 181.655 56.490 182.025 ;
        RECT 55.760 181.170 56.020 181.490 ;
        RECT 56.280 179.110 56.420 181.655 ;
        RECT 56.220 178.790 56.480 179.110 ;
        RECT 56.680 178.790 56.940 179.110 ;
        RECT 56.220 178.110 56.480 178.430 ;
        RECT 56.280 175.790 56.420 178.110 ;
        RECT 56.740 178.090 56.880 178.790 ;
        RECT 57.200 178.090 57.340 186.360 ;
        RECT 57.590 185.735 57.870 186.105 ;
        RECT 57.660 181.830 57.800 185.735 ;
        RECT 58.120 185.425 58.260 195.110 ;
        RECT 58.980 194.660 59.240 194.750 ;
        RECT 58.580 194.520 59.240 194.660 ;
        RECT 58.580 192.540 58.720 194.520 ;
        RECT 58.980 194.430 59.240 194.520 ;
        RECT 58.520 192.220 58.780 192.540 ;
        RECT 59.500 190.670 59.640 195.110 ;
        RECT 59.440 190.350 59.700 190.670 ;
        RECT 58.980 190.185 59.240 190.330 ;
        RECT 58.520 189.670 58.780 189.990 ;
        RECT 58.970 189.815 59.250 190.185 ;
        RECT 58.580 186.930 58.720 189.670 ;
        RECT 58.520 186.610 58.780 186.930 ;
        RECT 58.050 185.055 58.330 185.425 ;
        RECT 59.960 185.140 60.100 198.600 ;
        RECT 60.360 198.170 60.620 198.490 ;
        RECT 61.280 198.170 61.540 198.490 ;
        RECT 60.420 196.110 60.560 198.170 ;
        RECT 60.810 197.295 61.090 197.665 ;
        RECT 60.360 195.790 60.620 196.110 ;
        RECT 60.350 195.255 60.630 195.625 ;
        RECT 60.420 190.670 60.560 195.255 ;
        RECT 60.360 190.350 60.620 190.670 ;
        RECT 60.360 189.560 60.620 189.650 ;
        RECT 60.880 189.560 61.020 197.295 ;
        RECT 60.360 189.420 61.020 189.560 ;
        RECT 60.360 189.330 60.620 189.420 ;
        RECT 60.360 185.930 60.620 186.250 ;
        RECT 57.600 181.510 57.860 181.830 ;
        RECT 57.600 179.020 57.860 179.110 ;
        RECT 58.120 179.020 58.260 185.055 ;
        RECT 59.500 185.000 60.100 185.140 ;
        RECT 58.980 184.230 59.240 184.550 ;
        RECT 59.040 181.150 59.180 184.230 ;
        RECT 59.500 181.830 59.640 185.000 ;
        RECT 60.420 184.890 60.560 185.930 ;
        RECT 60.360 184.570 60.620 184.890 ;
        RECT 59.900 184.230 60.160 184.550 ;
        RECT 59.960 184.065 60.100 184.230 ;
        RECT 59.890 183.695 60.170 184.065 ;
        RECT 60.420 183.870 60.560 184.570 ;
        RECT 60.820 184.230 61.080 184.550 ;
        RECT 59.440 181.510 59.700 181.830 ;
        RECT 58.980 180.830 59.240 181.150 ;
        RECT 59.040 179.790 59.180 180.830 ;
        RECT 58.980 179.470 59.240 179.790 ;
        RECT 59.500 179.110 59.640 181.510 ;
        RECT 59.960 180.810 60.100 183.695 ;
        RECT 60.360 183.550 60.620 183.870 ;
        RECT 60.420 181.490 60.560 183.550 ;
        RECT 60.360 181.170 60.620 181.490 ;
        RECT 59.900 180.490 60.160 180.810 ;
        RECT 57.600 178.880 58.260 179.020 ;
        RECT 57.600 178.790 57.860 178.880 ;
        RECT 59.440 178.790 59.700 179.110 ;
        RECT 56.680 177.770 56.940 178.090 ;
        RECT 57.140 177.945 57.400 178.090 ;
        RECT 57.130 177.575 57.410 177.945 ;
        RECT 56.280 175.710 56.880 175.790 ;
        RECT 56.280 175.650 56.940 175.710 ;
        RECT 55.360 175.290 56.420 175.430 ;
        RECT 56.680 175.390 56.940 175.650 ;
        RECT 53.460 174.120 54.120 174.260 ;
        RECT 53.460 174.030 53.720 174.120 ;
        RECT 54.380 174.030 54.640 174.350 ;
        RECT 55.300 173.010 55.560 173.330 ;
        RECT 54.840 171.540 55.100 171.630 ;
        RECT 55.360 171.540 55.500 173.010 ;
        RECT 54.840 171.400 55.500 171.540 ;
        RECT 54.840 171.310 55.100 171.400 ;
        RECT 52.990 170.095 53.270 170.465 ;
        RECT 56.280 170.270 56.420 175.290 ;
        RECT 59.500 174.350 59.640 178.790 ;
        RECT 59.960 176.050 60.100 180.490 ;
        RECT 59.900 175.730 60.160 176.050 ;
        RECT 60.880 174.350 61.020 184.230 ;
        RECT 61.340 181.345 61.480 198.170 ;
        RECT 61.800 197.470 61.940 199.620 ;
        RECT 62.190 199.335 62.470 199.705 ;
        RECT 62.260 198.830 62.400 199.335 ;
        RECT 62.200 198.510 62.460 198.830 ;
        RECT 62.260 197.810 62.400 198.510 ;
        RECT 62.720 198.490 62.860 200.550 ;
        RECT 63.180 198.830 63.320 202.930 ;
        RECT 63.580 200.550 63.840 200.870 ;
        RECT 63.120 198.510 63.380 198.830 ;
        RECT 62.660 198.170 62.920 198.490 ;
        RECT 62.200 197.490 62.460 197.810 ;
        RECT 61.740 197.150 62.000 197.470 ;
        RECT 61.730 196.615 62.010 196.985 ;
        RECT 61.800 192.710 61.940 196.615 ;
        RECT 62.660 195.450 62.920 195.770 ;
        RECT 62.200 195.110 62.460 195.430 ;
        RECT 61.740 192.390 62.000 192.710 ;
        RECT 61.740 189.900 62.000 189.990 ;
        RECT 62.260 189.900 62.400 195.110 ;
        RECT 62.720 194.945 62.860 195.450 ;
        RECT 62.650 194.575 62.930 194.945 ;
        RECT 62.650 193.895 62.930 194.265 ;
        RECT 62.720 190.670 62.860 193.895 ;
        RECT 62.660 190.350 62.920 190.670 ;
        RECT 61.740 189.760 62.400 189.900 ;
        RECT 61.740 189.670 62.000 189.760 ;
        RECT 61.800 187.610 61.940 189.670 ;
        RECT 61.740 187.290 62.000 187.610 ;
        RECT 63.180 182.510 63.320 198.510 ;
        RECT 63.640 196.305 63.780 200.550 ;
        RECT 64.100 200.190 64.240 202.930 ;
        RECT 64.490 201.375 64.770 201.745 ;
        RECT 64.040 199.870 64.300 200.190 ;
        RECT 64.560 198.830 64.700 201.375 ;
        RECT 64.500 198.510 64.760 198.830 ;
        RECT 63.570 195.935 63.850 196.305 ;
        RECT 64.560 195.770 64.700 198.510 ;
        RECT 65.020 197.130 65.160 202.930 ;
        RECT 65.410 202.735 65.690 203.105 ;
        RECT 65.480 197.810 65.620 202.735 ;
        RECT 65.880 202.250 66.140 202.570 ;
        RECT 65.940 201.550 66.080 202.250 ;
        RECT 65.880 201.230 66.140 201.550 ;
        RECT 66.330 201.375 66.610 201.745 ;
        RECT 65.870 200.695 66.150 201.065 ;
        RECT 66.400 200.870 66.540 201.375 ;
        RECT 65.880 200.550 66.140 200.695 ;
        RECT 66.340 200.550 66.600 200.870 ;
        RECT 65.420 197.490 65.680 197.810 ;
        RECT 64.960 196.810 65.220 197.130 ;
        RECT 64.500 195.450 64.760 195.770 ;
        RECT 65.020 195.000 65.160 196.810 ;
        RECT 65.480 196.110 65.620 197.490 ;
        RECT 65.420 195.790 65.680 196.110 ;
        RECT 65.940 195.510 66.080 200.550 ;
        RECT 66.330 200.015 66.610 200.385 ;
        RECT 66.400 198.830 66.540 200.015 ;
        RECT 66.860 198.830 67.000 204.970 ;
        RECT 67.260 203.610 67.520 203.930 ;
        RECT 67.320 201.550 67.460 203.610 ;
        RECT 67.780 202.425 67.920 206.080 ;
        RECT 67.710 202.055 67.990 202.425 ;
        RECT 67.260 201.230 67.520 201.550 ;
        RECT 68.240 200.870 68.380 207.690 ;
        RECT 68.700 206.990 68.840 207.780 ;
        RECT 69.100 207.690 69.360 207.780 ;
        RECT 68.640 206.670 68.900 206.990 ;
        RECT 68.180 200.550 68.440 200.870 ;
        RECT 68.700 199.850 68.840 206.670 ;
        RECT 69.620 206.310 69.760 209.390 ;
        RECT 70.020 208.370 70.280 208.690 ;
        RECT 69.560 205.990 69.820 206.310 ;
        RECT 69.100 204.970 69.360 205.290 ;
        RECT 69.160 203.930 69.300 204.970 ;
        RECT 69.560 203.950 69.820 204.270 ;
        RECT 69.100 203.610 69.360 203.930 ;
        RECT 69.160 201.210 69.300 203.610 ;
        RECT 69.620 203.105 69.760 203.950 ;
        RECT 70.080 203.160 70.220 208.370 ;
        RECT 70.540 206.990 70.680 211.430 ;
        RECT 71.460 209.710 71.600 211.430 ;
        RECT 73.240 210.750 73.500 211.070 ;
        RECT 71.400 209.390 71.660 209.710 ;
        RECT 70.940 208.545 71.200 208.690 ;
        RECT 70.930 208.175 71.210 208.545 ;
        RECT 71.460 208.430 71.600 209.390 ;
        RECT 71.860 208.940 72.120 209.030 ;
        RECT 72.780 208.940 73.040 209.030 ;
        RECT 71.860 208.800 73.040 208.940 ;
        RECT 71.860 208.710 72.120 208.800 ;
        RECT 72.780 208.710 73.040 208.800 ;
        RECT 71.460 208.290 72.520 208.430 ;
        RECT 70.940 207.690 71.200 208.010 ;
        RECT 71.400 207.690 71.660 208.010 ;
        RECT 70.480 206.670 70.740 206.990 ;
        RECT 71.000 206.310 71.140 207.690 ;
        RECT 71.460 206.650 71.600 207.690 ;
        RECT 71.400 206.330 71.660 206.650 ;
        RECT 70.480 205.990 70.740 206.310 ;
        RECT 70.940 205.990 71.200 206.310 ;
        RECT 70.540 204.465 70.680 205.990 ;
        RECT 70.470 204.095 70.750 204.465 ;
        RECT 71.000 204.270 71.140 205.990 ;
        RECT 72.380 204.270 72.520 208.290 ;
        RECT 72.840 206.310 72.980 208.710 ;
        RECT 72.780 205.990 73.040 206.310 ;
        RECT 70.940 203.950 71.200 204.270 ;
        RECT 72.320 203.950 72.580 204.270 ;
        RECT 72.770 204.095 73.050 204.465 ;
        RECT 72.840 203.930 72.980 204.095 ;
        RECT 70.940 203.270 71.200 203.590 ;
        RECT 71.390 203.415 71.670 203.785 ;
        RECT 72.780 203.610 73.040 203.930 ;
        RECT 69.550 202.735 69.830 203.105 ;
        RECT 70.080 203.020 70.680 203.160 ;
        RECT 70.010 202.055 70.290 202.425 ;
        RECT 69.100 200.890 69.360 201.210 ;
        RECT 70.080 200.870 70.220 202.055 ;
        RECT 70.020 200.550 70.280 200.870 ;
        RECT 70.080 200.385 70.220 200.550 ;
        RECT 70.010 200.015 70.290 200.385 ;
        RECT 68.180 199.530 68.440 199.850 ;
        RECT 68.640 199.530 68.900 199.850 ;
        RECT 66.340 198.510 66.600 198.830 ;
        RECT 66.800 198.510 67.060 198.830 ;
        RECT 67.250 195.935 67.530 196.305 ;
        RECT 67.320 195.770 67.460 195.935 ;
        RECT 67.260 195.680 67.520 195.770 ;
        RECT 64.560 194.860 65.160 195.000 ;
        RECT 65.480 195.370 66.080 195.510 ;
        RECT 66.860 195.540 67.520 195.680 ;
        RECT 64.040 194.430 64.300 194.750 ;
        RECT 63.580 194.265 63.840 194.410 ;
        RECT 63.570 193.895 63.850 194.265 ;
        RECT 63.570 192.535 63.850 192.905 ;
        RECT 64.100 192.710 64.240 194.430 ;
        RECT 63.640 190.670 63.780 192.535 ;
        RECT 64.040 192.390 64.300 192.710 ;
        RECT 64.040 191.370 64.300 191.690 ;
        RECT 63.580 190.350 63.840 190.670 ;
        RECT 63.640 189.990 63.780 190.350 ;
        RECT 64.100 189.990 64.240 191.370 ;
        RECT 63.580 189.670 63.840 189.990 ;
        RECT 64.040 189.670 64.300 189.990 ;
        RECT 64.560 184.550 64.700 194.860 ;
        RECT 64.960 194.090 65.220 194.410 ;
        RECT 65.020 190.330 65.160 194.090 ;
        RECT 65.480 192.790 65.620 195.370 ;
        RECT 66.340 195.110 66.600 195.430 ;
        RECT 65.880 194.770 66.140 195.090 ;
        RECT 65.940 193.390 66.080 194.770 ;
        RECT 65.880 193.070 66.140 193.390 ;
        RECT 65.480 192.650 66.080 192.790 ;
        RECT 65.410 190.495 65.690 190.865 ;
        RECT 65.420 190.350 65.680 190.495 ;
        RECT 64.960 190.010 65.220 190.330 ;
        RECT 65.410 189.815 65.690 190.185 ;
        RECT 65.480 188.970 65.620 189.815 ;
        RECT 65.420 188.650 65.680 188.970 ;
        RECT 64.500 184.230 64.760 184.550 ;
        RECT 65.420 184.230 65.680 184.550 ;
        RECT 63.120 182.190 63.380 182.510 ;
        RECT 61.270 180.975 61.550 181.345 ;
        RECT 61.740 180.490 62.000 180.810 ;
        RECT 64.040 180.490 64.300 180.810 ;
        RECT 61.800 176.050 61.940 180.490 ;
        RECT 64.100 179.790 64.240 180.490 ;
        RECT 64.040 179.470 64.300 179.790 ;
        RECT 63.120 178.450 63.380 178.770 ;
        RECT 63.180 177.070 63.320 178.450 ;
        RECT 64.560 178.090 64.700 184.230 ;
        RECT 65.480 182.510 65.620 184.230 ;
        RECT 65.420 182.190 65.680 182.510 ;
        RECT 65.940 181.490 66.080 192.650 ;
        RECT 66.400 190.185 66.540 195.110 ;
        RECT 66.860 191.545 67.000 195.540 ;
        RECT 67.260 195.450 67.520 195.540 ;
        RECT 68.240 195.430 68.380 199.530 ;
        RECT 70.010 199.335 70.290 199.705 ;
        RECT 70.080 197.470 70.220 199.335 ;
        RECT 70.020 197.150 70.280 197.470 ;
        RECT 70.020 195.680 70.280 195.770 ;
        RECT 69.160 195.540 70.280 195.680 ;
        RECT 68.180 195.110 68.440 195.430 ;
        RECT 68.180 192.730 68.440 193.050 ;
        RECT 66.790 191.175 67.070 191.545 ;
        RECT 67.720 191.370 67.980 191.690 ;
        RECT 68.240 191.545 68.380 192.730 ;
        RECT 68.640 191.710 68.900 192.030 ;
        RECT 66.330 189.815 66.610 190.185 ;
        RECT 67.780 189.990 67.920 191.370 ;
        RECT 68.170 191.175 68.450 191.545 ;
        RECT 67.720 189.900 67.980 189.990 ;
        RECT 67.320 189.760 67.980 189.900 ;
        RECT 67.320 186.590 67.460 189.760 ;
        RECT 67.720 189.670 67.980 189.760 ;
        RECT 68.180 189.670 68.440 189.990 ;
        RECT 67.710 187.095 67.990 187.465 ;
        RECT 67.720 186.950 67.980 187.095 ;
        RECT 67.260 186.270 67.520 186.590 ;
        RECT 66.800 183.550 67.060 183.870 ;
        RECT 66.340 183.210 66.600 183.530 ;
        RECT 65.880 181.170 66.140 181.490 ;
        RECT 65.940 179.450 66.080 181.170 ;
        RECT 66.400 179.790 66.540 183.210 ;
        RECT 66.860 179.790 67.000 183.550 ;
        RECT 66.340 179.470 66.600 179.790 ;
        RECT 66.800 179.470 67.060 179.790 ;
        RECT 67.320 179.450 67.460 186.270 ;
        RECT 68.240 185.230 68.380 189.670 ;
        RECT 68.700 189.505 68.840 191.710 ;
        RECT 69.160 190.865 69.300 195.540 ;
        RECT 70.020 195.450 70.280 195.540 ;
        RECT 70.020 192.730 70.280 193.050 ;
        RECT 69.560 192.050 69.820 192.370 ;
        RECT 69.090 190.495 69.370 190.865 ;
        RECT 69.100 189.670 69.360 189.990 ;
        RECT 68.630 189.135 68.910 189.505 ;
        RECT 69.160 185.310 69.300 189.670 ;
        RECT 69.620 188.145 69.760 192.050 ;
        RECT 70.080 189.990 70.220 192.730 ;
        RECT 70.540 189.990 70.680 203.020 ;
        RECT 71.000 201.745 71.140 203.270 ;
        RECT 70.930 201.375 71.210 201.745 ;
        RECT 71.460 201.550 71.600 203.415 ;
        RECT 71.860 202.250 72.120 202.570 ;
        RECT 71.400 201.230 71.660 201.550 ;
        RECT 71.920 201.210 72.060 202.250 ;
        RECT 72.780 201.230 73.040 201.550 ;
        RECT 71.860 200.890 72.120 201.210 ;
        RECT 70.930 200.015 71.210 200.385 ;
        RECT 71.000 198.490 71.140 200.015 ;
        RECT 70.940 198.170 71.200 198.490 ;
        RECT 71.400 197.490 71.660 197.810 ;
        RECT 72.320 197.720 72.580 197.810 ;
        RECT 72.840 197.720 72.980 201.230 ;
        RECT 73.300 198.150 73.440 210.750 ;
        RECT 76.060 209.710 76.200 216.870 ;
        RECT 76.460 213.130 76.720 213.450 ;
        RECT 76.520 211.750 76.660 213.130 ;
        RECT 76.980 212.430 77.120 217.210 ;
        RECT 77.840 213.810 78.100 214.130 ;
        RECT 76.920 212.110 77.180 212.430 ;
        RECT 76.460 211.430 76.720 211.750 ;
        RECT 77.380 211.430 77.640 211.750 ;
        RECT 76.910 210.895 77.190 211.265 ;
        RECT 75.540 209.390 75.800 209.710 ;
        RECT 76.000 209.390 76.260 209.710 ;
        RECT 76.980 209.620 77.120 210.895 ;
        RECT 77.440 210.730 77.580 211.430 ;
        RECT 77.380 210.410 77.640 210.730 ;
        RECT 77.380 209.620 77.640 209.710 ;
        RECT 76.980 209.480 77.640 209.620 ;
        RECT 77.380 209.390 77.640 209.480 ;
        RECT 75.600 209.110 75.740 209.390 ;
        RECT 75.600 208.970 76.660 209.110 ;
        RECT 73.700 208.370 73.960 208.690 ;
        RECT 73.760 205.970 73.900 208.370 ;
        RECT 76.000 208.030 76.260 208.350 ;
        RECT 74.160 206.670 74.420 206.990 ;
        RECT 74.220 205.970 74.360 206.670 ;
        RECT 74.620 206.330 74.880 206.650 ;
        RECT 73.700 205.650 73.960 205.970 ;
        RECT 74.160 205.650 74.420 205.970 ;
        RECT 74.220 205.290 74.360 205.650 ;
        RECT 74.160 204.970 74.420 205.290 ;
        RECT 73.690 202.735 73.970 203.105 ;
        RECT 73.240 197.830 73.500 198.150 ;
        RECT 72.320 197.580 72.980 197.720 ;
        RECT 72.320 197.490 72.580 197.580 ;
        RECT 71.460 195.625 71.600 197.490 ;
        RECT 71.390 195.255 71.670 195.625 ;
        RECT 71.400 194.770 71.660 195.090 ;
        RECT 70.940 192.050 71.200 192.370 ;
        RECT 71.000 190.670 71.140 192.050 ;
        RECT 70.940 190.350 71.200 190.670 ;
        RECT 71.460 190.070 71.600 194.770 ;
        RECT 72.320 194.090 72.580 194.410 ;
        RECT 72.380 192.370 72.520 194.090 ;
        RECT 72.840 193.390 72.980 197.580 ;
        RECT 73.240 195.790 73.500 196.110 ;
        RECT 72.780 193.070 73.040 193.390 ;
        RECT 72.320 192.050 72.580 192.370 ;
        RECT 70.020 189.670 70.280 189.990 ;
        RECT 70.480 189.670 70.740 189.990 ;
        RECT 71.000 189.930 71.600 190.070 ;
        RECT 71.000 189.650 71.140 189.930 ;
        RECT 72.320 189.900 72.580 189.990 ;
        RECT 71.920 189.760 72.580 189.900 ;
        RECT 70.940 189.330 71.200 189.650 ;
        RECT 71.400 189.330 71.660 189.650 ;
        RECT 69.550 187.775 69.830 188.145 ;
        RECT 69.620 186.930 69.760 187.775 ;
        RECT 71.460 187.270 71.600 189.330 ;
        RECT 71.400 186.950 71.660 187.270 ;
        RECT 69.560 186.610 69.820 186.930 ;
        RECT 71.400 186.270 71.660 186.590 ;
        RECT 68.180 184.910 68.440 185.230 ;
        RECT 69.160 185.170 70.220 185.310 ;
        RECT 69.560 184.570 69.820 184.890 ;
        RECT 68.180 184.460 68.440 184.550 ;
        RECT 69.100 184.460 69.360 184.550 ;
        RECT 68.180 184.320 69.360 184.460 ;
        RECT 68.180 184.230 68.440 184.320 ;
        RECT 69.100 184.230 69.360 184.320 ;
        RECT 67.710 183.015 67.990 183.385 ;
        RECT 65.880 179.130 66.140 179.450 ;
        RECT 67.260 179.130 67.520 179.450 ;
        RECT 64.500 177.770 64.760 178.090 ;
        RECT 63.120 176.750 63.380 177.070 ;
        RECT 63.570 176.895 63.850 177.265 ;
        RECT 62.200 176.585 62.460 176.730 ;
        RECT 62.190 176.215 62.470 176.585 ;
        RECT 61.740 175.730 62.000 176.050 ;
        RECT 59.440 174.030 59.700 174.350 ;
        RECT 60.820 174.030 61.080 174.350 ;
        RECT 61.270 174.175 61.550 174.545 ;
        RECT 61.340 173.670 61.480 174.175 ;
        RECT 63.640 173.670 63.780 176.895 ;
        RECT 67.780 176.730 67.920 183.015 ;
        RECT 68.180 179.470 68.440 179.790 ;
        RECT 68.240 178.430 68.380 179.470 ;
        RECT 68.180 178.110 68.440 178.430 ;
        RECT 67.720 176.410 67.980 176.730 ;
        RECT 68.240 176.050 68.380 178.110 ;
        RECT 68.180 175.730 68.440 176.050 ;
        RECT 66.800 175.050 67.060 175.370 ;
        RECT 67.720 175.050 67.980 175.370 ;
        RECT 68.180 175.050 68.440 175.370 ;
        RECT 66.860 173.670 67.000 175.050 ;
        RECT 57.140 173.580 57.400 173.670 ;
        RECT 58.060 173.580 58.320 173.670 ;
        RECT 57.140 173.440 58.320 173.580 ;
        RECT 57.140 173.350 57.400 173.440 ;
        RECT 58.060 173.350 58.320 173.440 ;
        RECT 61.280 173.350 61.540 173.670 ;
        RECT 63.580 173.350 63.840 173.670 ;
        RECT 66.800 173.350 67.060 173.670 ;
        RECT 58.980 172.670 59.240 172.990 ;
        RECT 59.040 170.610 59.180 172.670 ;
        RECT 62.660 172.330 62.920 172.650 ;
        RECT 62.720 170.610 62.860 172.330 ;
        RECT 66.860 170.950 67.000 173.350 ;
        RECT 67.780 172.990 67.920 175.050 ;
        RECT 68.240 174.010 68.380 175.050 ;
        RECT 68.630 174.855 68.910 175.225 ;
        RECT 68.180 173.690 68.440 174.010 ;
        RECT 67.720 172.670 67.980 172.990 ;
        RECT 68.700 171.630 68.840 174.855 ;
        RECT 69.160 174.010 69.300 184.230 ;
        RECT 69.620 183.870 69.760 184.570 ;
        RECT 69.560 183.550 69.820 183.870 ;
        RECT 69.620 181.490 69.760 183.550 ;
        RECT 69.560 181.170 69.820 181.490 ;
        RECT 69.560 180.490 69.820 180.810 ;
        RECT 69.620 176.390 69.760 180.490 ;
        RECT 69.560 176.070 69.820 176.390 ;
        RECT 70.080 175.370 70.220 185.170 ;
        RECT 71.460 181.830 71.600 186.270 ;
        RECT 71.920 185.230 72.060 189.760 ;
        RECT 72.320 189.670 72.580 189.760 ;
        RECT 71.860 184.910 72.120 185.230 ;
        RECT 72.840 184.550 72.980 193.070 ;
        RECT 73.300 192.370 73.440 195.790 ;
        RECT 73.760 192.370 73.900 202.735 ;
        RECT 74.220 197.470 74.360 204.970 ;
        RECT 74.680 203.930 74.820 206.330 ;
        RECT 76.060 206.310 76.200 208.030 ;
        RECT 76.520 206.990 76.660 208.970 ;
        RECT 77.380 208.710 77.640 209.030 ;
        RECT 76.920 208.370 77.180 208.690 ;
        RECT 76.460 206.670 76.720 206.990 ;
        RECT 76.520 206.310 76.660 206.670 ;
        RECT 76.980 206.310 77.120 208.370 ;
        RECT 76.000 205.990 76.260 206.310 ;
        RECT 76.460 205.990 76.720 206.310 ;
        RECT 76.920 205.990 77.180 206.310 ;
        RECT 75.080 204.970 75.340 205.290 ;
        RECT 75.140 204.270 75.280 204.970 ;
        RECT 75.080 203.950 75.340 204.270 ;
        RECT 75.540 203.950 75.800 204.270 ;
        RECT 74.620 203.610 74.880 203.930 ;
        RECT 75.600 203.590 75.740 203.950 ;
        RECT 75.540 203.270 75.800 203.590 ;
        RECT 74.620 202.590 74.880 202.910 ;
        RECT 75.540 202.590 75.800 202.910 ;
        RECT 74.680 202.310 74.820 202.590 ;
        RECT 74.680 202.170 75.280 202.310 ;
        RECT 74.620 200.550 74.880 200.870 ;
        RECT 74.680 199.850 74.820 200.550 ;
        RECT 75.140 200.530 75.280 202.170 ;
        RECT 75.600 201.210 75.740 202.590 ;
        RECT 75.540 200.890 75.800 201.210 ;
        RECT 75.080 200.210 75.340 200.530 ;
        RECT 74.620 199.530 74.880 199.850 ;
        RECT 74.680 197.810 74.820 199.530 ;
        RECT 74.620 197.490 74.880 197.810 ;
        RECT 75.080 197.490 75.340 197.810 ;
        RECT 74.160 197.150 74.420 197.470 ;
        RECT 74.160 194.430 74.420 194.750 ;
        RECT 73.240 192.050 73.500 192.370 ;
        RECT 73.700 192.050 73.960 192.370 ;
        RECT 72.320 184.230 72.580 184.550 ;
        RECT 72.780 184.230 73.040 184.550 ;
        RECT 71.860 183.210 72.120 183.530 ;
        RECT 71.400 181.510 71.660 181.830 ;
        RECT 70.940 180.830 71.200 181.150 ;
        RECT 70.480 179.470 70.740 179.790 ;
        RECT 70.540 175.710 70.680 179.470 ;
        RECT 71.000 179.110 71.140 180.830 ;
        RECT 71.920 179.790 72.060 183.210 ;
        RECT 72.380 182.510 72.520 184.230 ;
        RECT 72.840 182.510 72.980 184.230 ;
        RECT 72.320 182.190 72.580 182.510 ;
        RECT 72.780 182.190 73.040 182.510 ;
        RECT 71.860 179.470 72.120 179.790 ;
        RECT 72.780 179.470 73.040 179.790 ;
        RECT 70.940 178.790 71.200 179.110 ;
        RECT 71.850 178.935 72.130 179.305 ;
        RECT 72.840 179.110 72.980 179.470 ;
        RECT 73.300 179.190 73.440 192.050 ;
        RECT 74.220 189.650 74.360 194.430 ;
        RECT 75.140 192.225 75.280 197.490 ;
        RECT 75.600 197.470 75.740 200.890 ;
        RECT 76.060 200.190 76.200 205.990 ;
        RECT 76.460 204.970 76.720 205.290 ;
        RECT 76.520 201.550 76.660 204.970 ;
        RECT 76.460 201.230 76.720 201.550 ;
        RECT 76.460 200.550 76.720 200.870 ;
        RECT 76.000 199.870 76.260 200.190 ;
        RECT 76.520 197.665 76.660 200.550 ;
        RECT 76.980 200.530 77.120 205.990 ;
        RECT 76.920 200.210 77.180 200.530 ;
        RECT 76.920 197.830 77.180 198.150 ;
        RECT 75.540 197.150 75.800 197.470 ;
        RECT 76.450 197.295 76.730 197.665 ;
        RECT 76.520 197.130 76.660 197.295 ;
        RECT 75.990 196.615 76.270 196.985 ;
        RECT 76.460 196.810 76.720 197.130 ;
        RECT 76.060 195.770 76.200 196.615 ;
        RECT 76.980 196.110 77.120 197.830 ;
        RECT 76.920 196.020 77.180 196.110 ;
        RECT 76.520 195.880 77.180 196.020 ;
        RECT 75.540 195.450 75.800 195.770 ;
        RECT 76.000 195.450 76.260 195.770 ;
        RECT 75.600 192.710 75.740 195.450 ;
        RECT 75.540 192.390 75.800 192.710 ;
        RECT 75.070 191.855 75.350 192.225 ;
        RECT 75.530 191.175 75.810 191.545 ;
        RECT 75.600 190.330 75.740 191.175 ;
        RECT 75.540 190.010 75.800 190.330 ;
        RECT 76.060 189.990 76.200 195.450 ;
        RECT 74.620 189.670 74.880 189.990 ;
        RECT 76.000 189.670 76.260 189.990 ;
        RECT 74.160 189.330 74.420 189.650 ;
        RECT 73.690 188.455 73.970 188.825 ;
        RECT 73.760 186.930 73.900 188.455 ;
        RECT 73.700 186.610 73.960 186.930 ;
        RECT 73.760 184.210 73.900 186.610 ;
        RECT 73.700 183.890 73.960 184.210 ;
        RECT 71.860 178.790 72.120 178.935 ;
        RECT 72.780 178.790 73.040 179.110 ;
        RECT 73.300 179.050 74.360 179.190 ;
        RECT 71.000 176.390 71.140 178.790 ;
        RECT 73.240 178.450 73.500 178.770 ;
        RECT 73.300 177.070 73.440 178.450 ;
        RECT 73.700 177.770 73.960 178.090 ;
        RECT 73.240 176.750 73.500 177.070 ;
        RECT 70.940 176.070 71.200 176.390 ;
        RECT 71.850 176.215 72.130 176.585 ;
        RECT 70.480 175.390 70.740 175.710 ;
        RECT 70.020 175.050 70.280 175.370 ;
        RECT 71.400 175.050 71.660 175.370 ;
        RECT 69.100 173.690 69.360 174.010 ;
        RECT 69.160 172.650 69.300 173.690 ;
        RECT 71.460 173.670 71.600 175.050 ;
        RECT 71.920 173.670 72.060 176.215 ;
        RECT 73.760 174.350 73.900 177.770 ;
        RECT 73.700 174.030 73.960 174.350 ;
        RECT 71.400 173.350 71.660 173.670 ;
        RECT 71.860 173.350 72.120 173.670 ;
        RECT 74.220 173.330 74.360 179.050 ;
        RECT 74.680 178.770 74.820 189.670 ;
        RECT 76.520 181.830 76.660 195.880 ;
        RECT 76.920 195.790 77.180 195.880 ;
        RECT 76.920 192.390 77.180 192.710 ;
        RECT 76.980 190.865 77.120 192.390 ;
        RECT 76.910 190.495 77.190 190.865 ;
        RECT 77.440 186.785 77.580 208.710 ;
        RECT 77.900 208.690 78.040 213.810 ;
        RECT 79.740 212.090 79.880 222.990 ;
        RECT 82.440 220.270 82.700 220.590 ;
        RECT 81.060 217.890 81.320 218.210 ;
        RECT 81.120 212.430 81.260 217.890 ;
        RECT 81.980 214.150 82.240 214.470 ;
        RECT 81.060 212.110 81.320 212.430 ;
        RECT 79.680 211.770 79.940 212.090 ;
        RECT 82.040 211.750 82.180 214.150 ;
        RECT 82.500 212.430 82.640 220.270 ;
        RECT 83.880 212.430 84.020 223.135 ;
        RECT 92.100 215.170 92.360 215.490 ;
        RECT 84.740 214.490 85.000 214.810 ;
        RECT 82.440 212.110 82.700 212.430 ;
        RECT 83.820 212.110 84.080 212.430 ;
        RECT 84.800 211.750 84.940 214.490 ;
        RECT 89.790 214.295 90.070 214.665 ;
        RECT 89.860 212.430 90.000 214.295 ;
        RECT 89.800 212.110 90.060 212.430 ;
        RECT 92.160 212.090 92.300 215.170 ;
        RECT 92.100 211.770 92.360 212.090 ;
        RECT 81.980 211.430 82.240 211.750 ;
        RECT 84.740 211.430 85.000 211.750 ;
        RECT 82.440 211.090 82.700 211.410 ;
        RECT 81.510 210.215 81.790 210.585 ;
        RECT 78.300 209.620 78.560 209.710 ;
        RECT 78.300 209.480 79.420 209.620 ;
        RECT 80.590 209.535 80.870 209.905 ;
        RECT 78.300 209.390 78.560 209.480 ;
        RECT 78.290 208.855 78.570 209.225 ;
        RECT 79.280 209.030 79.420 209.480 ;
        RECT 78.360 208.690 78.500 208.855 ;
        RECT 79.220 208.710 79.480 209.030 ;
        RECT 80.660 208.690 80.800 209.535 ;
        RECT 77.840 208.370 78.100 208.690 ;
        RECT 78.300 208.370 78.560 208.690 ;
        RECT 80.600 208.370 80.860 208.690 ;
        RECT 77.840 207.690 78.100 208.010 ;
        RECT 78.760 207.690 79.020 208.010 ;
        RECT 77.900 205.290 78.040 207.690 ;
        RECT 77.840 204.970 78.100 205.290 ;
        RECT 77.840 202.590 78.100 202.910 ;
        RECT 77.900 201.550 78.040 202.590 ;
        RECT 77.840 201.230 78.100 201.550 ;
        RECT 78.300 199.530 78.560 199.850 ;
        RECT 78.360 198.150 78.500 199.530 ;
        RECT 78.300 197.830 78.560 198.150 ;
        RECT 78.360 195.430 78.500 197.830 ;
        RECT 78.300 195.110 78.560 195.430 ;
        RECT 77.840 194.770 78.100 195.090 ;
        RECT 78.820 194.945 78.960 207.690 ;
        RECT 80.140 206.330 80.400 206.650 ;
        RECT 80.200 204.270 80.340 206.330 ;
        RECT 80.600 205.650 80.860 205.970 ;
        RECT 80.140 203.950 80.400 204.270 ;
        RECT 80.660 203.670 80.800 205.650 ;
        RECT 81.060 204.970 81.320 205.290 ;
        RECT 79.280 203.530 80.800 203.670 ;
        RECT 77.900 194.265 78.040 194.770 ;
        RECT 78.750 194.575 79.030 194.945 ;
        RECT 77.830 193.895 78.110 194.265 ;
        RECT 78.300 194.090 78.560 194.410 ;
        RECT 77.900 192.110 78.040 193.895 ;
        RECT 78.360 192.710 78.500 194.090 ;
        RECT 79.280 193.390 79.420 203.530 ;
        RECT 79.680 195.450 79.940 195.770 ;
        RECT 79.740 193.390 79.880 195.450 ;
        RECT 80.140 195.110 80.400 195.430 ;
        RECT 80.200 194.320 80.340 195.110 ;
        RECT 80.600 194.320 80.860 194.410 ;
        RECT 80.200 194.180 80.860 194.320 ;
        RECT 79.220 193.070 79.480 193.390 ;
        RECT 79.680 193.070 79.940 193.390 ;
        RECT 78.760 192.730 79.020 193.050 ;
        RECT 80.200 192.790 80.340 194.180 ;
        RECT 80.600 194.090 80.860 194.180 ;
        RECT 78.300 192.390 78.560 192.710 ;
        RECT 77.900 191.970 78.500 192.110 ;
        RECT 77.830 191.175 78.110 191.545 ;
        RECT 77.370 186.415 77.650 186.785 ;
        RECT 76.460 181.510 76.720 181.830 ;
        RECT 75.080 181.170 75.340 181.490 ;
        RECT 75.140 179.790 75.280 181.170 ;
        RECT 76.520 179.790 76.660 181.510 ;
        RECT 75.080 179.470 75.340 179.790 ;
        RECT 75.540 179.470 75.800 179.790 ;
        RECT 76.460 179.470 76.720 179.790 ;
        RECT 74.620 178.450 74.880 178.770 ;
        RECT 74.680 175.370 74.820 178.450 ;
        RECT 75.080 176.410 75.340 176.730 ;
        RECT 74.620 175.050 74.880 175.370 ;
        RECT 75.140 173.670 75.280 176.410 ;
        RECT 75.600 174.350 75.740 179.470 ;
        RECT 77.900 179.110 78.040 191.175 ;
        RECT 78.360 183.385 78.500 191.970 ;
        RECT 78.820 190.330 78.960 192.730 ;
        RECT 79.740 192.650 80.340 192.790 ;
        RECT 79.220 191.370 79.480 191.690 ;
        RECT 79.740 191.545 79.880 192.650 ;
        RECT 80.600 192.050 80.860 192.370 ;
        RECT 79.280 190.580 79.420 191.370 ;
        RECT 79.670 191.175 79.950 191.545 ;
        RECT 80.140 191.370 80.400 191.690 ;
        RECT 79.680 190.580 79.940 190.670 ;
        RECT 79.280 190.440 79.940 190.580 ;
        RECT 79.680 190.350 79.940 190.440 ;
        RECT 78.760 190.010 79.020 190.330 ;
        RECT 78.760 189.330 79.020 189.650 ;
        RECT 78.290 183.015 78.570 183.385 ;
        RECT 77.840 178.790 78.100 179.110 ;
        RECT 78.300 178.790 78.560 179.110 ;
        RECT 78.360 176.050 78.500 178.790 ;
        RECT 78.820 176.390 78.960 189.330 ;
        RECT 79.680 186.950 79.940 187.270 ;
        RECT 79.220 183.890 79.480 184.210 ;
        RECT 79.280 181.150 79.420 183.890 ;
        RECT 79.220 180.830 79.480 181.150 ;
        RECT 79.280 179.305 79.420 180.830 ;
        RECT 79.210 178.935 79.490 179.305 ;
        RECT 79.740 178.510 79.880 186.950 ;
        RECT 80.200 179.110 80.340 191.370 ;
        RECT 80.660 190.670 80.800 192.050 ;
        RECT 80.600 190.350 80.860 190.670 ;
        RECT 80.600 188.990 80.860 189.310 ;
        RECT 80.660 186.930 80.800 188.990 ;
        RECT 80.600 186.610 80.860 186.930 ;
        RECT 80.600 184.460 80.860 184.550 ;
        RECT 81.120 184.460 81.260 204.970 ;
        RECT 81.580 196.305 81.720 210.215 ;
        RECT 82.500 208.690 82.640 211.090 ;
        RECT 88.420 210.750 88.680 211.070 ;
        RECT 90.260 210.750 90.520 211.070 ;
        RECT 88.480 210.585 88.620 210.750 ;
        RECT 88.410 210.215 88.690 210.585 ;
        RECT 86.580 209.620 86.840 209.710 ;
        RECT 86.580 209.480 87.240 209.620 ;
        RECT 86.580 209.390 86.840 209.480 ;
        RECT 81.980 208.370 82.240 208.690 ;
        RECT 82.440 208.370 82.700 208.690 ;
        RECT 82.040 208.010 82.180 208.370 ;
        RECT 85.200 208.030 85.460 208.350 ;
        RECT 81.980 207.690 82.240 208.010 ;
        RECT 83.820 207.690 84.080 208.010 ;
        RECT 82.040 205.825 82.180 207.690 ;
        RECT 83.880 206.990 84.020 207.690 ;
        RECT 83.820 206.670 84.080 206.990 ;
        RECT 82.900 205.990 83.160 206.310 ;
        RECT 81.970 205.455 82.250 205.825 ;
        RECT 81.980 204.970 82.240 205.290 ;
        RECT 82.960 205.145 83.100 205.990 ;
        RECT 81.510 195.935 81.790 196.305 ;
        RECT 81.520 195.450 81.780 195.770 ;
        RECT 81.580 194.750 81.720 195.450 ;
        RECT 82.040 195.430 82.180 204.970 ;
        RECT 82.890 204.775 83.170 205.145 ;
        RECT 83.880 203.250 84.020 206.670 ;
        RECT 85.260 206.310 85.400 208.030 ;
        RECT 85.200 205.990 85.460 206.310 ;
        RECT 86.120 205.990 86.380 206.310 ;
        RECT 85.260 203.250 85.400 205.990 ;
        RECT 86.180 205.145 86.320 205.990 ;
        RECT 86.110 204.775 86.390 205.145 ;
        RECT 85.660 203.785 85.920 203.930 ;
        RECT 85.650 203.415 85.930 203.785 ;
        RECT 86.180 203.250 86.320 204.775 ;
        RECT 87.100 204.270 87.240 209.480 ;
        RECT 87.960 209.390 88.220 209.710 ;
        RECT 88.020 208.690 88.160 209.390 ;
        RECT 89.340 208.710 89.600 209.030 ;
        RECT 87.960 208.370 88.220 208.690 ;
        RECT 89.400 208.545 89.540 208.710 ;
        RECT 90.320 208.690 90.460 210.750 ;
        RECT 91.640 210.410 91.900 210.730 ;
        RECT 91.700 209.030 91.840 210.410 ;
        RECT 91.180 208.710 91.440 209.030 ;
        RECT 91.640 208.710 91.900 209.030 ;
        RECT 89.330 208.175 89.610 208.545 ;
        RECT 90.260 208.370 90.520 208.690 ;
        RECT 91.240 207.920 91.380 208.710 ;
        RECT 92.160 208.690 92.300 211.770 ;
        RECT 93.540 211.750 93.680 223.160 ;
        RECT 96.760 212.090 96.900 223.160 ;
        RECT 96.700 211.770 96.960 212.090 ;
        RECT 103.200 211.750 103.340 223.160 ;
        RECT 106.420 217.270 106.560 223.160 ;
        RECT 105.960 217.130 106.560 217.270 ;
        RECT 105.960 211.750 106.100 217.130 ;
        RECT 106.570 212.595 108.110 212.965 ;
        RECT 109.640 211.750 109.780 223.160 ;
        RECT 112.860 211.750 113.000 223.160 ;
        RECT 93.480 211.430 93.740 211.750 ;
        RECT 95.780 211.430 96.040 211.750 ;
        RECT 103.140 211.430 103.400 211.750 ;
        RECT 105.900 211.430 106.160 211.750 ;
        RECT 109.580 211.430 109.840 211.750 ;
        RECT 112.800 211.430 113.060 211.750 ;
        RECT 93.020 211.090 93.280 211.410 ;
        RECT 92.100 208.370 92.360 208.690 ;
        RECT 93.080 207.920 93.220 211.090 ;
        RECT 94.860 210.410 95.120 210.730 ;
        RECT 95.320 210.410 95.580 210.730 ;
        RECT 93.940 208.030 94.200 208.350 ;
        RECT 94.390 208.175 94.670 208.545 ;
        RECT 91.240 207.780 93.220 207.920 ;
        RECT 87.500 205.990 87.760 206.310 ;
        RECT 88.880 206.220 89.140 206.310 ;
        RECT 89.800 206.220 90.060 206.310 ;
        RECT 91.640 206.220 91.900 206.310 ;
        RECT 88.880 206.080 91.900 206.220 ;
        RECT 88.880 205.990 89.140 206.080 ;
        RECT 89.800 205.990 90.060 206.080 ;
        RECT 91.640 205.990 91.900 206.080 ;
        RECT 87.040 203.950 87.300 204.270 ;
        RECT 83.820 202.930 84.080 203.250 ;
        RECT 85.200 202.930 85.460 203.250 ;
        RECT 86.120 202.930 86.380 203.250 ;
        RECT 87.040 202.590 87.300 202.910 ;
        RECT 87.100 200.870 87.240 202.590 ;
        RECT 83.820 200.550 84.080 200.870 ;
        RECT 86.120 200.550 86.380 200.870 ;
        RECT 87.040 200.550 87.300 200.870 ;
        RECT 83.880 196.110 84.020 200.550 ;
        RECT 86.180 200.385 86.320 200.550 ;
        RECT 86.110 200.015 86.390 200.385 ;
        RECT 87.560 197.810 87.700 205.990 ;
        RECT 92.160 205.710 92.300 207.780 ;
        RECT 94.000 206.990 94.140 208.030 ;
        RECT 94.460 208.010 94.600 208.175 ;
        RECT 94.400 207.690 94.660 208.010 ;
        RECT 93.940 206.900 94.200 206.990 ;
        RECT 91.700 205.570 92.300 205.710 ;
        RECT 93.540 206.760 94.200 206.900 ;
        RECT 89.340 203.610 89.600 203.930 ;
        RECT 90.720 203.610 90.980 203.930 ;
        RECT 88.420 202.930 88.680 203.250 ;
        RECT 88.480 199.850 88.620 202.930 ;
        RECT 89.400 200.530 89.540 203.610 ;
        RECT 89.800 202.930 90.060 203.250 ;
        RECT 89.340 200.210 89.600 200.530 ;
        RECT 88.420 199.530 88.680 199.850 ;
        RECT 88.880 199.530 89.140 199.850 ;
        RECT 89.860 199.590 90.000 202.930 ;
        RECT 90.260 202.250 90.520 202.570 ;
        RECT 88.480 199.025 88.620 199.530 ;
        RECT 88.410 198.655 88.690 199.025 ;
        RECT 87.500 197.490 87.760 197.810 ;
        RECT 83.820 195.790 84.080 196.110 ;
        RECT 81.980 195.110 82.240 195.430 ;
        RECT 82.900 195.340 83.160 195.430 ;
        RECT 82.500 195.200 83.160 195.340 ;
        RECT 81.520 194.430 81.780 194.750 ;
        RECT 81.980 192.730 82.240 193.050 ;
        RECT 81.520 192.390 81.780 192.710 ;
        RECT 80.600 184.320 81.260 184.460 ;
        RECT 80.600 184.230 80.860 184.320 ;
        RECT 80.660 183.870 80.800 184.230 ;
        RECT 81.580 184.065 81.720 192.390 ;
        RECT 82.040 192.370 82.180 192.730 ;
        RECT 81.980 192.050 82.240 192.370 ;
        RECT 82.040 189.650 82.180 192.050 ;
        RECT 81.980 189.330 82.240 189.650 ;
        RECT 82.500 188.970 82.640 195.200 ;
        RECT 82.900 195.110 83.160 195.200 ;
        RECT 83.360 195.110 83.620 195.430 ;
        RECT 83.420 192.370 83.560 195.110 ;
        RECT 83.880 195.090 84.020 195.790 ;
        RECT 83.820 194.770 84.080 195.090 ;
        RECT 87.960 194.770 88.220 195.090 ;
        RECT 84.280 194.090 84.540 194.410 ;
        RECT 87.040 194.090 87.300 194.410 ;
        RECT 84.340 193.390 84.480 194.090 ;
        RECT 84.280 193.070 84.540 193.390 ;
        RECT 82.900 192.050 83.160 192.370 ;
        RECT 83.360 192.050 83.620 192.370 ;
        RECT 84.740 192.050 85.000 192.370 ;
        RECT 82.960 189.990 83.100 192.050 ;
        RECT 83.420 190.670 83.560 192.050 ;
        RECT 84.800 190.865 84.940 192.050 ;
        RECT 83.360 190.350 83.620 190.670 ;
        RECT 84.730 190.495 85.010 190.865 ;
        RECT 82.900 189.670 83.160 189.990 ;
        RECT 82.440 188.650 82.700 188.970 ;
        RECT 82.900 188.650 83.160 188.970 ;
        RECT 82.960 186.670 83.100 188.650 ;
        RECT 82.500 186.530 83.100 186.670 ;
        RECT 81.970 185.055 82.250 185.425 ;
        RECT 82.040 184.890 82.180 185.055 ;
        RECT 82.500 184.890 82.640 186.530 ;
        RECT 82.900 185.930 83.160 186.250 ;
        RECT 81.980 184.570 82.240 184.890 ;
        RECT 82.440 184.570 82.700 184.890 ;
        RECT 80.600 183.550 80.860 183.870 ;
        RECT 81.510 183.695 81.790 184.065 ;
        RECT 80.140 178.790 80.400 179.110 ;
        RECT 81.060 178.790 81.320 179.110 ;
        RECT 79.740 178.370 80.340 178.510 ;
        RECT 79.680 177.770 79.940 178.090 ;
        RECT 78.760 176.070 79.020 176.390 ;
        RECT 78.300 175.730 78.560 176.050 ;
        RECT 79.220 175.730 79.480 176.050 ;
        RECT 79.280 174.350 79.420 175.730 ;
        RECT 75.540 174.030 75.800 174.350 ;
        RECT 79.220 174.030 79.480 174.350 ;
        RECT 78.760 173.865 79.020 174.010 ;
        RECT 75.080 173.350 75.340 173.670 ;
        RECT 78.750 173.495 79.030 173.865 ;
        RECT 79.740 173.670 79.880 177.770 ;
        RECT 80.200 176.050 80.340 178.370 ;
        RECT 80.140 175.730 80.400 176.050 ;
        RECT 80.200 173.670 80.340 175.730 ;
        RECT 81.120 175.710 81.260 178.790 ;
        RECT 81.060 175.390 81.320 175.710 ;
        RECT 81.580 173.670 81.720 183.695 ;
        RECT 82.040 183.530 82.180 184.570 ;
        RECT 82.960 184.550 83.100 185.930 ;
        RECT 82.900 184.230 83.160 184.550 ;
        RECT 81.980 183.210 82.240 183.530 ;
        RECT 82.440 181.850 82.700 182.170 ;
        RECT 81.970 178.255 82.250 178.625 ;
        RECT 82.040 177.070 82.180 178.255 ;
        RECT 82.500 177.070 82.640 181.850 ;
        RECT 83.420 181.830 83.560 190.350 ;
        RECT 87.100 190.330 87.240 194.090 ;
        RECT 87.040 190.010 87.300 190.330 ;
        RECT 88.020 189.990 88.160 194.770 ;
        RECT 84.280 189.670 84.540 189.990 ;
        RECT 87.960 189.670 88.220 189.990 ;
        RECT 83.820 186.950 84.080 187.270 ;
        RECT 83.360 181.510 83.620 181.830 ;
        RECT 82.900 180.490 83.160 180.810 ;
        RECT 81.980 176.750 82.240 177.070 ;
        RECT 82.440 176.750 82.700 177.070 ;
        RECT 82.960 175.710 83.100 180.490 ;
        RECT 82.900 175.390 83.160 175.710 ;
        RECT 83.420 174.545 83.560 181.510 ;
        RECT 83.880 181.150 84.020 186.950 ;
        RECT 84.340 185.230 84.480 189.670 ;
        RECT 87.040 187.630 87.300 187.950 ;
        RECT 86.580 186.950 86.840 187.270 ;
        RECT 85.200 186.785 85.460 186.930 ;
        RECT 85.190 186.415 85.470 186.785 ;
        RECT 85.660 186.610 85.920 186.930 ;
        RECT 84.280 184.910 84.540 185.230 ;
        RECT 84.270 183.695 84.550 184.065 ;
        RECT 84.340 182.510 84.480 183.695 ;
        RECT 84.740 183.440 85.000 183.530 ;
        RECT 84.740 183.300 85.400 183.440 ;
        RECT 84.740 183.210 85.000 183.300 ;
        RECT 84.280 182.190 84.540 182.510 ;
        RECT 85.260 182.170 85.400 183.300 ;
        RECT 85.200 181.850 85.460 182.170 ;
        RECT 84.280 181.170 84.540 181.490 ;
        RECT 83.820 180.830 84.080 181.150 ;
        RECT 84.340 178.770 84.480 181.170 ;
        RECT 85.260 179.110 85.400 181.850 ;
        RECT 85.200 178.790 85.460 179.110 ;
        RECT 84.280 178.450 84.540 178.770 ;
        RECT 85.720 178.430 85.860 186.610 ;
        RECT 86.120 185.930 86.380 186.250 ;
        RECT 86.180 184.210 86.320 185.930 ;
        RECT 86.640 184.550 86.780 186.950 ;
        RECT 86.580 184.230 86.840 184.550 ;
        RECT 86.120 183.890 86.380 184.210 ;
        RECT 86.640 181.060 86.780 184.230 ;
        RECT 87.100 184.065 87.240 187.630 ;
        RECT 88.020 187.610 88.160 189.670 ;
        RECT 87.960 187.290 88.220 187.610 ;
        RECT 87.950 186.415 88.230 186.785 ;
        RECT 87.500 184.570 87.760 184.890 ;
        RECT 87.030 183.695 87.310 184.065 ;
        RECT 87.040 183.210 87.300 183.530 ;
        RECT 86.180 180.920 86.780 181.060 ;
        RECT 85.660 178.110 85.920 178.430 ;
        RECT 84.280 177.770 84.540 178.090 ;
        RECT 83.350 174.175 83.630 174.545 ;
        RECT 83.360 174.030 83.620 174.175 ;
        RECT 84.340 173.670 84.480 177.770 ;
        RECT 85.720 173.670 85.860 178.110 ;
        RECT 86.180 177.945 86.320 180.920 ;
        RECT 86.580 179.470 86.840 179.790 ;
        RECT 86.640 179.110 86.780 179.470 ;
        RECT 87.100 179.110 87.240 183.210 ;
        RECT 87.560 181.830 87.700 184.570 ;
        RECT 88.020 183.870 88.160 186.415 ;
        RECT 87.960 183.550 88.220 183.870 ;
        RECT 87.500 181.510 87.760 181.830 ;
        RECT 87.960 180.830 88.220 181.150 ;
        RECT 86.580 178.790 86.840 179.110 ;
        RECT 87.040 178.790 87.300 179.110 ;
        RECT 87.500 178.450 87.760 178.770 ;
        RECT 86.110 177.575 86.390 177.945 ;
        RECT 86.180 176.050 86.320 177.575 ;
        RECT 87.560 176.050 87.700 178.450 ;
        RECT 88.020 178.430 88.160 180.830 ;
        RECT 88.480 179.700 88.620 198.655 ;
        RECT 88.940 191.690 89.080 199.530 ;
        RECT 89.400 199.450 90.000 199.590 ;
        RECT 89.400 197.130 89.540 199.450 ;
        RECT 90.320 197.810 90.460 202.250 ;
        RECT 89.800 197.490 90.060 197.810 ;
        RECT 90.260 197.490 90.520 197.810 ;
        RECT 89.340 196.810 89.600 197.130 ;
        RECT 89.860 194.150 90.000 197.490 ;
        RECT 90.780 195.430 90.920 203.610 ;
        RECT 91.180 202.930 91.440 203.250 ;
        RECT 91.240 201.210 91.380 202.930 ;
        RECT 91.180 200.890 91.440 201.210 ;
        RECT 91.700 199.850 91.840 205.570 ;
        RECT 92.100 204.970 92.360 205.290 ;
        RECT 92.160 203.785 92.300 204.970 ;
        RECT 92.090 203.415 92.370 203.785 ;
        RECT 92.160 200.870 92.300 203.415 ;
        RECT 93.540 203.250 93.680 206.760 ;
        RECT 93.940 206.670 94.200 206.760 ;
        RECT 93.480 202.930 93.740 203.250 ;
        RECT 93.480 202.250 93.740 202.570 ;
        RECT 93.020 201.230 93.280 201.550 ;
        RECT 92.100 200.550 92.360 200.870 ;
        RECT 93.080 200.385 93.220 201.230 ;
        RECT 93.540 201.210 93.680 202.250 ;
        RECT 93.480 200.890 93.740 201.210 ;
        RECT 93.940 200.550 94.200 200.870 ;
        RECT 92.560 199.870 92.820 200.190 ;
        RECT 93.010 200.015 93.290 200.385 ;
        RECT 91.640 199.530 91.900 199.850 ;
        RECT 91.180 197.665 91.440 197.810 ;
        RECT 91.170 197.295 91.450 197.665 ;
        RECT 92.100 196.810 92.360 197.130 ;
        RECT 92.160 195.770 92.300 196.810 ;
        RECT 92.100 195.450 92.360 195.770 ;
        RECT 90.720 195.110 90.980 195.430 ;
        RECT 90.720 194.150 90.980 194.410 ;
        RECT 89.860 194.090 90.980 194.150 ;
        RECT 89.860 194.010 90.920 194.090 ;
        RECT 89.860 193.585 90.000 194.010 ;
        RECT 89.790 193.215 90.070 193.585 ;
        RECT 88.880 191.370 89.140 191.690 ;
        RECT 89.340 184.230 89.600 184.550 ;
        RECT 89.400 182.510 89.540 184.230 ;
        RECT 89.340 182.190 89.600 182.510 ;
        RECT 88.880 179.700 89.140 179.790 ;
        RECT 88.480 179.560 89.140 179.700 ;
        RECT 88.880 179.470 89.140 179.560 ;
        RECT 87.960 178.110 88.220 178.430 ;
        RECT 88.940 176.050 89.080 179.470 ;
        RECT 89.860 178.510 90.000 193.215 ;
        RECT 90.720 192.050 90.980 192.370 ;
        RECT 90.260 187.290 90.520 187.610 ;
        RECT 90.320 184.890 90.460 187.290 ;
        RECT 90.260 184.570 90.520 184.890 ;
        RECT 90.780 179.110 90.920 192.050 ;
        RECT 92.160 189.990 92.300 195.450 ;
        RECT 92.620 195.430 92.760 199.870 ;
        RECT 93.480 199.530 93.740 199.850 ;
        RECT 93.540 198.490 93.680 199.530 ;
        RECT 93.480 198.170 93.740 198.490 ;
        RECT 93.020 197.490 93.280 197.810 ;
        RECT 93.080 196.985 93.220 197.490 ;
        RECT 93.010 196.615 93.290 196.985 ;
        RECT 92.560 195.110 92.820 195.430 ;
        RECT 92.100 189.670 92.360 189.990 ;
        RECT 92.620 189.310 92.760 195.110 ;
        RECT 93.020 192.730 93.280 193.050 ;
        RECT 93.080 190.670 93.220 192.730 ;
        RECT 93.020 190.350 93.280 190.670 ;
        RECT 92.560 188.990 92.820 189.310 ;
        RECT 92.620 187.270 92.760 188.990 ;
        RECT 93.540 188.970 93.680 198.170 ;
        RECT 94.000 195.430 94.140 200.550 ;
        RECT 93.940 195.110 94.200 195.430 ;
        RECT 93.480 188.650 93.740 188.970 ;
        RECT 91.180 186.950 91.440 187.270 ;
        RECT 92.560 186.950 92.820 187.270 ;
        RECT 91.240 184.890 91.380 186.950 ;
        RECT 91.180 184.570 91.440 184.890 ;
        RECT 91.240 182.170 91.380 184.570 ;
        RECT 92.100 184.230 92.360 184.550 ;
        RECT 91.180 181.850 91.440 182.170 ;
        RECT 92.160 179.450 92.300 184.230 ;
        RECT 93.540 182.510 93.680 188.650 ;
        RECT 94.460 184.550 94.600 207.690 ;
        RECT 94.920 206.990 95.060 210.410 ;
        RECT 95.380 208.690 95.520 210.410 ;
        RECT 95.840 209.710 95.980 211.430 ;
        RECT 98.080 211.090 98.340 211.410 ;
        RECT 95.780 209.390 96.040 209.710 ;
        RECT 95.840 208.690 95.980 209.390 ;
        RECT 97.160 209.050 97.420 209.370 ;
        RECT 97.220 208.690 97.360 209.050 ;
        RECT 95.320 208.370 95.580 208.690 ;
        RECT 95.780 208.370 96.040 208.690 ;
        RECT 97.160 208.370 97.420 208.690 ;
        RECT 95.380 208.010 95.520 208.370 ;
        RECT 95.320 207.690 95.580 208.010 ;
        RECT 94.860 206.670 95.120 206.990 ;
        RECT 94.920 203.250 95.060 206.670 ;
        RECT 95.320 206.330 95.580 206.650 ;
        RECT 95.380 205.970 95.520 206.330 ;
        RECT 95.320 205.650 95.580 205.970 ;
        RECT 95.840 205.200 95.980 208.370 ;
        RECT 97.220 208.010 97.360 208.370 ;
        RECT 98.140 208.010 98.280 211.090 ;
        RECT 104.060 210.410 104.320 210.730 ;
        RECT 109.120 210.410 109.380 210.730 ;
        RECT 97.160 207.690 97.420 208.010 ;
        RECT 98.080 207.690 98.340 208.010 ;
        RECT 96.240 205.310 96.500 205.630 ;
        RECT 95.380 205.060 95.980 205.200 ;
        RECT 94.860 202.930 95.120 203.250 ;
        RECT 94.860 200.550 95.120 200.870 ;
        RECT 94.920 200.190 95.060 200.550 ;
        RECT 94.860 199.870 95.120 200.190 ;
        RECT 95.380 197.810 95.520 205.060 ;
        RECT 96.300 200.870 96.440 205.310 ;
        RECT 96.240 200.550 96.500 200.870 ;
        RECT 96.700 200.550 96.960 200.870 ;
        RECT 96.300 199.025 96.440 200.550 ;
        RECT 96.230 198.655 96.510 199.025 ;
        RECT 96.230 197.975 96.510 198.345 ;
        RECT 94.860 197.490 95.120 197.810 ;
        RECT 95.320 197.665 95.580 197.810 ;
        RECT 94.920 197.130 95.060 197.490 ;
        RECT 95.310 197.295 95.590 197.665 ;
        RECT 95.780 197.490 96.040 197.810 ;
        RECT 94.860 196.810 95.120 197.130 ;
        RECT 95.380 188.970 95.520 197.295 ;
        RECT 95.840 195.625 95.980 197.490 ;
        RECT 95.770 195.255 96.050 195.625 ;
        RECT 95.840 191.690 95.980 195.255 ;
        RECT 95.780 191.370 96.040 191.690 ;
        RECT 95.320 188.650 95.580 188.970 ;
        RECT 94.860 184.570 95.120 184.890 ;
        RECT 94.400 184.230 94.660 184.550 ;
        RECT 93.480 182.190 93.740 182.510 ;
        RECT 93.480 180.490 93.740 180.810 ;
        RECT 92.100 179.130 92.360 179.450 ;
        RECT 90.720 178.790 90.980 179.110 ;
        RECT 93.540 178.770 93.680 180.490 ;
        RECT 89.860 178.370 90.920 178.510 ;
        RECT 93.480 178.450 93.740 178.770 ;
        RECT 89.800 177.770 90.060 178.090 ;
        RECT 86.120 175.730 86.380 176.050 ;
        RECT 87.500 175.730 87.760 176.050 ;
        RECT 88.880 175.730 89.140 176.050 ;
        RECT 89.860 175.370 90.000 177.770 ;
        RECT 90.780 176.050 90.920 178.370 ;
        RECT 90.720 175.730 90.980 176.050 ;
        RECT 89.800 175.050 90.060 175.370 ;
        RECT 79.680 173.350 79.940 173.670 ;
        RECT 80.140 173.350 80.400 173.670 ;
        RECT 81.520 173.350 81.780 173.670 ;
        RECT 84.280 173.350 84.540 173.670 ;
        RECT 85.660 173.350 85.920 173.670 ;
        RECT 70.020 173.010 70.280 173.330 ;
        RECT 74.160 173.010 74.420 173.330 ;
        RECT 69.100 172.330 69.360 172.650 ;
        RECT 70.080 171.630 70.220 173.010 ;
        RECT 71.860 172.330 72.120 172.650 ;
        RECT 68.640 171.310 68.900 171.630 ;
        RECT 70.020 171.310 70.280 171.630 ;
        RECT 66.800 170.630 67.060 170.950 ;
        RECT 68.700 170.610 68.840 171.310 ;
        RECT 71.920 171.290 72.060 172.330 ;
        RECT 74.220 171.630 74.360 173.010 ;
        RECT 82.440 172.330 82.700 172.650 ;
        RECT 74.160 171.310 74.420 171.630 ;
        RECT 71.860 170.970 72.120 171.290 ;
        RECT 82.500 170.610 82.640 172.330 ;
        RECT 85.720 171.630 85.860 173.350 ;
        RECT 93.540 173.330 93.680 178.450 ;
        RECT 93.940 175.390 94.200 175.710 ;
        RECT 94.000 174.350 94.140 175.390 ;
        RECT 94.920 174.350 95.060 184.570 ;
        RECT 96.300 183.530 96.440 197.975 ;
        RECT 96.760 197.130 96.900 200.550 ;
        RECT 97.220 198.345 97.360 207.690 ;
        RECT 104.120 202.910 104.260 210.410 ;
        RECT 106.570 207.155 108.110 207.525 ;
        RECT 109.180 206.505 109.320 210.410 ;
        RECT 109.870 209.875 111.410 210.245 ;
        RECT 128.430 209.535 128.710 209.905 ;
        RECT 128.440 209.390 128.700 209.535 ;
        RECT 109.110 206.135 109.390 206.505 ;
        RECT 105.900 202.930 106.160 203.250 ;
        RECT 104.060 202.590 104.320 202.910 ;
        RECT 99.920 202.250 100.180 202.570 ;
        RECT 99.000 199.530 99.260 199.850 ;
        RECT 97.150 197.975 97.430 198.345 ;
        RECT 97.160 197.665 97.420 197.810 ;
        RECT 97.150 197.295 97.430 197.665 ;
        RECT 98.080 197.380 98.340 197.470 ;
        RECT 98.080 197.240 98.740 197.380 ;
        RECT 98.080 197.150 98.340 197.240 ;
        RECT 96.700 196.810 96.960 197.130 ;
        RECT 97.160 196.810 97.420 197.130 ;
        RECT 97.220 196.305 97.360 196.810 ;
        RECT 97.150 195.935 97.430 196.305 ;
        RECT 98.600 196.110 98.740 197.240 ;
        RECT 96.240 183.210 96.500 183.530 ;
        RECT 97.220 181.150 97.360 195.935 ;
        RECT 98.540 195.790 98.800 196.110 ;
        RECT 98.540 187.290 98.800 187.610 ;
        RECT 98.600 186.930 98.740 187.290 ;
        RECT 99.060 186.930 99.200 199.530 ;
        RECT 99.980 198.830 100.120 202.250 ;
        RECT 101.300 200.550 101.560 200.870 ;
        RECT 102.220 200.550 102.480 200.870 ;
        RECT 100.380 200.210 100.640 200.530 ;
        RECT 100.440 198.830 100.580 200.210 ;
        RECT 99.920 198.510 100.180 198.830 ;
        RECT 100.380 198.510 100.640 198.830 ;
        RECT 99.460 198.170 99.720 198.490 ;
        RECT 99.520 197.130 99.660 198.170 ;
        RECT 101.360 198.150 101.500 200.550 ;
        RECT 102.280 198.830 102.420 200.550 ;
        RECT 102.680 199.870 102.940 200.190 ;
        RECT 102.740 198.830 102.880 199.870 ;
        RECT 104.120 199.705 104.260 202.590 ;
        RECT 105.960 200.190 106.100 202.930 ;
        RECT 109.180 202.910 109.320 206.135 ;
        RECT 109.870 204.435 111.410 204.805 ;
        RECT 111.880 202.930 112.140 203.250 ;
        RECT 108.660 202.590 108.920 202.910 ;
        RECT 109.120 202.590 109.380 202.910 ;
        RECT 108.200 202.250 108.460 202.570 ;
        RECT 106.570 201.715 108.110 202.085 ;
        RECT 106.350 200.695 106.630 201.065 ;
        RECT 106.420 200.530 106.560 200.695 ;
        RECT 106.360 200.210 106.620 200.530 ;
        RECT 105.900 199.870 106.160 200.190 ;
        RECT 104.050 199.335 104.330 199.705 ;
        RECT 104.980 199.530 105.240 199.850 ;
        RECT 102.220 198.510 102.480 198.830 ;
        RECT 102.680 198.510 102.940 198.830 ;
        RECT 105.040 198.230 105.180 199.530 ;
        RECT 101.300 197.830 101.560 198.150 ;
        RECT 104.120 198.090 105.180 198.230 ;
        RECT 104.120 197.810 104.260 198.090 ;
        RECT 99.920 197.490 100.180 197.810 ;
        RECT 99.460 196.810 99.720 197.130 ;
        RECT 99.980 196.985 100.120 197.490 ;
        RECT 102.670 197.295 102.950 197.665 ;
        RECT 103.600 197.490 103.860 197.810 ;
        RECT 104.060 197.490 104.320 197.810 ;
        RECT 104.520 197.490 104.780 197.810 ;
        RECT 99.910 196.615 100.190 196.985 ;
        RECT 101.300 196.810 101.560 197.130 ;
        RECT 99.920 191.710 100.180 192.030 ;
        RECT 99.460 189.670 99.720 189.990 ;
        RECT 98.540 186.610 98.800 186.930 ;
        RECT 99.000 186.610 99.260 186.930 ;
        RECT 98.540 185.930 98.800 186.250 ;
        RECT 98.600 184.550 98.740 185.930 ;
        RECT 99.000 184.570 99.260 184.890 ;
        RECT 98.080 184.230 98.340 184.550 ;
        RECT 98.540 184.230 98.800 184.550 ;
        RECT 98.140 183.530 98.280 184.230 ;
        RECT 98.080 183.210 98.340 183.530 ;
        RECT 99.060 181.490 99.200 184.570 ;
        RECT 99.000 181.170 99.260 181.490 ;
        RECT 97.160 180.830 97.420 181.150 ;
        RECT 95.780 178.450 96.040 178.770 ;
        RECT 95.840 177.070 95.980 178.450 ;
        RECT 97.620 177.770 97.880 178.090 ;
        RECT 98.080 177.770 98.340 178.090 ;
        RECT 95.780 176.750 96.040 177.070 ;
        RECT 97.160 175.960 97.420 176.050 ;
        RECT 96.760 175.820 97.420 175.960 ;
        RECT 93.940 174.030 94.200 174.350 ;
        RECT 94.860 174.030 95.120 174.350 ;
        RECT 96.760 173.670 96.900 175.820 ;
        RECT 97.160 175.730 97.420 175.820 ;
        RECT 97.160 175.050 97.420 175.370 ;
        RECT 96.700 173.350 96.960 173.670 ;
        RECT 97.220 173.330 97.360 175.050 ;
        RECT 97.680 174.010 97.820 177.770 ;
        RECT 98.140 176.730 98.280 177.770 ;
        RECT 98.080 176.410 98.340 176.730 ;
        RECT 98.080 175.730 98.340 176.050 ;
        RECT 98.540 175.730 98.800 176.050 ;
        RECT 98.140 175.370 98.280 175.730 ;
        RECT 98.080 175.050 98.340 175.370 ;
        RECT 97.620 173.690 97.880 174.010 ;
        RECT 98.140 173.670 98.280 175.050 ;
        RECT 98.600 174.350 98.740 175.730 ;
        RECT 98.540 174.030 98.800 174.350 ;
        RECT 98.080 173.350 98.340 173.670 ;
        RECT 93.480 173.010 93.740 173.330 ;
        RECT 97.160 173.010 97.420 173.330 ;
        RECT 99.520 172.650 99.660 189.670 ;
        RECT 99.980 189.310 100.120 191.710 ;
        RECT 100.380 190.010 100.640 190.330 ;
        RECT 99.920 188.990 100.180 189.310 ;
        RECT 99.920 186.840 100.180 186.930 ;
        RECT 100.440 186.840 100.580 190.010 ;
        RECT 101.360 189.990 101.500 196.810 ;
        RECT 102.220 190.350 102.480 190.670 ;
        RECT 101.300 189.670 101.560 189.990 ;
        RECT 101.760 188.990 102.020 189.310 ;
        RECT 101.820 187.950 101.960 188.990 ;
        RECT 101.760 187.630 102.020 187.950 ;
        RECT 101.820 187.270 101.960 187.630 ;
        RECT 101.760 186.950 102.020 187.270 ;
        RECT 99.920 186.700 100.580 186.840 ;
        RECT 99.920 186.610 100.180 186.700 ;
        RECT 100.840 186.270 101.100 186.590 ;
        RECT 99.920 183.550 100.180 183.870 ;
        RECT 99.980 181.490 100.120 183.550 ;
        RECT 99.920 181.170 100.180 181.490 ;
        RECT 100.380 178.790 100.640 179.110 ;
        RECT 100.440 177.070 100.580 178.790 ;
        RECT 100.900 178.430 101.040 186.270 ;
        RECT 101.300 185.930 101.560 186.250 ;
        RECT 101.360 184.890 101.500 185.930 ;
        RECT 101.300 184.570 101.560 184.890 ;
        RECT 101.760 184.230 102.020 184.550 ;
        RECT 101.820 182.170 101.960 184.230 ;
        RECT 101.760 181.850 102.020 182.170 ;
        RECT 101.300 179.130 101.560 179.450 ;
        RECT 102.280 179.305 102.420 190.350 ;
        RECT 102.740 182.170 102.880 197.295 ;
        RECT 103.140 195.110 103.400 195.430 ;
        RECT 103.200 190.670 103.340 195.110 ;
        RECT 103.660 195.000 103.800 197.490 ;
        RECT 104.580 195.430 104.720 197.490 ;
        RECT 104.520 195.110 104.780 195.430 ;
        RECT 104.060 195.000 104.320 195.090 ;
        RECT 103.660 194.860 104.320 195.000 ;
        RECT 104.060 194.770 104.320 194.860 ;
        RECT 104.120 194.410 104.260 194.770 ;
        RECT 104.060 194.265 104.320 194.410 ;
        RECT 104.050 193.895 104.330 194.265 ;
        RECT 103.600 192.390 103.860 192.710 ;
        RECT 103.140 190.350 103.400 190.670 ;
        RECT 103.200 187.610 103.340 190.350 ;
        RECT 103.660 189.990 103.800 192.390 ;
        RECT 104.120 192.370 104.260 193.895 ;
        RECT 104.580 193.390 104.720 195.110 ;
        RECT 105.040 194.750 105.180 198.090 ;
        RECT 105.440 197.490 105.700 197.810 ;
        RECT 106.420 197.550 106.560 200.210 ;
        RECT 107.740 199.870 108.000 200.190 ;
        RECT 105.500 196.305 105.640 197.490 ;
        RECT 105.960 197.410 106.560 197.550 ;
        RECT 105.430 195.935 105.710 196.305 ;
        RECT 105.960 195.430 106.100 197.410 ;
        RECT 107.800 197.040 107.940 199.870 ;
        RECT 108.260 198.490 108.400 202.250 ;
        RECT 108.720 201.210 108.860 202.590 ;
        RECT 111.940 201.210 112.080 202.930 ;
        RECT 108.660 200.890 108.920 201.210 ;
        RECT 111.880 200.890 112.140 201.210 ;
        RECT 108.720 200.190 108.860 200.890 ;
        RECT 108.660 199.870 108.920 200.190 ;
        RECT 108.200 198.170 108.460 198.490 ;
        RECT 107.800 196.900 108.400 197.040 ;
        RECT 106.570 196.275 108.110 196.645 ;
        RECT 105.900 195.110 106.160 195.430 ;
        RECT 107.280 195.110 107.540 195.430 ;
        RECT 108.260 195.340 108.400 196.900 ;
        RECT 107.800 195.200 108.400 195.340 ;
        RECT 104.980 194.430 105.240 194.750 ;
        RECT 104.520 193.070 104.780 193.390 ;
        RECT 107.340 193.050 107.480 195.110 ;
        RECT 107.800 193.050 107.940 195.200 ;
        RECT 108.200 194.430 108.460 194.750 ;
        RECT 104.980 192.730 105.240 193.050 ;
        RECT 107.280 192.730 107.540 193.050 ;
        RECT 107.740 192.730 108.000 193.050 ;
        RECT 104.060 192.050 104.320 192.370 ;
        RECT 103.600 189.670 103.860 189.990 ;
        RECT 103.600 188.650 103.860 188.970 ;
        RECT 103.140 187.290 103.400 187.610 ;
        RECT 103.140 183.210 103.400 183.530 ;
        RECT 103.660 183.270 103.800 188.650 ;
        RECT 104.120 183.870 104.260 192.050 ;
        RECT 105.040 190.580 105.180 192.730 ;
        RECT 107.800 192.370 107.940 192.730 ;
        RECT 107.740 192.050 108.000 192.370 ;
        RECT 106.570 190.835 108.110 191.205 ;
        RECT 104.580 190.440 105.180 190.580 ;
        RECT 104.580 187.350 104.720 190.440 ;
        RECT 106.360 190.010 106.620 190.330 ;
        RECT 105.900 189.670 106.160 189.990 ;
        RECT 105.960 189.310 106.100 189.670 ;
        RECT 105.900 188.990 106.160 189.310 ;
        RECT 105.960 187.610 106.100 188.990 ;
        RECT 104.580 187.210 105.180 187.350 ;
        RECT 105.440 187.290 105.700 187.610 ;
        RECT 105.900 187.290 106.160 187.610 ;
        RECT 104.060 183.550 104.320 183.870 ;
        RECT 102.680 181.850 102.940 182.170 ;
        RECT 100.840 178.110 101.100 178.430 ;
        RECT 100.380 176.750 100.640 177.070 ;
        RECT 101.360 174.010 101.500 179.130 ;
        RECT 101.760 178.790 102.020 179.110 ;
        RECT 102.210 178.935 102.490 179.305 ;
        RECT 101.820 177.070 101.960 178.790 ;
        RECT 101.760 176.750 102.020 177.070 ;
        RECT 102.280 175.370 102.420 178.935 ;
        RECT 102.680 178.790 102.940 179.110 ;
        RECT 102.740 178.090 102.880 178.790 ;
        RECT 102.680 177.770 102.940 178.090 ;
        RECT 103.200 176.730 103.340 183.210 ;
        RECT 103.660 183.130 104.720 183.270 ;
        RECT 104.060 182.190 104.320 182.510 ;
        RECT 104.120 181.910 104.260 182.190 ;
        RECT 103.660 181.770 104.260 181.910 ;
        RECT 103.660 179.110 103.800 181.770 ;
        RECT 104.060 181.170 104.320 181.490 ;
        RECT 104.120 179.790 104.260 181.170 ;
        RECT 104.060 179.470 104.320 179.790 ;
        RECT 103.600 178.790 103.860 179.110 ;
        RECT 103.140 176.410 103.400 176.730 ;
        RECT 103.200 176.050 103.340 176.410 ;
        RECT 104.120 176.390 104.260 179.470 ;
        RECT 104.580 179.110 104.720 183.130 ;
        RECT 105.040 182.510 105.180 187.210 ;
        RECT 105.500 184.210 105.640 187.290 ;
        RECT 105.900 186.500 106.160 186.590 ;
        RECT 106.420 186.500 106.560 190.010 ;
        RECT 108.260 187.950 108.400 194.430 ;
        RECT 108.720 193.390 108.860 199.870 ;
        RECT 109.870 198.995 111.410 199.365 ;
        RECT 129.350 199.335 129.630 199.705 ;
        RECT 129.420 197.810 129.560 199.335 ;
        RECT 109.120 197.490 109.380 197.810 ;
        RECT 110.040 197.490 110.300 197.810 ;
        RECT 111.420 197.490 111.680 197.810 ;
        RECT 109.180 196.110 109.320 197.490 ;
        RECT 110.100 196.110 110.240 197.490 ;
        RECT 109.120 195.790 109.380 196.110 ;
        RECT 110.040 195.790 110.300 196.110 ;
        RECT 111.480 195.770 111.620 197.490 ;
        RECT 112.330 197.295 112.610 197.665 ;
        RECT 112.800 197.490 113.060 197.810 ;
        RECT 129.360 197.490 129.620 197.810 ;
        RECT 112.400 197.130 112.540 197.295 ;
        RECT 112.340 196.810 112.600 197.130 ;
        RECT 111.420 195.450 111.680 195.770 ;
        RECT 109.120 195.110 109.380 195.430 ;
        RECT 108.660 193.070 108.920 193.390 ;
        RECT 109.180 193.050 109.320 195.110 ;
        RECT 111.480 194.830 111.620 195.450 ;
        RECT 112.400 195.430 112.540 196.810 ;
        RECT 112.340 195.110 112.600 195.430 ;
        RECT 111.480 194.690 112.080 194.830 ;
        RECT 109.870 193.555 111.410 193.925 ;
        RECT 109.580 193.070 109.840 193.390 ;
        RECT 109.120 192.730 109.380 193.050 ;
        RECT 108.660 191.370 108.920 191.690 ;
        RECT 108.720 189.990 108.860 191.370 ;
        RECT 109.180 190.330 109.320 192.730 ;
        RECT 109.640 190.330 109.780 193.070 ;
        RECT 111.940 192.710 112.080 194.690 ;
        RECT 112.340 194.430 112.600 194.750 ;
        RECT 111.880 192.390 112.140 192.710 ;
        RECT 112.400 192.370 112.540 194.430 ;
        RECT 110.500 192.050 110.760 192.370 ;
        RECT 110.960 192.050 111.220 192.370 ;
        RECT 112.340 192.050 112.600 192.370 ;
        RECT 110.560 190.670 110.700 192.050 ;
        RECT 110.500 190.350 110.760 190.670 ;
        RECT 109.120 190.010 109.380 190.330 ;
        RECT 109.580 190.010 109.840 190.330 ;
        RECT 108.660 189.670 108.920 189.990 ;
        RECT 108.200 187.630 108.460 187.950 ;
        RECT 105.900 186.360 106.560 186.500 ;
        RECT 105.900 186.270 106.160 186.360 ;
        RECT 108.200 185.930 108.460 186.250 ;
        RECT 106.570 185.395 108.110 185.765 ;
        RECT 105.890 184.375 106.170 184.745 ;
        RECT 105.440 183.890 105.700 184.210 ;
        RECT 105.440 183.210 105.700 183.530 ;
        RECT 104.980 182.190 105.240 182.510 ;
        RECT 105.500 181.830 105.640 183.210 ;
        RECT 105.440 181.510 105.700 181.830 ;
        RECT 104.980 180.830 105.240 181.150 ;
        RECT 104.520 178.790 104.780 179.110 ;
        RECT 104.060 176.070 104.320 176.390 ;
        RECT 103.140 175.730 103.400 176.050 ;
        RECT 102.220 175.050 102.480 175.370 ;
        RECT 103.600 175.050 103.860 175.370 ;
        RECT 103.660 174.350 103.800 175.050 ;
        RECT 103.600 174.030 103.860 174.350 ;
        RECT 101.300 173.690 101.560 174.010 ;
        RECT 105.040 173.670 105.180 180.830 ;
        RECT 105.500 180.810 105.640 181.510 ;
        RECT 105.440 180.490 105.700 180.810 ;
        RECT 105.500 178.430 105.640 180.490 ;
        RECT 105.440 178.110 105.700 178.430 ;
        RECT 105.500 176.050 105.640 178.110 ;
        RECT 105.440 175.730 105.700 176.050 ;
        RECT 103.140 173.350 103.400 173.670 ;
        RECT 104.980 173.350 105.240 173.670 ;
        RECT 99.460 172.330 99.720 172.650 ;
        RECT 103.200 171.630 103.340 173.350 ;
        RECT 85.660 171.310 85.920 171.630 ;
        RECT 103.140 171.310 103.400 171.630 ;
        RECT 105.040 171.290 105.180 173.350 ;
        RECT 105.500 173.330 105.640 175.730 ;
        RECT 105.960 173.920 106.100 184.375 ;
        RECT 107.740 182.190 108.000 182.510 ;
        RECT 107.800 181.490 107.940 182.190 ;
        RECT 108.260 181.490 108.400 185.930 ;
        RECT 108.720 184.890 108.860 189.670 ;
        RECT 109.640 189.220 109.780 190.010 ;
        RECT 109.180 189.080 109.780 189.220 ;
        RECT 109.180 186.590 109.320 189.080 ;
        RECT 111.020 188.970 111.160 192.050 ;
        RECT 111.880 191.430 112.140 191.690 ;
        RECT 111.480 191.370 112.140 191.430 ;
        RECT 111.480 191.290 112.080 191.370 ;
        RECT 111.480 189.650 111.620 191.290 ;
        RECT 112.340 190.350 112.600 190.670 ;
        RECT 111.420 189.330 111.680 189.650 ;
        RECT 110.960 188.650 111.220 188.970 ;
        RECT 111.480 188.880 111.620 189.330 ;
        RECT 111.480 188.740 112.080 188.880 ;
        RECT 109.870 188.115 111.410 188.485 ;
        RECT 110.040 187.630 110.300 187.950 ;
        RECT 110.500 187.630 110.760 187.950 ;
        RECT 109.120 186.270 109.380 186.590 ;
        RECT 108.660 184.570 108.920 184.890 ;
        RECT 109.110 184.375 109.390 184.745 ;
        RECT 109.120 184.230 109.380 184.375 ;
        RECT 110.100 184.210 110.240 187.630 ;
        RECT 110.560 186.930 110.700 187.630 ;
        RECT 110.500 186.610 110.760 186.930 ;
        RECT 111.940 186.670 112.080 188.740 ;
        RECT 112.400 187.950 112.540 190.350 ;
        RECT 112.340 187.630 112.600 187.950 ;
        RECT 112.860 187.270 113.000 197.490 ;
        RECT 128.430 195.935 128.710 196.305 ;
        RECT 128.440 195.790 128.700 195.935 ;
        RECT 114.640 192.730 114.900 193.050 ;
        RECT 113.250 191.855 113.530 192.225 ;
        RECT 112.800 186.950 113.060 187.270 ;
        RECT 111.480 186.590 112.080 186.670 ;
        RECT 111.480 186.530 112.140 186.590 ;
        RECT 111.480 184.550 111.620 186.530 ;
        RECT 111.880 186.270 112.140 186.530 ;
        RECT 112.860 185.230 113.000 186.950 ;
        RECT 112.800 184.910 113.060 185.230 ;
        RECT 111.420 184.230 111.680 184.550 ;
        RECT 110.040 183.890 110.300 184.210 ;
        RECT 109.120 183.210 109.380 183.530 ;
        RECT 107.280 181.170 107.540 181.490 ;
        RECT 107.740 181.170 108.000 181.490 ;
        RECT 108.200 181.170 108.460 181.490 ;
        RECT 107.340 180.720 107.480 181.170 ;
        RECT 107.340 180.580 108.400 180.720 ;
        RECT 106.570 179.955 108.110 180.325 ;
        RECT 108.260 179.790 108.400 180.580 ;
        RECT 108.200 179.470 108.460 179.790 ;
        RECT 107.280 178.790 107.540 179.110 ;
        RECT 106.820 178.450 107.080 178.770 ;
        RECT 106.880 175.710 107.020 178.450 ;
        RECT 107.340 177.070 107.480 178.790 ;
        RECT 107.280 176.750 107.540 177.070 ;
        RECT 108.660 176.410 108.920 176.730 ;
        RECT 106.820 175.430 107.080 175.710 ;
        RECT 106.820 175.390 107.940 175.430 ;
        RECT 106.880 175.290 107.940 175.390 ;
        RECT 107.800 175.280 107.940 175.290 ;
        RECT 107.800 175.140 108.400 175.280 ;
        RECT 106.570 174.515 108.110 174.885 ;
        RECT 106.360 173.920 106.620 174.010 ;
        RECT 105.960 173.780 106.620 173.920 ;
        RECT 106.360 173.690 106.620 173.780 ;
        RECT 105.440 173.010 105.700 173.330 ;
        RECT 104.980 170.970 105.240 171.290 ;
        RECT 108.260 170.950 108.400 175.140 ;
        RECT 108.200 170.630 108.460 170.950 ;
        RECT 108.720 170.610 108.860 176.410 ;
        RECT 109.180 176.050 109.320 183.210 ;
        RECT 109.870 182.675 111.410 183.045 ;
        RECT 112.860 181.490 113.000 184.910 ;
        RECT 113.320 184.550 113.460 191.855 ;
        RECT 114.700 190.670 114.840 192.730 ;
        RECT 128.430 192.535 128.710 192.905 ;
        RECT 128.500 192.370 128.640 192.535 ;
        RECT 115.560 192.050 115.820 192.370 ;
        RECT 114.640 190.350 114.900 190.670 ;
        RECT 115.620 189.990 115.760 192.050 ;
        RECT 116.930 191.855 117.210 192.225 ;
        RECT 121.540 192.050 121.800 192.370 ;
        RECT 128.440 192.050 128.700 192.370 ;
        RECT 117.000 190.670 117.140 191.855 ;
        RECT 121.600 190.670 121.740 192.050 ;
        RECT 123.840 191.370 124.100 191.690 ;
        RECT 124.300 191.370 124.560 191.690 ;
        RECT 116.940 190.350 117.200 190.670 ;
        RECT 121.540 190.350 121.800 190.670 ;
        RECT 115.560 189.670 115.820 189.990 ;
        RECT 115.620 189.310 115.760 189.670 ;
        RECT 122.460 189.330 122.720 189.650 ;
        RECT 115.560 188.990 115.820 189.310 ;
        RECT 113.260 184.230 113.520 184.550 ;
        RECT 115.620 183.870 115.760 188.990 ;
        RECT 122.520 188.970 122.660 189.330 ;
        RECT 122.460 188.650 122.720 188.970 ;
        RECT 122.520 184.550 122.660 188.650 ;
        RECT 123.900 186.930 124.040 191.370 ;
        RECT 124.360 189.990 124.500 191.370 ;
        RECT 124.300 189.670 124.560 189.990 ;
        RECT 131.190 189.135 131.470 189.505 ;
        RECT 131.260 187.950 131.400 189.135 ;
        RECT 131.200 187.630 131.460 187.950 ;
        RECT 123.840 186.610 124.100 186.930 ;
        RECT 130.270 185.735 130.550 186.105 ;
        RECT 130.340 184.550 130.480 185.735 ;
        RECT 122.460 184.230 122.720 184.550 ;
        RECT 130.280 184.230 130.540 184.550 ;
        RECT 115.560 183.550 115.820 183.870 ;
        RECT 113.260 183.210 113.520 183.530 ;
        RECT 112.800 181.170 113.060 181.490 ;
        RECT 111.880 180.830 112.140 181.150 ;
        RECT 111.420 180.490 111.680 180.810 ;
        RECT 111.480 179.790 111.620 180.490 ;
        RECT 111.420 179.470 111.680 179.790 ;
        RECT 109.870 177.235 111.410 177.605 ;
        RECT 111.940 177.070 112.080 180.830 ;
        RECT 113.320 180.810 113.460 183.210 ;
        RECT 113.260 180.490 113.520 180.810 ;
        RECT 116.020 180.490 116.280 180.810 ;
        RECT 113.320 179.450 113.460 180.490 ;
        RECT 113.260 179.130 113.520 179.450 ;
        RECT 115.550 178.935 115.830 179.305 ;
        RECT 116.080 179.110 116.220 180.490 ;
        RECT 115.560 178.790 115.820 178.935 ;
        RECT 116.020 178.790 116.280 179.110 ;
        RECT 111.880 176.750 112.140 177.070 ;
        RECT 109.120 175.730 109.380 176.050 ;
        RECT 109.180 174.010 109.320 175.730 ;
        RECT 109.580 175.050 109.840 175.370 ;
        RECT 109.640 174.350 109.780 175.050 ;
        RECT 109.580 174.030 109.840 174.350 ;
        RECT 109.120 173.690 109.380 174.010 ;
        RECT 115.620 173.670 115.760 178.790 ;
        RECT 130.270 175.535 130.550 175.905 ;
        RECT 123.840 175.050 124.100 175.370 ;
        RECT 123.900 173.670 124.040 175.050 ;
        RECT 130.340 174.350 130.480 175.535 ;
        RECT 130.280 174.030 130.540 174.350 ;
        RECT 115.560 173.350 115.820 173.670 ;
        RECT 123.840 173.350 124.100 173.670 ;
        RECT 111.880 172.330 112.140 172.650 ;
        RECT 109.870 171.795 111.410 172.165 ;
        RECT 111.940 171.630 112.080 172.330 ;
        RECT 111.880 171.310 112.140 171.630 ;
        RECT 115.620 170.610 115.760 173.350 ;
        RECT 122.460 172.330 122.720 172.650 ;
        RECT 122.520 170.610 122.660 172.330 ;
        RECT 130.270 172.135 130.550 172.505 ;
        RECT 130.340 171.630 130.480 172.135 ;
        RECT 130.280 171.310 130.540 171.630 ;
        RECT 125.680 170.630 125.940 170.950 ;
        RECT 57.140 170.290 57.400 170.610 ;
        RECT 58.980 170.290 59.240 170.610 ;
        RECT 62.660 170.290 62.920 170.610 ;
        RECT 67.720 170.290 67.980 170.610 ;
        RECT 68.640 170.290 68.900 170.610 ;
        RECT 70.940 170.290 71.200 170.610 ;
        RECT 77.380 170.290 77.640 170.610 ;
        RECT 82.440 170.290 82.700 170.610 ;
        RECT 87.040 170.290 87.300 170.610 ;
        RECT 108.660 170.290 108.920 170.610 ;
        RECT 115.560 170.290 115.820 170.610 ;
        RECT 122.460 170.290 122.720 170.610 ;
        RECT 56.220 169.950 56.480 170.270 ;
        RECT 54.840 169.610 55.100 169.930 ;
        RECT 51.680 167.490 52.280 167.630 ;
        RECT 31.900 157.290 32.570 157.310 ;
        RECT 31.900 157.130 32.040 157.290 ;
        RECT 30.980 156.990 32.040 157.130 ;
        RECT 32.290 156.810 32.570 157.290 ;
        RECT 35.510 156.810 35.790 157.310 ;
        RECT 38.730 156.810 39.010 157.310 ;
        RECT 41.950 156.810 42.230 157.310 ;
        RECT 45.170 156.810 45.450 157.310 ;
        RECT 48.390 156.810 48.670 157.310 ;
        RECT 51.160 157.030 51.420 157.350 ;
        RECT 51.680 157.310 51.820 167.490 ;
        RECT 54.900 157.310 55.040 169.610 ;
        RECT 57.200 168.910 57.340 170.290 ;
        RECT 58.060 169.610 58.320 169.930 ;
        RECT 64.500 169.610 64.760 169.930 ;
        RECT 57.140 168.590 57.400 168.910 ;
        RECT 58.120 157.310 58.260 169.610 ;
        RECT 61.280 168.590 61.540 168.910 ;
        RECT 61.340 157.310 61.480 168.590 ;
        RECT 64.560 157.310 64.700 169.610 ;
        RECT 67.780 157.310 67.920 170.290 ;
        RECT 71.000 157.310 71.140 170.290 ;
        RECT 74.160 169.610 74.420 169.930 ;
        RECT 74.220 157.310 74.360 169.610 ;
        RECT 77.440 157.310 77.580 170.290 ;
        RECT 83.820 169.610 84.080 169.930 ;
        RECT 83.880 157.310 84.020 169.610 ;
        RECT 87.100 157.310 87.240 170.290 ;
        RECT 106.570 169.075 108.110 169.445 ;
        RECT 125.740 169.105 125.880 170.630 ;
        RECT 125.670 168.735 125.950 169.105 ;
        RECT 51.610 156.810 51.890 157.310 ;
        RECT 54.830 156.810 55.110 157.310 ;
        RECT 58.050 156.810 58.330 157.310 ;
        RECT 61.270 156.810 61.550 157.310 ;
        RECT 64.490 156.810 64.770 157.310 ;
        RECT 67.710 156.810 67.990 157.310 ;
        RECT 70.930 156.810 71.210 157.310 ;
        RECT 74.150 156.810 74.430 157.310 ;
        RECT 77.370 156.810 77.650 157.310 ;
        RECT 83.810 156.810 84.090 157.310 ;
        RECT 87.030 156.810 87.310 157.310 ;
        RECT 129.445 65.905 134.480 65.940 ;
        RECT 129.445 65.265 134.570 65.905 ;
        RECT 134.430 65.260 134.570 65.265 ;
        RECT 133.790 64.720 133.930 64.725 ;
        RECT 128.795 64.625 133.930 64.720 ;
        RECT 128.745 64.105 133.930 64.625 ;
        RECT 128.745 64.070 128.905 64.105 ;
        RECT 127.185 62.660 128.670 63.150 ;
        RECT 53.325 59.470 64.870 60.060 ;
        RECT 111.750 59.945 112.295 61.945 ;
        RECT 132.500 61.695 133.030 64.105 ;
        RECT 133.790 64.080 133.930 64.105 ;
        RECT 133.755 61.695 133.895 61.705 ;
        RECT 128.710 61.080 133.895 61.695 ;
        RECT 128.710 61.070 128.960 61.080 ;
        RECT 133.755 61.060 133.895 61.080 ;
        RECT 134.445 60.685 134.585 60.715 ;
        RECT 129.395 60.070 134.585 60.685 ;
        RECT 69.915 59.895 70.565 59.915 ;
        RECT 69.915 59.350 81.855 59.895 ;
        RECT 69.915 59.280 70.565 59.350 ;
        RECT 86.775 59.345 98.425 59.890 ;
        RECT 103.345 59.400 112.295 59.945 ;
        RECT 55.995 58.715 56.590 59.155 ;
        RECT 48.675 58.120 56.590 58.715 ;
        RECT 61.655 58.415 73.225 59.005 ;
        RECT 78.395 58.205 90.005 58.795 ;
        RECT 95.040 58.200 106.720 58.745 ;
        RECT 1.590 48.345 2.085 50.885 ;
        RECT 10.550 48.800 10.995 50.625 ;
        RECT 10.295 48.355 11.245 48.800 ;
        RECT 13.120 48.430 13.900 57.440 ;
        RECT 1.560 47.850 2.115 48.345 ;
        RECT 14.520 46.920 14.795 46.950 ;
        RECT 12.590 46.645 14.795 46.920 ;
        RECT 12.590 44.305 12.865 46.645 ;
        RECT 14.520 46.615 14.795 46.645 ;
        RECT 3.045 40.875 3.365 40.930 ;
        RECT 8.925 40.875 9.245 40.930 ;
        RECT 3.045 40.725 9.245 40.875 ;
        RECT 3.045 40.670 3.365 40.725 ;
        RECT 8.925 40.670 9.245 40.725 ;
        RECT 1.890 39.095 7.495 39.425 ;
        RECT 1.890 23.395 2.220 39.095 ;
        RECT 3.840 37.265 4.160 37.290 ;
        RECT 20.960 37.265 21.280 37.290 ;
        RECT 3.840 37.055 21.280 37.265 ;
        RECT 3.840 37.030 4.160 37.055 ;
        RECT 20.960 37.030 21.280 37.055 ;
        RECT 11.295 36.260 15.800 36.555 ;
        RECT 25.745 32.720 26.120 51.710 ;
        RECT 10.295 32.345 26.120 32.720 ;
        RECT 14.520 30.920 14.795 30.950 ;
        RECT 12.590 30.645 14.795 30.920 ;
        RECT 12.590 28.305 12.865 30.645 ;
        RECT 14.520 30.615 14.795 30.645 ;
        RECT 3.045 24.875 3.365 24.930 ;
        RECT 8.925 24.875 9.245 24.930 ;
        RECT 3.045 24.725 9.245 24.875 ;
        RECT 3.045 24.670 3.365 24.725 ;
        RECT 8.925 24.670 9.245 24.725 ;
        RECT 1.890 23.065 7.525 23.395 ;
        RECT 1.900 7.445 2.230 23.065 ;
        RECT 3.840 21.265 4.160 21.290 ;
        RECT 20.960 21.265 21.280 21.290 ;
        RECT 3.840 21.055 21.280 21.265 ;
        RECT 3.840 21.030 4.160 21.055 ;
        RECT 20.960 21.030 21.280 21.055 ;
        RECT 11.295 20.260 15.800 20.555 ;
        RECT 26.595 16.035 27.000 50.605 ;
        RECT 27.990 39.880 28.240 53.505 ;
        RECT 27.990 39.795 28.490 39.880 ;
        RECT 27.585 39.535 28.490 39.795 ;
        RECT 28.190 39.480 28.490 39.535 ;
        RECT 28.715 39.050 29.060 53.450 ;
        RECT 27.945 38.705 29.060 39.050 ;
        RECT 27.945 23.795 28.290 38.705 ;
        RECT 29.650 38.120 29.930 53.420 ;
        RECT 38.585 48.715 38.960 50.660 ;
        RECT 38.295 48.340 39.245 48.715 ;
        RECT 42.520 46.920 42.795 46.950 ;
        RECT 40.590 46.645 42.795 46.920 ;
        RECT 40.590 44.305 40.865 46.645 ;
        RECT 42.520 46.615 42.795 46.645 ;
        RECT 31.045 40.875 31.365 40.930 ;
        RECT 36.925 40.875 37.245 40.930 ;
        RECT 31.045 40.725 37.245 40.875 ;
        RECT 31.045 40.670 31.365 40.725 ;
        RECT 36.925 40.670 37.245 40.725 ;
        RECT 28.850 37.840 29.930 38.120 ;
        RECT 30.390 39.370 35.500 39.720 ;
        RECT 27.585 23.450 28.645 23.795 ;
        RECT 28.850 23.220 29.130 37.840 ;
        RECT 10.295 15.630 27.000 16.035 ;
        RECT 27.975 22.940 29.130 23.220 ;
        RECT 30.390 23.385 30.740 39.370 ;
        RECT 31.840 37.265 32.160 37.290 ;
        RECT 48.960 37.265 49.280 37.290 ;
        RECT 31.840 37.055 49.280 37.265 ;
        RECT 31.840 37.030 32.160 37.055 ;
        RECT 48.960 37.030 49.280 37.055 ;
        RECT 39.295 36.260 43.800 36.555 ;
        RECT 53.810 32.600 54.210 51.745 ;
        RECT 38.295 32.200 54.210 32.600 ;
        RECT 42.520 30.920 42.795 30.950 ;
        RECT 40.590 30.645 42.795 30.920 ;
        RECT 40.590 28.305 40.865 30.645 ;
        RECT 42.520 30.615 42.795 30.645 ;
        RECT 31.045 24.875 31.365 24.930 ;
        RECT 36.925 24.875 37.245 24.930 ;
        RECT 31.045 24.725 37.245 24.875 ;
        RECT 31.045 24.670 31.365 24.725 ;
        RECT 36.925 24.670 37.245 24.725 ;
        RECT 30.390 23.035 35.495 23.385 ;
        RECT 14.520 14.920 14.795 14.950 ;
        RECT 12.590 14.645 14.795 14.920 ;
        RECT 12.590 12.305 12.865 14.645 ;
        RECT 14.520 14.615 14.795 14.645 ;
        RECT 3.045 8.875 3.365 8.930 ;
        RECT 8.925 8.875 9.245 8.930 ;
        RECT 3.045 8.725 9.245 8.875 ;
        RECT 3.045 8.670 3.365 8.725 ;
        RECT 8.925 8.670 9.245 8.725 ;
        RECT 27.975 7.795 28.255 22.940 ;
        RECT 27.585 7.515 28.645 7.795 ;
        RECT 1.900 7.115 7.750 7.445 ;
        RECT 30.390 7.420 30.740 23.035 ;
        RECT 31.840 21.265 32.160 21.290 ;
        RECT 48.960 21.265 49.280 21.290 ;
        RECT 31.840 21.055 49.280 21.265 ;
        RECT 31.840 21.030 32.160 21.055 ;
        RECT 48.960 21.030 49.280 21.055 ;
        RECT 39.295 20.260 43.800 20.555 ;
        RECT 54.695 16.730 55.100 50.710 ;
        RECT 55.615 38.765 55.890 53.615 ;
        RECT 56.365 38.100 56.610 53.600 ;
        RECT 55.625 37.855 56.610 38.100 ;
        RECT 55.625 23.825 55.870 37.855 ;
        RECT 57.025 37.140 57.350 53.540 ;
        RECT 66.595 48.470 66.945 50.685 ;
        RECT 79.480 50.170 80.050 50.690 ;
        RECT 68.565 48.855 70.130 49.935 ;
        RECT 66.295 48.120 67.245 48.470 ;
        RECT 70.520 46.920 70.795 46.950 ;
        RECT 68.590 46.645 70.795 46.920 ;
        RECT 68.590 44.305 68.865 46.645 ;
        RECT 70.520 46.615 70.795 46.645 ;
        RECT 59.045 40.875 59.365 40.930 ;
        RECT 64.925 40.875 65.245 40.930 ;
        RECT 59.045 40.725 65.245 40.875 ;
        RECT 59.045 40.670 59.365 40.725 ;
        RECT 64.925 40.670 65.245 40.725 ;
        RECT 56.290 36.815 57.350 37.140 ;
        RECT 57.605 39.260 63.490 39.605 ;
        RECT 55.615 22.765 55.875 23.825 ;
        RECT 38.295 16.325 55.100 16.730 ;
        RECT 42.520 14.920 42.795 14.950 ;
        RECT 40.590 14.645 42.795 14.920 ;
        RECT 40.590 12.305 40.865 14.645 ;
        RECT 42.520 14.615 42.795 14.645 ;
        RECT 31.045 8.875 31.365 8.930 ;
        RECT 36.925 8.875 37.245 8.930 ;
        RECT 31.045 8.725 37.245 8.875 ;
        RECT 31.045 8.670 31.365 8.725 ;
        RECT 36.925 8.670 37.245 8.725 ;
        RECT 35.680 7.445 35.960 7.465 ;
        RECT 35.205 7.420 35.985 7.445 ;
        RECT 30.390 7.115 35.985 7.420 ;
        RECT 30.390 7.095 35.960 7.115 ;
        RECT 30.390 7.070 35.805 7.095 ;
        RECT 35.365 7.065 35.805 7.070 ;
        RECT 56.290 6.765 56.615 36.815 ;
        RECT 57.605 23.425 57.950 39.260 ;
        RECT 59.840 37.265 60.160 37.290 ;
        RECT 76.960 37.265 77.280 37.290 ;
        RECT 59.840 37.055 77.280 37.265 ;
        RECT 59.840 37.030 60.160 37.055 ;
        RECT 76.960 37.030 77.280 37.055 ;
        RECT 67.295 36.260 71.800 36.555 ;
        RECT 79.805 34.570 81.180 36.025 ;
        RECT 68.645 33.350 69.995 34.205 ;
        RECT 68.690 33.320 69.950 33.350 ;
        RECT 81.780 32.540 82.120 50.765 ;
        RECT 82.740 37.785 83.135 50.785 ;
        RECT 83.635 39.825 83.855 53.395 ;
        RECT 83.615 38.765 83.875 39.825 ;
        RECT 82.740 37.390 83.865 37.785 ;
        RECT 66.295 32.200 82.120 32.540 ;
        RECT 70.520 30.920 70.795 30.950 ;
        RECT 68.590 30.645 70.795 30.920 ;
        RECT 68.590 28.305 68.865 30.645 ;
        RECT 70.520 30.615 70.795 30.645 ;
        RECT 59.045 24.875 59.365 24.930 ;
        RECT 64.925 24.875 65.245 24.930 ;
        RECT 59.045 24.725 65.245 24.875 ;
        RECT 59.045 24.670 59.365 24.725 ;
        RECT 64.925 24.670 65.245 24.725 ;
        RECT 57.605 23.080 63.540 23.425 ;
        RECT 57.625 7.465 57.970 23.080 ;
        RECT 59.840 21.265 60.160 21.290 ;
        RECT 76.960 21.265 77.280 21.290 ;
        RECT 59.840 21.055 77.280 21.265 ;
        RECT 59.840 21.030 60.160 21.055 ;
        RECT 76.960 21.030 77.280 21.055 ;
        RECT 67.295 20.260 71.800 20.555 ;
        RECT 80.460 18.535 81.835 19.990 ;
        RECT 68.745 16.870 69.890 18.105 ;
        RECT 83.470 16.550 83.865 37.390 ;
        RECT 84.315 22.765 84.615 53.320 ;
        RECT 85.115 52.855 85.480 53.355 ;
        RECT 85.110 22.360 85.480 52.855 ;
        RECT 85.895 47.895 86.200 53.345 ;
        RECT 86.535 48.445 86.860 53.330 ;
        RECT 87.210 49.015 87.515 53.345 ;
        RECT 87.860 49.660 88.205 53.340 ;
        RECT 88.565 50.245 88.915 53.325 ;
        RECT 89.320 51.020 89.710 53.215 ;
        RECT 89.320 50.630 141.315 51.020 ;
        RECT 88.565 49.895 140.615 50.245 ;
        RECT 87.860 49.315 139.960 49.660 ;
        RECT 87.210 48.710 113.130 49.015 ;
        RECT 86.535 48.120 112.540 48.445 ;
        RECT 85.895 47.620 111.920 47.895 ;
        RECT 85.895 47.590 107.810 47.620 ;
        RECT 108.860 47.590 111.920 47.620 ;
        RECT 98.520 46.920 98.795 46.950 ;
        RECT 94.475 46.100 95.240 46.800 ;
        RECT 96.590 46.645 98.795 46.920 ;
        RECT 96.590 44.305 96.865 46.645 ;
        RECT 98.520 46.615 98.795 46.645 ;
        RECT 87.045 40.875 87.365 40.930 ;
        RECT 92.925 40.875 93.245 40.930 ;
        RECT 87.045 40.725 93.245 40.875 ;
        RECT 87.045 40.670 87.365 40.725 ;
        RECT 92.925 40.670 93.245 40.725 ;
        RECT 85.980 39.200 91.525 39.600 ;
        RECT 66.295 16.155 83.865 16.550 ;
        RECT 84.245 21.990 85.480 22.360 ;
        RECT 86.010 23.410 86.410 39.200 ;
        RECT 111.615 38.765 111.920 47.590 ;
        RECT 112.215 37.960 112.540 48.120 ;
        RECT 111.615 37.635 112.540 37.960 ;
        RECT 87.840 37.265 88.160 37.290 ;
        RECT 104.960 37.265 105.280 37.290 ;
        RECT 87.840 37.055 105.280 37.265 ;
        RECT 87.840 37.030 88.160 37.055 ;
        RECT 104.960 37.030 105.280 37.055 ;
        RECT 95.295 36.260 99.800 36.555 ;
        RECT 94.605 31.765 95.370 32.465 ;
        RECT 98.520 30.920 98.795 30.950 ;
        RECT 96.590 30.645 98.795 30.920 ;
        RECT 96.590 28.305 96.865 30.645 ;
        RECT 98.520 30.615 98.795 30.645 ;
        RECT 87.045 24.875 87.365 24.930 ;
        RECT 92.925 24.875 93.245 24.930 ;
        RECT 87.045 24.725 93.245 24.875 ;
        RECT 87.045 24.670 87.365 24.725 ;
        RECT 92.925 24.670 93.245 24.725 ;
        RECT 86.010 23.010 91.555 23.410 ;
        RECT 70.520 14.920 70.795 14.950 ;
        RECT 68.590 14.645 70.795 14.920 ;
        RECT 68.590 12.305 68.865 14.645 ;
        RECT 70.520 14.615 70.795 14.645 ;
        RECT 59.045 8.875 59.365 8.930 ;
        RECT 64.925 8.875 65.245 8.930 ;
        RECT 59.045 8.725 65.245 8.875 ;
        RECT 59.045 8.670 59.365 8.725 ;
        RECT 64.925 8.670 65.245 8.725 ;
        RECT 57.625 7.120 63.500 7.465 ;
        RECT 58.505 7.115 59.265 7.120 ;
        RECT 58.530 7.095 58.810 7.115 ;
        RECT 84.245 6.765 84.615 21.990 ;
        RECT 86.010 7.405 86.410 23.010 ;
        RECT 111.615 22.765 111.940 37.635 ;
        RECT 112.825 37.195 113.130 48.710 ;
        RECT 126.520 46.920 126.795 46.950 ;
        RECT 124.590 46.645 126.795 46.920 ;
        RECT 124.590 44.305 124.865 46.645 ;
        RECT 126.520 46.615 126.795 46.645 ;
        RECT 122.420 43.515 123.095 44.300 ;
        RECT 115.045 40.875 115.365 40.930 ;
        RECT 120.925 40.875 121.245 40.930 ;
        RECT 115.045 40.725 121.245 40.875 ;
        RECT 115.045 40.670 115.365 40.725 ;
        RECT 120.925 40.670 121.245 40.725 ;
        RECT 112.255 36.890 113.130 37.195 ;
        RECT 114.105 39.165 119.460 39.450 ;
        RECT 87.840 21.265 88.160 21.290 ;
        RECT 104.960 21.265 105.280 21.290 ;
        RECT 87.840 21.055 105.280 21.265 ;
        RECT 87.840 21.030 88.160 21.055 ;
        RECT 104.960 21.030 105.280 21.055 ;
        RECT 95.295 20.260 99.800 20.555 ;
        RECT 94.375 15.590 95.140 16.290 ;
        RECT 98.520 14.920 98.795 14.950 ;
        RECT 96.590 14.645 98.795 14.920 ;
        RECT 96.590 12.305 96.865 14.645 ;
        RECT 98.520 14.615 98.795 14.645 ;
        RECT 87.045 8.875 87.365 8.930 ;
        RECT 92.925 8.875 93.245 8.930 ;
        RECT 87.045 8.725 93.245 8.875 ;
        RECT 87.045 8.670 87.365 8.725 ;
        RECT 92.925 8.670 93.245 8.725 ;
        RECT 112.255 7.825 112.560 36.890 ;
        RECT 114.105 23.430 114.390 39.165 ;
        RECT 139.615 38.765 139.960 49.315 ;
        RECT 115.840 37.265 116.160 37.290 ;
        RECT 132.960 37.265 133.280 37.290 ;
        RECT 115.840 37.055 133.280 37.265 ;
        RECT 115.840 37.030 116.160 37.055 ;
        RECT 132.960 37.030 133.280 37.055 ;
        RECT 123.295 36.260 127.800 36.555 ;
        RECT 126.520 30.920 126.795 30.950 ;
        RECT 124.590 30.645 126.795 30.920 ;
        RECT 124.590 28.305 124.865 30.645 ;
        RECT 126.520 30.615 126.795 30.645 ;
        RECT 122.505 27.090 123.180 27.875 ;
        RECT 115.045 24.875 115.365 24.930 ;
        RECT 120.925 24.875 121.245 24.930 ;
        RECT 115.045 24.725 121.245 24.875 ;
        RECT 115.045 24.670 115.365 24.725 ;
        RECT 120.925 24.670 121.245 24.725 ;
        RECT 114.105 23.145 119.475 23.430 ;
        RECT 86.865 7.445 87.145 7.465 ;
        RECT 86.840 7.405 87.740 7.445 ;
        RECT 86.010 7.005 91.525 7.405 ;
        RECT 112.200 6.765 112.615 7.825 ;
        RECT 114.105 7.470 114.390 23.145 ;
        RECT 140.265 22.765 140.615 49.895 ;
        RECT 140.925 22.085 141.315 50.630 ;
        RECT 146.890 48.490 147.295 49.315 ;
        RECT 146.490 48.085 147.295 48.490 ;
        RECT 144.190 46.565 144.620 47.380 ;
        RECT 146.890 47.255 147.295 48.085 ;
        RECT 143.565 46.135 144.620 46.565 ;
        RECT 144.190 45.320 144.620 46.135 ;
        RECT 150.770 45.100 151.535 45.800 ;
        RECT 148.940 43.595 149.955 44.095 ;
        RECT 141.820 42.945 142.260 42.975 ;
        RECT 141.525 42.475 142.260 42.945 ;
        RECT 141.525 27.170 141.965 42.475 ;
        RECT 140.225 21.695 141.315 22.085 ;
        RECT 115.840 21.265 116.160 21.290 ;
        RECT 132.960 21.265 133.280 21.290 ;
        RECT 115.840 21.055 133.280 21.265 ;
        RECT 115.840 21.030 116.160 21.055 ;
        RECT 132.960 21.030 133.280 21.055 ;
        RECT 123.295 20.260 127.800 20.555 ;
        RECT 126.520 14.920 126.795 14.950 ;
        RECT 124.590 14.645 126.795 14.920 ;
        RECT 122.465 13.335 123.140 14.120 ;
        RECT 124.590 12.305 124.865 14.645 ;
        RECT 126.520 14.615 126.795 14.645 ;
        RECT 115.045 8.875 115.365 8.930 ;
        RECT 120.925 8.875 121.245 8.930 ;
        RECT 115.045 8.725 121.245 8.875 ;
        RECT 115.045 8.670 115.365 8.725 ;
        RECT 120.925 8.670 121.245 8.725 ;
        RECT 114.105 7.185 119.465 7.470 ;
        RECT 114.800 7.115 115.590 7.185 ;
        RECT 114.825 7.095 115.105 7.115 ;
        RECT 140.225 6.765 140.615 21.695 ;
        RECT 142.380 13.435 142.880 41.065 ;
        RECT 3.840 5.265 4.160 5.290 ;
        RECT 20.960 5.265 21.280 5.290 ;
        RECT 3.840 5.055 21.280 5.265 ;
        RECT 3.840 5.030 4.160 5.055 ;
        RECT 20.960 5.030 21.280 5.055 ;
        RECT 31.840 5.265 32.160 5.290 ;
        RECT 48.960 5.265 49.280 5.290 ;
        RECT 31.840 5.055 49.280 5.265 ;
        RECT 31.840 5.030 32.160 5.055 ;
        RECT 48.960 5.030 49.280 5.055 ;
        RECT 59.840 5.265 60.160 5.290 ;
        RECT 76.960 5.265 77.280 5.290 ;
        RECT 59.840 5.055 77.280 5.265 ;
        RECT 59.840 5.030 60.160 5.055 ;
        RECT 76.960 5.030 77.280 5.055 ;
        RECT 87.840 5.265 88.160 5.290 ;
        RECT 104.960 5.265 105.280 5.290 ;
        RECT 87.840 5.055 105.280 5.265 ;
        RECT 87.840 5.030 88.160 5.055 ;
        RECT 104.960 5.030 105.280 5.055 ;
        RECT 115.840 5.265 116.160 5.290 ;
        RECT 132.960 5.265 133.280 5.290 ;
        RECT 115.840 5.055 133.280 5.265 ;
        RECT 115.840 5.030 116.160 5.055 ;
        RECT 132.960 5.030 133.280 5.055 ;
        RECT 11.295 4.260 15.800 4.555 ;
        RECT 39.295 4.260 43.800 4.555 ;
        RECT 67.295 4.260 71.800 4.555 ;
        RECT 80.415 2.885 81.790 4.340 ;
        RECT 95.295 4.260 99.800 4.555 ;
        RECT 123.295 4.260 127.800 4.555 ;
      LAYER met3 ;
        RECT 8.720 223.470 9.220 223.620 ;
        RECT 83.785 223.470 84.115 223.485 ;
        RECT 8.720 223.170 84.115 223.470 ;
        RECT 8.720 223.020 9.220 223.170 ;
        RECT 83.785 223.155 84.115 223.170 ;
        RECT 8.720 220.070 9.220 220.220 ;
        RECT 16.165 220.070 16.495 220.085 ;
        RECT 8.720 219.770 16.495 220.070 ;
        RECT 8.720 219.620 9.220 219.770 ;
        RECT 16.165 219.755 16.495 219.770 ;
        RECT 8.720 216.670 9.220 216.820 ;
        RECT 8.720 216.370 22.230 216.670 ;
        RECT 8.720 216.220 9.220 216.370 ;
        RECT 21.930 214.630 22.230 216.370 ;
        RECT 89.765 214.630 90.095 214.645 ;
        RECT 21.930 214.330 90.095 214.630 ;
        RECT 89.765 214.315 90.095 214.330 ;
        RECT 8.720 213.270 9.220 213.420 ;
        RECT 23.985 213.270 24.315 213.285 ;
        RECT 8.720 212.970 24.315 213.270 ;
        RECT 8.720 212.820 9.220 212.970 ;
        RECT 23.985 212.955 24.315 212.970 ;
        RECT 106.550 212.615 108.130 212.945 ;
        RECT 17.545 211.230 17.875 211.245 ;
        RECT 22.350 211.230 22.730 211.240 ;
        RECT 17.545 210.930 22.730 211.230 ;
        RECT 17.545 210.915 17.875 210.930 ;
        RECT 22.350 210.920 22.730 210.930 ;
        RECT 55.725 211.230 56.055 211.245 ;
        RECT 76.885 211.230 77.215 211.245 ;
        RECT 55.725 210.930 77.215 211.230 ;
        RECT 55.725 210.915 56.055 210.930 ;
        RECT 76.885 210.915 77.215 210.930 ;
        RECT 18.005 210.550 18.335 210.565 ;
        RECT 56.390 210.550 56.770 210.560 ;
        RECT 18.005 210.250 56.770 210.550 ;
        RECT 18.005 210.235 18.335 210.250 ;
        RECT 56.390 210.240 56.770 210.250 ;
        RECT 81.485 210.550 81.815 210.565 ;
        RECT 88.385 210.550 88.715 210.565 ;
        RECT 81.485 210.250 88.715 210.550 ;
        RECT 81.485 210.235 81.815 210.250 ;
        RECT 88.385 210.235 88.715 210.250 ;
        RECT 8.720 209.870 9.220 210.020 ;
        RECT 109.850 209.895 111.430 210.225 ;
        RECT 80.565 209.870 80.895 209.885 ;
        RECT 8.720 209.570 80.895 209.870 ;
        RECT 8.720 209.420 9.220 209.570 ;
        RECT 80.565 209.555 80.895 209.570 ;
        RECT 128.405 209.870 128.735 209.885 ;
        RECT 131.980 209.870 132.480 210.020 ;
        RECT 128.405 209.570 132.480 209.870 ;
        RECT 128.405 209.555 128.735 209.570 ;
        RECT 131.980 209.420 132.480 209.570 ;
        RECT 38.910 209.190 39.290 209.200 ;
        RECT 64.925 209.190 65.255 209.205 ;
        RECT 78.265 209.190 78.595 209.205 ;
        RECT 21.930 208.890 78.595 209.190 ;
        RECT 20.305 207.830 20.635 207.845 ;
        RECT 21.930 207.830 22.230 208.890 ;
        RECT 38.910 208.880 39.290 208.890 ;
        RECT 64.925 208.875 65.255 208.890 ;
        RECT 78.265 208.875 78.595 208.890 ;
        RECT 61.245 208.510 61.575 208.525 ;
        RECT 70.905 208.510 71.235 208.525 ;
        RECT 61.245 208.210 71.235 208.510 ;
        RECT 61.245 208.195 61.575 208.210 ;
        RECT 70.905 208.195 71.235 208.210 ;
        RECT 89.305 208.510 89.635 208.525 ;
        RECT 94.365 208.510 94.695 208.525 ;
        RECT 89.305 208.210 94.695 208.510 ;
        RECT 89.305 208.195 89.635 208.210 ;
        RECT 94.365 208.195 94.695 208.210 ;
        RECT 20.305 207.530 22.230 207.830 ;
        RECT 41.005 207.830 41.335 207.845 ;
        RECT 65.845 207.830 66.175 207.845 ;
        RECT 41.005 207.530 66.175 207.830 ;
        RECT 20.305 207.515 20.635 207.530 ;
        RECT 41.005 207.515 41.335 207.530 ;
        RECT 65.845 207.515 66.175 207.530 ;
        RECT 106.550 207.175 108.130 207.505 ;
        RECT 56.645 207.150 56.975 207.165 ;
        RECT 67.685 207.150 68.015 207.165 ;
        RECT 56.645 206.850 68.015 207.150 ;
        RECT 56.645 206.835 56.975 206.850 ;
        RECT 67.685 206.835 68.015 206.850 ;
        RECT 8.720 206.470 9.220 206.620 ;
        RECT 60.785 206.470 61.115 206.485 ;
        RECT 8.720 206.170 61.115 206.470 ;
        RECT 8.720 206.020 9.220 206.170 ;
        RECT 60.785 206.155 61.115 206.170 ;
        RECT 62.165 206.470 62.495 206.485 ;
        RECT 109.085 206.470 109.415 206.485 ;
        RECT 62.165 206.170 109.415 206.470 ;
        RECT 62.165 206.155 62.495 206.170 ;
        RECT 109.085 206.155 109.415 206.170 ;
        RECT 54.805 205.800 55.135 205.805 ;
        RECT 54.550 205.790 55.135 205.800 ;
        RECT 66.305 205.790 66.635 205.805 ;
        RECT 81.945 205.790 82.275 205.805 ;
        RECT 54.550 205.490 55.360 205.790 ;
        RECT 66.305 205.490 82.275 205.790 ;
        RECT 54.550 205.480 55.135 205.490 ;
        RECT 54.805 205.475 55.135 205.480 ;
        RECT 66.305 205.475 66.635 205.490 ;
        RECT 81.945 205.475 82.275 205.490 ;
        RECT 47.445 205.110 47.775 205.125 ;
        RECT 52.045 205.110 52.375 205.125 ;
        RECT 82.865 205.110 83.195 205.125 ;
        RECT 86.085 205.110 86.415 205.125 ;
        RECT 47.445 204.810 86.415 205.110 ;
        RECT 47.445 204.795 47.775 204.810 ;
        RECT 52.045 204.795 52.375 204.810 ;
        RECT 82.865 204.795 83.195 204.810 ;
        RECT 86.085 204.795 86.415 204.810 ;
        RECT 109.850 204.455 111.430 204.785 ;
        RECT 36.865 204.430 37.195 204.445 ;
        RECT 59.865 204.430 60.195 204.445 ;
        RECT 36.865 204.130 60.195 204.430 ;
        RECT 36.865 204.115 37.195 204.130 ;
        RECT 59.865 204.115 60.195 204.130 ;
        RECT 64.925 204.430 65.255 204.445 ;
        RECT 70.445 204.430 70.775 204.445 ;
        RECT 72.745 204.430 73.075 204.445 ;
        RECT 64.925 204.130 73.075 204.430 ;
        RECT 64.925 204.115 65.255 204.130 ;
        RECT 70.445 204.115 70.775 204.130 ;
        RECT 72.745 204.115 73.075 204.130 ;
        RECT 41.925 203.750 42.255 203.765 ;
        RECT 50.205 203.750 50.535 203.765 ;
        RECT 41.925 203.450 50.535 203.750 ;
        RECT 41.925 203.435 42.255 203.450 ;
        RECT 50.205 203.435 50.535 203.450 ;
        RECT 51.125 203.750 51.455 203.765 ;
        RECT 71.365 203.750 71.695 203.765 ;
        RECT 51.125 203.450 71.695 203.750 ;
        RECT 51.125 203.435 51.455 203.450 ;
        RECT 71.365 203.435 71.695 203.450 ;
        RECT 85.625 203.750 85.955 203.765 ;
        RECT 92.065 203.750 92.395 203.765 ;
        RECT 85.625 203.450 92.395 203.750 ;
        RECT 85.625 203.435 85.955 203.450 ;
        RECT 92.065 203.435 92.395 203.450 ;
        RECT 8.720 203.070 9.220 203.220 ;
        RECT 65.385 203.070 65.715 203.085 ;
        RECT 8.720 202.770 65.715 203.070 ;
        RECT 8.720 202.620 9.220 202.770 ;
        RECT 65.385 202.755 65.715 202.770 ;
        RECT 69.525 203.070 69.855 203.085 ;
        RECT 73.665 203.070 73.995 203.085 ;
        RECT 69.525 202.770 73.995 203.070 ;
        RECT 69.525 202.755 69.855 202.770 ;
        RECT 73.665 202.755 73.995 202.770 ;
        RECT 52.505 202.400 52.835 202.405 ;
        RECT 52.505 202.390 53.090 202.400 ;
        RECT 52.280 202.090 53.090 202.390 ;
        RECT 52.505 202.080 53.090 202.090 ;
        RECT 53.630 202.390 54.010 202.400 ;
        RECT 54.345 202.390 54.675 202.405 ;
        RECT 53.630 202.090 54.675 202.390 ;
        RECT 53.630 202.080 54.010 202.090 ;
        RECT 52.505 202.075 52.835 202.080 ;
        RECT 54.345 202.075 54.675 202.090 ;
        RECT 67.685 202.390 68.015 202.405 ;
        RECT 69.985 202.390 70.315 202.405 ;
        RECT 67.685 202.090 70.315 202.390 ;
        RECT 67.685 202.075 68.015 202.090 ;
        RECT 69.985 202.075 70.315 202.090 ;
        RECT 106.550 201.735 108.130 202.065 ;
        RECT 45.145 201.710 45.475 201.725 ;
        RECT 64.465 201.710 64.795 201.725 ;
        RECT 45.145 201.410 64.795 201.710 ;
        RECT 45.145 201.395 45.475 201.410 ;
        RECT 64.465 201.395 64.795 201.410 ;
        RECT 66.305 201.710 66.635 201.725 ;
        RECT 70.905 201.710 71.235 201.725 ;
        RECT 66.305 201.410 71.235 201.710 ;
        RECT 66.305 201.395 66.635 201.410 ;
        RECT 70.905 201.395 71.235 201.410 ;
        RECT 42.385 201.030 42.715 201.045 ;
        RECT 58.485 201.030 58.815 201.045 ;
        RECT 42.385 200.730 58.815 201.030 ;
        RECT 42.385 200.715 42.715 200.730 ;
        RECT 58.485 200.715 58.815 200.730 ;
        RECT 60.990 201.030 61.370 201.040 ;
        RECT 61.705 201.030 62.035 201.045 ;
        RECT 60.990 200.730 62.035 201.030 ;
        RECT 60.990 200.720 61.370 200.730 ;
        RECT 61.705 200.715 62.035 200.730 ;
        RECT 65.845 201.030 66.175 201.045 ;
        RECT 106.325 201.030 106.655 201.045 ;
        RECT 65.845 200.730 106.655 201.030 ;
        RECT 65.845 200.715 66.175 200.730 ;
        RECT 106.325 200.715 106.655 200.730 ;
        RECT 45.605 200.350 45.935 200.365 ;
        RECT 66.305 200.350 66.635 200.365 ;
        RECT 45.605 200.050 66.635 200.350 ;
        RECT 45.605 200.035 45.935 200.050 ;
        RECT 66.305 200.035 66.635 200.050 ;
        RECT 69.985 200.350 70.315 200.365 ;
        RECT 70.905 200.350 71.235 200.365 ;
        RECT 86.085 200.360 86.415 200.365 ;
        RECT 69.985 200.050 71.235 200.350 ;
        RECT 69.985 200.035 70.315 200.050 ;
        RECT 70.905 200.035 71.235 200.050 ;
        RECT 85.830 200.350 86.415 200.360 ;
        RECT 92.985 200.350 93.315 200.365 ;
        RECT 85.830 200.050 93.315 200.350 ;
        RECT 85.830 200.040 86.415 200.050 ;
        RECT 86.085 200.035 86.415 200.040 ;
        RECT 92.985 200.035 93.315 200.050 ;
        RECT 8.720 199.670 9.220 199.820 ;
        RECT 62.165 199.670 62.495 199.685 ;
        RECT 8.720 199.370 62.495 199.670 ;
        RECT 8.720 199.220 9.220 199.370 ;
        RECT 62.165 199.355 62.495 199.370 ;
        RECT 69.985 199.670 70.315 199.685 ;
        RECT 104.025 199.670 104.355 199.685 ;
        RECT 69.985 199.370 104.355 199.670 ;
        RECT 69.985 199.355 70.315 199.370 ;
        RECT 104.025 199.355 104.355 199.370 ;
        RECT 129.325 199.670 129.655 199.685 ;
        RECT 131.980 199.670 132.480 199.820 ;
        RECT 129.325 199.370 132.480 199.670 ;
        RECT 129.325 199.355 129.655 199.370 ;
        RECT 109.850 199.015 111.430 199.345 ;
        RECT 131.980 199.220 132.480 199.370 ;
        RECT 37.785 198.990 38.115 199.005 ;
        RECT 46.985 198.990 47.315 199.005 ;
        RECT 56.645 198.990 56.975 199.005 ;
        RECT 37.785 198.690 56.975 198.990 ;
        RECT 37.785 198.675 38.115 198.690 ;
        RECT 46.985 198.675 47.315 198.690 ;
        RECT 56.645 198.675 56.975 198.690 ;
        RECT 88.385 198.990 88.715 199.005 ;
        RECT 96.205 198.990 96.535 199.005 ;
        RECT 88.385 198.690 96.535 198.990 ;
        RECT 88.385 198.675 88.715 198.690 ;
        RECT 96.205 198.675 96.535 198.690 ;
        RECT 46.985 198.310 47.315 198.325 ;
        RECT 47.905 198.310 48.235 198.325 ;
        RECT 53.885 198.310 54.215 198.325 ;
        RECT 46.985 198.010 54.215 198.310 ;
        RECT 46.985 197.995 47.315 198.010 ;
        RECT 47.905 197.995 48.235 198.010 ;
        RECT 53.885 197.995 54.215 198.010 ;
        RECT 55.725 198.310 56.055 198.325 ;
        RECT 58.230 198.310 58.610 198.320 ;
        RECT 58.945 198.310 59.275 198.325 ;
        RECT 55.725 198.010 59.275 198.310 ;
        RECT 55.725 197.995 56.055 198.010 ;
        RECT 58.230 198.000 58.610 198.010 ;
        RECT 58.945 197.995 59.275 198.010 ;
        RECT 96.205 198.310 96.535 198.325 ;
        RECT 97.125 198.310 97.455 198.325 ;
        RECT 96.205 198.010 97.455 198.310 ;
        RECT 96.205 197.995 96.535 198.010 ;
        RECT 97.125 197.995 97.455 198.010 ;
        RECT 23.985 197.630 24.315 197.645 ;
        RECT 42.590 197.630 42.970 197.640 ;
        RECT 23.985 197.330 42.970 197.630 ;
        RECT 23.985 197.315 24.315 197.330 ;
        RECT 42.590 197.320 42.970 197.330 ;
        RECT 47.905 197.630 48.235 197.645 ;
        RECT 49.285 197.630 49.615 197.645 ;
        RECT 52.505 197.630 52.835 197.645 ;
        RECT 47.905 197.330 52.835 197.630 ;
        RECT 47.905 197.315 48.235 197.330 ;
        RECT 49.285 197.315 49.615 197.330 ;
        RECT 52.505 197.315 52.835 197.330 ;
        RECT 55.265 197.630 55.595 197.645 ;
        RECT 60.785 197.630 61.115 197.645 ;
        RECT 76.425 197.630 76.755 197.645 ;
        RECT 55.265 197.330 76.755 197.630 ;
        RECT 55.265 197.315 55.595 197.330 ;
        RECT 60.785 197.315 61.115 197.330 ;
        RECT 76.425 197.315 76.755 197.330 ;
        RECT 91.145 197.630 91.475 197.645 ;
        RECT 95.285 197.630 95.615 197.645 ;
        RECT 91.145 197.330 95.615 197.630 ;
        RECT 91.145 197.315 91.475 197.330 ;
        RECT 95.285 197.315 95.615 197.330 ;
        RECT 97.125 197.630 97.455 197.645 ;
        RECT 102.645 197.630 102.975 197.645 ;
        RECT 112.305 197.630 112.635 197.645 ;
        RECT 97.125 197.330 112.635 197.630 ;
        RECT 97.125 197.315 97.455 197.330 ;
        RECT 102.645 197.315 102.975 197.330 ;
        RECT 112.305 197.315 112.635 197.330 ;
        RECT 41.465 196.950 41.795 196.965 ;
        RECT 61.705 196.950 62.035 196.965 ;
        RECT 75.965 196.950 76.295 196.965 ;
        RECT 41.465 196.650 76.295 196.950 ;
        RECT 41.465 196.635 41.795 196.650 ;
        RECT 61.705 196.635 62.035 196.650 ;
        RECT 75.965 196.635 76.295 196.650 ;
        RECT 92.985 196.950 93.315 196.965 ;
        RECT 99.885 196.950 100.215 196.965 ;
        RECT 92.985 196.650 100.215 196.950 ;
        RECT 92.985 196.635 93.315 196.650 ;
        RECT 99.885 196.635 100.215 196.650 ;
        RECT 8.720 196.270 9.220 196.420 ;
        RECT 106.550 196.295 108.130 196.625 ;
        RECT 63.545 196.270 63.875 196.285 ;
        RECT 8.720 195.970 63.875 196.270 ;
        RECT 8.720 195.820 9.220 195.970 ;
        RECT 63.545 195.955 63.875 195.970 ;
        RECT 67.225 196.270 67.555 196.285 ;
        RECT 81.485 196.270 81.815 196.285 ;
        RECT 67.225 195.970 81.815 196.270 ;
        RECT 67.225 195.955 67.555 195.970 ;
        RECT 81.485 195.955 81.815 195.970 ;
        RECT 97.125 196.270 97.455 196.285 ;
        RECT 105.405 196.270 105.735 196.285 ;
        RECT 97.125 195.970 105.735 196.270 ;
        RECT 97.125 195.955 97.455 195.970 ;
        RECT 105.405 195.955 105.735 195.970 ;
        RECT 128.405 196.270 128.735 196.285 ;
        RECT 131.980 196.270 132.480 196.420 ;
        RECT 128.405 195.970 132.480 196.270 ;
        RECT 128.405 195.955 128.735 195.970 ;
        RECT 131.980 195.820 132.480 195.970 ;
        RECT 39.830 195.590 40.210 195.600 ;
        RECT 42.385 195.590 42.715 195.605 ;
        RECT 39.830 195.290 42.715 195.590 ;
        RECT 39.830 195.280 40.210 195.290 ;
        RECT 42.385 195.275 42.715 195.290 ;
        RECT 46.065 195.590 46.395 195.605 ;
        RECT 49.745 195.590 50.075 195.605 ;
        RECT 46.065 195.290 50.075 195.590 ;
        RECT 46.065 195.275 46.395 195.290 ;
        RECT 49.745 195.275 50.075 195.290 ;
        RECT 56.390 195.590 56.770 195.600 ;
        RECT 60.325 195.590 60.655 195.605 ;
        RECT 56.390 195.290 60.655 195.590 ;
        RECT 56.390 195.280 56.770 195.290 ;
        RECT 60.325 195.275 60.655 195.290 ;
        RECT 61.910 195.590 62.290 195.600 ;
        RECT 71.365 195.590 71.695 195.605 ;
        RECT 95.745 195.590 96.075 195.605 ;
        RECT 61.910 195.290 96.075 195.590 ;
        RECT 61.910 195.280 62.290 195.290 ;
        RECT 71.365 195.275 71.695 195.290 ;
        RECT 95.745 195.275 96.075 195.290 ;
        RECT 17.545 194.910 17.875 194.925 ;
        RECT 62.625 194.910 62.955 194.925 ;
        RECT 78.725 194.910 79.055 194.925 ;
        RECT 17.545 194.610 79.055 194.910 ;
        RECT 17.545 194.595 17.875 194.610 ;
        RECT 62.625 194.595 62.955 194.610 ;
        RECT 78.725 194.595 79.055 194.610 ;
        RECT 42.590 194.230 42.970 194.240 ;
        RECT 62.625 194.230 62.955 194.245 ;
        RECT 42.590 193.930 62.955 194.230 ;
        RECT 42.590 193.920 42.970 193.930 ;
        RECT 62.625 193.915 62.955 193.930 ;
        RECT 63.545 194.240 63.875 194.245 ;
        RECT 63.545 194.230 64.130 194.240 ;
        RECT 77.805 194.230 78.135 194.245 ;
        RECT 104.025 194.230 104.355 194.245 ;
        RECT 63.545 193.930 64.330 194.230 ;
        RECT 77.805 193.930 104.355 194.230 ;
        RECT 63.545 193.920 64.130 193.930 ;
        RECT 63.545 193.915 63.875 193.920 ;
        RECT 77.805 193.915 78.135 193.930 ;
        RECT 104.025 193.915 104.355 193.930 ;
        RECT 109.850 193.575 111.430 193.905 ;
        RECT 38.245 193.560 38.575 193.565 ;
        RECT 37.990 193.550 38.575 193.560 ;
        RECT 37.790 193.250 38.575 193.550 ;
        RECT 37.990 193.240 38.575 193.250 ;
        RECT 38.245 193.235 38.575 193.240 ;
        RECT 39.165 193.550 39.495 193.565 ;
        RECT 49.030 193.550 49.410 193.560 ;
        RECT 39.165 193.250 49.410 193.550 ;
        RECT 39.165 193.235 39.495 193.250 ;
        RECT 49.030 193.240 49.410 193.250 ;
        RECT 52.505 193.550 52.835 193.565 ;
        RECT 89.765 193.550 90.095 193.565 ;
        RECT 52.505 193.250 90.095 193.550 ;
        RECT 52.505 193.235 52.835 193.250 ;
        RECT 89.765 193.235 90.095 193.250 ;
        RECT 8.720 192.870 9.220 193.020 ;
        RECT 63.545 192.870 63.875 192.885 ;
        RECT 8.720 192.570 63.875 192.870 ;
        RECT 8.720 192.420 9.220 192.570 ;
        RECT 63.545 192.555 63.875 192.570 ;
        RECT 128.405 192.870 128.735 192.885 ;
        RECT 131.980 192.870 132.480 193.020 ;
        RECT 128.405 192.570 132.480 192.870 ;
        RECT 128.405 192.555 128.735 192.570 ;
        RECT 131.980 192.420 132.480 192.570 ;
        RECT 18.465 192.190 18.795 192.205 ;
        RECT 32.725 192.190 33.055 192.205 ;
        RECT 18.465 191.890 33.055 192.190 ;
        RECT 18.465 191.875 18.795 191.890 ;
        RECT 32.725 191.875 33.055 191.890 ;
        RECT 37.785 192.190 38.115 192.205 ;
        RECT 39.625 192.190 39.955 192.205 ;
        RECT 41.925 192.190 42.255 192.205 ;
        RECT 37.785 191.890 42.255 192.190 ;
        RECT 37.785 191.875 38.115 191.890 ;
        RECT 39.625 191.875 39.955 191.890 ;
        RECT 41.925 191.875 42.255 191.890 ;
        RECT 51.585 192.190 51.915 192.205 ;
        RECT 57.565 192.200 57.895 192.205 ;
        RECT 53.630 192.190 54.010 192.200 ;
        RECT 51.585 191.890 54.010 192.190 ;
        RECT 51.585 191.875 51.915 191.890 ;
        RECT 53.630 191.880 54.010 191.890 ;
        RECT 57.310 192.190 57.895 192.200 ;
        RECT 75.045 192.190 75.375 192.205 ;
        RECT 113.225 192.190 113.555 192.205 ;
        RECT 116.905 192.190 117.235 192.205 ;
        RECT 57.310 191.890 58.120 192.190 ;
        RECT 75.045 191.890 117.235 192.190 ;
        RECT 57.310 191.880 57.895 191.890 ;
        RECT 57.565 191.875 57.895 191.880 ;
        RECT 75.045 191.875 75.375 191.890 ;
        RECT 113.225 191.875 113.555 191.890 ;
        RECT 116.905 191.875 117.235 191.890 ;
        RECT 17.085 191.510 17.415 191.525 ;
        RECT 66.765 191.510 67.095 191.525 ;
        RECT 17.085 191.210 67.095 191.510 ;
        RECT 17.085 191.195 17.415 191.210 ;
        RECT 66.765 191.195 67.095 191.210 ;
        RECT 68.145 191.510 68.475 191.525 ;
        RECT 75.505 191.510 75.835 191.525 ;
        RECT 68.145 191.210 75.835 191.510 ;
        RECT 68.145 191.195 68.475 191.210 ;
        RECT 75.505 191.195 75.835 191.210 ;
        RECT 77.805 191.510 78.135 191.525 ;
        RECT 79.645 191.510 79.975 191.525 ;
        RECT 77.805 191.210 79.975 191.510 ;
        RECT 77.805 191.195 78.135 191.210 ;
        RECT 79.645 191.195 79.975 191.210 ;
        RECT 106.550 190.855 108.130 191.185 ;
        RECT 28.125 190.830 28.455 190.845 ;
        RECT 65.385 190.830 65.715 190.845 ;
        RECT 69.065 190.830 69.395 190.845 ;
        RECT 28.125 190.530 69.395 190.830 ;
        RECT 28.125 190.515 28.455 190.530 ;
        RECT 65.385 190.515 65.715 190.530 ;
        RECT 69.065 190.515 69.395 190.530 ;
        RECT 76.885 190.830 77.215 190.845 ;
        RECT 84.705 190.830 85.035 190.845 ;
        RECT 76.885 190.530 85.035 190.830 ;
        RECT 76.885 190.515 77.215 190.530 ;
        RECT 84.705 190.515 85.035 190.530 ;
        RECT 27.665 190.150 27.995 190.165 ;
        RECT 51.125 190.150 51.455 190.165 ;
        RECT 27.665 189.850 51.455 190.150 ;
        RECT 27.665 189.835 27.995 189.850 ;
        RECT 51.125 189.835 51.455 189.850 ;
        RECT 58.945 190.150 59.275 190.165 ;
        RECT 61.910 190.150 62.290 190.160 ;
        RECT 58.945 189.850 62.290 190.150 ;
        RECT 58.945 189.835 59.275 189.850 ;
        RECT 61.910 189.840 62.290 189.850 ;
        RECT 65.385 190.150 65.715 190.165 ;
        RECT 66.305 190.150 66.635 190.165 ;
        RECT 65.385 189.850 66.635 190.150 ;
        RECT 65.385 189.835 65.715 189.850 ;
        RECT 66.305 189.835 66.635 189.850 ;
        RECT 8.720 189.470 9.220 189.620 ;
        RECT 48.365 189.470 48.695 189.485 ;
        RECT 49.285 189.480 49.615 189.485 ;
        RECT 8.720 189.170 48.695 189.470 ;
        RECT 8.720 189.020 9.220 189.170 ;
        RECT 48.365 189.155 48.695 189.170 ;
        RECT 49.030 189.470 49.615 189.480 ;
        RECT 50.665 189.470 50.995 189.485 ;
        RECT 68.605 189.470 68.935 189.485 ;
        RECT 49.030 189.170 49.840 189.470 ;
        RECT 50.665 189.170 68.935 189.470 ;
        RECT 49.030 189.160 49.615 189.170 ;
        RECT 49.285 189.155 49.615 189.160 ;
        RECT 50.665 189.155 50.995 189.170 ;
        RECT 68.605 189.155 68.935 189.170 ;
        RECT 131.165 189.470 131.495 189.485 ;
        RECT 131.980 189.470 132.480 189.620 ;
        RECT 131.165 189.170 132.480 189.470 ;
        RECT 131.165 189.155 131.495 189.170 ;
        RECT 131.980 189.020 132.480 189.170 ;
        RECT 22.605 188.790 22.935 188.805 ;
        RECT 50.205 188.790 50.535 188.805 ;
        RECT 22.605 188.490 50.535 188.790 ;
        RECT 22.605 188.475 22.935 188.490 ;
        RECT 50.205 188.475 50.535 188.490 ;
        RECT 52.965 188.790 53.295 188.805 ;
        RECT 54.550 188.790 54.930 188.800 ;
        RECT 52.965 188.490 54.930 188.790 ;
        RECT 52.965 188.475 53.295 188.490 ;
        RECT 54.550 188.480 54.930 188.490 ;
        RECT 55.725 188.790 56.055 188.805 ;
        RECT 73.665 188.790 73.995 188.805 ;
        RECT 55.725 188.490 73.995 188.790 ;
        RECT 55.725 188.475 56.055 188.490 ;
        RECT 73.665 188.475 73.995 188.490 ;
        RECT 109.850 188.135 111.430 188.465 ;
        RECT 45.145 188.110 45.475 188.125 ;
        RECT 52.045 188.110 52.375 188.125 ;
        RECT 45.145 187.810 52.375 188.110 ;
        RECT 45.145 187.795 45.475 187.810 ;
        RECT 52.045 187.795 52.375 187.810 ;
        RECT 57.105 188.110 57.435 188.125 ;
        RECT 69.525 188.110 69.855 188.125 ;
        RECT 57.105 187.810 69.855 188.110 ;
        RECT 57.105 187.795 57.435 187.810 ;
        RECT 69.525 187.795 69.855 187.810 ;
        RECT 20.305 187.430 20.635 187.445 ;
        RECT 67.685 187.430 68.015 187.445 ;
        RECT 20.305 187.130 68.015 187.430 ;
        RECT 20.305 187.115 20.635 187.130 ;
        RECT 67.685 187.115 68.015 187.130 ;
        RECT 36.865 186.750 37.195 186.765 ;
        RECT 77.345 186.750 77.675 186.765 ;
        RECT 36.865 186.450 77.675 186.750 ;
        RECT 36.865 186.435 37.195 186.450 ;
        RECT 77.345 186.435 77.675 186.450 ;
        RECT 85.165 186.750 85.495 186.765 ;
        RECT 87.925 186.750 88.255 186.765 ;
        RECT 85.165 186.450 88.255 186.750 ;
        RECT 85.165 186.435 85.495 186.450 ;
        RECT 87.925 186.435 88.255 186.450 ;
        RECT 8.720 186.070 9.220 186.220 ;
        RECT 57.565 186.070 57.895 186.085 ;
        RECT 8.720 185.770 57.895 186.070 ;
        RECT 8.720 185.620 9.220 185.770 ;
        RECT 57.565 185.755 57.895 185.770 ;
        RECT 130.245 186.070 130.575 186.085 ;
        RECT 131.980 186.070 132.480 186.220 ;
        RECT 130.245 185.770 132.480 186.070 ;
        RECT 130.245 185.755 130.575 185.770 ;
        RECT 106.550 185.415 108.130 185.745 ;
        RECT 131.980 185.620 132.480 185.770 ;
        RECT 34.105 185.390 34.435 185.405 ;
        RECT 42.385 185.390 42.715 185.405 ;
        RECT 34.105 185.090 42.715 185.390 ;
        RECT 34.105 185.075 34.435 185.090 ;
        RECT 42.385 185.075 42.715 185.090 ;
        RECT 44.225 185.390 44.555 185.405 ;
        RECT 45.605 185.390 45.935 185.405 ;
        RECT 52.505 185.400 52.835 185.405 ;
        RECT 52.505 185.390 53.090 185.400 ;
        RECT 44.225 185.090 45.935 185.390 ;
        RECT 52.280 185.090 53.090 185.390 ;
        RECT 44.225 185.075 44.555 185.090 ;
        RECT 45.605 185.075 45.935 185.090 ;
        RECT 52.505 185.080 53.090 185.090 ;
        RECT 58.025 185.390 58.355 185.405 ;
        RECT 81.945 185.390 82.275 185.405 ;
        RECT 58.025 185.090 82.275 185.390 ;
        RECT 52.505 185.075 52.835 185.080 ;
        RECT 58.025 185.075 58.355 185.090 ;
        RECT 81.945 185.075 82.275 185.090 ;
        RECT 29.045 184.710 29.375 184.725 ;
        RECT 33.185 184.710 33.515 184.725 ;
        RECT 105.865 184.710 106.195 184.725 ;
        RECT 109.085 184.710 109.415 184.725 ;
        RECT 29.045 184.410 109.415 184.710 ;
        RECT 29.045 184.395 29.375 184.410 ;
        RECT 33.185 184.395 33.515 184.410 ;
        RECT 105.865 184.395 106.195 184.410 ;
        RECT 109.085 184.395 109.415 184.410 ;
        RECT 38.910 184.030 39.290 184.040 ;
        RECT 39.625 184.030 39.955 184.045 ;
        RECT 38.910 183.730 39.955 184.030 ;
        RECT 38.910 183.720 39.290 183.730 ;
        RECT 39.625 183.715 39.955 183.730 ;
        RECT 41.005 184.030 41.335 184.045 ;
        RECT 42.385 184.030 42.715 184.045 ;
        RECT 46.065 184.030 46.395 184.045 ;
        RECT 41.005 183.730 46.395 184.030 ;
        RECT 41.005 183.715 41.335 183.730 ;
        RECT 42.385 183.715 42.715 183.730 ;
        RECT 46.065 183.715 46.395 183.730 ;
        RECT 48.365 184.030 48.695 184.045 ;
        RECT 57.310 184.030 57.690 184.040 ;
        RECT 48.365 183.730 57.690 184.030 ;
        RECT 48.365 183.715 48.695 183.730 ;
        RECT 57.310 183.720 57.690 183.730 ;
        RECT 59.865 184.030 60.195 184.045 ;
        RECT 81.485 184.030 81.815 184.045 ;
        RECT 59.865 183.730 81.815 184.030 ;
        RECT 23.985 183.350 24.315 183.365 ;
        RECT 49.745 183.350 50.075 183.365 ;
        RECT 56.185 183.350 56.515 183.365 ;
        RECT 23.985 183.050 56.515 183.350 ;
        RECT 57.350 183.350 57.650 183.720 ;
        RECT 59.865 183.715 60.195 183.730 ;
        RECT 81.485 183.715 81.815 183.730 ;
        RECT 84.245 184.030 84.575 184.045 ;
        RECT 87.005 184.030 87.335 184.045 ;
        RECT 84.245 183.730 87.335 184.030 ;
        RECT 84.245 183.715 84.575 183.730 ;
        RECT 87.005 183.715 87.335 183.730 ;
        RECT 67.685 183.350 68.015 183.365 ;
        RECT 78.265 183.350 78.595 183.365 ;
        RECT 57.350 183.050 78.595 183.350 ;
        RECT 23.985 183.035 24.315 183.050 ;
        RECT 49.745 183.035 50.075 183.050 ;
        RECT 56.185 183.035 56.515 183.050 ;
        RECT 67.685 183.035 68.015 183.050 ;
        RECT 78.265 183.035 78.595 183.050 ;
        RECT 8.720 182.670 9.220 182.820 ;
        RECT 109.850 182.695 111.430 183.025 ;
        RECT 10.185 182.670 10.515 182.685 ;
        RECT 46.525 182.670 46.855 182.685 ;
        RECT 8.720 182.370 10.515 182.670 ;
        RECT 8.720 182.220 9.220 182.370 ;
        RECT 10.185 182.355 10.515 182.370 ;
        RECT 21.930 182.370 46.855 182.670 ;
        RECT 17.545 181.990 17.875 182.005 ;
        RECT 21.930 181.990 22.230 182.370 ;
        RECT 46.525 182.355 46.855 182.370 ;
        RECT 47.190 182.670 47.570 182.680 ;
        RECT 47.905 182.670 48.235 182.685 ;
        RECT 47.190 182.370 48.235 182.670 ;
        RECT 47.190 182.360 47.570 182.370 ;
        RECT 47.905 182.355 48.235 182.370 ;
        RECT 49.285 182.670 49.615 182.685 ;
        RECT 63.750 182.670 64.130 182.680 ;
        RECT 49.285 182.370 64.130 182.670 ;
        RECT 49.285 182.355 49.615 182.370 ;
        RECT 63.750 182.360 64.130 182.370 ;
        RECT 17.545 181.690 22.230 181.990 ;
        RECT 25.825 181.990 26.155 182.005 ;
        RECT 49.285 181.990 49.615 182.005 ;
        RECT 25.825 181.690 49.615 181.990 ;
        RECT 17.545 181.675 17.875 181.690 ;
        RECT 25.825 181.675 26.155 181.690 ;
        RECT 49.285 181.675 49.615 181.690 ;
        RECT 56.185 181.990 56.515 182.005 ;
        RECT 58.230 181.990 58.610 182.000 ;
        RECT 56.185 181.690 58.610 181.990 ;
        RECT 56.185 181.675 56.515 181.690 ;
        RECT 58.230 181.680 58.610 181.690 ;
        RECT 22.605 181.310 22.935 181.325 ;
        RECT 33.645 181.310 33.975 181.325 ;
        RECT 22.605 181.010 33.975 181.310 ;
        RECT 22.605 180.995 22.935 181.010 ;
        RECT 33.645 180.995 33.975 181.010 ;
        RECT 39.625 181.310 39.955 181.325 ;
        RECT 61.245 181.310 61.575 181.325 ;
        RECT 39.625 181.010 61.575 181.310 ;
        RECT 39.625 180.995 39.955 181.010 ;
        RECT 61.245 180.995 61.575 181.010 ;
        RECT 27.665 180.630 27.995 180.645 ;
        RECT 60.990 180.630 61.370 180.640 ;
        RECT 27.665 180.330 61.370 180.630 ;
        RECT 27.665 180.315 27.995 180.330 ;
        RECT 60.990 180.320 61.370 180.330 ;
        RECT 106.550 179.975 108.130 180.305 ;
        RECT 37.785 179.950 38.115 179.965 ;
        RECT 41.005 179.950 41.335 179.965 ;
        RECT 52.505 179.950 52.835 179.965 ;
        RECT 54.345 179.950 54.675 179.965 ;
        RECT 37.785 179.650 54.675 179.950 ;
        RECT 37.785 179.635 38.115 179.650 ;
        RECT 41.005 179.635 41.335 179.650 ;
        RECT 52.505 179.635 52.835 179.650 ;
        RECT 54.345 179.635 54.675 179.650 ;
        RECT 8.720 179.270 9.220 179.420 ;
        RECT 21.685 179.270 22.015 179.285 ;
        RECT 48.825 179.280 49.155 179.285 ;
        RECT 47.190 179.270 47.570 179.280 ;
        RECT 8.720 178.970 15.330 179.270 ;
        RECT 8.720 178.820 9.220 178.970 ;
        RECT 15.030 177.230 15.330 178.970 ;
        RECT 21.685 178.970 47.570 179.270 ;
        RECT 21.685 178.955 22.015 178.970 ;
        RECT 47.190 178.960 47.570 178.970 ;
        RECT 48.825 179.270 49.410 179.280 ;
        RECT 50.205 179.270 50.535 179.285 ;
        RECT 71.825 179.270 72.155 179.285 ;
        RECT 79.185 179.270 79.515 179.285 ;
        RECT 48.825 178.970 49.610 179.270 ;
        RECT 50.205 178.970 79.515 179.270 ;
        RECT 48.825 178.960 49.410 178.970 ;
        RECT 48.825 178.955 49.155 178.960 ;
        RECT 50.205 178.955 50.535 178.970 ;
        RECT 71.825 178.955 72.155 178.970 ;
        RECT 79.185 178.955 79.515 178.970 ;
        RECT 102.185 179.270 102.515 179.285 ;
        RECT 115.525 179.270 115.855 179.285 ;
        RECT 102.185 178.970 115.855 179.270 ;
        RECT 102.185 178.955 102.515 178.970 ;
        RECT 115.525 178.955 115.855 178.970 ;
        RECT 37.325 178.590 37.655 178.605 ;
        RECT 81.945 178.590 82.275 178.605 ;
        RECT 37.325 178.290 82.275 178.590 ;
        RECT 37.325 178.275 37.655 178.290 ;
        RECT 81.945 178.275 82.275 178.290 ;
        RECT 16.625 177.910 16.955 177.925 ;
        RECT 43.765 177.910 44.095 177.925 ;
        RECT 45.605 177.920 45.935 177.925 ;
        RECT 16.625 177.610 44.095 177.910 ;
        RECT 16.625 177.595 16.955 177.610 ;
        RECT 43.765 177.595 44.095 177.610 ;
        RECT 45.350 177.910 45.935 177.920 ;
        RECT 53.425 177.910 53.755 177.925 ;
        RECT 57.105 177.910 57.435 177.925 ;
        RECT 86.085 177.910 86.415 177.925 ;
        RECT 45.350 177.610 46.160 177.910 ;
        RECT 53.425 177.610 86.415 177.910 ;
        RECT 45.350 177.600 45.935 177.610 ;
        RECT 45.605 177.595 45.935 177.600 ;
        RECT 53.425 177.595 53.755 177.610 ;
        RECT 57.105 177.595 57.435 177.610 ;
        RECT 86.085 177.595 86.415 177.610 ;
        RECT 109.850 177.255 111.430 177.585 ;
        RECT 46.065 177.230 46.395 177.245 ;
        RECT 15.030 176.930 46.395 177.230 ;
        RECT 46.065 176.915 46.395 176.930 ;
        RECT 46.985 176.915 47.315 177.245 ;
        RECT 49.030 177.230 49.410 177.240 ;
        RECT 63.545 177.230 63.875 177.245 ;
        RECT 49.030 176.930 63.875 177.230 ;
        RECT 49.030 176.920 49.410 176.930 ;
        RECT 63.545 176.915 63.875 176.930 ;
        RECT 41.465 176.550 41.795 176.565 ;
        RECT 45.350 176.550 45.730 176.560 ;
        RECT 47.000 176.550 47.300 176.915 ;
        RECT 41.465 176.250 45.730 176.550 ;
        RECT 41.465 176.235 41.795 176.250 ;
        RECT 45.350 176.240 45.730 176.250 ;
        RECT 46.310 176.250 47.300 176.550 ;
        RECT 47.905 176.550 48.235 176.565 ;
        RECT 53.425 176.550 53.755 176.565 ;
        RECT 47.905 176.250 53.755 176.550 ;
        RECT 8.720 175.870 9.220 176.020 ;
        RECT 43.765 175.870 44.095 175.885 ;
        RECT 46.310 175.870 46.610 176.250 ;
        RECT 47.905 176.235 48.235 176.250 ;
        RECT 53.425 176.235 53.755 176.250 ;
        RECT 62.165 176.550 62.495 176.565 ;
        RECT 71.825 176.550 72.155 176.565 ;
        RECT 62.165 176.250 72.155 176.550 ;
        RECT 62.165 176.235 62.495 176.250 ;
        RECT 71.825 176.235 72.155 176.250 ;
        RECT 8.720 175.570 42.930 175.870 ;
        RECT 8.720 175.420 9.220 175.570 ;
        RECT 18.005 175.190 18.335 175.205 ;
        RECT 22.350 175.190 22.730 175.200 ;
        RECT 18.005 174.890 22.730 175.190 ;
        RECT 18.005 174.875 18.335 174.890 ;
        RECT 22.350 174.880 22.730 174.890 ;
        RECT 39.830 175.190 40.210 175.200 ;
        RECT 41.465 175.190 41.795 175.205 ;
        RECT 39.830 174.890 41.795 175.190 ;
        RECT 42.630 175.190 42.930 175.570 ;
        RECT 43.765 175.570 46.610 175.870 ;
        RECT 46.985 175.870 47.315 175.885 ;
        RECT 85.830 175.870 86.210 175.880 ;
        RECT 46.985 175.570 86.210 175.870 ;
        RECT 43.765 175.555 44.095 175.570 ;
        RECT 46.985 175.555 47.315 175.570 ;
        RECT 85.830 175.560 86.210 175.570 ;
        RECT 130.245 175.870 130.575 175.885 ;
        RECT 131.980 175.870 132.480 176.020 ;
        RECT 130.245 175.570 132.480 175.870 ;
        RECT 130.245 175.555 130.575 175.570 ;
        RECT 131.980 175.420 132.480 175.570 ;
        RECT 68.605 175.190 68.935 175.205 ;
        RECT 42.630 174.890 68.935 175.190 ;
        RECT 39.830 174.880 40.210 174.890 ;
        RECT 41.465 174.875 41.795 174.890 ;
        RECT 68.605 174.875 68.935 174.890 ;
        RECT 106.550 174.535 108.130 174.865 ;
        RECT 36.405 174.510 36.735 174.525 ;
        RECT 51.585 174.510 51.915 174.525 ;
        RECT 36.405 174.210 51.915 174.510 ;
        RECT 36.405 174.195 36.735 174.210 ;
        RECT 51.585 174.195 51.915 174.210 ;
        RECT 61.245 174.510 61.575 174.525 ;
        RECT 83.325 174.510 83.655 174.525 ;
        RECT 61.245 174.210 83.655 174.510 ;
        RECT 61.245 174.195 61.575 174.210 ;
        RECT 83.325 174.195 83.655 174.210 ;
        RECT 30.425 173.830 30.755 173.845 ;
        RECT 78.725 173.830 79.055 173.845 ;
        RECT 30.425 173.530 79.055 173.830 ;
        RECT 30.425 173.515 30.755 173.530 ;
        RECT 78.725 173.515 79.055 173.530 ;
        RECT 37.990 173.150 38.370 173.160 ;
        RECT 42.385 173.150 42.715 173.165 ;
        RECT 37.990 172.850 42.715 173.150 ;
        RECT 37.990 172.840 38.370 172.850 ;
        RECT 42.385 172.835 42.715 172.850 ;
        RECT 8.720 172.470 9.220 172.620 ;
        RECT 33.185 172.470 33.515 172.485 ;
        RECT 8.720 172.170 33.515 172.470 ;
        RECT 8.720 172.020 9.220 172.170 ;
        RECT 33.185 172.155 33.515 172.170 ;
        RECT 130.245 172.470 130.575 172.485 ;
        RECT 131.980 172.470 132.480 172.620 ;
        RECT 130.245 172.170 132.480 172.470 ;
        RECT 130.245 172.155 130.575 172.170 ;
        RECT 109.850 171.815 111.430 172.145 ;
        RECT 131.980 172.020 132.480 172.170 ;
        RECT 23.065 171.790 23.395 171.805 ;
        RECT 48.365 171.790 48.695 171.805 ;
        RECT 23.065 171.490 48.695 171.790 ;
        RECT 23.065 171.475 23.395 171.490 ;
        RECT 48.365 171.475 48.695 171.490 ;
        RECT 26.285 171.110 26.615 171.125 ;
        RECT 45.145 171.110 45.475 171.125 ;
        RECT 26.285 170.810 45.475 171.110 ;
        RECT 26.285 170.795 26.615 170.810 ;
        RECT 45.145 170.795 45.475 170.810 ;
        RECT 20.305 170.430 20.635 170.445 ;
        RECT 52.965 170.430 53.295 170.445 ;
        RECT 20.305 170.130 53.295 170.430 ;
        RECT 20.305 170.115 20.635 170.130 ;
        RECT 52.965 170.115 53.295 170.130 ;
        RECT 19.845 169.750 20.175 169.765 ;
        RECT 48.825 169.750 49.155 169.765 ;
        RECT 19.845 169.450 49.155 169.750 ;
        RECT 19.845 169.435 20.175 169.450 ;
        RECT 48.825 169.435 49.155 169.450 ;
        RECT 8.720 169.070 9.220 169.220 ;
        RECT 106.550 169.095 108.130 169.425 ;
        RECT 44.685 169.070 45.015 169.085 ;
        RECT 8.720 168.770 45.015 169.070 ;
        RECT 8.720 168.620 9.220 168.770 ;
        RECT 44.685 168.755 45.015 168.770 ;
        RECT 125.645 169.070 125.975 169.085 ;
        RECT 131.980 169.070 132.480 169.220 ;
        RECT 125.645 168.770 132.480 169.070 ;
        RECT 125.645 168.755 125.975 168.770 ;
        RECT 131.980 168.620 132.480 168.770 ;
        RECT 25.825 168.390 26.155 168.405 ;
        RECT 51.585 168.390 51.915 168.405 ;
        RECT 25.825 168.090 51.915 168.390 ;
        RECT 25.825 168.075 26.155 168.090 ;
        RECT 51.585 168.075 51.915 168.090 ;
        RECT 8.720 165.670 9.220 165.820 ;
        RECT 38.705 165.670 39.035 165.685 ;
        RECT 8.720 165.370 39.035 165.670 ;
        RECT 8.720 165.220 9.220 165.370 ;
        RECT 38.705 165.355 39.035 165.370 ;
        RECT 28.125 164.310 28.455 164.325 ;
        RECT 41.925 164.310 42.255 164.325 ;
        RECT 28.125 164.010 42.255 164.310 ;
        RECT 28.125 163.995 28.455 164.010 ;
        RECT 41.925 163.995 42.255 164.010 ;
        RECT 26.745 163.630 27.075 163.645 ;
        RECT 38.705 163.630 39.035 163.645 ;
        RECT 26.745 163.330 39.035 163.630 ;
        RECT 26.745 163.315 27.075 163.330 ;
        RECT 38.705 163.315 39.035 163.330 ;
        RECT 8.720 162.270 9.220 162.420 ;
        RECT 43.765 162.270 44.095 162.285 ;
        RECT 8.720 161.970 44.095 162.270 ;
        RECT 8.720 161.820 9.220 161.970 ;
        RECT 43.765 161.955 44.095 161.970 ;
        RECT 8.720 158.870 9.220 159.020 ;
        RECT 11.105 158.870 11.435 158.885 ;
        RECT 8.720 158.570 11.435 158.870 ;
        RECT 8.720 158.420 9.220 158.570 ;
        RECT 11.105 158.555 11.435 158.570 ;
        RECT 79.480 50.170 80.050 50.690 ;
        RECT 68.665 49.870 69.975 49.875 ;
        RECT 68.635 48.950 70.005 49.870 ;
        RECT 68.665 48.945 69.975 48.950 ;
        RECT 146.510 48.490 146.965 48.515 ;
        RECT 94.645 48.085 146.965 48.490 ;
        RECT 94.645 46.215 95.050 48.085 ;
        RECT 146.510 48.060 146.965 48.085 ;
        RECT 143.585 46.565 144.065 46.590 ;
        RECT 95.565 46.470 107.495 46.565 ;
        RECT 109.175 46.470 144.065 46.565 ;
        RECT 95.565 46.135 144.065 46.470 ;
        RECT 79.805 34.570 81.180 36.025 ;
        RECT 68.665 34.225 69.975 34.230 ;
        RECT 68.635 33.330 70.005 34.225 ;
        RECT 68.665 33.325 69.975 33.330 ;
        RECT 95.565 32.295 95.995 46.135 ;
        RECT 143.585 46.110 144.065 46.135 ;
        RECT 150.825 45.680 151.375 45.705 ;
        RECT 94.695 31.865 95.995 32.295 ;
        RECT 96.770 45.180 151.375 45.680 ;
        RECT 80.460 18.535 81.835 19.990 ;
        RECT 68.660 16.800 69.980 18.180 ;
        RECT 96.770 16.190 97.270 45.180 ;
        RECT 150.825 45.155 151.375 45.180 ;
        RECT 148.960 44.095 149.510 44.120 ;
        RECT 122.495 43.595 149.510 44.095 ;
        RECT 148.960 43.570 149.510 43.595 ;
        RECT 141.500 27.655 141.990 27.680 ;
        RECT 122.590 27.215 141.990 27.655 ;
        RECT 141.500 27.190 141.990 27.215 ;
        RECT 94.530 15.690 97.270 16.190 ;
        RECT 142.355 13.980 142.905 14.005 ;
        RECT 122.560 13.480 142.905 13.980 ;
        RECT 142.355 13.455 142.905 13.480 ;
        RECT 7.350 7.445 7.730 7.470 ;
        RECT 7.350 7.115 142.905 7.445 ;
        RECT 7.350 7.090 7.730 7.115 ;
        RECT 80.415 2.885 81.790 4.340 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 22.375 210.915 22.705 211.245 ;
        RECT 22.390 175.205 22.690 210.915 ;
        RECT 56.415 210.235 56.745 210.565 ;
        RECT 38.935 208.875 39.265 209.205 ;
        RECT 38.015 193.235 38.345 193.565 ;
        RECT 22.375 174.875 22.705 175.205 ;
        RECT 38.030 173.165 38.330 193.235 ;
        RECT 38.950 184.045 39.250 208.875 ;
        RECT 54.575 205.475 54.905 205.805 ;
        RECT 52.735 202.075 53.065 202.405 ;
        RECT 53.655 202.075 53.985 202.405 ;
        RECT 42.615 197.315 42.945 197.645 ;
        RECT 39.855 195.275 40.185 195.605 ;
        RECT 38.935 183.715 39.265 184.045 ;
        RECT 39.870 175.205 40.170 195.275 ;
        RECT 42.630 194.245 42.930 197.315 ;
        RECT 42.615 193.915 42.945 194.245 ;
        RECT 49.055 193.235 49.385 193.565 ;
        RECT 49.070 189.485 49.370 193.235 ;
        RECT 49.055 189.155 49.385 189.485 ;
        RECT 52.750 185.405 53.050 202.075 ;
        RECT 53.670 192.205 53.970 202.075 ;
        RECT 53.655 191.875 53.985 192.205 ;
        RECT 54.590 188.805 54.890 205.475 ;
        RECT 56.430 195.605 56.730 210.235 ;
        RECT 61.015 200.715 61.345 201.045 ;
        RECT 58.255 197.995 58.585 198.325 ;
        RECT 56.415 195.275 56.745 195.605 ;
        RECT 57.335 191.875 57.665 192.205 ;
        RECT 54.575 188.475 54.905 188.805 ;
        RECT 52.735 185.075 53.065 185.405 ;
        RECT 57.350 184.045 57.650 191.875 ;
        RECT 57.335 183.715 57.665 184.045 ;
        RECT 47.215 182.355 47.545 182.685 ;
        RECT 47.230 179.285 47.530 182.355 ;
        RECT 58.270 182.005 58.570 197.995 ;
        RECT 58.255 181.675 58.585 182.005 ;
        RECT 61.030 180.645 61.330 200.715 ;
        RECT 85.855 200.035 86.185 200.365 ;
        RECT 61.935 195.275 62.265 195.605 ;
        RECT 61.950 190.165 62.250 195.275 ;
        RECT 63.775 193.915 64.105 194.245 ;
        RECT 61.935 189.835 62.265 190.165 ;
        RECT 63.790 182.685 64.090 193.915 ;
        RECT 63.775 182.355 64.105 182.685 ;
        RECT 61.015 180.315 61.345 180.645 ;
        RECT 47.215 178.955 47.545 179.285 ;
        RECT 49.055 178.955 49.385 179.285 ;
        RECT 45.375 177.595 45.705 177.925 ;
        RECT 45.390 176.565 45.690 177.595 ;
        RECT 49.070 177.245 49.370 178.955 ;
        RECT 49.055 176.915 49.385 177.245 ;
        RECT 45.375 176.235 45.705 176.565 ;
        RECT 85.870 175.885 86.170 200.035 ;
        RECT 85.855 175.555 86.185 175.885 ;
        RECT 39.855 174.875 40.185 175.205 ;
        RECT 38.015 172.835 38.345 173.165 ;
        RECT 106.540 169.020 108.140 213.020 ;
        RECT 109.840 169.020 111.440 213.020 ;
        RECT 80.525 50.625 81.705 50.740 ;
        RECT 79.535 50.230 81.705 50.625 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 68.660 18.155 69.980 49.875 ;
        RECT 80.525 35.855 81.705 50.230 ;
        RECT 79.870 34.675 81.705 35.855 ;
        RECT 68.655 16.825 69.985 18.155 ;
        RECT 80.525 4.270 81.705 34.675 ;
        RECT 80.495 3.030 81.735 4.270 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

