VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 1.290 52.730 13.780 58.190 ;
        RECT 1.290 50.380 31.720 52.730 ;
        RECT 43.310 50.380 61.780 52.730 ;
        RECT 67.310 50.380 85.780 52.730 ;
      LAYER nwell ;
        RECT 27.290 49.600 29.790 49.880 ;
        RECT 55.790 49.600 58.290 49.880 ;
        RECT 83.290 49.600 85.790 49.880 ;
        RECT 111.790 49.600 114.290 49.880 ;
        RECT 5.410 49.355 12.800 49.585 ;
        RECT 1.290 47.890 12.800 49.355 ;
        RECT 26.050 49.355 29.790 49.600 ;
        RECT 33.410 49.355 40.800 49.585 ;
        RECT 26.050 47.890 40.800 49.355 ;
        RECT 54.050 49.355 58.290 49.600 ;
        RECT 61.410 49.355 68.800 49.585 ;
        RECT 54.050 47.890 68.800 49.355 ;
        RECT 82.050 49.355 85.790 49.600 ;
        RECT 89.410 49.355 96.800 49.585 ;
        RECT 82.050 47.890 96.800 49.355 ;
        RECT 110.050 49.355 114.290 49.600 ;
        RECT 117.410 49.355 124.800 49.585 ;
        RECT 110.050 47.890 124.800 49.355 ;
        RECT 1.290 45.580 21.135 47.890 ;
        RECT 26.050 45.595 49.135 47.890 ;
        RECT 54.050 45.595 77.135 47.890 ;
        RECT 82.050 45.595 105.135 47.890 ;
        RECT 110.050 45.595 133.135 47.890 ;
        RECT 138.050 45.595 140.160 49.600 ;
        RECT 24.025 45.580 49.135 45.595 ;
        RECT 52.025 45.580 77.135 45.595 ;
        RECT 80.025 45.580 105.135 45.595 ;
        RECT 108.025 45.580 133.135 45.595 ;
        RECT 136.025 45.580 140.160 45.595 ;
        RECT 1.290 39.410 140.160 45.580 ;
      LAYER pwell ;
        RECT 143.290 44.730 149.800 50.190 ;
        RECT 143.290 40.560 155.780 44.730 ;
      LAYER nwell ;
        RECT 1.290 39.405 26.135 39.410 ;
        RECT 27.440 39.405 54.135 39.410 ;
        RECT 55.790 39.405 82.135 39.410 ;
        RECT 84.280 39.405 110.135 39.410 ;
        RECT 111.790 39.405 138.135 39.410 ;
        RECT 1.290 39.395 24.110 39.405 ;
        RECT 12.720 39.390 24.110 39.395 ;
        RECT 27.545 39.395 52.110 39.405 ;
        RECT 27.545 39.390 29.790 39.395 ;
        RECT 40.720 39.390 52.110 39.395 ;
        RECT 55.790 39.395 80.110 39.405 ;
        RECT 55.790 39.380 58.290 39.395 ;
        RECT 68.720 39.390 80.110 39.395 ;
        RECT 84.850 39.395 108.110 39.405 ;
        RECT 84.850 39.380 85.790 39.395 ;
        RECT 96.720 39.390 108.110 39.395 ;
        RECT 111.790 39.395 136.110 39.405 ;
        RECT 111.790 39.380 114.290 39.395 ;
        RECT 124.720 39.390 136.110 39.395 ;
      LAYER pwell ;
        RECT 26.135 39.020 28.245 39.025 ;
        RECT 54.135 39.020 56.245 39.025 ;
        RECT 82.135 39.020 84.245 39.025 ;
        RECT 110.135 39.020 112.245 39.025 ;
        RECT 138.135 39.020 140.245 39.025 ;
        RECT 24.110 39.015 28.245 39.020 ;
        RECT 52.110 39.015 56.245 39.020 ;
        RECT 80.110 39.015 84.245 39.020 ;
        RECT 108.110 39.015 112.245 39.020 ;
        RECT 136.110 39.015 140.245 39.020 ;
        RECT 1.950 35.920 28.245 39.015 ;
        RECT 1.950 34.915 24.200 35.920 ;
        RECT 26.135 34.925 28.245 35.920 ;
        RECT 29.950 35.920 56.245 39.015 ;
        RECT 29.950 34.915 52.200 35.920 ;
        RECT 54.135 34.925 56.245 35.920 ;
        RECT 57.950 35.920 84.245 39.015 ;
        RECT 57.950 34.915 80.200 35.920 ;
        RECT 82.135 34.925 84.245 35.920 ;
        RECT 85.950 35.920 112.245 39.015 ;
        RECT 85.950 34.915 108.200 35.920 ;
        RECT 110.135 34.925 112.245 35.920 ;
        RECT 113.950 35.920 140.245 39.015 ;
        RECT 113.950 34.915 136.200 35.920 ;
        RECT 138.135 34.925 140.245 35.920 ;
      LAYER nwell ;
        RECT 27.290 33.600 29.790 33.880 ;
        RECT 55.290 33.600 57.790 33.880 ;
        RECT 83.790 33.600 86.290 33.880 ;
        RECT 111.790 33.600 114.290 33.880 ;
        RECT 5.410 33.355 12.800 33.585 ;
        RECT 1.290 31.890 12.800 33.355 ;
        RECT 26.050 33.355 29.790 33.600 ;
        RECT 33.410 33.355 40.800 33.585 ;
        RECT 26.050 31.890 40.800 33.355 ;
        RECT 54.050 33.355 57.790 33.600 ;
        RECT 61.410 33.355 68.800 33.585 ;
        RECT 54.050 31.890 68.800 33.355 ;
        RECT 82.050 33.355 86.290 33.600 ;
        RECT 89.410 33.355 96.800 33.585 ;
        RECT 82.050 31.890 96.800 33.355 ;
        RECT 110.050 33.355 114.290 33.600 ;
        RECT 117.410 33.355 124.800 33.585 ;
        RECT 110.050 31.890 124.800 33.355 ;
        RECT 1.290 29.580 21.135 31.890 ;
        RECT 26.050 29.595 49.135 31.890 ;
        RECT 54.050 29.595 77.135 31.890 ;
        RECT 82.050 29.595 105.135 31.890 ;
        RECT 110.050 29.595 133.135 31.890 ;
        RECT 138.050 29.595 140.160 33.600 ;
        RECT 24.025 29.580 49.135 29.595 ;
        RECT 52.025 29.580 77.135 29.595 ;
        RECT 80.025 29.580 105.135 29.595 ;
        RECT 108.025 29.580 133.135 29.595 ;
        RECT 136.025 29.580 140.160 29.595 ;
        RECT 1.290 23.410 140.160 29.580 ;
        RECT 1.290 23.405 26.135 23.410 ;
        RECT 28.755 23.405 54.135 23.410 ;
        RECT 56.840 23.405 82.135 23.410 ;
        RECT 83.790 23.405 110.135 23.410 ;
        RECT 111.790 23.405 138.135 23.410 ;
        RECT 1.290 23.395 24.110 23.405 ;
        RECT 12.720 23.390 24.110 23.395 ;
        RECT 28.755 23.395 52.110 23.405 ;
        RECT 28.755 23.380 29.790 23.395 ;
        RECT 40.720 23.390 52.110 23.395 ;
        RECT 56.840 23.395 80.110 23.405 ;
        RECT 56.840 23.380 57.790 23.395 ;
        RECT 68.720 23.390 80.110 23.395 ;
        RECT 83.790 23.395 108.110 23.405 ;
        RECT 83.790 23.380 86.290 23.395 ;
        RECT 96.720 23.390 108.110 23.395 ;
        RECT 111.790 23.395 136.110 23.405 ;
        RECT 111.790 23.380 114.290 23.395 ;
        RECT 124.720 23.390 136.110 23.395 ;
      LAYER pwell ;
        RECT 26.135 23.020 28.245 23.025 ;
        RECT 54.135 23.020 56.245 23.025 ;
        RECT 82.135 23.020 84.245 23.025 ;
        RECT 110.135 23.020 112.245 23.025 ;
        RECT 138.135 23.020 140.245 23.025 ;
        RECT 24.110 23.015 28.245 23.020 ;
        RECT 52.110 23.015 56.245 23.020 ;
        RECT 80.110 23.015 84.245 23.020 ;
        RECT 108.110 23.015 112.245 23.020 ;
        RECT 136.110 23.015 140.245 23.020 ;
        RECT 1.950 19.920 28.245 23.015 ;
        RECT 1.950 18.915 24.200 19.920 ;
        RECT 26.135 18.925 28.245 19.920 ;
        RECT 29.950 19.920 56.245 23.015 ;
        RECT 29.950 18.915 52.200 19.920 ;
        RECT 54.135 18.925 56.245 19.920 ;
        RECT 57.950 19.920 84.245 23.015 ;
        RECT 57.950 18.915 80.200 19.920 ;
        RECT 82.135 18.925 84.245 19.920 ;
        RECT 85.950 19.920 112.245 23.015 ;
        RECT 85.950 18.915 108.200 19.920 ;
        RECT 110.135 18.925 112.245 19.920 ;
        RECT 113.950 19.920 140.245 23.015 ;
        RECT 113.950 18.915 136.200 19.920 ;
        RECT 138.135 18.925 140.245 19.920 ;
      LAYER nwell ;
        RECT 27.790 17.600 30.290 17.880 ;
        RECT 55.290 17.600 57.790 17.880 ;
        RECT 83.790 17.600 86.290 17.880 ;
        RECT 111.790 17.600 114.290 17.880 ;
        RECT 5.410 17.355 12.800 17.585 ;
        RECT 1.290 15.890 12.800 17.355 ;
        RECT 26.050 17.355 30.290 17.600 ;
        RECT 33.410 17.355 40.800 17.585 ;
        RECT 26.050 15.890 40.800 17.355 ;
        RECT 54.050 17.355 57.790 17.600 ;
        RECT 61.410 17.355 68.800 17.585 ;
        RECT 54.050 15.890 68.800 17.355 ;
        RECT 82.050 17.355 86.290 17.600 ;
        RECT 89.410 17.355 96.800 17.585 ;
        RECT 82.050 15.890 96.800 17.355 ;
        RECT 110.050 17.355 114.290 17.600 ;
        RECT 117.410 17.355 124.800 17.585 ;
        RECT 110.050 15.890 124.800 17.355 ;
        RECT 1.290 13.580 21.135 15.890 ;
        RECT 26.050 13.595 49.135 15.890 ;
        RECT 54.050 13.595 77.135 15.890 ;
        RECT 82.050 13.595 105.135 15.890 ;
        RECT 110.050 13.595 133.135 15.890 ;
        RECT 138.050 13.595 140.160 17.600 ;
        RECT 24.025 13.580 49.135 13.595 ;
        RECT 52.025 13.580 77.135 13.595 ;
        RECT 80.025 13.580 105.135 13.595 ;
        RECT 108.025 13.580 133.135 13.595 ;
        RECT 136.025 13.580 140.160 13.595 ;
        RECT 1.290 7.410 140.160 13.580 ;
        RECT 1.290 7.405 26.135 7.410 ;
        RECT 27.790 7.405 54.135 7.410 ;
        RECT 55.495 7.405 82.135 7.410 ;
        RECT 83.790 7.405 110.135 7.410 ;
        RECT 111.790 7.405 138.135 7.410 ;
        RECT 1.290 7.395 24.110 7.405 ;
        RECT 12.720 7.390 24.110 7.395 ;
        RECT 27.790 7.395 52.110 7.405 ;
        RECT 57.115 7.400 80.110 7.405 ;
        RECT 57.290 7.395 80.110 7.400 ;
        RECT 27.790 7.380 30.290 7.395 ;
        RECT 40.720 7.390 52.110 7.395 ;
        RECT 68.720 7.390 80.110 7.395 ;
        RECT 83.790 7.395 108.110 7.405 ;
        RECT 83.790 7.380 86.290 7.395 ;
        RECT 96.720 7.390 108.110 7.395 ;
        RECT 111.790 7.395 136.110 7.405 ;
        RECT 111.790 7.380 114.290 7.395 ;
        RECT 124.720 7.390 136.110 7.395 ;
      LAYER pwell ;
        RECT 26.135 7.020 28.245 7.025 ;
        RECT 54.135 7.020 56.245 7.025 ;
        RECT 82.135 7.020 84.245 7.025 ;
        RECT 110.135 7.020 112.245 7.025 ;
        RECT 138.135 7.020 140.245 7.025 ;
        RECT 24.110 7.015 28.245 7.020 ;
        RECT 52.110 7.015 56.245 7.020 ;
        RECT 80.110 7.015 84.245 7.020 ;
        RECT 108.110 7.015 112.245 7.020 ;
        RECT 136.110 7.015 140.245 7.020 ;
        RECT 1.950 3.920 28.245 7.015 ;
        RECT 1.950 2.915 24.200 3.920 ;
        RECT 26.135 2.925 28.245 3.920 ;
        RECT 29.950 3.920 56.245 7.015 ;
        RECT 29.950 2.915 52.200 3.920 ;
        RECT 54.135 2.925 56.245 3.920 ;
        RECT 57.950 3.920 84.245 7.015 ;
        RECT 57.950 2.915 80.200 3.920 ;
        RECT 82.135 2.925 84.245 3.920 ;
        RECT 85.950 3.920 112.245 7.015 ;
        RECT 85.950 2.915 108.200 3.920 ;
        RECT 110.135 2.925 112.245 3.920 ;
        RECT 113.950 3.920 140.245 7.015 ;
        RECT 113.950 2.915 136.200 3.920 ;
        RECT 138.135 2.925 140.245 3.920 ;
      LAYER li1 ;
        RECT 1.470 57.840 13.600 58.010 ;
        RECT 1.470 56.190 1.640 57.840 ;
        RECT 2.120 56.670 4.280 57.360 ;
        RECT 4.810 56.670 6.970 57.360 ;
        RECT 7.450 56.190 7.620 57.840 ;
        RECT 8.100 56.670 10.260 57.360 ;
        RECT 10.790 56.670 12.950 57.360 ;
        RECT 13.430 56.190 13.600 57.840 ;
        RECT 1.470 56.020 13.600 56.190 ;
        RECT 1.470 54.370 1.640 56.020 ;
        RECT 2.120 54.850 4.280 55.540 ;
        RECT 4.810 54.850 6.970 55.540 ;
        RECT 7.450 54.370 7.620 56.020 ;
        RECT 8.100 54.850 10.260 55.540 ;
        RECT 10.790 54.850 12.950 55.540 ;
        RECT 13.430 54.370 13.600 56.020 ;
        RECT 1.470 54.200 13.600 54.370 ;
        RECT 1.470 52.550 1.640 54.200 ;
        RECT 2.120 53.030 4.280 53.720 ;
        RECT 4.810 53.030 6.970 53.720 ;
        RECT 7.450 52.550 7.620 54.200 ;
        RECT 8.100 53.030 10.260 53.720 ;
        RECT 10.790 53.030 12.950 53.720 ;
        RECT 13.430 52.550 13.600 54.200 ;
        RECT 1.470 52.380 31.540 52.550 ;
        RECT 1.470 50.855 1.640 52.380 ;
        RECT 2.120 51.210 4.280 51.900 ;
        RECT 4.810 51.210 6.970 51.900 ;
        RECT 7.450 50.855 7.620 52.380 ;
        RECT 8.100 51.210 10.260 51.900 ;
        RECT 10.790 51.210 12.950 51.900 ;
        RECT 1.470 50.730 9.960 50.855 ;
        RECT 13.430 50.730 13.600 52.380 ;
        RECT 14.080 51.210 16.240 51.900 ;
        RECT 16.770 51.210 18.930 51.900 ;
        RECT 19.410 50.730 19.580 52.380 ;
        RECT 20.060 51.210 22.220 51.900 ;
        RECT 22.750 51.210 24.910 51.900 ;
        RECT 25.390 50.730 25.560 52.380 ;
        RECT 26.040 51.210 28.200 51.900 ;
        RECT 28.730 51.210 30.890 51.900 ;
        RECT 31.370 50.730 31.540 52.380 ;
        RECT 1.470 50.560 31.540 50.730 ;
        RECT 43.490 52.540 61.600 52.550 ;
        RECT 67.490 52.540 85.600 52.550 ;
        RECT 43.490 52.380 85.600 52.540 ;
        RECT 43.490 50.730 43.660 52.380 ;
        RECT 44.140 51.210 46.300 51.900 ;
        RECT 46.830 51.210 48.990 51.900 ;
        RECT 49.470 50.730 49.640 52.380 ;
        RECT 50.120 51.210 52.280 51.900 ;
        RECT 52.810 51.210 54.970 51.900 ;
        RECT 55.450 50.730 55.620 52.380 ;
        RECT 61.430 52.090 67.670 52.380 ;
        RECT 56.100 51.210 58.260 51.900 ;
        RECT 58.790 51.210 60.950 51.900 ;
        RECT 61.430 50.730 61.600 52.090 ;
        RECT 43.490 50.560 61.600 50.730 ;
        RECT 67.490 50.730 67.660 52.090 ;
        RECT 68.140 51.210 70.300 51.900 ;
        RECT 70.830 51.210 72.990 51.900 ;
        RECT 73.470 50.730 73.640 52.380 ;
        RECT 74.120 51.210 76.280 51.900 ;
        RECT 76.810 51.210 78.970 51.900 ;
        RECT 79.450 50.730 79.620 52.380 ;
        RECT 80.100 51.210 82.260 51.900 ;
        RECT 82.790 51.210 84.950 51.900 ;
        RECT 85.430 50.730 85.600 52.380 ;
        RECT 67.490 50.560 85.600 50.730 ;
        RECT 1.585 50.360 9.960 50.560 ;
        RECT 77.790 50.170 80.360 50.560 ;
        RECT 1.450 49.480 27.925 49.960 ;
        RECT 29.450 49.480 55.925 49.960 ;
        RECT 57.450 49.480 83.925 49.960 ;
        RECT 85.450 49.480 111.925 49.960 ;
        RECT 113.450 49.480 139.925 49.960 ;
        RECT 1.435 49.420 27.925 49.480 ;
        RECT 29.435 49.420 55.925 49.480 ;
        RECT 57.435 49.420 83.925 49.480 ;
        RECT 85.435 49.420 111.925 49.480 ;
        RECT 113.435 49.420 139.925 49.480 ;
        RECT 143.470 49.840 149.620 50.010 ;
        RECT 1.435 49.260 27.980 49.420 ;
        RECT 1.435 49.235 14.180 49.260 ;
        RECT 1.435 49.005 5.760 49.235 ;
        RECT 1.470 39.745 1.640 49.005 ;
        RECT 2.365 48.435 4.405 48.605 ;
        RECT 1.980 40.375 2.150 48.375 ;
        RECT 4.620 40.375 4.790 48.375 ;
        RECT 2.365 40.145 4.405 40.315 ;
        RECT 5.130 39.745 5.300 49.005 ;
        RECT 1.470 39.575 5.300 39.745 ;
        RECT 5.590 39.745 5.760 49.005 ;
        RECT 6.390 48.725 8.390 48.895 ;
        RECT 6.160 40.470 6.330 48.510 ;
        RECT 8.450 40.470 8.620 48.510 ;
        RECT 6.390 40.085 8.390 40.255 ;
        RECT 9.020 39.745 9.190 49.235 ;
        RECT 9.820 48.725 11.820 48.895 ;
        RECT 9.590 40.470 9.760 48.510 ;
        RECT 11.880 40.470 12.050 48.510 ;
        RECT 12.450 47.665 14.180 49.235 ;
        RECT 26.230 49.250 27.980 49.260 ;
        RECT 12.450 47.495 20.915 47.665 ;
        RECT 12.450 46.085 14.255 47.495 ;
        RECT 14.595 46.625 14.765 46.955 ;
        RECT 14.980 46.925 20.020 47.095 ;
        RECT 14.980 46.485 20.020 46.655 ;
        RECT 20.235 46.625 20.405 46.955 ;
        RECT 20.745 46.085 20.915 47.495 ;
        RECT 12.450 45.915 20.915 46.085 ;
        RECT 12.450 45.400 14.180 45.915 ;
        RECT 12.450 45.285 23.930 45.400 ;
        RECT 9.820 40.085 11.820 40.255 ;
        RECT 12.450 39.745 12.620 45.285 ;
        RECT 5.590 39.575 12.620 39.745 ;
        RECT 12.900 45.230 23.930 45.285 ;
        RECT 12.900 39.740 13.070 45.230 ;
        RECT 13.700 44.720 17.700 44.890 ;
        RECT 13.470 40.465 13.640 44.505 ;
        RECT 17.760 40.465 17.930 44.505 ;
        RECT 13.700 40.080 17.700 40.250 ;
        RECT 18.330 39.740 18.500 45.230 ;
        RECT 19.130 44.720 23.130 44.890 ;
        RECT 18.900 40.465 19.070 44.505 ;
        RECT 23.190 40.465 23.360 44.505 ;
        RECT 19.130 40.080 23.130 40.250 ;
        RECT 23.760 39.740 23.930 45.230 ;
        RECT 12.900 39.570 23.930 39.740 ;
        RECT 24.205 45.245 25.955 45.415 ;
        RECT 24.205 39.755 24.375 45.245 ;
        RECT 24.915 44.735 25.245 44.905 ;
        RECT 24.775 40.480 24.945 44.520 ;
        RECT 25.215 40.480 25.385 44.520 ;
        RECT 24.915 40.095 25.245 40.265 ;
        RECT 25.785 39.755 25.955 45.245 ;
        RECT 24.205 39.585 25.955 39.755 ;
        RECT 26.230 39.760 26.400 49.250 ;
        RECT 26.940 48.740 27.270 48.910 ;
        RECT 26.800 40.485 26.970 48.525 ;
        RECT 27.240 40.485 27.410 48.525 ;
        RECT 26.940 40.100 27.270 40.270 ;
        RECT 27.810 39.760 27.980 49.250 ;
        RECT 29.435 49.260 55.980 49.420 ;
        RECT 29.435 49.235 42.180 49.260 ;
        RECT 29.435 49.005 33.760 49.235 ;
        RECT 26.230 39.590 27.980 39.760 ;
        RECT 29.470 39.745 29.640 49.005 ;
        RECT 30.365 48.435 32.405 48.605 ;
        RECT 29.980 40.375 30.150 48.375 ;
        RECT 32.620 40.375 32.790 48.375 ;
        RECT 30.365 40.145 32.405 40.315 ;
        RECT 33.130 39.745 33.300 49.005 ;
        RECT 29.470 39.575 33.300 39.745 ;
        RECT 33.590 39.745 33.760 49.005 ;
        RECT 34.390 48.725 36.390 48.895 ;
        RECT 34.160 40.470 34.330 48.510 ;
        RECT 36.450 40.470 36.620 48.510 ;
        RECT 34.390 40.085 36.390 40.255 ;
        RECT 37.020 39.745 37.190 49.235 ;
        RECT 37.820 48.725 39.820 48.895 ;
        RECT 37.590 40.470 37.760 48.510 ;
        RECT 39.880 40.470 40.050 48.510 ;
        RECT 40.450 47.665 42.180 49.235 ;
        RECT 54.230 49.250 55.980 49.260 ;
        RECT 40.450 47.495 48.915 47.665 ;
        RECT 40.450 46.085 42.255 47.495 ;
        RECT 42.595 46.625 42.765 46.955 ;
        RECT 42.980 46.925 48.020 47.095 ;
        RECT 42.980 46.485 48.020 46.655 ;
        RECT 48.235 46.625 48.405 46.955 ;
        RECT 48.745 46.085 48.915 47.495 ;
        RECT 40.450 45.915 48.915 46.085 ;
        RECT 40.450 45.400 42.180 45.915 ;
        RECT 40.450 45.285 51.930 45.400 ;
        RECT 37.820 40.085 39.820 40.255 ;
        RECT 40.450 39.745 40.620 45.285 ;
        RECT 33.590 39.575 40.620 39.745 ;
        RECT 40.900 45.230 51.930 45.285 ;
        RECT 40.900 39.740 41.070 45.230 ;
        RECT 41.700 44.720 45.700 44.890 ;
        RECT 41.470 40.465 41.640 44.505 ;
        RECT 45.760 40.465 45.930 44.505 ;
        RECT 41.700 40.080 45.700 40.250 ;
        RECT 46.330 39.740 46.500 45.230 ;
        RECT 47.130 44.720 51.130 44.890 ;
        RECT 46.900 40.465 47.070 44.505 ;
        RECT 51.190 40.465 51.360 44.505 ;
        RECT 47.130 40.080 51.130 40.250 ;
        RECT 51.760 39.740 51.930 45.230 ;
        RECT 40.900 39.570 51.930 39.740 ;
        RECT 52.205 45.245 53.955 45.415 ;
        RECT 52.205 39.755 52.375 45.245 ;
        RECT 52.915 44.735 53.245 44.905 ;
        RECT 52.775 40.480 52.945 44.520 ;
        RECT 53.215 40.480 53.385 44.520 ;
        RECT 52.915 40.095 53.245 40.265 ;
        RECT 53.785 39.755 53.955 45.245 ;
        RECT 52.205 39.585 53.955 39.755 ;
        RECT 54.230 39.760 54.400 49.250 ;
        RECT 54.940 48.740 55.270 48.910 ;
        RECT 54.800 40.485 54.970 48.525 ;
        RECT 55.240 40.485 55.410 48.525 ;
        RECT 54.940 40.100 55.270 40.270 ;
        RECT 55.810 39.760 55.980 49.250 ;
        RECT 57.435 49.260 83.980 49.420 ;
        RECT 57.435 49.235 70.180 49.260 ;
        RECT 57.435 49.005 61.760 49.235 ;
        RECT 54.230 39.590 55.980 39.760 ;
        RECT 57.470 39.745 57.640 49.005 ;
        RECT 58.365 48.435 60.405 48.605 ;
        RECT 57.980 40.375 58.150 48.375 ;
        RECT 60.620 40.375 60.790 48.375 ;
        RECT 58.365 40.145 60.405 40.315 ;
        RECT 61.130 39.745 61.300 49.005 ;
        RECT 57.470 39.575 61.300 39.745 ;
        RECT 61.590 39.745 61.760 49.005 ;
        RECT 62.390 48.725 64.390 48.895 ;
        RECT 62.160 40.470 62.330 48.510 ;
        RECT 64.450 40.470 64.620 48.510 ;
        RECT 62.390 40.085 64.390 40.255 ;
        RECT 65.020 39.745 65.190 49.235 ;
        RECT 65.820 48.725 67.820 48.895 ;
        RECT 65.590 40.470 65.760 48.510 ;
        RECT 67.880 40.470 68.050 48.510 ;
        RECT 68.450 47.665 70.180 49.235 ;
        RECT 82.230 49.250 83.980 49.260 ;
        RECT 68.450 47.495 76.915 47.665 ;
        RECT 68.450 46.085 70.255 47.495 ;
        RECT 70.595 46.625 70.765 46.955 ;
        RECT 70.980 46.925 76.020 47.095 ;
        RECT 70.980 46.485 76.020 46.655 ;
        RECT 76.235 46.625 76.405 46.955 ;
        RECT 76.745 46.085 76.915 47.495 ;
        RECT 68.450 45.915 76.915 46.085 ;
        RECT 68.450 45.400 70.180 45.915 ;
        RECT 68.450 45.285 79.930 45.400 ;
        RECT 65.820 40.085 67.820 40.255 ;
        RECT 68.450 39.745 68.620 45.285 ;
        RECT 61.590 39.575 68.620 39.745 ;
        RECT 68.900 45.230 79.930 45.285 ;
        RECT 68.900 39.740 69.070 45.230 ;
        RECT 69.700 44.720 73.700 44.890 ;
        RECT 69.470 40.465 69.640 44.505 ;
        RECT 73.760 40.465 73.930 44.505 ;
        RECT 69.700 40.080 73.700 40.250 ;
        RECT 74.330 39.740 74.500 45.230 ;
        RECT 75.130 44.720 79.130 44.890 ;
        RECT 74.900 40.465 75.070 44.505 ;
        RECT 79.190 40.465 79.360 44.505 ;
        RECT 75.130 40.080 79.130 40.250 ;
        RECT 79.760 39.740 79.930 45.230 ;
        RECT 68.900 39.570 79.930 39.740 ;
        RECT 80.205 45.245 81.955 45.415 ;
        RECT 80.205 39.755 80.375 45.245 ;
        RECT 80.915 44.735 81.245 44.905 ;
        RECT 80.775 40.480 80.945 44.520 ;
        RECT 81.215 40.480 81.385 44.520 ;
        RECT 80.915 40.095 81.245 40.265 ;
        RECT 81.785 39.755 81.955 45.245 ;
        RECT 80.205 39.585 81.955 39.755 ;
        RECT 82.230 39.760 82.400 49.250 ;
        RECT 82.940 48.740 83.270 48.910 ;
        RECT 82.800 40.485 82.970 48.525 ;
        RECT 83.240 40.485 83.410 48.525 ;
        RECT 82.940 40.100 83.270 40.270 ;
        RECT 83.810 39.760 83.980 49.250 ;
        RECT 85.435 49.260 111.980 49.420 ;
        RECT 85.435 49.235 98.180 49.260 ;
        RECT 85.435 49.005 89.760 49.235 ;
        RECT 82.230 39.590 83.980 39.760 ;
        RECT 85.470 39.745 85.640 49.005 ;
        RECT 86.365 48.435 88.405 48.605 ;
        RECT 85.980 40.375 86.150 48.375 ;
        RECT 88.620 40.375 88.790 48.375 ;
        RECT 86.365 40.145 88.405 40.315 ;
        RECT 89.130 39.745 89.300 49.005 ;
        RECT 85.470 39.575 89.300 39.745 ;
        RECT 89.590 39.745 89.760 49.005 ;
        RECT 90.390 48.725 92.390 48.895 ;
        RECT 90.160 40.470 90.330 48.510 ;
        RECT 92.450 40.470 92.620 48.510 ;
        RECT 90.390 40.085 92.390 40.255 ;
        RECT 93.020 39.745 93.190 49.235 ;
        RECT 93.820 48.725 95.820 48.895 ;
        RECT 93.590 40.470 93.760 48.510 ;
        RECT 95.880 40.470 96.050 48.510 ;
        RECT 96.450 47.665 98.180 49.235 ;
        RECT 110.230 49.250 111.980 49.260 ;
        RECT 96.450 47.495 104.915 47.665 ;
        RECT 96.450 46.085 98.255 47.495 ;
        RECT 98.595 46.625 98.765 46.955 ;
        RECT 98.980 46.925 104.020 47.095 ;
        RECT 98.980 46.485 104.020 46.655 ;
        RECT 104.235 46.625 104.405 46.955 ;
        RECT 104.745 46.085 104.915 47.495 ;
        RECT 96.450 45.915 104.915 46.085 ;
        RECT 96.450 45.400 98.180 45.915 ;
        RECT 96.450 45.285 107.930 45.400 ;
        RECT 93.820 40.085 95.820 40.255 ;
        RECT 96.450 39.745 96.620 45.285 ;
        RECT 89.590 39.575 96.620 39.745 ;
        RECT 96.900 45.230 107.930 45.285 ;
        RECT 96.900 39.740 97.070 45.230 ;
        RECT 97.700 44.720 101.700 44.890 ;
        RECT 97.470 40.465 97.640 44.505 ;
        RECT 101.760 40.465 101.930 44.505 ;
        RECT 97.700 40.080 101.700 40.250 ;
        RECT 102.330 39.740 102.500 45.230 ;
        RECT 103.130 44.720 107.130 44.890 ;
        RECT 102.900 40.465 103.070 44.505 ;
        RECT 107.190 40.465 107.360 44.505 ;
        RECT 103.130 40.080 107.130 40.250 ;
        RECT 107.760 39.740 107.930 45.230 ;
        RECT 96.900 39.570 107.930 39.740 ;
        RECT 108.205 45.245 109.955 45.415 ;
        RECT 108.205 39.755 108.375 45.245 ;
        RECT 108.915 44.735 109.245 44.905 ;
        RECT 108.775 40.480 108.945 44.520 ;
        RECT 109.215 40.480 109.385 44.520 ;
        RECT 108.915 40.095 109.245 40.265 ;
        RECT 109.785 39.755 109.955 45.245 ;
        RECT 108.205 39.585 109.955 39.755 ;
        RECT 110.230 39.760 110.400 49.250 ;
        RECT 110.940 48.740 111.270 48.910 ;
        RECT 110.800 40.485 110.970 48.525 ;
        RECT 111.240 40.485 111.410 48.525 ;
        RECT 110.940 40.100 111.270 40.270 ;
        RECT 111.810 39.760 111.980 49.250 ;
        RECT 113.435 49.260 139.980 49.420 ;
        RECT 113.435 49.235 126.180 49.260 ;
        RECT 113.435 49.005 117.760 49.235 ;
        RECT 110.230 39.590 111.980 39.760 ;
        RECT 113.470 39.745 113.640 49.005 ;
        RECT 114.365 48.435 116.405 48.605 ;
        RECT 113.980 40.375 114.150 48.375 ;
        RECT 116.620 40.375 116.790 48.375 ;
        RECT 114.365 40.145 116.405 40.315 ;
        RECT 117.130 39.745 117.300 49.005 ;
        RECT 113.470 39.575 117.300 39.745 ;
        RECT 117.590 39.745 117.760 49.005 ;
        RECT 118.390 48.725 120.390 48.895 ;
        RECT 118.160 40.470 118.330 48.510 ;
        RECT 120.450 40.470 120.620 48.510 ;
        RECT 118.390 40.085 120.390 40.255 ;
        RECT 121.020 39.745 121.190 49.235 ;
        RECT 121.820 48.725 123.820 48.895 ;
        RECT 121.590 40.470 121.760 48.510 ;
        RECT 123.880 40.470 124.050 48.510 ;
        RECT 124.450 47.665 126.180 49.235 ;
        RECT 138.230 49.250 139.980 49.260 ;
        RECT 124.450 47.495 132.915 47.665 ;
        RECT 124.450 46.085 126.255 47.495 ;
        RECT 126.595 46.625 126.765 46.955 ;
        RECT 126.980 46.925 132.020 47.095 ;
        RECT 126.980 46.485 132.020 46.655 ;
        RECT 132.235 46.625 132.405 46.955 ;
        RECT 132.745 46.085 132.915 47.495 ;
        RECT 124.450 45.915 132.915 46.085 ;
        RECT 124.450 45.400 126.180 45.915 ;
        RECT 124.450 45.285 135.930 45.400 ;
        RECT 121.820 40.085 123.820 40.255 ;
        RECT 124.450 39.745 124.620 45.285 ;
        RECT 117.590 39.575 124.620 39.745 ;
        RECT 124.900 45.230 135.930 45.285 ;
        RECT 124.900 39.740 125.070 45.230 ;
        RECT 125.700 44.720 129.700 44.890 ;
        RECT 125.470 40.465 125.640 44.505 ;
        RECT 129.760 40.465 129.930 44.505 ;
        RECT 125.700 40.080 129.700 40.250 ;
        RECT 130.330 39.740 130.500 45.230 ;
        RECT 131.130 44.720 135.130 44.890 ;
        RECT 130.900 40.465 131.070 44.505 ;
        RECT 135.190 40.465 135.360 44.505 ;
        RECT 131.130 40.080 135.130 40.250 ;
        RECT 135.760 39.740 135.930 45.230 ;
        RECT 124.900 39.570 135.930 39.740 ;
        RECT 136.205 45.245 137.955 45.415 ;
        RECT 136.205 39.755 136.375 45.245 ;
        RECT 136.915 44.735 137.245 44.905 ;
        RECT 136.775 40.480 136.945 44.520 ;
        RECT 137.215 40.480 137.385 44.520 ;
        RECT 136.915 40.095 137.245 40.265 ;
        RECT 137.785 39.755 137.955 45.245 ;
        RECT 136.205 39.585 137.955 39.755 ;
        RECT 138.230 39.760 138.400 49.250 ;
        RECT 138.940 48.740 139.270 48.910 ;
        RECT 138.800 40.485 138.970 48.525 ;
        RECT 139.240 40.485 139.410 48.525 ;
        RECT 138.940 40.100 139.270 40.270 ;
        RECT 139.810 39.760 139.980 49.250 ;
        RECT 143.470 48.190 143.640 49.840 ;
        RECT 144.120 48.670 146.280 49.360 ;
        RECT 146.810 48.670 148.970 49.360 ;
        RECT 149.450 48.190 149.620 49.840 ;
        RECT 143.470 48.020 149.620 48.190 ;
        RECT 143.470 46.370 143.640 48.020 ;
        RECT 144.120 46.850 146.280 47.540 ;
        RECT 146.810 46.850 148.970 47.540 ;
        RECT 149.450 46.370 149.620 48.020 ;
        RECT 143.470 46.200 149.620 46.370 ;
        RECT 143.470 44.550 143.640 46.200 ;
        RECT 144.120 45.030 146.280 45.720 ;
        RECT 146.810 45.030 148.970 45.720 ;
        RECT 149.450 44.550 149.620 46.200 ;
        RECT 143.470 44.380 155.600 44.550 ;
        RECT 143.470 42.730 143.640 44.380 ;
        RECT 144.120 43.210 146.280 43.900 ;
        RECT 146.810 43.210 148.970 43.900 ;
        RECT 149.450 42.730 149.620 44.380 ;
        RECT 150.100 43.210 152.260 43.900 ;
        RECT 152.790 43.210 154.950 43.900 ;
        RECT 155.430 42.730 155.600 44.380 ;
        RECT 143.470 42.560 155.600 42.730 ;
        RECT 143.470 40.910 143.640 42.560 ;
        RECT 144.120 41.390 146.280 42.080 ;
        RECT 146.810 41.390 148.970 42.080 ;
        RECT 149.450 40.910 149.620 42.560 ;
        RECT 150.100 41.390 152.260 42.080 ;
        RECT 152.790 41.390 154.950 42.080 ;
        RECT 155.430 40.910 155.600 42.560 ;
        RECT 143.470 40.740 155.600 40.910 ;
        RECT 150.780 40.250 154.340 40.740 ;
        RECT 138.230 39.590 139.980 39.760 ;
        RECT 2.130 38.665 24.020 38.835 ;
        RECT 2.130 35.265 2.300 38.665 ;
        RECT 2.930 38.155 6.930 38.325 ;
        RECT 2.700 35.945 2.870 37.985 ;
        RECT 6.990 35.945 7.160 37.985 ;
        RECT 2.930 35.605 6.930 35.775 ;
        RECT 7.560 35.265 7.730 38.665 ;
        RECT 8.360 38.155 12.360 38.325 ;
        RECT 8.130 35.945 8.300 37.985 ;
        RECT 12.420 35.945 12.590 37.985 ;
        RECT 8.360 35.605 12.360 35.775 ;
        RECT 12.990 35.265 13.160 38.665 ;
        RECT 13.790 38.155 17.790 38.325 ;
        RECT 13.560 35.945 13.730 37.985 ;
        RECT 17.850 35.945 18.020 37.985 ;
        RECT 13.790 35.605 17.790 35.775 ;
        RECT 18.420 35.265 18.590 38.665 ;
        RECT 19.220 38.155 23.220 38.325 ;
        RECT 18.990 35.945 19.160 37.985 ;
        RECT 23.280 35.945 23.450 37.985 ;
        RECT 23.850 36.240 24.020 38.665 ;
        RECT 24.290 38.670 26.040 38.840 ;
        RECT 24.290 36.270 24.460 38.670 ;
        RECT 25.000 38.160 25.330 38.330 ;
        RECT 24.860 36.950 25.030 37.990 ;
        RECT 25.300 36.950 25.470 37.990 ;
        RECT 25.000 36.610 25.330 36.780 ;
        RECT 25.870 36.270 26.040 38.670 ;
        RECT 24.290 36.240 26.040 36.270 ;
        RECT 26.315 38.675 28.065 38.845 ;
        RECT 26.315 36.240 26.485 38.675 ;
        RECT 27.025 38.165 27.355 38.335 ;
        RECT 19.220 35.605 23.220 35.775 ;
        RECT 23.850 35.275 26.485 36.240 ;
        RECT 26.885 35.955 27.055 37.995 ;
        RECT 27.325 35.955 27.495 37.995 ;
        RECT 27.025 35.615 27.355 35.785 ;
        RECT 27.895 35.275 28.065 38.675 ;
        RECT 23.850 35.265 28.065 35.275 ;
        RECT 2.130 35.245 28.065 35.265 ;
        RECT 30.130 38.665 52.020 38.835 ;
        RECT 30.130 35.265 30.300 38.665 ;
        RECT 30.930 38.155 34.930 38.325 ;
        RECT 30.700 35.945 30.870 37.985 ;
        RECT 34.990 35.945 35.160 37.985 ;
        RECT 30.930 35.605 34.930 35.775 ;
        RECT 35.560 35.265 35.730 38.665 ;
        RECT 36.360 38.155 40.360 38.325 ;
        RECT 36.130 35.945 36.300 37.985 ;
        RECT 40.420 35.945 40.590 37.985 ;
        RECT 36.360 35.605 40.360 35.775 ;
        RECT 40.990 35.265 41.160 38.665 ;
        RECT 41.790 38.155 45.790 38.325 ;
        RECT 41.560 35.945 41.730 37.985 ;
        RECT 45.850 35.945 46.020 37.985 ;
        RECT 41.790 35.605 45.790 35.775 ;
        RECT 46.420 35.265 46.590 38.665 ;
        RECT 47.220 38.155 51.220 38.325 ;
        RECT 46.990 35.945 47.160 37.985 ;
        RECT 51.280 35.945 51.450 37.985 ;
        RECT 51.850 36.240 52.020 38.665 ;
        RECT 52.290 38.670 54.040 38.840 ;
        RECT 52.290 36.270 52.460 38.670 ;
        RECT 53.000 38.160 53.330 38.330 ;
        RECT 52.860 36.950 53.030 37.990 ;
        RECT 53.300 36.950 53.470 37.990 ;
        RECT 53.000 36.610 53.330 36.780 ;
        RECT 53.870 36.270 54.040 38.670 ;
        RECT 52.290 36.240 54.040 36.270 ;
        RECT 54.315 38.675 56.065 38.845 ;
        RECT 54.315 36.240 54.485 38.675 ;
        RECT 55.025 38.165 55.355 38.335 ;
        RECT 47.220 35.605 51.220 35.775 ;
        RECT 51.850 35.275 54.485 36.240 ;
        RECT 54.885 35.955 55.055 37.995 ;
        RECT 55.325 35.955 55.495 37.995 ;
        RECT 55.025 35.615 55.355 35.785 ;
        RECT 55.895 35.275 56.065 38.675 ;
        RECT 51.850 35.265 56.065 35.275 ;
        RECT 30.130 35.245 56.065 35.265 ;
        RECT 58.130 38.665 80.020 38.835 ;
        RECT 58.130 35.265 58.300 38.665 ;
        RECT 58.930 38.155 62.930 38.325 ;
        RECT 58.700 35.945 58.870 37.985 ;
        RECT 62.990 35.945 63.160 37.985 ;
        RECT 58.930 35.605 62.930 35.775 ;
        RECT 63.560 35.265 63.730 38.665 ;
        RECT 64.360 38.155 68.360 38.325 ;
        RECT 64.130 35.945 64.300 37.985 ;
        RECT 68.420 35.945 68.590 37.985 ;
        RECT 64.360 35.605 68.360 35.775 ;
        RECT 68.990 35.265 69.160 38.665 ;
        RECT 69.790 38.155 73.790 38.325 ;
        RECT 69.560 35.945 69.730 37.985 ;
        RECT 73.850 35.945 74.020 37.985 ;
        RECT 69.790 35.605 73.790 35.775 ;
        RECT 74.420 35.265 74.590 38.665 ;
        RECT 75.220 38.155 79.220 38.325 ;
        RECT 74.990 35.945 75.160 37.985 ;
        RECT 79.280 35.945 79.450 37.985 ;
        RECT 79.850 36.240 80.020 38.665 ;
        RECT 80.290 38.670 82.040 38.840 ;
        RECT 80.290 36.270 80.460 38.670 ;
        RECT 81.000 38.160 81.330 38.330 ;
        RECT 80.860 36.950 81.030 37.990 ;
        RECT 81.300 36.950 81.470 37.990 ;
        RECT 81.000 36.610 81.330 36.780 ;
        RECT 81.870 36.270 82.040 38.670 ;
        RECT 80.290 36.240 82.040 36.270 ;
        RECT 82.315 38.675 84.065 38.845 ;
        RECT 82.315 36.240 82.485 38.675 ;
        RECT 83.025 38.165 83.355 38.335 ;
        RECT 75.220 35.605 79.220 35.775 ;
        RECT 79.850 35.275 82.485 36.240 ;
        RECT 82.885 35.955 83.055 37.995 ;
        RECT 83.325 35.955 83.495 37.995 ;
        RECT 83.025 35.615 83.355 35.785 ;
        RECT 83.895 35.275 84.065 38.675 ;
        RECT 79.850 35.265 84.065 35.275 ;
        RECT 58.130 35.245 84.065 35.265 ;
        RECT 86.130 38.665 108.020 38.835 ;
        RECT 86.130 35.265 86.300 38.665 ;
        RECT 86.930 38.155 90.930 38.325 ;
        RECT 86.700 35.945 86.870 37.985 ;
        RECT 90.990 35.945 91.160 37.985 ;
        RECT 86.930 35.605 90.930 35.775 ;
        RECT 91.560 35.265 91.730 38.665 ;
        RECT 92.360 38.155 96.360 38.325 ;
        RECT 92.130 35.945 92.300 37.985 ;
        RECT 96.420 35.945 96.590 37.985 ;
        RECT 92.360 35.605 96.360 35.775 ;
        RECT 96.990 35.265 97.160 38.665 ;
        RECT 97.790 38.155 101.790 38.325 ;
        RECT 97.560 35.945 97.730 37.985 ;
        RECT 101.850 35.945 102.020 37.985 ;
        RECT 97.790 35.605 101.790 35.775 ;
        RECT 102.420 35.265 102.590 38.665 ;
        RECT 103.220 38.155 107.220 38.325 ;
        RECT 102.990 35.945 103.160 37.985 ;
        RECT 107.280 35.945 107.450 37.985 ;
        RECT 107.850 36.240 108.020 38.665 ;
        RECT 108.290 38.670 110.040 38.840 ;
        RECT 108.290 36.270 108.460 38.670 ;
        RECT 109.000 38.160 109.330 38.330 ;
        RECT 108.860 36.950 109.030 37.990 ;
        RECT 109.300 36.950 109.470 37.990 ;
        RECT 109.000 36.610 109.330 36.780 ;
        RECT 109.870 36.270 110.040 38.670 ;
        RECT 108.290 36.240 110.040 36.270 ;
        RECT 110.315 38.675 112.065 38.845 ;
        RECT 110.315 36.240 110.485 38.675 ;
        RECT 111.025 38.165 111.355 38.335 ;
        RECT 103.220 35.605 107.220 35.775 ;
        RECT 107.850 35.275 110.485 36.240 ;
        RECT 110.885 35.955 111.055 37.995 ;
        RECT 111.325 35.955 111.495 37.995 ;
        RECT 111.025 35.615 111.355 35.785 ;
        RECT 111.895 35.275 112.065 38.675 ;
        RECT 107.850 35.265 112.065 35.275 ;
        RECT 86.130 35.245 112.065 35.265 ;
        RECT 114.130 38.665 136.020 38.835 ;
        RECT 114.130 35.265 114.300 38.665 ;
        RECT 114.930 38.155 118.930 38.325 ;
        RECT 114.700 35.945 114.870 37.985 ;
        RECT 118.990 35.945 119.160 37.985 ;
        RECT 114.930 35.605 118.930 35.775 ;
        RECT 119.560 35.265 119.730 38.665 ;
        RECT 120.360 38.155 124.360 38.325 ;
        RECT 120.130 35.945 120.300 37.985 ;
        RECT 124.420 35.945 124.590 37.985 ;
        RECT 120.360 35.605 124.360 35.775 ;
        RECT 124.990 35.265 125.160 38.665 ;
        RECT 125.790 38.155 129.790 38.325 ;
        RECT 125.560 35.945 125.730 37.985 ;
        RECT 129.850 35.945 130.020 37.985 ;
        RECT 125.790 35.605 129.790 35.775 ;
        RECT 130.420 35.265 130.590 38.665 ;
        RECT 131.220 38.155 135.220 38.325 ;
        RECT 130.990 35.945 131.160 37.985 ;
        RECT 135.280 35.945 135.450 37.985 ;
        RECT 135.850 36.240 136.020 38.665 ;
        RECT 136.290 38.670 138.040 38.840 ;
        RECT 136.290 36.270 136.460 38.670 ;
        RECT 137.000 38.160 137.330 38.330 ;
        RECT 136.860 36.950 137.030 37.990 ;
        RECT 137.300 36.950 137.470 37.990 ;
        RECT 137.000 36.610 137.330 36.780 ;
        RECT 137.870 36.270 138.040 38.670 ;
        RECT 136.290 36.240 138.040 36.270 ;
        RECT 138.315 38.675 140.065 38.845 ;
        RECT 138.315 36.240 138.485 38.675 ;
        RECT 139.025 38.165 139.355 38.335 ;
        RECT 131.220 35.605 135.220 35.775 ;
        RECT 135.850 35.275 138.485 36.240 ;
        RECT 138.885 35.955 139.055 37.995 ;
        RECT 139.325 35.955 139.495 37.995 ;
        RECT 139.025 35.615 139.355 35.785 ;
        RECT 139.895 35.275 140.065 38.675 ;
        RECT 135.850 35.265 140.065 35.275 ;
        RECT 114.130 35.245 140.065 35.265 ;
        RECT 1.475 35.105 28.065 35.245 ;
        RECT 29.475 35.105 56.065 35.245 ;
        RECT 57.475 35.105 84.065 35.245 ;
        RECT 85.475 35.105 112.065 35.245 ;
        RECT 113.475 35.105 140.065 35.245 ;
        RECT 1.475 34.380 28.055 35.105 ;
        RECT 29.475 34.380 56.055 35.105 ;
        RECT 57.475 34.380 84.055 35.105 ;
        RECT 85.475 34.380 112.055 35.105 ;
        RECT 113.475 34.380 140.055 35.105 ;
        RECT 1.450 33.480 27.925 33.960 ;
        RECT 29.450 33.480 55.925 33.960 ;
        RECT 57.450 33.480 83.925 33.960 ;
        RECT 85.450 33.480 111.925 33.960 ;
        RECT 113.450 33.480 139.925 33.960 ;
        RECT 1.435 33.420 27.925 33.480 ;
        RECT 29.435 33.420 55.925 33.480 ;
        RECT 57.435 33.420 83.925 33.480 ;
        RECT 85.435 33.420 111.925 33.480 ;
        RECT 113.435 33.420 139.925 33.480 ;
        RECT 1.435 33.260 27.980 33.420 ;
        RECT 1.435 33.235 14.180 33.260 ;
        RECT 1.435 33.005 5.760 33.235 ;
        RECT 1.470 23.745 1.640 33.005 ;
        RECT 2.365 32.435 4.405 32.605 ;
        RECT 1.980 24.375 2.150 32.375 ;
        RECT 4.620 24.375 4.790 32.375 ;
        RECT 2.365 24.145 4.405 24.315 ;
        RECT 5.130 23.745 5.300 33.005 ;
        RECT 1.470 23.575 5.300 23.745 ;
        RECT 5.590 23.745 5.760 33.005 ;
        RECT 6.390 32.725 8.390 32.895 ;
        RECT 6.160 24.470 6.330 32.510 ;
        RECT 8.450 24.470 8.620 32.510 ;
        RECT 6.390 24.085 8.390 24.255 ;
        RECT 9.020 23.745 9.190 33.235 ;
        RECT 9.820 32.725 11.820 32.895 ;
        RECT 9.590 24.470 9.760 32.510 ;
        RECT 11.880 24.470 12.050 32.510 ;
        RECT 12.450 31.665 14.180 33.235 ;
        RECT 26.230 33.250 27.980 33.260 ;
        RECT 12.450 31.495 20.915 31.665 ;
        RECT 12.450 30.085 14.255 31.495 ;
        RECT 14.595 30.625 14.765 30.955 ;
        RECT 14.980 30.925 20.020 31.095 ;
        RECT 14.980 30.485 20.020 30.655 ;
        RECT 20.235 30.625 20.405 30.955 ;
        RECT 20.745 30.085 20.915 31.495 ;
        RECT 12.450 29.915 20.915 30.085 ;
        RECT 12.450 29.400 14.180 29.915 ;
        RECT 12.450 29.285 23.930 29.400 ;
        RECT 9.820 24.085 11.820 24.255 ;
        RECT 12.450 23.745 12.620 29.285 ;
        RECT 5.590 23.575 12.620 23.745 ;
        RECT 12.900 29.230 23.930 29.285 ;
        RECT 12.900 23.740 13.070 29.230 ;
        RECT 13.700 28.720 17.700 28.890 ;
        RECT 13.470 24.465 13.640 28.505 ;
        RECT 17.760 24.465 17.930 28.505 ;
        RECT 13.700 24.080 17.700 24.250 ;
        RECT 18.330 23.740 18.500 29.230 ;
        RECT 19.130 28.720 23.130 28.890 ;
        RECT 18.900 24.465 19.070 28.505 ;
        RECT 23.190 24.465 23.360 28.505 ;
        RECT 19.130 24.080 23.130 24.250 ;
        RECT 23.760 23.740 23.930 29.230 ;
        RECT 12.900 23.570 23.930 23.740 ;
        RECT 24.205 29.245 25.955 29.415 ;
        RECT 24.205 23.755 24.375 29.245 ;
        RECT 24.915 28.735 25.245 28.905 ;
        RECT 24.775 24.480 24.945 28.520 ;
        RECT 25.215 24.480 25.385 28.520 ;
        RECT 24.915 24.095 25.245 24.265 ;
        RECT 25.785 23.755 25.955 29.245 ;
        RECT 24.205 23.585 25.955 23.755 ;
        RECT 26.230 23.760 26.400 33.250 ;
        RECT 26.940 32.740 27.270 32.910 ;
        RECT 26.800 24.485 26.970 32.525 ;
        RECT 27.240 24.485 27.410 32.525 ;
        RECT 26.940 24.100 27.270 24.270 ;
        RECT 27.810 23.760 27.980 33.250 ;
        RECT 29.435 33.260 55.980 33.420 ;
        RECT 29.435 33.235 42.180 33.260 ;
        RECT 29.435 33.005 33.760 33.235 ;
        RECT 26.230 23.590 27.980 23.760 ;
        RECT 29.470 23.745 29.640 33.005 ;
        RECT 30.365 32.435 32.405 32.605 ;
        RECT 29.980 24.375 30.150 32.375 ;
        RECT 32.620 24.375 32.790 32.375 ;
        RECT 30.365 24.145 32.405 24.315 ;
        RECT 33.130 23.745 33.300 33.005 ;
        RECT 29.470 23.575 33.300 23.745 ;
        RECT 33.590 23.745 33.760 33.005 ;
        RECT 34.390 32.725 36.390 32.895 ;
        RECT 34.160 24.470 34.330 32.510 ;
        RECT 36.450 24.470 36.620 32.510 ;
        RECT 34.390 24.085 36.390 24.255 ;
        RECT 37.020 23.745 37.190 33.235 ;
        RECT 37.820 32.725 39.820 32.895 ;
        RECT 37.590 24.470 37.760 32.510 ;
        RECT 39.880 24.470 40.050 32.510 ;
        RECT 40.450 31.665 42.180 33.235 ;
        RECT 54.230 33.250 55.980 33.260 ;
        RECT 40.450 31.495 48.915 31.665 ;
        RECT 40.450 30.085 42.255 31.495 ;
        RECT 42.595 30.625 42.765 30.955 ;
        RECT 42.980 30.925 48.020 31.095 ;
        RECT 42.980 30.485 48.020 30.655 ;
        RECT 48.235 30.625 48.405 30.955 ;
        RECT 48.745 30.085 48.915 31.495 ;
        RECT 40.450 29.915 48.915 30.085 ;
        RECT 40.450 29.400 42.180 29.915 ;
        RECT 40.450 29.285 51.930 29.400 ;
        RECT 37.820 24.085 39.820 24.255 ;
        RECT 40.450 23.745 40.620 29.285 ;
        RECT 33.590 23.575 40.620 23.745 ;
        RECT 40.900 29.230 51.930 29.285 ;
        RECT 40.900 23.740 41.070 29.230 ;
        RECT 41.700 28.720 45.700 28.890 ;
        RECT 41.470 24.465 41.640 28.505 ;
        RECT 45.760 24.465 45.930 28.505 ;
        RECT 41.700 24.080 45.700 24.250 ;
        RECT 46.330 23.740 46.500 29.230 ;
        RECT 47.130 28.720 51.130 28.890 ;
        RECT 46.900 24.465 47.070 28.505 ;
        RECT 51.190 24.465 51.360 28.505 ;
        RECT 47.130 24.080 51.130 24.250 ;
        RECT 51.760 23.740 51.930 29.230 ;
        RECT 40.900 23.570 51.930 23.740 ;
        RECT 52.205 29.245 53.955 29.415 ;
        RECT 52.205 23.755 52.375 29.245 ;
        RECT 52.915 28.735 53.245 28.905 ;
        RECT 52.775 24.480 52.945 28.520 ;
        RECT 53.215 24.480 53.385 28.520 ;
        RECT 52.915 24.095 53.245 24.265 ;
        RECT 53.785 23.755 53.955 29.245 ;
        RECT 52.205 23.585 53.955 23.755 ;
        RECT 54.230 23.760 54.400 33.250 ;
        RECT 54.940 32.740 55.270 32.910 ;
        RECT 54.800 24.485 54.970 32.525 ;
        RECT 55.240 24.485 55.410 32.525 ;
        RECT 54.940 24.100 55.270 24.270 ;
        RECT 55.810 23.760 55.980 33.250 ;
        RECT 57.435 33.260 83.980 33.420 ;
        RECT 57.435 33.235 70.180 33.260 ;
        RECT 57.435 33.005 61.760 33.235 ;
        RECT 54.230 23.590 55.980 23.760 ;
        RECT 57.470 23.745 57.640 33.005 ;
        RECT 58.365 32.435 60.405 32.605 ;
        RECT 57.980 24.375 58.150 32.375 ;
        RECT 60.620 24.375 60.790 32.375 ;
        RECT 58.365 24.145 60.405 24.315 ;
        RECT 61.130 23.745 61.300 33.005 ;
        RECT 57.470 23.575 61.300 23.745 ;
        RECT 61.590 23.745 61.760 33.005 ;
        RECT 62.390 32.725 64.390 32.895 ;
        RECT 62.160 24.470 62.330 32.510 ;
        RECT 64.450 24.470 64.620 32.510 ;
        RECT 62.390 24.085 64.390 24.255 ;
        RECT 65.020 23.745 65.190 33.235 ;
        RECT 65.820 32.725 67.820 32.895 ;
        RECT 65.590 24.470 65.760 32.510 ;
        RECT 67.880 24.470 68.050 32.510 ;
        RECT 68.450 31.665 70.180 33.235 ;
        RECT 82.230 33.250 83.980 33.260 ;
        RECT 68.450 31.495 76.915 31.665 ;
        RECT 68.450 30.085 70.255 31.495 ;
        RECT 70.595 30.625 70.765 30.955 ;
        RECT 70.980 30.925 76.020 31.095 ;
        RECT 70.980 30.485 76.020 30.655 ;
        RECT 76.235 30.625 76.405 30.955 ;
        RECT 76.745 30.085 76.915 31.495 ;
        RECT 68.450 29.915 76.915 30.085 ;
        RECT 68.450 29.400 70.180 29.915 ;
        RECT 68.450 29.285 79.930 29.400 ;
        RECT 65.820 24.085 67.820 24.255 ;
        RECT 68.450 23.745 68.620 29.285 ;
        RECT 61.590 23.575 68.620 23.745 ;
        RECT 68.900 29.230 79.930 29.285 ;
        RECT 68.900 23.740 69.070 29.230 ;
        RECT 69.700 28.720 73.700 28.890 ;
        RECT 69.470 24.465 69.640 28.505 ;
        RECT 73.760 24.465 73.930 28.505 ;
        RECT 69.700 24.080 73.700 24.250 ;
        RECT 74.330 23.740 74.500 29.230 ;
        RECT 75.130 28.720 79.130 28.890 ;
        RECT 74.900 24.465 75.070 28.505 ;
        RECT 79.190 24.465 79.360 28.505 ;
        RECT 75.130 24.080 79.130 24.250 ;
        RECT 79.760 23.740 79.930 29.230 ;
        RECT 68.900 23.570 79.930 23.740 ;
        RECT 80.205 29.245 81.955 29.415 ;
        RECT 80.205 23.755 80.375 29.245 ;
        RECT 80.915 28.735 81.245 28.905 ;
        RECT 80.775 24.480 80.945 28.520 ;
        RECT 81.215 24.480 81.385 28.520 ;
        RECT 80.915 24.095 81.245 24.265 ;
        RECT 81.785 23.755 81.955 29.245 ;
        RECT 80.205 23.585 81.955 23.755 ;
        RECT 82.230 23.760 82.400 33.250 ;
        RECT 82.940 32.740 83.270 32.910 ;
        RECT 82.800 24.485 82.970 32.525 ;
        RECT 83.240 24.485 83.410 32.525 ;
        RECT 82.940 24.100 83.270 24.270 ;
        RECT 83.810 23.760 83.980 33.250 ;
        RECT 85.435 33.260 111.980 33.420 ;
        RECT 85.435 33.235 98.180 33.260 ;
        RECT 85.435 33.005 89.760 33.235 ;
        RECT 82.230 23.590 83.980 23.760 ;
        RECT 85.470 23.745 85.640 33.005 ;
        RECT 86.365 32.435 88.405 32.605 ;
        RECT 85.980 24.375 86.150 32.375 ;
        RECT 88.620 24.375 88.790 32.375 ;
        RECT 86.365 24.145 88.405 24.315 ;
        RECT 89.130 23.745 89.300 33.005 ;
        RECT 85.470 23.575 89.300 23.745 ;
        RECT 89.590 23.745 89.760 33.005 ;
        RECT 90.390 32.725 92.390 32.895 ;
        RECT 90.160 24.470 90.330 32.510 ;
        RECT 92.450 24.470 92.620 32.510 ;
        RECT 90.390 24.085 92.390 24.255 ;
        RECT 93.020 23.745 93.190 33.235 ;
        RECT 93.820 32.725 95.820 32.895 ;
        RECT 93.590 24.470 93.760 32.510 ;
        RECT 95.880 24.470 96.050 32.510 ;
        RECT 96.450 31.665 98.180 33.235 ;
        RECT 110.230 33.250 111.980 33.260 ;
        RECT 96.450 31.495 104.915 31.665 ;
        RECT 96.450 30.085 98.255 31.495 ;
        RECT 98.595 30.625 98.765 30.955 ;
        RECT 98.980 30.925 104.020 31.095 ;
        RECT 98.980 30.485 104.020 30.655 ;
        RECT 104.235 30.625 104.405 30.955 ;
        RECT 104.745 30.085 104.915 31.495 ;
        RECT 96.450 29.915 104.915 30.085 ;
        RECT 96.450 29.400 98.180 29.915 ;
        RECT 96.450 29.285 107.930 29.400 ;
        RECT 93.820 24.085 95.820 24.255 ;
        RECT 96.450 23.745 96.620 29.285 ;
        RECT 89.590 23.575 96.620 23.745 ;
        RECT 96.900 29.230 107.930 29.285 ;
        RECT 96.900 23.740 97.070 29.230 ;
        RECT 97.700 28.720 101.700 28.890 ;
        RECT 97.470 24.465 97.640 28.505 ;
        RECT 101.760 24.465 101.930 28.505 ;
        RECT 97.700 24.080 101.700 24.250 ;
        RECT 102.330 23.740 102.500 29.230 ;
        RECT 103.130 28.720 107.130 28.890 ;
        RECT 102.900 24.465 103.070 28.505 ;
        RECT 107.190 24.465 107.360 28.505 ;
        RECT 103.130 24.080 107.130 24.250 ;
        RECT 107.760 23.740 107.930 29.230 ;
        RECT 96.900 23.570 107.930 23.740 ;
        RECT 108.205 29.245 109.955 29.415 ;
        RECT 108.205 23.755 108.375 29.245 ;
        RECT 108.915 28.735 109.245 28.905 ;
        RECT 108.775 24.480 108.945 28.520 ;
        RECT 109.215 24.480 109.385 28.520 ;
        RECT 108.915 24.095 109.245 24.265 ;
        RECT 109.785 23.755 109.955 29.245 ;
        RECT 108.205 23.585 109.955 23.755 ;
        RECT 110.230 23.760 110.400 33.250 ;
        RECT 110.940 32.740 111.270 32.910 ;
        RECT 110.800 24.485 110.970 32.525 ;
        RECT 111.240 24.485 111.410 32.525 ;
        RECT 110.940 24.100 111.270 24.270 ;
        RECT 111.810 23.760 111.980 33.250 ;
        RECT 113.435 33.260 139.980 33.420 ;
        RECT 113.435 33.235 126.180 33.260 ;
        RECT 113.435 33.005 117.760 33.235 ;
        RECT 110.230 23.590 111.980 23.760 ;
        RECT 113.470 23.745 113.640 33.005 ;
        RECT 114.365 32.435 116.405 32.605 ;
        RECT 113.980 24.375 114.150 32.375 ;
        RECT 116.620 24.375 116.790 32.375 ;
        RECT 114.365 24.145 116.405 24.315 ;
        RECT 117.130 23.745 117.300 33.005 ;
        RECT 113.470 23.575 117.300 23.745 ;
        RECT 117.590 23.745 117.760 33.005 ;
        RECT 118.390 32.725 120.390 32.895 ;
        RECT 118.160 24.470 118.330 32.510 ;
        RECT 120.450 24.470 120.620 32.510 ;
        RECT 118.390 24.085 120.390 24.255 ;
        RECT 121.020 23.745 121.190 33.235 ;
        RECT 121.820 32.725 123.820 32.895 ;
        RECT 121.590 24.470 121.760 32.510 ;
        RECT 123.880 24.470 124.050 32.510 ;
        RECT 124.450 31.665 126.180 33.235 ;
        RECT 138.230 33.250 139.980 33.260 ;
        RECT 124.450 31.495 132.915 31.665 ;
        RECT 124.450 30.085 126.255 31.495 ;
        RECT 126.595 30.625 126.765 30.955 ;
        RECT 126.980 30.925 132.020 31.095 ;
        RECT 126.980 30.485 132.020 30.655 ;
        RECT 132.235 30.625 132.405 30.955 ;
        RECT 132.745 30.085 132.915 31.495 ;
        RECT 124.450 29.915 132.915 30.085 ;
        RECT 124.450 29.400 126.180 29.915 ;
        RECT 124.450 29.285 135.930 29.400 ;
        RECT 121.820 24.085 123.820 24.255 ;
        RECT 124.450 23.745 124.620 29.285 ;
        RECT 117.590 23.575 124.620 23.745 ;
        RECT 124.900 29.230 135.930 29.285 ;
        RECT 124.900 23.740 125.070 29.230 ;
        RECT 125.700 28.720 129.700 28.890 ;
        RECT 125.470 24.465 125.640 28.505 ;
        RECT 129.760 24.465 129.930 28.505 ;
        RECT 125.700 24.080 129.700 24.250 ;
        RECT 130.330 23.740 130.500 29.230 ;
        RECT 131.130 28.720 135.130 28.890 ;
        RECT 130.900 24.465 131.070 28.505 ;
        RECT 135.190 24.465 135.360 28.505 ;
        RECT 131.130 24.080 135.130 24.250 ;
        RECT 135.760 23.740 135.930 29.230 ;
        RECT 124.900 23.570 135.930 23.740 ;
        RECT 136.205 29.245 137.955 29.415 ;
        RECT 136.205 23.755 136.375 29.245 ;
        RECT 136.915 28.735 137.245 28.905 ;
        RECT 136.775 24.480 136.945 28.520 ;
        RECT 137.215 24.480 137.385 28.520 ;
        RECT 136.915 24.095 137.245 24.265 ;
        RECT 137.785 23.755 137.955 29.245 ;
        RECT 136.205 23.585 137.955 23.755 ;
        RECT 138.230 23.760 138.400 33.250 ;
        RECT 138.940 32.740 139.270 32.910 ;
        RECT 138.800 24.485 138.970 32.525 ;
        RECT 139.240 24.485 139.410 32.525 ;
        RECT 138.940 24.100 139.270 24.270 ;
        RECT 139.810 23.760 139.980 33.250 ;
        RECT 138.230 23.590 139.980 23.760 ;
        RECT 2.130 22.665 24.020 22.835 ;
        RECT 2.130 19.265 2.300 22.665 ;
        RECT 2.930 22.155 6.930 22.325 ;
        RECT 2.700 19.945 2.870 21.985 ;
        RECT 6.990 19.945 7.160 21.985 ;
        RECT 2.930 19.605 6.930 19.775 ;
        RECT 7.560 19.265 7.730 22.665 ;
        RECT 8.360 22.155 12.360 22.325 ;
        RECT 8.130 19.945 8.300 21.985 ;
        RECT 12.420 19.945 12.590 21.985 ;
        RECT 8.360 19.605 12.360 19.775 ;
        RECT 12.990 19.265 13.160 22.665 ;
        RECT 13.790 22.155 17.790 22.325 ;
        RECT 13.560 19.945 13.730 21.985 ;
        RECT 17.850 19.945 18.020 21.985 ;
        RECT 13.790 19.605 17.790 19.775 ;
        RECT 18.420 19.265 18.590 22.665 ;
        RECT 19.220 22.155 23.220 22.325 ;
        RECT 18.990 19.945 19.160 21.985 ;
        RECT 23.280 19.945 23.450 21.985 ;
        RECT 23.850 20.240 24.020 22.665 ;
        RECT 24.290 22.670 26.040 22.840 ;
        RECT 24.290 20.270 24.460 22.670 ;
        RECT 25.000 22.160 25.330 22.330 ;
        RECT 24.860 20.950 25.030 21.990 ;
        RECT 25.300 20.950 25.470 21.990 ;
        RECT 25.000 20.610 25.330 20.780 ;
        RECT 25.870 20.270 26.040 22.670 ;
        RECT 24.290 20.240 26.040 20.270 ;
        RECT 26.315 22.675 28.065 22.845 ;
        RECT 26.315 20.240 26.485 22.675 ;
        RECT 27.025 22.165 27.355 22.335 ;
        RECT 19.220 19.605 23.220 19.775 ;
        RECT 23.850 19.275 26.485 20.240 ;
        RECT 26.885 19.955 27.055 21.995 ;
        RECT 27.325 19.955 27.495 21.995 ;
        RECT 27.025 19.615 27.355 19.785 ;
        RECT 27.895 19.275 28.065 22.675 ;
        RECT 23.850 19.265 28.065 19.275 ;
        RECT 2.130 19.245 28.065 19.265 ;
        RECT 30.130 22.665 52.020 22.835 ;
        RECT 30.130 19.265 30.300 22.665 ;
        RECT 30.930 22.155 34.930 22.325 ;
        RECT 30.700 19.945 30.870 21.985 ;
        RECT 34.990 19.945 35.160 21.985 ;
        RECT 30.930 19.605 34.930 19.775 ;
        RECT 35.560 19.265 35.730 22.665 ;
        RECT 36.360 22.155 40.360 22.325 ;
        RECT 36.130 19.945 36.300 21.985 ;
        RECT 40.420 19.945 40.590 21.985 ;
        RECT 36.360 19.605 40.360 19.775 ;
        RECT 40.990 19.265 41.160 22.665 ;
        RECT 41.790 22.155 45.790 22.325 ;
        RECT 41.560 19.945 41.730 21.985 ;
        RECT 45.850 19.945 46.020 21.985 ;
        RECT 41.790 19.605 45.790 19.775 ;
        RECT 46.420 19.265 46.590 22.665 ;
        RECT 47.220 22.155 51.220 22.325 ;
        RECT 46.990 19.945 47.160 21.985 ;
        RECT 51.280 19.945 51.450 21.985 ;
        RECT 51.850 20.240 52.020 22.665 ;
        RECT 52.290 22.670 54.040 22.840 ;
        RECT 52.290 20.270 52.460 22.670 ;
        RECT 53.000 22.160 53.330 22.330 ;
        RECT 52.860 20.950 53.030 21.990 ;
        RECT 53.300 20.950 53.470 21.990 ;
        RECT 53.000 20.610 53.330 20.780 ;
        RECT 53.870 20.270 54.040 22.670 ;
        RECT 52.290 20.240 54.040 20.270 ;
        RECT 54.315 22.675 56.065 22.845 ;
        RECT 54.315 20.240 54.485 22.675 ;
        RECT 55.025 22.165 55.355 22.335 ;
        RECT 47.220 19.605 51.220 19.775 ;
        RECT 51.850 19.275 54.485 20.240 ;
        RECT 54.885 19.955 55.055 21.995 ;
        RECT 55.325 19.955 55.495 21.995 ;
        RECT 55.025 19.615 55.355 19.785 ;
        RECT 55.895 19.275 56.065 22.675 ;
        RECT 51.850 19.265 56.065 19.275 ;
        RECT 30.130 19.245 56.065 19.265 ;
        RECT 58.130 22.665 80.020 22.835 ;
        RECT 58.130 19.265 58.300 22.665 ;
        RECT 58.930 22.155 62.930 22.325 ;
        RECT 58.700 19.945 58.870 21.985 ;
        RECT 62.990 19.945 63.160 21.985 ;
        RECT 58.930 19.605 62.930 19.775 ;
        RECT 63.560 19.265 63.730 22.665 ;
        RECT 64.360 22.155 68.360 22.325 ;
        RECT 64.130 19.945 64.300 21.985 ;
        RECT 68.420 19.945 68.590 21.985 ;
        RECT 64.360 19.605 68.360 19.775 ;
        RECT 68.990 19.265 69.160 22.665 ;
        RECT 69.790 22.155 73.790 22.325 ;
        RECT 69.560 19.945 69.730 21.985 ;
        RECT 73.850 19.945 74.020 21.985 ;
        RECT 69.790 19.605 73.790 19.775 ;
        RECT 74.420 19.265 74.590 22.665 ;
        RECT 75.220 22.155 79.220 22.325 ;
        RECT 74.990 19.945 75.160 21.985 ;
        RECT 79.280 19.945 79.450 21.985 ;
        RECT 79.850 20.240 80.020 22.665 ;
        RECT 80.290 22.670 82.040 22.840 ;
        RECT 80.290 20.270 80.460 22.670 ;
        RECT 81.000 22.160 81.330 22.330 ;
        RECT 80.860 20.950 81.030 21.990 ;
        RECT 81.300 20.950 81.470 21.990 ;
        RECT 81.000 20.610 81.330 20.780 ;
        RECT 81.870 20.270 82.040 22.670 ;
        RECT 80.290 20.240 82.040 20.270 ;
        RECT 82.315 22.675 84.065 22.845 ;
        RECT 82.315 20.240 82.485 22.675 ;
        RECT 83.025 22.165 83.355 22.335 ;
        RECT 75.220 19.605 79.220 19.775 ;
        RECT 79.850 19.275 82.485 20.240 ;
        RECT 82.885 19.955 83.055 21.995 ;
        RECT 83.325 19.955 83.495 21.995 ;
        RECT 83.025 19.615 83.355 19.785 ;
        RECT 83.895 19.275 84.065 22.675 ;
        RECT 79.850 19.265 84.065 19.275 ;
        RECT 58.130 19.245 84.065 19.265 ;
        RECT 86.130 22.665 108.020 22.835 ;
        RECT 86.130 19.265 86.300 22.665 ;
        RECT 86.930 22.155 90.930 22.325 ;
        RECT 86.700 19.945 86.870 21.985 ;
        RECT 90.990 19.945 91.160 21.985 ;
        RECT 86.930 19.605 90.930 19.775 ;
        RECT 91.560 19.265 91.730 22.665 ;
        RECT 92.360 22.155 96.360 22.325 ;
        RECT 92.130 19.945 92.300 21.985 ;
        RECT 96.420 19.945 96.590 21.985 ;
        RECT 92.360 19.605 96.360 19.775 ;
        RECT 96.990 19.265 97.160 22.665 ;
        RECT 97.790 22.155 101.790 22.325 ;
        RECT 97.560 19.945 97.730 21.985 ;
        RECT 101.850 19.945 102.020 21.985 ;
        RECT 97.790 19.605 101.790 19.775 ;
        RECT 102.420 19.265 102.590 22.665 ;
        RECT 103.220 22.155 107.220 22.325 ;
        RECT 102.990 19.945 103.160 21.985 ;
        RECT 107.280 19.945 107.450 21.985 ;
        RECT 107.850 20.240 108.020 22.665 ;
        RECT 108.290 22.670 110.040 22.840 ;
        RECT 108.290 20.270 108.460 22.670 ;
        RECT 109.000 22.160 109.330 22.330 ;
        RECT 108.860 20.950 109.030 21.990 ;
        RECT 109.300 20.950 109.470 21.990 ;
        RECT 109.000 20.610 109.330 20.780 ;
        RECT 109.870 20.270 110.040 22.670 ;
        RECT 108.290 20.240 110.040 20.270 ;
        RECT 110.315 22.675 112.065 22.845 ;
        RECT 110.315 20.240 110.485 22.675 ;
        RECT 111.025 22.165 111.355 22.335 ;
        RECT 103.220 19.605 107.220 19.775 ;
        RECT 107.850 19.275 110.485 20.240 ;
        RECT 110.885 19.955 111.055 21.995 ;
        RECT 111.325 19.955 111.495 21.995 ;
        RECT 111.025 19.615 111.355 19.785 ;
        RECT 111.895 19.275 112.065 22.675 ;
        RECT 107.850 19.265 112.065 19.275 ;
        RECT 86.130 19.245 112.065 19.265 ;
        RECT 114.130 22.665 136.020 22.835 ;
        RECT 114.130 19.265 114.300 22.665 ;
        RECT 114.930 22.155 118.930 22.325 ;
        RECT 114.700 19.945 114.870 21.985 ;
        RECT 118.990 19.945 119.160 21.985 ;
        RECT 114.930 19.605 118.930 19.775 ;
        RECT 119.560 19.265 119.730 22.665 ;
        RECT 120.360 22.155 124.360 22.325 ;
        RECT 120.130 19.945 120.300 21.985 ;
        RECT 124.420 19.945 124.590 21.985 ;
        RECT 120.360 19.605 124.360 19.775 ;
        RECT 124.990 19.265 125.160 22.665 ;
        RECT 125.790 22.155 129.790 22.325 ;
        RECT 125.560 19.945 125.730 21.985 ;
        RECT 129.850 19.945 130.020 21.985 ;
        RECT 125.790 19.605 129.790 19.775 ;
        RECT 130.420 19.265 130.590 22.665 ;
        RECT 131.220 22.155 135.220 22.325 ;
        RECT 130.990 19.945 131.160 21.985 ;
        RECT 135.280 19.945 135.450 21.985 ;
        RECT 135.850 20.240 136.020 22.665 ;
        RECT 136.290 22.670 138.040 22.840 ;
        RECT 136.290 20.270 136.460 22.670 ;
        RECT 137.000 22.160 137.330 22.330 ;
        RECT 136.860 20.950 137.030 21.990 ;
        RECT 137.300 20.950 137.470 21.990 ;
        RECT 137.000 20.610 137.330 20.780 ;
        RECT 137.870 20.270 138.040 22.670 ;
        RECT 136.290 20.240 138.040 20.270 ;
        RECT 138.315 22.675 140.065 22.845 ;
        RECT 138.315 20.240 138.485 22.675 ;
        RECT 139.025 22.165 139.355 22.335 ;
        RECT 131.220 19.605 135.220 19.775 ;
        RECT 135.850 19.275 138.485 20.240 ;
        RECT 138.885 19.955 139.055 21.995 ;
        RECT 139.325 19.955 139.495 21.995 ;
        RECT 139.025 19.615 139.355 19.785 ;
        RECT 139.895 19.275 140.065 22.675 ;
        RECT 135.850 19.265 140.065 19.275 ;
        RECT 114.130 19.245 140.065 19.265 ;
        RECT 1.475 19.105 28.065 19.245 ;
        RECT 29.475 19.105 56.065 19.245 ;
        RECT 57.475 19.105 84.065 19.245 ;
        RECT 85.475 19.105 112.065 19.245 ;
        RECT 113.475 19.105 140.065 19.245 ;
        RECT 1.475 18.380 28.055 19.105 ;
        RECT 29.475 18.380 56.055 19.105 ;
        RECT 57.475 18.380 84.055 19.105 ;
        RECT 85.475 18.380 112.055 19.105 ;
        RECT 113.475 18.380 140.055 19.105 ;
        RECT 1.450 17.480 27.925 17.960 ;
        RECT 29.450 17.480 55.925 17.960 ;
        RECT 57.450 17.480 83.925 17.960 ;
        RECT 85.450 17.480 111.925 17.960 ;
        RECT 113.450 17.480 139.925 17.960 ;
        RECT 1.435 17.420 27.925 17.480 ;
        RECT 29.435 17.420 55.925 17.480 ;
        RECT 57.435 17.420 83.925 17.480 ;
        RECT 85.435 17.420 111.925 17.480 ;
        RECT 113.435 17.420 139.925 17.480 ;
        RECT 1.435 17.260 27.980 17.420 ;
        RECT 1.435 17.235 14.180 17.260 ;
        RECT 1.435 17.005 5.760 17.235 ;
        RECT 1.470 7.745 1.640 17.005 ;
        RECT 2.365 16.435 4.405 16.605 ;
        RECT 1.980 8.375 2.150 16.375 ;
        RECT 4.620 8.375 4.790 16.375 ;
        RECT 2.365 8.145 4.405 8.315 ;
        RECT 5.130 7.745 5.300 17.005 ;
        RECT 1.470 7.575 5.300 7.745 ;
        RECT 5.590 7.745 5.760 17.005 ;
        RECT 6.390 16.725 8.390 16.895 ;
        RECT 6.160 8.470 6.330 16.510 ;
        RECT 8.450 8.470 8.620 16.510 ;
        RECT 6.390 8.085 8.390 8.255 ;
        RECT 9.020 7.745 9.190 17.235 ;
        RECT 9.820 16.725 11.820 16.895 ;
        RECT 9.590 8.470 9.760 16.510 ;
        RECT 11.880 8.470 12.050 16.510 ;
        RECT 12.450 15.665 14.180 17.235 ;
        RECT 26.230 17.250 27.980 17.260 ;
        RECT 12.450 15.495 20.915 15.665 ;
        RECT 12.450 14.085 14.255 15.495 ;
        RECT 14.595 14.625 14.765 14.955 ;
        RECT 14.980 14.925 20.020 15.095 ;
        RECT 14.980 14.485 20.020 14.655 ;
        RECT 20.235 14.625 20.405 14.955 ;
        RECT 20.745 14.085 20.915 15.495 ;
        RECT 12.450 13.915 20.915 14.085 ;
        RECT 12.450 13.400 14.180 13.915 ;
        RECT 12.450 13.285 23.930 13.400 ;
        RECT 9.820 8.085 11.820 8.255 ;
        RECT 12.450 7.745 12.620 13.285 ;
        RECT 5.590 7.575 12.620 7.745 ;
        RECT 12.900 13.230 23.930 13.285 ;
        RECT 12.900 7.740 13.070 13.230 ;
        RECT 13.700 12.720 17.700 12.890 ;
        RECT 13.470 8.465 13.640 12.505 ;
        RECT 17.760 8.465 17.930 12.505 ;
        RECT 13.700 8.080 17.700 8.250 ;
        RECT 18.330 7.740 18.500 13.230 ;
        RECT 19.130 12.720 23.130 12.890 ;
        RECT 18.900 8.465 19.070 12.505 ;
        RECT 23.190 8.465 23.360 12.505 ;
        RECT 19.130 8.080 23.130 8.250 ;
        RECT 23.760 7.740 23.930 13.230 ;
        RECT 12.900 7.570 23.930 7.740 ;
        RECT 24.205 13.245 25.955 13.415 ;
        RECT 24.205 7.755 24.375 13.245 ;
        RECT 24.915 12.735 25.245 12.905 ;
        RECT 24.775 8.480 24.945 12.520 ;
        RECT 25.215 8.480 25.385 12.520 ;
        RECT 24.915 8.095 25.245 8.265 ;
        RECT 25.785 7.755 25.955 13.245 ;
        RECT 24.205 7.585 25.955 7.755 ;
        RECT 26.230 7.760 26.400 17.250 ;
        RECT 26.940 16.740 27.270 16.910 ;
        RECT 26.800 8.485 26.970 16.525 ;
        RECT 27.240 8.485 27.410 16.525 ;
        RECT 26.940 8.100 27.270 8.270 ;
        RECT 27.810 7.760 27.980 17.250 ;
        RECT 29.435 17.260 55.980 17.420 ;
        RECT 29.435 17.235 42.180 17.260 ;
        RECT 29.435 17.005 33.760 17.235 ;
        RECT 26.230 7.590 27.980 7.760 ;
        RECT 29.470 7.745 29.640 17.005 ;
        RECT 30.365 16.435 32.405 16.605 ;
        RECT 29.980 8.375 30.150 16.375 ;
        RECT 32.620 8.375 32.790 16.375 ;
        RECT 30.365 8.145 32.405 8.315 ;
        RECT 33.130 7.745 33.300 17.005 ;
        RECT 29.470 7.575 33.300 7.745 ;
        RECT 33.590 7.745 33.760 17.005 ;
        RECT 34.390 16.725 36.390 16.895 ;
        RECT 34.160 8.470 34.330 16.510 ;
        RECT 36.450 8.470 36.620 16.510 ;
        RECT 34.390 8.085 36.390 8.255 ;
        RECT 37.020 7.745 37.190 17.235 ;
        RECT 37.820 16.725 39.820 16.895 ;
        RECT 37.590 8.470 37.760 16.510 ;
        RECT 39.880 8.470 40.050 16.510 ;
        RECT 40.450 15.665 42.180 17.235 ;
        RECT 54.230 17.250 55.980 17.260 ;
        RECT 40.450 15.495 48.915 15.665 ;
        RECT 40.450 14.085 42.255 15.495 ;
        RECT 42.595 14.625 42.765 14.955 ;
        RECT 42.980 14.925 48.020 15.095 ;
        RECT 42.980 14.485 48.020 14.655 ;
        RECT 48.235 14.625 48.405 14.955 ;
        RECT 48.745 14.085 48.915 15.495 ;
        RECT 40.450 13.915 48.915 14.085 ;
        RECT 40.450 13.400 42.180 13.915 ;
        RECT 40.450 13.285 51.930 13.400 ;
        RECT 37.820 8.085 39.820 8.255 ;
        RECT 40.450 7.745 40.620 13.285 ;
        RECT 33.590 7.575 40.620 7.745 ;
        RECT 40.900 13.230 51.930 13.285 ;
        RECT 40.900 7.740 41.070 13.230 ;
        RECT 41.700 12.720 45.700 12.890 ;
        RECT 41.470 8.465 41.640 12.505 ;
        RECT 45.760 8.465 45.930 12.505 ;
        RECT 41.700 8.080 45.700 8.250 ;
        RECT 46.330 7.740 46.500 13.230 ;
        RECT 47.130 12.720 51.130 12.890 ;
        RECT 46.900 8.465 47.070 12.505 ;
        RECT 51.190 8.465 51.360 12.505 ;
        RECT 47.130 8.080 51.130 8.250 ;
        RECT 51.760 7.740 51.930 13.230 ;
        RECT 40.900 7.570 51.930 7.740 ;
        RECT 52.205 13.245 53.955 13.415 ;
        RECT 52.205 7.755 52.375 13.245 ;
        RECT 52.915 12.735 53.245 12.905 ;
        RECT 52.775 8.480 52.945 12.520 ;
        RECT 53.215 8.480 53.385 12.520 ;
        RECT 52.915 8.095 53.245 8.265 ;
        RECT 53.785 7.755 53.955 13.245 ;
        RECT 52.205 7.585 53.955 7.755 ;
        RECT 54.230 7.760 54.400 17.250 ;
        RECT 54.940 16.740 55.270 16.910 ;
        RECT 54.800 8.485 54.970 16.525 ;
        RECT 55.240 8.485 55.410 16.525 ;
        RECT 54.940 8.100 55.270 8.270 ;
        RECT 55.810 7.760 55.980 17.250 ;
        RECT 57.435 17.260 83.980 17.420 ;
        RECT 57.435 17.235 70.180 17.260 ;
        RECT 57.435 17.005 61.760 17.235 ;
        RECT 54.230 7.590 55.980 7.760 ;
        RECT 57.470 7.745 57.640 17.005 ;
        RECT 58.365 16.435 60.405 16.605 ;
        RECT 57.980 8.375 58.150 16.375 ;
        RECT 60.620 8.375 60.790 16.375 ;
        RECT 58.365 8.145 60.405 8.315 ;
        RECT 61.130 7.745 61.300 17.005 ;
        RECT 57.470 7.575 61.300 7.745 ;
        RECT 61.590 7.745 61.760 17.005 ;
        RECT 62.390 16.725 64.390 16.895 ;
        RECT 62.160 8.470 62.330 16.510 ;
        RECT 64.450 8.470 64.620 16.510 ;
        RECT 62.390 8.085 64.390 8.255 ;
        RECT 65.020 7.745 65.190 17.235 ;
        RECT 65.820 16.725 67.820 16.895 ;
        RECT 65.590 8.470 65.760 16.510 ;
        RECT 67.880 8.470 68.050 16.510 ;
        RECT 68.450 15.665 70.180 17.235 ;
        RECT 82.230 17.250 83.980 17.260 ;
        RECT 68.450 15.495 76.915 15.665 ;
        RECT 68.450 14.085 70.255 15.495 ;
        RECT 70.595 14.625 70.765 14.955 ;
        RECT 70.980 14.925 76.020 15.095 ;
        RECT 70.980 14.485 76.020 14.655 ;
        RECT 76.235 14.625 76.405 14.955 ;
        RECT 76.745 14.085 76.915 15.495 ;
        RECT 68.450 13.915 76.915 14.085 ;
        RECT 68.450 13.400 70.180 13.915 ;
        RECT 68.450 13.285 79.930 13.400 ;
        RECT 65.820 8.085 67.820 8.255 ;
        RECT 68.450 7.745 68.620 13.285 ;
        RECT 61.590 7.575 68.620 7.745 ;
        RECT 68.900 13.230 79.930 13.285 ;
        RECT 68.900 7.740 69.070 13.230 ;
        RECT 69.700 12.720 73.700 12.890 ;
        RECT 69.470 8.465 69.640 12.505 ;
        RECT 73.760 8.465 73.930 12.505 ;
        RECT 69.700 8.080 73.700 8.250 ;
        RECT 74.330 7.740 74.500 13.230 ;
        RECT 75.130 12.720 79.130 12.890 ;
        RECT 74.900 8.465 75.070 12.505 ;
        RECT 79.190 8.465 79.360 12.505 ;
        RECT 75.130 8.080 79.130 8.250 ;
        RECT 79.760 7.740 79.930 13.230 ;
        RECT 68.900 7.570 79.930 7.740 ;
        RECT 80.205 13.245 81.955 13.415 ;
        RECT 80.205 7.755 80.375 13.245 ;
        RECT 80.915 12.735 81.245 12.905 ;
        RECT 80.775 8.480 80.945 12.520 ;
        RECT 81.215 8.480 81.385 12.520 ;
        RECT 80.915 8.095 81.245 8.265 ;
        RECT 81.785 7.755 81.955 13.245 ;
        RECT 80.205 7.585 81.955 7.755 ;
        RECT 82.230 7.760 82.400 17.250 ;
        RECT 82.940 16.740 83.270 16.910 ;
        RECT 82.800 8.485 82.970 16.525 ;
        RECT 83.240 8.485 83.410 16.525 ;
        RECT 82.940 8.100 83.270 8.270 ;
        RECT 83.810 7.760 83.980 17.250 ;
        RECT 85.435 17.260 111.980 17.420 ;
        RECT 85.435 17.235 98.180 17.260 ;
        RECT 85.435 17.005 89.760 17.235 ;
        RECT 82.230 7.590 83.980 7.760 ;
        RECT 85.470 7.745 85.640 17.005 ;
        RECT 86.365 16.435 88.405 16.605 ;
        RECT 85.980 8.375 86.150 16.375 ;
        RECT 88.620 8.375 88.790 16.375 ;
        RECT 86.365 8.145 88.405 8.315 ;
        RECT 89.130 7.745 89.300 17.005 ;
        RECT 85.470 7.575 89.300 7.745 ;
        RECT 89.590 7.745 89.760 17.005 ;
        RECT 90.390 16.725 92.390 16.895 ;
        RECT 90.160 8.470 90.330 16.510 ;
        RECT 92.450 8.470 92.620 16.510 ;
        RECT 90.390 8.085 92.390 8.255 ;
        RECT 93.020 7.745 93.190 17.235 ;
        RECT 93.820 16.725 95.820 16.895 ;
        RECT 93.590 8.470 93.760 16.510 ;
        RECT 95.880 8.470 96.050 16.510 ;
        RECT 96.450 15.665 98.180 17.235 ;
        RECT 110.230 17.250 111.980 17.260 ;
        RECT 96.450 15.495 104.915 15.665 ;
        RECT 96.450 14.085 98.255 15.495 ;
        RECT 98.595 14.625 98.765 14.955 ;
        RECT 98.980 14.925 104.020 15.095 ;
        RECT 98.980 14.485 104.020 14.655 ;
        RECT 104.235 14.625 104.405 14.955 ;
        RECT 104.745 14.085 104.915 15.495 ;
        RECT 96.450 13.915 104.915 14.085 ;
        RECT 96.450 13.400 98.180 13.915 ;
        RECT 96.450 13.285 107.930 13.400 ;
        RECT 93.820 8.085 95.820 8.255 ;
        RECT 96.450 7.745 96.620 13.285 ;
        RECT 89.590 7.575 96.620 7.745 ;
        RECT 96.900 13.230 107.930 13.285 ;
        RECT 96.900 7.740 97.070 13.230 ;
        RECT 97.700 12.720 101.700 12.890 ;
        RECT 97.470 8.465 97.640 12.505 ;
        RECT 101.760 8.465 101.930 12.505 ;
        RECT 97.700 8.080 101.700 8.250 ;
        RECT 102.330 7.740 102.500 13.230 ;
        RECT 103.130 12.720 107.130 12.890 ;
        RECT 102.900 8.465 103.070 12.505 ;
        RECT 107.190 8.465 107.360 12.505 ;
        RECT 103.130 8.080 107.130 8.250 ;
        RECT 107.760 7.740 107.930 13.230 ;
        RECT 96.900 7.570 107.930 7.740 ;
        RECT 108.205 13.245 109.955 13.415 ;
        RECT 108.205 7.755 108.375 13.245 ;
        RECT 108.915 12.735 109.245 12.905 ;
        RECT 108.775 8.480 108.945 12.520 ;
        RECT 109.215 8.480 109.385 12.520 ;
        RECT 108.915 8.095 109.245 8.265 ;
        RECT 109.785 7.755 109.955 13.245 ;
        RECT 108.205 7.585 109.955 7.755 ;
        RECT 110.230 7.760 110.400 17.250 ;
        RECT 110.940 16.740 111.270 16.910 ;
        RECT 110.800 8.485 110.970 16.525 ;
        RECT 111.240 8.485 111.410 16.525 ;
        RECT 110.940 8.100 111.270 8.270 ;
        RECT 111.810 7.760 111.980 17.250 ;
        RECT 113.435 17.260 139.980 17.420 ;
        RECT 113.435 17.235 126.180 17.260 ;
        RECT 113.435 17.005 117.760 17.235 ;
        RECT 110.230 7.590 111.980 7.760 ;
        RECT 113.470 7.745 113.640 17.005 ;
        RECT 114.365 16.435 116.405 16.605 ;
        RECT 113.980 8.375 114.150 16.375 ;
        RECT 116.620 8.375 116.790 16.375 ;
        RECT 114.365 8.145 116.405 8.315 ;
        RECT 117.130 7.745 117.300 17.005 ;
        RECT 113.470 7.575 117.300 7.745 ;
        RECT 117.590 7.745 117.760 17.005 ;
        RECT 118.390 16.725 120.390 16.895 ;
        RECT 118.160 8.470 118.330 16.510 ;
        RECT 120.450 8.470 120.620 16.510 ;
        RECT 118.390 8.085 120.390 8.255 ;
        RECT 121.020 7.745 121.190 17.235 ;
        RECT 121.820 16.725 123.820 16.895 ;
        RECT 121.590 8.470 121.760 16.510 ;
        RECT 123.880 8.470 124.050 16.510 ;
        RECT 124.450 15.665 126.180 17.235 ;
        RECT 138.230 17.250 139.980 17.260 ;
        RECT 124.450 15.495 132.915 15.665 ;
        RECT 124.450 14.085 126.255 15.495 ;
        RECT 126.595 14.625 126.765 14.955 ;
        RECT 126.980 14.925 132.020 15.095 ;
        RECT 126.980 14.485 132.020 14.655 ;
        RECT 132.235 14.625 132.405 14.955 ;
        RECT 132.745 14.085 132.915 15.495 ;
        RECT 124.450 13.915 132.915 14.085 ;
        RECT 124.450 13.400 126.180 13.915 ;
        RECT 124.450 13.285 135.930 13.400 ;
        RECT 121.820 8.085 123.820 8.255 ;
        RECT 124.450 7.745 124.620 13.285 ;
        RECT 117.590 7.575 124.620 7.745 ;
        RECT 124.900 13.230 135.930 13.285 ;
        RECT 124.900 7.740 125.070 13.230 ;
        RECT 125.700 12.720 129.700 12.890 ;
        RECT 125.470 8.465 125.640 12.505 ;
        RECT 129.760 8.465 129.930 12.505 ;
        RECT 125.700 8.080 129.700 8.250 ;
        RECT 130.330 7.740 130.500 13.230 ;
        RECT 131.130 12.720 135.130 12.890 ;
        RECT 130.900 8.465 131.070 12.505 ;
        RECT 135.190 8.465 135.360 12.505 ;
        RECT 131.130 8.080 135.130 8.250 ;
        RECT 135.760 7.740 135.930 13.230 ;
        RECT 124.900 7.570 135.930 7.740 ;
        RECT 136.205 13.245 137.955 13.415 ;
        RECT 136.205 7.755 136.375 13.245 ;
        RECT 136.915 12.735 137.245 12.905 ;
        RECT 136.775 8.480 136.945 12.520 ;
        RECT 137.215 8.480 137.385 12.520 ;
        RECT 136.915 8.095 137.245 8.265 ;
        RECT 137.785 7.755 137.955 13.245 ;
        RECT 136.205 7.585 137.955 7.755 ;
        RECT 138.230 7.760 138.400 17.250 ;
        RECT 138.940 16.740 139.270 16.910 ;
        RECT 138.800 8.485 138.970 16.525 ;
        RECT 139.240 8.485 139.410 16.525 ;
        RECT 138.940 8.100 139.270 8.270 ;
        RECT 139.810 7.760 139.980 17.250 ;
        RECT 138.230 7.590 139.980 7.760 ;
        RECT 2.130 6.665 24.020 6.835 ;
        RECT 2.130 3.265 2.300 6.665 ;
        RECT 2.930 6.155 6.930 6.325 ;
        RECT 2.700 3.945 2.870 5.985 ;
        RECT 6.990 3.945 7.160 5.985 ;
        RECT 2.930 3.605 6.930 3.775 ;
        RECT 7.560 3.265 7.730 6.665 ;
        RECT 8.360 6.155 12.360 6.325 ;
        RECT 8.130 3.945 8.300 5.985 ;
        RECT 12.420 3.945 12.590 5.985 ;
        RECT 8.360 3.605 12.360 3.775 ;
        RECT 12.990 3.265 13.160 6.665 ;
        RECT 13.790 6.155 17.790 6.325 ;
        RECT 13.560 3.945 13.730 5.985 ;
        RECT 17.850 3.945 18.020 5.985 ;
        RECT 13.790 3.605 17.790 3.775 ;
        RECT 18.420 3.265 18.590 6.665 ;
        RECT 19.220 6.155 23.220 6.325 ;
        RECT 18.990 3.945 19.160 5.985 ;
        RECT 23.280 3.945 23.450 5.985 ;
        RECT 23.850 4.240 24.020 6.665 ;
        RECT 24.290 6.670 26.040 6.840 ;
        RECT 24.290 4.270 24.460 6.670 ;
        RECT 25.000 6.160 25.330 6.330 ;
        RECT 24.860 4.950 25.030 5.990 ;
        RECT 25.300 4.950 25.470 5.990 ;
        RECT 25.000 4.610 25.330 4.780 ;
        RECT 25.870 4.270 26.040 6.670 ;
        RECT 24.290 4.240 26.040 4.270 ;
        RECT 26.315 6.675 28.065 6.845 ;
        RECT 26.315 4.240 26.485 6.675 ;
        RECT 27.025 6.165 27.355 6.335 ;
        RECT 19.220 3.605 23.220 3.775 ;
        RECT 23.850 3.275 26.485 4.240 ;
        RECT 26.885 3.955 27.055 5.995 ;
        RECT 27.325 3.955 27.495 5.995 ;
        RECT 27.025 3.615 27.355 3.785 ;
        RECT 27.895 3.275 28.065 6.675 ;
        RECT 23.850 3.265 28.065 3.275 ;
        RECT 2.130 3.245 28.065 3.265 ;
        RECT 30.130 6.665 52.020 6.835 ;
        RECT 30.130 3.265 30.300 6.665 ;
        RECT 30.930 6.155 34.930 6.325 ;
        RECT 30.700 3.945 30.870 5.985 ;
        RECT 34.990 3.945 35.160 5.985 ;
        RECT 30.930 3.605 34.930 3.775 ;
        RECT 35.560 3.265 35.730 6.665 ;
        RECT 36.360 6.155 40.360 6.325 ;
        RECT 36.130 3.945 36.300 5.985 ;
        RECT 40.420 3.945 40.590 5.985 ;
        RECT 36.360 3.605 40.360 3.775 ;
        RECT 40.990 3.265 41.160 6.665 ;
        RECT 41.790 6.155 45.790 6.325 ;
        RECT 41.560 3.945 41.730 5.985 ;
        RECT 45.850 3.945 46.020 5.985 ;
        RECT 41.790 3.605 45.790 3.775 ;
        RECT 46.420 3.265 46.590 6.665 ;
        RECT 47.220 6.155 51.220 6.325 ;
        RECT 46.990 3.945 47.160 5.985 ;
        RECT 51.280 3.945 51.450 5.985 ;
        RECT 51.850 4.240 52.020 6.665 ;
        RECT 52.290 6.670 54.040 6.840 ;
        RECT 52.290 4.270 52.460 6.670 ;
        RECT 53.000 6.160 53.330 6.330 ;
        RECT 52.860 4.950 53.030 5.990 ;
        RECT 53.300 4.950 53.470 5.990 ;
        RECT 53.000 4.610 53.330 4.780 ;
        RECT 53.870 4.270 54.040 6.670 ;
        RECT 52.290 4.240 54.040 4.270 ;
        RECT 54.315 6.675 56.065 6.845 ;
        RECT 54.315 4.240 54.485 6.675 ;
        RECT 55.025 6.165 55.355 6.335 ;
        RECT 47.220 3.605 51.220 3.775 ;
        RECT 51.850 3.275 54.485 4.240 ;
        RECT 54.885 3.955 55.055 5.995 ;
        RECT 55.325 3.955 55.495 5.995 ;
        RECT 55.025 3.615 55.355 3.785 ;
        RECT 55.895 3.275 56.065 6.675 ;
        RECT 51.850 3.265 56.065 3.275 ;
        RECT 30.130 3.245 56.065 3.265 ;
        RECT 58.130 6.665 80.020 6.835 ;
        RECT 58.130 3.265 58.300 6.665 ;
        RECT 58.930 6.155 62.930 6.325 ;
        RECT 58.700 3.945 58.870 5.985 ;
        RECT 62.990 3.945 63.160 5.985 ;
        RECT 58.930 3.605 62.930 3.775 ;
        RECT 63.560 3.265 63.730 6.665 ;
        RECT 64.360 6.155 68.360 6.325 ;
        RECT 64.130 3.945 64.300 5.985 ;
        RECT 68.420 3.945 68.590 5.985 ;
        RECT 64.360 3.605 68.360 3.775 ;
        RECT 68.990 3.265 69.160 6.665 ;
        RECT 69.790 6.155 73.790 6.325 ;
        RECT 69.560 3.945 69.730 5.985 ;
        RECT 73.850 3.945 74.020 5.985 ;
        RECT 69.790 3.605 73.790 3.775 ;
        RECT 74.420 3.265 74.590 6.665 ;
        RECT 75.220 6.155 79.220 6.325 ;
        RECT 74.990 3.945 75.160 5.985 ;
        RECT 79.280 3.945 79.450 5.985 ;
        RECT 79.850 4.240 80.020 6.665 ;
        RECT 80.290 6.670 82.040 6.840 ;
        RECT 80.290 4.270 80.460 6.670 ;
        RECT 81.000 6.160 81.330 6.330 ;
        RECT 80.860 4.950 81.030 5.990 ;
        RECT 81.300 4.950 81.470 5.990 ;
        RECT 81.000 4.610 81.330 4.780 ;
        RECT 81.870 4.270 82.040 6.670 ;
        RECT 80.290 4.240 82.040 4.270 ;
        RECT 82.315 6.675 84.065 6.845 ;
        RECT 82.315 4.240 82.485 6.675 ;
        RECT 83.025 6.165 83.355 6.335 ;
        RECT 75.220 3.605 79.220 3.775 ;
        RECT 79.850 3.275 82.485 4.240 ;
        RECT 82.885 3.955 83.055 5.995 ;
        RECT 83.325 3.955 83.495 5.995 ;
        RECT 83.025 3.615 83.355 3.785 ;
        RECT 83.895 3.275 84.065 6.675 ;
        RECT 79.850 3.265 84.065 3.275 ;
        RECT 58.130 3.245 84.065 3.265 ;
        RECT 86.130 6.665 108.020 6.835 ;
        RECT 86.130 3.265 86.300 6.665 ;
        RECT 86.930 6.155 90.930 6.325 ;
        RECT 86.700 3.945 86.870 5.985 ;
        RECT 90.990 3.945 91.160 5.985 ;
        RECT 86.930 3.605 90.930 3.775 ;
        RECT 91.560 3.265 91.730 6.665 ;
        RECT 92.360 6.155 96.360 6.325 ;
        RECT 92.130 3.945 92.300 5.985 ;
        RECT 96.420 3.945 96.590 5.985 ;
        RECT 92.360 3.605 96.360 3.775 ;
        RECT 96.990 3.265 97.160 6.665 ;
        RECT 97.790 6.155 101.790 6.325 ;
        RECT 97.560 3.945 97.730 5.985 ;
        RECT 101.850 3.945 102.020 5.985 ;
        RECT 97.790 3.605 101.790 3.775 ;
        RECT 102.420 3.265 102.590 6.665 ;
        RECT 103.220 6.155 107.220 6.325 ;
        RECT 102.990 3.945 103.160 5.985 ;
        RECT 107.280 3.945 107.450 5.985 ;
        RECT 107.850 4.240 108.020 6.665 ;
        RECT 108.290 6.670 110.040 6.840 ;
        RECT 108.290 4.270 108.460 6.670 ;
        RECT 109.000 6.160 109.330 6.330 ;
        RECT 108.860 4.950 109.030 5.990 ;
        RECT 109.300 4.950 109.470 5.990 ;
        RECT 109.000 4.610 109.330 4.780 ;
        RECT 109.870 4.270 110.040 6.670 ;
        RECT 108.290 4.240 110.040 4.270 ;
        RECT 110.315 6.675 112.065 6.845 ;
        RECT 110.315 4.240 110.485 6.675 ;
        RECT 111.025 6.165 111.355 6.335 ;
        RECT 103.220 3.605 107.220 3.775 ;
        RECT 107.850 3.275 110.485 4.240 ;
        RECT 110.885 3.955 111.055 5.995 ;
        RECT 111.325 3.955 111.495 5.995 ;
        RECT 111.025 3.615 111.355 3.785 ;
        RECT 111.895 3.275 112.065 6.675 ;
        RECT 107.850 3.265 112.065 3.275 ;
        RECT 86.130 3.245 112.065 3.265 ;
        RECT 114.130 6.665 136.020 6.835 ;
        RECT 114.130 3.265 114.300 6.665 ;
        RECT 114.930 6.155 118.930 6.325 ;
        RECT 114.700 3.945 114.870 5.985 ;
        RECT 118.990 3.945 119.160 5.985 ;
        RECT 114.930 3.605 118.930 3.775 ;
        RECT 119.560 3.265 119.730 6.665 ;
        RECT 120.360 6.155 124.360 6.325 ;
        RECT 120.130 3.945 120.300 5.985 ;
        RECT 124.420 3.945 124.590 5.985 ;
        RECT 120.360 3.605 124.360 3.775 ;
        RECT 124.990 3.265 125.160 6.665 ;
        RECT 125.790 6.155 129.790 6.325 ;
        RECT 125.560 3.945 125.730 5.985 ;
        RECT 129.850 3.945 130.020 5.985 ;
        RECT 125.790 3.605 129.790 3.775 ;
        RECT 130.420 3.265 130.590 6.665 ;
        RECT 131.220 6.155 135.220 6.325 ;
        RECT 130.990 3.945 131.160 5.985 ;
        RECT 135.280 3.945 135.450 5.985 ;
        RECT 135.850 4.240 136.020 6.665 ;
        RECT 136.290 6.670 138.040 6.840 ;
        RECT 136.290 4.270 136.460 6.670 ;
        RECT 137.000 6.160 137.330 6.330 ;
        RECT 136.860 4.950 137.030 5.990 ;
        RECT 137.300 4.950 137.470 5.990 ;
        RECT 137.000 4.610 137.330 4.780 ;
        RECT 137.870 4.270 138.040 6.670 ;
        RECT 136.290 4.240 138.040 4.270 ;
        RECT 138.315 6.675 140.065 6.845 ;
        RECT 138.315 4.240 138.485 6.675 ;
        RECT 139.025 6.165 139.355 6.335 ;
        RECT 131.220 3.605 135.220 3.775 ;
        RECT 135.850 3.275 138.485 4.240 ;
        RECT 138.885 3.955 139.055 5.995 ;
        RECT 139.325 3.955 139.495 5.995 ;
        RECT 139.025 3.615 139.355 3.785 ;
        RECT 139.895 3.275 140.065 6.675 ;
        RECT 135.850 3.265 140.065 3.275 ;
        RECT 114.130 3.245 140.065 3.265 ;
        RECT 1.475 3.105 28.065 3.245 ;
        RECT 29.475 3.105 56.065 3.245 ;
        RECT 57.475 3.105 84.065 3.245 ;
        RECT 85.475 3.105 112.065 3.245 ;
        RECT 113.475 3.105 140.065 3.245 ;
        RECT 1.475 2.380 28.055 3.105 ;
        RECT 29.475 2.380 56.055 3.105 ;
        RECT 57.475 2.380 84.055 3.105 ;
        RECT 85.475 2.380 112.055 3.105 ;
        RECT 113.475 2.380 140.055 3.105 ;
      LAYER met1 ;
        RECT 10.970 57.310 13.930 57.410 ;
        RECT 2.150 57.280 4.255 57.310 ;
        RECT 2.090 56.720 4.255 57.280 ;
        RECT 4.835 57.280 6.940 57.310 ;
        RECT 8.130 57.280 10.235 57.310 ;
        RECT 4.835 56.720 10.235 57.280 ;
        RECT 10.815 56.720 13.930 57.310 ;
        RECT 2.090 55.490 3.990 56.720 ;
        RECT 4.890 56.680 10.190 56.720 ;
        RECT 10.970 56.630 13.930 56.720 ;
        RECT 2.090 54.900 4.255 55.490 ;
        RECT 4.835 55.480 6.940 55.490 ;
        RECT 8.130 55.480 10.235 55.490 ;
        RECT 4.835 54.900 10.235 55.480 ;
        RECT 10.815 54.900 12.920 55.490 ;
        RECT 2.090 54.880 3.990 54.900 ;
        RECT 4.890 54.880 10.190 54.900 ;
        RECT 2.290 53.670 4.190 53.680 ;
        RECT 4.890 53.670 10.190 53.680 ;
        RECT 10.890 53.670 12.790 54.900 ;
        RECT 2.150 53.080 4.255 53.670 ;
        RECT 4.835 53.080 10.235 53.670 ;
        RECT 10.815 53.080 12.920 53.670 ;
        RECT 2.290 51.850 4.190 53.080 ;
        RECT 61.420 52.540 61.630 52.570 ;
        RECT 61.420 52.090 67.670 52.540 ;
        RECT 61.420 52.060 61.630 52.090 ;
        RECT 10.890 51.875 13.215 51.880 ;
        RECT 10.890 51.850 16.180 51.875 ;
        RECT 25.745 51.850 26.120 51.945 ;
        RECT 41.065 51.875 46.190 51.880 ;
        RECT 28.820 51.850 46.190 51.875 ;
        RECT 46.890 51.850 52.190 51.980 ;
        RECT 52.890 51.850 58.190 51.880 ;
        RECT 58.890 51.850 70.290 51.880 ;
        RECT 70.890 51.850 76.190 51.880 ;
        RECT 76.890 51.850 82.190 51.880 ;
        RECT 2.150 51.260 4.255 51.850 ;
        RECT 4.835 51.780 6.940 51.850 ;
        RECT 8.130 51.780 10.235 51.850 ;
        RECT 4.835 51.260 10.235 51.780 ;
        RECT 10.815 51.260 16.215 51.850 ;
        RECT 16.795 51.260 22.195 51.850 ;
        RECT 22.775 51.810 24.880 51.850 ;
        RECT 25.745 51.810 28.175 51.850 ;
        RECT 22.775 51.260 28.175 51.810 ;
        RECT 28.755 51.270 46.275 51.850 ;
        RECT 28.755 51.260 30.860 51.270 ;
        RECT 41.065 51.260 46.275 51.270 ;
        RECT 46.855 51.280 52.255 51.850 ;
        RECT 46.855 51.260 48.960 51.280 ;
        RECT 50.150 51.260 52.255 51.280 ;
        RECT 52.835 51.260 58.235 51.850 ;
        RECT 58.815 51.260 70.290 51.850 ;
        RECT 70.855 51.260 76.255 51.850 ;
        RECT 76.835 51.280 82.235 51.850 ;
        RECT 76.835 51.260 78.940 51.280 ;
        RECT 80.130 51.260 82.235 51.280 ;
        RECT 82.815 51.260 84.920 51.850 ;
        RECT 4.890 51.180 10.190 51.260 ;
        RECT 10.890 51.180 16.180 51.260 ;
        RECT 16.840 51.255 22.160 51.260 ;
        RECT 12.720 51.170 16.180 51.180 ;
        RECT 1.560 50.360 9.985 50.855 ;
        RECT 10.520 50.500 11.025 50.595 ;
        RECT 17.030 50.500 17.285 51.255 ;
        RECT 22.810 51.215 28.130 51.260 ;
        RECT 28.855 50.575 29.260 51.260 ;
        RECT 41.065 51.180 46.190 51.260 ;
        RECT 47.135 50.630 47.510 51.260 ;
        RECT 52.890 51.180 58.190 51.260 ;
        RECT 58.890 51.180 70.290 51.260 ;
        RECT 70.890 51.180 76.190 51.260 ;
        RECT 59.065 50.680 59.470 51.180 ;
        RECT 10.520 50.245 17.285 50.500 ;
        RECT 10.520 50.150 11.025 50.245 ;
        RECT 26.565 50.170 29.260 50.575 ;
        RECT 38.555 50.255 47.510 50.630 ;
        RECT 54.665 50.275 59.470 50.680 ;
        RECT 71.015 50.655 71.365 51.180 ;
        RECT 81.780 50.735 82.120 51.260 ;
        RECT 82.970 51.160 84.910 51.260 ;
        RECT 83.130 50.755 83.525 51.160 ;
        RECT 66.565 50.305 71.365 50.655 ;
        RECT 77.790 50.170 80.360 50.690 ;
        RECT 81.750 50.395 82.150 50.735 ;
        RECT 82.710 50.360 83.525 50.755 ;
        RECT 84.470 51.100 84.910 51.160 ;
        RECT 144.190 51.100 146.190 51.180 ;
        RECT 84.470 50.660 146.190 51.100 ;
        RECT 27.490 49.960 30.190 49.980 ;
        RECT 55.390 49.960 58.090 49.980 ;
        RECT 83.490 49.960 85.790 49.980 ;
        RECT 111.590 49.960 113.890 49.980 ;
        RECT 1.450 49.280 139.925 49.960 ;
        RECT 144.190 49.310 146.190 50.660 ;
        RECT 1.450 49.260 27.925 49.280 ;
        RECT 29.450 49.260 55.925 49.280 ;
        RECT 57.450 49.260 83.925 49.280 ;
        RECT 85.450 49.260 111.925 49.280 ;
        RECT 113.450 49.260 139.925 49.280 ;
        RECT 2.420 48.635 4.330 49.260 ;
        RECT 6.420 48.925 8.305 48.930 ;
        RECT 9.865 48.925 11.750 48.930 ;
        RECT 6.410 48.695 8.370 48.925 ;
        RECT 9.840 48.695 11.800 48.925 ;
        RECT 2.385 48.405 4.385 48.635 ;
        RECT 6.130 48.410 6.360 48.490 ;
        RECT 1.590 48.355 2.085 48.375 ;
        RECT 1.590 45.060 2.180 48.355 ;
        RECT 4.590 48.275 4.820 48.355 ;
        RECT 4.560 45.060 4.820 48.275 ;
        RECT 1.590 43.245 4.820 45.060 ;
        RECT 1.590 40.395 2.180 43.245 ;
        RECT 3.075 40.640 3.335 40.960 ;
        RECT 4.560 40.645 4.820 43.245 ;
        RECT 5.890 40.990 6.360 48.410 ;
        RECT 6.850 41.775 7.740 48.695 ;
        RECT 8.420 48.390 8.650 48.490 ;
        RECT 8.420 48.380 8.775 48.390 ;
        RECT 9.560 48.380 9.790 48.490 ;
        RECT 3.130 40.480 3.280 40.640 ;
        RECT 1.590 35.255 2.085 40.395 ;
        RECT 3.105 40.345 3.310 40.480 ;
        RECT 4.590 40.395 4.820 40.645 ;
        RECT 5.610 40.550 6.360 40.990 ;
        RECT 6.780 40.775 7.795 41.775 ;
        RECT 2.385 40.115 4.385 40.345 ;
        RECT 5.610 38.355 5.980 40.550 ;
        RECT 6.130 40.490 6.360 40.550 ;
        RECT 6.850 40.285 7.740 40.775 ;
        RECT 8.420 40.580 9.790 48.380 ;
        RECT 10.325 43.635 11.215 48.695 ;
        RECT 11.850 48.410 12.080 48.490 ;
        RECT 10.320 42.015 11.220 43.635 ;
        RECT 10.325 41.605 11.215 42.015 ;
        RECT 10.250 40.605 11.280 41.605 ;
        RECT 11.850 40.625 12.225 48.410 ;
        RECT 12.500 48.025 14.180 49.260 ;
        RECT 15.015 48.025 19.940 48.035 ;
        RECT 12.500 47.545 19.940 48.025 ;
        RECT 12.500 45.285 14.180 47.545 ;
        RECT 15.015 47.125 19.940 47.545 ;
        RECT 14.520 46.935 14.775 46.960 ;
        RECT 14.520 46.920 14.795 46.935 ;
        RECT 14.490 46.645 14.825 46.920 ;
        RECT 15.000 46.895 20.000 47.125 ;
        RECT 20.210 46.935 20.465 46.960 ;
        RECT 14.520 46.630 14.775 46.645 ;
        RECT 15.000 46.455 20.000 46.685 ;
        RECT 20.205 46.645 20.465 46.935 ;
        RECT 20.210 46.630 20.465 46.645 ;
        RECT 15.045 46.445 19.900 46.455 ;
        RECT 15.045 44.920 17.690 44.925 ;
        RECT 13.720 44.720 17.690 44.920 ;
        RECT 13.720 44.690 17.680 44.720 ;
        RECT 12.560 44.335 12.895 44.610 ;
        RECT 13.440 44.440 13.670 44.485 ;
        RECT 8.420 40.560 8.775 40.580 ;
        RECT 8.420 40.490 8.650 40.560 ;
        RECT 9.560 40.490 9.790 40.580 ;
        RECT 10.320 40.465 11.230 40.605 ;
        RECT 11.850 40.490 12.240 40.625 ;
        RECT 10.310 40.285 11.320 40.465 ;
        RECT 6.410 40.055 8.370 40.285 ;
        RECT 9.840 40.055 11.800 40.285 ;
        RECT 7.135 39.065 7.465 40.055 ;
        RECT 9.865 40.050 11.750 40.055 ;
        RECT 12.045 38.355 12.240 40.490 ;
        RECT 12.630 38.830 12.820 44.335 ;
        RECT 13.250 43.105 13.670 44.440 ;
        RECT 14.975 43.105 16.320 44.690 ;
        RECT 13.250 41.720 16.320 43.105 ;
        RECT 13.250 40.990 13.670 41.720 ;
        RECT 13.245 40.485 13.670 40.990 ;
        RECT 12.630 38.640 12.945 38.830 ;
        RECT 2.950 38.125 6.910 38.355 ;
        RECT 8.380 38.125 12.340 38.355 ;
        RECT 12.755 38.130 12.945 38.640 ;
        RECT 2.670 37.515 2.900 37.965 ;
        RECT 4.150 37.515 4.940 38.125 ;
        RECT 2.670 37.210 4.940 37.515 ;
        RECT 2.615 37.195 4.940 37.210 ;
        RECT 2.530 36.350 4.940 37.195 ;
        RECT 2.530 35.975 2.900 36.350 ;
        RECT 2.670 35.965 2.900 35.975 ;
        RECT 4.150 35.805 4.940 36.350 ;
        RECT 6.960 37.880 7.190 37.965 ;
        RECT 8.100 37.880 8.330 37.965 ;
        RECT 6.960 36.055 8.330 37.880 ;
        RECT 6.960 35.965 7.190 36.055 ;
        RECT 2.950 35.575 6.910 35.805 ;
        RECT 2.530 35.255 2.755 35.265 ;
        RECT 7.430 35.255 7.920 36.055 ;
        RECT 8.100 35.965 8.330 36.055 ;
        RECT 9.815 37.745 11.155 38.125 ;
        RECT 12.390 37.745 12.620 37.965 ;
        RECT 9.815 36.150 12.620 37.745 ;
        RECT 9.815 35.805 11.155 36.150 ;
        RECT 12.390 35.965 12.620 36.150 ;
        RECT 8.380 35.575 12.340 35.805 ;
        RECT 12.770 35.785 12.945 38.130 ;
        RECT 13.245 37.965 13.540 40.485 ;
        RECT 14.975 40.280 16.320 41.720 ;
        RECT 17.730 44.390 17.960 44.485 ;
        RECT 18.205 44.390 18.695 46.445 ;
        RECT 19.265 44.920 19.900 44.925 ;
        RECT 19.150 44.690 23.110 44.920 ;
        RECT 18.870 44.390 19.100 44.485 ;
        RECT 17.730 40.565 19.100 44.390 ;
        RECT 17.730 40.485 17.960 40.565 ;
        RECT 18.870 40.485 19.100 40.565 ;
        RECT 20.525 40.280 21.870 44.690 ;
        RECT 23.160 44.420 23.390 44.485 ;
        RECT 24.045 44.425 24.520 49.260 ;
        RECT 25.845 48.455 26.525 49.260 ;
        RECT 26.945 48.735 27.280 48.985 ;
        RECT 26.960 48.710 27.250 48.735 ;
        RECT 30.420 48.635 32.330 49.260 ;
        RECT 34.420 48.925 36.305 48.930 ;
        RECT 37.865 48.925 39.750 48.930 ;
        RECT 34.410 48.695 36.370 48.925 ;
        RECT 37.840 48.695 39.800 48.925 ;
        RECT 26.770 48.455 27.000 48.505 ;
        RECT 25.845 47.955 27.000 48.455 ;
        RECT 24.915 44.735 25.250 44.985 ;
        RECT 24.935 44.705 25.225 44.735 ;
        RECT 24.745 44.425 24.975 44.500 ;
        RECT 23.160 40.485 23.615 44.420 ;
        RECT 24.045 43.680 24.975 44.425 ;
        RECT 24.380 40.565 24.975 43.680 ;
        RECT 24.745 40.500 24.975 40.565 ;
        RECT 25.185 44.475 25.415 44.500 ;
        RECT 25.185 40.920 25.695 44.475 ;
        RECT 25.185 40.550 25.880 40.920 ;
        RECT 26.380 40.600 27.000 47.955 ;
        RECT 25.185 40.500 25.415 40.550 ;
        RECT 13.720 40.250 17.680 40.280 ;
        RECT 19.150 40.250 23.110 40.280 ;
        RECT 13.720 40.090 23.110 40.250 ;
        RECT 13.720 40.050 17.680 40.090 ;
        RECT 19.150 40.050 23.110 40.090 ;
        RECT 23.275 38.660 23.615 40.485 ;
        RECT 24.925 38.660 25.345 40.305 ;
        RECT 23.275 38.505 25.345 38.660 ;
        RECT 23.350 38.390 25.345 38.505 ;
        RECT 13.810 38.125 17.770 38.355 ;
        RECT 19.240 38.125 23.200 38.355 ;
        RECT 13.245 37.205 13.760 37.965 ;
        RECT 13.315 36.025 13.760 37.205 ;
        RECT 13.530 35.965 13.760 36.025 ;
        RECT 15.190 35.805 16.145 38.125 ;
        RECT 17.820 37.900 18.050 37.965 ;
        RECT 18.960 37.900 19.190 37.965 ;
        RECT 17.820 36.030 19.190 37.900 ;
        RECT 17.820 35.965 18.050 36.030 ;
        RECT 12.755 35.255 12.945 35.785 ;
        RECT 13.810 35.575 17.770 35.805 ;
        RECT 18.225 35.255 18.780 36.030 ;
        RECT 18.960 35.965 19.190 36.030 ;
        RECT 20.635 35.805 21.590 38.125 ;
        RECT 23.350 37.970 23.615 38.390 ;
        RECT 24.925 38.115 25.345 38.390 ;
        RECT 25.580 39.355 25.880 40.550 ;
        RECT 26.770 40.505 27.000 40.600 ;
        RECT 27.210 48.430 27.440 48.505 ;
        RECT 27.210 41.110 27.985 48.430 ;
        RECT 30.385 48.405 32.385 48.635 ;
        RECT 34.130 48.410 34.360 48.490 ;
        RECT 29.950 45.060 30.180 48.355 ;
        RECT 32.590 48.275 32.820 48.355 ;
        RECT 32.560 45.060 32.820 48.275 ;
        RECT 29.950 43.245 32.820 45.060 ;
        RECT 27.210 40.580 28.060 41.110 ;
        RECT 29.950 40.825 30.180 43.245 ;
        RECT 27.210 40.505 27.440 40.580 ;
        RECT 26.875 39.825 27.390 40.315 ;
        RECT 27.690 39.825 28.060 40.580 ;
        RECT 29.590 40.395 30.180 40.825 ;
        RECT 31.075 40.640 31.335 40.960 ;
        RECT 32.560 40.645 32.820 43.245 ;
        RECT 33.890 40.990 34.360 48.410 ;
        RECT 34.850 41.775 35.740 48.695 ;
        RECT 36.420 48.390 36.650 48.490 ;
        RECT 36.420 48.380 36.775 48.390 ;
        RECT 37.560 48.380 37.790 48.490 ;
        RECT 31.130 40.480 31.280 40.640 ;
        RECT 26.875 39.360 27.385 39.825 ;
        RECT 26.510 39.355 27.385 39.360 ;
        RECT 25.580 38.950 27.385 39.355 ;
        RECT 25.580 38.110 25.880 38.950 ;
        RECT 26.510 38.935 27.385 38.950 ;
        RECT 26.875 38.825 27.385 38.935 ;
        RECT 26.875 38.125 27.390 38.825 ;
        RECT 27.615 38.795 28.615 39.825 ;
        RECT 23.275 37.965 23.615 37.970 ;
        RECT 23.250 36.020 23.615 37.965 ;
        RECT 24.830 37.900 25.060 37.970 ;
        RECT 24.335 37.230 25.060 37.900 ;
        RECT 24.325 37.040 25.060 37.230 ;
        RECT 24.325 36.240 24.680 37.040 ;
        RECT 24.830 36.970 25.060 37.040 ;
        RECT 25.270 37.925 25.500 37.970 ;
        RECT 25.640 37.925 25.880 38.110 ;
        RECT 25.270 37.595 25.880 37.925 ;
        RECT 26.855 37.870 27.085 37.975 ;
        RECT 25.270 37.040 25.765 37.595 ;
        RECT 25.270 36.970 25.500 37.040 ;
        RECT 25.020 36.785 25.310 36.810 ;
        RECT 25.005 36.535 25.340 36.785 ;
        RECT 26.625 36.765 27.085 37.870 ;
        RECT 26.305 36.240 27.085 36.765 ;
        RECT 23.885 36.060 27.085 36.240 ;
        RECT 23.250 35.965 23.480 36.020 ;
        RECT 19.240 35.575 23.200 35.805 ;
        RECT 23.885 35.620 26.690 36.060 ;
        RECT 26.855 35.975 27.085 36.060 ;
        RECT 27.295 37.910 27.525 37.975 ;
        RECT 27.690 37.910 28.060 38.795 ;
        RECT 27.295 37.585 28.060 37.910 ;
        RECT 27.295 36.045 28.055 37.585 ;
        RECT 27.295 35.975 27.525 36.045 ;
        RECT 27.045 35.795 27.335 35.815 ;
        RECT 23.885 35.255 26.350 35.620 ;
        RECT 27.020 35.545 27.355 35.795 ;
        RECT 29.590 35.280 30.085 40.395 ;
        RECT 31.105 40.345 31.310 40.480 ;
        RECT 32.590 40.395 32.820 40.645 ;
        RECT 33.610 40.550 34.360 40.990 ;
        RECT 34.780 40.775 35.795 41.775 ;
        RECT 30.385 40.115 32.385 40.345 ;
        RECT 33.610 38.355 33.980 40.550 ;
        RECT 34.130 40.490 34.360 40.550 ;
        RECT 34.850 40.285 35.740 40.775 ;
        RECT 36.420 40.580 37.790 48.380 ;
        RECT 38.325 43.635 39.215 48.695 ;
        RECT 39.850 48.410 40.080 48.490 ;
        RECT 38.320 42.015 39.220 43.635 ;
        RECT 38.325 41.605 39.215 42.015 ;
        RECT 38.250 40.605 39.280 41.605 ;
        RECT 39.850 40.625 40.225 48.410 ;
        RECT 40.500 48.025 42.180 49.260 ;
        RECT 43.015 48.025 47.940 48.035 ;
        RECT 40.500 47.545 47.940 48.025 ;
        RECT 40.500 45.285 42.180 47.545 ;
        RECT 43.015 47.125 47.940 47.545 ;
        RECT 42.520 46.935 42.775 46.960 ;
        RECT 42.520 46.920 42.795 46.935 ;
        RECT 42.490 46.645 42.825 46.920 ;
        RECT 43.000 46.895 48.000 47.125 ;
        RECT 48.210 46.935 48.465 46.960 ;
        RECT 42.520 46.630 42.775 46.645 ;
        RECT 43.000 46.455 48.000 46.685 ;
        RECT 48.205 46.645 48.465 46.935 ;
        RECT 48.210 46.630 48.465 46.645 ;
        RECT 43.045 46.445 47.900 46.455 ;
        RECT 43.045 44.920 45.690 44.925 ;
        RECT 41.720 44.720 45.690 44.920 ;
        RECT 41.720 44.690 45.680 44.720 ;
        RECT 40.560 44.335 40.895 44.610 ;
        RECT 41.440 44.440 41.670 44.485 ;
        RECT 36.420 40.560 36.775 40.580 ;
        RECT 36.420 40.490 36.650 40.560 ;
        RECT 37.560 40.490 37.790 40.580 ;
        RECT 38.320 40.465 39.230 40.605 ;
        RECT 39.850 40.490 40.240 40.625 ;
        RECT 38.310 40.285 39.320 40.465 ;
        RECT 34.410 40.055 36.370 40.285 ;
        RECT 37.840 40.055 39.800 40.285 ;
        RECT 35.120 39.340 35.470 40.055 ;
        RECT 37.865 40.050 39.750 40.055 ;
        RECT 40.045 38.355 40.240 40.490 ;
        RECT 40.630 38.830 40.820 44.335 ;
        RECT 41.250 43.105 41.670 44.440 ;
        RECT 42.975 43.105 44.320 44.690 ;
        RECT 41.250 41.720 44.320 43.105 ;
        RECT 41.250 40.990 41.670 41.720 ;
        RECT 41.245 40.485 41.670 40.990 ;
        RECT 40.630 38.640 40.945 38.830 ;
        RECT 30.950 38.125 34.910 38.355 ;
        RECT 36.380 38.125 40.340 38.355 ;
        RECT 40.755 38.130 40.945 38.640 ;
        RECT 30.670 37.515 30.900 37.965 ;
        RECT 32.150 37.515 32.940 38.125 ;
        RECT 30.670 37.210 32.940 37.515 ;
        RECT 30.615 37.195 32.940 37.210 ;
        RECT 30.530 36.350 32.940 37.195 ;
        RECT 30.530 35.975 30.900 36.350 ;
        RECT 30.670 35.965 30.900 35.975 ;
        RECT 32.150 35.805 32.940 36.350 ;
        RECT 34.960 37.880 35.190 37.965 ;
        RECT 36.100 37.880 36.330 37.965 ;
        RECT 34.960 36.055 36.330 37.880 ;
        RECT 34.960 35.965 35.190 36.055 ;
        RECT 30.950 35.575 34.910 35.805 ;
        RECT 27.990 35.255 30.085 35.280 ;
        RECT 30.530 35.255 30.755 35.265 ;
        RECT 35.430 35.255 35.920 36.055 ;
        RECT 36.100 35.965 36.330 36.055 ;
        RECT 37.815 37.745 39.155 38.125 ;
        RECT 40.390 37.745 40.620 37.965 ;
        RECT 37.815 36.150 40.620 37.745 ;
        RECT 37.815 35.805 39.155 36.150 ;
        RECT 40.390 35.965 40.620 36.150 ;
        RECT 36.380 35.575 40.340 35.805 ;
        RECT 40.770 35.785 40.945 38.130 ;
        RECT 41.245 37.965 41.540 40.485 ;
        RECT 42.975 40.280 44.320 41.720 ;
        RECT 45.730 44.390 45.960 44.485 ;
        RECT 46.205 44.390 46.695 46.445 ;
        RECT 47.265 44.920 47.900 44.925 ;
        RECT 47.150 44.690 51.110 44.920 ;
        RECT 46.870 44.390 47.100 44.485 ;
        RECT 45.730 40.565 47.100 44.390 ;
        RECT 45.730 40.485 45.960 40.565 ;
        RECT 46.870 40.485 47.100 40.565 ;
        RECT 48.525 40.280 49.870 44.690 ;
        RECT 51.160 44.420 51.390 44.485 ;
        RECT 52.045 44.425 52.520 49.260 ;
        RECT 53.845 48.455 54.525 49.260 ;
        RECT 54.945 48.735 55.280 48.985 ;
        RECT 54.960 48.710 55.250 48.735 ;
        RECT 58.420 48.635 60.330 49.260 ;
        RECT 62.420 48.925 64.305 48.930 ;
        RECT 65.865 48.925 67.750 48.930 ;
        RECT 62.410 48.695 64.370 48.925 ;
        RECT 65.840 48.695 67.800 48.925 ;
        RECT 54.770 48.455 55.000 48.505 ;
        RECT 53.845 47.955 55.000 48.455 ;
        RECT 52.915 44.735 53.250 44.985 ;
        RECT 52.935 44.705 53.225 44.735 ;
        RECT 52.745 44.425 52.975 44.500 ;
        RECT 51.160 40.485 51.615 44.420 ;
        RECT 52.045 43.680 52.975 44.425 ;
        RECT 52.380 40.565 52.975 43.680 ;
        RECT 52.745 40.500 52.975 40.565 ;
        RECT 53.185 44.475 53.415 44.500 ;
        RECT 53.185 40.920 53.695 44.475 ;
        RECT 53.185 40.550 53.880 40.920 ;
        RECT 54.380 40.600 55.000 47.955 ;
        RECT 53.185 40.500 53.415 40.550 ;
        RECT 41.720 40.250 45.680 40.280 ;
        RECT 47.150 40.250 51.110 40.280 ;
        RECT 41.720 40.090 51.110 40.250 ;
        RECT 41.720 40.050 45.680 40.090 ;
        RECT 47.150 40.050 51.110 40.090 ;
        RECT 51.275 38.660 51.615 40.485 ;
        RECT 52.925 38.660 53.345 40.305 ;
        RECT 51.275 38.505 53.345 38.660 ;
        RECT 51.350 38.390 53.345 38.505 ;
        RECT 41.810 38.125 45.770 38.355 ;
        RECT 47.240 38.125 51.200 38.355 ;
        RECT 41.245 37.205 41.760 37.965 ;
        RECT 41.315 36.025 41.760 37.205 ;
        RECT 41.530 35.965 41.760 36.025 ;
        RECT 43.190 35.805 44.145 38.125 ;
        RECT 45.820 37.900 46.050 37.965 ;
        RECT 46.960 37.900 47.190 37.965 ;
        RECT 45.820 36.030 47.190 37.900 ;
        RECT 45.820 35.965 46.050 36.030 ;
        RECT 40.755 35.255 40.945 35.785 ;
        RECT 41.810 35.575 45.770 35.805 ;
        RECT 46.225 35.255 46.780 36.030 ;
        RECT 46.960 35.965 47.190 36.030 ;
        RECT 48.635 35.805 49.590 38.125 ;
        RECT 51.350 37.970 51.615 38.390 ;
        RECT 52.925 38.115 53.345 38.390 ;
        RECT 53.580 39.355 53.880 40.550 ;
        RECT 54.770 40.505 55.000 40.600 ;
        RECT 55.210 48.430 55.440 48.505 ;
        RECT 55.210 41.110 55.985 48.430 ;
        RECT 58.385 48.405 60.385 48.635 ;
        RECT 62.130 48.410 62.360 48.490 ;
        RECT 57.950 45.060 58.180 48.355 ;
        RECT 60.590 48.275 60.820 48.355 ;
        RECT 60.560 45.060 60.820 48.275 ;
        RECT 57.950 43.245 60.820 45.060 ;
        RECT 55.210 40.580 56.060 41.110 ;
        RECT 57.950 40.825 58.180 43.245 ;
        RECT 55.210 40.505 55.440 40.580 ;
        RECT 54.875 39.825 55.390 40.315 ;
        RECT 54.875 39.360 55.385 39.825 ;
        RECT 55.690 39.795 56.060 40.580 ;
        RECT 57.590 40.395 58.180 40.825 ;
        RECT 59.075 40.640 59.335 40.960 ;
        RECT 60.560 40.645 60.820 43.245 ;
        RECT 61.890 40.990 62.360 48.410 ;
        RECT 62.850 41.775 63.740 48.695 ;
        RECT 64.420 48.390 64.650 48.490 ;
        RECT 64.420 48.380 64.775 48.390 ;
        RECT 65.560 48.380 65.790 48.490 ;
        RECT 59.130 40.480 59.280 40.640 ;
        RECT 54.510 39.355 55.385 39.360 ;
        RECT 53.580 38.950 55.385 39.355 ;
        RECT 53.580 38.110 53.880 38.950 ;
        RECT 54.510 38.935 55.385 38.950 ;
        RECT 54.875 38.825 55.385 38.935 ;
        RECT 54.875 38.125 55.390 38.825 ;
        RECT 55.585 38.795 56.615 39.795 ;
        RECT 51.275 37.965 51.615 37.970 ;
        RECT 51.250 36.020 51.615 37.965 ;
        RECT 52.830 37.900 53.060 37.970 ;
        RECT 52.335 37.230 53.060 37.900 ;
        RECT 52.325 37.040 53.060 37.230 ;
        RECT 52.325 36.240 52.680 37.040 ;
        RECT 52.830 36.970 53.060 37.040 ;
        RECT 53.270 37.925 53.500 37.970 ;
        RECT 53.640 37.925 53.880 38.110 ;
        RECT 53.270 37.595 53.880 37.925 ;
        RECT 54.855 37.870 55.085 37.975 ;
        RECT 53.270 37.040 53.765 37.595 ;
        RECT 53.270 36.970 53.500 37.040 ;
        RECT 53.020 36.785 53.310 36.810 ;
        RECT 53.005 36.535 53.340 36.785 ;
        RECT 54.625 36.765 55.085 37.870 ;
        RECT 54.305 36.240 55.085 36.765 ;
        RECT 51.885 36.060 55.085 36.240 ;
        RECT 51.250 35.965 51.480 36.020 ;
        RECT 47.240 35.575 51.200 35.805 ;
        RECT 51.885 35.620 54.690 36.060 ;
        RECT 54.855 35.975 55.085 36.060 ;
        RECT 55.295 37.910 55.525 37.975 ;
        RECT 55.690 37.910 56.060 38.795 ;
        RECT 55.295 37.585 56.060 37.910 ;
        RECT 55.295 36.045 56.055 37.585 ;
        RECT 55.295 35.975 55.525 36.045 ;
        RECT 55.045 35.795 55.335 35.815 ;
        RECT 51.885 35.255 54.350 35.620 ;
        RECT 55.020 35.545 55.355 35.795 ;
        RECT 57.590 35.280 58.085 40.395 ;
        RECT 59.105 40.345 59.310 40.480 ;
        RECT 60.590 40.395 60.820 40.645 ;
        RECT 61.610 40.550 62.360 40.990 ;
        RECT 62.780 40.775 63.795 41.775 ;
        RECT 58.385 40.115 60.385 40.345 ;
        RECT 61.610 38.355 61.980 40.550 ;
        RECT 62.130 40.490 62.360 40.550 ;
        RECT 62.850 40.285 63.740 40.775 ;
        RECT 64.420 40.580 65.790 48.380 ;
        RECT 66.325 43.635 67.215 48.695 ;
        RECT 67.850 48.410 68.080 48.490 ;
        RECT 66.320 42.015 67.220 43.635 ;
        RECT 66.325 41.605 67.215 42.015 ;
        RECT 66.250 40.605 67.280 41.605 ;
        RECT 67.850 40.625 68.225 48.410 ;
        RECT 68.500 48.025 70.180 49.260 ;
        RECT 71.015 48.025 75.940 48.035 ;
        RECT 68.500 47.545 75.940 48.025 ;
        RECT 68.500 45.285 70.180 47.545 ;
        RECT 71.015 47.125 75.940 47.545 ;
        RECT 70.520 46.935 70.775 46.960 ;
        RECT 70.520 46.920 70.795 46.935 ;
        RECT 70.490 46.645 70.825 46.920 ;
        RECT 71.000 46.895 76.000 47.125 ;
        RECT 76.210 46.935 76.465 46.960 ;
        RECT 70.520 46.630 70.775 46.645 ;
        RECT 71.000 46.455 76.000 46.685 ;
        RECT 76.205 46.645 76.465 46.935 ;
        RECT 76.210 46.630 76.465 46.645 ;
        RECT 71.045 46.445 75.900 46.455 ;
        RECT 71.045 44.920 73.690 44.925 ;
        RECT 69.720 44.720 73.690 44.920 ;
        RECT 69.720 44.690 73.680 44.720 ;
        RECT 68.560 44.335 68.895 44.610 ;
        RECT 69.440 44.440 69.670 44.485 ;
        RECT 64.420 40.560 64.775 40.580 ;
        RECT 64.420 40.490 64.650 40.560 ;
        RECT 65.560 40.490 65.790 40.580 ;
        RECT 66.320 40.465 67.230 40.605 ;
        RECT 67.850 40.490 68.240 40.625 ;
        RECT 66.310 40.285 67.320 40.465 ;
        RECT 62.410 40.055 64.370 40.285 ;
        RECT 65.840 40.055 67.800 40.285 ;
        RECT 63.115 39.230 63.460 40.055 ;
        RECT 65.865 40.050 67.750 40.055 ;
        RECT 68.045 38.355 68.240 40.490 ;
        RECT 68.630 38.830 68.820 44.335 ;
        RECT 69.250 43.105 69.670 44.440 ;
        RECT 70.975 43.105 72.320 44.690 ;
        RECT 69.250 41.720 72.320 43.105 ;
        RECT 69.250 40.990 69.670 41.720 ;
        RECT 69.245 40.485 69.670 40.990 ;
        RECT 68.630 38.640 68.945 38.830 ;
        RECT 58.950 38.125 62.910 38.355 ;
        RECT 64.380 38.125 68.340 38.355 ;
        RECT 68.755 38.130 68.945 38.640 ;
        RECT 58.670 37.515 58.900 37.965 ;
        RECT 60.150 37.515 60.940 38.125 ;
        RECT 58.670 37.210 60.940 37.515 ;
        RECT 58.615 37.195 60.940 37.210 ;
        RECT 58.530 36.350 60.940 37.195 ;
        RECT 58.530 35.975 58.900 36.350 ;
        RECT 58.670 35.965 58.900 35.975 ;
        RECT 60.150 35.805 60.940 36.350 ;
        RECT 62.960 37.880 63.190 37.965 ;
        RECT 64.100 37.880 64.330 37.965 ;
        RECT 62.960 36.055 64.330 37.880 ;
        RECT 62.960 35.965 63.190 36.055 ;
        RECT 58.950 35.575 62.910 35.805 ;
        RECT 55.590 35.255 58.085 35.280 ;
        RECT 58.530 35.255 58.755 35.265 ;
        RECT 63.430 35.255 63.920 36.055 ;
        RECT 64.100 35.965 64.330 36.055 ;
        RECT 65.815 37.745 67.155 38.125 ;
        RECT 68.390 37.745 68.620 37.965 ;
        RECT 65.815 36.150 68.620 37.745 ;
        RECT 65.815 35.805 67.155 36.150 ;
        RECT 68.390 35.965 68.620 36.150 ;
        RECT 64.380 35.575 68.340 35.805 ;
        RECT 68.770 35.785 68.945 38.130 ;
        RECT 69.245 37.965 69.540 40.485 ;
        RECT 70.975 40.280 72.320 41.720 ;
        RECT 73.730 44.390 73.960 44.485 ;
        RECT 74.205 44.390 74.695 46.445 ;
        RECT 75.265 44.920 75.900 44.925 ;
        RECT 75.150 44.690 79.110 44.920 ;
        RECT 74.870 44.390 75.100 44.485 ;
        RECT 73.730 40.565 75.100 44.390 ;
        RECT 73.730 40.485 73.960 40.565 ;
        RECT 74.870 40.485 75.100 40.565 ;
        RECT 76.525 40.280 77.870 44.690 ;
        RECT 79.160 44.420 79.390 44.485 ;
        RECT 80.045 44.425 80.520 49.260 ;
        RECT 81.845 48.455 82.525 49.260 ;
        RECT 82.945 48.735 83.280 48.985 ;
        RECT 82.960 48.710 83.250 48.735 ;
        RECT 86.420 48.635 88.330 49.260 ;
        RECT 90.420 48.925 92.305 48.930 ;
        RECT 93.865 48.925 95.750 48.930 ;
        RECT 90.410 48.695 92.370 48.925 ;
        RECT 93.840 48.695 95.800 48.925 ;
        RECT 82.770 48.455 83.000 48.505 ;
        RECT 81.845 47.955 83.000 48.455 ;
        RECT 80.915 44.735 81.250 44.985 ;
        RECT 80.935 44.705 81.225 44.735 ;
        RECT 80.745 44.425 80.975 44.500 ;
        RECT 79.160 40.485 79.615 44.420 ;
        RECT 80.045 43.680 80.975 44.425 ;
        RECT 80.380 40.565 80.975 43.680 ;
        RECT 80.745 40.500 80.975 40.565 ;
        RECT 81.185 44.475 81.415 44.500 ;
        RECT 81.185 40.920 81.695 44.475 ;
        RECT 81.185 40.550 81.880 40.920 ;
        RECT 82.380 40.600 83.000 47.955 ;
        RECT 81.185 40.500 81.415 40.550 ;
        RECT 69.720 40.250 73.680 40.280 ;
        RECT 75.150 40.250 79.110 40.280 ;
        RECT 69.720 40.090 79.110 40.250 ;
        RECT 69.720 40.050 73.680 40.090 ;
        RECT 75.150 40.050 79.110 40.090 ;
        RECT 79.275 38.660 79.615 40.485 ;
        RECT 80.925 38.660 81.345 40.305 ;
        RECT 79.275 38.505 81.345 38.660 ;
        RECT 79.350 38.390 81.345 38.505 ;
        RECT 69.810 38.125 73.770 38.355 ;
        RECT 75.240 38.125 79.200 38.355 ;
        RECT 69.245 37.205 69.760 37.965 ;
        RECT 69.315 36.025 69.760 37.205 ;
        RECT 69.530 35.965 69.760 36.025 ;
        RECT 71.190 35.805 72.145 38.125 ;
        RECT 73.820 37.900 74.050 37.965 ;
        RECT 74.960 37.900 75.190 37.965 ;
        RECT 73.820 36.030 75.190 37.900 ;
        RECT 73.820 35.965 74.050 36.030 ;
        RECT 68.755 35.255 68.945 35.785 ;
        RECT 69.810 35.575 73.770 35.805 ;
        RECT 74.225 35.255 74.780 36.030 ;
        RECT 74.960 35.965 75.190 36.030 ;
        RECT 76.635 35.805 77.590 38.125 ;
        RECT 79.350 37.970 79.615 38.390 ;
        RECT 80.925 38.115 81.345 38.390 ;
        RECT 81.580 39.355 81.880 40.550 ;
        RECT 82.770 40.505 83.000 40.600 ;
        RECT 83.210 48.430 83.440 48.505 ;
        RECT 83.210 41.110 83.985 48.430 ;
        RECT 86.385 48.405 88.385 48.635 ;
        RECT 90.130 48.410 90.360 48.490 ;
        RECT 85.950 45.060 86.180 48.355 ;
        RECT 88.590 48.275 88.820 48.355 ;
        RECT 88.560 45.060 88.820 48.275 ;
        RECT 85.950 43.245 88.820 45.060 ;
        RECT 83.210 40.580 84.060 41.110 ;
        RECT 85.950 40.825 86.180 43.245 ;
        RECT 83.210 40.505 83.440 40.580 ;
        RECT 82.875 39.825 83.390 40.315 ;
        RECT 82.875 39.360 83.385 39.825 ;
        RECT 83.690 39.795 84.060 40.580 ;
        RECT 85.590 40.395 86.180 40.825 ;
        RECT 87.075 40.640 87.335 40.960 ;
        RECT 88.560 40.645 88.820 43.245 ;
        RECT 89.890 40.990 90.360 48.410 ;
        RECT 90.850 41.775 91.740 48.695 ;
        RECT 92.420 48.390 92.650 48.490 ;
        RECT 92.420 48.380 92.775 48.390 ;
        RECT 93.560 48.380 93.790 48.490 ;
        RECT 87.130 40.480 87.280 40.640 ;
        RECT 82.510 39.355 83.385 39.360 ;
        RECT 81.580 38.950 83.385 39.355 ;
        RECT 81.580 38.110 81.880 38.950 ;
        RECT 82.510 38.935 83.385 38.950 ;
        RECT 82.875 38.825 83.385 38.935 ;
        RECT 82.875 38.125 83.390 38.825 ;
        RECT 83.585 38.795 84.615 39.795 ;
        RECT 79.275 37.965 79.615 37.970 ;
        RECT 79.250 36.020 79.615 37.965 ;
        RECT 80.830 37.900 81.060 37.970 ;
        RECT 80.335 37.230 81.060 37.900 ;
        RECT 80.325 37.040 81.060 37.230 ;
        RECT 80.325 36.240 80.680 37.040 ;
        RECT 80.830 36.970 81.060 37.040 ;
        RECT 81.270 37.925 81.500 37.970 ;
        RECT 81.640 37.925 81.880 38.110 ;
        RECT 81.270 37.595 81.880 37.925 ;
        RECT 82.855 37.870 83.085 37.975 ;
        RECT 81.270 37.040 81.765 37.595 ;
        RECT 81.270 36.970 81.500 37.040 ;
        RECT 81.020 36.785 81.310 36.810 ;
        RECT 81.005 36.535 81.340 36.785 ;
        RECT 82.625 36.765 83.085 37.870 ;
        RECT 82.305 36.240 83.085 36.765 ;
        RECT 79.885 36.060 83.085 36.240 ;
        RECT 79.250 35.965 79.480 36.020 ;
        RECT 79.885 35.960 82.690 36.060 ;
        RECT 82.855 35.975 83.085 36.060 ;
        RECT 83.295 37.910 83.525 37.975 ;
        RECT 83.690 37.910 84.060 38.795 ;
        RECT 83.295 37.585 84.060 37.910 ;
        RECT 83.295 36.045 84.055 37.585 ;
        RECT 83.295 35.975 83.525 36.045 ;
        RECT 75.240 35.575 79.200 35.805 ;
        RECT 79.830 35.785 82.690 35.960 ;
        RECT 83.045 35.795 83.335 35.815 ;
        RECT 79.870 35.620 82.690 35.785 ;
        RECT 79.870 35.255 82.350 35.620 ;
        RECT 83.020 35.545 83.355 35.795 ;
        RECT 85.590 35.280 86.085 40.395 ;
        RECT 87.105 40.345 87.310 40.480 ;
        RECT 88.590 40.395 88.820 40.645 ;
        RECT 89.610 40.550 90.360 40.990 ;
        RECT 90.780 40.775 91.795 41.775 ;
        RECT 86.385 40.115 88.385 40.345 ;
        RECT 89.610 38.355 89.980 40.550 ;
        RECT 90.130 40.490 90.360 40.550 ;
        RECT 90.850 40.285 91.740 40.775 ;
        RECT 92.420 40.580 93.790 48.380 ;
        RECT 94.325 43.635 95.215 48.695 ;
        RECT 95.850 48.410 96.080 48.490 ;
        RECT 94.320 42.015 95.220 43.635 ;
        RECT 94.325 41.605 95.215 42.015 ;
        RECT 94.250 40.605 95.280 41.605 ;
        RECT 95.850 40.625 96.225 48.410 ;
        RECT 96.500 48.025 98.180 49.260 ;
        RECT 99.015 48.025 103.940 48.035 ;
        RECT 96.500 47.545 103.940 48.025 ;
        RECT 96.500 45.285 98.180 47.545 ;
        RECT 99.015 47.125 103.940 47.545 ;
        RECT 98.520 46.935 98.775 46.960 ;
        RECT 98.520 46.920 98.795 46.935 ;
        RECT 98.490 46.645 98.825 46.920 ;
        RECT 99.000 46.895 104.000 47.125 ;
        RECT 104.210 46.935 104.465 46.960 ;
        RECT 98.520 46.630 98.775 46.645 ;
        RECT 99.000 46.455 104.000 46.685 ;
        RECT 104.205 46.645 104.465 46.935 ;
        RECT 104.210 46.630 104.465 46.645 ;
        RECT 99.045 46.445 103.900 46.455 ;
        RECT 99.045 44.920 101.690 44.925 ;
        RECT 97.720 44.720 101.690 44.920 ;
        RECT 97.720 44.690 101.680 44.720 ;
        RECT 96.560 44.335 96.895 44.610 ;
        RECT 97.440 44.440 97.670 44.485 ;
        RECT 92.420 40.560 92.775 40.580 ;
        RECT 92.420 40.490 92.650 40.560 ;
        RECT 93.560 40.490 93.790 40.580 ;
        RECT 94.320 40.465 95.230 40.605 ;
        RECT 95.850 40.490 96.240 40.625 ;
        RECT 94.310 40.285 95.320 40.465 ;
        RECT 90.410 40.055 92.370 40.285 ;
        RECT 93.840 40.055 95.800 40.285 ;
        RECT 91.095 39.170 91.495 40.055 ;
        RECT 93.865 40.050 95.750 40.055 ;
        RECT 96.045 38.355 96.240 40.490 ;
        RECT 96.630 38.830 96.820 44.335 ;
        RECT 97.250 43.105 97.670 44.440 ;
        RECT 98.975 43.105 100.320 44.690 ;
        RECT 97.250 41.720 100.320 43.105 ;
        RECT 97.250 40.990 97.670 41.720 ;
        RECT 97.245 40.485 97.670 40.990 ;
        RECT 96.630 38.640 96.945 38.830 ;
        RECT 86.950 38.125 90.910 38.355 ;
        RECT 92.380 38.125 96.340 38.355 ;
        RECT 96.755 38.130 96.945 38.640 ;
        RECT 86.670 37.515 86.900 37.965 ;
        RECT 88.150 37.515 88.940 38.125 ;
        RECT 86.670 37.210 88.940 37.515 ;
        RECT 86.615 37.195 88.940 37.210 ;
        RECT 86.530 36.350 88.940 37.195 ;
        RECT 86.530 35.975 86.900 36.350 ;
        RECT 86.670 35.965 86.900 35.975 ;
        RECT 88.150 35.805 88.940 36.350 ;
        RECT 90.960 37.880 91.190 37.965 ;
        RECT 92.100 37.880 92.330 37.965 ;
        RECT 90.960 36.055 92.330 37.880 ;
        RECT 90.960 35.965 91.190 36.055 ;
        RECT 86.950 35.575 90.910 35.805 ;
        RECT 83.590 35.255 86.085 35.280 ;
        RECT 86.530 35.255 86.755 35.265 ;
        RECT 91.430 35.255 91.920 36.055 ;
        RECT 92.100 35.965 92.330 36.055 ;
        RECT 93.815 37.745 95.155 38.125 ;
        RECT 96.390 37.745 96.620 37.965 ;
        RECT 93.815 36.150 96.620 37.745 ;
        RECT 93.815 35.805 95.155 36.150 ;
        RECT 96.390 35.965 96.620 36.150 ;
        RECT 92.380 35.575 96.340 35.805 ;
        RECT 96.770 35.785 96.945 38.130 ;
        RECT 97.245 37.965 97.540 40.485 ;
        RECT 98.975 40.280 100.320 41.720 ;
        RECT 101.730 44.390 101.960 44.485 ;
        RECT 102.205 44.390 102.695 46.445 ;
        RECT 103.265 44.920 103.900 44.925 ;
        RECT 103.150 44.690 107.110 44.920 ;
        RECT 102.870 44.390 103.100 44.485 ;
        RECT 101.730 40.565 103.100 44.390 ;
        RECT 101.730 40.485 101.960 40.565 ;
        RECT 102.870 40.485 103.100 40.565 ;
        RECT 104.525 40.280 105.870 44.690 ;
        RECT 107.160 44.420 107.390 44.485 ;
        RECT 108.045 44.425 108.520 49.260 ;
        RECT 109.845 48.455 110.525 49.260 ;
        RECT 110.945 48.735 111.280 48.985 ;
        RECT 110.960 48.710 111.250 48.735 ;
        RECT 114.420 48.635 116.330 49.260 ;
        RECT 118.420 48.925 120.305 48.930 ;
        RECT 121.865 48.925 123.750 48.930 ;
        RECT 118.410 48.695 120.370 48.925 ;
        RECT 121.840 48.695 123.800 48.925 ;
        RECT 110.770 48.455 111.000 48.505 ;
        RECT 109.845 47.955 111.000 48.455 ;
        RECT 108.915 44.735 109.250 44.985 ;
        RECT 108.935 44.705 109.225 44.735 ;
        RECT 108.745 44.425 108.975 44.500 ;
        RECT 107.160 40.485 107.615 44.420 ;
        RECT 108.045 43.680 108.975 44.425 ;
        RECT 108.380 40.565 108.975 43.680 ;
        RECT 108.745 40.500 108.975 40.565 ;
        RECT 109.185 44.475 109.415 44.500 ;
        RECT 109.185 40.920 109.695 44.475 ;
        RECT 109.185 40.550 109.880 40.920 ;
        RECT 110.380 40.600 111.000 47.955 ;
        RECT 109.185 40.500 109.415 40.550 ;
        RECT 97.720 40.250 101.680 40.280 ;
        RECT 103.150 40.250 107.110 40.280 ;
        RECT 97.720 40.090 107.110 40.250 ;
        RECT 97.720 40.050 101.680 40.090 ;
        RECT 103.150 40.050 107.110 40.090 ;
        RECT 107.275 38.660 107.615 40.485 ;
        RECT 108.925 38.660 109.345 40.305 ;
        RECT 107.275 38.505 109.345 38.660 ;
        RECT 107.350 38.390 109.345 38.505 ;
        RECT 97.810 38.125 101.770 38.355 ;
        RECT 103.240 38.125 107.200 38.355 ;
        RECT 97.245 37.205 97.760 37.965 ;
        RECT 97.315 36.025 97.760 37.205 ;
        RECT 97.530 35.965 97.760 36.025 ;
        RECT 99.190 35.805 100.145 38.125 ;
        RECT 101.820 37.900 102.050 37.965 ;
        RECT 102.960 37.900 103.190 37.965 ;
        RECT 101.820 36.030 103.190 37.900 ;
        RECT 101.820 35.965 102.050 36.030 ;
        RECT 96.755 35.255 96.945 35.785 ;
        RECT 97.810 35.575 101.770 35.805 ;
        RECT 102.225 35.255 102.780 36.030 ;
        RECT 102.960 35.965 103.190 36.030 ;
        RECT 104.635 35.805 105.590 38.125 ;
        RECT 107.350 37.970 107.615 38.390 ;
        RECT 108.925 38.115 109.345 38.390 ;
        RECT 109.580 39.355 109.880 40.550 ;
        RECT 110.770 40.505 111.000 40.600 ;
        RECT 111.210 48.430 111.440 48.505 ;
        RECT 111.210 41.110 111.985 48.430 ;
        RECT 114.385 48.405 116.385 48.635 ;
        RECT 118.130 48.410 118.360 48.490 ;
        RECT 113.950 45.060 114.180 48.355 ;
        RECT 116.590 48.275 116.820 48.355 ;
        RECT 116.560 45.060 116.820 48.275 ;
        RECT 113.950 43.245 116.820 45.060 ;
        RECT 111.210 40.580 112.060 41.110 ;
        RECT 113.950 40.825 114.180 43.245 ;
        RECT 111.210 40.505 111.440 40.580 ;
        RECT 110.875 39.825 111.390 40.315 ;
        RECT 110.875 39.360 111.385 39.825 ;
        RECT 111.690 39.795 112.060 40.580 ;
        RECT 113.590 40.395 114.180 40.825 ;
        RECT 115.075 40.640 115.335 40.960 ;
        RECT 116.560 40.645 116.820 43.245 ;
        RECT 117.890 40.990 118.360 48.410 ;
        RECT 118.850 41.775 119.740 48.695 ;
        RECT 120.420 48.390 120.650 48.490 ;
        RECT 120.420 48.380 120.775 48.390 ;
        RECT 121.560 48.380 121.790 48.490 ;
        RECT 115.130 40.480 115.280 40.640 ;
        RECT 110.510 39.355 111.385 39.360 ;
        RECT 109.580 38.950 111.385 39.355 ;
        RECT 109.580 38.110 109.880 38.950 ;
        RECT 110.510 38.935 111.385 38.950 ;
        RECT 110.875 38.825 111.385 38.935 ;
        RECT 110.875 38.125 111.390 38.825 ;
        RECT 111.585 38.795 112.615 39.795 ;
        RECT 107.275 37.965 107.615 37.970 ;
        RECT 107.250 36.020 107.615 37.965 ;
        RECT 108.830 37.900 109.060 37.970 ;
        RECT 108.335 37.230 109.060 37.900 ;
        RECT 108.325 37.040 109.060 37.230 ;
        RECT 108.325 36.240 108.680 37.040 ;
        RECT 108.830 36.970 109.060 37.040 ;
        RECT 109.270 37.925 109.500 37.970 ;
        RECT 109.640 37.925 109.880 38.110 ;
        RECT 109.270 37.595 109.880 37.925 ;
        RECT 110.855 37.870 111.085 37.975 ;
        RECT 109.270 37.040 109.765 37.595 ;
        RECT 109.270 36.970 109.500 37.040 ;
        RECT 109.020 36.785 109.310 36.810 ;
        RECT 109.005 36.535 109.340 36.785 ;
        RECT 110.625 36.765 111.085 37.870 ;
        RECT 110.305 36.240 111.085 36.765 ;
        RECT 107.885 36.060 111.085 36.240 ;
        RECT 107.250 35.965 107.480 36.020 ;
        RECT 103.240 35.575 107.200 35.805 ;
        RECT 107.885 35.620 110.690 36.060 ;
        RECT 110.855 35.975 111.085 36.060 ;
        RECT 111.295 37.910 111.525 37.975 ;
        RECT 111.690 37.910 112.060 38.795 ;
        RECT 111.295 37.585 112.060 37.910 ;
        RECT 111.295 36.045 112.055 37.585 ;
        RECT 111.295 35.975 111.525 36.045 ;
        RECT 111.045 35.795 111.335 35.815 ;
        RECT 107.885 35.255 110.350 35.620 ;
        RECT 111.020 35.545 111.355 35.795 ;
        RECT 113.590 35.280 114.085 40.395 ;
        RECT 115.105 40.345 115.310 40.480 ;
        RECT 116.590 40.395 116.820 40.645 ;
        RECT 117.610 40.550 118.360 40.990 ;
        RECT 118.780 40.775 119.795 41.775 ;
        RECT 114.385 40.115 116.385 40.345 ;
        RECT 117.610 38.355 117.980 40.550 ;
        RECT 118.130 40.490 118.360 40.550 ;
        RECT 118.850 40.285 119.740 40.775 ;
        RECT 120.420 40.580 121.790 48.380 ;
        RECT 122.325 43.635 123.215 48.695 ;
        RECT 123.850 48.410 124.080 48.490 ;
        RECT 122.320 42.015 123.220 43.635 ;
        RECT 122.325 41.605 123.215 42.015 ;
        RECT 122.250 40.605 123.280 41.605 ;
        RECT 123.850 40.625 124.225 48.410 ;
        RECT 124.500 48.025 126.180 49.260 ;
        RECT 127.015 48.025 131.940 48.035 ;
        RECT 124.500 47.545 131.940 48.025 ;
        RECT 124.500 45.285 126.180 47.545 ;
        RECT 127.015 47.125 131.940 47.545 ;
        RECT 126.520 46.935 126.775 46.960 ;
        RECT 126.520 46.920 126.795 46.935 ;
        RECT 126.490 46.645 126.825 46.920 ;
        RECT 127.000 46.895 132.000 47.125 ;
        RECT 132.210 46.935 132.465 46.960 ;
        RECT 126.520 46.630 126.775 46.645 ;
        RECT 127.000 46.455 132.000 46.685 ;
        RECT 132.205 46.645 132.465 46.935 ;
        RECT 132.210 46.630 132.465 46.645 ;
        RECT 127.045 46.445 131.900 46.455 ;
        RECT 127.045 44.920 129.690 44.925 ;
        RECT 125.720 44.720 129.690 44.920 ;
        RECT 125.720 44.690 129.680 44.720 ;
        RECT 124.560 44.335 124.895 44.610 ;
        RECT 125.440 44.440 125.670 44.485 ;
        RECT 120.420 40.560 120.775 40.580 ;
        RECT 120.420 40.490 120.650 40.560 ;
        RECT 121.560 40.490 121.790 40.580 ;
        RECT 122.320 40.465 123.230 40.605 ;
        RECT 123.850 40.490 124.240 40.625 ;
        RECT 122.310 40.285 123.320 40.465 ;
        RECT 118.410 40.055 120.370 40.285 ;
        RECT 121.840 40.055 123.800 40.285 ;
        RECT 119.145 39.135 119.430 40.055 ;
        RECT 121.865 40.050 123.750 40.055 ;
        RECT 124.045 38.355 124.240 40.490 ;
        RECT 124.630 38.830 124.820 44.335 ;
        RECT 125.250 43.105 125.670 44.440 ;
        RECT 126.975 43.105 128.320 44.690 ;
        RECT 125.250 41.720 128.320 43.105 ;
        RECT 125.250 40.990 125.670 41.720 ;
        RECT 125.245 40.485 125.670 40.990 ;
        RECT 124.630 38.640 124.945 38.830 ;
        RECT 114.950 38.125 118.910 38.355 ;
        RECT 120.380 38.125 124.340 38.355 ;
        RECT 124.755 38.130 124.945 38.640 ;
        RECT 114.670 37.515 114.900 37.965 ;
        RECT 116.150 37.515 116.940 38.125 ;
        RECT 114.670 37.210 116.940 37.515 ;
        RECT 114.615 37.195 116.940 37.210 ;
        RECT 114.530 36.350 116.940 37.195 ;
        RECT 114.530 35.975 114.900 36.350 ;
        RECT 114.670 35.965 114.900 35.975 ;
        RECT 116.150 35.805 116.940 36.350 ;
        RECT 118.960 37.880 119.190 37.965 ;
        RECT 120.100 37.880 120.330 37.965 ;
        RECT 118.960 36.055 120.330 37.880 ;
        RECT 118.960 35.965 119.190 36.055 ;
        RECT 114.950 35.575 118.910 35.805 ;
        RECT 111.490 35.255 114.190 35.280 ;
        RECT 114.530 35.255 114.755 35.265 ;
        RECT 119.430 35.255 119.920 36.055 ;
        RECT 120.100 35.965 120.330 36.055 ;
        RECT 121.815 37.745 123.155 38.125 ;
        RECT 124.390 37.745 124.620 37.965 ;
        RECT 121.815 36.150 124.620 37.745 ;
        RECT 121.815 35.805 123.155 36.150 ;
        RECT 124.390 35.965 124.620 36.150 ;
        RECT 120.380 35.575 124.340 35.805 ;
        RECT 124.770 35.785 124.945 38.130 ;
        RECT 125.245 37.965 125.540 40.485 ;
        RECT 126.975 40.280 128.320 41.720 ;
        RECT 129.730 44.390 129.960 44.485 ;
        RECT 130.205 44.390 130.695 46.445 ;
        RECT 131.265 44.920 131.900 44.925 ;
        RECT 131.150 44.690 135.110 44.920 ;
        RECT 130.870 44.390 131.100 44.485 ;
        RECT 129.730 40.565 131.100 44.390 ;
        RECT 129.730 40.485 129.960 40.565 ;
        RECT 130.870 40.485 131.100 40.565 ;
        RECT 132.525 40.280 133.870 44.690 ;
        RECT 135.160 44.420 135.390 44.485 ;
        RECT 136.045 44.425 136.520 49.260 ;
        RECT 137.845 48.455 138.525 49.260 ;
        RECT 138.945 48.735 139.280 48.985 ;
        RECT 138.960 48.710 139.250 48.735 ;
        RECT 144.150 48.720 146.255 49.310 ;
        RECT 146.835 48.720 148.940 49.310 ;
        RECT 138.770 48.455 139.000 48.505 ;
        RECT 137.845 47.955 139.000 48.455 ;
        RECT 136.915 44.735 137.250 44.985 ;
        RECT 136.935 44.705 137.225 44.735 ;
        RECT 136.745 44.425 136.975 44.500 ;
        RECT 135.160 40.485 135.615 44.420 ;
        RECT 136.045 43.680 136.975 44.425 ;
        RECT 136.380 40.565 136.975 43.680 ;
        RECT 136.745 40.500 136.975 40.565 ;
        RECT 137.185 44.475 137.415 44.500 ;
        RECT 137.185 40.920 137.695 44.475 ;
        RECT 137.185 40.550 137.880 40.920 ;
        RECT 138.380 40.600 139.000 47.955 ;
        RECT 137.185 40.500 137.415 40.550 ;
        RECT 125.720 40.250 129.680 40.280 ;
        RECT 131.150 40.250 135.110 40.280 ;
        RECT 125.720 40.090 135.110 40.250 ;
        RECT 125.720 40.050 129.680 40.090 ;
        RECT 131.150 40.050 135.110 40.090 ;
        RECT 135.275 38.660 135.615 40.485 ;
        RECT 136.925 38.660 137.345 40.305 ;
        RECT 135.275 38.505 137.345 38.660 ;
        RECT 135.350 38.390 137.345 38.505 ;
        RECT 125.810 38.125 129.770 38.355 ;
        RECT 131.240 38.125 135.200 38.355 ;
        RECT 125.245 37.205 125.760 37.965 ;
        RECT 125.315 36.025 125.760 37.205 ;
        RECT 125.530 35.965 125.760 36.025 ;
        RECT 127.190 35.805 128.145 38.125 ;
        RECT 129.820 37.900 130.050 37.965 ;
        RECT 130.960 37.900 131.190 37.965 ;
        RECT 129.820 36.030 131.190 37.900 ;
        RECT 129.820 35.965 130.050 36.030 ;
        RECT 124.755 35.255 124.945 35.785 ;
        RECT 125.810 35.575 129.770 35.805 ;
        RECT 130.225 35.255 130.780 36.030 ;
        RECT 130.960 35.965 131.190 36.030 ;
        RECT 132.635 35.805 133.590 38.125 ;
        RECT 135.350 37.970 135.615 38.390 ;
        RECT 136.925 38.115 137.345 38.390 ;
        RECT 137.580 39.355 137.880 40.550 ;
        RECT 138.770 40.505 139.000 40.600 ;
        RECT 139.210 48.430 139.440 48.505 ;
        RECT 139.210 41.110 139.985 48.430 ;
        RECT 146.860 47.490 148.890 48.720 ;
        RECT 144.150 46.900 146.255 47.490 ;
        RECT 146.835 46.900 148.940 47.490 ;
        RECT 144.160 45.670 146.190 46.900 ;
        RECT 146.890 46.880 148.890 46.900 ;
        RECT 146.890 45.670 154.890 45.680 ;
        RECT 144.150 45.080 146.255 45.670 ;
        RECT 146.835 45.180 154.890 45.670 ;
        RECT 146.835 45.080 148.940 45.180 ;
        RECT 144.190 43.850 146.190 43.880 ;
        RECT 144.150 43.260 146.255 43.850 ;
        RECT 146.835 43.780 148.940 43.850 ;
        RECT 149.425 43.780 149.925 44.125 ;
        RECT 152.890 43.850 154.890 45.180 ;
        RECT 150.130 43.780 152.235 43.850 ;
        RECT 146.835 43.280 152.235 43.780 ;
        RECT 146.835 43.260 148.940 43.280 ;
        RECT 150.130 43.260 152.235 43.280 ;
        RECT 152.815 43.260 154.920 43.850 ;
        RECT 144.190 42.945 146.190 43.260 ;
        RECT 141.790 42.505 146.190 42.945 ;
        RECT 144.190 42.030 146.190 42.505 ;
        RECT 144.150 41.440 146.255 42.030 ;
        RECT 146.835 41.980 148.940 42.030 ;
        RECT 150.130 41.980 152.235 42.030 ;
        RECT 146.835 41.480 152.235 41.980 ;
        RECT 146.835 41.440 148.940 41.480 ;
        RECT 149.530 41.440 152.235 41.480 ;
        RECT 152.815 41.440 154.920 42.030 ;
        RECT 149.530 41.240 150.310 41.440 ;
        RECT 139.210 40.580 140.060 41.110 ;
        RECT 149.530 41.035 150.030 41.240 ;
        RECT 139.210 40.505 139.440 40.580 ;
        RECT 138.875 39.825 139.390 40.315 ;
        RECT 138.875 39.360 139.385 39.825 ;
        RECT 139.690 39.795 140.060 40.580 ;
        RECT 142.350 40.535 150.030 41.035 ;
        RECT 153.565 40.995 154.355 41.440 ;
        RECT 150.785 40.205 154.355 40.995 ;
        RECT 150.785 40.055 151.575 40.205 ;
        RECT 138.510 39.355 139.385 39.360 ;
        RECT 137.580 38.950 139.385 39.355 ;
        RECT 137.580 38.110 137.880 38.950 ;
        RECT 138.510 38.935 139.385 38.950 ;
        RECT 138.875 38.825 139.385 38.935 ;
        RECT 138.875 38.125 139.390 38.825 ;
        RECT 139.585 38.795 140.615 39.795 ;
        RECT 141.105 39.265 151.575 40.055 ;
        RECT 135.275 37.965 135.615 37.970 ;
        RECT 135.250 36.020 135.615 37.965 ;
        RECT 136.830 37.900 137.060 37.970 ;
        RECT 136.335 37.230 137.060 37.900 ;
        RECT 136.325 37.040 137.060 37.230 ;
        RECT 136.325 36.240 136.680 37.040 ;
        RECT 136.830 36.970 137.060 37.040 ;
        RECT 137.270 37.925 137.500 37.970 ;
        RECT 137.640 37.925 137.880 38.110 ;
        RECT 137.270 37.595 137.880 37.925 ;
        RECT 138.855 37.870 139.085 37.975 ;
        RECT 137.270 37.040 137.765 37.595 ;
        RECT 137.270 36.970 137.500 37.040 ;
        RECT 137.020 36.785 137.310 36.810 ;
        RECT 137.005 36.535 137.340 36.785 ;
        RECT 138.625 36.765 139.085 37.870 ;
        RECT 138.305 36.240 139.085 36.765 ;
        RECT 135.885 36.060 139.085 36.240 ;
        RECT 135.250 35.965 135.480 36.020 ;
        RECT 131.240 35.575 135.200 35.805 ;
        RECT 135.885 35.620 138.690 36.060 ;
        RECT 138.855 35.975 139.085 36.060 ;
        RECT 139.295 37.910 139.525 37.975 ;
        RECT 139.690 37.910 140.060 38.795 ;
        RECT 139.295 37.585 140.060 37.910 ;
        RECT 139.295 36.045 140.055 37.585 ;
        RECT 139.295 35.975 139.525 36.045 ;
        RECT 139.045 35.795 139.335 35.815 ;
        RECT 135.885 35.335 138.350 35.620 ;
        RECT 139.020 35.545 139.355 35.795 ;
        RECT 141.105 35.335 141.895 39.265 ;
        RECT 135.885 35.255 141.895 35.335 ;
        RECT 1.475 34.545 141.895 35.255 ;
        RECT 1.475 34.380 140.080 34.545 ;
        RECT 27.790 33.960 30.490 33.980 ;
        RECT 55.390 33.960 57.990 33.980 ;
        RECT 83.390 33.960 86.290 33.980 ;
        RECT 111.190 33.960 114.190 33.980 ;
        RECT 1.450 33.280 139.925 33.960 ;
        RECT 1.450 33.260 27.925 33.280 ;
        RECT 29.450 33.260 83.925 33.280 ;
        RECT 85.450 33.260 111.925 33.280 ;
        RECT 113.450 33.260 139.925 33.280 ;
        RECT 2.420 32.635 4.330 33.260 ;
        RECT 6.420 32.925 8.305 32.930 ;
        RECT 9.865 32.925 11.750 32.930 ;
        RECT 6.410 32.695 8.370 32.925 ;
        RECT 9.840 32.695 11.800 32.925 ;
        RECT 2.385 32.405 4.385 32.635 ;
        RECT 6.130 32.410 6.360 32.490 ;
        RECT 1.950 29.060 2.180 32.355 ;
        RECT 4.590 32.275 4.820 32.355 ;
        RECT 4.560 29.060 4.820 32.275 ;
        RECT 1.950 27.245 4.820 29.060 ;
        RECT 1.950 24.825 2.180 27.245 ;
        RECT 1.590 24.395 2.180 24.825 ;
        RECT 3.075 24.640 3.335 24.960 ;
        RECT 4.560 24.645 4.820 27.245 ;
        RECT 5.890 24.990 6.360 32.410 ;
        RECT 6.850 25.775 7.740 32.695 ;
        RECT 8.420 32.390 8.650 32.490 ;
        RECT 8.420 32.380 8.775 32.390 ;
        RECT 9.560 32.380 9.790 32.490 ;
        RECT 3.130 24.480 3.280 24.640 ;
        RECT 1.590 19.255 2.085 24.395 ;
        RECT 3.105 24.345 3.310 24.480 ;
        RECT 4.590 24.395 4.820 24.645 ;
        RECT 5.610 24.550 6.360 24.990 ;
        RECT 6.780 24.775 7.795 25.775 ;
        RECT 2.385 24.115 4.385 24.345 ;
        RECT 5.610 22.355 5.980 24.550 ;
        RECT 6.130 24.490 6.360 24.550 ;
        RECT 6.850 24.285 7.740 24.775 ;
        RECT 8.420 24.580 9.790 32.380 ;
        RECT 10.325 27.635 11.215 32.695 ;
        RECT 11.850 32.410 12.080 32.490 ;
        RECT 10.320 26.015 11.220 27.635 ;
        RECT 10.325 25.605 11.215 26.015 ;
        RECT 10.250 24.605 11.280 25.605 ;
        RECT 11.850 24.625 12.225 32.410 ;
        RECT 12.500 32.025 14.180 33.260 ;
        RECT 15.015 32.025 19.940 32.035 ;
        RECT 12.500 31.545 19.940 32.025 ;
        RECT 12.500 29.285 14.180 31.545 ;
        RECT 15.015 31.125 19.940 31.545 ;
        RECT 14.520 30.935 14.775 30.960 ;
        RECT 14.520 30.920 14.795 30.935 ;
        RECT 14.490 30.645 14.825 30.920 ;
        RECT 15.000 30.895 20.000 31.125 ;
        RECT 20.210 30.935 20.465 30.960 ;
        RECT 14.520 30.630 14.775 30.645 ;
        RECT 15.000 30.455 20.000 30.685 ;
        RECT 20.205 30.645 20.465 30.935 ;
        RECT 20.210 30.630 20.465 30.645 ;
        RECT 15.045 30.445 19.900 30.455 ;
        RECT 15.045 28.920 17.690 28.925 ;
        RECT 13.720 28.720 17.690 28.920 ;
        RECT 13.720 28.690 17.680 28.720 ;
        RECT 12.560 28.335 12.895 28.610 ;
        RECT 13.440 28.440 13.670 28.485 ;
        RECT 8.420 24.560 8.775 24.580 ;
        RECT 8.420 24.490 8.650 24.560 ;
        RECT 9.560 24.490 9.790 24.580 ;
        RECT 10.320 24.465 11.230 24.605 ;
        RECT 11.850 24.490 12.240 24.625 ;
        RECT 10.310 24.285 11.320 24.465 ;
        RECT 6.410 24.055 8.370 24.285 ;
        RECT 9.840 24.055 11.800 24.285 ;
        RECT 7.165 23.035 7.495 24.055 ;
        RECT 9.865 24.050 11.750 24.055 ;
        RECT 12.045 22.355 12.240 24.490 ;
        RECT 12.630 22.830 12.820 28.335 ;
        RECT 13.250 27.105 13.670 28.440 ;
        RECT 14.975 27.105 16.320 28.690 ;
        RECT 13.250 25.720 16.320 27.105 ;
        RECT 13.250 24.990 13.670 25.720 ;
        RECT 13.245 24.485 13.670 24.990 ;
        RECT 12.630 22.640 12.945 22.830 ;
        RECT 2.950 22.125 6.910 22.355 ;
        RECT 8.380 22.125 12.340 22.355 ;
        RECT 12.755 22.130 12.945 22.640 ;
        RECT 2.670 21.515 2.900 21.965 ;
        RECT 4.150 21.515 4.940 22.125 ;
        RECT 2.670 21.210 4.940 21.515 ;
        RECT 2.615 21.195 4.940 21.210 ;
        RECT 2.530 20.350 4.940 21.195 ;
        RECT 2.530 19.975 2.900 20.350 ;
        RECT 2.670 19.965 2.900 19.975 ;
        RECT 4.150 19.805 4.940 20.350 ;
        RECT 6.960 21.880 7.190 21.965 ;
        RECT 8.100 21.880 8.330 21.965 ;
        RECT 6.960 20.055 8.330 21.880 ;
        RECT 6.960 19.965 7.190 20.055 ;
        RECT 2.950 19.575 6.910 19.805 ;
        RECT 2.530 19.255 2.755 19.265 ;
        RECT 7.430 19.255 7.920 20.055 ;
        RECT 8.100 19.965 8.330 20.055 ;
        RECT 9.815 21.745 11.155 22.125 ;
        RECT 12.390 21.745 12.620 21.965 ;
        RECT 9.815 20.150 12.620 21.745 ;
        RECT 9.815 19.805 11.155 20.150 ;
        RECT 12.390 19.965 12.620 20.150 ;
        RECT 8.380 19.575 12.340 19.805 ;
        RECT 12.770 19.785 12.945 22.130 ;
        RECT 13.245 21.965 13.540 24.485 ;
        RECT 14.975 24.280 16.320 25.720 ;
        RECT 17.730 28.390 17.960 28.485 ;
        RECT 18.205 28.390 18.695 30.445 ;
        RECT 19.265 28.920 19.900 28.925 ;
        RECT 19.150 28.690 23.110 28.920 ;
        RECT 18.870 28.390 19.100 28.485 ;
        RECT 17.730 24.565 19.100 28.390 ;
        RECT 17.730 24.485 17.960 24.565 ;
        RECT 18.870 24.485 19.100 24.565 ;
        RECT 20.525 24.280 21.870 28.690 ;
        RECT 23.160 28.420 23.390 28.485 ;
        RECT 24.045 28.425 24.520 33.260 ;
        RECT 25.845 32.455 26.525 33.260 ;
        RECT 26.945 32.735 27.280 32.985 ;
        RECT 26.960 32.710 27.250 32.735 ;
        RECT 30.420 32.635 32.330 33.260 ;
        RECT 34.420 32.925 36.305 32.930 ;
        RECT 37.865 32.925 39.750 32.930 ;
        RECT 34.410 32.695 36.370 32.925 ;
        RECT 37.840 32.695 39.800 32.925 ;
        RECT 26.770 32.455 27.000 32.505 ;
        RECT 25.845 31.955 27.000 32.455 ;
        RECT 24.915 28.735 25.250 28.985 ;
        RECT 24.935 28.705 25.225 28.735 ;
        RECT 24.745 28.425 24.975 28.500 ;
        RECT 23.160 24.485 23.615 28.420 ;
        RECT 24.045 27.680 24.975 28.425 ;
        RECT 24.380 24.565 24.975 27.680 ;
        RECT 24.745 24.500 24.975 24.565 ;
        RECT 25.185 28.475 25.415 28.500 ;
        RECT 25.185 24.920 25.695 28.475 ;
        RECT 25.185 24.550 25.880 24.920 ;
        RECT 26.380 24.600 27.000 31.955 ;
        RECT 25.185 24.500 25.415 24.550 ;
        RECT 13.720 24.250 17.680 24.280 ;
        RECT 19.150 24.250 23.110 24.280 ;
        RECT 13.720 24.090 23.110 24.250 ;
        RECT 13.720 24.050 17.680 24.090 ;
        RECT 19.150 24.050 23.110 24.090 ;
        RECT 23.275 22.660 23.615 24.485 ;
        RECT 24.925 22.660 25.345 24.305 ;
        RECT 23.275 22.505 25.345 22.660 ;
        RECT 23.350 22.390 25.345 22.505 ;
        RECT 13.810 22.125 17.770 22.355 ;
        RECT 19.240 22.125 23.200 22.355 ;
        RECT 13.245 21.205 13.760 21.965 ;
        RECT 13.315 20.025 13.760 21.205 ;
        RECT 13.530 19.965 13.760 20.025 ;
        RECT 15.190 19.805 16.145 22.125 ;
        RECT 17.820 21.900 18.050 21.965 ;
        RECT 18.960 21.900 19.190 21.965 ;
        RECT 17.820 20.030 19.190 21.900 ;
        RECT 17.820 19.965 18.050 20.030 ;
        RECT 12.755 19.255 12.945 19.785 ;
        RECT 13.810 19.575 17.770 19.805 ;
        RECT 18.225 19.255 18.780 20.030 ;
        RECT 18.960 19.965 19.190 20.030 ;
        RECT 20.635 19.805 21.590 22.125 ;
        RECT 23.350 21.970 23.615 22.390 ;
        RECT 24.925 22.115 25.345 22.390 ;
        RECT 25.580 23.355 25.880 24.550 ;
        RECT 26.770 24.505 27.000 24.600 ;
        RECT 27.210 32.430 27.440 32.505 ;
        RECT 27.210 25.110 27.985 32.430 ;
        RECT 30.385 32.405 32.385 32.635 ;
        RECT 34.130 32.410 34.360 32.490 ;
        RECT 29.950 29.060 30.180 32.355 ;
        RECT 32.590 32.275 32.820 32.355 ;
        RECT 32.560 29.060 32.820 32.275 ;
        RECT 29.950 27.245 32.820 29.060 ;
        RECT 27.210 24.580 28.060 25.110 ;
        RECT 29.950 24.825 30.180 27.245 ;
        RECT 27.210 24.505 27.440 24.580 ;
        RECT 26.875 23.825 27.390 24.315 ;
        RECT 27.690 23.825 28.060 24.580 ;
        RECT 29.590 24.395 30.180 24.825 ;
        RECT 31.075 24.640 31.335 24.960 ;
        RECT 32.560 24.645 32.820 27.245 ;
        RECT 33.890 24.990 34.360 32.410 ;
        RECT 34.850 25.775 35.740 32.695 ;
        RECT 36.420 32.390 36.650 32.490 ;
        RECT 36.420 32.380 36.775 32.390 ;
        RECT 37.560 32.380 37.790 32.490 ;
        RECT 31.130 24.480 31.280 24.640 ;
        RECT 26.875 23.360 27.385 23.825 ;
        RECT 26.510 23.355 27.385 23.360 ;
        RECT 25.580 22.950 27.385 23.355 ;
        RECT 25.580 22.110 25.880 22.950 ;
        RECT 26.510 22.935 27.385 22.950 ;
        RECT 26.875 22.825 27.385 22.935 ;
        RECT 26.875 22.125 27.390 22.825 ;
        RECT 27.615 22.795 28.615 23.825 ;
        RECT 23.275 21.965 23.615 21.970 ;
        RECT 23.250 20.020 23.615 21.965 ;
        RECT 24.830 21.900 25.060 21.970 ;
        RECT 24.335 21.230 25.060 21.900 ;
        RECT 24.325 21.040 25.060 21.230 ;
        RECT 24.325 20.240 24.680 21.040 ;
        RECT 24.830 20.970 25.060 21.040 ;
        RECT 25.270 21.925 25.500 21.970 ;
        RECT 25.640 21.925 25.880 22.110 ;
        RECT 25.270 21.595 25.880 21.925 ;
        RECT 26.855 21.870 27.085 21.975 ;
        RECT 25.270 21.040 25.765 21.595 ;
        RECT 25.270 20.970 25.500 21.040 ;
        RECT 25.020 20.785 25.310 20.810 ;
        RECT 25.005 20.535 25.340 20.785 ;
        RECT 26.625 20.765 27.085 21.870 ;
        RECT 26.305 20.240 27.085 20.765 ;
        RECT 23.885 20.060 27.085 20.240 ;
        RECT 23.250 19.965 23.480 20.020 ;
        RECT 19.240 19.575 23.200 19.805 ;
        RECT 23.885 19.620 26.690 20.060 ;
        RECT 26.855 19.975 27.085 20.060 ;
        RECT 27.295 21.910 27.525 21.975 ;
        RECT 27.690 21.910 28.060 22.795 ;
        RECT 27.295 21.585 28.060 21.910 ;
        RECT 27.295 20.045 28.055 21.585 ;
        RECT 27.295 19.975 27.525 20.045 ;
        RECT 27.045 19.795 27.335 19.815 ;
        RECT 23.885 19.255 26.350 19.620 ;
        RECT 27.020 19.545 27.355 19.795 ;
        RECT 29.590 19.280 30.085 24.395 ;
        RECT 31.105 24.345 31.310 24.480 ;
        RECT 32.590 24.395 32.820 24.645 ;
        RECT 33.610 24.550 34.360 24.990 ;
        RECT 34.780 24.775 35.795 25.775 ;
        RECT 30.385 24.115 32.385 24.345 ;
        RECT 33.610 22.355 33.980 24.550 ;
        RECT 34.130 24.490 34.360 24.550 ;
        RECT 34.850 24.285 35.740 24.775 ;
        RECT 36.420 24.580 37.790 32.380 ;
        RECT 38.325 27.635 39.215 32.695 ;
        RECT 39.850 32.410 40.080 32.490 ;
        RECT 38.320 26.015 39.220 27.635 ;
        RECT 38.325 25.605 39.215 26.015 ;
        RECT 38.250 24.605 39.280 25.605 ;
        RECT 39.850 24.625 40.225 32.410 ;
        RECT 40.500 32.025 42.180 33.260 ;
        RECT 43.015 32.025 47.940 32.035 ;
        RECT 40.500 31.545 47.940 32.025 ;
        RECT 40.500 29.285 42.180 31.545 ;
        RECT 43.015 31.125 47.940 31.545 ;
        RECT 42.520 30.935 42.775 30.960 ;
        RECT 42.520 30.920 42.795 30.935 ;
        RECT 42.490 30.645 42.825 30.920 ;
        RECT 43.000 30.895 48.000 31.125 ;
        RECT 48.210 30.935 48.465 30.960 ;
        RECT 42.520 30.630 42.775 30.645 ;
        RECT 43.000 30.455 48.000 30.685 ;
        RECT 48.205 30.645 48.465 30.935 ;
        RECT 48.210 30.630 48.465 30.645 ;
        RECT 43.045 30.445 47.900 30.455 ;
        RECT 43.045 28.920 45.690 28.925 ;
        RECT 41.720 28.720 45.690 28.920 ;
        RECT 41.720 28.690 45.680 28.720 ;
        RECT 40.560 28.335 40.895 28.610 ;
        RECT 41.440 28.440 41.670 28.485 ;
        RECT 36.420 24.560 36.775 24.580 ;
        RECT 36.420 24.490 36.650 24.560 ;
        RECT 37.560 24.490 37.790 24.580 ;
        RECT 38.320 24.465 39.230 24.605 ;
        RECT 39.850 24.490 40.240 24.625 ;
        RECT 38.310 24.285 39.320 24.465 ;
        RECT 34.410 24.055 36.370 24.285 ;
        RECT 37.840 24.055 39.800 24.285 ;
        RECT 35.115 23.005 35.465 24.055 ;
        RECT 37.865 24.050 39.750 24.055 ;
        RECT 40.045 22.355 40.240 24.490 ;
        RECT 40.630 22.830 40.820 28.335 ;
        RECT 41.250 27.105 41.670 28.440 ;
        RECT 42.975 27.105 44.320 28.690 ;
        RECT 41.250 25.720 44.320 27.105 ;
        RECT 41.250 24.990 41.670 25.720 ;
        RECT 41.245 24.485 41.670 24.990 ;
        RECT 40.630 22.640 40.945 22.830 ;
        RECT 30.950 22.125 34.910 22.355 ;
        RECT 36.380 22.125 40.340 22.355 ;
        RECT 40.755 22.130 40.945 22.640 ;
        RECT 30.670 21.515 30.900 21.965 ;
        RECT 32.150 21.515 32.940 22.125 ;
        RECT 30.670 21.210 32.940 21.515 ;
        RECT 30.615 21.195 32.940 21.210 ;
        RECT 30.530 20.350 32.940 21.195 ;
        RECT 30.530 19.975 30.900 20.350 ;
        RECT 30.670 19.965 30.900 19.975 ;
        RECT 32.150 19.805 32.940 20.350 ;
        RECT 34.960 21.880 35.190 21.965 ;
        RECT 36.100 21.880 36.330 21.965 ;
        RECT 34.960 20.055 36.330 21.880 ;
        RECT 34.960 19.965 35.190 20.055 ;
        RECT 30.950 19.575 34.910 19.805 ;
        RECT 27.890 19.255 30.085 19.280 ;
        RECT 30.530 19.255 30.755 19.265 ;
        RECT 35.430 19.255 35.920 20.055 ;
        RECT 36.100 19.965 36.330 20.055 ;
        RECT 37.815 21.745 39.155 22.125 ;
        RECT 40.390 21.745 40.620 21.965 ;
        RECT 37.815 20.150 40.620 21.745 ;
        RECT 37.815 19.805 39.155 20.150 ;
        RECT 40.390 19.965 40.620 20.150 ;
        RECT 36.380 19.575 40.340 19.805 ;
        RECT 40.770 19.785 40.945 22.130 ;
        RECT 41.245 21.965 41.540 24.485 ;
        RECT 42.975 24.280 44.320 25.720 ;
        RECT 45.730 28.390 45.960 28.485 ;
        RECT 46.205 28.390 46.695 30.445 ;
        RECT 47.265 28.920 47.900 28.925 ;
        RECT 47.150 28.690 51.110 28.920 ;
        RECT 46.870 28.390 47.100 28.485 ;
        RECT 45.730 24.565 47.100 28.390 ;
        RECT 45.730 24.485 45.960 24.565 ;
        RECT 46.870 24.485 47.100 24.565 ;
        RECT 48.525 24.280 49.870 28.690 ;
        RECT 51.160 28.420 51.390 28.485 ;
        RECT 52.045 28.425 52.520 33.260 ;
        RECT 53.845 32.455 54.525 33.260 ;
        RECT 55.390 33.180 57.990 33.260 ;
        RECT 54.945 32.735 55.280 32.985 ;
        RECT 54.960 32.710 55.250 32.735 ;
        RECT 58.420 32.635 60.330 33.260 ;
        RECT 62.420 32.925 64.305 32.930 ;
        RECT 65.865 32.925 67.750 32.930 ;
        RECT 62.410 32.695 64.370 32.925 ;
        RECT 65.840 32.695 67.800 32.925 ;
        RECT 54.770 32.455 55.000 32.505 ;
        RECT 53.845 31.955 55.000 32.455 ;
        RECT 52.915 28.735 53.250 28.985 ;
        RECT 52.935 28.705 53.225 28.735 ;
        RECT 52.745 28.425 52.975 28.500 ;
        RECT 51.160 24.485 51.615 28.420 ;
        RECT 52.045 27.680 52.975 28.425 ;
        RECT 52.380 24.565 52.975 27.680 ;
        RECT 52.745 24.500 52.975 24.565 ;
        RECT 53.185 28.475 53.415 28.500 ;
        RECT 53.185 24.920 53.695 28.475 ;
        RECT 53.185 24.550 53.880 24.920 ;
        RECT 54.380 24.600 55.000 31.955 ;
        RECT 53.185 24.500 53.415 24.550 ;
        RECT 41.720 24.250 45.680 24.280 ;
        RECT 47.150 24.250 51.110 24.280 ;
        RECT 41.720 24.090 51.110 24.250 ;
        RECT 41.720 24.050 45.680 24.090 ;
        RECT 47.150 24.050 51.110 24.090 ;
        RECT 51.275 22.660 51.615 24.485 ;
        RECT 52.925 22.660 53.345 24.305 ;
        RECT 51.275 22.505 53.345 22.660 ;
        RECT 51.350 22.390 53.345 22.505 ;
        RECT 41.810 22.125 45.770 22.355 ;
        RECT 47.240 22.125 51.200 22.355 ;
        RECT 41.245 21.205 41.760 21.965 ;
        RECT 41.315 20.025 41.760 21.205 ;
        RECT 41.530 19.965 41.760 20.025 ;
        RECT 43.190 19.805 44.145 22.125 ;
        RECT 45.820 21.900 46.050 21.965 ;
        RECT 46.960 21.900 47.190 21.965 ;
        RECT 45.820 20.030 47.190 21.900 ;
        RECT 45.820 19.965 46.050 20.030 ;
        RECT 40.755 19.255 40.945 19.785 ;
        RECT 41.810 19.575 45.770 19.805 ;
        RECT 46.225 19.255 46.780 20.030 ;
        RECT 46.960 19.965 47.190 20.030 ;
        RECT 48.635 19.805 49.590 22.125 ;
        RECT 51.350 21.970 51.615 22.390 ;
        RECT 52.925 22.115 53.345 22.390 ;
        RECT 53.580 23.355 53.880 24.550 ;
        RECT 54.770 24.505 55.000 24.600 ;
        RECT 55.210 32.430 55.440 32.505 ;
        RECT 55.210 25.110 55.985 32.430 ;
        RECT 58.385 32.405 60.385 32.635 ;
        RECT 62.130 32.410 62.360 32.490 ;
        RECT 57.950 29.060 58.180 32.355 ;
        RECT 60.590 32.275 60.820 32.355 ;
        RECT 60.560 29.060 60.820 32.275 ;
        RECT 57.950 27.245 60.820 29.060 ;
        RECT 55.210 24.580 56.060 25.110 ;
        RECT 57.950 24.825 58.180 27.245 ;
        RECT 55.210 24.505 55.440 24.580 ;
        RECT 54.875 23.825 55.390 24.315 ;
        RECT 54.875 23.360 55.385 23.825 ;
        RECT 55.690 23.795 56.060 24.580 ;
        RECT 57.590 24.395 58.180 24.825 ;
        RECT 59.075 24.640 59.335 24.960 ;
        RECT 60.560 24.645 60.820 27.245 ;
        RECT 61.890 24.990 62.360 32.410 ;
        RECT 62.850 25.775 63.740 32.695 ;
        RECT 64.420 32.390 64.650 32.490 ;
        RECT 64.420 32.380 64.775 32.390 ;
        RECT 65.560 32.380 65.790 32.490 ;
        RECT 59.130 24.480 59.280 24.640 ;
        RECT 54.510 23.355 55.385 23.360 ;
        RECT 53.580 22.950 55.385 23.355 ;
        RECT 53.580 22.110 53.880 22.950 ;
        RECT 54.510 22.935 55.385 22.950 ;
        RECT 54.875 22.825 55.385 22.935 ;
        RECT 54.875 22.125 55.390 22.825 ;
        RECT 55.585 22.795 56.615 23.795 ;
        RECT 51.275 21.965 51.615 21.970 ;
        RECT 51.250 20.020 51.615 21.965 ;
        RECT 52.830 21.900 53.060 21.970 ;
        RECT 52.335 21.230 53.060 21.900 ;
        RECT 52.325 21.040 53.060 21.230 ;
        RECT 52.325 20.240 52.680 21.040 ;
        RECT 52.830 20.970 53.060 21.040 ;
        RECT 53.270 21.925 53.500 21.970 ;
        RECT 53.640 21.925 53.880 22.110 ;
        RECT 53.270 21.595 53.880 21.925 ;
        RECT 54.855 21.870 55.085 21.975 ;
        RECT 53.270 21.040 53.765 21.595 ;
        RECT 53.270 20.970 53.500 21.040 ;
        RECT 53.020 20.785 53.310 20.810 ;
        RECT 53.005 20.535 53.340 20.785 ;
        RECT 54.625 20.765 55.085 21.870 ;
        RECT 54.305 20.240 55.085 20.765 ;
        RECT 51.885 20.060 55.085 20.240 ;
        RECT 51.250 19.965 51.480 20.020 ;
        RECT 47.240 19.575 51.200 19.805 ;
        RECT 51.885 19.620 54.690 20.060 ;
        RECT 54.855 19.975 55.085 20.060 ;
        RECT 55.295 21.910 55.525 21.975 ;
        RECT 55.690 21.910 56.060 22.795 ;
        RECT 55.295 21.585 56.060 21.910 ;
        RECT 55.295 20.045 56.055 21.585 ;
        RECT 55.295 19.975 55.525 20.045 ;
        RECT 55.045 19.795 55.335 19.815 ;
        RECT 51.885 19.255 54.350 19.620 ;
        RECT 55.020 19.545 55.355 19.795 ;
        RECT 57.590 19.280 58.085 24.395 ;
        RECT 59.105 24.345 59.310 24.480 ;
        RECT 60.590 24.395 60.820 24.645 ;
        RECT 61.610 24.550 62.360 24.990 ;
        RECT 62.780 24.775 63.795 25.775 ;
        RECT 58.385 24.115 60.385 24.345 ;
        RECT 61.610 22.355 61.980 24.550 ;
        RECT 62.130 24.490 62.360 24.550 ;
        RECT 62.850 24.285 63.740 24.775 ;
        RECT 64.420 24.580 65.790 32.380 ;
        RECT 66.325 27.635 67.215 32.695 ;
        RECT 67.850 32.410 68.080 32.490 ;
        RECT 66.320 26.015 67.220 27.635 ;
        RECT 66.325 25.605 67.215 26.015 ;
        RECT 66.250 24.605 67.280 25.605 ;
        RECT 67.850 24.625 68.225 32.410 ;
        RECT 68.500 32.025 70.180 33.260 ;
        RECT 71.015 32.025 75.940 32.035 ;
        RECT 68.500 31.545 75.940 32.025 ;
        RECT 68.500 29.285 70.180 31.545 ;
        RECT 71.015 31.125 75.940 31.545 ;
        RECT 70.520 30.935 70.775 30.960 ;
        RECT 70.520 30.920 70.795 30.935 ;
        RECT 70.490 30.645 70.825 30.920 ;
        RECT 71.000 30.895 76.000 31.125 ;
        RECT 76.210 30.935 76.465 30.960 ;
        RECT 70.520 30.630 70.775 30.645 ;
        RECT 71.000 30.455 76.000 30.685 ;
        RECT 76.205 30.645 76.465 30.935 ;
        RECT 76.210 30.630 76.465 30.645 ;
        RECT 71.045 30.445 75.900 30.455 ;
        RECT 71.045 28.920 73.690 28.925 ;
        RECT 69.720 28.720 73.690 28.920 ;
        RECT 69.720 28.690 73.680 28.720 ;
        RECT 68.560 28.335 68.895 28.610 ;
        RECT 69.440 28.440 69.670 28.485 ;
        RECT 64.420 24.560 64.775 24.580 ;
        RECT 64.420 24.490 64.650 24.560 ;
        RECT 65.560 24.490 65.790 24.580 ;
        RECT 66.320 24.465 67.230 24.605 ;
        RECT 67.850 24.490 68.240 24.625 ;
        RECT 66.310 24.285 67.320 24.465 ;
        RECT 62.410 24.055 64.370 24.285 ;
        RECT 65.840 24.055 67.800 24.285 ;
        RECT 63.165 23.050 63.510 24.055 ;
        RECT 65.865 24.050 67.750 24.055 ;
        RECT 68.045 22.355 68.240 24.490 ;
        RECT 68.630 22.830 68.820 28.335 ;
        RECT 69.250 27.105 69.670 28.440 ;
        RECT 70.975 27.105 72.320 28.690 ;
        RECT 69.250 25.720 72.320 27.105 ;
        RECT 69.250 24.990 69.670 25.720 ;
        RECT 69.245 24.485 69.670 24.990 ;
        RECT 68.630 22.640 68.945 22.830 ;
        RECT 58.950 22.125 62.910 22.355 ;
        RECT 64.380 22.125 68.340 22.355 ;
        RECT 68.755 22.130 68.945 22.640 ;
        RECT 58.670 21.515 58.900 21.965 ;
        RECT 60.150 21.515 60.940 22.125 ;
        RECT 58.670 21.210 60.940 21.515 ;
        RECT 58.615 21.195 60.940 21.210 ;
        RECT 58.530 20.350 60.940 21.195 ;
        RECT 58.530 19.975 58.900 20.350 ;
        RECT 58.670 19.965 58.900 19.975 ;
        RECT 60.150 19.805 60.940 20.350 ;
        RECT 62.960 21.880 63.190 21.965 ;
        RECT 64.100 21.880 64.330 21.965 ;
        RECT 62.960 20.055 64.330 21.880 ;
        RECT 62.960 19.965 63.190 20.055 ;
        RECT 58.950 19.575 62.910 19.805 ;
        RECT 55.490 19.255 58.085 19.280 ;
        RECT 58.530 19.255 58.755 19.265 ;
        RECT 63.430 19.255 63.920 20.055 ;
        RECT 64.100 19.965 64.330 20.055 ;
        RECT 65.815 21.745 67.155 22.125 ;
        RECT 68.390 21.745 68.620 21.965 ;
        RECT 65.815 20.150 68.620 21.745 ;
        RECT 65.815 19.805 67.155 20.150 ;
        RECT 68.390 19.965 68.620 20.150 ;
        RECT 64.380 19.575 68.340 19.805 ;
        RECT 68.770 19.785 68.945 22.130 ;
        RECT 69.245 21.965 69.540 24.485 ;
        RECT 70.975 24.280 72.320 25.720 ;
        RECT 73.730 28.390 73.960 28.485 ;
        RECT 74.205 28.390 74.695 30.445 ;
        RECT 75.265 28.920 75.900 28.925 ;
        RECT 75.150 28.690 79.110 28.920 ;
        RECT 74.870 28.390 75.100 28.485 ;
        RECT 73.730 24.565 75.100 28.390 ;
        RECT 73.730 24.485 73.960 24.565 ;
        RECT 74.870 24.485 75.100 24.565 ;
        RECT 76.525 24.280 77.870 28.690 ;
        RECT 79.160 28.420 79.390 28.485 ;
        RECT 80.045 28.425 80.520 33.260 ;
        RECT 81.845 32.455 82.525 33.260 ;
        RECT 82.945 32.735 83.280 32.985 ;
        RECT 82.960 32.710 83.250 32.735 ;
        RECT 86.420 32.635 88.330 33.260 ;
        RECT 90.420 32.925 92.305 32.930 ;
        RECT 93.865 32.925 95.750 32.930 ;
        RECT 90.410 32.695 92.370 32.925 ;
        RECT 93.840 32.695 95.800 32.925 ;
        RECT 82.770 32.455 83.000 32.505 ;
        RECT 81.845 31.955 83.000 32.455 ;
        RECT 80.915 28.735 81.250 28.985 ;
        RECT 80.935 28.705 81.225 28.735 ;
        RECT 80.745 28.425 80.975 28.500 ;
        RECT 79.160 24.485 79.615 28.420 ;
        RECT 80.045 27.680 80.975 28.425 ;
        RECT 80.380 24.565 80.975 27.680 ;
        RECT 80.745 24.500 80.975 24.565 ;
        RECT 81.185 28.475 81.415 28.500 ;
        RECT 81.185 24.920 81.695 28.475 ;
        RECT 81.185 24.550 81.880 24.920 ;
        RECT 82.380 24.600 83.000 31.955 ;
        RECT 81.185 24.500 81.415 24.550 ;
        RECT 69.720 24.250 73.680 24.280 ;
        RECT 75.150 24.250 79.110 24.280 ;
        RECT 69.720 24.090 79.110 24.250 ;
        RECT 69.720 24.050 73.680 24.090 ;
        RECT 75.150 24.050 79.110 24.090 ;
        RECT 79.275 22.660 79.615 24.485 ;
        RECT 80.925 22.660 81.345 24.305 ;
        RECT 79.275 22.505 81.345 22.660 ;
        RECT 79.350 22.390 81.345 22.505 ;
        RECT 69.810 22.125 73.770 22.355 ;
        RECT 75.240 22.125 79.200 22.355 ;
        RECT 69.245 21.205 69.760 21.965 ;
        RECT 69.315 20.025 69.760 21.205 ;
        RECT 69.530 19.965 69.760 20.025 ;
        RECT 71.190 19.805 72.145 22.125 ;
        RECT 73.820 21.900 74.050 21.965 ;
        RECT 74.960 21.900 75.190 21.965 ;
        RECT 73.820 20.030 75.190 21.900 ;
        RECT 73.820 19.965 74.050 20.030 ;
        RECT 68.755 19.255 68.945 19.785 ;
        RECT 69.810 19.575 73.770 19.805 ;
        RECT 74.225 19.255 74.780 20.030 ;
        RECT 74.960 19.965 75.190 20.030 ;
        RECT 76.635 19.805 77.590 22.125 ;
        RECT 79.350 21.970 79.615 22.390 ;
        RECT 80.925 22.115 81.345 22.390 ;
        RECT 81.580 23.355 81.880 24.550 ;
        RECT 82.770 24.505 83.000 24.600 ;
        RECT 83.210 32.430 83.440 32.505 ;
        RECT 83.210 25.110 83.985 32.430 ;
        RECT 86.385 32.405 88.385 32.635 ;
        RECT 90.130 32.410 90.360 32.490 ;
        RECT 85.950 29.060 86.180 32.355 ;
        RECT 88.590 32.275 88.820 32.355 ;
        RECT 88.560 29.060 88.820 32.275 ;
        RECT 85.950 27.245 88.820 29.060 ;
        RECT 83.210 24.580 84.060 25.110 ;
        RECT 85.950 24.825 86.180 27.245 ;
        RECT 83.210 24.505 83.440 24.580 ;
        RECT 82.875 23.825 83.390 24.315 ;
        RECT 82.875 23.360 83.385 23.825 ;
        RECT 83.690 23.795 84.060 24.580 ;
        RECT 85.590 24.395 86.180 24.825 ;
        RECT 87.075 24.640 87.335 24.960 ;
        RECT 88.560 24.645 88.820 27.245 ;
        RECT 89.890 24.990 90.360 32.410 ;
        RECT 90.850 25.775 91.740 32.695 ;
        RECT 92.420 32.390 92.650 32.490 ;
        RECT 92.420 32.380 92.775 32.390 ;
        RECT 93.560 32.380 93.790 32.490 ;
        RECT 87.130 24.480 87.280 24.640 ;
        RECT 82.510 23.355 83.385 23.360 ;
        RECT 81.580 22.950 83.385 23.355 ;
        RECT 81.580 22.110 81.880 22.950 ;
        RECT 82.510 22.935 83.385 22.950 ;
        RECT 82.875 22.825 83.385 22.935 ;
        RECT 82.875 22.125 83.390 22.825 ;
        RECT 83.615 22.795 84.645 23.795 ;
        RECT 79.275 21.965 79.615 21.970 ;
        RECT 79.250 20.020 79.615 21.965 ;
        RECT 80.830 21.900 81.060 21.970 ;
        RECT 80.335 21.230 81.060 21.900 ;
        RECT 80.325 21.040 81.060 21.230 ;
        RECT 80.325 20.240 80.680 21.040 ;
        RECT 80.830 20.970 81.060 21.040 ;
        RECT 81.270 21.925 81.500 21.970 ;
        RECT 81.640 21.925 81.880 22.110 ;
        RECT 81.270 21.595 81.880 21.925 ;
        RECT 82.855 21.870 83.085 21.975 ;
        RECT 81.270 21.040 81.765 21.595 ;
        RECT 81.270 20.970 81.500 21.040 ;
        RECT 81.020 20.785 81.310 20.810 ;
        RECT 81.005 20.535 81.340 20.785 ;
        RECT 82.625 20.765 83.085 21.870 ;
        RECT 82.305 20.240 83.085 20.765 ;
        RECT 79.885 20.060 83.085 20.240 ;
        RECT 79.250 19.965 79.480 20.020 ;
        RECT 75.240 19.575 79.200 19.805 ;
        RECT 79.885 19.620 82.690 20.060 ;
        RECT 82.855 19.975 83.085 20.060 ;
        RECT 83.295 21.910 83.525 21.975 ;
        RECT 83.690 21.910 84.060 22.795 ;
        RECT 83.295 21.585 84.060 21.910 ;
        RECT 83.295 20.045 84.055 21.585 ;
        RECT 83.295 19.975 83.525 20.045 ;
        RECT 83.045 19.795 83.335 19.815 ;
        RECT 79.885 19.255 82.350 19.620 ;
        RECT 83.020 19.545 83.355 19.795 ;
        RECT 85.590 19.280 86.085 24.395 ;
        RECT 87.105 24.345 87.310 24.480 ;
        RECT 88.590 24.395 88.820 24.645 ;
        RECT 89.610 24.550 90.360 24.990 ;
        RECT 90.780 24.775 91.795 25.775 ;
        RECT 86.385 24.115 88.385 24.345 ;
        RECT 89.610 22.355 89.980 24.550 ;
        RECT 90.130 24.490 90.360 24.550 ;
        RECT 90.850 24.285 91.740 24.775 ;
        RECT 92.420 24.580 93.790 32.380 ;
        RECT 94.325 27.635 95.215 32.695 ;
        RECT 95.850 32.410 96.080 32.490 ;
        RECT 94.320 26.015 95.220 27.635 ;
        RECT 94.325 25.605 95.215 26.015 ;
        RECT 94.250 24.605 95.280 25.605 ;
        RECT 95.850 24.625 96.225 32.410 ;
        RECT 96.500 32.025 98.180 33.260 ;
        RECT 99.015 32.025 103.940 32.035 ;
        RECT 96.500 31.545 103.940 32.025 ;
        RECT 96.500 29.285 98.180 31.545 ;
        RECT 99.015 31.125 103.940 31.545 ;
        RECT 98.520 30.935 98.775 30.960 ;
        RECT 98.520 30.920 98.795 30.935 ;
        RECT 98.490 30.645 98.825 30.920 ;
        RECT 99.000 30.895 104.000 31.125 ;
        RECT 104.210 30.935 104.465 30.960 ;
        RECT 98.520 30.630 98.775 30.645 ;
        RECT 99.000 30.455 104.000 30.685 ;
        RECT 104.205 30.645 104.465 30.935 ;
        RECT 104.210 30.630 104.465 30.645 ;
        RECT 99.045 30.445 103.900 30.455 ;
        RECT 99.045 28.920 101.690 28.925 ;
        RECT 97.720 28.720 101.690 28.920 ;
        RECT 97.720 28.690 101.680 28.720 ;
        RECT 96.560 28.335 96.895 28.610 ;
        RECT 97.440 28.440 97.670 28.485 ;
        RECT 92.420 24.560 92.775 24.580 ;
        RECT 92.420 24.490 92.650 24.560 ;
        RECT 93.560 24.490 93.790 24.580 ;
        RECT 94.320 24.465 95.230 24.605 ;
        RECT 95.850 24.490 96.240 24.625 ;
        RECT 94.310 24.285 95.320 24.465 ;
        RECT 90.410 24.055 92.370 24.285 ;
        RECT 93.840 24.055 95.800 24.285 ;
        RECT 91.125 22.980 91.525 24.055 ;
        RECT 93.865 24.050 95.750 24.055 ;
        RECT 96.045 22.355 96.240 24.490 ;
        RECT 96.630 22.830 96.820 28.335 ;
        RECT 97.250 27.105 97.670 28.440 ;
        RECT 98.975 27.105 100.320 28.690 ;
        RECT 97.250 25.720 100.320 27.105 ;
        RECT 97.250 24.990 97.670 25.720 ;
        RECT 97.245 24.485 97.670 24.990 ;
        RECT 96.630 22.640 96.945 22.830 ;
        RECT 86.950 22.125 90.910 22.355 ;
        RECT 92.380 22.125 96.340 22.355 ;
        RECT 96.755 22.130 96.945 22.640 ;
        RECT 86.670 21.515 86.900 21.965 ;
        RECT 88.150 21.515 88.940 22.125 ;
        RECT 86.670 21.210 88.940 21.515 ;
        RECT 86.615 21.195 88.940 21.210 ;
        RECT 86.530 20.350 88.940 21.195 ;
        RECT 86.530 19.975 86.900 20.350 ;
        RECT 86.670 19.965 86.900 19.975 ;
        RECT 88.150 19.805 88.940 20.350 ;
        RECT 90.960 21.880 91.190 21.965 ;
        RECT 92.100 21.880 92.330 21.965 ;
        RECT 90.960 20.055 92.330 21.880 ;
        RECT 90.960 19.965 91.190 20.055 ;
        RECT 86.950 19.575 90.910 19.805 ;
        RECT 83.790 19.255 86.085 19.280 ;
        RECT 86.530 19.255 86.755 19.265 ;
        RECT 91.430 19.255 91.920 20.055 ;
        RECT 92.100 19.965 92.330 20.055 ;
        RECT 93.815 21.745 95.155 22.125 ;
        RECT 96.390 21.745 96.620 21.965 ;
        RECT 93.815 20.150 96.620 21.745 ;
        RECT 93.815 19.805 95.155 20.150 ;
        RECT 96.390 19.965 96.620 20.150 ;
        RECT 92.380 19.575 96.340 19.805 ;
        RECT 96.770 19.785 96.945 22.130 ;
        RECT 97.245 21.965 97.540 24.485 ;
        RECT 98.975 24.280 100.320 25.720 ;
        RECT 101.730 28.390 101.960 28.485 ;
        RECT 102.205 28.390 102.695 30.445 ;
        RECT 103.265 28.920 103.900 28.925 ;
        RECT 103.150 28.690 107.110 28.920 ;
        RECT 102.870 28.390 103.100 28.485 ;
        RECT 101.730 24.565 103.100 28.390 ;
        RECT 101.730 24.485 101.960 24.565 ;
        RECT 102.870 24.485 103.100 24.565 ;
        RECT 104.525 24.280 105.870 28.690 ;
        RECT 107.160 28.420 107.390 28.485 ;
        RECT 108.045 28.425 108.520 33.260 ;
        RECT 109.845 32.455 110.525 33.260 ;
        RECT 110.945 32.735 111.280 32.985 ;
        RECT 110.960 32.710 111.250 32.735 ;
        RECT 114.420 32.635 116.330 33.260 ;
        RECT 118.420 32.925 120.305 32.930 ;
        RECT 121.865 32.925 123.750 32.930 ;
        RECT 118.410 32.695 120.370 32.925 ;
        RECT 121.840 32.695 123.800 32.925 ;
        RECT 110.770 32.455 111.000 32.505 ;
        RECT 109.845 31.955 111.000 32.455 ;
        RECT 108.915 28.735 109.250 28.985 ;
        RECT 108.935 28.705 109.225 28.735 ;
        RECT 108.745 28.425 108.975 28.500 ;
        RECT 107.160 24.485 107.615 28.420 ;
        RECT 108.045 27.680 108.975 28.425 ;
        RECT 108.380 24.565 108.975 27.680 ;
        RECT 108.745 24.500 108.975 24.565 ;
        RECT 109.185 28.475 109.415 28.500 ;
        RECT 109.185 24.920 109.695 28.475 ;
        RECT 109.185 24.550 109.880 24.920 ;
        RECT 110.380 24.600 111.000 31.955 ;
        RECT 109.185 24.500 109.415 24.550 ;
        RECT 97.720 24.250 101.680 24.280 ;
        RECT 103.150 24.250 107.110 24.280 ;
        RECT 97.720 24.090 107.110 24.250 ;
        RECT 97.720 24.050 101.680 24.090 ;
        RECT 103.150 24.050 107.110 24.090 ;
        RECT 107.275 22.660 107.615 24.485 ;
        RECT 108.925 22.660 109.345 24.305 ;
        RECT 107.275 22.505 109.345 22.660 ;
        RECT 107.350 22.390 109.345 22.505 ;
        RECT 97.810 22.125 101.770 22.355 ;
        RECT 103.240 22.125 107.200 22.355 ;
        RECT 97.245 21.205 97.760 21.965 ;
        RECT 97.315 20.025 97.760 21.205 ;
        RECT 97.530 19.965 97.760 20.025 ;
        RECT 99.190 19.805 100.145 22.125 ;
        RECT 101.820 21.900 102.050 21.965 ;
        RECT 102.960 21.900 103.190 21.965 ;
        RECT 101.820 20.030 103.190 21.900 ;
        RECT 101.820 19.965 102.050 20.030 ;
        RECT 96.755 19.255 96.945 19.785 ;
        RECT 97.810 19.575 101.770 19.805 ;
        RECT 102.225 19.255 102.780 20.030 ;
        RECT 102.960 19.965 103.190 20.030 ;
        RECT 104.635 19.805 105.590 22.125 ;
        RECT 107.350 21.970 107.615 22.390 ;
        RECT 108.925 22.115 109.345 22.390 ;
        RECT 109.580 23.355 109.880 24.550 ;
        RECT 110.770 24.505 111.000 24.600 ;
        RECT 111.210 32.430 111.440 32.505 ;
        RECT 111.210 25.110 111.985 32.430 ;
        RECT 114.385 32.405 116.385 32.635 ;
        RECT 118.130 32.410 118.360 32.490 ;
        RECT 113.950 29.060 114.180 32.355 ;
        RECT 116.590 32.275 116.820 32.355 ;
        RECT 116.560 29.060 116.820 32.275 ;
        RECT 113.950 27.245 116.820 29.060 ;
        RECT 111.210 24.580 112.060 25.110 ;
        RECT 113.950 24.825 114.180 27.245 ;
        RECT 111.210 24.505 111.440 24.580 ;
        RECT 110.875 23.825 111.390 24.315 ;
        RECT 110.875 23.360 111.385 23.825 ;
        RECT 111.690 23.795 112.060 24.580 ;
        RECT 113.590 24.395 114.180 24.825 ;
        RECT 115.075 24.640 115.335 24.960 ;
        RECT 116.560 24.645 116.820 27.245 ;
        RECT 117.890 24.990 118.360 32.410 ;
        RECT 118.850 25.775 119.740 32.695 ;
        RECT 120.420 32.390 120.650 32.490 ;
        RECT 120.420 32.380 120.775 32.390 ;
        RECT 121.560 32.380 121.790 32.490 ;
        RECT 115.130 24.480 115.280 24.640 ;
        RECT 110.510 23.355 111.385 23.360 ;
        RECT 109.580 22.950 111.385 23.355 ;
        RECT 109.580 22.110 109.880 22.950 ;
        RECT 110.510 22.935 111.385 22.950 ;
        RECT 110.875 22.825 111.385 22.935 ;
        RECT 110.875 22.125 111.390 22.825 ;
        RECT 111.585 22.795 112.615 23.795 ;
        RECT 107.275 21.965 107.615 21.970 ;
        RECT 107.250 20.020 107.615 21.965 ;
        RECT 108.830 21.900 109.060 21.970 ;
        RECT 108.335 21.230 109.060 21.900 ;
        RECT 108.325 21.040 109.060 21.230 ;
        RECT 108.325 20.240 108.680 21.040 ;
        RECT 108.830 20.970 109.060 21.040 ;
        RECT 109.270 21.925 109.500 21.970 ;
        RECT 109.640 21.925 109.880 22.110 ;
        RECT 109.270 21.595 109.880 21.925 ;
        RECT 110.855 21.870 111.085 21.975 ;
        RECT 109.270 21.040 109.765 21.595 ;
        RECT 109.270 20.970 109.500 21.040 ;
        RECT 109.020 20.785 109.310 20.810 ;
        RECT 109.005 20.535 109.340 20.785 ;
        RECT 110.625 20.765 111.085 21.870 ;
        RECT 110.305 20.240 111.085 20.765 ;
        RECT 107.885 20.060 111.085 20.240 ;
        RECT 107.250 19.965 107.480 20.020 ;
        RECT 103.240 19.575 107.200 19.805 ;
        RECT 107.885 19.620 110.690 20.060 ;
        RECT 110.855 19.975 111.085 20.060 ;
        RECT 111.295 21.910 111.525 21.975 ;
        RECT 111.690 21.910 112.060 22.795 ;
        RECT 111.295 21.585 112.060 21.910 ;
        RECT 111.295 20.045 112.055 21.585 ;
        RECT 111.295 19.975 111.525 20.045 ;
        RECT 111.045 19.795 111.335 19.815 ;
        RECT 107.885 19.255 110.350 19.620 ;
        RECT 111.020 19.545 111.355 19.795 ;
        RECT 113.590 19.255 114.085 24.395 ;
        RECT 115.105 24.345 115.310 24.480 ;
        RECT 116.590 24.395 116.820 24.645 ;
        RECT 117.610 24.550 118.360 24.990 ;
        RECT 118.780 24.775 119.795 25.775 ;
        RECT 114.385 24.115 116.385 24.345 ;
        RECT 117.610 22.355 117.980 24.550 ;
        RECT 118.130 24.490 118.360 24.550 ;
        RECT 118.850 24.285 119.740 24.775 ;
        RECT 120.420 24.580 121.790 32.380 ;
        RECT 122.325 27.635 123.215 32.695 ;
        RECT 123.850 32.410 124.080 32.490 ;
        RECT 122.320 26.015 123.220 27.635 ;
        RECT 122.325 25.605 123.215 26.015 ;
        RECT 122.250 24.605 123.280 25.605 ;
        RECT 123.850 24.625 124.225 32.410 ;
        RECT 124.500 32.025 126.180 33.260 ;
        RECT 127.015 32.025 131.940 32.035 ;
        RECT 124.500 31.545 131.940 32.025 ;
        RECT 124.500 29.285 126.180 31.545 ;
        RECT 127.015 31.125 131.940 31.545 ;
        RECT 126.520 30.935 126.775 30.960 ;
        RECT 126.520 30.920 126.795 30.935 ;
        RECT 126.490 30.645 126.825 30.920 ;
        RECT 127.000 30.895 132.000 31.125 ;
        RECT 132.210 30.935 132.465 30.960 ;
        RECT 126.520 30.630 126.775 30.645 ;
        RECT 127.000 30.455 132.000 30.685 ;
        RECT 132.205 30.645 132.465 30.935 ;
        RECT 132.210 30.630 132.465 30.645 ;
        RECT 127.045 30.445 131.900 30.455 ;
        RECT 127.045 28.920 129.690 28.925 ;
        RECT 125.720 28.720 129.690 28.920 ;
        RECT 125.720 28.690 129.680 28.720 ;
        RECT 124.560 28.335 124.895 28.610 ;
        RECT 125.440 28.440 125.670 28.485 ;
        RECT 120.420 24.560 120.775 24.580 ;
        RECT 120.420 24.490 120.650 24.560 ;
        RECT 121.560 24.490 121.790 24.580 ;
        RECT 122.320 24.465 123.230 24.605 ;
        RECT 123.850 24.490 124.240 24.625 ;
        RECT 122.310 24.285 123.320 24.465 ;
        RECT 118.410 24.055 120.370 24.285 ;
        RECT 121.840 24.055 123.800 24.285 ;
        RECT 119.160 23.115 119.445 24.055 ;
        RECT 121.865 24.050 123.750 24.055 ;
        RECT 124.045 22.355 124.240 24.490 ;
        RECT 124.630 22.830 124.820 28.335 ;
        RECT 125.250 27.105 125.670 28.440 ;
        RECT 126.975 27.105 128.320 28.690 ;
        RECT 125.250 25.720 128.320 27.105 ;
        RECT 125.250 24.990 125.670 25.720 ;
        RECT 125.245 24.485 125.670 24.990 ;
        RECT 124.630 22.640 124.945 22.830 ;
        RECT 114.950 22.125 118.910 22.355 ;
        RECT 120.380 22.125 124.340 22.355 ;
        RECT 124.755 22.130 124.945 22.640 ;
        RECT 114.670 21.515 114.900 21.965 ;
        RECT 116.150 21.515 116.940 22.125 ;
        RECT 114.670 21.210 116.940 21.515 ;
        RECT 114.615 21.195 116.940 21.210 ;
        RECT 114.530 20.350 116.940 21.195 ;
        RECT 114.530 19.975 114.900 20.350 ;
        RECT 114.670 19.965 114.900 19.975 ;
        RECT 116.150 19.805 116.940 20.350 ;
        RECT 118.960 21.880 119.190 21.965 ;
        RECT 120.100 21.880 120.330 21.965 ;
        RECT 118.960 20.055 120.330 21.880 ;
        RECT 118.960 19.965 119.190 20.055 ;
        RECT 114.950 19.575 118.910 19.805 ;
        RECT 114.530 19.255 114.755 19.265 ;
        RECT 119.430 19.255 119.920 20.055 ;
        RECT 120.100 19.965 120.330 20.055 ;
        RECT 121.815 21.745 123.155 22.125 ;
        RECT 124.390 21.745 124.620 21.965 ;
        RECT 121.815 20.150 124.620 21.745 ;
        RECT 121.815 19.805 123.155 20.150 ;
        RECT 124.390 19.965 124.620 20.150 ;
        RECT 120.380 19.575 124.340 19.805 ;
        RECT 124.770 19.785 124.945 22.130 ;
        RECT 125.245 21.965 125.540 24.485 ;
        RECT 126.975 24.280 128.320 25.720 ;
        RECT 129.730 28.390 129.960 28.485 ;
        RECT 130.205 28.390 130.695 30.445 ;
        RECT 131.265 28.920 131.900 28.925 ;
        RECT 131.150 28.690 135.110 28.920 ;
        RECT 130.870 28.390 131.100 28.485 ;
        RECT 129.730 24.565 131.100 28.390 ;
        RECT 129.730 24.485 129.960 24.565 ;
        RECT 130.870 24.485 131.100 24.565 ;
        RECT 132.525 24.280 133.870 28.690 ;
        RECT 135.160 28.420 135.390 28.485 ;
        RECT 136.045 28.425 136.520 33.260 ;
        RECT 137.845 32.455 138.525 33.260 ;
        RECT 138.945 32.735 139.280 32.985 ;
        RECT 138.960 32.710 139.250 32.735 ;
        RECT 138.770 32.455 139.000 32.505 ;
        RECT 137.845 31.955 139.000 32.455 ;
        RECT 136.915 28.735 137.250 28.985 ;
        RECT 136.935 28.705 137.225 28.735 ;
        RECT 136.745 28.425 136.975 28.500 ;
        RECT 135.160 24.485 135.615 28.420 ;
        RECT 136.045 27.680 136.975 28.425 ;
        RECT 136.380 24.565 136.975 27.680 ;
        RECT 136.745 24.500 136.975 24.565 ;
        RECT 137.185 28.475 137.415 28.500 ;
        RECT 137.185 24.920 137.695 28.475 ;
        RECT 137.185 24.550 137.880 24.920 ;
        RECT 138.380 24.600 139.000 31.955 ;
        RECT 137.185 24.500 137.415 24.550 ;
        RECT 125.720 24.250 129.680 24.280 ;
        RECT 131.150 24.250 135.110 24.280 ;
        RECT 125.720 24.090 135.110 24.250 ;
        RECT 125.720 24.050 129.680 24.090 ;
        RECT 131.150 24.050 135.110 24.090 ;
        RECT 135.275 22.660 135.615 24.485 ;
        RECT 136.925 22.660 137.345 24.305 ;
        RECT 135.275 22.505 137.345 22.660 ;
        RECT 135.350 22.390 137.345 22.505 ;
        RECT 125.810 22.125 129.770 22.355 ;
        RECT 131.240 22.125 135.200 22.355 ;
        RECT 125.245 21.205 125.760 21.965 ;
        RECT 125.315 20.025 125.760 21.205 ;
        RECT 125.530 19.965 125.760 20.025 ;
        RECT 127.190 19.805 128.145 22.125 ;
        RECT 129.820 21.900 130.050 21.965 ;
        RECT 130.960 21.900 131.190 21.965 ;
        RECT 129.820 20.030 131.190 21.900 ;
        RECT 129.820 19.965 130.050 20.030 ;
        RECT 124.755 19.255 124.945 19.785 ;
        RECT 125.810 19.575 129.770 19.805 ;
        RECT 130.225 19.255 130.780 20.030 ;
        RECT 130.960 19.965 131.190 20.030 ;
        RECT 132.635 19.805 133.590 22.125 ;
        RECT 135.350 21.970 135.615 22.390 ;
        RECT 136.925 22.115 137.345 22.390 ;
        RECT 137.580 23.355 137.880 24.550 ;
        RECT 138.770 24.505 139.000 24.600 ;
        RECT 139.210 32.430 139.440 32.505 ;
        RECT 139.210 25.110 139.985 32.430 ;
        RECT 139.210 24.580 140.060 25.110 ;
        RECT 139.210 24.505 139.440 24.580 ;
        RECT 138.875 23.825 139.390 24.315 ;
        RECT 138.875 23.360 139.385 23.825 ;
        RECT 139.690 23.795 140.060 24.580 ;
        RECT 138.510 23.355 139.385 23.360 ;
        RECT 137.580 22.950 139.385 23.355 ;
        RECT 137.580 22.110 137.880 22.950 ;
        RECT 138.510 22.935 139.385 22.950 ;
        RECT 138.875 22.825 139.385 22.935 ;
        RECT 138.875 22.125 139.390 22.825 ;
        RECT 139.615 22.795 140.645 23.795 ;
        RECT 135.275 21.965 135.615 21.970 ;
        RECT 135.250 20.020 135.615 21.965 ;
        RECT 136.830 21.900 137.060 21.970 ;
        RECT 136.335 21.230 137.060 21.900 ;
        RECT 136.325 21.040 137.060 21.230 ;
        RECT 136.325 20.240 136.680 21.040 ;
        RECT 136.830 20.970 137.060 21.040 ;
        RECT 137.270 21.925 137.500 21.970 ;
        RECT 137.640 21.925 137.880 22.110 ;
        RECT 137.270 21.595 137.880 21.925 ;
        RECT 138.855 21.870 139.085 21.975 ;
        RECT 137.270 21.040 137.765 21.595 ;
        RECT 137.270 20.970 137.500 21.040 ;
        RECT 137.020 20.785 137.310 20.810 ;
        RECT 137.005 20.535 137.340 20.785 ;
        RECT 138.625 20.765 139.085 21.870 ;
        RECT 138.305 20.240 139.085 20.765 ;
        RECT 135.885 20.060 139.085 20.240 ;
        RECT 135.250 19.965 135.480 20.020 ;
        RECT 131.240 19.575 135.200 19.805 ;
        RECT 135.885 19.620 138.690 20.060 ;
        RECT 138.855 19.975 139.085 20.060 ;
        RECT 139.295 21.910 139.525 21.975 ;
        RECT 139.690 21.910 140.060 22.795 ;
        RECT 139.295 21.585 140.060 21.910 ;
        RECT 139.295 20.045 140.055 21.585 ;
        RECT 139.295 19.975 139.525 20.045 ;
        RECT 139.045 19.795 139.335 19.815 ;
        RECT 135.885 19.255 138.350 19.620 ;
        RECT 139.020 19.545 139.355 19.795 ;
        RECT 1.475 18.380 112.080 19.255 ;
        RECT 113.475 18.380 140.080 19.255 ;
        RECT 27.790 17.960 30.690 17.980 ;
        RECT 55.390 17.960 57.890 17.980 ;
        RECT 68.845 17.960 69.785 17.985 ;
        RECT 83.690 17.960 86.190 17.980 ;
        RECT 1.450 17.280 111.925 17.960 ;
        RECT 1.450 17.260 27.925 17.280 ;
        RECT 29.450 17.260 55.925 17.280 ;
        RECT 57.450 17.260 83.925 17.280 ;
        RECT 85.450 17.260 111.925 17.280 ;
        RECT 113.450 17.260 139.925 17.960 ;
        RECT 2.420 16.635 4.330 17.260 ;
        RECT 6.420 16.925 8.305 16.930 ;
        RECT 9.865 16.925 11.750 16.930 ;
        RECT 6.410 16.695 8.370 16.925 ;
        RECT 9.840 16.695 11.800 16.925 ;
        RECT 2.385 16.405 4.385 16.635 ;
        RECT 6.130 16.410 6.360 16.490 ;
        RECT 1.950 13.060 2.180 16.355 ;
        RECT 4.590 16.275 4.820 16.355 ;
        RECT 4.560 13.060 4.820 16.275 ;
        RECT 1.950 11.245 4.820 13.060 ;
        RECT 1.950 8.825 2.180 11.245 ;
        RECT 1.590 8.395 2.180 8.825 ;
        RECT 3.075 8.640 3.335 8.960 ;
        RECT 4.560 8.645 4.820 11.245 ;
        RECT 5.890 8.990 6.360 16.410 ;
        RECT 6.850 9.775 7.740 16.695 ;
        RECT 8.420 16.390 8.650 16.490 ;
        RECT 8.420 16.380 8.775 16.390 ;
        RECT 9.560 16.380 9.790 16.490 ;
        RECT 3.130 8.480 3.280 8.640 ;
        RECT 1.590 3.255 2.085 8.395 ;
        RECT 3.105 8.345 3.310 8.480 ;
        RECT 4.590 8.395 4.820 8.645 ;
        RECT 5.610 8.550 6.360 8.990 ;
        RECT 6.780 8.775 7.795 9.775 ;
        RECT 2.385 8.115 4.385 8.345 ;
        RECT 5.610 6.355 5.980 8.550 ;
        RECT 6.130 8.490 6.360 8.550 ;
        RECT 6.850 8.285 7.740 8.775 ;
        RECT 8.420 8.580 9.790 16.380 ;
        RECT 10.325 11.635 11.215 16.695 ;
        RECT 11.850 16.410 12.080 16.490 ;
        RECT 10.320 10.015 11.220 11.635 ;
        RECT 10.325 9.605 11.215 10.015 ;
        RECT 10.250 8.605 11.280 9.605 ;
        RECT 11.850 8.625 12.225 16.410 ;
        RECT 12.500 16.025 14.180 17.260 ;
        RECT 15.015 16.025 19.940 16.035 ;
        RECT 12.500 15.545 19.940 16.025 ;
        RECT 12.500 13.285 14.180 15.545 ;
        RECT 15.015 15.125 19.940 15.545 ;
        RECT 14.520 14.935 14.775 14.960 ;
        RECT 14.520 14.920 14.795 14.935 ;
        RECT 14.490 14.645 14.825 14.920 ;
        RECT 15.000 14.895 20.000 15.125 ;
        RECT 20.210 14.935 20.465 14.960 ;
        RECT 14.520 14.630 14.775 14.645 ;
        RECT 15.000 14.455 20.000 14.685 ;
        RECT 20.205 14.645 20.465 14.935 ;
        RECT 20.210 14.630 20.465 14.645 ;
        RECT 15.045 14.445 19.900 14.455 ;
        RECT 15.045 12.920 17.690 12.925 ;
        RECT 13.720 12.720 17.690 12.920 ;
        RECT 13.720 12.690 17.680 12.720 ;
        RECT 12.560 12.335 12.895 12.610 ;
        RECT 13.440 12.440 13.670 12.485 ;
        RECT 8.420 8.560 8.775 8.580 ;
        RECT 8.420 8.490 8.650 8.560 ;
        RECT 9.560 8.490 9.790 8.580 ;
        RECT 10.320 8.465 11.230 8.605 ;
        RECT 11.850 8.490 12.240 8.625 ;
        RECT 10.310 8.285 11.320 8.465 ;
        RECT 6.410 8.055 8.370 8.285 ;
        RECT 9.840 8.055 11.800 8.285 ;
        RECT 7.130 7.085 7.460 8.055 ;
        RECT 9.865 8.050 11.750 8.055 ;
        RECT 12.045 6.355 12.240 8.490 ;
        RECT 12.630 6.830 12.820 12.335 ;
        RECT 13.250 11.105 13.670 12.440 ;
        RECT 14.975 11.105 16.320 12.690 ;
        RECT 13.250 9.720 16.320 11.105 ;
        RECT 13.250 8.990 13.670 9.720 ;
        RECT 13.245 8.485 13.670 8.990 ;
        RECT 12.630 6.640 12.945 6.830 ;
        RECT 2.950 6.125 6.910 6.355 ;
        RECT 8.380 6.125 12.340 6.355 ;
        RECT 12.755 6.130 12.945 6.640 ;
        RECT 2.670 5.515 2.900 5.965 ;
        RECT 4.150 5.515 4.940 6.125 ;
        RECT 2.670 5.210 4.940 5.515 ;
        RECT 2.615 5.195 4.940 5.210 ;
        RECT 2.530 4.350 4.940 5.195 ;
        RECT 2.530 3.975 2.900 4.350 ;
        RECT 2.670 3.965 2.900 3.975 ;
        RECT 4.150 3.805 4.940 4.350 ;
        RECT 6.960 5.880 7.190 5.965 ;
        RECT 8.100 5.880 8.330 5.965 ;
        RECT 6.960 4.055 8.330 5.880 ;
        RECT 6.960 3.965 7.190 4.055 ;
        RECT 2.950 3.575 6.910 3.805 ;
        RECT 2.530 3.255 2.755 3.265 ;
        RECT 7.430 3.255 7.920 4.055 ;
        RECT 8.100 3.965 8.330 4.055 ;
        RECT 9.815 5.745 11.155 6.125 ;
        RECT 12.390 5.745 12.620 5.965 ;
        RECT 9.815 4.150 12.620 5.745 ;
        RECT 9.815 3.805 11.155 4.150 ;
        RECT 12.390 3.965 12.620 4.150 ;
        RECT 8.380 3.575 12.340 3.805 ;
        RECT 12.770 3.785 12.945 6.130 ;
        RECT 13.245 5.965 13.540 8.485 ;
        RECT 14.975 8.280 16.320 9.720 ;
        RECT 17.730 12.390 17.960 12.485 ;
        RECT 18.205 12.390 18.695 14.445 ;
        RECT 19.265 12.920 19.900 12.925 ;
        RECT 19.150 12.690 23.110 12.920 ;
        RECT 18.870 12.390 19.100 12.485 ;
        RECT 17.730 8.565 19.100 12.390 ;
        RECT 17.730 8.485 17.960 8.565 ;
        RECT 18.870 8.485 19.100 8.565 ;
        RECT 20.525 8.280 21.870 12.690 ;
        RECT 23.160 12.420 23.390 12.485 ;
        RECT 24.045 12.425 24.520 17.260 ;
        RECT 25.845 16.455 26.525 17.260 ;
        RECT 26.945 16.735 27.280 16.985 ;
        RECT 26.960 16.710 27.250 16.735 ;
        RECT 30.420 16.635 32.330 17.260 ;
        RECT 34.420 16.925 36.305 16.930 ;
        RECT 37.865 16.925 39.750 16.930 ;
        RECT 34.410 16.695 36.370 16.925 ;
        RECT 37.840 16.695 39.800 16.925 ;
        RECT 26.770 16.455 27.000 16.505 ;
        RECT 25.845 15.955 27.000 16.455 ;
        RECT 24.915 12.735 25.250 12.985 ;
        RECT 24.935 12.705 25.225 12.735 ;
        RECT 24.745 12.425 24.975 12.500 ;
        RECT 23.160 8.485 23.615 12.420 ;
        RECT 24.045 11.680 24.975 12.425 ;
        RECT 24.380 8.565 24.975 11.680 ;
        RECT 24.745 8.500 24.975 8.565 ;
        RECT 25.185 12.475 25.415 12.500 ;
        RECT 25.185 8.920 25.695 12.475 ;
        RECT 25.185 8.550 25.880 8.920 ;
        RECT 26.380 8.600 27.000 15.955 ;
        RECT 25.185 8.500 25.415 8.550 ;
        RECT 13.720 8.250 17.680 8.280 ;
        RECT 19.150 8.250 23.110 8.280 ;
        RECT 13.720 8.090 23.110 8.250 ;
        RECT 13.720 8.050 17.680 8.090 ;
        RECT 19.150 8.050 23.110 8.090 ;
        RECT 23.275 6.660 23.615 8.485 ;
        RECT 24.925 6.660 25.345 8.305 ;
        RECT 23.275 6.505 25.345 6.660 ;
        RECT 23.350 6.390 25.345 6.505 ;
        RECT 13.810 6.125 17.770 6.355 ;
        RECT 19.240 6.125 23.200 6.355 ;
        RECT 13.245 5.205 13.760 5.965 ;
        RECT 13.315 4.025 13.760 5.205 ;
        RECT 13.530 3.965 13.760 4.025 ;
        RECT 15.190 3.805 16.145 6.125 ;
        RECT 17.820 5.900 18.050 5.965 ;
        RECT 18.960 5.900 19.190 5.965 ;
        RECT 17.820 4.030 19.190 5.900 ;
        RECT 17.820 3.965 18.050 4.030 ;
        RECT 12.755 3.255 12.945 3.785 ;
        RECT 13.810 3.575 17.770 3.805 ;
        RECT 18.225 3.255 18.780 4.030 ;
        RECT 18.960 3.965 19.190 4.030 ;
        RECT 20.635 3.805 21.590 6.125 ;
        RECT 23.350 5.970 23.615 6.390 ;
        RECT 24.925 6.115 25.345 6.390 ;
        RECT 25.580 7.355 25.880 8.550 ;
        RECT 26.770 8.505 27.000 8.600 ;
        RECT 27.210 16.430 27.440 16.505 ;
        RECT 27.210 9.110 27.985 16.430 ;
        RECT 30.385 16.405 32.385 16.635 ;
        RECT 34.130 16.410 34.360 16.490 ;
        RECT 29.950 13.060 30.180 16.355 ;
        RECT 32.590 16.275 32.820 16.355 ;
        RECT 32.560 13.060 32.820 16.275 ;
        RECT 29.950 11.245 32.820 13.060 ;
        RECT 27.210 8.580 28.060 9.110 ;
        RECT 29.950 8.825 30.180 11.245 ;
        RECT 27.210 8.505 27.440 8.580 ;
        RECT 26.875 7.825 27.390 8.315 ;
        RECT 27.690 7.825 28.060 8.580 ;
        RECT 29.590 8.395 30.180 8.825 ;
        RECT 31.075 8.640 31.335 8.960 ;
        RECT 32.560 8.645 32.820 11.245 ;
        RECT 33.890 8.990 34.360 16.410 ;
        RECT 34.850 9.775 35.740 16.695 ;
        RECT 36.420 16.390 36.650 16.490 ;
        RECT 36.420 16.380 36.775 16.390 ;
        RECT 37.560 16.380 37.790 16.490 ;
        RECT 31.130 8.480 31.280 8.640 ;
        RECT 26.875 7.360 27.385 7.825 ;
        RECT 26.510 7.355 27.385 7.360 ;
        RECT 25.580 6.950 27.385 7.355 ;
        RECT 25.580 6.110 25.880 6.950 ;
        RECT 26.510 6.935 27.385 6.950 ;
        RECT 26.875 6.825 27.385 6.935 ;
        RECT 26.875 6.125 27.390 6.825 ;
        RECT 27.615 6.795 28.615 7.825 ;
        RECT 23.275 5.965 23.615 5.970 ;
        RECT 23.250 4.020 23.615 5.965 ;
        RECT 24.830 5.900 25.060 5.970 ;
        RECT 24.335 5.230 25.060 5.900 ;
        RECT 24.325 5.040 25.060 5.230 ;
        RECT 24.325 4.240 24.680 5.040 ;
        RECT 24.830 4.970 25.060 5.040 ;
        RECT 25.270 5.925 25.500 5.970 ;
        RECT 25.640 5.925 25.880 6.110 ;
        RECT 25.270 5.595 25.880 5.925 ;
        RECT 26.855 5.870 27.085 5.975 ;
        RECT 25.270 5.040 25.765 5.595 ;
        RECT 25.270 4.970 25.500 5.040 ;
        RECT 25.020 4.785 25.310 4.810 ;
        RECT 25.005 4.535 25.340 4.785 ;
        RECT 26.625 4.765 27.085 5.870 ;
        RECT 26.305 4.240 27.085 4.765 ;
        RECT 23.885 4.060 27.085 4.240 ;
        RECT 23.250 3.965 23.480 4.020 ;
        RECT 19.240 3.575 23.200 3.805 ;
        RECT 23.885 3.620 26.690 4.060 ;
        RECT 26.855 3.975 27.085 4.060 ;
        RECT 27.295 5.910 27.525 5.975 ;
        RECT 27.690 5.910 28.060 6.795 ;
        RECT 27.295 5.585 28.060 5.910 ;
        RECT 27.295 4.045 28.055 5.585 ;
        RECT 27.295 3.975 27.525 4.045 ;
        RECT 27.045 3.795 27.335 3.815 ;
        RECT 23.885 3.255 26.350 3.620 ;
        RECT 27.020 3.545 27.355 3.795 ;
        RECT 29.590 3.280 30.085 8.395 ;
        RECT 31.105 8.345 31.310 8.480 ;
        RECT 32.590 8.395 32.820 8.645 ;
        RECT 33.610 8.550 34.360 8.990 ;
        RECT 34.780 8.775 35.795 9.775 ;
        RECT 30.385 8.115 32.385 8.345 ;
        RECT 33.610 6.355 33.980 8.550 ;
        RECT 34.130 8.490 34.360 8.550 ;
        RECT 34.850 8.285 35.740 8.775 ;
        RECT 36.420 8.580 37.790 16.380 ;
        RECT 38.325 11.635 39.215 16.695 ;
        RECT 39.850 16.410 40.080 16.490 ;
        RECT 38.320 10.015 39.220 11.635 ;
        RECT 38.325 9.605 39.215 10.015 ;
        RECT 38.250 8.605 39.280 9.605 ;
        RECT 39.850 8.625 40.225 16.410 ;
        RECT 40.500 16.025 42.180 17.260 ;
        RECT 43.015 16.025 47.940 16.035 ;
        RECT 40.500 15.545 47.940 16.025 ;
        RECT 40.500 13.285 42.180 15.545 ;
        RECT 43.015 15.125 47.940 15.545 ;
        RECT 42.520 14.935 42.775 14.960 ;
        RECT 42.520 14.920 42.795 14.935 ;
        RECT 42.490 14.645 42.825 14.920 ;
        RECT 43.000 14.895 48.000 15.125 ;
        RECT 48.210 14.935 48.465 14.960 ;
        RECT 42.520 14.630 42.775 14.645 ;
        RECT 43.000 14.455 48.000 14.685 ;
        RECT 48.205 14.645 48.465 14.935 ;
        RECT 48.210 14.630 48.465 14.645 ;
        RECT 43.045 14.445 47.900 14.455 ;
        RECT 43.045 12.920 45.690 12.925 ;
        RECT 41.720 12.720 45.690 12.920 ;
        RECT 41.720 12.690 45.680 12.720 ;
        RECT 40.560 12.335 40.895 12.610 ;
        RECT 41.440 12.440 41.670 12.485 ;
        RECT 36.420 8.560 36.775 8.580 ;
        RECT 36.420 8.490 36.650 8.560 ;
        RECT 37.560 8.490 37.790 8.580 ;
        RECT 38.320 8.465 39.230 8.605 ;
        RECT 39.850 8.490 40.240 8.625 ;
        RECT 38.310 8.285 39.320 8.465 ;
        RECT 34.410 8.055 36.370 8.285 ;
        RECT 37.840 8.055 39.800 8.285 ;
        RECT 35.210 7.040 35.560 8.055 ;
        RECT 37.865 8.050 39.750 8.055 ;
        RECT 40.045 6.355 40.240 8.490 ;
        RECT 40.630 6.830 40.820 12.335 ;
        RECT 41.250 11.105 41.670 12.440 ;
        RECT 42.975 11.105 44.320 12.690 ;
        RECT 41.250 9.720 44.320 11.105 ;
        RECT 41.250 8.990 41.670 9.720 ;
        RECT 41.245 8.485 41.670 8.990 ;
        RECT 40.630 6.640 40.945 6.830 ;
        RECT 30.950 6.125 34.910 6.355 ;
        RECT 36.380 6.125 40.340 6.355 ;
        RECT 40.755 6.130 40.945 6.640 ;
        RECT 30.670 5.515 30.900 5.965 ;
        RECT 32.150 5.515 32.940 6.125 ;
        RECT 30.670 5.210 32.940 5.515 ;
        RECT 30.615 5.195 32.940 5.210 ;
        RECT 30.530 4.350 32.940 5.195 ;
        RECT 30.530 3.975 30.900 4.350 ;
        RECT 30.670 3.965 30.900 3.975 ;
        RECT 32.150 3.805 32.940 4.350 ;
        RECT 34.960 5.880 35.190 5.965 ;
        RECT 36.100 5.880 36.330 5.965 ;
        RECT 34.960 4.055 36.330 5.880 ;
        RECT 34.960 3.965 35.190 4.055 ;
        RECT 30.950 3.575 34.910 3.805 ;
        RECT 27.990 3.255 30.090 3.280 ;
        RECT 30.530 3.255 30.755 3.265 ;
        RECT 35.430 3.255 35.920 4.055 ;
        RECT 36.100 3.965 36.330 4.055 ;
        RECT 37.815 5.745 39.155 6.125 ;
        RECT 40.390 5.745 40.620 5.965 ;
        RECT 37.815 4.150 40.620 5.745 ;
        RECT 37.815 3.805 39.155 4.150 ;
        RECT 40.390 3.965 40.620 4.150 ;
        RECT 36.380 3.575 40.340 3.805 ;
        RECT 40.770 3.785 40.945 6.130 ;
        RECT 41.245 5.965 41.540 8.485 ;
        RECT 42.975 8.280 44.320 9.720 ;
        RECT 45.730 12.390 45.960 12.485 ;
        RECT 46.205 12.390 46.695 14.445 ;
        RECT 47.265 12.920 47.900 12.925 ;
        RECT 47.150 12.690 51.110 12.920 ;
        RECT 46.870 12.390 47.100 12.485 ;
        RECT 45.730 8.565 47.100 12.390 ;
        RECT 45.730 8.485 45.960 8.565 ;
        RECT 46.870 8.485 47.100 8.565 ;
        RECT 48.525 8.280 49.870 12.690 ;
        RECT 51.160 12.420 51.390 12.485 ;
        RECT 52.045 12.425 52.520 17.260 ;
        RECT 53.845 16.455 54.525 17.260 ;
        RECT 54.945 16.735 55.280 16.985 ;
        RECT 54.960 16.710 55.250 16.735 ;
        RECT 58.420 16.635 60.330 17.260 ;
        RECT 62.420 16.925 64.305 16.930 ;
        RECT 65.865 16.925 67.750 16.930 ;
        RECT 62.410 16.695 64.370 16.925 ;
        RECT 65.840 16.695 67.800 16.925 ;
        RECT 54.770 16.455 55.000 16.505 ;
        RECT 53.845 15.955 55.000 16.455 ;
        RECT 52.915 12.735 53.250 12.985 ;
        RECT 52.935 12.705 53.225 12.735 ;
        RECT 52.745 12.425 52.975 12.500 ;
        RECT 51.160 8.485 51.615 12.420 ;
        RECT 52.045 11.680 52.975 12.425 ;
        RECT 52.380 8.565 52.975 11.680 ;
        RECT 52.745 8.500 52.975 8.565 ;
        RECT 53.185 12.475 53.415 12.500 ;
        RECT 53.185 8.920 53.695 12.475 ;
        RECT 53.185 8.550 53.880 8.920 ;
        RECT 54.380 8.600 55.000 15.955 ;
        RECT 53.185 8.500 53.415 8.550 ;
        RECT 41.720 8.250 45.680 8.280 ;
        RECT 47.150 8.250 51.110 8.280 ;
        RECT 41.720 8.090 51.110 8.250 ;
        RECT 41.720 8.050 45.680 8.090 ;
        RECT 47.150 8.050 51.110 8.090 ;
        RECT 51.275 6.660 51.615 8.485 ;
        RECT 52.925 6.660 53.345 8.305 ;
        RECT 51.275 6.505 53.345 6.660 ;
        RECT 51.350 6.390 53.345 6.505 ;
        RECT 41.810 6.125 45.770 6.355 ;
        RECT 47.240 6.125 51.200 6.355 ;
        RECT 41.245 5.205 41.760 5.965 ;
        RECT 41.315 4.025 41.760 5.205 ;
        RECT 41.530 3.965 41.760 4.025 ;
        RECT 43.190 3.805 44.145 6.125 ;
        RECT 45.820 5.900 46.050 5.965 ;
        RECT 46.960 5.900 47.190 5.965 ;
        RECT 45.820 4.030 47.190 5.900 ;
        RECT 45.820 3.965 46.050 4.030 ;
        RECT 40.755 3.255 40.945 3.785 ;
        RECT 41.810 3.575 45.770 3.805 ;
        RECT 46.225 3.255 46.780 4.030 ;
        RECT 46.960 3.965 47.190 4.030 ;
        RECT 48.635 3.805 49.590 6.125 ;
        RECT 51.350 5.970 51.615 6.390 ;
        RECT 52.925 6.115 53.345 6.390 ;
        RECT 53.580 7.355 53.880 8.550 ;
        RECT 54.770 8.505 55.000 8.600 ;
        RECT 55.210 16.430 55.440 16.505 ;
        RECT 55.210 9.110 55.985 16.430 ;
        RECT 58.385 16.405 60.385 16.635 ;
        RECT 62.130 16.410 62.360 16.490 ;
        RECT 57.950 13.060 58.180 16.355 ;
        RECT 60.590 16.275 60.820 16.355 ;
        RECT 60.560 13.060 60.820 16.275 ;
        RECT 57.950 11.245 60.820 13.060 ;
        RECT 55.210 8.580 56.060 9.110 ;
        RECT 57.950 8.825 58.180 11.245 ;
        RECT 55.210 8.505 55.440 8.580 ;
        RECT 54.875 7.825 55.390 8.315 ;
        RECT 54.875 7.360 55.385 7.825 ;
        RECT 55.690 7.795 56.060 8.580 ;
        RECT 57.590 8.395 58.180 8.825 ;
        RECT 59.075 8.640 59.335 8.960 ;
        RECT 60.560 8.645 60.820 11.245 ;
        RECT 61.890 8.990 62.360 16.410 ;
        RECT 62.850 9.775 63.740 16.695 ;
        RECT 64.420 16.390 64.650 16.490 ;
        RECT 64.420 16.380 64.775 16.390 ;
        RECT 65.560 16.380 65.790 16.490 ;
        RECT 59.130 8.480 59.280 8.640 ;
        RECT 54.510 7.355 55.385 7.360 ;
        RECT 53.580 6.950 55.385 7.355 ;
        RECT 53.580 6.110 53.880 6.950 ;
        RECT 54.510 6.935 55.385 6.950 ;
        RECT 54.875 6.825 55.385 6.935 ;
        RECT 54.875 6.125 55.390 6.825 ;
        RECT 55.615 6.795 56.645 7.795 ;
        RECT 51.275 5.965 51.615 5.970 ;
        RECT 51.250 4.020 51.615 5.965 ;
        RECT 52.830 5.900 53.060 5.970 ;
        RECT 52.335 5.230 53.060 5.900 ;
        RECT 52.325 5.040 53.060 5.230 ;
        RECT 52.325 4.240 52.680 5.040 ;
        RECT 52.830 4.970 53.060 5.040 ;
        RECT 53.270 5.925 53.500 5.970 ;
        RECT 53.640 5.925 53.880 6.110 ;
        RECT 53.270 5.595 53.880 5.925 ;
        RECT 54.855 5.870 55.085 5.975 ;
        RECT 53.270 5.040 53.765 5.595 ;
        RECT 53.270 4.970 53.500 5.040 ;
        RECT 53.020 4.785 53.310 4.810 ;
        RECT 53.005 4.535 53.340 4.785 ;
        RECT 54.625 4.765 55.085 5.870 ;
        RECT 54.305 4.240 55.085 4.765 ;
        RECT 51.885 4.060 55.085 4.240 ;
        RECT 51.250 3.965 51.480 4.020 ;
        RECT 47.240 3.575 51.200 3.805 ;
        RECT 51.885 3.620 54.690 4.060 ;
        RECT 54.855 3.975 55.085 4.060 ;
        RECT 55.295 5.910 55.525 5.975 ;
        RECT 55.690 5.910 56.060 6.795 ;
        RECT 55.295 5.585 56.060 5.910 ;
        RECT 55.295 4.045 56.055 5.585 ;
        RECT 55.295 3.975 55.525 4.045 ;
        RECT 55.045 3.795 55.335 3.815 ;
        RECT 51.885 3.255 54.350 3.620 ;
        RECT 55.020 3.545 55.355 3.795 ;
        RECT 57.590 3.280 58.085 8.395 ;
        RECT 59.105 8.345 59.310 8.480 ;
        RECT 60.590 8.395 60.820 8.645 ;
        RECT 61.610 8.550 62.360 8.990 ;
        RECT 62.780 8.775 63.795 9.775 ;
        RECT 58.385 8.115 60.385 8.345 ;
        RECT 61.610 6.355 61.980 8.550 ;
        RECT 62.130 8.490 62.360 8.550 ;
        RECT 62.850 8.285 63.740 8.775 ;
        RECT 64.420 8.580 65.790 16.380 ;
        RECT 66.325 11.635 67.215 16.695 ;
        RECT 67.850 16.410 68.080 16.490 ;
        RECT 66.320 10.015 67.220 11.635 ;
        RECT 66.325 9.605 67.215 10.015 ;
        RECT 66.250 8.605 67.280 9.605 ;
        RECT 67.850 8.625 68.225 16.410 ;
        RECT 68.500 16.025 70.180 17.260 ;
        RECT 71.015 16.025 75.940 16.035 ;
        RECT 68.500 15.545 75.940 16.025 ;
        RECT 68.500 13.285 70.180 15.545 ;
        RECT 71.015 15.125 75.940 15.545 ;
        RECT 70.520 14.935 70.775 14.960 ;
        RECT 70.520 14.920 70.795 14.935 ;
        RECT 70.490 14.645 70.825 14.920 ;
        RECT 71.000 14.895 76.000 15.125 ;
        RECT 76.210 14.935 76.465 14.960 ;
        RECT 70.520 14.630 70.775 14.645 ;
        RECT 71.000 14.455 76.000 14.685 ;
        RECT 76.205 14.645 76.465 14.935 ;
        RECT 76.210 14.630 76.465 14.645 ;
        RECT 71.045 14.445 75.900 14.455 ;
        RECT 71.045 12.920 73.690 12.925 ;
        RECT 69.720 12.720 73.690 12.920 ;
        RECT 69.720 12.690 73.680 12.720 ;
        RECT 68.560 12.335 68.895 12.610 ;
        RECT 69.440 12.440 69.670 12.485 ;
        RECT 64.420 8.560 64.775 8.580 ;
        RECT 64.420 8.490 64.650 8.560 ;
        RECT 65.560 8.490 65.790 8.580 ;
        RECT 66.320 8.465 67.230 8.605 ;
        RECT 67.850 8.490 68.240 8.625 ;
        RECT 66.310 8.285 67.320 8.465 ;
        RECT 62.410 8.055 64.370 8.285 ;
        RECT 65.840 8.055 67.800 8.285 ;
        RECT 63.125 7.090 63.470 8.055 ;
        RECT 65.865 8.050 67.750 8.055 ;
        RECT 68.045 6.355 68.240 8.490 ;
        RECT 68.630 6.830 68.820 12.335 ;
        RECT 69.250 11.105 69.670 12.440 ;
        RECT 70.975 11.105 72.320 12.690 ;
        RECT 69.250 9.720 72.320 11.105 ;
        RECT 69.250 8.990 69.670 9.720 ;
        RECT 69.245 8.485 69.670 8.990 ;
        RECT 68.630 6.640 68.945 6.830 ;
        RECT 58.950 6.125 62.910 6.355 ;
        RECT 64.380 6.125 68.340 6.355 ;
        RECT 68.755 6.130 68.945 6.640 ;
        RECT 58.670 5.515 58.900 5.965 ;
        RECT 60.150 5.515 60.940 6.125 ;
        RECT 58.670 5.210 60.940 5.515 ;
        RECT 58.615 5.195 60.940 5.210 ;
        RECT 58.530 4.350 60.940 5.195 ;
        RECT 58.530 3.975 58.900 4.350 ;
        RECT 58.670 3.965 58.900 3.975 ;
        RECT 60.150 3.805 60.940 4.350 ;
        RECT 62.960 5.880 63.190 5.965 ;
        RECT 64.100 5.880 64.330 5.965 ;
        RECT 62.960 4.055 64.330 5.880 ;
        RECT 62.960 3.965 63.190 4.055 ;
        RECT 58.950 3.575 62.910 3.805 ;
        RECT 55.790 3.255 58.085 3.280 ;
        RECT 58.530 3.255 58.755 3.265 ;
        RECT 63.430 3.255 63.920 4.055 ;
        RECT 64.100 3.965 64.330 4.055 ;
        RECT 65.815 5.745 67.155 6.125 ;
        RECT 68.390 5.745 68.620 5.965 ;
        RECT 65.815 4.150 68.620 5.745 ;
        RECT 65.815 3.805 67.155 4.150 ;
        RECT 68.390 3.965 68.620 4.150 ;
        RECT 64.380 3.575 68.340 3.805 ;
        RECT 68.770 3.785 68.945 6.130 ;
        RECT 69.245 5.965 69.540 8.485 ;
        RECT 70.975 8.280 72.320 9.720 ;
        RECT 73.730 12.390 73.960 12.485 ;
        RECT 74.205 12.390 74.695 14.445 ;
        RECT 75.265 12.920 75.900 12.925 ;
        RECT 75.150 12.690 79.110 12.920 ;
        RECT 74.870 12.390 75.100 12.485 ;
        RECT 73.730 8.565 75.100 12.390 ;
        RECT 73.730 8.485 73.960 8.565 ;
        RECT 74.870 8.485 75.100 8.565 ;
        RECT 76.525 8.280 77.870 12.690 ;
        RECT 79.160 12.420 79.390 12.485 ;
        RECT 80.045 12.425 80.520 17.260 ;
        RECT 81.845 16.455 82.525 17.260 ;
        RECT 82.945 16.735 83.280 16.985 ;
        RECT 82.960 16.710 83.250 16.735 ;
        RECT 86.420 16.635 88.330 17.260 ;
        RECT 90.420 16.925 92.305 16.930 ;
        RECT 93.865 16.925 95.750 16.930 ;
        RECT 90.410 16.695 92.370 16.925 ;
        RECT 93.840 16.695 95.800 16.925 ;
        RECT 82.770 16.455 83.000 16.505 ;
        RECT 81.845 15.955 83.000 16.455 ;
        RECT 80.915 12.735 81.250 12.985 ;
        RECT 80.935 12.705 81.225 12.735 ;
        RECT 80.745 12.425 80.975 12.500 ;
        RECT 79.160 8.485 79.615 12.420 ;
        RECT 80.045 11.680 80.975 12.425 ;
        RECT 80.380 8.565 80.975 11.680 ;
        RECT 80.745 8.500 80.975 8.565 ;
        RECT 81.185 12.475 81.415 12.500 ;
        RECT 81.185 8.920 81.695 12.475 ;
        RECT 81.185 8.550 81.880 8.920 ;
        RECT 82.380 8.600 83.000 15.955 ;
        RECT 81.185 8.500 81.415 8.550 ;
        RECT 69.720 8.250 73.680 8.280 ;
        RECT 75.150 8.250 79.110 8.280 ;
        RECT 69.720 8.090 79.110 8.250 ;
        RECT 69.720 8.050 73.680 8.090 ;
        RECT 75.150 8.050 79.110 8.090 ;
        RECT 79.275 6.660 79.615 8.485 ;
        RECT 80.925 6.660 81.345 8.305 ;
        RECT 79.275 6.505 81.345 6.660 ;
        RECT 79.350 6.390 81.345 6.505 ;
        RECT 69.810 6.125 73.770 6.355 ;
        RECT 75.240 6.125 79.200 6.355 ;
        RECT 69.245 5.205 69.760 5.965 ;
        RECT 69.315 4.025 69.760 5.205 ;
        RECT 69.530 3.965 69.760 4.025 ;
        RECT 71.190 3.805 72.145 6.125 ;
        RECT 73.820 5.900 74.050 5.965 ;
        RECT 74.960 5.900 75.190 5.965 ;
        RECT 73.820 4.030 75.190 5.900 ;
        RECT 73.820 3.965 74.050 4.030 ;
        RECT 68.755 3.255 68.945 3.785 ;
        RECT 69.810 3.575 73.770 3.805 ;
        RECT 74.225 3.255 74.780 4.030 ;
        RECT 74.960 3.965 75.190 4.030 ;
        RECT 76.635 3.805 77.590 6.125 ;
        RECT 79.350 5.970 79.615 6.390 ;
        RECT 80.925 6.115 81.345 6.390 ;
        RECT 81.580 7.355 81.880 8.550 ;
        RECT 82.770 8.505 83.000 8.600 ;
        RECT 83.210 16.430 83.440 16.505 ;
        RECT 83.210 9.110 83.985 16.430 ;
        RECT 86.385 16.405 88.385 16.635 ;
        RECT 90.130 16.410 90.360 16.490 ;
        RECT 85.950 13.060 86.180 16.355 ;
        RECT 88.590 16.275 88.820 16.355 ;
        RECT 88.560 13.060 88.820 16.275 ;
        RECT 85.950 11.245 88.820 13.060 ;
        RECT 83.210 8.580 84.060 9.110 ;
        RECT 85.950 8.825 86.180 11.245 ;
        RECT 83.210 8.505 83.440 8.580 ;
        RECT 82.875 7.825 83.390 8.315 ;
        RECT 82.875 7.360 83.385 7.825 ;
        RECT 83.690 7.795 84.060 8.580 ;
        RECT 85.590 8.395 86.180 8.825 ;
        RECT 87.075 8.640 87.335 8.960 ;
        RECT 88.560 8.645 88.820 11.245 ;
        RECT 89.890 8.990 90.360 16.410 ;
        RECT 90.850 9.775 91.740 16.695 ;
        RECT 92.420 16.390 92.650 16.490 ;
        RECT 92.420 16.380 92.775 16.390 ;
        RECT 93.560 16.380 93.790 16.490 ;
        RECT 87.130 8.480 87.280 8.640 ;
        RECT 82.510 7.355 83.385 7.360 ;
        RECT 81.580 6.950 83.385 7.355 ;
        RECT 81.580 6.110 81.880 6.950 ;
        RECT 82.510 6.935 83.385 6.950 ;
        RECT 82.875 6.825 83.385 6.935 ;
        RECT 82.875 6.125 83.390 6.825 ;
        RECT 83.615 6.795 84.645 7.795 ;
        RECT 79.275 5.965 79.615 5.970 ;
        RECT 79.250 4.020 79.615 5.965 ;
        RECT 80.830 5.900 81.060 5.970 ;
        RECT 80.335 5.230 81.060 5.900 ;
        RECT 80.325 5.040 81.060 5.230 ;
        RECT 80.325 4.240 80.680 5.040 ;
        RECT 80.830 4.970 81.060 5.040 ;
        RECT 81.270 5.925 81.500 5.970 ;
        RECT 81.640 5.925 81.880 6.110 ;
        RECT 81.270 5.595 81.880 5.925 ;
        RECT 82.855 5.870 83.085 5.975 ;
        RECT 81.270 5.040 81.765 5.595 ;
        RECT 81.270 4.970 81.500 5.040 ;
        RECT 81.020 4.785 81.310 4.810 ;
        RECT 81.005 4.535 81.340 4.785 ;
        RECT 82.625 4.765 83.085 5.870 ;
        RECT 82.305 4.240 83.085 4.765 ;
        RECT 79.885 4.060 83.085 4.240 ;
        RECT 79.250 3.965 79.480 4.020 ;
        RECT 75.240 3.575 79.200 3.805 ;
        RECT 79.885 3.620 82.690 4.060 ;
        RECT 82.855 3.975 83.085 4.060 ;
        RECT 83.295 5.910 83.525 5.975 ;
        RECT 83.690 5.910 84.060 6.795 ;
        RECT 83.295 5.585 84.060 5.910 ;
        RECT 83.295 4.045 84.055 5.585 ;
        RECT 83.295 3.975 83.525 4.045 ;
        RECT 83.045 3.795 83.335 3.815 ;
        RECT 79.885 3.255 82.350 3.620 ;
        RECT 83.020 3.545 83.355 3.795 ;
        RECT 85.590 3.280 86.085 8.395 ;
        RECT 87.105 8.345 87.310 8.480 ;
        RECT 88.590 8.395 88.820 8.645 ;
        RECT 89.610 8.550 90.360 8.990 ;
        RECT 90.780 8.775 91.795 9.775 ;
        RECT 86.385 8.115 88.385 8.345 ;
        RECT 89.610 6.355 89.980 8.550 ;
        RECT 90.130 8.490 90.360 8.550 ;
        RECT 90.850 8.285 91.740 8.775 ;
        RECT 92.420 8.580 93.790 16.380 ;
        RECT 94.325 11.635 95.215 16.695 ;
        RECT 95.850 16.410 96.080 16.490 ;
        RECT 94.320 10.015 95.220 11.635 ;
        RECT 94.325 9.605 95.215 10.015 ;
        RECT 94.250 8.605 95.280 9.605 ;
        RECT 95.850 8.625 96.225 16.410 ;
        RECT 96.500 16.025 98.180 17.260 ;
        RECT 99.015 16.025 103.940 16.035 ;
        RECT 96.500 15.545 103.940 16.025 ;
        RECT 96.500 13.285 98.180 15.545 ;
        RECT 99.015 15.125 103.940 15.545 ;
        RECT 98.520 14.935 98.775 14.960 ;
        RECT 98.520 14.920 98.795 14.935 ;
        RECT 98.490 14.645 98.825 14.920 ;
        RECT 99.000 14.895 104.000 15.125 ;
        RECT 104.210 14.935 104.465 14.960 ;
        RECT 98.520 14.630 98.775 14.645 ;
        RECT 99.000 14.455 104.000 14.685 ;
        RECT 104.205 14.645 104.465 14.935 ;
        RECT 104.210 14.630 104.465 14.645 ;
        RECT 99.045 14.445 103.900 14.455 ;
        RECT 99.045 12.920 101.690 12.925 ;
        RECT 97.720 12.720 101.690 12.920 ;
        RECT 97.720 12.690 101.680 12.720 ;
        RECT 96.560 12.335 96.895 12.610 ;
        RECT 97.440 12.440 97.670 12.485 ;
        RECT 92.420 8.560 92.775 8.580 ;
        RECT 92.420 8.490 92.650 8.560 ;
        RECT 93.560 8.490 93.790 8.580 ;
        RECT 94.320 8.465 95.230 8.605 ;
        RECT 95.850 8.490 96.240 8.625 ;
        RECT 94.310 8.285 95.320 8.465 ;
        RECT 90.410 8.055 92.370 8.285 ;
        RECT 93.840 8.055 95.800 8.285 ;
        RECT 91.095 6.975 91.495 8.055 ;
        RECT 93.865 8.050 95.750 8.055 ;
        RECT 96.045 6.355 96.240 8.490 ;
        RECT 96.630 6.830 96.820 12.335 ;
        RECT 97.250 11.105 97.670 12.440 ;
        RECT 98.975 11.105 100.320 12.690 ;
        RECT 97.250 9.720 100.320 11.105 ;
        RECT 97.250 8.990 97.670 9.720 ;
        RECT 97.245 8.485 97.670 8.990 ;
        RECT 96.630 6.640 96.945 6.830 ;
        RECT 86.950 6.125 90.910 6.355 ;
        RECT 92.380 6.125 96.340 6.355 ;
        RECT 96.755 6.130 96.945 6.640 ;
        RECT 86.670 5.515 86.900 5.965 ;
        RECT 88.150 5.515 88.940 6.125 ;
        RECT 86.670 5.210 88.940 5.515 ;
        RECT 86.615 5.195 88.940 5.210 ;
        RECT 86.530 4.350 88.940 5.195 ;
        RECT 86.530 3.975 86.900 4.350 ;
        RECT 86.670 3.965 86.900 3.975 ;
        RECT 88.150 3.805 88.940 4.350 ;
        RECT 90.960 5.880 91.190 5.965 ;
        RECT 92.100 5.880 92.330 5.965 ;
        RECT 90.960 4.055 92.330 5.880 ;
        RECT 90.960 3.965 91.190 4.055 ;
        RECT 86.950 3.575 90.910 3.805 ;
        RECT 83.890 3.255 86.085 3.280 ;
        RECT 86.530 3.255 86.755 3.265 ;
        RECT 91.430 3.255 91.920 4.055 ;
        RECT 92.100 3.965 92.330 4.055 ;
        RECT 93.815 5.745 95.155 6.125 ;
        RECT 96.390 5.745 96.620 5.965 ;
        RECT 93.815 4.150 96.620 5.745 ;
        RECT 93.815 3.805 95.155 4.150 ;
        RECT 96.390 3.965 96.620 4.150 ;
        RECT 92.380 3.575 96.340 3.805 ;
        RECT 96.770 3.785 96.945 6.130 ;
        RECT 97.245 5.965 97.540 8.485 ;
        RECT 98.975 8.280 100.320 9.720 ;
        RECT 101.730 12.390 101.960 12.485 ;
        RECT 102.205 12.390 102.695 14.445 ;
        RECT 103.265 12.920 103.900 12.925 ;
        RECT 103.150 12.690 107.110 12.920 ;
        RECT 102.870 12.390 103.100 12.485 ;
        RECT 101.730 8.565 103.100 12.390 ;
        RECT 101.730 8.485 101.960 8.565 ;
        RECT 102.870 8.485 103.100 8.565 ;
        RECT 104.525 8.280 105.870 12.690 ;
        RECT 107.160 12.420 107.390 12.485 ;
        RECT 108.045 12.425 108.520 17.260 ;
        RECT 109.845 16.455 110.525 17.260 ;
        RECT 110.945 16.735 111.280 16.985 ;
        RECT 110.960 16.710 111.250 16.735 ;
        RECT 114.420 16.635 116.330 17.260 ;
        RECT 118.420 16.925 120.305 16.930 ;
        RECT 121.865 16.925 123.750 16.930 ;
        RECT 118.410 16.695 120.370 16.925 ;
        RECT 121.840 16.695 123.800 16.925 ;
        RECT 110.770 16.455 111.000 16.505 ;
        RECT 109.845 15.955 111.000 16.455 ;
        RECT 108.915 12.735 109.250 12.985 ;
        RECT 108.935 12.705 109.225 12.735 ;
        RECT 108.745 12.425 108.975 12.500 ;
        RECT 107.160 8.485 107.615 12.420 ;
        RECT 108.045 11.680 108.975 12.425 ;
        RECT 108.380 8.565 108.975 11.680 ;
        RECT 108.745 8.500 108.975 8.565 ;
        RECT 109.185 12.475 109.415 12.500 ;
        RECT 109.185 8.920 109.695 12.475 ;
        RECT 109.185 8.550 109.880 8.920 ;
        RECT 110.380 8.600 111.000 15.955 ;
        RECT 109.185 8.500 109.415 8.550 ;
        RECT 97.720 8.250 101.680 8.280 ;
        RECT 103.150 8.250 107.110 8.280 ;
        RECT 97.720 8.090 107.110 8.250 ;
        RECT 97.720 8.050 101.680 8.090 ;
        RECT 103.150 8.050 107.110 8.090 ;
        RECT 107.275 6.660 107.615 8.485 ;
        RECT 108.925 6.660 109.345 8.305 ;
        RECT 107.275 6.505 109.345 6.660 ;
        RECT 107.350 6.390 109.345 6.505 ;
        RECT 97.810 6.125 101.770 6.355 ;
        RECT 103.240 6.125 107.200 6.355 ;
        RECT 97.245 5.205 97.760 5.965 ;
        RECT 97.315 4.025 97.760 5.205 ;
        RECT 97.530 3.965 97.760 4.025 ;
        RECT 99.190 3.805 100.145 6.125 ;
        RECT 101.820 5.900 102.050 5.965 ;
        RECT 102.960 5.900 103.190 5.965 ;
        RECT 101.820 4.030 103.190 5.900 ;
        RECT 101.820 3.965 102.050 4.030 ;
        RECT 96.755 3.255 96.945 3.785 ;
        RECT 97.810 3.575 101.770 3.805 ;
        RECT 102.225 3.255 102.780 4.030 ;
        RECT 102.960 3.965 103.190 4.030 ;
        RECT 104.635 3.805 105.590 6.125 ;
        RECT 107.350 5.970 107.615 6.390 ;
        RECT 108.925 6.115 109.345 6.390 ;
        RECT 109.580 7.355 109.880 8.550 ;
        RECT 110.770 8.505 111.000 8.600 ;
        RECT 111.210 16.430 111.440 16.505 ;
        RECT 111.210 9.110 111.985 16.430 ;
        RECT 114.385 16.405 116.385 16.635 ;
        RECT 118.130 16.410 118.360 16.490 ;
        RECT 113.950 13.060 114.180 16.355 ;
        RECT 116.590 16.275 116.820 16.355 ;
        RECT 116.560 13.060 116.820 16.275 ;
        RECT 113.950 11.245 116.820 13.060 ;
        RECT 111.210 8.580 112.060 9.110 ;
        RECT 113.950 8.825 114.180 11.245 ;
        RECT 111.210 8.505 111.440 8.580 ;
        RECT 110.875 7.825 111.390 8.315 ;
        RECT 110.875 7.360 111.385 7.825 ;
        RECT 111.690 7.795 112.060 8.580 ;
        RECT 113.590 8.395 114.180 8.825 ;
        RECT 115.075 8.640 115.335 8.960 ;
        RECT 116.560 8.645 116.820 11.245 ;
        RECT 117.890 8.990 118.360 16.410 ;
        RECT 118.850 9.775 119.740 16.695 ;
        RECT 120.420 16.390 120.650 16.490 ;
        RECT 120.420 16.380 120.775 16.390 ;
        RECT 121.560 16.380 121.790 16.490 ;
        RECT 115.130 8.480 115.280 8.640 ;
        RECT 110.510 7.355 111.385 7.360 ;
        RECT 109.580 6.950 111.385 7.355 ;
        RECT 109.580 6.110 109.880 6.950 ;
        RECT 110.510 6.935 111.385 6.950 ;
        RECT 110.875 6.825 111.385 6.935 ;
        RECT 110.875 6.125 111.390 6.825 ;
        RECT 111.615 6.795 112.645 7.795 ;
        RECT 107.275 5.965 107.615 5.970 ;
        RECT 107.250 4.020 107.615 5.965 ;
        RECT 108.830 5.900 109.060 5.970 ;
        RECT 108.335 5.230 109.060 5.900 ;
        RECT 108.325 5.040 109.060 5.230 ;
        RECT 108.325 4.240 108.680 5.040 ;
        RECT 108.830 4.970 109.060 5.040 ;
        RECT 109.270 5.925 109.500 5.970 ;
        RECT 109.640 5.925 109.880 6.110 ;
        RECT 109.270 5.595 109.880 5.925 ;
        RECT 110.855 5.870 111.085 5.975 ;
        RECT 109.270 5.040 109.765 5.595 ;
        RECT 109.270 4.970 109.500 5.040 ;
        RECT 109.020 4.785 109.310 4.810 ;
        RECT 109.005 4.535 109.340 4.785 ;
        RECT 110.625 4.765 111.085 5.870 ;
        RECT 110.305 4.240 111.085 4.765 ;
        RECT 107.885 4.060 111.085 4.240 ;
        RECT 107.250 3.965 107.480 4.020 ;
        RECT 103.240 3.575 107.200 3.805 ;
        RECT 107.885 3.620 110.690 4.060 ;
        RECT 110.855 3.975 111.085 4.060 ;
        RECT 111.295 5.910 111.525 5.975 ;
        RECT 111.690 5.910 112.060 6.795 ;
        RECT 111.295 5.585 112.060 5.910 ;
        RECT 111.295 4.045 112.055 5.585 ;
        RECT 111.295 3.975 111.525 4.045 ;
        RECT 111.045 3.795 111.335 3.815 ;
        RECT 107.885 3.255 110.350 3.620 ;
        RECT 111.020 3.545 111.355 3.795 ;
        RECT 113.590 3.280 114.085 8.395 ;
        RECT 115.105 8.345 115.310 8.480 ;
        RECT 116.590 8.395 116.820 8.645 ;
        RECT 117.610 8.550 118.360 8.990 ;
        RECT 118.780 8.775 119.795 9.775 ;
        RECT 114.385 8.115 116.385 8.345 ;
        RECT 117.610 6.355 117.980 8.550 ;
        RECT 118.130 8.490 118.360 8.550 ;
        RECT 118.850 8.285 119.740 8.775 ;
        RECT 120.420 8.580 121.790 16.380 ;
        RECT 122.325 11.635 123.215 16.695 ;
        RECT 123.850 16.410 124.080 16.490 ;
        RECT 122.320 10.015 123.220 11.635 ;
        RECT 122.325 9.605 123.215 10.015 ;
        RECT 122.250 8.605 123.280 9.605 ;
        RECT 123.850 8.625 124.225 16.410 ;
        RECT 124.500 16.025 126.180 17.260 ;
        RECT 127.015 16.025 131.940 16.035 ;
        RECT 124.500 15.545 131.940 16.025 ;
        RECT 124.500 13.285 126.180 15.545 ;
        RECT 127.015 15.125 131.940 15.545 ;
        RECT 126.520 14.935 126.775 14.960 ;
        RECT 126.520 14.920 126.795 14.935 ;
        RECT 126.490 14.645 126.825 14.920 ;
        RECT 127.000 14.895 132.000 15.125 ;
        RECT 132.210 14.935 132.465 14.960 ;
        RECT 126.520 14.630 126.775 14.645 ;
        RECT 127.000 14.455 132.000 14.685 ;
        RECT 132.205 14.645 132.465 14.935 ;
        RECT 132.210 14.630 132.465 14.645 ;
        RECT 127.045 14.445 131.900 14.455 ;
        RECT 127.045 12.920 129.690 12.925 ;
        RECT 125.720 12.720 129.690 12.920 ;
        RECT 125.720 12.690 129.680 12.720 ;
        RECT 124.560 12.335 124.895 12.610 ;
        RECT 125.440 12.440 125.670 12.485 ;
        RECT 120.420 8.560 120.775 8.580 ;
        RECT 120.420 8.490 120.650 8.560 ;
        RECT 121.560 8.490 121.790 8.580 ;
        RECT 122.320 8.465 123.230 8.605 ;
        RECT 123.850 8.490 124.240 8.625 ;
        RECT 122.310 8.285 123.320 8.465 ;
        RECT 118.410 8.055 120.370 8.285 ;
        RECT 121.840 8.055 123.800 8.285 ;
        RECT 119.150 7.155 119.435 8.055 ;
        RECT 121.865 8.050 123.750 8.055 ;
        RECT 124.045 6.355 124.240 8.490 ;
        RECT 124.630 6.830 124.820 12.335 ;
        RECT 125.250 11.105 125.670 12.440 ;
        RECT 126.975 11.105 128.320 12.690 ;
        RECT 125.250 9.720 128.320 11.105 ;
        RECT 125.250 8.990 125.670 9.720 ;
        RECT 125.245 8.485 125.670 8.990 ;
        RECT 124.630 6.640 124.945 6.830 ;
        RECT 114.950 6.125 118.910 6.355 ;
        RECT 120.380 6.125 124.340 6.355 ;
        RECT 124.755 6.130 124.945 6.640 ;
        RECT 114.670 5.515 114.900 5.965 ;
        RECT 116.150 5.515 116.940 6.125 ;
        RECT 114.670 5.210 116.940 5.515 ;
        RECT 114.615 5.195 116.940 5.210 ;
        RECT 114.530 4.350 116.940 5.195 ;
        RECT 114.530 3.975 114.900 4.350 ;
        RECT 114.670 3.965 114.900 3.975 ;
        RECT 116.150 3.805 116.940 4.350 ;
        RECT 118.960 5.880 119.190 5.965 ;
        RECT 120.100 5.880 120.330 5.965 ;
        RECT 118.960 4.055 120.330 5.880 ;
        RECT 118.960 3.965 119.190 4.055 ;
        RECT 114.950 3.575 118.910 3.805 ;
        RECT 111.590 3.255 114.085 3.280 ;
        RECT 114.530 3.255 114.755 3.265 ;
        RECT 119.430 3.255 119.920 4.055 ;
        RECT 120.100 3.965 120.330 4.055 ;
        RECT 121.815 5.745 123.155 6.125 ;
        RECT 124.390 5.745 124.620 5.965 ;
        RECT 121.815 4.150 124.620 5.745 ;
        RECT 121.815 3.805 123.155 4.150 ;
        RECT 124.390 3.965 124.620 4.150 ;
        RECT 120.380 3.575 124.340 3.805 ;
        RECT 124.770 3.785 124.945 6.130 ;
        RECT 125.245 5.965 125.540 8.485 ;
        RECT 126.975 8.280 128.320 9.720 ;
        RECT 129.730 12.390 129.960 12.485 ;
        RECT 130.205 12.390 130.695 14.445 ;
        RECT 131.265 12.920 131.900 12.925 ;
        RECT 131.150 12.690 135.110 12.920 ;
        RECT 130.870 12.390 131.100 12.485 ;
        RECT 129.730 8.565 131.100 12.390 ;
        RECT 129.730 8.485 129.960 8.565 ;
        RECT 130.870 8.485 131.100 8.565 ;
        RECT 132.525 8.280 133.870 12.690 ;
        RECT 135.160 12.420 135.390 12.485 ;
        RECT 136.045 12.425 136.520 17.260 ;
        RECT 137.845 16.455 138.525 17.260 ;
        RECT 138.945 16.735 139.280 16.985 ;
        RECT 138.960 16.710 139.250 16.735 ;
        RECT 138.770 16.455 139.000 16.505 ;
        RECT 137.845 15.955 139.000 16.455 ;
        RECT 136.915 12.735 137.250 12.985 ;
        RECT 136.935 12.705 137.225 12.735 ;
        RECT 136.745 12.425 136.975 12.500 ;
        RECT 135.160 8.485 135.615 12.420 ;
        RECT 136.045 11.680 136.975 12.425 ;
        RECT 136.380 8.565 136.975 11.680 ;
        RECT 136.745 8.500 136.975 8.565 ;
        RECT 137.185 12.475 137.415 12.500 ;
        RECT 137.185 8.920 137.695 12.475 ;
        RECT 137.185 8.550 137.880 8.920 ;
        RECT 138.380 8.600 139.000 15.955 ;
        RECT 137.185 8.500 137.415 8.550 ;
        RECT 125.720 8.250 129.680 8.280 ;
        RECT 131.150 8.250 135.110 8.280 ;
        RECT 125.720 8.090 135.110 8.250 ;
        RECT 125.720 8.050 129.680 8.090 ;
        RECT 131.150 8.050 135.110 8.090 ;
        RECT 135.275 6.660 135.615 8.485 ;
        RECT 136.925 6.660 137.345 8.305 ;
        RECT 135.275 6.505 137.345 6.660 ;
        RECT 135.350 6.390 137.345 6.505 ;
        RECT 125.810 6.125 129.770 6.355 ;
        RECT 131.240 6.125 135.200 6.355 ;
        RECT 125.245 5.205 125.760 5.965 ;
        RECT 125.315 4.025 125.760 5.205 ;
        RECT 125.530 3.965 125.760 4.025 ;
        RECT 127.190 3.805 128.145 6.125 ;
        RECT 129.820 5.900 130.050 5.965 ;
        RECT 130.960 5.900 131.190 5.965 ;
        RECT 129.820 4.030 131.190 5.900 ;
        RECT 129.820 3.965 130.050 4.030 ;
        RECT 124.755 3.255 124.945 3.785 ;
        RECT 125.810 3.575 129.770 3.805 ;
        RECT 130.225 3.255 130.780 4.030 ;
        RECT 130.960 3.965 131.190 4.030 ;
        RECT 132.635 3.805 133.590 6.125 ;
        RECT 135.350 5.970 135.615 6.390 ;
        RECT 136.925 6.115 137.345 6.390 ;
        RECT 137.580 7.355 137.880 8.550 ;
        RECT 138.770 8.505 139.000 8.600 ;
        RECT 139.210 16.430 139.440 16.505 ;
        RECT 139.210 9.110 139.985 16.430 ;
        RECT 139.210 8.580 140.060 9.110 ;
        RECT 139.210 8.505 139.440 8.580 ;
        RECT 138.875 7.825 139.390 8.315 ;
        RECT 138.875 7.360 139.385 7.825 ;
        RECT 139.690 7.795 140.060 8.580 ;
        RECT 138.510 7.355 139.385 7.360 ;
        RECT 137.580 6.950 139.385 7.355 ;
        RECT 137.580 6.110 137.880 6.950 ;
        RECT 138.510 6.935 139.385 6.950 ;
        RECT 138.875 6.825 139.385 6.935 ;
        RECT 138.875 6.125 139.390 6.825 ;
        RECT 139.615 6.795 140.645 7.795 ;
        RECT 135.275 5.965 135.615 5.970 ;
        RECT 135.250 4.020 135.615 5.965 ;
        RECT 136.830 5.900 137.060 5.970 ;
        RECT 136.335 5.230 137.060 5.900 ;
        RECT 136.325 5.040 137.060 5.230 ;
        RECT 136.325 4.240 136.680 5.040 ;
        RECT 136.830 4.970 137.060 5.040 ;
        RECT 137.270 5.925 137.500 5.970 ;
        RECT 137.640 5.925 137.880 6.110 ;
        RECT 137.270 5.595 137.880 5.925 ;
        RECT 138.855 5.870 139.085 5.975 ;
        RECT 137.270 5.040 137.765 5.595 ;
        RECT 137.270 4.970 137.500 5.040 ;
        RECT 137.020 4.785 137.310 4.810 ;
        RECT 137.005 4.535 137.340 4.785 ;
        RECT 138.625 4.765 139.085 5.870 ;
        RECT 138.305 4.240 139.085 4.765 ;
        RECT 135.885 4.060 139.085 4.240 ;
        RECT 135.250 3.965 135.480 4.020 ;
        RECT 131.240 3.575 135.200 3.805 ;
        RECT 135.885 3.620 138.690 4.060 ;
        RECT 138.855 3.975 139.085 4.060 ;
        RECT 139.295 5.910 139.525 5.975 ;
        RECT 139.690 5.910 140.060 6.795 ;
        RECT 139.295 5.585 140.060 5.910 ;
        RECT 139.295 4.045 140.055 5.585 ;
        RECT 139.295 3.975 139.525 4.045 ;
        RECT 139.045 3.795 139.335 3.815 ;
        RECT 135.885 3.255 138.350 3.620 ;
        RECT 139.020 3.545 139.355 3.795 ;
        RECT 1.475 2.380 140.080 3.255 ;
      LAYER met2 ;
        RECT 1.590 48.345 2.085 50.885 ;
        RECT 10.550 48.800 10.995 50.625 ;
        RECT 10.295 48.355 11.245 48.800 ;
        RECT 13.120 48.430 13.900 57.440 ;
        RECT 1.560 47.850 2.115 48.345 ;
        RECT 14.520 46.920 14.795 46.950 ;
        RECT 12.590 46.645 14.795 46.920 ;
        RECT 12.590 44.305 12.865 46.645 ;
        RECT 14.520 46.615 14.795 46.645 ;
        RECT 3.045 40.875 3.365 40.930 ;
        RECT 8.925 40.875 9.245 40.930 ;
        RECT 3.045 40.725 9.245 40.875 ;
        RECT 3.045 40.670 3.365 40.725 ;
        RECT 8.925 40.670 9.245 40.725 ;
        RECT 1.890 39.095 7.495 39.425 ;
        RECT 1.890 23.395 2.220 39.095 ;
        RECT 3.840 37.265 4.160 37.290 ;
        RECT 20.960 37.265 21.280 37.290 ;
        RECT 3.840 37.055 21.280 37.265 ;
        RECT 3.840 37.030 4.160 37.055 ;
        RECT 20.960 37.030 21.280 37.055 ;
        RECT 11.295 36.260 15.800 36.555 ;
        RECT 25.745 32.720 26.120 51.710 ;
        RECT 10.295 32.345 26.120 32.720 ;
        RECT 14.520 30.920 14.795 30.950 ;
        RECT 12.590 30.645 14.795 30.920 ;
        RECT 12.590 28.305 12.865 30.645 ;
        RECT 14.520 30.615 14.795 30.645 ;
        RECT 3.045 24.875 3.365 24.930 ;
        RECT 8.925 24.875 9.245 24.930 ;
        RECT 3.045 24.725 9.245 24.875 ;
        RECT 3.045 24.670 3.365 24.725 ;
        RECT 8.925 24.670 9.245 24.725 ;
        RECT 1.890 23.065 7.525 23.395 ;
        RECT 1.900 7.445 2.230 23.065 ;
        RECT 3.840 21.265 4.160 21.290 ;
        RECT 20.960 21.265 21.280 21.290 ;
        RECT 3.840 21.055 21.280 21.265 ;
        RECT 3.840 21.030 4.160 21.055 ;
        RECT 20.960 21.030 21.280 21.055 ;
        RECT 11.295 20.260 15.800 20.555 ;
        RECT 26.595 16.035 27.000 50.605 ;
        RECT 27.990 39.880 28.240 53.505 ;
        RECT 27.990 39.795 28.490 39.880 ;
        RECT 27.585 39.535 28.490 39.795 ;
        RECT 28.190 39.480 28.490 39.535 ;
        RECT 28.715 39.050 29.060 53.450 ;
        RECT 27.945 38.705 29.060 39.050 ;
        RECT 27.945 23.795 28.290 38.705 ;
        RECT 29.650 38.120 29.930 53.420 ;
        RECT 38.585 48.715 38.960 50.660 ;
        RECT 38.295 48.340 39.245 48.715 ;
        RECT 42.520 46.920 42.795 46.950 ;
        RECT 40.590 46.645 42.795 46.920 ;
        RECT 40.590 44.305 40.865 46.645 ;
        RECT 42.520 46.615 42.795 46.645 ;
        RECT 31.045 40.875 31.365 40.930 ;
        RECT 36.925 40.875 37.245 40.930 ;
        RECT 31.045 40.725 37.245 40.875 ;
        RECT 31.045 40.670 31.365 40.725 ;
        RECT 36.925 40.670 37.245 40.725 ;
        RECT 28.850 37.840 29.930 38.120 ;
        RECT 30.390 39.370 35.500 39.720 ;
        RECT 27.585 23.450 28.645 23.795 ;
        RECT 28.850 23.220 29.130 37.840 ;
        RECT 10.295 15.630 27.000 16.035 ;
        RECT 27.975 22.940 29.130 23.220 ;
        RECT 30.390 23.385 30.740 39.370 ;
        RECT 31.840 37.265 32.160 37.290 ;
        RECT 48.960 37.265 49.280 37.290 ;
        RECT 31.840 37.055 49.280 37.265 ;
        RECT 31.840 37.030 32.160 37.055 ;
        RECT 48.960 37.030 49.280 37.055 ;
        RECT 39.295 36.260 43.800 36.555 ;
        RECT 53.810 32.600 54.210 51.745 ;
        RECT 38.295 32.200 54.210 32.600 ;
        RECT 42.520 30.920 42.795 30.950 ;
        RECT 40.590 30.645 42.795 30.920 ;
        RECT 40.590 28.305 40.865 30.645 ;
        RECT 42.520 30.615 42.795 30.645 ;
        RECT 31.045 24.875 31.365 24.930 ;
        RECT 36.925 24.875 37.245 24.930 ;
        RECT 31.045 24.725 37.245 24.875 ;
        RECT 31.045 24.670 31.365 24.725 ;
        RECT 36.925 24.670 37.245 24.725 ;
        RECT 30.390 23.035 35.495 23.385 ;
        RECT 14.520 14.920 14.795 14.950 ;
        RECT 12.590 14.645 14.795 14.920 ;
        RECT 12.590 12.305 12.865 14.645 ;
        RECT 14.520 14.615 14.795 14.645 ;
        RECT 3.045 8.875 3.365 8.930 ;
        RECT 8.925 8.875 9.245 8.930 ;
        RECT 3.045 8.725 9.245 8.875 ;
        RECT 3.045 8.670 3.365 8.725 ;
        RECT 8.925 8.670 9.245 8.725 ;
        RECT 27.975 7.795 28.255 22.940 ;
        RECT 27.585 7.515 28.645 7.795 ;
        RECT 1.900 7.115 7.750 7.445 ;
        RECT 30.390 7.420 30.740 23.035 ;
        RECT 31.840 21.265 32.160 21.290 ;
        RECT 48.960 21.265 49.280 21.290 ;
        RECT 31.840 21.055 49.280 21.265 ;
        RECT 31.840 21.030 32.160 21.055 ;
        RECT 48.960 21.030 49.280 21.055 ;
        RECT 39.295 20.260 43.800 20.555 ;
        RECT 54.695 16.730 55.100 50.710 ;
        RECT 55.615 38.765 55.890 53.615 ;
        RECT 56.365 38.100 56.610 53.600 ;
        RECT 55.625 37.855 56.610 38.100 ;
        RECT 55.625 23.825 55.870 37.855 ;
        RECT 57.025 37.140 57.350 53.540 ;
        RECT 66.595 48.470 66.945 50.685 ;
        RECT 79.480 50.170 80.050 50.690 ;
        RECT 68.565 48.855 70.130 49.935 ;
        RECT 66.295 48.120 67.245 48.470 ;
        RECT 70.520 46.920 70.795 46.950 ;
        RECT 68.590 46.645 70.795 46.920 ;
        RECT 68.590 44.305 68.865 46.645 ;
        RECT 70.520 46.615 70.795 46.645 ;
        RECT 59.045 40.875 59.365 40.930 ;
        RECT 64.925 40.875 65.245 40.930 ;
        RECT 59.045 40.725 65.245 40.875 ;
        RECT 59.045 40.670 59.365 40.725 ;
        RECT 64.925 40.670 65.245 40.725 ;
        RECT 56.290 36.815 57.350 37.140 ;
        RECT 57.605 39.260 63.490 39.605 ;
        RECT 55.615 22.765 55.875 23.825 ;
        RECT 38.295 16.325 55.100 16.730 ;
        RECT 42.520 14.920 42.795 14.950 ;
        RECT 40.590 14.645 42.795 14.920 ;
        RECT 40.590 12.305 40.865 14.645 ;
        RECT 42.520 14.615 42.795 14.645 ;
        RECT 31.045 8.875 31.365 8.930 ;
        RECT 36.925 8.875 37.245 8.930 ;
        RECT 31.045 8.725 37.245 8.875 ;
        RECT 31.045 8.670 31.365 8.725 ;
        RECT 36.925 8.670 37.245 8.725 ;
        RECT 35.680 7.445 35.960 7.465 ;
        RECT 35.205 7.420 35.985 7.445 ;
        RECT 30.390 7.115 35.985 7.420 ;
        RECT 30.390 7.095 35.960 7.115 ;
        RECT 30.390 7.070 35.805 7.095 ;
        RECT 35.365 7.065 35.805 7.070 ;
        RECT 56.290 6.765 56.615 36.815 ;
        RECT 57.605 23.425 57.950 39.260 ;
        RECT 59.840 37.265 60.160 37.290 ;
        RECT 76.960 37.265 77.280 37.290 ;
        RECT 59.840 37.055 77.280 37.265 ;
        RECT 59.840 37.030 60.160 37.055 ;
        RECT 76.960 37.030 77.280 37.055 ;
        RECT 67.295 36.260 71.800 36.555 ;
        RECT 79.805 34.570 81.180 36.025 ;
        RECT 68.645 33.350 69.995 34.205 ;
        RECT 68.690 33.320 69.950 33.350 ;
        RECT 81.780 32.540 82.120 50.765 ;
        RECT 82.740 37.785 83.135 50.785 ;
        RECT 83.635 39.825 83.855 53.395 ;
        RECT 83.615 38.765 83.875 39.825 ;
        RECT 82.740 37.390 83.865 37.785 ;
        RECT 66.295 32.200 82.120 32.540 ;
        RECT 70.520 30.920 70.795 30.950 ;
        RECT 68.590 30.645 70.795 30.920 ;
        RECT 68.590 28.305 68.865 30.645 ;
        RECT 70.520 30.615 70.795 30.645 ;
        RECT 59.045 24.875 59.365 24.930 ;
        RECT 64.925 24.875 65.245 24.930 ;
        RECT 59.045 24.725 65.245 24.875 ;
        RECT 59.045 24.670 59.365 24.725 ;
        RECT 64.925 24.670 65.245 24.725 ;
        RECT 57.605 23.080 63.540 23.425 ;
        RECT 57.625 7.465 57.970 23.080 ;
        RECT 59.840 21.265 60.160 21.290 ;
        RECT 76.960 21.265 77.280 21.290 ;
        RECT 59.840 21.055 77.280 21.265 ;
        RECT 59.840 21.030 60.160 21.055 ;
        RECT 76.960 21.030 77.280 21.055 ;
        RECT 67.295 20.260 71.800 20.555 ;
        RECT 80.460 18.535 81.835 19.990 ;
        RECT 68.745 16.870 69.890 18.105 ;
        RECT 83.470 16.550 83.865 37.390 ;
        RECT 84.315 22.765 84.615 53.320 ;
        RECT 85.115 52.855 85.480 53.355 ;
        RECT 85.110 22.360 85.480 52.855 ;
        RECT 85.895 47.895 86.200 53.345 ;
        RECT 86.535 48.445 86.860 53.330 ;
        RECT 87.210 49.015 87.515 53.345 ;
        RECT 87.860 49.660 88.205 53.340 ;
        RECT 88.565 50.245 88.915 53.325 ;
        RECT 89.320 51.020 89.710 53.215 ;
        RECT 89.320 50.630 141.315 51.020 ;
        RECT 88.565 49.895 140.615 50.245 ;
        RECT 87.860 49.315 139.960 49.660 ;
        RECT 87.210 48.710 113.130 49.015 ;
        RECT 86.535 48.120 112.540 48.445 ;
        RECT 85.895 47.620 111.920 47.895 ;
        RECT 85.895 47.590 107.810 47.620 ;
        RECT 108.860 47.590 111.920 47.620 ;
        RECT 98.520 46.920 98.795 46.950 ;
        RECT 94.475 46.100 95.240 46.800 ;
        RECT 96.590 46.645 98.795 46.920 ;
        RECT 96.590 44.305 96.865 46.645 ;
        RECT 98.520 46.615 98.795 46.645 ;
        RECT 87.045 40.875 87.365 40.930 ;
        RECT 92.925 40.875 93.245 40.930 ;
        RECT 87.045 40.725 93.245 40.875 ;
        RECT 87.045 40.670 87.365 40.725 ;
        RECT 92.925 40.670 93.245 40.725 ;
        RECT 85.980 39.200 91.525 39.600 ;
        RECT 66.295 16.155 83.865 16.550 ;
        RECT 84.245 21.990 85.480 22.360 ;
        RECT 86.010 23.410 86.410 39.200 ;
        RECT 111.615 38.765 111.920 47.590 ;
        RECT 112.215 37.960 112.540 48.120 ;
        RECT 111.615 37.635 112.540 37.960 ;
        RECT 87.840 37.265 88.160 37.290 ;
        RECT 104.960 37.265 105.280 37.290 ;
        RECT 87.840 37.055 105.280 37.265 ;
        RECT 87.840 37.030 88.160 37.055 ;
        RECT 104.960 37.030 105.280 37.055 ;
        RECT 95.295 36.260 99.800 36.555 ;
        RECT 94.605 31.765 95.370 32.465 ;
        RECT 98.520 30.920 98.795 30.950 ;
        RECT 96.590 30.645 98.795 30.920 ;
        RECT 96.590 28.305 96.865 30.645 ;
        RECT 98.520 30.615 98.795 30.645 ;
        RECT 87.045 24.875 87.365 24.930 ;
        RECT 92.925 24.875 93.245 24.930 ;
        RECT 87.045 24.725 93.245 24.875 ;
        RECT 87.045 24.670 87.365 24.725 ;
        RECT 92.925 24.670 93.245 24.725 ;
        RECT 86.010 23.010 91.555 23.410 ;
        RECT 70.520 14.920 70.795 14.950 ;
        RECT 68.590 14.645 70.795 14.920 ;
        RECT 68.590 12.305 68.865 14.645 ;
        RECT 70.520 14.615 70.795 14.645 ;
        RECT 59.045 8.875 59.365 8.930 ;
        RECT 64.925 8.875 65.245 8.930 ;
        RECT 59.045 8.725 65.245 8.875 ;
        RECT 59.045 8.670 59.365 8.725 ;
        RECT 64.925 8.670 65.245 8.725 ;
        RECT 57.625 7.120 63.500 7.465 ;
        RECT 58.505 7.115 59.265 7.120 ;
        RECT 58.530 7.095 58.810 7.115 ;
        RECT 84.245 6.765 84.615 21.990 ;
        RECT 86.010 7.405 86.410 23.010 ;
        RECT 111.615 22.765 111.940 37.635 ;
        RECT 112.825 37.195 113.130 48.710 ;
        RECT 126.520 46.920 126.795 46.950 ;
        RECT 124.590 46.645 126.795 46.920 ;
        RECT 124.590 44.305 124.865 46.645 ;
        RECT 126.520 46.615 126.795 46.645 ;
        RECT 122.420 43.515 123.095 44.300 ;
        RECT 115.045 40.875 115.365 40.930 ;
        RECT 120.925 40.875 121.245 40.930 ;
        RECT 115.045 40.725 121.245 40.875 ;
        RECT 115.045 40.670 115.365 40.725 ;
        RECT 120.925 40.670 121.245 40.725 ;
        RECT 112.255 36.890 113.130 37.195 ;
        RECT 114.105 39.165 119.460 39.450 ;
        RECT 87.840 21.265 88.160 21.290 ;
        RECT 104.960 21.265 105.280 21.290 ;
        RECT 87.840 21.055 105.280 21.265 ;
        RECT 87.840 21.030 88.160 21.055 ;
        RECT 104.960 21.030 105.280 21.055 ;
        RECT 95.295 20.260 99.800 20.555 ;
        RECT 94.375 15.590 95.140 16.290 ;
        RECT 98.520 14.920 98.795 14.950 ;
        RECT 96.590 14.645 98.795 14.920 ;
        RECT 96.590 12.305 96.865 14.645 ;
        RECT 98.520 14.615 98.795 14.645 ;
        RECT 87.045 8.875 87.365 8.930 ;
        RECT 92.925 8.875 93.245 8.930 ;
        RECT 87.045 8.725 93.245 8.875 ;
        RECT 87.045 8.670 87.365 8.725 ;
        RECT 92.925 8.670 93.245 8.725 ;
        RECT 112.255 7.825 112.560 36.890 ;
        RECT 114.105 23.430 114.390 39.165 ;
        RECT 139.615 38.765 139.960 49.315 ;
        RECT 115.840 37.265 116.160 37.290 ;
        RECT 132.960 37.265 133.280 37.290 ;
        RECT 115.840 37.055 133.280 37.265 ;
        RECT 115.840 37.030 116.160 37.055 ;
        RECT 132.960 37.030 133.280 37.055 ;
        RECT 123.295 36.260 127.800 36.555 ;
        RECT 126.520 30.920 126.795 30.950 ;
        RECT 124.590 30.645 126.795 30.920 ;
        RECT 124.590 28.305 124.865 30.645 ;
        RECT 126.520 30.615 126.795 30.645 ;
        RECT 122.505 27.090 123.180 27.875 ;
        RECT 115.045 24.875 115.365 24.930 ;
        RECT 120.925 24.875 121.245 24.930 ;
        RECT 115.045 24.725 121.245 24.875 ;
        RECT 115.045 24.670 115.365 24.725 ;
        RECT 120.925 24.670 121.245 24.725 ;
        RECT 114.105 23.145 119.475 23.430 ;
        RECT 86.865 7.445 87.145 7.465 ;
        RECT 86.840 7.405 87.740 7.445 ;
        RECT 86.010 7.005 91.525 7.405 ;
        RECT 112.200 6.765 112.615 7.825 ;
        RECT 114.105 7.470 114.390 23.145 ;
        RECT 140.265 22.765 140.615 49.895 ;
        RECT 140.925 22.085 141.315 50.630 ;
        RECT 146.890 48.490 147.295 49.315 ;
        RECT 146.490 48.085 147.295 48.490 ;
        RECT 144.190 46.565 144.620 47.380 ;
        RECT 146.890 47.255 147.295 48.085 ;
        RECT 143.565 46.135 144.620 46.565 ;
        RECT 144.190 45.320 144.620 46.135 ;
        RECT 150.770 45.100 151.535 45.800 ;
        RECT 148.940 43.595 149.955 44.095 ;
        RECT 141.820 42.945 142.260 42.975 ;
        RECT 141.525 42.475 142.260 42.945 ;
        RECT 141.525 27.170 141.965 42.475 ;
        RECT 140.225 21.695 141.315 22.085 ;
        RECT 115.840 21.265 116.160 21.290 ;
        RECT 132.960 21.265 133.280 21.290 ;
        RECT 115.840 21.055 133.280 21.265 ;
        RECT 115.840 21.030 116.160 21.055 ;
        RECT 132.960 21.030 133.280 21.055 ;
        RECT 123.295 20.260 127.800 20.555 ;
        RECT 126.520 14.920 126.795 14.950 ;
        RECT 124.590 14.645 126.795 14.920 ;
        RECT 122.465 13.335 123.140 14.120 ;
        RECT 124.590 12.305 124.865 14.645 ;
        RECT 126.520 14.615 126.795 14.645 ;
        RECT 115.045 8.875 115.365 8.930 ;
        RECT 120.925 8.875 121.245 8.930 ;
        RECT 115.045 8.725 121.245 8.875 ;
        RECT 115.045 8.670 115.365 8.725 ;
        RECT 120.925 8.670 121.245 8.725 ;
        RECT 114.105 7.185 119.465 7.470 ;
        RECT 114.800 7.115 115.590 7.185 ;
        RECT 114.825 7.095 115.105 7.115 ;
        RECT 140.225 6.765 140.615 21.695 ;
        RECT 142.380 13.435 142.880 41.065 ;
        RECT 3.840 5.265 4.160 5.290 ;
        RECT 20.960 5.265 21.280 5.290 ;
        RECT 3.840 5.055 21.280 5.265 ;
        RECT 3.840 5.030 4.160 5.055 ;
        RECT 20.960 5.030 21.280 5.055 ;
        RECT 31.840 5.265 32.160 5.290 ;
        RECT 48.960 5.265 49.280 5.290 ;
        RECT 31.840 5.055 49.280 5.265 ;
        RECT 31.840 5.030 32.160 5.055 ;
        RECT 48.960 5.030 49.280 5.055 ;
        RECT 59.840 5.265 60.160 5.290 ;
        RECT 76.960 5.265 77.280 5.290 ;
        RECT 59.840 5.055 77.280 5.265 ;
        RECT 59.840 5.030 60.160 5.055 ;
        RECT 76.960 5.030 77.280 5.055 ;
        RECT 87.840 5.265 88.160 5.290 ;
        RECT 104.960 5.265 105.280 5.290 ;
        RECT 87.840 5.055 105.280 5.265 ;
        RECT 87.840 5.030 88.160 5.055 ;
        RECT 104.960 5.030 105.280 5.055 ;
        RECT 115.840 5.265 116.160 5.290 ;
        RECT 132.960 5.265 133.280 5.290 ;
        RECT 115.840 5.055 133.280 5.265 ;
        RECT 115.840 5.030 116.160 5.055 ;
        RECT 132.960 5.030 133.280 5.055 ;
        RECT 11.295 4.260 15.800 4.555 ;
        RECT 39.295 4.260 43.800 4.555 ;
        RECT 67.295 4.260 71.800 4.555 ;
        RECT 80.415 2.885 81.790 4.340 ;
        RECT 95.295 4.260 99.800 4.555 ;
        RECT 123.295 4.260 127.800 4.555 ;
      LAYER met3 ;
        RECT 79.480 50.170 80.050 50.690 ;
        RECT 68.665 49.870 69.975 49.875 ;
        RECT 68.635 48.950 70.005 49.870 ;
        RECT 68.665 48.945 69.975 48.950 ;
        RECT 146.510 48.490 146.965 48.515 ;
        RECT 94.645 48.085 146.965 48.490 ;
        RECT 94.645 46.215 95.050 48.085 ;
        RECT 146.510 48.060 146.965 48.085 ;
        RECT 143.585 46.565 144.065 46.590 ;
        RECT 95.565 46.470 107.495 46.565 ;
        RECT 109.175 46.470 144.065 46.565 ;
        RECT 95.565 46.135 144.065 46.470 ;
        RECT 79.805 34.570 81.180 36.025 ;
        RECT 68.665 34.225 69.975 34.230 ;
        RECT 68.635 33.330 70.005 34.225 ;
        RECT 68.665 33.325 69.975 33.330 ;
        RECT 95.565 32.295 95.995 46.135 ;
        RECT 143.585 46.110 144.065 46.135 ;
        RECT 150.825 45.680 151.375 45.705 ;
        RECT 94.695 31.865 95.995 32.295 ;
        RECT 96.770 45.180 151.375 45.680 ;
        RECT 80.460 18.535 81.835 19.990 ;
        RECT 68.660 16.800 69.980 18.180 ;
        RECT 96.770 16.190 97.270 45.180 ;
        RECT 150.825 45.155 151.375 45.180 ;
        RECT 148.960 44.095 149.510 44.120 ;
        RECT 122.495 43.595 149.510 44.095 ;
        RECT 148.960 43.570 149.510 43.595 ;
        RECT 141.500 27.655 141.990 27.680 ;
        RECT 122.590 27.215 141.990 27.655 ;
        RECT 141.500 27.190 141.990 27.215 ;
        RECT 94.530 15.690 97.270 16.190 ;
        RECT 142.355 13.980 142.905 14.005 ;
        RECT 122.560 13.480 142.905 13.980 ;
        RECT 142.355 13.455 142.905 13.480 ;
        RECT 7.350 7.445 7.730 7.470 ;
        RECT 7.350 7.115 142.905 7.445 ;
        RECT 7.350 7.090 7.730 7.115 ;
        RECT 80.415 2.885 81.790 4.340 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 80.525 50.625 81.705 50.740 ;
        RECT 79.535 50.230 81.705 50.625 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 68.660 18.155 69.980 49.875 ;
        RECT 80.525 35.855 81.705 50.230 ;
        RECT 79.870 34.675 81.705 35.855 ;
        RECT 68.655 16.825 69.985 18.155 ;
        RECT 80.525 4.270 81.705 34.675 ;
        RECT 80.495 3.030 81.735 4.270 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

