magic
tech sky130A
magscale 1 2
timestamp 1757914993
<< pwell >>
rect 7519 -21472 7606 -20305
<< locali >>
rect 3840 -19826 15792 -19798
rect 3840 -19914 3864 -19826
rect 15764 -19888 15792 -19826
rect 15764 -19912 15804 -19888
rect 3796 -19930 3864 -19914
rect 3796 -20020 3824 -19930
rect 4120 -19962 5476 -19934
rect 4120 -20020 4138 -19962
rect 3796 -20044 4138 -20020
rect 5454 -20014 5476 -19962
rect 5772 -19962 7106 -19934
rect 5772 -20014 5796 -19962
rect 5454 -20038 5796 -20014
rect 7082 -20016 7106 -19962
rect 7474 -19962 8816 -19934
rect 7474 -20016 7506 -19962
rect 8784 -19992 8816 -19962
rect 9112 -19962 10494 -19934
rect 9112 -19992 9164 -19962
rect 8784 -20002 9164 -19992
rect 8798 -20016 9140 -20002
rect 10472 -20010 10494 -19962
rect 10790 -19962 12156 -19934
rect 10790 -20010 10814 -19962
rect 7082 -20018 7142 -20016
rect 7438 -20018 7506 -20016
rect 7082 -20040 7506 -20018
rect 10472 -20024 10814 -20010
rect 12138 -20004 12156 -19962
rect 12452 -19962 13818 -19934
rect 12452 -20004 12480 -19962
rect 12138 -20024 12480 -20004
rect 13796 -19990 13818 -19962
rect 14114 -19962 15482 -19934
rect 14114 -19990 14138 -19962
rect 13796 -20020 14138 -19990
rect 15462 -20002 15482 -19962
rect 15778 -20002 15804 -19912
rect 15462 -20018 15804 -20002
rect 7082 -20056 7502 -20040
rect 2937 -22431 16660 -22403
rect 2937 -22551 2980 -22431
rect 16622 -22551 16660 -22431
rect 2937 -22578 16660 -22551
<< viali >>
rect 3864 -19912 15764 -19826
rect 3864 -19930 15778 -19912
rect 3824 -19934 15778 -19930
rect 3824 -20020 4120 -19934
rect 5476 -20014 5772 -19934
rect 7106 -20016 7474 -19934
rect 8816 -19992 9112 -19934
rect 10494 -20010 10790 -19934
rect 7142 -20018 7438 -20016
rect 12156 -20004 12452 -19934
rect 13818 -19990 14114 -19934
rect 15482 -20002 15778 -19934
rect 2980 -22551 16622 -22431
<< metal1 >>
rect 9188 -19769 9316 -19768
rect 3809 -19770 9316 -19769
rect 9914 -19769 10060 -19768
rect 9914 -19770 15830 -19769
rect 3809 -19826 15830 -19770
rect 3809 -19877 3864 -19826
rect 3748 -19930 3864 -19877
rect 15764 -19912 15830 -19826
rect 3748 -20020 3824 -19930
rect 4120 -20014 5476 -19934
rect 5772 -20014 7106 -19934
rect 4120 -20016 7106 -20014
rect 7474 -19992 8816 -19934
rect 9112 -19992 10494 -19934
rect 7474 -20010 10494 -19992
rect 10790 -20004 12156 -19934
rect 12452 -19990 13818 -19934
rect 14114 -19990 15482 -19934
rect 12452 -20002 15482 -19990
rect 15778 -20002 15830 -19912
rect 12452 -20004 15830 -20002
rect 10790 -20010 15830 -20004
rect 7474 -20016 15830 -20010
rect 4120 -20018 7142 -20016
rect 7438 -20017 15830 -20016
rect 7438 -20018 8878 -20017
rect 4120 -20020 8878 -20018
rect 3748 -20050 8878 -20020
rect 9076 -20050 15830 -20017
rect 3085 -20548 3541 -20157
rect 3748 -20203 3840 -20050
rect 3940 -20153 4003 -20095
rect 3748 -20337 3944 -20203
rect 4089 -20206 4487 -20203
rect 3073 -21753 3198 -20749
rect 3436 -21749 3561 -20745
rect 3830 -21378 3944 -20337
rect 4001 -20560 4487 -20206
rect 4789 -20520 5187 -20163
rect 5407 -20203 5499 -20050
rect 5600 -20148 5663 -20090
rect 5735 -20202 6133 -20186
rect 5407 -20369 5587 -20203
rect 4001 -20882 4172 -20560
rect 4001 -21373 4197 -20882
rect 4406 -21074 4804 -20717
rect 3942 -21486 4008 -21434
rect 3942 -21520 3994 -21486
rect 3875 -21720 4075 -21520
rect 3942 -21827 4008 -21720
rect 3053 -22403 3198 -21898
rect 3440 -22065 3556 -21900
rect 3812 -22031 3932 -21874
rect 4122 -21876 4197 -21373
rect 4396 -21733 4794 -21376
rect 5093 -21736 5199 -20747
rect 5473 -21378 5587 -20369
rect 5668 -20543 6133 -20202
rect 5668 -20859 5839 -20543
rect 6427 -20553 6825 -20196
rect 7074 -20207 7166 -20050
rect 7263 -20153 7326 -20095
rect 8749 -20179 8841 -20050
rect 8936 -20128 8999 -20070
rect 7327 -20201 7498 -20197
rect 7074 -20367 7258 -20207
rect 5668 -21369 5875 -20859
rect 6064 -21091 6462 -20734
rect 5598 -21521 5664 -21438
rect 5532 -21721 5732 -21521
rect 5598 -21831 5664 -21721
rect 3440 -22194 3559 -22065
rect 3440 -22319 3559 -22313
rect 3740 -22248 3932 -22031
rect 3999 -22240 4202 -21876
rect 5800 -21878 5875 -21369
rect 6064 -21725 6462 -21368
rect 6762 -21753 6887 -20749
rect 7144 -21382 7258 -20367
rect 7326 -20564 7786 -20201
rect 8060 -20548 8520 -20185
rect 8749 -20291 8927 -20179
rect 7327 -20884 7498 -20564
rect 7327 -21364 7513 -20884
rect 7705 -21076 8165 -20713
rect 7256 -21544 7308 -21434
rect 7204 -21744 7404 -21544
rect 7256 -21826 7308 -21744
rect 4373 -21919 4485 -21883
rect 4370 -21925 4488 -21919
rect 4898 -21920 5017 -21905
rect 4370 -22049 4488 -22043
rect 3440 -22403 3559 -22401
rect 3740 -22403 3832 -22248
rect 3937 -22351 4000 -22293
rect 4373 -22294 4485 -22049
rect 4771 -22112 5169 -21920
rect 5489 -22001 5609 -21880
rect 4771 -22231 4898 -22112
rect 5017 -22231 5169 -22112
rect 4771 -22277 5169 -22231
rect 5425 -22254 5609 -22001
rect 5655 -22216 5875 -21878
rect 7438 -21881 7513 -21364
rect 7705 -21737 8165 -21374
rect 8423 -21745 8548 -20741
rect 8813 -21354 8927 -20291
rect 8998 -20197 9169 -20187
rect 8998 -20560 9471 -20197
rect 9765 -20536 10225 -20173
rect 10434 -20197 10526 -20050
rect 10617 -20145 10680 -20087
rect 10434 -20295 10622 -20197
rect 10680 -20207 11140 -20185
rect 8998 -20874 9169 -20560
rect 8998 -21354 9194 -20874
rect 9394 -21096 9854 -20733
rect 8941 -21512 8991 -21424
rect 8884 -21712 9084 -21512
rect 8941 -21821 8991 -21712
rect 6039 -22130 6148 -21907
rect 6549 -21925 6667 -21919
rect 6417 -22043 6549 -21932
rect 6667 -22043 6815 -21932
rect 7134 -21999 7254 -21882
rect 6036 -22136 6154 -22130
rect 5655 -22242 5858 -22216
rect 5425 -22403 5517 -22254
rect 6036 -22260 6154 -22254
rect 5598 -22349 5661 -22291
rect 6039 -22305 6148 -22260
rect 6417 -22289 6815 -22043
rect 7064 -22256 7254 -21999
rect 7314 -22245 7517 -21881
rect 7693 -21958 7802 -21911
rect 7064 -22403 7156 -22256
rect 7258 -22356 7321 -22298
rect 7693 -22309 7802 -22069
rect 8060 -22136 8520 -21930
rect 8809 -21971 8929 -21874
rect 9119 -21876 9194 -21354
rect 9386 -21757 9846 -21394
rect 10108 -21760 10232 -20696
rect 10508 -21372 10622 -20295
rect 10674 -20548 11140 -20207
rect 11418 -20540 11878 -20177
rect 12125 -20187 12217 -20050
rect 12280 -20138 12343 -20080
rect 12125 -20351 12273 -20187
rect 12346 -20201 12517 -20200
rect 10674 -20887 10845 -20548
rect 10674 -21374 10890 -20887
rect 11063 -21088 11523 -20725
rect 10616 -21520 10666 -21427
rect 10573 -21720 10773 -21520
rect 10616 -21824 10666 -21720
rect 8745 -21981 8929 -21971
rect 8060 -22254 8220 -22136
rect 8338 -22254 8520 -22136
rect 8060 -22293 8520 -22254
rect 8715 -22248 8929 -21981
rect 8991 -22240 9194 -21876
rect 9389 -21922 9498 -21899
rect 9384 -22178 9502 -21922
rect 8715 -22395 8837 -22248
rect 8931 -22351 8994 -22293
rect 9753 -21958 10213 -21926
rect 9753 -22067 9955 -21958
rect 10064 -22067 10213 -21958
rect 10482 -21969 10592 -21878
rect 10815 -21886 10890 -21374
rect 11063 -21741 11523 -21378
rect 11773 -21745 11898 -20741
rect 12159 -21362 12273 -20351
rect 12337 -20564 12797 -20201
rect 13087 -20544 13547 -20181
rect 13773 -20195 13865 -20050
rect 13941 -20143 14004 -20085
rect 13773 -20341 13929 -20195
rect 14022 -20205 14482 -20201
rect 12346 -20882 12517 -20564
rect 12346 -21367 12556 -20882
rect 12740 -21096 13200 -20733
rect 12283 -21523 12333 -21429
rect 12227 -21723 12427 -21523
rect 12283 -21826 12333 -21723
rect 9753 -22289 10213 -22067
rect 10394 -22258 10592 -21969
rect 10664 -22244 10890 -21886
rect 11060 -21959 11169 -21881
rect 10664 -22250 10867 -22244
rect 9384 -22302 9502 -22296
rect 8546 -22403 8837 -22395
rect 10394 -22403 10486 -22258
rect 11060 -22285 11169 -22068
rect 11418 -22178 11878 -21922
rect 12163 -21967 12273 -21874
rect 12481 -21888 12556 -21367
rect 12724 -21745 13184 -21382
rect 13437 -21737 13562 -20733
rect 13815 -21370 13929 -20341
rect 14002 -20564 14482 -20205
rect 14752 -20544 15212 -20181
rect 15428 -20195 15520 -20050
rect 15604 -20140 15667 -20082
rect 15428 -20387 15592 -20195
rect 14002 -20862 14173 -20564
rect 14002 -21372 14200 -20862
rect 14397 -21096 14857 -20733
rect 13933 -21517 14002 -21419
rect 13888 -21717 14088 -21517
rect 13933 -21826 14002 -21717
rect 11418 -22285 11576 -22178
rect 10602 -22349 10665 -22291
rect 11694 -22285 11878 -22178
rect 12081 -22254 12273 -21967
rect 12336 -22239 12556 -21888
rect 12713 -22188 12822 -21897
rect 12336 -22252 12539 -22239
rect 11576 -22302 11694 -22296
rect 12081 -22403 12173 -22254
rect 13075 -21959 13535 -21922
rect 13075 -22068 13269 -21959
rect 13378 -22068 13535 -21959
rect 13825 -21975 13935 -21876
rect 14125 -21881 14200 -21372
rect 14397 -21745 14857 -21382
rect 15110 -21741 15235 -20737
rect 15478 -21370 15592 -20387
rect 15672 -20705 15809 -20188
rect 16054 -20544 16514 -20181
rect 15667 -21068 16127 -20705
rect 15672 -21221 15809 -21068
rect 15672 -21368 15817 -21221
rect 15638 -21437 15705 -21436
rect 15612 -21438 15705 -21437
rect 15596 -21525 15705 -21438
rect 15751 -21484 15817 -21368
rect 16001 -21398 16201 -21198
rect 15506 -21725 15706 -21525
rect 15765 -21684 15817 -21484
rect 15596 -21818 15705 -21725
rect 15760 -21743 15817 -21684
rect 16023 -21554 16166 -21398
rect 16023 -21663 16049 -21554
rect 16158 -21663 16166 -21554
rect 16023 -21735 16166 -21663
rect 16388 -21733 16513 -20729
rect 16049 -21742 16158 -21735
rect 15596 -21820 15691 -21818
rect 15612 -21823 15691 -21820
rect 13075 -22285 13535 -22068
rect 13739 -22256 13935 -21975
rect 13989 -22219 14200 -21881
rect 14374 -21948 14483 -21901
rect 13989 -22245 14192 -22219
rect 12286 -22356 12349 -22298
rect 12713 -22303 12822 -22297
rect 13739 -22403 13831 -22256
rect 13941 -22349 14004 -22291
rect 14374 -22305 14483 -22057
rect 14756 -22188 15216 -21910
rect 15494 -21957 15604 -21870
rect 15751 -21873 15817 -21743
rect 14756 -22273 14928 -22188
rect 15037 -22273 15216 -22188
rect 15410 -22250 15604 -21957
rect 15665 -22172 15817 -21873
rect 15665 -22249 15772 -22172
rect 14928 -22303 15037 -22297
rect 15410 -22403 15502 -22250
rect 16050 -22277 16510 -21914
rect 15597 -22351 15660 -22293
rect 2937 -22431 16660 -22403
rect 2937 -22499 2980 -22431
rect 2935 -22551 2980 -22499
rect 16622 -22499 16660 -22431
rect 16622 -22551 16661 -22499
rect 2935 -22615 16661 -22551
<< via1 >>
rect 3440 -22313 3559 -22194
rect 4370 -22043 4488 -21925
rect 4898 -22231 5017 -22112
rect 6549 -22043 6667 -21925
rect 6036 -22254 6154 -22136
rect 7693 -22069 7802 -21958
rect 8220 -22254 8338 -22136
rect 9384 -22296 9502 -22178
rect 9955 -22067 10064 -21958
rect 11060 -22068 11169 -21959
rect 11576 -22296 11694 -22178
rect 12713 -22297 12822 -22188
rect 13269 -22068 13378 -21959
rect 16049 -21663 16158 -21554
rect 14374 -22057 14483 -21948
rect 14928 -22297 15037 -22188
<< metal2 >>
rect 16049 -21554 16158 -21548
rect 4364 -22043 4370 -21925
rect 4488 -22043 6549 -21925
rect 6667 -22043 6673 -21925
rect 16049 -21948 16158 -21663
rect 7682 -21958 7812 -21954
rect 7682 -22069 7693 -21958
rect 7802 -22067 9955 -21958
rect 10064 -22067 10070 -21958
rect 7802 -22069 7812 -22067
rect 11054 -22068 11060 -21959
rect 11169 -22068 13269 -21959
rect 13378 -22068 13384 -21959
rect 14368 -22057 14374 -21948
rect 14483 -22057 16158 -21948
rect 7682 -22081 7812 -22069
rect 4898 -22112 5017 -22106
rect 3434 -22313 3440 -22194
rect 3559 -22231 4898 -22194
rect 3559 -22313 5017 -22231
rect 6030 -22254 6036 -22136
rect 6154 -22254 8220 -22136
rect 8338 -22254 8344 -22136
rect 9378 -22296 9384 -22178
rect 9502 -22296 11576 -22178
rect 11694 -22296 11700 -22178
rect 12707 -22297 12713 -22188
rect 12822 -22297 14928 -22188
rect 15037 -22297 15043 -22188
use sky130_fd_pr__nfet_01v8_ATLS57  XM1
timestamp 1757903622
transform 1 0 3966 0 1 -22062
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM2
timestamp 1757903622
transform 1 0 3970 0 1 -20794
box -211 -819 211 819
use sky130_fd_pr__nfet_01v8_ATLS57  XM3
timestamp 1757903622
transform 1 0 5627 0 1 -22062
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM4
timestamp 1757903622
transform 1 0 5629 0 1 -20791
box -211 -819 211 819
use sky130_fd_pr__nfet_01v8_ATLS57  XM5
timestamp 1757903622
transform 1 0 7279 0 1 -22062
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM6
timestamp 1757903622
transform 1 0 7292 0 1 -20793
box -211 -819 211 819
use sky130_fd_pr__nfet_01v8_ATLS57  XM7
timestamp 1757903622
transform 1 0 10633 0 1 -22062
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM8
timestamp 1757903622
transform 1 0 10646 0 1 -20788
box -211 -819 211 819
use sky130_fd_pr__nfet_01v8_ATLS57  XM9
timestamp 1757903622
transform 1 0 8963 0 1 -22058
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM10
timestamp 1757903622
transform 1 0 8968 0 1 -20773
box -211 -819 211 819
use sky130_fd_pr__nfet_01v8_ATLS57  XM11
timestamp 1757903622
transform 1 0 13958 0 1 -22061
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM12
timestamp 1757903622
transform 1 0 13971 0 1 -20780
box -211 -819 211 819
use sky130_fd_pr__nfet_01v8_ATLS57  XM13
timestamp 1757903622
transform 1 0 12310 0 1 -22063
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM14
timestamp 1757903622
transform 1 0 12312 0 1 -20783
box -211 -819 211 819
use sky130_fd_pr__nfet_01v8_ATLS57  XM15
timestamp 1757903622
transform 1 0 15631 0 1 -22061
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_XGA5KQ  XM16
timestamp 1757903622
transform 1 0 15631 0 1 -20784
box -211 -819 211 819
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR1
timestamp 1757903622
transform -1 0 6823 0 -1 -20625
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR2
timestamp 1757903622
transform -1 0 6459 0 -1 -20625
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR3
timestamp 1757903622
transform 1 0 3500 0 1 -20626
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR4
timestamp 1757903622
transform 1 0 3136 0 1 -21822
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR5
timestamp 1757903622
transform -1 0 6095 0 -1 -20625
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR6
timestamp 1757903622
transform 1 0 3500 0 1 -21822
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR7
timestamp 1757903622
transform -1 0 5157 0 -1 -20623
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR8
timestamp 1757903622
transform -1 0 6823 0 -1 -21821
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR9
timestamp 1757903622
transform -1 0 4793 0 -1 -20623
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR10
timestamp 1757903622
transform -1 0 4429 0 -1 -20623
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR11
timestamp 1757903622
transform -1 0 5157 0 -1 -21819
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR12
timestamp 1757903622
transform -1 0 4793 0 -1 -21819
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR13
timestamp 1757903622
transform -1 0 4429 0 -1 -21819
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR14
timestamp 1757903622
transform -1 0 6459 0 -1 -21821
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR15
timestamp 1757903622
transform -1 0 6095 0 -1 -21821
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR16
timestamp 1757903622
transform -1 0 8482 0 -1 -21823
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR17
timestamp 1757903622
transform -1 0 8118 0 -1 -21823
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR18
timestamp 1757903622
transform -1 0 7754 0 -1 -21823
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR19
timestamp 1757903622
transform -1 0 8482 0 -1 -20627
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR20
timestamp 1757903622
transform -1 0 8118 0 -1 -20627
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR21
timestamp 1757903622
transform -1 0 7754 0 -1 -20627
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR22
timestamp 1757903622
transform -1 0 11837 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR23
timestamp 1757903622
transform -1 0 11473 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR24
timestamp 1757903622
transform -1 0 11109 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR25
timestamp 1757903622
transform -1 0 11837 0 -1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR26
timestamp 1757903622
transform -1 0 11473 0 -1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR27
timestamp 1757903622
transform -1 0 11109 0 -1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR28
timestamp 1757903622
transform 1 0 13139 0 1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR29
timestamp 1757903622
transform 1 0 13503 0 1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR30
timestamp 1757903622
transform -1 0 12775 0 -1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR31
timestamp 1757903622
transform -1 0 13503 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR32
timestamp 1757903622
transform -1 0 13139 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR33
timestamp 1757903622
transform -1 0 12775 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR34
timestamp 1757903622
transform -1 0 10171 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR35
timestamp 1757903622
transform -1 0 9807 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR36
timestamp 1757903622
transform -1 0 9443 0 -1 -20624
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR37
timestamp 1757903622
transform -1 0 10171 0 -1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR38
timestamp 1757903622
transform -1 0 9807 0 -1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR39
timestamp 1757903622
transform -1 0 9443 0 -1 -21820
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR40
timestamp 1757903622
transform -1 0 15164 0 -1 -20625
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR41
timestamp 1757903622
transform -1 0 14800 0 -1 -20625
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR42
timestamp 1757903622
transform -1 0 14436 0 -1 -20625
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR43
timestamp 1757903622
transform -1 0 15164 0 -1 -21821
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR44
timestamp 1757903622
transform -1 0 14800 0 -1 -21821
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR45
timestamp 1757903622
transform -1 0 14436 0 -1 -21821
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR46
timestamp 1757903622
transform 1 0 16096 0 1 -21819
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR47
timestamp 1757903622
transform 1 0 16096 0 1 -20623
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR48
timestamp 1757903622
transform 1 0 16460 0 1 -21819
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR49
timestamp 1757903622
transform 1 0 16460 0 1 -20623
box -235 -651 235 651
use sky130_fd_pr__res_high_po_0p69_ZKG2N9  XR76
timestamp 1757903622
transform 1 0 3136 0 1 -20626
box -235 -651 235 651
<< labels >>
flabel metal1 7204 -21744 7404 -21544 0 FreeSans 256 0 0 0 B2
port 6 nsew
flabel metal1 5532 -21721 5732 -21521 0 FreeSans 256 0 0 0 B1
port 7 nsew
flabel metal1 10573 -21720 10773 -21520 0 FreeSans 256 0 0 0 B4
port 4 nsew
flabel metal1 3875 -21720 4075 -21520 0 FreeSans 256 0 0 0 B0
port 8 nsew
flabel metal1 12227 -21723 12427 -21523 0 FreeSans 256 0 0 0 B5
port 3 nsew
flabel metal1 8884 -21712 9084 -21512 0 FreeSans 256 0 0 0 B3
port 5 nsew
flabel metal1 13888 -21717 14088 -21517 0 FreeSans 256 0 0 0 B6
port 2 nsew
flabel metal1 15506 -21725 15706 -21525 0 FreeSans 256 0 0 0 B7
port 1 nsew
flabel metal1 8546 -22595 8746 -22395 0 FreeSans 256 0 0 0 VSS
port 10 nsew
flabel metal1 8512 -20026 8712 -19826 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 16001 -21398 16201 -21198 0 FreeSans 256 0 0 0 OUT
port 9 nsew
<< end >>
