VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adc_dac_tern_alu
  CLASS BLOCK ;
  FOREIGN tt_um_adc_dac_tern_alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 88.130 100.100 93.400 100.145 ;
        RECT 87.135 100.085 93.400 100.100 ;
        RECT 77.510 97.125 93.400 100.085 ;
        RECT 87.620 97.110 93.400 97.125 ;
      LAYER pwell ;
        RECT 79.770 93.945 87.730 96.965 ;
        RECT 77.790 93.855 87.750 93.945 ;
        RECT 71.780 90.895 87.750 93.855 ;
        RECT 77.790 90.845 87.750 90.895 ;
      LAYER nwell ;
        RECT 78.310 90.295 81.270 90.395 ;
        RECT 78.110 90.215 81.270 90.295 ;
        RECT 77.165 90.210 81.270 90.215 ;
        RECT 88.130 90.210 93.400 97.110 ;
        RECT 77.165 90.205 82.955 90.210 ;
        RECT 71.900 90.175 82.955 90.205 ;
        RECT 87.035 90.175 93.400 90.210 ;
        RECT 71.900 86.245 93.400 90.175 ;
        RECT 77.305 86.235 93.400 86.245 ;
        RECT 78.310 86.215 93.400 86.235 ;
        RECT 78.310 86.205 82.685 86.215 ;
        RECT 87.635 86.210 93.400 86.215 ;
        RECT 81.210 86.190 82.685 86.205 ;
      LAYER pwell ;
        RECT 71.880 77.915 87.830 85.875 ;
      LAYER nwell ;
        RECT 88.130 77.955 93.400 86.210 ;
      LAYER pwell ;
        RECT 93.550 77.965 95.660 100.065 ;
      LAYER nwell ;
        RECT 96.070 90.705 100.260 93.075 ;
        RECT 96.070 90.125 100.365 90.705 ;
        RECT 95.940 86.165 101.790 90.125 ;
      LAYER pwell ;
        RECT 96.090 77.975 101.760 85.935 ;
        RECT 79.780 61.570 83.950 74.060 ;
      LAYER nwell ;
        RECT 84.070 65.870 86.180 74.060 ;
      LAYER pwell ;
        RECT 84.050 61.575 86.160 65.675 ;
        RECT 86.245 61.585 92.235 74.075 ;
      LAYER nwell ;
        RECT 92.365 65.885 94.475 74.075 ;
      LAYER pwell ;
        RECT 92.355 61.575 94.465 65.675 ;
        RECT 94.575 61.575 100.565 74.065 ;
      LAYER nwell ;
        RECT 100.680 65.875 102.790 74.065 ;
      LAYER pwell ;
        RECT 100.615 61.575 102.725 65.675 ;
        RECT 102.870 61.565 108.860 74.055 ;
      LAYER nwell ;
        RECT 109.060 65.975 111.170 74.165 ;
      LAYER pwell ;
        RECT 109.035 61.595 111.145 65.695 ;
        RECT 111.315 61.580 117.305 74.070 ;
      LAYER nwell ;
        RECT 117.450 65.900 119.560 74.090 ;
      LAYER pwell ;
        RECT 117.385 61.575 119.495 65.675 ;
        RECT 119.645 61.580 125.635 74.070 ;
      LAYER nwell ;
        RECT 125.780 65.925 127.890 74.115 ;
      LAYER pwell ;
        RECT 125.770 61.570 127.880 65.670 ;
        RECT 127.975 61.580 133.965 74.070 ;
      LAYER nwell ;
        RECT 134.075 65.940 136.185 74.130 ;
      LAYER pwell ;
        RECT 134.010 61.580 136.120 65.680 ;
        RECT 136.280 61.575 142.270 74.065 ;
      LAYER nwell ;
        RECT 142.375 65.920 144.485 74.110 ;
      LAYER pwell ;
        RECT 142.375 61.580 144.485 65.680 ;
        RECT 144.580 61.585 148.750 74.075 ;
        RECT 1.710 52.730 14.200 58.190 ;
        RECT 1.710 50.380 32.140 52.730 ;
        RECT 43.730 50.380 62.200 52.730 ;
        RECT 67.730 50.380 86.200 52.730 ;
      LAYER nwell ;
        RECT 27.710 49.600 30.210 49.880 ;
        RECT 56.210 49.600 58.710 49.880 ;
        RECT 83.710 49.600 86.210 49.880 ;
        RECT 112.210 49.600 114.710 49.880 ;
        RECT 5.830 49.355 13.220 49.585 ;
        RECT 1.710 47.890 13.220 49.355 ;
        RECT 26.470 49.355 30.210 49.600 ;
        RECT 33.830 49.355 41.220 49.585 ;
        RECT 26.470 47.890 41.220 49.355 ;
        RECT 54.470 49.355 58.710 49.600 ;
        RECT 61.830 49.355 69.220 49.585 ;
        RECT 54.470 47.890 69.220 49.355 ;
        RECT 82.470 49.355 86.210 49.600 ;
        RECT 89.830 49.355 97.220 49.585 ;
        RECT 82.470 47.890 97.220 49.355 ;
        RECT 110.470 49.355 114.710 49.600 ;
        RECT 117.830 49.355 125.220 49.585 ;
        RECT 110.470 47.890 125.220 49.355 ;
        RECT 1.710 45.580 21.555 47.890 ;
        RECT 26.470 45.595 49.555 47.890 ;
        RECT 54.470 45.595 77.555 47.890 ;
        RECT 82.470 45.595 105.555 47.890 ;
        RECT 110.470 45.595 133.555 47.890 ;
        RECT 138.470 45.595 140.580 49.600 ;
        RECT 24.445 45.580 49.555 45.595 ;
        RECT 52.445 45.580 77.555 45.595 ;
        RECT 80.445 45.580 105.555 45.595 ;
        RECT 108.445 45.580 133.555 45.595 ;
        RECT 136.445 45.580 140.580 45.595 ;
        RECT 1.710 39.410 140.580 45.580 ;
      LAYER pwell ;
        RECT 143.710 44.730 150.220 50.190 ;
        RECT 143.710 40.560 156.200 44.730 ;
      LAYER nwell ;
        RECT 1.710 39.405 26.555 39.410 ;
        RECT 27.860 39.405 54.555 39.410 ;
        RECT 56.210 39.405 82.555 39.410 ;
        RECT 84.700 39.405 110.555 39.410 ;
        RECT 112.210 39.405 138.555 39.410 ;
        RECT 1.710 39.395 24.530 39.405 ;
        RECT 13.140 39.390 24.530 39.395 ;
        RECT 27.965 39.395 52.530 39.405 ;
        RECT 27.965 39.390 30.210 39.395 ;
        RECT 41.140 39.390 52.530 39.395 ;
        RECT 56.210 39.395 80.530 39.405 ;
        RECT 56.210 39.380 58.710 39.395 ;
        RECT 69.140 39.390 80.530 39.395 ;
        RECT 85.270 39.395 108.530 39.405 ;
        RECT 85.270 39.380 86.210 39.395 ;
        RECT 97.140 39.390 108.530 39.395 ;
        RECT 112.210 39.395 136.530 39.405 ;
        RECT 112.210 39.380 114.710 39.395 ;
        RECT 125.140 39.390 136.530 39.395 ;
      LAYER pwell ;
        RECT 26.555 39.020 28.665 39.025 ;
        RECT 54.555 39.020 56.665 39.025 ;
        RECT 82.555 39.020 84.665 39.025 ;
        RECT 110.555 39.020 112.665 39.025 ;
        RECT 138.555 39.020 140.665 39.025 ;
        RECT 24.530 39.015 28.665 39.020 ;
        RECT 52.530 39.015 56.665 39.020 ;
        RECT 80.530 39.015 84.665 39.020 ;
        RECT 108.530 39.015 112.665 39.020 ;
        RECT 136.530 39.015 140.665 39.020 ;
        RECT 2.370 35.920 28.665 39.015 ;
        RECT 2.370 34.915 24.620 35.920 ;
        RECT 26.555 34.925 28.665 35.920 ;
        RECT 30.370 35.920 56.665 39.015 ;
        RECT 30.370 34.915 52.620 35.920 ;
        RECT 54.555 34.925 56.665 35.920 ;
        RECT 58.370 35.920 84.665 39.015 ;
        RECT 58.370 34.915 80.620 35.920 ;
        RECT 82.555 34.925 84.665 35.920 ;
        RECT 86.370 35.920 112.665 39.015 ;
        RECT 86.370 34.915 108.620 35.920 ;
        RECT 110.555 34.925 112.665 35.920 ;
        RECT 114.370 35.920 140.665 39.015 ;
        RECT 114.370 34.915 136.620 35.920 ;
        RECT 138.555 34.925 140.665 35.920 ;
      LAYER nwell ;
        RECT 27.710 33.600 30.210 33.880 ;
        RECT 55.710 33.600 58.210 33.880 ;
        RECT 84.210 33.600 86.710 33.880 ;
        RECT 112.210 33.600 114.710 33.880 ;
        RECT 5.830 33.355 13.220 33.585 ;
        RECT 1.710 31.890 13.220 33.355 ;
        RECT 26.470 33.355 30.210 33.600 ;
        RECT 33.830 33.355 41.220 33.585 ;
        RECT 26.470 31.890 41.220 33.355 ;
        RECT 54.470 33.355 58.210 33.600 ;
        RECT 61.830 33.355 69.220 33.585 ;
        RECT 54.470 31.890 69.220 33.355 ;
        RECT 82.470 33.355 86.710 33.600 ;
        RECT 89.830 33.355 97.220 33.585 ;
        RECT 82.470 31.890 97.220 33.355 ;
        RECT 110.470 33.355 114.710 33.600 ;
        RECT 117.830 33.355 125.220 33.585 ;
        RECT 110.470 31.890 125.220 33.355 ;
        RECT 1.710 29.580 21.555 31.890 ;
        RECT 26.470 29.595 49.555 31.890 ;
        RECT 54.470 29.595 77.555 31.890 ;
        RECT 82.470 29.595 105.555 31.890 ;
        RECT 110.470 29.595 133.555 31.890 ;
        RECT 138.470 29.595 140.580 33.600 ;
        RECT 24.445 29.580 49.555 29.595 ;
        RECT 52.445 29.580 77.555 29.595 ;
        RECT 80.445 29.580 105.555 29.595 ;
        RECT 108.445 29.580 133.555 29.595 ;
        RECT 136.445 29.580 140.580 29.595 ;
        RECT 1.710 23.410 140.580 29.580 ;
        RECT 1.710 23.405 26.555 23.410 ;
        RECT 29.175 23.405 54.555 23.410 ;
        RECT 57.260 23.405 82.555 23.410 ;
        RECT 84.210 23.405 110.555 23.410 ;
        RECT 112.210 23.405 138.555 23.410 ;
        RECT 1.710 23.395 24.530 23.405 ;
        RECT 13.140 23.390 24.530 23.395 ;
        RECT 29.175 23.395 52.530 23.405 ;
        RECT 29.175 23.380 30.210 23.395 ;
        RECT 41.140 23.390 52.530 23.395 ;
        RECT 57.260 23.395 80.530 23.405 ;
        RECT 57.260 23.380 58.210 23.395 ;
        RECT 69.140 23.390 80.530 23.395 ;
        RECT 84.210 23.395 108.530 23.405 ;
        RECT 84.210 23.380 86.710 23.395 ;
        RECT 97.140 23.390 108.530 23.395 ;
        RECT 112.210 23.395 136.530 23.405 ;
        RECT 112.210 23.380 114.710 23.395 ;
        RECT 125.140 23.390 136.530 23.395 ;
      LAYER pwell ;
        RECT 26.555 23.020 28.665 23.025 ;
        RECT 54.555 23.020 56.665 23.025 ;
        RECT 82.555 23.020 84.665 23.025 ;
        RECT 110.555 23.020 112.665 23.025 ;
        RECT 138.555 23.020 140.665 23.025 ;
        RECT 24.530 23.015 28.665 23.020 ;
        RECT 52.530 23.015 56.665 23.020 ;
        RECT 80.530 23.015 84.665 23.020 ;
        RECT 108.530 23.015 112.665 23.020 ;
        RECT 136.530 23.015 140.665 23.020 ;
        RECT 2.370 19.920 28.665 23.015 ;
        RECT 2.370 18.915 24.620 19.920 ;
        RECT 26.555 18.925 28.665 19.920 ;
        RECT 30.370 19.920 56.665 23.015 ;
        RECT 30.370 18.915 52.620 19.920 ;
        RECT 54.555 18.925 56.665 19.920 ;
        RECT 58.370 19.920 84.665 23.015 ;
        RECT 58.370 18.915 80.620 19.920 ;
        RECT 82.555 18.925 84.665 19.920 ;
        RECT 86.370 19.920 112.665 23.015 ;
        RECT 86.370 18.915 108.620 19.920 ;
        RECT 110.555 18.925 112.665 19.920 ;
        RECT 114.370 19.920 140.665 23.015 ;
        RECT 114.370 18.915 136.620 19.920 ;
        RECT 138.555 18.925 140.665 19.920 ;
      LAYER nwell ;
        RECT 28.210 17.600 30.710 17.880 ;
        RECT 55.710 17.600 58.210 17.880 ;
        RECT 84.210 17.600 86.710 17.880 ;
        RECT 112.210 17.600 114.710 17.880 ;
        RECT 5.830 17.355 13.220 17.585 ;
        RECT 1.710 15.890 13.220 17.355 ;
        RECT 26.470 17.355 30.710 17.600 ;
        RECT 33.830 17.355 41.220 17.585 ;
        RECT 26.470 15.890 41.220 17.355 ;
        RECT 54.470 17.355 58.210 17.600 ;
        RECT 61.830 17.355 69.220 17.585 ;
        RECT 54.470 15.890 69.220 17.355 ;
        RECT 82.470 17.355 86.710 17.600 ;
        RECT 89.830 17.355 97.220 17.585 ;
        RECT 82.470 15.890 97.220 17.355 ;
        RECT 110.470 17.355 114.710 17.600 ;
        RECT 117.830 17.355 125.220 17.585 ;
        RECT 110.470 15.890 125.220 17.355 ;
        RECT 1.710 13.580 21.555 15.890 ;
        RECT 26.470 13.595 49.555 15.890 ;
        RECT 54.470 13.595 77.555 15.890 ;
        RECT 82.470 13.595 105.555 15.890 ;
        RECT 110.470 13.595 133.555 15.890 ;
        RECT 138.470 13.595 140.580 17.600 ;
        RECT 24.445 13.580 49.555 13.595 ;
        RECT 52.445 13.580 77.555 13.595 ;
        RECT 80.445 13.580 105.555 13.595 ;
        RECT 108.445 13.580 133.555 13.595 ;
        RECT 136.445 13.580 140.580 13.595 ;
        RECT 1.710 7.410 140.580 13.580 ;
        RECT 1.710 7.405 26.555 7.410 ;
        RECT 28.210 7.405 54.555 7.410 ;
        RECT 55.915 7.405 82.555 7.410 ;
        RECT 84.210 7.405 110.555 7.410 ;
        RECT 112.210 7.405 138.555 7.410 ;
        RECT 1.710 7.395 24.530 7.405 ;
        RECT 13.140 7.390 24.530 7.395 ;
        RECT 28.210 7.395 52.530 7.405 ;
        RECT 57.535 7.400 80.530 7.405 ;
        RECT 57.710 7.395 80.530 7.400 ;
        RECT 28.210 7.380 30.710 7.395 ;
        RECT 41.140 7.390 52.530 7.395 ;
        RECT 69.140 7.390 80.530 7.395 ;
        RECT 84.210 7.395 108.530 7.405 ;
        RECT 84.210 7.380 86.710 7.395 ;
        RECT 97.140 7.390 108.530 7.395 ;
        RECT 112.210 7.395 136.530 7.405 ;
        RECT 112.210 7.380 114.710 7.395 ;
        RECT 125.140 7.390 136.530 7.395 ;
      LAYER pwell ;
        RECT 26.555 7.020 28.665 7.025 ;
        RECT 54.555 7.020 56.665 7.025 ;
        RECT 82.555 7.020 84.665 7.025 ;
        RECT 110.555 7.020 112.665 7.025 ;
        RECT 138.555 7.020 140.665 7.025 ;
        RECT 24.530 7.015 28.665 7.020 ;
        RECT 52.530 7.015 56.665 7.020 ;
        RECT 80.530 7.015 84.665 7.020 ;
        RECT 108.530 7.015 112.665 7.020 ;
        RECT 136.530 7.015 140.665 7.020 ;
        RECT 2.370 3.920 28.665 7.015 ;
        RECT 2.370 2.915 24.620 3.920 ;
        RECT 26.555 2.925 28.665 3.920 ;
        RECT 30.370 3.920 56.665 7.015 ;
        RECT 30.370 2.915 52.620 3.920 ;
        RECT 54.555 2.925 56.665 3.920 ;
        RECT 58.370 3.920 84.665 7.015 ;
        RECT 58.370 2.915 80.620 3.920 ;
        RECT 82.555 2.925 84.665 3.920 ;
        RECT 86.370 3.920 112.665 7.015 ;
        RECT 86.370 2.915 108.620 3.920 ;
        RECT 110.555 2.925 112.665 3.920 ;
        RECT 114.370 3.920 140.665 7.015 ;
        RECT 114.370 2.915 136.620 3.920 ;
        RECT 138.555 2.925 140.665 3.920 ;
      LAYER li1 ;
        RECT 88.310 99.905 93.220 99.965 ;
        RECT 77.690 99.795 93.220 99.905 ;
        RECT 77.690 99.735 88.480 99.795 ;
        RECT 77.690 97.475 77.860 99.735 ;
        RECT 78.585 99.165 86.625 99.335 ;
        RECT 78.200 98.105 78.370 99.105 ;
        RECT 86.840 98.105 87.010 99.105 ;
        RECT 78.585 97.875 86.625 98.045 ;
        RECT 87.350 97.475 88.480 99.735 ;
        RECT 89.020 99.285 89.350 99.455 ;
        RECT 77.690 97.330 88.480 97.475 ;
        RECT 77.690 97.305 87.520 97.330 ;
        RECT 79.950 96.615 87.550 96.785 ;
        RECT 79.950 94.215 80.120 96.615 ;
        RECT 80.750 96.105 86.750 96.275 ;
        RECT 80.520 94.895 80.690 95.935 ;
        RECT 86.810 94.895 86.980 95.935 ;
        RECT 80.750 94.555 86.750 94.725 ;
        RECT 87.380 94.215 87.550 96.615 ;
        RECT 79.950 94.045 87.550 94.215 ;
        RECT 80.000 93.765 87.540 94.045 ;
        RECT 71.960 93.670 77.700 93.675 ;
        RECT 77.970 93.670 87.570 93.765 ;
        RECT 71.960 93.595 87.570 93.670 ;
        RECT 71.960 93.505 78.140 93.595 ;
        RECT 71.960 91.245 72.130 93.505 ;
        RECT 72.810 92.935 76.850 93.105 ;
        RECT 72.470 91.875 72.640 92.875 ;
        RECT 77.020 91.875 77.190 92.875 ;
        RECT 72.810 91.645 76.850 91.815 ;
        RECT 77.530 91.245 78.140 93.505 ;
        RECT 78.770 93.085 86.770 93.255 ;
        RECT 78.540 91.875 78.710 92.915 ;
        RECT 86.830 91.875 87.000 92.915 ;
        RECT 78.770 91.535 86.770 91.705 ;
        RECT 71.960 91.195 78.140 91.245 ;
        RECT 87.400 91.195 87.570 93.595 ;
        RECT 71.960 91.075 87.570 91.195 ;
        RECT 77.540 91.035 87.570 91.075 ;
        RECT 77.590 91.030 87.570 91.035 ;
        RECT 77.970 91.025 87.570 91.030 ;
        RECT 78.490 90.045 81.090 90.215 ;
        RECT 72.080 90.005 78.195 90.025 ;
        RECT 78.490 90.005 78.660 90.045 ;
        RECT 72.080 89.855 78.660 90.005 ;
        RECT 72.080 86.595 72.250 89.855 ;
        RECT 72.975 89.285 74.015 89.455 ;
        RECT 72.590 87.225 72.760 89.225 ;
        RECT 74.230 87.225 74.400 89.225 ;
        RECT 72.975 86.995 74.015 87.165 ;
        RECT 74.740 86.595 74.910 89.855 ;
        RECT 75.635 89.285 76.675 89.455 ;
        RECT 75.250 87.225 75.420 89.225 ;
        RECT 76.890 87.225 77.060 89.225 ;
        RECT 75.635 86.995 76.675 87.165 ;
        RECT 77.400 86.595 78.660 89.855 ;
        RECT 80.920 89.990 81.090 90.045 ;
        RECT 82.160 89.990 87.650 89.995 ;
        RECT 80.920 89.825 87.650 89.990 ;
        RECT 79.290 89.535 80.290 89.705 ;
        RECT 79.060 87.280 79.230 89.320 ;
        RECT 80.350 87.280 80.520 89.320 ;
        RECT 79.290 86.895 80.290 87.065 ;
        RECT 72.080 86.555 78.660 86.595 ;
        RECT 80.920 86.565 82.365 89.825 ;
        RECT 83.055 89.255 84.095 89.425 ;
        RECT 82.670 87.195 82.840 89.195 ;
        RECT 84.310 87.195 84.480 89.195 ;
        RECT 83.055 86.965 84.095 87.135 ;
        RECT 84.820 86.565 84.990 89.825 ;
        RECT 85.715 89.255 86.755 89.425 ;
        RECT 85.330 87.195 85.500 89.195 ;
        RECT 86.970 87.195 87.140 89.195 ;
        RECT 85.715 86.965 86.755 87.135 ;
        RECT 87.480 86.565 87.650 89.825 ;
        RECT 80.920 86.555 87.650 86.565 ;
        RECT 72.080 86.455 87.650 86.555 ;
        RECT 72.080 86.425 77.570 86.455 ;
        RECT 78.490 86.405 87.650 86.455 ;
        RECT 78.490 86.385 81.090 86.405 ;
        RECT 82.160 86.395 87.650 86.405 ;
        RECT 72.060 85.525 87.650 85.695 ;
        RECT 72.060 78.275 72.230 85.525 ;
        RECT 72.910 84.955 73.950 85.125 ;
        RECT 72.570 78.895 72.740 84.895 ;
        RECT 74.120 78.895 74.290 84.895 ;
        RECT 72.910 78.665 73.950 78.835 ;
        RECT 74.630 78.275 74.800 85.525 ;
        RECT 75.480 84.955 76.520 85.125 ;
        RECT 75.140 78.895 75.310 84.895 ;
        RECT 76.690 78.895 76.860 84.895 ;
        RECT 75.480 78.665 76.520 78.835 ;
        RECT 77.200 78.275 77.370 85.525 ;
        RECT 78.050 84.955 79.090 85.125 ;
        RECT 77.710 78.895 77.880 84.895 ;
        RECT 79.260 78.895 79.430 84.895 ;
        RECT 78.050 78.665 79.090 78.835 ;
        RECT 79.770 78.275 79.940 85.525 ;
        RECT 80.620 84.955 81.660 85.125 ;
        RECT 80.280 78.895 80.450 84.895 ;
        RECT 81.830 78.895 82.000 84.895 ;
        RECT 80.620 78.665 81.660 78.835 ;
        RECT 82.340 78.275 82.510 85.525 ;
        RECT 83.190 84.955 84.230 85.125 ;
        RECT 82.850 78.895 83.020 84.895 ;
        RECT 84.400 78.895 84.570 84.895 ;
        RECT 83.190 78.665 84.230 78.835 ;
        RECT 84.910 78.275 85.080 85.525 ;
        RECT 85.760 84.955 86.800 85.125 ;
        RECT 85.420 78.895 85.590 84.895 ;
        RECT 86.970 78.895 87.140 84.895 ;
        RECT 85.760 78.665 86.800 78.835 ;
        RECT 87.480 78.275 87.650 85.525 ;
        RECT 88.310 78.305 88.480 97.330 ;
        RECT 88.880 79.030 89.050 99.070 ;
        RECT 89.320 79.030 89.490 99.070 ;
        RECT 89.020 78.645 89.350 78.815 ;
        RECT 89.890 78.305 90.060 99.795 ;
        RECT 90.600 99.285 90.930 99.455 ;
        RECT 90.460 79.030 90.630 99.070 ;
        RECT 90.900 79.030 91.070 99.070 ;
        RECT 90.600 78.645 90.930 78.815 ;
        RECT 91.470 78.305 91.640 99.795 ;
        RECT 92.180 99.285 92.510 99.455 ;
        RECT 92.040 79.030 92.210 99.070 ;
        RECT 92.480 79.030 92.650 99.070 ;
        RECT 92.180 78.645 92.510 78.815 ;
        RECT 93.050 78.305 93.220 99.795 ;
        RECT 72.055 77.830 87.655 78.275 ;
        RECT 88.310 78.135 93.220 78.305 ;
        RECT 93.730 99.715 95.480 99.885 ;
        RECT 93.730 78.315 93.900 99.715 ;
        RECT 94.440 99.205 94.770 99.375 ;
        RECT 94.300 78.995 94.470 99.035 ;
        RECT 94.740 78.995 94.910 99.035 ;
        RECT 95.310 85.765 95.480 99.715 ;
        RECT 96.300 92.895 99.080 93.380 ;
        RECT 96.250 92.725 100.080 92.895 ;
        RECT 96.250 90.485 96.420 92.725 ;
        RECT 97.145 92.155 99.185 92.325 ;
        RECT 96.760 91.095 96.930 92.095 ;
        RECT 99.400 91.095 99.570 92.095 ;
        RECT 97.145 90.865 99.185 91.035 ;
        RECT 99.910 90.485 100.080 92.725 ;
        RECT 96.250 90.295 100.125 90.485 ;
        RECT 96.255 89.945 100.125 90.295 ;
        RECT 96.120 89.775 101.610 89.945 ;
        RECT 96.120 86.515 96.290 89.775 ;
        RECT 97.015 89.205 98.055 89.375 ;
        RECT 96.630 87.145 96.800 89.145 ;
        RECT 98.270 87.145 98.440 89.145 ;
        RECT 97.015 86.915 98.055 87.085 ;
        RECT 98.780 86.515 98.950 89.775 ;
        RECT 99.675 89.205 100.715 89.375 ;
        RECT 99.290 87.145 99.460 89.145 ;
        RECT 100.930 87.145 101.100 89.145 ;
        RECT 99.675 86.915 100.715 87.085 ;
        RECT 101.440 86.515 101.610 89.775 ;
        RECT 96.120 86.345 101.610 86.515 ;
        RECT 95.310 85.755 96.435 85.765 ;
        RECT 95.310 85.585 101.580 85.755 ;
        RECT 94.440 78.655 94.770 78.825 ;
        RECT 95.310 78.325 96.440 85.585 ;
        RECT 97.120 85.015 98.160 85.185 ;
        RECT 96.780 78.955 96.950 84.955 ;
        RECT 98.330 78.955 98.500 84.955 ;
        RECT 97.120 78.725 98.160 78.895 ;
        RECT 98.840 78.325 99.010 85.585 ;
        RECT 99.690 85.015 100.730 85.185 ;
        RECT 99.350 78.955 99.520 84.955 ;
        RECT 100.900 78.955 101.070 84.955 ;
        RECT 99.690 78.725 100.730 78.895 ;
        RECT 101.410 78.325 101.580 85.585 ;
        RECT 95.310 78.315 101.580 78.325 ;
        RECT 93.730 78.195 101.580 78.315 ;
        RECT 93.670 78.155 101.580 78.195 ;
        RECT 93.670 77.830 101.555 78.155 ;
        RECT 72.055 76.990 101.555 77.830 ;
        RECT 72.055 76.920 94.120 76.990 ;
        RECT 72.055 76.870 87.655 76.920 ;
        RECT 84.475 74.495 144.235 74.945 ;
        RECT 84.475 74.365 144.295 74.495 ;
        RECT 84.255 74.125 144.295 74.365 ;
        RECT 84.255 73.880 85.965 74.125 ;
        RECT 92.545 73.895 94.255 74.125 ;
        RECT 79.960 73.710 83.770 73.880 ;
        RECT 79.960 67.900 80.130 73.710 ;
        RECT 80.610 71.070 81.300 73.230 ;
        RECT 80.610 68.380 81.300 70.540 ;
        RECT 81.780 67.900 81.950 73.710 ;
        RECT 82.430 71.070 83.120 73.230 ;
        RECT 82.430 68.380 83.120 70.540 ;
        RECT 83.600 67.900 83.770 73.710 ;
        RECT 79.960 67.730 83.770 67.900 ;
        RECT 79.960 61.920 80.130 67.730 ;
        RECT 80.610 65.090 81.300 67.250 ;
        RECT 80.610 62.400 81.300 64.560 ;
        RECT 81.780 61.920 81.950 67.730 ;
        RECT 82.430 65.090 83.120 67.250 ;
        RECT 82.430 62.400 83.120 64.560 ;
        RECT 83.600 61.920 83.770 67.730 ;
        RECT 84.250 73.710 86.000 73.880 ;
        RECT 84.250 66.220 84.420 73.710 ;
        RECT 84.960 73.200 85.290 73.370 ;
        RECT 84.820 66.945 84.990 72.985 ;
        RECT 85.260 66.945 85.430 72.985 ;
        RECT 84.960 66.560 85.290 66.730 ;
        RECT 85.830 66.220 86.000 73.710 ;
        RECT 84.250 66.050 86.000 66.220 ;
        RECT 86.425 73.725 92.055 73.895 ;
        RECT 86.425 67.915 86.595 73.725 ;
        RECT 87.075 71.085 87.765 73.245 ;
        RECT 87.075 68.395 87.765 70.555 ;
        RECT 88.245 67.915 88.415 73.725 ;
        RECT 88.895 71.085 89.585 73.245 ;
        RECT 88.895 68.395 89.585 70.555 ;
        RECT 90.065 67.915 90.235 73.725 ;
        RECT 90.715 71.085 91.405 73.245 ;
        RECT 90.715 68.395 91.405 70.555 ;
        RECT 91.885 67.915 92.055 73.725 ;
        RECT 86.425 67.745 92.055 67.915 ;
        RECT 84.230 65.325 85.980 65.495 ;
        RECT 84.230 61.925 84.400 65.325 ;
        RECT 84.940 64.815 85.270 64.985 ;
        RECT 84.800 62.605 84.970 64.645 ;
        RECT 85.240 62.605 85.410 64.645 ;
        RECT 84.940 62.265 85.270 62.435 ;
        RECT 85.810 61.925 85.980 65.325 ;
        RECT 84.230 61.920 85.980 61.925 ;
        RECT 86.425 61.935 86.595 67.745 ;
        RECT 87.075 65.105 87.765 67.265 ;
        RECT 87.075 62.415 87.765 64.575 ;
        RECT 88.245 61.935 88.415 67.745 ;
        RECT 88.895 65.105 89.585 67.265 ;
        RECT 88.895 62.415 89.585 64.575 ;
        RECT 90.065 61.935 90.235 67.745 ;
        RECT 90.715 65.105 91.405 67.265 ;
        RECT 90.715 62.415 91.405 64.575 ;
        RECT 91.885 61.935 92.055 67.745 ;
        RECT 92.545 73.725 94.295 73.895 ;
        RECT 92.545 66.235 92.715 73.725 ;
        RECT 93.255 73.215 93.585 73.385 ;
        RECT 93.115 66.960 93.285 73.000 ;
        RECT 93.555 66.960 93.725 73.000 ;
        RECT 93.255 66.575 93.585 66.745 ;
        RECT 94.125 66.235 94.295 73.725 ;
        RECT 92.545 66.065 94.295 66.235 ;
        RECT 94.755 73.715 100.385 73.885 ;
        RECT 94.755 67.905 94.925 73.715 ;
        RECT 95.405 71.075 96.095 73.235 ;
        RECT 95.405 68.385 96.095 70.545 ;
        RECT 96.575 67.905 96.745 73.715 ;
        RECT 97.225 71.075 97.915 73.235 ;
        RECT 97.225 68.385 97.915 70.545 ;
        RECT 98.395 67.905 98.565 73.715 ;
        RECT 99.045 71.075 99.735 73.235 ;
        RECT 99.045 68.385 99.735 70.545 ;
        RECT 100.215 67.905 100.385 73.715 ;
        RECT 100.685 73.735 102.805 74.125 ;
        RECT 109.195 73.925 111.095 74.125 ;
        RECT 100.685 73.655 102.785 73.735 ;
        RECT 103.050 73.705 108.680 73.875 ;
        RECT 94.755 67.735 100.385 67.905 ;
        RECT 86.425 61.920 92.055 61.935 ;
        RECT 92.535 65.325 94.285 65.495 ;
        RECT 92.535 61.925 92.705 65.325 ;
        RECT 93.245 64.815 93.575 64.985 ;
        RECT 93.105 62.605 93.275 64.645 ;
        RECT 93.545 62.605 93.715 64.645 ;
        RECT 93.245 62.265 93.575 62.435 ;
        RECT 94.115 61.925 94.285 65.325 ;
        RECT 92.535 61.920 94.285 61.925 ;
        RECT 94.755 61.925 94.925 67.735 ;
        RECT 95.405 65.095 96.095 67.255 ;
        RECT 95.405 62.405 96.095 64.565 ;
        RECT 96.575 61.925 96.745 67.735 ;
        RECT 97.225 65.095 97.915 67.255 ;
        RECT 97.225 62.405 97.915 64.565 ;
        RECT 98.395 61.925 98.565 67.735 ;
        RECT 99.045 65.095 99.735 67.255 ;
        RECT 99.045 62.405 99.735 64.565 ;
        RECT 100.215 61.925 100.385 67.735 ;
        RECT 100.860 66.225 101.030 73.655 ;
        RECT 101.570 73.205 101.900 73.375 ;
        RECT 101.430 66.950 101.600 72.990 ;
        RECT 101.870 66.950 102.040 72.990 ;
        RECT 101.570 66.565 101.900 66.735 ;
        RECT 102.440 66.225 102.610 73.655 ;
        RECT 100.860 66.055 102.610 66.225 ;
        RECT 103.050 67.895 103.220 73.705 ;
        RECT 103.700 71.065 104.390 73.225 ;
        RECT 103.700 68.375 104.390 70.535 ;
        RECT 104.870 67.895 105.040 73.705 ;
        RECT 105.520 71.065 106.210 73.225 ;
        RECT 105.520 68.375 106.210 70.535 ;
        RECT 106.690 67.895 106.860 73.705 ;
        RECT 107.340 71.065 108.030 73.225 ;
        RECT 107.340 68.375 108.030 70.535 ;
        RECT 108.510 67.895 108.680 73.705 ;
        RECT 103.050 67.725 108.680 67.895 ;
        RECT 94.755 61.920 100.385 61.925 ;
        RECT 100.795 65.325 102.545 65.495 ;
        RECT 100.795 61.925 100.965 65.325 ;
        RECT 101.505 64.815 101.835 64.985 ;
        RECT 101.365 62.605 101.535 64.645 ;
        RECT 101.805 62.605 101.975 64.645 ;
        RECT 101.505 62.265 101.835 62.435 ;
        RECT 102.375 61.925 102.545 65.325 ;
        RECT 100.795 61.920 102.545 61.925 ;
        RECT 103.050 61.920 103.220 67.725 ;
        RECT 103.700 65.085 104.390 67.245 ;
        RECT 103.700 62.395 104.390 64.555 ;
        RECT 104.870 61.920 105.040 67.725 ;
        RECT 105.520 65.085 106.210 67.245 ;
        RECT 105.520 62.395 106.210 64.555 ;
        RECT 106.690 61.920 106.860 67.725 ;
        RECT 107.340 65.085 108.030 67.245 ;
        RECT 107.340 62.395 108.030 64.555 ;
        RECT 108.510 61.920 108.680 67.725 ;
        RECT 109.240 73.815 110.990 73.925 ;
        RECT 117.635 73.910 119.345 74.125 ;
        RECT 125.965 73.935 127.675 74.125 ;
        RECT 134.255 73.950 135.965 74.125 ;
        RECT 109.240 66.325 109.410 73.815 ;
        RECT 109.950 73.305 110.280 73.475 ;
        RECT 109.810 67.050 109.980 73.090 ;
        RECT 110.250 67.050 110.420 73.090 ;
        RECT 109.950 66.665 110.280 66.835 ;
        RECT 110.820 66.325 110.990 73.815 ;
        RECT 109.240 66.155 110.990 66.325 ;
        RECT 111.495 73.720 117.125 73.890 ;
        RECT 111.495 67.910 111.665 73.720 ;
        RECT 112.145 71.080 112.835 73.240 ;
        RECT 112.145 68.390 112.835 70.550 ;
        RECT 113.315 67.910 113.485 73.720 ;
        RECT 113.965 71.080 114.655 73.240 ;
        RECT 113.965 68.390 114.655 70.550 ;
        RECT 115.135 67.910 115.305 73.720 ;
        RECT 115.785 71.080 116.475 73.240 ;
        RECT 115.785 68.390 116.475 70.550 ;
        RECT 116.955 67.910 117.125 73.720 ;
        RECT 111.495 67.740 117.125 67.910 ;
        RECT 109.215 65.345 110.965 65.515 ;
        RECT 109.215 61.945 109.385 65.345 ;
        RECT 109.925 64.835 110.255 65.005 ;
        RECT 109.785 62.625 109.955 64.665 ;
        RECT 110.225 62.625 110.395 64.665 ;
        RECT 109.925 62.285 110.255 62.455 ;
        RECT 110.795 61.945 110.965 65.345 ;
        RECT 109.215 61.920 110.965 61.945 ;
        RECT 111.495 61.930 111.665 67.740 ;
        RECT 112.145 65.100 112.835 67.260 ;
        RECT 112.145 62.410 112.835 64.570 ;
        RECT 113.315 61.930 113.485 67.740 ;
        RECT 113.965 65.100 114.655 67.260 ;
        RECT 113.965 62.410 114.655 64.570 ;
        RECT 115.135 61.930 115.305 67.740 ;
        RECT 115.785 65.100 116.475 67.260 ;
        RECT 115.785 62.410 116.475 64.570 ;
        RECT 116.955 61.930 117.125 67.740 ;
        RECT 117.630 73.740 119.380 73.910 ;
        RECT 117.630 66.250 117.800 73.740 ;
        RECT 118.340 73.230 118.670 73.400 ;
        RECT 118.200 66.975 118.370 73.015 ;
        RECT 118.640 66.975 118.810 73.015 ;
        RECT 118.340 66.590 118.670 66.760 ;
        RECT 119.210 66.250 119.380 73.740 ;
        RECT 117.630 66.080 119.380 66.250 ;
        RECT 119.825 73.720 125.455 73.890 ;
        RECT 119.825 67.910 119.995 73.720 ;
        RECT 120.475 71.080 121.165 73.240 ;
        RECT 120.475 68.390 121.165 70.550 ;
        RECT 121.645 67.910 121.815 73.720 ;
        RECT 122.295 71.080 122.985 73.240 ;
        RECT 122.295 68.390 122.985 70.550 ;
        RECT 123.465 67.910 123.635 73.720 ;
        RECT 124.115 71.080 124.805 73.240 ;
        RECT 124.115 68.390 124.805 70.550 ;
        RECT 125.285 67.910 125.455 73.720 ;
        RECT 119.825 67.740 125.455 67.910 ;
        RECT 111.495 61.920 117.125 61.930 ;
        RECT 117.565 65.325 119.315 65.495 ;
        RECT 117.565 61.925 117.735 65.325 ;
        RECT 118.275 64.815 118.605 64.985 ;
        RECT 118.135 62.605 118.305 64.645 ;
        RECT 118.575 62.605 118.745 64.645 ;
        RECT 118.275 62.265 118.605 62.435 ;
        RECT 119.145 61.925 119.315 65.325 ;
        RECT 117.565 61.920 119.315 61.925 ;
        RECT 119.825 61.930 119.995 67.740 ;
        RECT 120.475 65.100 121.165 67.260 ;
        RECT 120.475 62.410 121.165 64.570 ;
        RECT 121.645 61.930 121.815 67.740 ;
        RECT 122.295 65.100 122.985 67.260 ;
        RECT 122.295 62.410 122.985 64.570 ;
        RECT 123.465 61.930 123.635 67.740 ;
        RECT 124.115 65.100 124.805 67.260 ;
        RECT 124.115 62.410 124.805 64.570 ;
        RECT 125.285 61.930 125.455 67.740 ;
        RECT 125.960 73.765 127.710 73.935 ;
        RECT 125.960 66.275 126.130 73.765 ;
        RECT 126.670 73.255 127.000 73.425 ;
        RECT 126.530 67.000 126.700 73.040 ;
        RECT 126.970 67.000 127.140 73.040 ;
        RECT 126.670 66.615 127.000 66.785 ;
        RECT 127.540 66.275 127.710 73.765 ;
        RECT 125.960 66.105 127.710 66.275 ;
        RECT 128.155 73.720 133.785 73.890 ;
        RECT 128.155 67.910 128.325 73.720 ;
        RECT 128.805 71.080 129.495 73.240 ;
        RECT 128.805 68.390 129.495 70.550 ;
        RECT 129.975 67.910 130.145 73.720 ;
        RECT 130.625 71.080 131.315 73.240 ;
        RECT 130.625 68.390 131.315 70.550 ;
        RECT 131.795 67.910 131.965 73.720 ;
        RECT 132.445 71.080 133.135 73.240 ;
        RECT 132.445 68.390 133.135 70.550 ;
        RECT 133.615 67.910 133.785 73.720 ;
        RECT 128.155 67.740 133.785 67.910 ;
        RECT 119.825 61.920 125.455 61.930 ;
        RECT 125.950 65.320 127.700 65.490 ;
        RECT 125.950 61.920 126.120 65.320 ;
        RECT 126.660 64.810 126.990 64.980 ;
        RECT 126.520 62.600 126.690 64.640 ;
        RECT 126.960 62.600 127.130 64.640 ;
        RECT 126.660 62.260 126.990 62.430 ;
        RECT 127.530 61.920 127.700 65.320 ;
        RECT 128.155 61.930 128.325 67.740 ;
        RECT 128.805 65.100 129.495 67.260 ;
        RECT 128.805 62.410 129.495 64.570 ;
        RECT 129.975 61.930 130.145 67.740 ;
        RECT 130.625 65.100 131.315 67.260 ;
        RECT 130.625 62.410 131.315 64.570 ;
        RECT 131.795 61.930 131.965 67.740 ;
        RECT 132.445 65.100 133.135 67.260 ;
        RECT 132.445 62.410 133.135 64.570 ;
        RECT 133.615 61.930 133.785 67.740 ;
        RECT 134.255 73.780 136.005 73.950 ;
        RECT 142.585 73.930 144.295 74.125 ;
        RECT 134.255 66.290 134.425 73.780 ;
        RECT 134.965 73.270 135.295 73.440 ;
        RECT 134.825 67.015 134.995 73.055 ;
        RECT 135.265 67.015 135.435 73.055 ;
        RECT 134.965 66.630 135.295 66.800 ;
        RECT 135.835 66.290 136.005 73.780 ;
        RECT 134.255 66.120 136.005 66.290 ;
        RECT 136.460 73.715 142.090 73.885 ;
        RECT 136.460 67.905 136.630 73.715 ;
        RECT 137.110 71.075 137.800 73.235 ;
        RECT 137.110 68.385 137.800 70.545 ;
        RECT 138.280 67.905 138.450 73.715 ;
        RECT 138.930 71.075 139.620 73.235 ;
        RECT 138.930 68.385 139.620 70.545 ;
        RECT 140.100 67.905 140.270 73.715 ;
        RECT 140.750 71.075 141.440 73.235 ;
        RECT 140.750 68.385 141.440 70.545 ;
        RECT 141.920 67.905 142.090 73.715 ;
        RECT 136.460 67.735 142.090 67.905 ;
        RECT 128.155 61.920 133.785 61.930 ;
        RECT 134.190 65.330 135.940 65.500 ;
        RECT 134.190 61.930 134.360 65.330 ;
        RECT 134.900 64.820 135.230 64.990 ;
        RECT 134.760 62.610 134.930 64.650 ;
        RECT 135.200 62.610 135.370 64.650 ;
        RECT 134.900 62.270 135.230 62.440 ;
        RECT 135.770 61.930 135.940 65.330 ;
        RECT 134.190 61.920 135.940 61.930 ;
        RECT 136.460 61.925 136.630 67.735 ;
        RECT 137.110 65.095 137.800 67.255 ;
        RECT 137.110 62.405 137.800 64.565 ;
        RECT 138.280 61.925 138.450 67.735 ;
        RECT 138.930 65.095 139.620 67.255 ;
        RECT 138.930 62.405 139.620 64.565 ;
        RECT 140.100 61.925 140.270 67.735 ;
        RECT 140.750 65.095 141.440 67.255 ;
        RECT 140.750 62.405 141.440 64.565 ;
        RECT 141.920 61.925 142.090 67.735 ;
        RECT 142.555 73.760 144.305 73.930 ;
        RECT 142.555 66.270 142.725 73.760 ;
        RECT 143.265 73.250 143.595 73.420 ;
        RECT 143.125 66.995 143.295 73.035 ;
        RECT 143.565 66.995 143.735 73.035 ;
        RECT 143.265 66.610 143.595 66.780 ;
        RECT 144.135 66.270 144.305 73.760 ;
        RECT 142.555 66.100 144.305 66.270 ;
        RECT 144.760 73.725 148.570 73.895 ;
        RECT 144.760 67.915 144.930 73.725 ;
        RECT 145.410 71.085 146.100 73.245 ;
        RECT 145.410 68.395 146.100 70.555 ;
        RECT 146.580 67.915 146.750 73.725 ;
        RECT 147.230 71.085 147.920 73.245 ;
        RECT 147.230 68.395 147.920 70.555 ;
        RECT 148.400 67.915 148.570 73.725 ;
        RECT 144.760 67.745 148.570 67.915 ;
        RECT 136.460 61.920 142.090 61.925 ;
        RECT 142.555 65.330 144.305 65.500 ;
        RECT 142.555 61.930 142.725 65.330 ;
        RECT 143.265 64.820 143.595 64.990 ;
        RECT 143.125 62.610 143.295 64.650 ;
        RECT 143.565 62.610 143.735 64.650 ;
        RECT 143.265 62.270 143.595 62.440 ;
        RECT 144.135 61.930 144.305 65.330 ;
        RECT 142.555 61.920 144.305 61.930 ;
        RECT 144.760 61.935 144.930 67.745 ;
        RECT 145.410 65.105 146.100 67.265 ;
        RECT 145.410 62.415 146.100 64.575 ;
        RECT 146.580 61.935 146.750 67.745 ;
        RECT 147.230 65.105 147.920 67.265 ;
        RECT 147.230 62.415 147.920 64.575 ;
        RECT 148.400 61.935 148.570 67.745 ;
        RECT 144.760 61.920 148.570 61.935 ;
        RECT 79.960 61.045 148.575 61.920 ;
        RECT 1.890 57.840 14.020 58.010 ;
        RECT 1.890 56.190 2.060 57.840 ;
        RECT 2.540 56.670 4.700 57.360 ;
        RECT 5.230 56.670 7.390 57.360 ;
        RECT 7.870 56.190 8.040 57.840 ;
        RECT 8.520 56.670 10.680 57.360 ;
        RECT 11.210 56.670 13.370 57.360 ;
        RECT 13.850 56.190 14.020 57.840 ;
        RECT 1.890 56.020 14.020 56.190 ;
        RECT 1.890 54.370 2.060 56.020 ;
        RECT 2.540 54.850 4.700 55.540 ;
        RECT 5.230 54.850 7.390 55.540 ;
        RECT 7.870 54.370 8.040 56.020 ;
        RECT 8.520 54.850 10.680 55.540 ;
        RECT 11.210 54.850 13.370 55.540 ;
        RECT 13.850 54.370 14.020 56.020 ;
        RECT 1.890 54.200 14.020 54.370 ;
        RECT 1.890 52.550 2.060 54.200 ;
        RECT 2.540 53.030 4.700 53.720 ;
        RECT 5.230 53.030 7.390 53.720 ;
        RECT 7.870 52.550 8.040 54.200 ;
        RECT 8.520 53.030 10.680 53.720 ;
        RECT 11.210 53.030 13.370 53.720 ;
        RECT 13.850 52.550 14.020 54.200 ;
        RECT 1.890 52.380 31.960 52.550 ;
        RECT 1.890 50.855 2.060 52.380 ;
        RECT 2.540 51.210 4.700 51.900 ;
        RECT 5.230 51.210 7.390 51.900 ;
        RECT 7.870 50.855 8.040 52.380 ;
        RECT 8.520 51.210 10.680 51.900 ;
        RECT 11.210 51.210 13.370 51.900 ;
        RECT 1.890 50.730 10.380 50.855 ;
        RECT 13.850 50.730 14.020 52.380 ;
        RECT 14.500 51.210 16.660 51.900 ;
        RECT 17.190 51.210 19.350 51.900 ;
        RECT 19.830 50.730 20.000 52.380 ;
        RECT 20.480 51.210 22.640 51.900 ;
        RECT 23.170 51.210 25.330 51.900 ;
        RECT 25.810 50.730 25.980 52.380 ;
        RECT 26.460 51.210 28.620 51.900 ;
        RECT 29.150 51.210 31.310 51.900 ;
        RECT 31.790 50.730 31.960 52.380 ;
        RECT 1.890 50.560 31.960 50.730 ;
        RECT 43.910 52.540 62.020 52.550 ;
        RECT 67.910 52.540 86.020 52.550 ;
        RECT 43.910 52.380 86.020 52.540 ;
        RECT 43.910 50.730 44.080 52.380 ;
        RECT 44.560 51.210 46.720 51.900 ;
        RECT 47.250 51.210 49.410 51.900 ;
        RECT 49.890 50.730 50.060 52.380 ;
        RECT 50.540 51.210 52.700 51.900 ;
        RECT 53.230 51.210 55.390 51.900 ;
        RECT 55.870 50.730 56.040 52.380 ;
        RECT 61.850 52.090 68.090 52.380 ;
        RECT 56.520 51.210 58.680 51.900 ;
        RECT 59.210 51.210 61.370 51.900 ;
        RECT 61.850 50.730 62.020 52.090 ;
        RECT 43.910 50.560 62.020 50.730 ;
        RECT 67.910 50.730 68.080 52.090 ;
        RECT 68.560 51.210 70.720 51.900 ;
        RECT 71.250 51.210 73.410 51.900 ;
        RECT 73.890 50.730 74.060 52.380 ;
        RECT 74.540 51.210 76.700 51.900 ;
        RECT 77.230 51.210 79.390 51.900 ;
        RECT 79.870 50.730 80.040 52.380 ;
        RECT 80.520 51.210 82.680 51.900 ;
        RECT 83.210 51.210 85.370 51.900 ;
        RECT 85.850 50.730 86.020 52.380 ;
        RECT 67.910 50.560 86.020 50.730 ;
        RECT 2.005 50.360 10.380 50.560 ;
        RECT 78.210 50.170 80.780 50.560 ;
        RECT 1.870 49.480 28.345 49.960 ;
        RECT 29.870 49.480 56.345 49.960 ;
        RECT 57.870 49.480 84.345 49.960 ;
        RECT 85.870 49.480 112.345 49.960 ;
        RECT 113.870 49.480 140.345 49.960 ;
        RECT 1.855 49.420 28.345 49.480 ;
        RECT 29.855 49.420 56.345 49.480 ;
        RECT 57.855 49.420 84.345 49.480 ;
        RECT 85.855 49.420 112.345 49.480 ;
        RECT 113.855 49.420 140.345 49.480 ;
        RECT 143.890 49.840 150.040 50.010 ;
        RECT 1.855 49.260 28.400 49.420 ;
        RECT 1.855 49.235 14.600 49.260 ;
        RECT 1.855 49.005 6.180 49.235 ;
        RECT 1.890 39.745 2.060 49.005 ;
        RECT 2.785 48.435 4.825 48.605 ;
        RECT 2.400 40.375 2.570 48.375 ;
        RECT 5.040 40.375 5.210 48.375 ;
        RECT 2.785 40.145 4.825 40.315 ;
        RECT 5.550 39.745 5.720 49.005 ;
        RECT 1.890 39.575 5.720 39.745 ;
        RECT 6.010 39.745 6.180 49.005 ;
        RECT 6.810 48.725 8.810 48.895 ;
        RECT 6.580 40.470 6.750 48.510 ;
        RECT 8.870 40.470 9.040 48.510 ;
        RECT 6.810 40.085 8.810 40.255 ;
        RECT 9.440 39.745 9.610 49.235 ;
        RECT 10.240 48.725 12.240 48.895 ;
        RECT 10.010 40.470 10.180 48.510 ;
        RECT 12.300 40.470 12.470 48.510 ;
        RECT 12.870 47.665 14.600 49.235 ;
        RECT 26.650 49.250 28.400 49.260 ;
        RECT 12.870 47.495 21.335 47.665 ;
        RECT 12.870 46.085 14.675 47.495 ;
        RECT 15.015 46.625 15.185 46.955 ;
        RECT 15.400 46.925 20.440 47.095 ;
        RECT 15.400 46.485 20.440 46.655 ;
        RECT 20.655 46.625 20.825 46.955 ;
        RECT 21.165 46.085 21.335 47.495 ;
        RECT 12.870 45.915 21.335 46.085 ;
        RECT 12.870 45.400 14.600 45.915 ;
        RECT 12.870 45.285 24.350 45.400 ;
        RECT 10.240 40.085 12.240 40.255 ;
        RECT 12.870 39.745 13.040 45.285 ;
        RECT 6.010 39.575 13.040 39.745 ;
        RECT 13.320 45.230 24.350 45.285 ;
        RECT 13.320 39.740 13.490 45.230 ;
        RECT 14.120 44.720 18.120 44.890 ;
        RECT 13.890 40.465 14.060 44.505 ;
        RECT 18.180 40.465 18.350 44.505 ;
        RECT 14.120 40.080 18.120 40.250 ;
        RECT 18.750 39.740 18.920 45.230 ;
        RECT 19.550 44.720 23.550 44.890 ;
        RECT 19.320 40.465 19.490 44.505 ;
        RECT 23.610 40.465 23.780 44.505 ;
        RECT 19.550 40.080 23.550 40.250 ;
        RECT 24.180 39.740 24.350 45.230 ;
        RECT 13.320 39.570 24.350 39.740 ;
        RECT 24.625 45.245 26.375 45.415 ;
        RECT 24.625 39.755 24.795 45.245 ;
        RECT 25.335 44.735 25.665 44.905 ;
        RECT 25.195 40.480 25.365 44.520 ;
        RECT 25.635 40.480 25.805 44.520 ;
        RECT 25.335 40.095 25.665 40.265 ;
        RECT 26.205 39.755 26.375 45.245 ;
        RECT 24.625 39.585 26.375 39.755 ;
        RECT 26.650 39.760 26.820 49.250 ;
        RECT 27.360 48.740 27.690 48.910 ;
        RECT 27.220 40.485 27.390 48.525 ;
        RECT 27.660 40.485 27.830 48.525 ;
        RECT 27.360 40.100 27.690 40.270 ;
        RECT 28.230 39.760 28.400 49.250 ;
        RECT 29.855 49.260 56.400 49.420 ;
        RECT 29.855 49.235 42.600 49.260 ;
        RECT 29.855 49.005 34.180 49.235 ;
        RECT 26.650 39.590 28.400 39.760 ;
        RECT 29.890 39.745 30.060 49.005 ;
        RECT 30.785 48.435 32.825 48.605 ;
        RECT 30.400 40.375 30.570 48.375 ;
        RECT 33.040 40.375 33.210 48.375 ;
        RECT 30.785 40.145 32.825 40.315 ;
        RECT 33.550 39.745 33.720 49.005 ;
        RECT 29.890 39.575 33.720 39.745 ;
        RECT 34.010 39.745 34.180 49.005 ;
        RECT 34.810 48.725 36.810 48.895 ;
        RECT 34.580 40.470 34.750 48.510 ;
        RECT 36.870 40.470 37.040 48.510 ;
        RECT 34.810 40.085 36.810 40.255 ;
        RECT 37.440 39.745 37.610 49.235 ;
        RECT 38.240 48.725 40.240 48.895 ;
        RECT 38.010 40.470 38.180 48.510 ;
        RECT 40.300 40.470 40.470 48.510 ;
        RECT 40.870 47.665 42.600 49.235 ;
        RECT 54.650 49.250 56.400 49.260 ;
        RECT 40.870 47.495 49.335 47.665 ;
        RECT 40.870 46.085 42.675 47.495 ;
        RECT 43.015 46.625 43.185 46.955 ;
        RECT 43.400 46.925 48.440 47.095 ;
        RECT 43.400 46.485 48.440 46.655 ;
        RECT 48.655 46.625 48.825 46.955 ;
        RECT 49.165 46.085 49.335 47.495 ;
        RECT 40.870 45.915 49.335 46.085 ;
        RECT 40.870 45.400 42.600 45.915 ;
        RECT 40.870 45.285 52.350 45.400 ;
        RECT 38.240 40.085 40.240 40.255 ;
        RECT 40.870 39.745 41.040 45.285 ;
        RECT 34.010 39.575 41.040 39.745 ;
        RECT 41.320 45.230 52.350 45.285 ;
        RECT 41.320 39.740 41.490 45.230 ;
        RECT 42.120 44.720 46.120 44.890 ;
        RECT 41.890 40.465 42.060 44.505 ;
        RECT 46.180 40.465 46.350 44.505 ;
        RECT 42.120 40.080 46.120 40.250 ;
        RECT 46.750 39.740 46.920 45.230 ;
        RECT 47.550 44.720 51.550 44.890 ;
        RECT 47.320 40.465 47.490 44.505 ;
        RECT 51.610 40.465 51.780 44.505 ;
        RECT 47.550 40.080 51.550 40.250 ;
        RECT 52.180 39.740 52.350 45.230 ;
        RECT 41.320 39.570 52.350 39.740 ;
        RECT 52.625 45.245 54.375 45.415 ;
        RECT 52.625 39.755 52.795 45.245 ;
        RECT 53.335 44.735 53.665 44.905 ;
        RECT 53.195 40.480 53.365 44.520 ;
        RECT 53.635 40.480 53.805 44.520 ;
        RECT 53.335 40.095 53.665 40.265 ;
        RECT 54.205 39.755 54.375 45.245 ;
        RECT 52.625 39.585 54.375 39.755 ;
        RECT 54.650 39.760 54.820 49.250 ;
        RECT 55.360 48.740 55.690 48.910 ;
        RECT 55.220 40.485 55.390 48.525 ;
        RECT 55.660 40.485 55.830 48.525 ;
        RECT 55.360 40.100 55.690 40.270 ;
        RECT 56.230 39.760 56.400 49.250 ;
        RECT 57.855 49.260 84.400 49.420 ;
        RECT 57.855 49.235 70.600 49.260 ;
        RECT 57.855 49.005 62.180 49.235 ;
        RECT 54.650 39.590 56.400 39.760 ;
        RECT 57.890 39.745 58.060 49.005 ;
        RECT 58.785 48.435 60.825 48.605 ;
        RECT 58.400 40.375 58.570 48.375 ;
        RECT 61.040 40.375 61.210 48.375 ;
        RECT 58.785 40.145 60.825 40.315 ;
        RECT 61.550 39.745 61.720 49.005 ;
        RECT 57.890 39.575 61.720 39.745 ;
        RECT 62.010 39.745 62.180 49.005 ;
        RECT 62.810 48.725 64.810 48.895 ;
        RECT 62.580 40.470 62.750 48.510 ;
        RECT 64.870 40.470 65.040 48.510 ;
        RECT 62.810 40.085 64.810 40.255 ;
        RECT 65.440 39.745 65.610 49.235 ;
        RECT 66.240 48.725 68.240 48.895 ;
        RECT 66.010 40.470 66.180 48.510 ;
        RECT 68.300 40.470 68.470 48.510 ;
        RECT 68.870 47.665 70.600 49.235 ;
        RECT 82.650 49.250 84.400 49.260 ;
        RECT 68.870 47.495 77.335 47.665 ;
        RECT 68.870 46.085 70.675 47.495 ;
        RECT 71.015 46.625 71.185 46.955 ;
        RECT 71.400 46.925 76.440 47.095 ;
        RECT 71.400 46.485 76.440 46.655 ;
        RECT 76.655 46.625 76.825 46.955 ;
        RECT 77.165 46.085 77.335 47.495 ;
        RECT 68.870 45.915 77.335 46.085 ;
        RECT 68.870 45.400 70.600 45.915 ;
        RECT 68.870 45.285 80.350 45.400 ;
        RECT 66.240 40.085 68.240 40.255 ;
        RECT 68.870 39.745 69.040 45.285 ;
        RECT 62.010 39.575 69.040 39.745 ;
        RECT 69.320 45.230 80.350 45.285 ;
        RECT 69.320 39.740 69.490 45.230 ;
        RECT 70.120 44.720 74.120 44.890 ;
        RECT 69.890 40.465 70.060 44.505 ;
        RECT 74.180 40.465 74.350 44.505 ;
        RECT 70.120 40.080 74.120 40.250 ;
        RECT 74.750 39.740 74.920 45.230 ;
        RECT 75.550 44.720 79.550 44.890 ;
        RECT 75.320 40.465 75.490 44.505 ;
        RECT 79.610 40.465 79.780 44.505 ;
        RECT 75.550 40.080 79.550 40.250 ;
        RECT 80.180 39.740 80.350 45.230 ;
        RECT 69.320 39.570 80.350 39.740 ;
        RECT 80.625 45.245 82.375 45.415 ;
        RECT 80.625 39.755 80.795 45.245 ;
        RECT 81.335 44.735 81.665 44.905 ;
        RECT 81.195 40.480 81.365 44.520 ;
        RECT 81.635 40.480 81.805 44.520 ;
        RECT 81.335 40.095 81.665 40.265 ;
        RECT 82.205 39.755 82.375 45.245 ;
        RECT 80.625 39.585 82.375 39.755 ;
        RECT 82.650 39.760 82.820 49.250 ;
        RECT 83.360 48.740 83.690 48.910 ;
        RECT 83.220 40.485 83.390 48.525 ;
        RECT 83.660 40.485 83.830 48.525 ;
        RECT 83.360 40.100 83.690 40.270 ;
        RECT 84.230 39.760 84.400 49.250 ;
        RECT 85.855 49.260 112.400 49.420 ;
        RECT 85.855 49.235 98.600 49.260 ;
        RECT 85.855 49.005 90.180 49.235 ;
        RECT 82.650 39.590 84.400 39.760 ;
        RECT 85.890 39.745 86.060 49.005 ;
        RECT 86.785 48.435 88.825 48.605 ;
        RECT 86.400 40.375 86.570 48.375 ;
        RECT 89.040 40.375 89.210 48.375 ;
        RECT 86.785 40.145 88.825 40.315 ;
        RECT 89.550 39.745 89.720 49.005 ;
        RECT 85.890 39.575 89.720 39.745 ;
        RECT 90.010 39.745 90.180 49.005 ;
        RECT 90.810 48.725 92.810 48.895 ;
        RECT 90.580 40.470 90.750 48.510 ;
        RECT 92.870 40.470 93.040 48.510 ;
        RECT 90.810 40.085 92.810 40.255 ;
        RECT 93.440 39.745 93.610 49.235 ;
        RECT 94.240 48.725 96.240 48.895 ;
        RECT 94.010 40.470 94.180 48.510 ;
        RECT 96.300 40.470 96.470 48.510 ;
        RECT 96.870 47.665 98.600 49.235 ;
        RECT 110.650 49.250 112.400 49.260 ;
        RECT 96.870 47.495 105.335 47.665 ;
        RECT 96.870 46.085 98.675 47.495 ;
        RECT 99.015 46.625 99.185 46.955 ;
        RECT 99.400 46.925 104.440 47.095 ;
        RECT 99.400 46.485 104.440 46.655 ;
        RECT 104.655 46.625 104.825 46.955 ;
        RECT 105.165 46.085 105.335 47.495 ;
        RECT 96.870 45.915 105.335 46.085 ;
        RECT 96.870 45.400 98.600 45.915 ;
        RECT 96.870 45.285 108.350 45.400 ;
        RECT 94.240 40.085 96.240 40.255 ;
        RECT 96.870 39.745 97.040 45.285 ;
        RECT 90.010 39.575 97.040 39.745 ;
        RECT 97.320 45.230 108.350 45.285 ;
        RECT 97.320 39.740 97.490 45.230 ;
        RECT 98.120 44.720 102.120 44.890 ;
        RECT 97.890 40.465 98.060 44.505 ;
        RECT 102.180 40.465 102.350 44.505 ;
        RECT 98.120 40.080 102.120 40.250 ;
        RECT 102.750 39.740 102.920 45.230 ;
        RECT 103.550 44.720 107.550 44.890 ;
        RECT 103.320 40.465 103.490 44.505 ;
        RECT 107.610 40.465 107.780 44.505 ;
        RECT 103.550 40.080 107.550 40.250 ;
        RECT 108.180 39.740 108.350 45.230 ;
        RECT 97.320 39.570 108.350 39.740 ;
        RECT 108.625 45.245 110.375 45.415 ;
        RECT 108.625 39.755 108.795 45.245 ;
        RECT 109.335 44.735 109.665 44.905 ;
        RECT 109.195 40.480 109.365 44.520 ;
        RECT 109.635 40.480 109.805 44.520 ;
        RECT 109.335 40.095 109.665 40.265 ;
        RECT 110.205 39.755 110.375 45.245 ;
        RECT 108.625 39.585 110.375 39.755 ;
        RECT 110.650 39.760 110.820 49.250 ;
        RECT 111.360 48.740 111.690 48.910 ;
        RECT 111.220 40.485 111.390 48.525 ;
        RECT 111.660 40.485 111.830 48.525 ;
        RECT 111.360 40.100 111.690 40.270 ;
        RECT 112.230 39.760 112.400 49.250 ;
        RECT 113.855 49.260 140.400 49.420 ;
        RECT 113.855 49.235 126.600 49.260 ;
        RECT 113.855 49.005 118.180 49.235 ;
        RECT 110.650 39.590 112.400 39.760 ;
        RECT 113.890 39.745 114.060 49.005 ;
        RECT 114.785 48.435 116.825 48.605 ;
        RECT 114.400 40.375 114.570 48.375 ;
        RECT 117.040 40.375 117.210 48.375 ;
        RECT 114.785 40.145 116.825 40.315 ;
        RECT 117.550 39.745 117.720 49.005 ;
        RECT 113.890 39.575 117.720 39.745 ;
        RECT 118.010 39.745 118.180 49.005 ;
        RECT 118.810 48.725 120.810 48.895 ;
        RECT 118.580 40.470 118.750 48.510 ;
        RECT 120.870 40.470 121.040 48.510 ;
        RECT 118.810 40.085 120.810 40.255 ;
        RECT 121.440 39.745 121.610 49.235 ;
        RECT 122.240 48.725 124.240 48.895 ;
        RECT 122.010 40.470 122.180 48.510 ;
        RECT 124.300 40.470 124.470 48.510 ;
        RECT 124.870 47.665 126.600 49.235 ;
        RECT 138.650 49.250 140.400 49.260 ;
        RECT 124.870 47.495 133.335 47.665 ;
        RECT 124.870 46.085 126.675 47.495 ;
        RECT 127.015 46.625 127.185 46.955 ;
        RECT 127.400 46.925 132.440 47.095 ;
        RECT 127.400 46.485 132.440 46.655 ;
        RECT 132.655 46.625 132.825 46.955 ;
        RECT 133.165 46.085 133.335 47.495 ;
        RECT 124.870 45.915 133.335 46.085 ;
        RECT 124.870 45.400 126.600 45.915 ;
        RECT 124.870 45.285 136.350 45.400 ;
        RECT 122.240 40.085 124.240 40.255 ;
        RECT 124.870 39.745 125.040 45.285 ;
        RECT 118.010 39.575 125.040 39.745 ;
        RECT 125.320 45.230 136.350 45.285 ;
        RECT 125.320 39.740 125.490 45.230 ;
        RECT 126.120 44.720 130.120 44.890 ;
        RECT 125.890 40.465 126.060 44.505 ;
        RECT 130.180 40.465 130.350 44.505 ;
        RECT 126.120 40.080 130.120 40.250 ;
        RECT 130.750 39.740 130.920 45.230 ;
        RECT 131.550 44.720 135.550 44.890 ;
        RECT 131.320 40.465 131.490 44.505 ;
        RECT 135.610 40.465 135.780 44.505 ;
        RECT 131.550 40.080 135.550 40.250 ;
        RECT 136.180 39.740 136.350 45.230 ;
        RECT 125.320 39.570 136.350 39.740 ;
        RECT 136.625 45.245 138.375 45.415 ;
        RECT 136.625 39.755 136.795 45.245 ;
        RECT 137.335 44.735 137.665 44.905 ;
        RECT 137.195 40.480 137.365 44.520 ;
        RECT 137.635 40.480 137.805 44.520 ;
        RECT 137.335 40.095 137.665 40.265 ;
        RECT 138.205 39.755 138.375 45.245 ;
        RECT 136.625 39.585 138.375 39.755 ;
        RECT 138.650 39.760 138.820 49.250 ;
        RECT 139.360 48.740 139.690 48.910 ;
        RECT 139.220 40.485 139.390 48.525 ;
        RECT 139.660 40.485 139.830 48.525 ;
        RECT 139.360 40.100 139.690 40.270 ;
        RECT 140.230 39.760 140.400 49.250 ;
        RECT 143.890 48.190 144.060 49.840 ;
        RECT 144.540 48.670 146.700 49.360 ;
        RECT 147.230 48.670 149.390 49.360 ;
        RECT 149.870 48.190 150.040 49.840 ;
        RECT 143.890 48.020 150.040 48.190 ;
        RECT 143.890 46.370 144.060 48.020 ;
        RECT 144.540 46.850 146.700 47.540 ;
        RECT 147.230 46.850 149.390 47.540 ;
        RECT 149.870 46.370 150.040 48.020 ;
        RECT 143.890 46.200 150.040 46.370 ;
        RECT 143.890 44.550 144.060 46.200 ;
        RECT 144.540 45.030 146.700 45.720 ;
        RECT 147.230 45.030 149.390 45.720 ;
        RECT 149.870 44.550 150.040 46.200 ;
        RECT 143.890 44.380 156.020 44.550 ;
        RECT 143.890 42.730 144.060 44.380 ;
        RECT 144.540 43.210 146.700 43.900 ;
        RECT 147.230 43.210 149.390 43.900 ;
        RECT 149.870 42.730 150.040 44.380 ;
        RECT 150.520 43.210 152.680 43.900 ;
        RECT 153.210 43.210 155.370 43.900 ;
        RECT 155.850 42.730 156.020 44.380 ;
        RECT 143.890 42.560 156.020 42.730 ;
        RECT 143.890 40.910 144.060 42.560 ;
        RECT 144.540 41.390 146.700 42.080 ;
        RECT 147.230 41.390 149.390 42.080 ;
        RECT 149.870 40.910 150.040 42.560 ;
        RECT 150.520 41.390 152.680 42.080 ;
        RECT 153.210 41.390 155.370 42.080 ;
        RECT 155.850 40.910 156.020 42.560 ;
        RECT 143.890 40.740 156.020 40.910 ;
        RECT 151.200 40.250 154.760 40.740 ;
        RECT 138.650 39.590 140.400 39.760 ;
        RECT 2.550 38.665 24.440 38.835 ;
        RECT 2.550 35.265 2.720 38.665 ;
        RECT 3.350 38.155 7.350 38.325 ;
        RECT 3.120 35.945 3.290 37.985 ;
        RECT 7.410 35.945 7.580 37.985 ;
        RECT 3.350 35.605 7.350 35.775 ;
        RECT 7.980 35.265 8.150 38.665 ;
        RECT 8.780 38.155 12.780 38.325 ;
        RECT 8.550 35.945 8.720 37.985 ;
        RECT 12.840 35.945 13.010 37.985 ;
        RECT 8.780 35.605 12.780 35.775 ;
        RECT 13.410 35.265 13.580 38.665 ;
        RECT 14.210 38.155 18.210 38.325 ;
        RECT 13.980 35.945 14.150 37.985 ;
        RECT 18.270 35.945 18.440 37.985 ;
        RECT 14.210 35.605 18.210 35.775 ;
        RECT 18.840 35.265 19.010 38.665 ;
        RECT 19.640 38.155 23.640 38.325 ;
        RECT 19.410 35.945 19.580 37.985 ;
        RECT 23.700 35.945 23.870 37.985 ;
        RECT 24.270 36.240 24.440 38.665 ;
        RECT 24.710 38.670 26.460 38.840 ;
        RECT 24.710 36.270 24.880 38.670 ;
        RECT 25.420 38.160 25.750 38.330 ;
        RECT 25.280 36.950 25.450 37.990 ;
        RECT 25.720 36.950 25.890 37.990 ;
        RECT 25.420 36.610 25.750 36.780 ;
        RECT 26.290 36.270 26.460 38.670 ;
        RECT 24.710 36.240 26.460 36.270 ;
        RECT 26.735 38.675 28.485 38.845 ;
        RECT 26.735 36.240 26.905 38.675 ;
        RECT 27.445 38.165 27.775 38.335 ;
        RECT 19.640 35.605 23.640 35.775 ;
        RECT 24.270 35.275 26.905 36.240 ;
        RECT 27.305 35.955 27.475 37.995 ;
        RECT 27.745 35.955 27.915 37.995 ;
        RECT 27.445 35.615 27.775 35.785 ;
        RECT 28.315 35.275 28.485 38.675 ;
        RECT 24.270 35.265 28.485 35.275 ;
        RECT 2.550 35.245 28.485 35.265 ;
        RECT 30.550 38.665 52.440 38.835 ;
        RECT 30.550 35.265 30.720 38.665 ;
        RECT 31.350 38.155 35.350 38.325 ;
        RECT 31.120 35.945 31.290 37.985 ;
        RECT 35.410 35.945 35.580 37.985 ;
        RECT 31.350 35.605 35.350 35.775 ;
        RECT 35.980 35.265 36.150 38.665 ;
        RECT 36.780 38.155 40.780 38.325 ;
        RECT 36.550 35.945 36.720 37.985 ;
        RECT 40.840 35.945 41.010 37.985 ;
        RECT 36.780 35.605 40.780 35.775 ;
        RECT 41.410 35.265 41.580 38.665 ;
        RECT 42.210 38.155 46.210 38.325 ;
        RECT 41.980 35.945 42.150 37.985 ;
        RECT 46.270 35.945 46.440 37.985 ;
        RECT 42.210 35.605 46.210 35.775 ;
        RECT 46.840 35.265 47.010 38.665 ;
        RECT 47.640 38.155 51.640 38.325 ;
        RECT 47.410 35.945 47.580 37.985 ;
        RECT 51.700 35.945 51.870 37.985 ;
        RECT 52.270 36.240 52.440 38.665 ;
        RECT 52.710 38.670 54.460 38.840 ;
        RECT 52.710 36.270 52.880 38.670 ;
        RECT 53.420 38.160 53.750 38.330 ;
        RECT 53.280 36.950 53.450 37.990 ;
        RECT 53.720 36.950 53.890 37.990 ;
        RECT 53.420 36.610 53.750 36.780 ;
        RECT 54.290 36.270 54.460 38.670 ;
        RECT 52.710 36.240 54.460 36.270 ;
        RECT 54.735 38.675 56.485 38.845 ;
        RECT 54.735 36.240 54.905 38.675 ;
        RECT 55.445 38.165 55.775 38.335 ;
        RECT 47.640 35.605 51.640 35.775 ;
        RECT 52.270 35.275 54.905 36.240 ;
        RECT 55.305 35.955 55.475 37.995 ;
        RECT 55.745 35.955 55.915 37.995 ;
        RECT 55.445 35.615 55.775 35.785 ;
        RECT 56.315 35.275 56.485 38.675 ;
        RECT 52.270 35.265 56.485 35.275 ;
        RECT 30.550 35.245 56.485 35.265 ;
        RECT 58.550 38.665 80.440 38.835 ;
        RECT 58.550 35.265 58.720 38.665 ;
        RECT 59.350 38.155 63.350 38.325 ;
        RECT 59.120 35.945 59.290 37.985 ;
        RECT 63.410 35.945 63.580 37.985 ;
        RECT 59.350 35.605 63.350 35.775 ;
        RECT 63.980 35.265 64.150 38.665 ;
        RECT 64.780 38.155 68.780 38.325 ;
        RECT 64.550 35.945 64.720 37.985 ;
        RECT 68.840 35.945 69.010 37.985 ;
        RECT 64.780 35.605 68.780 35.775 ;
        RECT 69.410 35.265 69.580 38.665 ;
        RECT 70.210 38.155 74.210 38.325 ;
        RECT 69.980 35.945 70.150 37.985 ;
        RECT 74.270 35.945 74.440 37.985 ;
        RECT 70.210 35.605 74.210 35.775 ;
        RECT 74.840 35.265 75.010 38.665 ;
        RECT 75.640 38.155 79.640 38.325 ;
        RECT 75.410 35.945 75.580 37.985 ;
        RECT 79.700 35.945 79.870 37.985 ;
        RECT 80.270 36.240 80.440 38.665 ;
        RECT 80.710 38.670 82.460 38.840 ;
        RECT 80.710 36.270 80.880 38.670 ;
        RECT 81.420 38.160 81.750 38.330 ;
        RECT 81.280 36.950 81.450 37.990 ;
        RECT 81.720 36.950 81.890 37.990 ;
        RECT 81.420 36.610 81.750 36.780 ;
        RECT 82.290 36.270 82.460 38.670 ;
        RECT 80.710 36.240 82.460 36.270 ;
        RECT 82.735 38.675 84.485 38.845 ;
        RECT 82.735 36.240 82.905 38.675 ;
        RECT 83.445 38.165 83.775 38.335 ;
        RECT 75.640 35.605 79.640 35.775 ;
        RECT 80.270 35.275 82.905 36.240 ;
        RECT 83.305 35.955 83.475 37.995 ;
        RECT 83.745 35.955 83.915 37.995 ;
        RECT 83.445 35.615 83.775 35.785 ;
        RECT 84.315 35.275 84.485 38.675 ;
        RECT 80.270 35.265 84.485 35.275 ;
        RECT 58.550 35.245 84.485 35.265 ;
        RECT 86.550 38.665 108.440 38.835 ;
        RECT 86.550 35.265 86.720 38.665 ;
        RECT 87.350 38.155 91.350 38.325 ;
        RECT 87.120 35.945 87.290 37.985 ;
        RECT 91.410 35.945 91.580 37.985 ;
        RECT 87.350 35.605 91.350 35.775 ;
        RECT 91.980 35.265 92.150 38.665 ;
        RECT 92.780 38.155 96.780 38.325 ;
        RECT 92.550 35.945 92.720 37.985 ;
        RECT 96.840 35.945 97.010 37.985 ;
        RECT 92.780 35.605 96.780 35.775 ;
        RECT 97.410 35.265 97.580 38.665 ;
        RECT 98.210 38.155 102.210 38.325 ;
        RECT 97.980 35.945 98.150 37.985 ;
        RECT 102.270 35.945 102.440 37.985 ;
        RECT 98.210 35.605 102.210 35.775 ;
        RECT 102.840 35.265 103.010 38.665 ;
        RECT 103.640 38.155 107.640 38.325 ;
        RECT 103.410 35.945 103.580 37.985 ;
        RECT 107.700 35.945 107.870 37.985 ;
        RECT 108.270 36.240 108.440 38.665 ;
        RECT 108.710 38.670 110.460 38.840 ;
        RECT 108.710 36.270 108.880 38.670 ;
        RECT 109.420 38.160 109.750 38.330 ;
        RECT 109.280 36.950 109.450 37.990 ;
        RECT 109.720 36.950 109.890 37.990 ;
        RECT 109.420 36.610 109.750 36.780 ;
        RECT 110.290 36.270 110.460 38.670 ;
        RECT 108.710 36.240 110.460 36.270 ;
        RECT 110.735 38.675 112.485 38.845 ;
        RECT 110.735 36.240 110.905 38.675 ;
        RECT 111.445 38.165 111.775 38.335 ;
        RECT 103.640 35.605 107.640 35.775 ;
        RECT 108.270 35.275 110.905 36.240 ;
        RECT 111.305 35.955 111.475 37.995 ;
        RECT 111.745 35.955 111.915 37.995 ;
        RECT 111.445 35.615 111.775 35.785 ;
        RECT 112.315 35.275 112.485 38.675 ;
        RECT 108.270 35.265 112.485 35.275 ;
        RECT 86.550 35.245 112.485 35.265 ;
        RECT 114.550 38.665 136.440 38.835 ;
        RECT 114.550 35.265 114.720 38.665 ;
        RECT 115.350 38.155 119.350 38.325 ;
        RECT 115.120 35.945 115.290 37.985 ;
        RECT 119.410 35.945 119.580 37.985 ;
        RECT 115.350 35.605 119.350 35.775 ;
        RECT 119.980 35.265 120.150 38.665 ;
        RECT 120.780 38.155 124.780 38.325 ;
        RECT 120.550 35.945 120.720 37.985 ;
        RECT 124.840 35.945 125.010 37.985 ;
        RECT 120.780 35.605 124.780 35.775 ;
        RECT 125.410 35.265 125.580 38.665 ;
        RECT 126.210 38.155 130.210 38.325 ;
        RECT 125.980 35.945 126.150 37.985 ;
        RECT 130.270 35.945 130.440 37.985 ;
        RECT 126.210 35.605 130.210 35.775 ;
        RECT 130.840 35.265 131.010 38.665 ;
        RECT 131.640 38.155 135.640 38.325 ;
        RECT 131.410 35.945 131.580 37.985 ;
        RECT 135.700 35.945 135.870 37.985 ;
        RECT 136.270 36.240 136.440 38.665 ;
        RECT 136.710 38.670 138.460 38.840 ;
        RECT 136.710 36.270 136.880 38.670 ;
        RECT 137.420 38.160 137.750 38.330 ;
        RECT 137.280 36.950 137.450 37.990 ;
        RECT 137.720 36.950 137.890 37.990 ;
        RECT 137.420 36.610 137.750 36.780 ;
        RECT 138.290 36.270 138.460 38.670 ;
        RECT 136.710 36.240 138.460 36.270 ;
        RECT 138.735 38.675 140.485 38.845 ;
        RECT 138.735 36.240 138.905 38.675 ;
        RECT 139.445 38.165 139.775 38.335 ;
        RECT 131.640 35.605 135.640 35.775 ;
        RECT 136.270 35.275 138.905 36.240 ;
        RECT 139.305 35.955 139.475 37.995 ;
        RECT 139.745 35.955 139.915 37.995 ;
        RECT 139.445 35.615 139.775 35.785 ;
        RECT 140.315 35.275 140.485 38.675 ;
        RECT 136.270 35.265 140.485 35.275 ;
        RECT 114.550 35.245 140.485 35.265 ;
        RECT 1.895 35.105 28.485 35.245 ;
        RECT 29.895 35.105 56.485 35.245 ;
        RECT 57.895 35.105 84.485 35.245 ;
        RECT 85.895 35.105 112.485 35.245 ;
        RECT 113.895 35.105 140.485 35.245 ;
        RECT 1.895 34.380 28.475 35.105 ;
        RECT 29.895 34.380 56.475 35.105 ;
        RECT 57.895 34.380 84.475 35.105 ;
        RECT 85.895 34.380 112.475 35.105 ;
        RECT 113.895 34.380 140.475 35.105 ;
        RECT 1.870 33.480 28.345 33.960 ;
        RECT 29.870 33.480 56.345 33.960 ;
        RECT 57.870 33.480 84.345 33.960 ;
        RECT 85.870 33.480 112.345 33.960 ;
        RECT 113.870 33.480 140.345 33.960 ;
        RECT 1.855 33.420 28.345 33.480 ;
        RECT 29.855 33.420 56.345 33.480 ;
        RECT 57.855 33.420 84.345 33.480 ;
        RECT 85.855 33.420 112.345 33.480 ;
        RECT 113.855 33.420 140.345 33.480 ;
        RECT 1.855 33.260 28.400 33.420 ;
        RECT 1.855 33.235 14.600 33.260 ;
        RECT 1.855 33.005 6.180 33.235 ;
        RECT 1.890 23.745 2.060 33.005 ;
        RECT 2.785 32.435 4.825 32.605 ;
        RECT 2.400 24.375 2.570 32.375 ;
        RECT 5.040 24.375 5.210 32.375 ;
        RECT 2.785 24.145 4.825 24.315 ;
        RECT 5.550 23.745 5.720 33.005 ;
        RECT 1.890 23.575 5.720 23.745 ;
        RECT 6.010 23.745 6.180 33.005 ;
        RECT 6.810 32.725 8.810 32.895 ;
        RECT 6.580 24.470 6.750 32.510 ;
        RECT 8.870 24.470 9.040 32.510 ;
        RECT 6.810 24.085 8.810 24.255 ;
        RECT 9.440 23.745 9.610 33.235 ;
        RECT 10.240 32.725 12.240 32.895 ;
        RECT 10.010 24.470 10.180 32.510 ;
        RECT 12.300 24.470 12.470 32.510 ;
        RECT 12.870 31.665 14.600 33.235 ;
        RECT 26.650 33.250 28.400 33.260 ;
        RECT 12.870 31.495 21.335 31.665 ;
        RECT 12.870 30.085 14.675 31.495 ;
        RECT 15.015 30.625 15.185 30.955 ;
        RECT 15.400 30.925 20.440 31.095 ;
        RECT 15.400 30.485 20.440 30.655 ;
        RECT 20.655 30.625 20.825 30.955 ;
        RECT 21.165 30.085 21.335 31.495 ;
        RECT 12.870 29.915 21.335 30.085 ;
        RECT 12.870 29.400 14.600 29.915 ;
        RECT 12.870 29.285 24.350 29.400 ;
        RECT 10.240 24.085 12.240 24.255 ;
        RECT 12.870 23.745 13.040 29.285 ;
        RECT 6.010 23.575 13.040 23.745 ;
        RECT 13.320 29.230 24.350 29.285 ;
        RECT 13.320 23.740 13.490 29.230 ;
        RECT 14.120 28.720 18.120 28.890 ;
        RECT 13.890 24.465 14.060 28.505 ;
        RECT 18.180 24.465 18.350 28.505 ;
        RECT 14.120 24.080 18.120 24.250 ;
        RECT 18.750 23.740 18.920 29.230 ;
        RECT 19.550 28.720 23.550 28.890 ;
        RECT 19.320 24.465 19.490 28.505 ;
        RECT 23.610 24.465 23.780 28.505 ;
        RECT 19.550 24.080 23.550 24.250 ;
        RECT 24.180 23.740 24.350 29.230 ;
        RECT 13.320 23.570 24.350 23.740 ;
        RECT 24.625 29.245 26.375 29.415 ;
        RECT 24.625 23.755 24.795 29.245 ;
        RECT 25.335 28.735 25.665 28.905 ;
        RECT 25.195 24.480 25.365 28.520 ;
        RECT 25.635 24.480 25.805 28.520 ;
        RECT 25.335 24.095 25.665 24.265 ;
        RECT 26.205 23.755 26.375 29.245 ;
        RECT 24.625 23.585 26.375 23.755 ;
        RECT 26.650 23.760 26.820 33.250 ;
        RECT 27.360 32.740 27.690 32.910 ;
        RECT 27.220 24.485 27.390 32.525 ;
        RECT 27.660 24.485 27.830 32.525 ;
        RECT 27.360 24.100 27.690 24.270 ;
        RECT 28.230 23.760 28.400 33.250 ;
        RECT 29.855 33.260 56.400 33.420 ;
        RECT 29.855 33.235 42.600 33.260 ;
        RECT 29.855 33.005 34.180 33.235 ;
        RECT 26.650 23.590 28.400 23.760 ;
        RECT 29.890 23.745 30.060 33.005 ;
        RECT 30.785 32.435 32.825 32.605 ;
        RECT 30.400 24.375 30.570 32.375 ;
        RECT 33.040 24.375 33.210 32.375 ;
        RECT 30.785 24.145 32.825 24.315 ;
        RECT 33.550 23.745 33.720 33.005 ;
        RECT 29.890 23.575 33.720 23.745 ;
        RECT 34.010 23.745 34.180 33.005 ;
        RECT 34.810 32.725 36.810 32.895 ;
        RECT 34.580 24.470 34.750 32.510 ;
        RECT 36.870 24.470 37.040 32.510 ;
        RECT 34.810 24.085 36.810 24.255 ;
        RECT 37.440 23.745 37.610 33.235 ;
        RECT 38.240 32.725 40.240 32.895 ;
        RECT 38.010 24.470 38.180 32.510 ;
        RECT 40.300 24.470 40.470 32.510 ;
        RECT 40.870 31.665 42.600 33.235 ;
        RECT 54.650 33.250 56.400 33.260 ;
        RECT 40.870 31.495 49.335 31.665 ;
        RECT 40.870 30.085 42.675 31.495 ;
        RECT 43.015 30.625 43.185 30.955 ;
        RECT 43.400 30.925 48.440 31.095 ;
        RECT 43.400 30.485 48.440 30.655 ;
        RECT 48.655 30.625 48.825 30.955 ;
        RECT 49.165 30.085 49.335 31.495 ;
        RECT 40.870 29.915 49.335 30.085 ;
        RECT 40.870 29.400 42.600 29.915 ;
        RECT 40.870 29.285 52.350 29.400 ;
        RECT 38.240 24.085 40.240 24.255 ;
        RECT 40.870 23.745 41.040 29.285 ;
        RECT 34.010 23.575 41.040 23.745 ;
        RECT 41.320 29.230 52.350 29.285 ;
        RECT 41.320 23.740 41.490 29.230 ;
        RECT 42.120 28.720 46.120 28.890 ;
        RECT 41.890 24.465 42.060 28.505 ;
        RECT 46.180 24.465 46.350 28.505 ;
        RECT 42.120 24.080 46.120 24.250 ;
        RECT 46.750 23.740 46.920 29.230 ;
        RECT 47.550 28.720 51.550 28.890 ;
        RECT 47.320 24.465 47.490 28.505 ;
        RECT 51.610 24.465 51.780 28.505 ;
        RECT 47.550 24.080 51.550 24.250 ;
        RECT 52.180 23.740 52.350 29.230 ;
        RECT 41.320 23.570 52.350 23.740 ;
        RECT 52.625 29.245 54.375 29.415 ;
        RECT 52.625 23.755 52.795 29.245 ;
        RECT 53.335 28.735 53.665 28.905 ;
        RECT 53.195 24.480 53.365 28.520 ;
        RECT 53.635 24.480 53.805 28.520 ;
        RECT 53.335 24.095 53.665 24.265 ;
        RECT 54.205 23.755 54.375 29.245 ;
        RECT 52.625 23.585 54.375 23.755 ;
        RECT 54.650 23.760 54.820 33.250 ;
        RECT 55.360 32.740 55.690 32.910 ;
        RECT 55.220 24.485 55.390 32.525 ;
        RECT 55.660 24.485 55.830 32.525 ;
        RECT 55.360 24.100 55.690 24.270 ;
        RECT 56.230 23.760 56.400 33.250 ;
        RECT 57.855 33.260 84.400 33.420 ;
        RECT 57.855 33.235 70.600 33.260 ;
        RECT 57.855 33.005 62.180 33.235 ;
        RECT 54.650 23.590 56.400 23.760 ;
        RECT 57.890 23.745 58.060 33.005 ;
        RECT 58.785 32.435 60.825 32.605 ;
        RECT 58.400 24.375 58.570 32.375 ;
        RECT 61.040 24.375 61.210 32.375 ;
        RECT 58.785 24.145 60.825 24.315 ;
        RECT 61.550 23.745 61.720 33.005 ;
        RECT 57.890 23.575 61.720 23.745 ;
        RECT 62.010 23.745 62.180 33.005 ;
        RECT 62.810 32.725 64.810 32.895 ;
        RECT 62.580 24.470 62.750 32.510 ;
        RECT 64.870 24.470 65.040 32.510 ;
        RECT 62.810 24.085 64.810 24.255 ;
        RECT 65.440 23.745 65.610 33.235 ;
        RECT 66.240 32.725 68.240 32.895 ;
        RECT 66.010 24.470 66.180 32.510 ;
        RECT 68.300 24.470 68.470 32.510 ;
        RECT 68.870 31.665 70.600 33.235 ;
        RECT 82.650 33.250 84.400 33.260 ;
        RECT 68.870 31.495 77.335 31.665 ;
        RECT 68.870 30.085 70.675 31.495 ;
        RECT 71.015 30.625 71.185 30.955 ;
        RECT 71.400 30.925 76.440 31.095 ;
        RECT 71.400 30.485 76.440 30.655 ;
        RECT 76.655 30.625 76.825 30.955 ;
        RECT 77.165 30.085 77.335 31.495 ;
        RECT 68.870 29.915 77.335 30.085 ;
        RECT 68.870 29.400 70.600 29.915 ;
        RECT 68.870 29.285 80.350 29.400 ;
        RECT 66.240 24.085 68.240 24.255 ;
        RECT 68.870 23.745 69.040 29.285 ;
        RECT 62.010 23.575 69.040 23.745 ;
        RECT 69.320 29.230 80.350 29.285 ;
        RECT 69.320 23.740 69.490 29.230 ;
        RECT 70.120 28.720 74.120 28.890 ;
        RECT 69.890 24.465 70.060 28.505 ;
        RECT 74.180 24.465 74.350 28.505 ;
        RECT 70.120 24.080 74.120 24.250 ;
        RECT 74.750 23.740 74.920 29.230 ;
        RECT 75.550 28.720 79.550 28.890 ;
        RECT 75.320 24.465 75.490 28.505 ;
        RECT 79.610 24.465 79.780 28.505 ;
        RECT 75.550 24.080 79.550 24.250 ;
        RECT 80.180 23.740 80.350 29.230 ;
        RECT 69.320 23.570 80.350 23.740 ;
        RECT 80.625 29.245 82.375 29.415 ;
        RECT 80.625 23.755 80.795 29.245 ;
        RECT 81.335 28.735 81.665 28.905 ;
        RECT 81.195 24.480 81.365 28.520 ;
        RECT 81.635 24.480 81.805 28.520 ;
        RECT 81.335 24.095 81.665 24.265 ;
        RECT 82.205 23.755 82.375 29.245 ;
        RECT 80.625 23.585 82.375 23.755 ;
        RECT 82.650 23.760 82.820 33.250 ;
        RECT 83.360 32.740 83.690 32.910 ;
        RECT 83.220 24.485 83.390 32.525 ;
        RECT 83.660 24.485 83.830 32.525 ;
        RECT 83.360 24.100 83.690 24.270 ;
        RECT 84.230 23.760 84.400 33.250 ;
        RECT 85.855 33.260 112.400 33.420 ;
        RECT 85.855 33.235 98.600 33.260 ;
        RECT 85.855 33.005 90.180 33.235 ;
        RECT 82.650 23.590 84.400 23.760 ;
        RECT 85.890 23.745 86.060 33.005 ;
        RECT 86.785 32.435 88.825 32.605 ;
        RECT 86.400 24.375 86.570 32.375 ;
        RECT 89.040 24.375 89.210 32.375 ;
        RECT 86.785 24.145 88.825 24.315 ;
        RECT 89.550 23.745 89.720 33.005 ;
        RECT 85.890 23.575 89.720 23.745 ;
        RECT 90.010 23.745 90.180 33.005 ;
        RECT 90.810 32.725 92.810 32.895 ;
        RECT 90.580 24.470 90.750 32.510 ;
        RECT 92.870 24.470 93.040 32.510 ;
        RECT 90.810 24.085 92.810 24.255 ;
        RECT 93.440 23.745 93.610 33.235 ;
        RECT 94.240 32.725 96.240 32.895 ;
        RECT 94.010 24.470 94.180 32.510 ;
        RECT 96.300 24.470 96.470 32.510 ;
        RECT 96.870 31.665 98.600 33.235 ;
        RECT 110.650 33.250 112.400 33.260 ;
        RECT 96.870 31.495 105.335 31.665 ;
        RECT 96.870 30.085 98.675 31.495 ;
        RECT 99.015 30.625 99.185 30.955 ;
        RECT 99.400 30.925 104.440 31.095 ;
        RECT 99.400 30.485 104.440 30.655 ;
        RECT 104.655 30.625 104.825 30.955 ;
        RECT 105.165 30.085 105.335 31.495 ;
        RECT 96.870 29.915 105.335 30.085 ;
        RECT 96.870 29.400 98.600 29.915 ;
        RECT 96.870 29.285 108.350 29.400 ;
        RECT 94.240 24.085 96.240 24.255 ;
        RECT 96.870 23.745 97.040 29.285 ;
        RECT 90.010 23.575 97.040 23.745 ;
        RECT 97.320 29.230 108.350 29.285 ;
        RECT 97.320 23.740 97.490 29.230 ;
        RECT 98.120 28.720 102.120 28.890 ;
        RECT 97.890 24.465 98.060 28.505 ;
        RECT 102.180 24.465 102.350 28.505 ;
        RECT 98.120 24.080 102.120 24.250 ;
        RECT 102.750 23.740 102.920 29.230 ;
        RECT 103.550 28.720 107.550 28.890 ;
        RECT 103.320 24.465 103.490 28.505 ;
        RECT 107.610 24.465 107.780 28.505 ;
        RECT 103.550 24.080 107.550 24.250 ;
        RECT 108.180 23.740 108.350 29.230 ;
        RECT 97.320 23.570 108.350 23.740 ;
        RECT 108.625 29.245 110.375 29.415 ;
        RECT 108.625 23.755 108.795 29.245 ;
        RECT 109.335 28.735 109.665 28.905 ;
        RECT 109.195 24.480 109.365 28.520 ;
        RECT 109.635 24.480 109.805 28.520 ;
        RECT 109.335 24.095 109.665 24.265 ;
        RECT 110.205 23.755 110.375 29.245 ;
        RECT 108.625 23.585 110.375 23.755 ;
        RECT 110.650 23.760 110.820 33.250 ;
        RECT 111.360 32.740 111.690 32.910 ;
        RECT 111.220 24.485 111.390 32.525 ;
        RECT 111.660 24.485 111.830 32.525 ;
        RECT 111.360 24.100 111.690 24.270 ;
        RECT 112.230 23.760 112.400 33.250 ;
        RECT 113.855 33.260 140.400 33.420 ;
        RECT 113.855 33.235 126.600 33.260 ;
        RECT 113.855 33.005 118.180 33.235 ;
        RECT 110.650 23.590 112.400 23.760 ;
        RECT 113.890 23.745 114.060 33.005 ;
        RECT 114.785 32.435 116.825 32.605 ;
        RECT 114.400 24.375 114.570 32.375 ;
        RECT 117.040 24.375 117.210 32.375 ;
        RECT 114.785 24.145 116.825 24.315 ;
        RECT 117.550 23.745 117.720 33.005 ;
        RECT 113.890 23.575 117.720 23.745 ;
        RECT 118.010 23.745 118.180 33.005 ;
        RECT 118.810 32.725 120.810 32.895 ;
        RECT 118.580 24.470 118.750 32.510 ;
        RECT 120.870 24.470 121.040 32.510 ;
        RECT 118.810 24.085 120.810 24.255 ;
        RECT 121.440 23.745 121.610 33.235 ;
        RECT 122.240 32.725 124.240 32.895 ;
        RECT 122.010 24.470 122.180 32.510 ;
        RECT 124.300 24.470 124.470 32.510 ;
        RECT 124.870 31.665 126.600 33.235 ;
        RECT 138.650 33.250 140.400 33.260 ;
        RECT 124.870 31.495 133.335 31.665 ;
        RECT 124.870 30.085 126.675 31.495 ;
        RECT 127.015 30.625 127.185 30.955 ;
        RECT 127.400 30.925 132.440 31.095 ;
        RECT 127.400 30.485 132.440 30.655 ;
        RECT 132.655 30.625 132.825 30.955 ;
        RECT 133.165 30.085 133.335 31.495 ;
        RECT 124.870 29.915 133.335 30.085 ;
        RECT 124.870 29.400 126.600 29.915 ;
        RECT 124.870 29.285 136.350 29.400 ;
        RECT 122.240 24.085 124.240 24.255 ;
        RECT 124.870 23.745 125.040 29.285 ;
        RECT 118.010 23.575 125.040 23.745 ;
        RECT 125.320 29.230 136.350 29.285 ;
        RECT 125.320 23.740 125.490 29.230 ;
        RECT 126.120 28.720 130.120 28.890 ;
        RECT 125.890 24.465 126.060 28.505 ;
        RECT 130.180 24.465 130.350 28.505 ;
        RECT 126.120 24.080 130.120 24.250 ;
        RECT 130.750 23.740 130.920 29.230 ;
        RECT 131.550 28.720 135.550 28.890 ;
        RECT 131.320 24.465 131.490 28.505 ;
        RECT 135.610 24.465 135.780 28.505 ;
        RECT 131.550 24.080 135.550 24.250 ;
        RECT 136.180 23.740 136.350 29.230 ;
        RECT 125.320 23.570 136.350 23.740 ;
        RECT 136.625 29.245 138.375 29.415 ;
        RECT 136.625 23.755 136.795 29.245 ;
        RECT 137.335 28.735 137.665 28.905 ;
        RECT 137.195 24.480 137.365 28.520 ;
        RECT 137.635 24.480 137.805 28.520 ;
        RECT 137.335 24.095 137.665 24.265 ;
        RECT 138.205 23.755 138.375 29.245 ;
        RECT 136.625 23.585 138.375 23.755 ;
        RECT 138.650 23.760 138.820 33.250 ;
        RECT 139.360 32.740 139.690 32.910 ;
        RECT 139.220 24.485 139.390 32.525 ;
        RECT 139.660 24.485 139.830 32.525 ;
        RECT 139.360 24.100 139.690 24.270 ;
        RECT 140.230 23.760 140.400 33.250 ;
        RECT 138.650 23.590 140.400 23.760 ;
        RECT 2.550 22.665 24.440 22.835 ;
        RECT 2.550 19.265 2.720 22.665 ;
        RECT 3.350 22.155 7.350 22.325 ;
        RECT 3.120 19.945 3.290 21.985 ;
        RECT 7.410 19.945 7.580 21.985 ;
        RECT 3.350 19.605 7.350 19.775 ;
        RECT 7.980 19.265 8.150 22.665 ;
        RECT 8.780 22.155 12.780 22.325 ;
        RECT 8.550 19.945 8.720 21.985 ;
        RECT 12.840 19.945 13.010 21.985 ;
        RECT 8.780 19.605 12.780 19.775 ;
        RECT 13.410 19.265 13.580 22.665 ;
        RECT 14.210 22.155 18.210 22.325 ;
        RECT 13.980 19.945 14.150 21.985 ;
        RECT 18.270 19.945 18.440 21.985 ;
        RECT 14.210 19.605 18.210 19.775 ;
        RECT 18.840 19.265 19.010 22.665 ;
        RECT 19.640 22.155 23.640 22.325 ;
        RECT 19.410 19.945 19.580 21.985 ;
        RECT 23.700 19.945 23.870 21.985 ;
        RECT 24.270 20.240 24.440 22.665 ;
        RECT 24.710 22.670 26.460 22.840 ;
        RECT 24.710 20.270 24.880 22.670 ;
        RECT 25.420 22.160 25.750 22.330 ;
        RECT 25.280 20.950 25.450 21.990 ;
        RECT 25.720 20.950 25.890 21.990 ;
        RECT 25.420 20.610 25.750 20.780 ;
        RECT 26.290 20.270 26.460 22.670 ;
        RECT 24.710 20.240 26.460 20.270 ;
        RECT 26.735 22.675 28.485 22.845 ;
        RECT 26.735 20.240 26.905 22.675 ;
        RECT 27.445 22.165 27.775 22.335 ;
        RECT 19.640 19.605 23.640 19.775 ;
        RECT 24.270 19.275 26.905 20.240 ;
        RECT 27.305 19.955 27.475 21.995 ;
        RECT 27.745 19.955 27.915 21.995 ;
        RECT 27.445 19.615 27.775 19.785 ;
        RECT 28.315 19.275 28.485 22.675 ;
        RECT 24.270 19.265 28.485 19.275 ;
        RECT 2.550 19.245 28.485 19.265 ;
        RECT 30.550 22.665 52.440 22.835 ;
        RECT 30.550 19.265 30.720 22.665 ;
        RECT 31.350 22.155 35.350 22.325 ;
        RECT 31.120 19.945 31.290 21.985 ;
        RECT 35.410 19.945 35.580 21.985 ;
        RECT 31.350 19.605 35.350 19.775 ;
        RECT 35.980 19.265 36.150 22.665 ;
        RECT 36.780 22.155 40.780 22.325 ;
        RECT 36.550 19.945 36.720 21.985 ;
        RECT 40.840 19.945 41.010 21.985 ;
        RECT 36.780 19.605 40.780 19.775 ;
        RECT 41.410 19.265 41.580 22.665 ;
        RECT 42.210 22.155 46.210 22.325 ;
        RECT 41.980 19.945 42.150 21.985 ;
        RECT 46.270 19.945 46.440 21.985 ;
        RECT 42.210 19.605 46.210 19.775 ;
        RECT 46.840 19.265 47.010 22.665 ;
        RECT 47.640 22.155 51.640 22.325 ;
        RECT 47.410 19.945 47.580 21.985 ;
        RECT 51.700 19.945 51.870 21.985 ;
        RECT 52.270 20.240 52.440 22.665 ;
        RECT 52.710 22.670 54.460 22.840 ;
        RECT 52.710 20.270 52.880 22.670 ;
        RECT 53.420 22.160 53.750 22.330 ;
        RECT 53.280 20.950 53.450 21.990 ;
        RECT 53.720 20.950 53.890 21.990 ;
        RECT 53.420 20.610 53.750 20.780 ;
        RECT 54.290 20.270 54.460 22.670 ;
        RECT 52.710 20.240 54.460 20.270 ;
        RECT 54.735 22.675 56.485 22.845 ;
        RECT 54.735 20.240 54.905 22.675 ;
        RECT 55.445 22.165 55.775 22.335 ;
        RECT 47.640 19.605 51.640 19.775 ;
        RECT 52.270 19.275 54.905 20.240 ;
        RECT 55.305 19.955 55.475 21.995 ;
        RECT 55.745 19.955 55.915 21.995 ;
        RECT 55.445 19.615 55.775 19.785 ;
        RECT 56.315 19.275 56.485 22.675 ;
        RECT 52.270 19.265 56.485 19.275 ;
        RECT 30.550 19.245 56.485 19.265 ;
        RECT 58.550 22.665 80.440 22.835 ;
        RECT 58.550 19.265 58.720 22.665 ;
        RECT 59.350 22.155 63.350 22.325 ;
        RECT 59.120 19.945 59.290 21.985 ;
        RECT 63.410 19.945 63.580 21.985 ;
        RECT 59.350 19.605 63.350 19.775 ;
        RECT 63.980 19.265 64.150 22.665 ;
        RECT 64.780 22.155 68.780 22.325 ;
        RECT 64.550 19.945 64.720 21.985 ;
        RECT 68.840 19.945 69.010 21.985 ;
        RECT 64.780 19.605 68.780 19.775 ;
        RECT 69.410 19.265 69.580 22.665 ;
        RECT 70.210 22.155 74.210 22.325 ;
        RECT 69.980 19.945 70.150 21.985 ;
        RECT 74.270 19.945 74.440 21.985 ;
        RECT 70.210 19.605 74.210 19.775 ;
        RECT 74.840 19.265 75.010 22.665 ;
        RECT 75.640 22.155 79.640 22.325 ;
        RECT 75.410 19.945 75.580 21.985 ;
        RECT 79.700 19.945 79.870 21.985 ;
        RECT 80.270 20.240 80.440 22.665 ;
        RECT 80.710 22.670 82.460 22.840 ;
        RECT 80.710 20.270 80.880 22.670 ;
        RECT 81.420 22.160 81.750 22.330 ;
        RECT 81.280 20.950 81.450 21.990 ;
        RECT 81.720 20.950 81.890 21.990 ;
        RECT 81.420 20.610 81.750 20.780 ;
        RECT 82.290 20.270 82.460 22.670 ;
        RECT 80.710 20.240 82.460 20.270 ;
        RECT 82.735 22.675 84.485 22.845 ;
        RECT 82.735 20.240 82.905 22.675 ;
        RECT 83.445 22.165 83.775 22.335 ;
        RECT 75.640 19.605 79.640 19.775 ;
        RECT 80.270 19.275 82.905 20.240 ;
        RECT 83.305 19.955 83.475 21.995 ;
        RECT 83.745 19.955 83.915 21.995 ;
        RECT 83.445 19.615 83.775 19.785 ;
        RECT 84.315 19.275 84.485 22.675 ;
        RECT 80.270 19.265 84.485 19.275 ;
        RECT 58.550 19.245 84.485 19.265 ;
        RECT 86.550 22.665 108.440 22.835 ;
        RECT 86.550 19.265 86.720 22.665 ;
        RECT 87.350 22.155 91.350 22.325 ;
        RECT 87.120 19.945 87.290 21.985 ;
        RECT 91.410 19.945 91.580 21.985 ;
        RECT 87.350 19.605 91.350 19.775 ;
        RECT 91.980 19.265 92.150 22.665 ;
        RECT 92.780 22.155 96.780 22.325 ;
        RECT 92.550 19.945 92.720 21.985 ;
        RECT 96.840 19.945 97.010 21.985 ;
        RECT 92.780 19.605 96.780 19.775 ;
        RECT 97.410 19.265 97.580 22.665 ;
        RECT 98.210 22.155 102.210 22.325 ;
        RECT 97.980 19.945 98.150 21.985 ;
        RECT 102.270 19.945 102.440 21.985 ;
        RECT 98.210 19.605 102.210 19.775 ;
        RECT 102.840 19.265 103.010 22.665 ;
        RECT 103.640 22.155 107.640 22.325 ;
        RECT 103.410 19.945 103.580 21.985 ;
        RECT 107.700 19.945 107.870 21.985 ;
        RECT 108.270 20.240 108.440 22.665 ;
        RECT 108.710 22.670 110.460 22.840 ;
        RECT 108.710 20.270 108.880 22.670 ;
        RECT 109.420 22.160 109.750 22.330 ;
        RECT 109.280 20.950 109.450 21.990 ;
        RECT 109.720 20.950 109.890 21.990 ;
        RECT 109.420 20.610 109.750 20.780 ;
        RECT 110.290 20.270 110.460 22.670 ;
        RECT 108.710 20.240 110.460 20.270 ;
        RECT 110.735 22.675 112.485 22.845 ;
        RECT 110.735 20.240 110.905 22.675 ;
        RECT 111.445 22.165 111.775 22.335 ;
        RECT 103.640 19.605 107.640 19.775 ;
        RECT 108.270 19.275 110.905 20.240 ;
        RECT 111.305 19.955 111.475 21.995 ;
        RECT 111.745 19.955 111.915 21.995 ;
        RECT 111.445 19.615 111.775 19.785 ;
        RECT 112.315 19.275 112.485 22.675 ;
        RECT 108.270 19.265 112.485 19.275 ;
        RECT 86.550 19.245 112.485 19.265 ;
        RECT 114.550 22.665 136.440 22.835 ;
        RECT 114.550 19.265 114.720 22.665 ;
        RECT 115.350 22.155 119.350 22.325 ;
        RECT 115.120 19.945 115.290 21.985 ;
        RECT 119.410 19.945 119.580 21.985 ;
        RECT 115.350 19.605 119.350 19.775 ;
        RECT 119.980 19.265 120.150 22.665 ;
        RECT 120.780 22.155 124.780 22.325 ;
        RECT 120.550 19.945 120.720 21.985 ;
        RECT 124.840 19.945 125.010 21.985 ;
        RECT 120.780 19.605 124.780 19.775 ;
        RECT 125.410 19.265 125.580 22.665 ;
        RECT 126.210 22.155 130.210 22.325 ;
        RECT 125.980 19.945 126.150 21.985 ;
        RECT 130.270 19.945 130.440 21.985 ;
        RECT 126.210 19.605 130.210 19.775 ;
        RECT 130.840 19.265 131.010 22.665 ;
        RECT 131.640 22.155 135.640 22.325 ;
        RECT 131.410 19.945 131.580 21.985 ;
        RECT 135.700 19.945 135.870 21.985 ;
        RECT 136.270 20.240 136.440 22.665 ;
        RECT 136.710 22.670 138.460 22.840 ;
        RECT 136.710 20.270 136.880 22.670 ;
        RECT 137.420 22.160 137.750 22.330 ;
        RECT 137.280 20.950 137.450 21.990 ;
        RECT 137.720 20.950 137.890 21.990 ;
        RECT 137.420 20.610 137.750 20.780 ;
        RECT 138.290 20.270 138.460 22.670 ;
        RECT 136.710 20.240 138.460 20.270 ;
        RECT 138.735 22.675 140.485 22.845 ;
        RECT 138.735 20.240 138.905 22.675 ;
        RECT 139.445 22.165 139.775 22.335 ;
        RECT 131.640 19.605 135.640 19.775 ;
        RECT 136.270 19.275 138.905 20.240 ;
        RECT 139.305 19.955 139.475 21.995 ;
        RECT 139.745 19.955 139.915 21.995 ;
        RECT 139.445 19.615 139.775 19.785 ;
        RECT 140.315 19.275 140.485 22.675 ;
        RECT 136.270 19.265 140.485 19.275 ;
        RECT 114.550 19.245 140.485 19.265 ;
        RECT 1.895 19.105 28.485 19.245 ;
        RECT 29.895 19.105 56.485 19.245 ;
        RECT 57.895 19.105 84.485 19.245 ;
        RECT 85.895 19.105 112.485 19.245 ;
        RECT 113.895 19.105 140.485 19.245 ;
        RECT 1.895 18.380 28.475 19.105 ;
        RECT 29.895 18.380 56.475 19.105 ;
        RECT 57.895 18.380 84.475 19.105 ;
        RECT 85.895 18.380 112.475 19.105 ;
        RECT 113.895 18.380 140.475 19.105 ;
        RECT 1.870 17.480 28.345 17.960 ;
        RECT 29.870 17.480 56.345 17.960 ;
        RECT 57.870 17.480 84.345 17.960 ;
        RECT 85.870 17.480 112.345 17.960 ;
        RECT 113.870 17.480 140.345 17.960 ;
        RECT 1.855 17.420 28.345 17.480 ;
        RECT 29.855 17.420 56.345 17.480 ;
        RECT 57.855 17.420 84.345 17.480 ;
        RECT 85.855 17.420 112.345 17.480 ;
        RECT 113.855 17.420 140.345 17.480 ;
        RECT 1.855 17.260 28.400 17.420 ;
        RECT 1.855 17.235 14.600 17.260 ;
        RECT 1.855 17.005 6.180 17.235 ;
        RECT 1.890 7.745 2.060 17.005 ;
        RECT 2.785 16.435 4.825 16.605 ;
        RECT 2.400 8.375 2.570 16.375 ;
        RECT 5.040 8.375 5.210 16.375 ;
        RECT 2.785 8.145 4.825 8.315 ;
        RECT 5.550 7.745 5.720 17.005 ;
        RECT 1.890 7.575 5.720 7.745 ;
        RECT 6.010 7.745 6.180 17.005 ;
        RECT 6.810 16.725 8.810 16.895 ;
        RECT 6.580 8.470 6.750 16.510 ;
        RECT 8.870 8.470 9.040 16.510 ;
        RECT 6.810 8.085 8.810 8.255 ;
        RECT 9.440 7.745 9.610 17.235 ;
        RECT 10.240 16.725 12.240 16.895 ;
        RECT 10.010 8.470 10.180 16.510 ;
        RECT 12.300 8.470 12.470 16.510 ;
        RECT 12.870 15.665 14.600 17.235 ;
        RECT 26.650 17.250 28.400 17.260 ;
        RECT 12.870 15.495 21.335 15.665 ;
        RECT 12.870 14.085 14.675 15.495 ;
        RECT 15.015 14.625 15.185 14.955 ;
        RECT 15.400 14.925 20.440 15.095 ;
        RECT 15.400 14.485 20.440 14.655 ;
        RECT 20.655 14.625 20.825 14.955 ;
        RECT 21.165 14.085 21.335 15.495 ;
        RECT 12.870 13.915 21.335 14.085 ;
        RECT 12.870 13.400 14.600 13.915 ;
        RECT 12.870 13.285 24.350 13.400 ;
        RECT 10.240 8.085 12.240 8.255 ;
        RECT 12.870 7.745 13.040 13.285 ;
        RECT 6.010 7.575 13.040 7.745 ;
        RECT 13.320 13.230 24.350 13.285 ;
        RECT 13.320 7.740 13.490 13.230 ;
        RECT 14.120 12.720 18.120 12.890 ;
        RECT 13.890 8.465 14.060 12.505 ;
        RECT 18.180 8.465 18.350 12.505 ;
        RECT 14.120 8.080 18.120 8.250 ;
        RECT 18.750 7.740 18.920 13.230 ;
        RECT 19.550 12.720 23.550 12.890 ;
        RECT 19.320 8.465 19.490 12.505 ;
        RECT 23.610 8.465 23.780 12.505 ;
        RECT 19.550 8.080 23.550 8.250 ;
        RECT 24.180 7.740 24.350 13.230 ;
        RECT 13.320 7.570 24.350 7.740 ;
        RECT 24.625 13.245 26.375 13.415 ;
        RECT 24.625 7.755 24.795 13.245 ;
        RECT 25.335 12.735 25.665 12.905 ;
        RECT 25.195 8.480 25.365 12.520 ;
        RECT 25.635 8.480 25.805 12.520 ;
        RECT 25.335 8.095 25.665 8.265 ;
        RECT 26.205 7.755 26.375 13.245 ;
        RECT 24.625 7.585 26.375 7.755 ;
        RECT 26.650 7.760 26.820 17.250 ;
        RECT 27.360 16.740 27.690 16.910 ;
        RECT 27.220 8.485 27.390 16.525 ;
        RECT 27.660 8.485 27.830 16.525 ;
        RECT 27.360 8.100 27.690 8.270 ;
        RECT 28.230 7.760 28.400 17.250 ;
        RECT 29.855 17.260 56.400 17.420 ;
        RECT 29.855 17.235 42.600 17.260 ;
        RECT 29.855 17.005 34.180 17.235 ;
        RECT 26.650 7.590 28.400 7.760 ;
        RECT 29.890 7.745 30.060 17.005 ;
        RECT 30.785 16.435 32.825 16.605 ;
        RECT 30.400 8.375 30.570 16.375 ;
        RECT 33.040 8.375 33.210 16.375 ;
        RECT 30.785 8.145 32.825 8.315 ;
        RECT 33.550 7.745 33.720 17.005 ;
        RECT 29.890 7.575 33.720 7.745 ;
        RECT 34.010 7.745 34.180 17.005 ;
        RECT 34.810 16.725 36.810 16.895 ;
        RECT 34.580 8.470 34.750 16.510 ;
        RECT 36.870 8.470 37.040 16.510 ;
        RECT 34.810 8.085 36.810 8.255 ;
        RECT 37.440 7.745 37.610 17.235 ;
        RECT 38.240 16.725 40.240 16.895 ;
        RECT 38.010 8.470 38.180 16.510 ;
        RECT 40.300 8.470 40.470 16.510 ;
        RECT 40.870 15.665 42.600 17.235 ;
        RECT 54.650 17.250 56.400 17.260 ;
        RECT 40.870 15.495 49.335 15.665 ;
        RECT 40.870 14.085 42.675 15.495 ;
        RECT 43.015 14.625 43.185 14.955 ;
        RECT 43.400 14.925 48.440 15.095 ;
        RECT 43.400 14.485 48.440 14.655 ;
        RECT 48.655 14.625 48.825 14.955 ;
        RECT 49.165 14.085 49.335 15.495 ;
        RECT 40.870 13.915 49.335 14.085 ;
        RECT 40.870 13.400 42.600 13.915 ;
        RECT 40.870 13.285 52.350 13.400 ;
        RECT 38.240 8.085 40.240 8.255 ;
        RECT 40.870 7.745 41.040 13.285 ;
        RECT 34.010 7.575 41.040 7.745 ;
        RECT 41.320 13.230 52.350 13.285 ;
        RECT 41.320 7.740 41.490 13.230 ;
        RECT 42.120 12.720 46.120 12.890 ;
        RECT 41.890 8.465 42.060 12.505 ;
        RECT 46.180 8.465 46.350 12.505 ;
        RECT 42.120 8.080 46.120 8.250 ;
        RECT 46.750 7.740 46.920 13.230 ;
        RECT 47.550 12.720 51.550 12.890 ;
        RECT 47.320 8.465 47.490 12.505 ;
        RECT 51.610 8.465 51.780 12.505 ;
        RECT 47.550 8.080 51.550 8.250 ;
        RECT 52.180 7.740 52.350 13.230 ;
        RECT 41.320 7.570 52.350 7.740 ;
        RECT 52.625 13.245 54.375 13.415 ;
        RECT 52.625 7.755 52.795 13.245 ;
        RECT 53.335 12.735 53.665 12.905 ;
        RECT 53.195 8.480 53.365 12.520 ;
        RECT 53.635 8.480 53.805 12.520 ;
        RECT 53.335 8.095 53.665 8.265 ;
        RECT 54.205 7.755 54.375 13.245 ;
        RECT 52.625 7.585 54.375 7.755 ;
        RECT 54.650 7.760 54.820 17.250 ;
        RECT 55.360 16.740 55.690 16.910 ;
        RECT 55.220 8.485 55.390 16.525 ;
        RECT 55.660 8.485 55.830 16.525 ;
        RECT 55.360 8.100 55.690 8.270 ;
        RECT 56.230 7.760 56.400 17.250 ;
        RECT 57.855 17.260 84.400 17.420 ;
        RECT 57.855 17.235 70.600 17.260 ;
        RECT 57.855 17.005 62.180 17.235 ;
        RECT 54.650 7.590 56.400 7.760 ;
        RECT 57.890 7.745 58.060 17.005 ;
        RECT 58.785 16.435 60.825 16.605 ;
        RECT 58.400 8.375 58.570 16.375 ;
        RECT 61.040 8.375 61.210 16.375 ;
        RECT 58.785 8.145 60.825 8.315 ;
        RECT 61.550 7.745 61.720 17.005 ;
        RECT 57.890 7.575 61.720 7.745 ;
        RECT 62.010 7.745 62.180 17.005 ;
        RECT 62.810 16.725 64.810 16.895 ;
        RECT 62.580 8.470 62.750 16.510 ;
        RECT 64.870 8.470 65.040 16.510 ;
        RECT 62.810 8.085 64.810 8.255 ;
        RECT 65.440 7.745 65.610 17.235 ;
        RECT 66.240 16.725 68.240 16.895 ;
        RECT 66.010 8.470 66.180 16.510 ;
        RECT 68.300 8.470 68.470 16.510 ;
        RECT 68.870 15.665 70.600 17.235 ;
        RECT 82.650 17.250 84.400 17.260 ;
        RECT 68.870 15.495 77.335 15.665 ;
        RECT 68.870 14.085 70.675 15.495 ;
        RECT 71.015 14.625 71.185 14.955 ;
        RECT 71.400 14.925 76.440 15.095 ;
        RECT 71.400 14.485 76.440 14.655 ;
        RECT 76.655 14.625 76.825 14.955 ;
        RECT 77.165 14.085 77.335 15.495 ;
        RECT 68.870 13.915 77.335 14.085 ;
        RECT 68.870 13.400 70.600 13.915 ;
        RECT 68.870 13.285 80.350 13.400 ;
        RECT 66.240 8.085 68.240 8.255 ;
        RECT 68.870 7.745 69.040 13.285 ;
        RECT 62.010 7.575 69.040 7.745 ;
        RECT 69.320 13.230 80.350 13.285 ;
        RECT 69.320 7.740 69.490 13.230 ;
        RECT 70.120 12.720 74.120 12.890 ;
        RECT 69.890 8.465 70.060 12.505 ;
        RECT 74.180 8.465 74.350 12.505 ;
        RECT 70.120 8.080 74.120 8.250 ;
        RECT 74.750 7.740 74.920 13.230 ;
        RECT 75.550 12.720 79.550 12.890 ;
        RECT 75.320 8.465 75.490 12.505 ;
        RECT 79.610 8.465 79.780 12.505 ;
        RECT 75.550 8.080 79.550 8.250 ;
        RECT 80.180 7.740 80.350 13.230 ;
        RECT 69.320 7.570 80.350 7.740 ;
        RECT 80.625 13.245 82.375 13.415 ;
        RECT 80.625 7.755 80.795 13.245 ;
        RECT 81.335 12.735 81.665 12.905 ;
        RECT 81.195 8.480 81.365 12.520 ;
        RECT 81.635 8.480 81.805 12.520 ;
        RECT 81.335 8.095 81.665 8.265 ;
        RECT 82.205 7.755 82.375 13.245 ;
        RECT 80.625 7.585 82.375 7.755 ;
        RECT 82.650 7.760 82.820 17.250 ;
        RECT 83.360 16.740 83.690 16.910 ;
        RECT 83.220 8.485 83.390 16.525 ;
        RECT 83.660 8.485 83.830 16.525 ;
        RECT 83.360 8.100 83.690 8.270 ;
        RECT 84.230 7.760 84.400 17.250 ;
        RECT 85.855 17.260 112.400 17.420 ;
        RECT 85.855 17.235 98.600 17.260 ;
        RECT 85.855 17.005 90.180 17.235 ;
        RECT 82.650 7.590 84.400 7.760 ;
        RECT 85.890 7.745 86.060 17.005 ;
        RECT 86.785 16.435 88.825 16.605 ;
        RECT 86.400 8.375 86.570 16.375 ;
        RECT 89.040 8.375 89.210 16.375 ;
        RECT 86.785 8.145 88.825 8.315 ;
        RECT 89.550 7.745 89.720 17.005 ;
        RECT 85.890 7.575 89.720 7.745 ;
        RECT 90.010 7.745 90.180 17.005 ;
        RECT 90.810 16.725 92.810 16.895 ;
        RECT 90.580 8.470 90.750 16.510 ;
        RECT 92.870 8.470 93.040 16.510 ;
        RECT 90.810 8.085 92.810 8.255 ;
        RECT 93.440 7.745 93.610 17.235 ;
        RECT 94.240 16.725 96.240 16.895 ;
        RECT 94.010 8.470 94.180 16.510 ;
        RECT 96.300 8.470 96.470 16.510 ;
        RECT 96.870 15.665 98.600 17.235 ;
        RECT 110.650 17.250 112.400 17.260 ;
        RECT 96.870 15.495 105.335 15.665 ;
        RECT 96.870 14.085 98.675 15.495 ;
        RECT 99.015 14.625 99.185 14.955 ;
        RECT 99.400 14.925 104.440 15.095 ;
        RECT 99.400 14.485 104.440 14.655 ;
        RECT 104.655 14.625 104.825 14.955 ;
        RECT 105.165 14.085 105.335 15.495 ;
        RECT 96.870 13.915 105.335 14.085 ;
        RECT 96.870 13.400 98.600 13.915 ;
        RECT 96.870 13.285 108.350 13.400 ;
        RECT 94.240 8.085 96.240 8.255 ;
        RECT 96.870 7.745 97.040 13.285 ;
        RECT 90.010 7.575 97.040 7.745 ;
        RECT 97.320 13.230 108.350 13.285 ;
        RECT 97.320 7.740 97.490 13.230 ;
        RECT 98.120 12.720 102.120 12.890 ;
        RECT 97.890 8.465 98.060 12.505 ;
        RECT 102.180 8.465 102.350 12.505 ;
        RECT 98.120 8.080 102.120 8.250 ;
        RECT 102.750 7.740 102.920 13.230 ;
        RECT 103.550 12.720 107.550 12.890 ;
        RECT 103.320 8.465 103.490 12.505 ;
        RECT 107.610 8.465 107.780 12.505 ;
        RECT 103.550 8.080 107.550 8.250 ;
        RECT 108.180 7.740 108.350 13.230 ;
        RECT 97.320 7.570 108.350 7.740 ;
        RECT 108.625 13.245 110.375 13.415 ;
        RECT 108.625 7.755 108.795 13.245 ;
        RECT 109.335 12.735 109.665 12.905 ;
        RECT 109.195 8.480 109.365 12.520 ;
        RECT 109.635 8.480 109.805 12.520 ;
        RECT 109.335 8.095 109.665 8.265 ;
        RECT 110.205 7.755 110.375 13.245 ;
        RECT 108.625 7.585 110.375 7.755 ;
        RECT 110.650 7.760 110.820 17.250 ;
        RECT 111.360 16.740 111.690 16.910 ;
        RECT 111.220 8.485 111.390 16.525 ;
        RECT 111.660 8.485 111.830 16.525 ;
        RECT 111.360 8.100 111.690 8.270 ;
        RECT 112.230 7.760 112.400 17.250 ;
        RECT 113.855 17.260 140.400 17.420 ;
        RECT 113.855 17.235 126.600 17.260 ;
        RECT 113.855 17.005 118.180 17.235 ;
        RECT 110.650 7.590 112.400 7.760 ;
        RECT 113.890 7.745 114.060 17.005 ;
        RECT 114.785 16.435 116.825 16.605 ;
        RECT 114.400 8.375 114.570 16.375 ;
        RECT 117.040 8.375 117.210 16.375 ;
        RECT 114.785 8.145 116.825 8.315 ;
        RECT 117.550 7.745 117.720 17.005 ;
        RECT 113.890 7.575 117.720 7.745 ;
        RECT 118.010 7.745 118.180 17.005 ;
        RECT 118.810 16.725 120.810 16.895 ;
        RECT 118.580 8.470 118.750 16.510 ;
        RECT 120.870 8.470 121.040 16.510 ;
        RECT 118.810 8.085 120.810 8.255 ;
        RECT 121.440 7.745 121.610 17.235 ;
        RECT 122.240 16.725 124.240 16.895 ;
        RECT 122.010 8.470 122.180 16.510 ;
        RECT 124.300 8.470 124.470 16.510 ;
        RECT 124.870 15.665 126.600 17.235 ;
        RECT 138.650 17.250 140.400 17.260 ;
        RECT 124.870 15.495 133.335 15.665 ;
        RECT 124.870 14.085 126.675 15.495 ;
        RECT 127.015 14.625 127.185 14.955 ;
        RECT 127.400 14.925 132.440 15.095 ;
        RECT 127.400 14.485 132.440 14.655 ;
        RECT 132.655 14.625 132.825 14.955 ;
        RECT 133.165 14.085 133.335 15.495 ;
        RECT 124.870 13.915 133.335 14.085 ;
        RECT 124.870 13.400 126.600 13.915 ;
        RECT 124.870 13.285 136.350 13.400 ;
        RECT 122.240 8.085 124.240 8.255 ;
        RECT 124.870 7.745 125.040 13.285 ;
        RECT 118.010 7.575 125.040 7.745 ;
        RECT 125.320 13.230 136.350 13.285 ;
        RECT 125.320 7.740 125.490 13.230 ;
        RECT 126.120 12.720 130.120 12.890 ;
        RECT 125.890 8.465 126.060 12.505 ;
        RECT 130.180 8.465 130.350 12.505 ;
        RECT 126.120 8.080 130.120 8.250 ;
        RECT 130.750 7.740 130.920 13.230 ;
        RECT 131.550 12.720 135.550 12.890 ;
        RECT 131.320 8.465 131.490 12.505 ;
        RECT 135.610 8.465 135.780 12.505 ;
        RECT 131.550 8.080 135.550 8.250 ;
        RECT 136.180 7.740 136.350 13.230 ;
        RECT 125.320 7.570 136.350 7.740 ;
        RECT 136.625 13.245 138.375 13.415 ;
        RECT 136.625 7.755 136.795 13.245 ;
        RECT 137.335 12.735 137.665 12.905 ;
        RECT 137.195 8.480 137.365 12.520 ;
        RECT 137.635 8.480 137.805 12.520 ;
        RECT 137.335 8.095 137.665 8.265 ;
        RECT 138.205 7.755 138.375 13.245 ;
        RECT 136.625 7.585 138.375 7.755 ;
        RECT 138.650 7.760 138.820 17.250 ;
        RECT 139.360 16.740 139.690 16.910 ;
        RECT 139.220 8.485 139.390 16.525 ;
        RECT 139.660 8.485 139.830 16.525 ;
        RECT 139.360 8.100 139.690 8.270 ;
        RECT 140.230 7.760 140.400 17.250 ;
        RECT 138.650 7.590 140.400 7.760 ;
        RECT 2.550 6.665 24.440 6.835 ;
        RECT 2.550 3.265 2.720 6.665 ;
        RECT 3.350 6.155 7.350 6.325 ;
        RECT 3.120 3.945 3.290 5.985 ;
        RECT 7.410 3.945 7.580 5.985 ;
        RECT 3.350 3.605 7.350 3.775 ;
        RECT 7.980 3.265 8.150 6.665 ;
        RECT 8.780 6.155 12.780 6.325 ;
        RECT 8.550 3.945 8.720 5.985 ;
        RECT 12.840 3.945 13.010 5.985 ;
        RECT 8.780 3.605 12.780 3.775 ;
        RECT 13.410 3.265 13.580 6.665 ;
        RECT 14.210 6.155 18.210 6.325 ;
        RECT 13.980 3.945 14.150 5.985 ;
        RECT 18.270 3.945 18.440 5.985 ;
        RECT 14.210 3.605 18.210 3.775 ;
        RECT 18.840 3.265 19.010 6.665 ;
        RECT 19.640 6.155 23.640 6.325 ;
        RECT 19.410 3.945 19.580 5.985 ;
        RECT 23.700 3.945 23.870 5.985 ;
        RECT 24.270 4.240 24.440 6.665 ;
        RECT 24.710 6.670 26.460 6.840 ;
        RECT 24.710 4.270 24.880 6.670 ;
        RECT 25.420 6.160 25.750 6.330 ;
        RECT 25.280 4.950 25.450 5.990 ;
        RECT 25.720 4.950 25.890 5.990 ;
        RECT 25.420 4.610 25.750 4.780 ;
        RECT 26.290 4.270 26.460 6.670 ;
        RECT 24.710 4.240 26.460 4.270 ;
        RECT 26.735 6.675 28.485 6.845 ;
        RECT 26.735 4.240 26.905 6.675 ;
        RECT 27.445 6.165 27.775 6.335 ;
        RECT 19.640 3.605 23.640 3.775 ;
        RECT 24.270 3.275 26.905 4.240 ;
        RECT 27.305 3.955 27.475 5.995 ;
        RECT 27.745 3.955 27.915 5.995 ;
        RECT 27.445 3.615 27.775 3.785 ;
        RECT 28.315 3.275 28.485 6.675 ;
        RECT 24.270 3.265 28.485 3.275 ;
        RECT 2.550 3.245 28.485 3.265 ;
        RECT 30.550 6.665 52.440 6.835 ;
        RECT 30.550 3.265 30.720 6.665 ;
        RECT 31.350 6.155 35.350 6.325 ;
        RECT 31.120 3.945 31.290 5.985 ;
        RECT 35.410 3.945 35.580 5.985 ;
        RECT 31.350 3.605 35.350 3.775 ;
        RECT 35.980 3.265 36.150 6.665 ;
        RECT 36.780 6.155 40.780 6.325 ;
        RECT 36.550 3.945 36.720 5.985 ;
        RECT 40.840 3.945 41.010 5.985 ;
        RECT 36.780 3.605 40.780 3.775 ;
        RECT 41.410 3.265 41.580 6.665 ;
        RECT 42.210 6.155 46.210 6.325 ;
        RECT 41.980 3.945 42.150 5.985 ;
        RECT 46.270 3.945 46.440 5.985 ;
        RECT 42.210 3.605 46.210 3.775 ;
        RECT 46.840 3.265 47.010 6.665 ;
        RECT 47.640 6.155 51.640 6.325 ;
        RECT 47.410 3.945 47.580 5.985 ;
        RECT 51.700 3.945 51.870 5.985 ;
        RECT 52.270 4.240 52.440 6.665 ;
        RECT 52.710 6.670 54.460 6.840 ;
        RECT 52.710 4.270 52.880 6.670 ;
        RECT 53.420 6.160 53.750 6.330 ;
        RECT 53.280 4.950 53.450 5.990 ;
        RECT 53.720 4.950 53.890 5.990 ;
        RECT 53.420 4.610 53.750 4.780 ;
        RECT 54.290 4.270 54.460 6.670 ;
        RECT 52.710 4.240 54.460 4.270 ;
        RECT 54.735 6.675 56.485 6.845 ;
        RECT 54.735 4.240 54.905 6.675 ;
        RECT 55.445 6.165 55.775 6.335 ;
        RECT 47.640 3.605 51.640 3.775 ;
        RECT 52.270 3.275 54.905 4.240 ;
        RECT 55.305 3.955 55.475 5.995 ;
        RECT 55.745 3.955 55.915 5.995 ;
        RECT 55.445 3.615 55.775 3.785 ;
        RECT 56.315 3.275 56.485 6.675 ;
        RECT 52.270 3.265 56.485 3.275 ;
        RECT 30.550 3.245 56.485 3.265 ;
        RECT 58.550 6.665 80.440 6.835 ;
        RECT 58.550 3.265 58.720 6.665 ;
        RECT 59.350 6.155 63.350 6.325 ;
        RECT 59.120 3.945 59.290 5.985 ;
        RECT 63.410 3.945 63.580 5.985 ;
        RECT 59.350 3.605 63.350 3.775 ;
        RECT 63.980 3.265 64.150 6.665 ;
        RECT 64.780 6.155 68.780 6.325 ;
        RECT 64.550 3.945 64.720 5.985 ;
        RECT 68.840 3.945 69.010 5.985 ;
        RECT 64.780 3.605 68.780 3.775 ;
        RECT 69.410 3.265 69.580 6.665 ;
        RECT 70.210 6.155 74.210 6.325 ;
        RECT 69.980 3.945 70.150 5.985 ;
        RECT 74.270 3.945 74.440 5.985 ;
        RECT 70.210 3.605 74.210 3.775 ;
        RECT 74.840 3.265 75.010 6.665 ;
        RECT 75.640 6.155 79.640 6.325 ;
        RECT 75.410 3.945 75.580 5.985 ;
        RECT 79.700 3.945 79.870 5.985 ;
        RECT 80.270 4.240 80.440 6.665 ;
        RECT 80.710 6.670 82.460 6.840 ;
        RECT 80.710 4.270 80.880 6.670 ;
        RECT 81.420 6.160 81.750 6.330 ;
        RECT 81.280 4.950 81.450 5.990 ;
        RECT 81.720 4.950 81.890 5.990 ;
        RECT 81.420 4.610 81.750 4.780 ;
        RECT 82.290 4.270 82.460 6.670 ;
        RECT 80.710 4.240 82.460 4.270 ;
        RECT 82.735 6.675 84.485 6.845 ;
        RECT 82.735 4.240 82.905 6.675 ;
        RECT 83.445 6.165 83.775 6.335 ;
        RECT 75.640 3.605 79.640 3.775 ;
        RECT 80.270 3.275 82.905 4.240 ;
        RECT 83.305 3.955 83.475 5.995 ;
        RECT 83.745 3.955 83.915 5.995 ;
        RECT 83.445 3.615 83.775 3.785 ;
        RECT 84.315 3.275 84.485 6.675 ;
        RECT 80.270 3.265 84.485 3.275 ;
        RECT 58.550 3.245 84.485 3.265 ;
        RECT 86.550 6.665 108.440 6.835 ;
        RECT 86.550 3.265 86.720 6.665 ;
        RECT 87.350 6.155 91.350 6.325 ;
        RECT 87.120 3.945 87.290 5.985 ;
        RECT 91.410 3.945 91.580 5.985 ;
        RECT 87.350 3.605 91.350 3.775 ;
        RECT 91.980 3.265 92.150 6.665 ;
        RECT 92.780 6.155 96.780 6.325 ;
        RECT 92.550 3.945 92.720 5.985 ;
        RECT 96.840 3.945 97.010 5.985 ;
        RECT 92.780 3.605 96.780 3.775 ;
        RECT 97.410 3.265 97.580 6.665 ;
        RECT 98.210 6.155 102.210 6.325 ;
        RECT 97.980 3.945 98.150 5.985 ;
        RECT 102.270 3.945 102.440 5.985 ;
        RECT 98.210 3.605 102.210 3.775 ;
        RECT 102.840 3.265 103.010 6.665 ;
        RECT 103.640 6.155 107.640 6.325 ;
        RECT 103.410 3.945 103.580 5.985 ;
        RECT 107.700 3.945 107.870 5.985 ;
        RECT 108.270 4.240 108.440 6.665 ;
        RECT 108.710 6.670 110.460 6.840 ;
        RECT 108.710 4.270 108.880 6.670 ;
        RECT 109.420 6.160 109.750 6.330 ;
        RECT 109.280 4.950 109.450 5.990 ;
        RECT 109.720 4.950 109.890 5.990 ;
        RECT 109.420 4.610 109.750 4.780 ;
        RECT 110.290 4.270 110.460 6.670 ;
        RECT 108.710 4.240 110.460 4.270 ;
        RECT 110.735 6.675 112.485 6.845 ;
        RECT 110.735 4.240 110.905 6.675 ;
        RECT 111.445 6.165 111.775 6.335 ;
        RECT 103.640 3.605 107.640 3.775 ;
        RECT 108.270 3.275 110.905 4.240 ;
        RECT 111.305 3.955 111.475 5.995 ;
        RECT 111.745 3.955 111.915 5.995 ;
        RECT 111.445 3.615 111.775 3.785 ;
        RECT 112.315 3.275 112.485 6.675 ;
        RECT 108.270 3.265 112.485 3.275 ;
        RECT 86.550 3.245 112.485 3.265 ;
        RECT 114.550 6.665 136.440 6.835 ;
        RECT 114.550 3.265 114.720 6.665 ;
        RECT 115.350 6.155 119.350 6.325 ;
        RECT 115.120 3.945 115.290 5.985 ;
        RECT 119.410 3.945 119.580 5.985 ;
        RECT 115.350 3.605 119.350 3.775 ;
        RECT 119.980 3.265 120.150 6.665 ;
        RECT 120.780 6.155 124.780 6.325 ;
        RECT 120.550 3.945 120.720 5.985 ;
        RECT 124.840 3.945 125.010 5.985 ;
        RECT 120.780 3.605 124.780 3.775 ;
        RECT 125.410 3.265 125.580 6.665 ;
        RECT 126.210 6.155 130.210 6.325 ;
        RECT 125.980 3.945 126.150 5.985 ;
        RECT 130.270 3.945 130.440 5.985 ;
        RECT 126.210 3.605 130.210 3.775 ;
        RECT 130.840 3.265 131.010 6.665 ;
        RECT 131.640 6.155 135.640 6.325 ;
        RECT 131.410 3.945 131.580 5.985 ;
        RECT 135.700 3.945 135.870 5.985 ;
        RECT 136.270 4.240 136.440 6.665 ;
        RECT 136.710 6.670 138.460 6.840 ;
        RECT 136.710 4.270 136.880 6.670 ;
        RECT 137.420 6.160 137.750 6.330 ;
        RECT 137.280 4.950 137.450 5.990 ;
        RECT 137.720 4.950 137.890 5.990 ;
        RECT 137.420 4.610 137.750 4.780 ;
        RECT 138.290 4.270 138.460 6.670 ;
        RECT 136.710 4.240 138.460 4.270 ;
        RECT 138.735 6.675 140.485 6.845 ;
        RECT 138.735 4.240 138.905 6.675 ;
        RECT 139.445 6.165 139.775 6.335 ;
        RECT 131.640 3.605 135.640 3.775 ;
        RECT 136.270 3.275 138.905 4.240 ;
        RECT 139.305 3.955 139.475 5.995 ;
        RECT 139.745 3.955 139.915 5.995 ;
        RECT 139.445 3.615 139.775 3.785 ;
        RECT 140.315 3.275 140.485 6.675 ;
        RECT 136.270 3.265 140.485 3.275 ;
        RECT 114.550 3.245 140.485 3.265 ;
        RECT 1.895 3.105 28.485 3.245 ;
        RECT 29.895 3.105 56.485 3.245 ;
        RECT 57.895 3.105 84.485 3.245 ;
        RECT 85.895 3.105 112.485 3.245 ;
        RECT 113.895 3.105 140.485 3.245 ;
        RECT 1.895 2.380 28.475 3.105 ;
        RECT 29.895 2.380 56.475 3.105 ;
        RECT 57.895 2.380 84.475 3.105 ;
        RECT 85.895 2.380 112.475 3.105 ;
        RECT 113.895 2.380 140.475 3.105 ;
      LAYER met1 ;
        RECT 95.140 100.385 96.200 100.395 ;
        RECT 77.490 100.380 96.200 100.385 ;
        RECT 77.490 99.765 96.240 100.380 ;
        RECT 78.645 99.430 88.475 99.765 ;
        RECT 95.140 99.735 96.240 99.765 ;
        RECT 78.645 99.365 86.675 99.430 ;
        RECT 78.605 99.205 86.675 99.365 ;
        RECT 78.605 99.135 86.605 99.205 ;
        RECT 78.170 99.070 78.400 99.085 ;
        RECT 78.130 98.975 78.400 99.070 ;
        RECT 86.810 98.975 87.040 99.085 ;
        RECT 78.130 98.250 87.040 98.975 ;
        RECT 78.170 98.220 87.040 98.250 ;
        RECT 78.170 98.125 78.400 98.220 ;
        RECT 86.810 98.125 87.040 98.220 ;
        RECT 87.380 98.965 88.475 99.430 ;
        RECT 89.040 99.260 89.370 99.540 ;
        RECT 90.590 99.265 90.920 99.545 ;
        RECT 89.040 99.255 89.330 99.260 ;
        RECT 90.620 99.255 90.910 99.265 ;
        RECT 92.180 99.260 92.510 99.540 ;
        RECT 92.200 99.255 92.490 99.260 ;
        RECT 94.430 99.195 94.760 99.475 ;
        RECT 94.460 99.175 94.750 99.195 ;
        RECT 88.850 98.965 89.080 99.050 ;
        RECT 78.605 97.845 86.605 98.075 ;
        RECT 78.665 97.560 86.600 97.845 ;
        RECT 79.830 95.920 80.415 97.560 ;
        RECT 87.380 97.330 89.080 98.965 ;
        RECT 87.900 97.080 89.080 97.330 ;
        RECT 80.770 96.075 86.730 96.305 ;
        RECT 79.830 95.915 80.550 95.920 ;
        RECT 79.830 95.885 80.720 95.915 ;
        RECT 80.915 95.885 86.545 96.075 ;
        RECT 79.830 95.230 86.545 95.885 ;
        RECT 86.780 95.875 87.010 95.915 ;
        RECT 80.185 95.015 86.545 95.230 ;
        RECT 80.490 94.985 86.545 95.015 ;
        RECT 86.765 95.000 87.490 95.875 ;
        RECT 80.490 94.915 80.720 94.985 ;
        RECT 80.915 94.755 86.545 94.985 ;
        RECT 86.780 94.915 87.455 95.000 ;
        RECT 86.900 94.890 87.455 94.915 ;
        RECT 80.770 94.525 86.730 94.755 ;
        RECT 77.920 93.685 78.470 93.695 ;
        RECT 72.905 93.610 76.835 93.630 ;
        RECT 77.720 93.610 78.470 93.685 ;
        RECT 72.905 93.145 78.575 93.610 ;
        RECT 72.905 93.135 76.980 93.145 ;
        RECT 72.830 93.090 76.980 93.135 ;
        RECT 72.830 92.920 76.835 93.090 ;
        RECT 72.830 92.905 76.830 92.920 ;
        RECT 77.545 92.895 78.525 93.145 ;
        RECT 78.790 93.055 86.750 93.285 ;
        RECT 72.440 92.710 72.670 92.855 ;
        RECT 76.990 92.710 77.220 92.855 ;
        RECT 72.440 92.010 77.220 92.710 ;
        RECT 72.440 91.895 72.670 92.010 ;
        RECT 76.990 91.895 77.220 92.010 ;
        RECT 77.545 91.975 78.740 92.895 ;
        RECT 72.830 91.615 76.830 91.845 ;
        RECT 72.925 91.295 76.790 91.615 ;
        RECT 77.545 91.570 78.360 91.975 ;
        RECT 78.510 91.895 78.740 91.975 ;
        RECT 78.965 91.735 86.555 93.055 ;
        RECT 87.120 92.955 87.455 94.890 ;
        RECT 86.920 92.895 87.455 92.955 ;
        RECT 86.800 92.885 87.455 92.895 ;
        RECT 86.800 92.690 87.560 92.885 ;
        RECT 86.800 92.220 87.900 92.690 ;
        RECT 86.800 92.010 87.560 92.220 ;
        RECT 86.800 91.895 87.030 92.010 ;
        RECT 77.710 91.535 78.360 91.570 ;
        RECT 72.925 91.290 77.245 91.295 ;
        RECT 72.925 91.055 77.380 91.290 ;
        RECT 73.905 90.870 77.380 91.055 ;
        RECT 77.825 91.190 78.315 91.535 ;
        RECT 78.790 91.505 86.750 91.735 ;
        RECT 77.825 91.050 79.120 91.190 ;
        RECT 78.050 90.925 80.015 91.050 ;
        RECT 81.195 91.045 82.090 91.505 ;
        RECT 76.935 90.675 77.380 90.870 ;
        RECT 78.905 90.835 80.015 90.925 ;
        RECT 78.905 90.675 80.245 90.835 ;
        RECT 76.935 90.585 78.005 90.675 ;
        RECT 76.950 90.460 78.005 90.585 ;
        RECT 76.950 90.265 78.720 90.460 ;
        RECT 75.700 90.200 76.585 90.230 ;
        RECT 73.000 90.070 76.635 90.200 ;
        RECT 73.000 89.700 76.640 90.070 ;
        RECT 77.560 89.970 78.720 90.265 ;
        RECT 77.560 89.745 78.860 89.970 ;
        RECT 73.010 89.485 73.950 89.700 ;
        RECT 75.700 89.485 76.640 89.700 ;
        RECT 78.245 89.690 78.860 89.745 ;
        RECT 79.310 89.735 80.245 90.675 ;
        RECT 81.175 90.545 82.090 91.045 ;
        RECT 81.175 90.100 86.740 90.545 ;
        RECT 81.195 89.980 86.740 90.100 ;
        RECT 72.995 89.255 73.995 89.485 ;
        RECT 75.655 89.255 76.655 89.485 ;
        RECT 78.245 89.355 78.870 89.690 ;
        RECT 79.310 89.505 80.270 89.735 ;
        RECT 81.195 89.690 86.825 89.980 ;
        RECT 79.310 89.450 80.245 89.505 ;
        RECT 72.560 89.020 72.790 89.205 ;
        RECT 74.200 89.020 74.430 89.205 ;
        RECT 72.560 87.410 74.430 89.020 ;
        RECT 72.560 87.245 72.790 87.410 ;
        RECT 72.940 87.195 73.915 87.410 ;
        RECT 74.200 87.245 74.430 87.410 ;
        RECT 75.220 89.000 75.450 89.205 ;
        RECT 75.875 89.000 76.265 89.005 ;
        RECT 76.860 89.000 77.090 89.205 ;
        RECT 78.455 89.110 78.870 89.355 ;
        RECT 79.030 89.110 79.260 89.300 ;
        RECT 75.220 87.390 77.090 89.000 ;
        RECT 78.420 89.065 79.260 89.110 ;
        RECT 75.220 87.245 75.450 87.390 ;
        RECT 75.590 87.245 77.090 87.390 ;
        RECT 72.940 86.965 73.995 87.195 ;
        RECT 75.590 87.190 76.935 87.245 ;
        RECT 75.590 86.995 76.795 87.190 ;
        RECT 75.590 86.965 76.655 86.995 ;
        RECT 72.940 86.125 73.950 86.965 ;
        RECT 72.940 85.615 73.940 86.125 ;
        RECT 72.940 85.580 73.925 85.615 ;
        RECT 72.940 85.155 73.915 85.580 ;
        RECT 75.590 85.155 76.565 86.965 ;
        RECT 77.530 86.450 78.235 88.275 ;
        RECT 78.420 87.350 79.270 89.065 ;
        RECT 78.420 87.300 79.260 87.350 ;
        RECT 78.420 87.285 79.200 87.300 ;
        RECT 79.425 87.095 80.170 89.450 ;
        RECT 80.320 89.120 80.550 89.300 ;
        RECT 81.195 89.120 82.090 89.690 ;
        RECT 83.155 89.650 86.825 89.690 ;
        RECT 83.155 89.455 84.160 89.650 ;
        RECT 85.820 89.455 86.825 89.650 ;
        RECT 83.075 89.310 84.160 89.455 ;
        RECT 85.735 89.315 86.825 89.455 ;
        RECT 83.075 89.225 84.075 89.310 ;
        RECT 85.735 89.225 86.735 89.315 ;
        RECT 80.320 87.485 82.235 89.120 ;
        RECT 82.640 89.070 82.870 89.175 ;
        RECT 84.280 89.070 84.510 89.175 ;
        RECT 80.320 87.300 82.335 87.485 ;
        RECT 80.380 87.295 82.335 87.300 ;
        RECT 79.310 86.865 80.270 87.095 ;
        RECT 79.425 86.850 80.170 86.865 ;
        RECT 80.995 86.450 82.335 87.295 ;
        RECT 82.640 87.400 84.510 89.070 ;
        RECT 82.640 87.215 82.870 87.400 ;
        RECT 83.205 87.165 84.125 87.400 ;
        RECT 84.280 87.215 84.510 87.400 ;
        RECT 85.300 89.065 85.530 89.175 ;
        RECT 86.940 89.065 87.170 89.175 ;
        RECT 85.300 87.395 87.190 89.065 ;
        RECT 85.300 87.215 85.530 87.395 ;
        RECT 85.845 87.165 86.765 87.395 ;
        RECT 86.940 87.215 87.170 87.395 ;
        RECT 83.075 87.140 84.125 87.165 ;
        RECT 83.075 86.935 84.140 87.140 ;
        RECT 85.735 86.935 86.765 87.165 ;
        RECT 83.205 86.665 84.140 86.935 ;
        RECT 77.530 86.420 82.335 86.450 ;
        RECT 77.530 86.055 82.320 86.420 ;
        RECT 77.615 86.015 82.320 86.055 ;
        RECT 83.220 86.170 84.140 86.665 ;
        RECT 85.840 86.555 86.765 86.935 ;
        RECT 72.930 84.925 73.930 85.155 ;
        RECT 75.500 85.050 76.565 85.155 ;
        RECT 77.060 85.105 79.075 85.415 ;
        RECT 79.710 85.130 80.350 86.015 ;
        RECT 83.220 85.635 84.575 86.170 ;
        RECT 80.695 85.430 82.610 85.565 ;
        RECT 80.695 85.155 82.620 85.430 ;
        RECT 83.220 85.155 84.140 85.635 ;
        RECT 85.840 85.155 86.760 86.555 ;
        RECT 87.425 85.605 88.035 86.210 ;
        RECT 75.500 84.925 76.500 85.050 ;
        RECT 77.060 85.045 77.500 85.105 ;
        RECT 77.060 84.885 77.370 85.045 ;
        RECT 78.050 85.025 79.075 85.105 ;
        RECT 78.070 84.925 79.070 85.025 ;
        RECT 72.540 84.785 72.770 84.875 ;
        RECT 74.090 84.785 74.320 84.875 ;
        RECT 72.540 79.100 74.320 84.785 ;
        RECT 72.540 78.915 72.770 79.100 ;
        RECT 74.090 78.915 74.320 79.100 ;
        RECT 75.110 84.775 75.340 84.875 ;
        RECT 76.660 84.775 76.890 84.875 ;
        RECT 75.110 79.090 76.890 84.775 ;
        RECT 75.110 78.915 75.340 79.090 ;
        RECT 76.660 78.915 76.890 79.090 ;
        RECT 72.930 78.760 73.930 78.865 ;
        RECT 72.930 78.635 73.940 78.760 ;
        RECT 75.500 78.755 76.500 78.865 ;
        RECT 72.960 78.620 73.940 78.635 ;
        RECT 75.415 78.730 76.500 78.755 ;
        RECT 77.060 78.735 77.330 84.885 ;
        RECT 79.675 84.875 80.350 85.130 ;
        RECT 80.640 85.140 82.620 85.155 ;
        RECT 80.640 84.925 81.640 85.140 ;
        RECT 82.275 85.115 82.620 85.140 ;
        RECT 77.680 84.765 77.910 84.875 ;
        RECT 79.230 84.765 79.460 84.875 ;
        RECT 77.680 84.665 79.460 84.765 ;
        RECT 79.675 84.765 80.480 84.875 ;
        RECT 81.800 84.765 82.030 84.875 ;
        RECT 79.675 84.665 82.030 84.765 ;
        RECT 77.680 79.090 82.030 84.665 ;
        RECT 77.680 79.080 79.460 79.090 ;
        RECT 79.985 79.085 82.030 79.090 ;
        RECT 77.680 78.915 77.910 79.080 ;
        RECT 79.230 78.915 79.460 79.080 ;
        RECT 80.250 79.080 82.030 79.085 ;
        RECT 80.250 78.915 80.480 79.080 ;
        RECT 81.800 78.915 82.030 79.080 ;
        RECT 78.070 78.775 79.070 78.865 ;
        RECT 75.415 78.620 76.560 78.730 ;
        RECT 77.060 78.620 77.500 78.735 ;
        RECT 78.010 78.635 79.070 78.775 ;
        RECT 80.640 78.635 81.640 78.865 ;
        RECT 82.310 78.675 82.620 85.115 ;
        RECT 82.805 84.875 83.000 84.970 ;
        RECT 83.210 84.925 84.210 85.155 ;
        RECT 85.780 84.925 86.780 85.155 ;
        RECT 82.805 84.755 83.050 84.875 ;
        RECT 84.370 84.755 84.600 84.875 ;
        RECT 82.805 84.190 84.600 84.755 ;
        RECT 82.820 79.070 84.600 84.190 ;
        RECT 82.820 78.915 83.050 79.070 ;
        RECT 84.370 78.915 84.600 79.070 ;
        RECT 85.390 84.765 85.620 84.875 ;
        RECT 86.940 84.765 87.170 84.875 ;
        RECT 85.390 79.080 87.170 84.765 ;
        RECT 85.390 78.915 85.620 79.080 ;
        RECT 86.940 78.915 87.170 79.080 ;
        RECT 72.960 78.470 77.545 78.620 ;
        RECT 72.950 78.080 77.545 78.470 ;
        RECT 78.010 78.470 79.020 78.635 ;
        RECT 78.010 78.400 79.030 78.470 ;
        RECT 78.010 78.080 79.035 78.400 ;
        RECT 78.075 77.800 79.035 78.080 ;
        RECT 80.685 77.800 81.555 78.635 ;
        RECT 82.275 78.470 82.620 78.675 ;
        RECT 83.210 78.635 84.210 78.865 ;
        RECT 85.780 78.635 86.780 78.865 ;
        RECT 87.510 78.815 87.985 85.605 ;
        RECT 88.270 79.120 89.080 97.080 ;
        RECT 88.850 79.050 89.080 79.120 ;
        RECT 89.290 99.005 89.520 99.050 ;
        RECT 90.430 99.005 90.660 99.050 ;
        RECT 89.290 79.115 89.830 99.005 ;
        RECT 90.080 79.115 90.660 99.005 ;
        RECT 89.290 79.050 89.520 79.115 ;
        RECT 90.430 79.050 90.660 79.115 ;
        RECT 90.870 99.005 91.100 99.050 ;
        RECT 92.010 99.020 92.240 99.050 ;
        RECT 90.870 79.115 91.440 99.005 ;
        RECT 91.640 79.130 92.240 99.020 ;
        RECT 90.870 79.050 91.100 79.115 ;
        RECT 92.010 79.050 92.240 79.130 ;
        RECT 92.450 99.010 92.680 99.050 ;
        RECT 92.450 98.915 93.035 99.010 ;
        RECT 94.270 98.970 94.500 99.015 ;
        RECT 93.895 98.915 94.500 98.970 ;
        RECT 92.450 79.105 94.500 98.915 ;
        RECT 92.450 79.080 92.875 79.105 ;
        RECT 93.895 79.080 94.500 79.105 ;
        RECT 92.450 79.050 92.680 79.080 ;
        RECT 94.270 79.015 94.500 79.080 ;
        RECT 94.710 98.975 94.940 99.015 ;
        RECT 94.710 91.885 95.280 98.975 ;
        RECT 95.695 93.385 96.240 99.735 ;
        RECT 98.845 93.385 99.250 93.430 ;
        RECT 95.695 92.850 99.250 93.385 ;
        RECT 95.695 92.840 99.115 92.850 ;
        RECT 97.185 92.355 99.115 92.840 ;
        RECT 97.165 92.125 99.165 92.355 ;
        RECT 96.730 91.905 96.960 92.075 ;
        RECT 99.370 91.905 99.600 92.075 ;
        RECT 96.730 91.885 99.600 91.905 ;
        RECT 94.710 91.360 99.600 91.885 ;
        RECT 94.710 85.700 95.280 91.360 ;
        RECT 96.730 91.325 99.600 91.360 ;
        RECT 96.730 91.115 96.960 91.325 ;
        RECT 99.370 91.115 99.600 91.325 ;
        RECT 97.230 91.065 99.110 91.075 ;
        RECT 97.165 90.835 99.165 91.065 ;
        RECT 97.230 90.125 99.110 90.835 ;
        RECT 97.230 89.835 100.685 90.125 ;
        RECT 97.230 89.790 100.735 89.835 ;
        RECT 97.250 89.715 100.735 89.790 ;
        RECT 97.250 89.405 98.155 89.715 ;
        RECT 99.830 89.405 100.735 89.715 ;
        RECT 97.035 89.305 98.155 89.405 ;
        RECT 97.035 89.175 98.035 89.305 ;
        RECT 99.695 89.285 100.735 89.405 ;
        RECT 99.695 89.175 100.695 89.285 ;
        RECT 96.600 88.970 96.830 89.125 ;
        RECT 98.240 88.970 98.470 89.125 ;
        RECT 96.600 88.455 98.555 88.970 ;
        RECT 96.310 87.995 98.555 88.455 ;
        RECT 96.600 87.480 98.555 87.995 ;
        RECT 99.260 88.935 99.490 89.125 ;
        RECT 100.900 88.935 101.130 89.125 ;
        RECT 96.600 87.165 96.830 87.480 ;
        RECT 98.240 87.165 98.470 87.480 ;
        RECT 99.260 87.445 101.235 88.935 ;
        RECT 99.260 87.165 99.490 87.445 ;
        RECT 100.900 87.165 101.130 87.445 ;
        RECT 99.770 87.115 100.705 87.160 ;
        RECT 97.035 87.110 98.035 87.115 ;
        RECT 97.035 86.885 98.100 87.110 ;
        RECT 99.695 86.885 100.705 87.115 ;
        RECT 94.710 85.575 96.365 85.700 ;
        RECT 94.710 79.115 96.400 85.575 ;
        RECT 97.165 85.215 98.100 86.885 ;
        RECT 99.770 85.215 100.705 86.885 ;
        RECT 97.140 84.985 98.140 85.215 ;
        RECT 99.710 84.985 100.710 85.215 ;
        RECT 94.710 79.085 95.150 79.115 ;
        RECT 94.710 79.015 94.940 79.085 ;
        RECT 95.450 78.910 96.400 79.115 ;
        RECT 96.750 84.730 96.980 84.935 ;
        RECT 97.205 84.730 98.110 84.985 ;
        RECT 98.300 84.730 98.530 84.935 ;
        RECT 96.750 79.130 98.530 84.730 ;
        RECT 99.320 84.755 99.550 84.935 ;
        RECT 99.800 84.755 100.705 84.985 ;
        RECT 100.870 84.755 101.100 84.935 ;
        RECT 99.320 80.450 101.100 84.755 ;
        RECT 96.750 78.975 96.980 79.130 ;
        RECT 98.300 78.975 98.530 79.130 ;
        RECT 99.195 79.155 101.100 80.450 ;
        RECT 99.195 79.085 99.550 79.155 ;
        RECT 99.160 78.975 99.550 79.085 ;
        RECT 100.870 78.975 101.100 79.155 ;
        RECT 89.030 78.815 89.360 78.895 ;
        RECT 90.610 78.815 90.940 78.845 ;
        RECT 92.195 78.815 92.525 78.845 ;
        RECT 83.240 78.470 84.135 78.635 ;
        RECT 85.825 78.470 86.720 78.635 ;
        RECT 82.275 78.135 86.720 78.470 ;
        RECT 82.275 78.130 82.620 78.135 ;
        RECT 87.510 78.095 92.530 78.815 ;
        RECT 94.370 78.465 95.005 78.860 ;
        RECT 95.320 78.310 96.400 78.910 ;
        RECT 97.140 78.695 98.140 78.925 ;
        RECT 99.160 78.825 99.480 78.975 ;
        RECT 99.710 78.695 100.710 78.925 ;
        RECT 97.205 78.310 98.055 78.695 ;
        RECT 99.750 78.310 100.600 78.695 ;
        RECT 95.320 77.800 101.555 78.310 ;
        RECT 72.020 76.905 101.575 77.800 ;
        RECT 111.215 75.090 111.855 75.095 ;
        RECT 84.320 75.085 111.855 75.090 ;
        RECT 114.845 75.090 115.575 75.095 ;
        RECT 114.845 75.085 144.425 75.090 ;
        RECT 84.320 74.550 144.425 75.085 ;
        RECT 84.015 73.850 144.425 74.550 ;
        RECT 84.015 73.685 109.665 73.850 ;
        RECT 110.655 73.685 144.425 73.850 ;
        RECT 80.660 73.150 81.250 73.200 ;
        RECT 82.480 73.150 83.070 73.200 ;
        RECT 80.660 71.195 83.070 73.150 ;
        RECT 84.015 72.920 84.475 73.685 ;
        RECT 84.975 73.170 85.290 73.460 ;
        RECT 84.790 72.920 85.020 72.965 ;
        RECT 84.015 72.250 85.020 72.920 ;
        RECT 80.660 71.095 81.250 71.195 ;
        RECT 82.480 71.095 83.070 71.195 ;
        RECT 80.660 70.190 81.250 70.515 ;
        RECT 82.480 70.210 83.070 70.515 ;
        RECT 80.640 65.170 81.265 70.190 ;
        RECT 82.455 65.190 83.080 70.210 ;
        RECT 84.425 67.045 85.020 72.250 ;
        RECT 84.790 66.965 85.020 67.045 ;
        RECT 85.230 72.905 85.460 72.965 ;
        RECT 87.125 72.920 87.715 73.215 ;
        RECT 85.720 72.905 87.715 72.920 ;
        RECT 85.230 71.135 87.715 72.905 ;
        RECT 85.230 69.525 86.135 71.135 ;
        RECT 87.125 71.110 87.715 71.135 ;
        RECT 88.945 73.120 89.535 73.215 ;
        RECT 90.765 73.120 91.355 73.215 ;
        RECT 88.945 71.335 91.355 73.120 ;
        RECT 92.310 72.920 92.770 73.685 ;
        RECT 93.275 73.195 93.590 73.485 ;
        RECT 93.275 73.185 93.565 73.195 ;
        RECT 95.455 73.005 96.045 73.205 ;
        RECT 93.085 72.920 93.315 72.980 ;
        RECT 92.310 72.090 93.315 72.920 ;
        RECT 88.945 71.110 89.535 71.335 ;
        RECT 90.765 71.110 91.355 71.335 ;
        RECT 87.125 70.350 87.715 70.530 ;
        RECT 88.945 70.350 89.535 70.530 ;
        RECT 85.230 67.070 86.260 69.525 ;
        RECT 87.125 68.565 89.535 70.350 ;
        RECT 90.765 70.200 91.355 70.530 ;
        RECT 87.125 68.425 87.715 68.565 ;
        RECT 88.945 68.425 89.535 68.565 ;
        RECT 90.740 68.425 91.355 70.200 ;
        RECT 90.740 67.235 91.270 68.425 ;
        RECT 85.230 66.965 85.460 67.070 ;
        RECT 84.985 66.760 85.315 66.765 ;
        RECT 84.980 66.530 85.315 66.760 ;
        RECT 84.985 66.505 85.315 66.530 ;
        RECT 84.985 66.335 85.245 66.505 ;
        RECT 84.650 65.335 85.650 66.335 ;
        RECT 80.660 65.115 81.250 65.170 ;
        RECT 82.480 65.115 83.070 65.190 ;
        RECT 84.985 65.015 85.315 65.335 ;
        RECT 84.960 64.800 85.315 65.015 ;
        RECT 84.960 64.785 85.250 64.800 ;
        RECT 84.770 64.565 85.000 64.625 ;
        RECT 80.660 64.445 81.250 64.535 ;
        RECT 80.540 61.920 81.265 64.445 ;
        RECT 82.480 64.435 83.070 64.535 ;
        RECT 82.475 62.340 83.070 64.435 ;
        RECT 84.335 63.780 85.000 64.565 ;
        RECT 83.975 62.695 85.000 63.780 ;
        RECT 82.475 61.920 83.070 61.930 ;
        RECT 83.975 61.920 84.435 62.695 ;
        RECT 84.770 62.625 85.000 62.695 ;
        RECT 85.210 64.555 85.440 64.625 ;
        RECT 85.885 64.555 86.260 67.070 ;
        RECT 87.125 67.055 87.715 67.235 ;
        RECT 88.945 67.055 89.535 67.235 ;
        RECT 87.125 65.270 89.535 67.055 ;
        RECT 87.125 65.130 87.715 65.270 ;
        RECT 88.945 65.130 89.535 65.270 ;
        RECT 90.740 65.255 91.355 67.235 ;
        RECT 92.640 67.045 93.315 72.090 ;
        RECT 93.085 66.980 93.315 67.045 ;
        RECT 93.525 72.925 93.755 72.980 ;
        RECT 93.950 72.925 96.045 73.005 ;
        RECT 93.525 71.220 96.045 72.925 ;
        RECT 93.525 69.640 94.470 71.220 ;
        RECT 95.455 71.100 96.045 71.220 ;
        RECT 97.275 72.955 97.865 73.205 ;
        RECT 99.095 72.955 99.685 73.205 ;
        RECT 97.275 71.170 99.685 72.955 ;
        RECT 100.645 72.900 101.105 73.685 ;
        RECT 101.590 73.170 101.905 73.460 ;
        RECT 101.400 72.900 101.630 72.970 ;
        RECT 100.645 72.100 101.630 72.900 ;
        RECT 97.275 71.100 97.865 71.170 ;
        RECT 99.095 71.100 99.685 71.170 ;
        RECT 95.455 70.265 96.045 70.520 ;
        RECT 97.275 70.265 97.865 70.520 ;
        RECT 93.525 67.090 94.650 69.640 ;
        RECT 95.455 68.480 97.865 70.265 ;
        RECT 99.095 70.190 99.685 70.520 ;
        RECT 95.455 68.415 96.045 68.480 ;
        RECT 97.275 68.415 97.865 68.480 ;
        RECT 93.525 66.980 93.755 67.090 ;
        RECT 93.275 66.745 93.565 66.775 ;
        RECT 93.265 66.330 93.595 66.745 ;
        RECT 92.935 65.330 93.935 66.330 ;
        RECT 90.765 65.130 91.355 65.255 ;
        RECT 93.265 64.780 93.595 65.330 ;
        RECT 85.210 62.735 86.285 64.555 ;
        RECT 85.210 62.625 85.440 62.735 ;
        RECT 84.960 62.180 85.275 62.470 ;
        RECT 87.125 62.445 87.715 64.550 ;
        RECT 88.945 64.335 89.535 64.550 ;
        RECT 89.765 64.335 90.360 64.410 ;
        RECT 90.765 64.335 91.355 64.550 ;
        RECT 93.075 64.535 93.305 64.625 ;
        RECT 93.515 64.545 93.745 64.625 ;
        RECT 94.275 64.545 94.650 67.090 ;
        RECT 95.455 67.095 96.045 67.225 ;
        RECT 97.275 67.095 97.865 67.225 ;
        RECT 95.455 65.310 97.865 67.095 ;
        RECT 95.455 65.120 96.045 65.310 ;
        RECT 97.275 65.120 97.865 65.310 ;
        RECT 99.085 65.170 99.710 70.190 ;
        RECT 100.995 67.025 101.630 72.100 ;
        RECT 101.400 66.970 101.630 67.025 ;
        RECT 101.840 72.950 102.070 72.970 ;
        RECT 101.840 72.930 102.765 72.950 ;
        RECT 103.750 72.930 104.340 73.195 ;
        RECT 101.840 71.115 104.340 72.930 ;
        RECT 101.840 69.515 102.765 71.115 ;
        RECT 103.750 71.090 104.340 71.115 ;
        RECT 105.570 73.010 106.160 73.195 ;
        RECT 107.390 73.010 107.980 73.195 ;
        RECT 105.570 71.195 107.980 73.010 ;
        RECT 109.020 73.040 109.480 73.685 ;
        RECT 109.955 73.295 110.270 73.585 ;
        RECT 109.970 73.275 110.260 73.295 ;
        RECT 109.780 73.040 110.010 73.070 ;
        RECT 109.020 72.480 110.010 73.040 ;
        RECT 105.570 71.090 106.160 71.195 ;
        RECT 107.390 71.090 107.980 71.195 ;
        RECT 103.750 70.370 104.340 70.510 ;
        RECT 105.570 70.370 106.160 70.510 ;
        RECT 101.840 67.115 102.840 69.515 ;
        RECT 103.750 68.555 106.160 70.370 ;
        RECT 103.750 68.405 104.340 68.555 ;
        RECT 105.570 68.405 106.160 68.555 ;
        RECT 107.390 70.230 107.980 70.510 ;
        RECT 101.840 66.970 102.070 67.115 ;
        RECT 101.555 66.535 101.880 66.765 ;
        RECT 101.555 66.215 101.815 66.535 ;
        RECT 101.295 65.215 102.295 66.215 ;
        RECT 99.095 65.120 99.685 65.170 ;
        RECT 101.555 65.015 101.815 65.215 ;
        RECT 101.525 64.785 101.815 65.015 ;
        RECT 88.945 62.550 91.355 64.335 ;
        RECT 92.720 63.930 93.320 64.535 ;
        RECT 88.945 62.445 89.535 62.550 ;
        RECT 90.765 62.445 91.355 62.550 ;
        RECT 92.400 62.665 93.320 63.930 ;
        RECT 93.515 62.855 94.650 64.545 ;
        RECT 93.515 62.725 94.565 62.855 ;
        RECT 92.400 61.920 92.860 62.665 ;
        RECT 93.075 62.625 93.305 62.665 ;
        RECT 93.515 62.625 93.745 62.725 ;
        RECT 93.265 62.190 93.580 62.480 ;
        RECT 95.455 62.435 96.045 64.540 ;
        RECT 97.275 64.275 97.865 64.540 ;
        RECT 98.020 64.275 98.610 64.340 ;
        RECT 99.095 64.275 99.685 64.540 ;
        RECT 101.335 64.525 101.565 64.625 ;
        RECT 97.275 62.490 99.685 64.275 ;
        RECT 100.945 63.940 101.565 64.525 ;
        RECT 97.275 62.435 97.865 62.490 ;
        RECT 99.095 62.435 99.685 62.490 ;
        RECT 100.595 62.655 101.565 63.940 ;
        RECT 95.470 62.410 96.015 62.435 ;
        RECT 100.595 61.920 101.055 62.655 ;
        RECT 101.335 62.625 101.565 62.655 ;
        RECT 101.775 64.530 102.005 64.625 ;
        RECT 102.465 64.530 102.840 67.115 ;
        RECT 103.750 67.065 104.340 67.215 ;
        RECT 105.570 67.065 106.160 67.215 ;
        RECT 103.750 65.250 106.160 67.065 ;
        RECT 103.750 65.110 104.340 65.250 ;
        RECT 105.570 65.110 106.160 65.250 ;
        RECT 107.390 65.210 108.015 70.230 ;
        RECT 109.340 67.165 110.010 72.480 ;
        RECT 109.780 67.070 110.010 67.165 ;
        RECT 110.220 73.000 110.450 73.070 ;
        RECT 110.220 72.950 111.120 73.000 ;
        RECT 112.195 72.950 112.785 73.210 ;
        RECT 110.220 71.135 112.785 72.950 ;
        RECT 110.220 69.565 111.120 71.135 ;
        RECT 112.195 71.105 112.785 71.135 ;
        RECT 114.015 73.070 114.605 73.210 ;
        RECT 115.835 73.070 116.425 73.210 ;
        RECT 114.015 71.255 116.425 73.070 ;
        RECT 117.445 72.950 117.905 73.685 ;
        RECT 118.360 73.210 118.675 73.500 ;
        RECT 118.360 73.200 118.650 73.210 ;
        RECT 120.525 73.010 121.115 73.210 ;
        RECT 118.675 72.995 121.115 73.010 ;
        RECT 118.170 72.950 118.400 72.995 ;
        RECT 117.445 72.460 118.400 72.950 ;
        RECT 114.015 71.105 114.605 71.255 ;
        RECT 115.835 71.105 116.425 71.255 ;
        RECT 112.195 70.270 112.785 70.525 ;
        RECT 114.015 70.270 114.605 70.525 ;
        RECT 115.835 70.455 116.425 70.525 ;
        RECT 110.220 67.165 111.245 69.565 ;
        RECT 112.195 68.455 114.605 70.270 ;
        RECT 112.195 68.420 112.785 68.455 ;
        RECT 114.015 68.420 114.605 68.455 ;
        RECT 110.220 67.070 110.450 67.165 ;
        RECT 109.970 66.635 110.260 66.865 ;
        RECT 109.980 66.375 110.230 66.635 ;
        RECT 109.695 65.375 110.695 66.375 ;
        RECT 107.390 65.110 107.980 65.210 ;
        RECT 109.980 65.035 110.230 65.375 ;
        RECT 109.945 64.805 110.235 65.035 ;
        RECT 109.755 64.565 109.985 64.645 ;
        RECT 101.775 62.710 102.860 64.530 ;
        RECT 103.750 64.380 104.340 64.530 ;
        RECT 101.775 62.625 102.005 62.710 ;
        RECT 101.525 62.445 101.815 62.465 ;
        RECT 101.525 62.235 101.880 62.445 ;
        RECT 103.740 62.425 104.340 64.380 ;
        RECT 105.570 64.285 106.160 64.530 ;
        RECT 107.390 64.285 107.980 64.530 ;
        RECT 105.570 62.470 107.980 64.285 ;
        RECT 109.320 64.080 109.985 64.565 ;
        RECT 109.000 64.030 109.985 64.080 ;
        RECT 105.570 62.425 106.160 62.470 ;
        RECT 107.390 62.425 107.980 62.470 ;
        RECT 108.850 62.695 109.985 64.030 ;
        RECT 103.740 62.390 104.285 62.425 ;
        RECT 101.565 62.155 101.880 62.235 ;
        RECT 108.850 61.960 109.460 62.695 ;
        RECT 109.755 62.645 109.985 62.695 ;
        RECT 110.195 64.555 110.425 64.645 ;
        RECT 110.870 64.555 111.245 67.165 ;
        RECT 112.195 66.965 112.785 67.230 ;
        RECT 114.015 66.965 114.605 67.230 ;
        RECT 112.195 65.150 114.605 66.965 ;
        RECT 112.195 65.125 112.785 65.150 ;
        RECT 114.015 65.125 114.605 65.150 ;
        RECT 115.815 65.135 116.435 70.455 ;
        RECT 117.815 67.075 118.400 72.460 ;
        RECT 118.170 66.995 118.400 67.075 ;
        RECT 118.610 71.195 121.115 72.995 ;
        RECT 118.610 69.500 119.500 71.195 ;
        RECT 120.525 71.105 121.115 71.195 ;
        RECT 122.345 73.050 122.935 73.210 ;
        RECT 124.165 73.050 124.755 73.210 ;
        RECT 122.345 71.235 124.755 73.050 ;
        RECT 125.900 73.000 126.360 73.685 ;
        RECT 126.675 73.245 126.990 73.535 ;
        RECT 126.690 73.225 126.980 73.245 ;
        RECT 126.500 73.000 126.730 73.020 ;
        RECT 125.900 72.180 126.730 73.000 ;
        RECT 122.345 71.105 122.935 71.235 ;
        RECT 124.165 71.105 124.755 71.235 ;
        RECT 120.525 70.310 121.115 70.525 ;
        RECT 122.345 70.310 122.935 70.525 ;
        RECT 118.610 67.065 119.725 69.500 ;
        RECT 120.525 68.495 122.935 70.310 ;
        RECT 124.165 70.230 124.755 70.525 ;
        RECT 120.525 68.420 121.115 68.495 ;
        RECT 122.345 68.420 122.935 68.495 ;
        RECT 118.610 66.995 118.840 67.065 ;
        RECT 118.355 66.790 118.605 66.800 ;
        RECT 118.355 66.560 118.650 66.790 ;
        RECT 118.355 66.335 118.605 66.560 ;
        RECT 118.140 65.335 119.140 66.335 ;
        RECT 115.835 65.125 116.425 65.135 ;
        RECT 118.355 65.015 118.605 65.335 ;
        RECT 118.295 64.815 118.605 65.015 ;
        RECT 118.295 64.785 118.585 64.815 ;
        RECT 110.195 62.735 111.245 64.555 ;
        RECT 118.105 64.545 118.335 64.625 ;
        RECT 110.195 62.645 110.425 62.735 ;
        RECT 109.945 62.470 110.235 62.485 ;
        RECT 109.930 62.180 110.245 62.470 ;
        RECT 112.195 62.425 112.785 64.545 ;
        RECT 114.015 64.305 114.605 64.545 ;
        RECT 115.835 64.305 116.425 64.545 ;
        RECT 114.015 62.490 116.425 64.305 ;
        RECT 117.685 64.090 118.335 64.545 ;
        RECT 114.015 62.440 114.605 62.490 ;
        RECT 115.835 62.440 116.425 62.490 ;
        RECT 117.245 62.645 118.335 64.090 ;
        RECT 108.005 61.920 109.460 61.960 ;
        RECT 117.245 61.920 117.705 62.645 ;
        RECT 118.105 62.625 118.335 62.645 ;
        RECT 118.545 64.505 118.775 64.625 ;
        RECT 119.350 64.505 119.725 67.065 ;
        RECT 120.525 67.045 121.115 67.230 ;
        RECT 122.345 67.045 122.935 67.230 ;
        RECT 120.525 65.230 122.935 67.045 ;
        RECT 120.525 65.125 121.115 65.230 ;
        RECT 122.345 65.125 122.935 65.230 ;
        RECT 124.140 65.210 124.765 70.230 ;
        RECT 126.070 67.125 126.730 72.180 ;
        RECT 126.500 67.020 126.730 67.125 ;
        RECT 126.940 72.935 127.170 73.020 ;
        RECT 126.940 72.930 127.860 72.935 ;
        RECT 128.855 72.930 129.445 73.210 ;
        RECT 126.940 71.115 129.445 72.930 ;
        RECT 126.940 69.525 127.860 71.115 ;
        RECT 128.855 71.105 129.445 71.115 ;
        RECT 130.675 73.030 131.265 73.210 ;
        RECT 132.495 73.030 133.085 73.210 ;
        RECT 130.675 71.215 133.085 73.030 ;
        RECT 134.140 72.960 134.600 73.685 ;
        RECT 134.980 73.220 135.295 73.510 ;
        RECT 134.795 72.960 135.025 73.035 ;
        RECT 134.140 72.230 135.025 72.960 ;
        RECT 130.675 71.105 131.265 71.215 ;
        RECT 132.495 71.105 133.085 71.215 ;
        RECT 128.855 70.270 129.445 70.525 ;
        RECT 130.675 70.270 131.265 70.525 ;
        RECT 132.495 70.270 133.085 70.525 ;
        RECT 126.940 67.100 128.055 69.525 ;
        RECT 128.855 68.455 131.275 70.270 ;
        RECT 128.855 68.420 129.445 68.455 ;
        RECT 130.675 68.420 131.265 68.455 ;
        RECT 126.940 67.020 127.170 67.100 ;
        RECT 126.690 66.585 126.980 66.815 ;
        RECT 126.690 66.320 126.940 66.585 ;
        RECT 126.410 65.320 127.410 66.320 ;
        RECT 124.165 65.125 124.755 65.210 ;
        RECT 126.690 65.010 126.940 65.320 ;
        RECT 126.680 64.780 126.970 65.010 ;
        RECT 126.490 64.565 126.720 64.620 ;
        RECT 118.545 62.715 119.725 64.505 ;
        RECT 120.525 64.530 121.115 64.545 ;
        RECT 118.545 62.685 119.610 62.715 ;
        RECT 118.545 62.625 118.775 62.685 ;
        RECT 120.525 62.510 121.120 64.530 ;
        RECT 122.345 64.325 122.935 64.545 ;
        RECT 124.165 64.325 124.755 64.545 ;
        RECT 122.345 62.510 124.755 64.325 ;
        RECT 126.090 64.100 126.720 64.565 ;
        RECT 118.285 62.190 118.600 62.480 ;
        RECT 120.525 62.440 121.115 62.510 ;
        RECT 122.345 62.440 122.935 62.510 ;
        RECT 123.155 62.425 123.745 62.510 ;
        RECT 124.165 62.440 124.755 62.510 ;
        RECT 125.680 62.665 126.720 64.100 ;
        RECT 125.680 61.920 126.140 62.665 ;
        RECT 126.490 62.620 126.720 62.665 ;
        RECT 126.930 64.495 127.160 64.620 ;
        RECT 127.680 64.495 128.055 67.100 ;
        RECT 128.855 67.025 129.445 67.230 ;
        RECT 130.675 67.025 131.265 67.230 ;
        RECT 128.855 65.210 131.265 67.025 ;
        RECT 132.460 65.250 133.085 70.270 ;
        RECT 134.350 67.085 135.025 72.230 ;
        RECT 134.795 67.035 135.025 67.085 ;
        RECT 135.235 72.930 135.465 73.035 ;
        RECT 137.160 72.930 137.750 73.205 ;
        RECT 135.235 71.115 137.750 72.930 ;
        RECT 135.235 69.625 136.140 71.115 ;
        RECT 137.160 71.100 137.750 71.115 ;
        RECT 138.980 73.030 139.570 73.205 ;
        RECT 140.800 73.030 141.390 73.205 ;
        RECT 138.980 71.215 141.390 73.030 ;
        RECT 142.415 72.960 142.875 73.685 ;
        RECT 143.295 73.450 143.610 73.525 ;
        RECT 143.285 73.235 143.610 73.450 ;
        RECT 143.285 73.220 143.575 73.235 ;
        RECT 145.460 73.030 146.050 73.215 ;
        RECT 147.280 73.030 147.870 73.215 ;
        RECT 143.095 72.960 143.325 73.015 ;
        RECT 142.415 72.000 143.325 72.960 ;
        RECT 138.980 71.100 139.570 71.215 ;
        RECT 140.800 71.100 141.390 71.215 ;
        RECT 137.160 70.270 137.750 70.520 ;
        RECT 138.980 70.270 139.570 70.520 ;
        RECT 135.235 67.075 136.275 69.625 ;
        RECT 137.160 68.455 139.570 70.270 ;
        RECT 137.160 68.415 137.750 68.455 ;
        RECT 138.980 68.415 139.570 68.455 ;
        RECT 140.800 70.250 141.390 70.520 ;
        RECT 140.800 68.415 141.450 70.250 ;
        RECT 140.825 67.225 141.450 68.415 ;
        RECT 135.235 67.035 135.465 67.075 ;
        RECT 134.940 66.350 135.285 66.840 ;
        RECT 134.715 65.350 135.715 66.350 ;
        RECT 128.855 65.125 129.445 65.210 ;
        RECT 130.675 65.125 131.265 65.210 ;
        RECT 132.495 65.125 133.085 65.250 ;
        RECT 134.940 65.020 135.285 65.350 ;
        RECT 134.920 64.805 135.285 65.020 ;
        RECT 134.920 64.790 135.210 64.805 ;
        RECT 134.730 64.555 134.960 64.630 ;
        RECT 126.930 62.740 128.055 64.495 ;
        RECT 128.855 64.450 129.445 64.545 ;
        RECT 126.930 62.675 127.970 62.740 ;
        RECT 126.930 62.620 127.160 62.675 ;
        RECT 126.680 62.445 126.970 62.460 ;
        RECT 126.680 62.230 127.020 62.445 ;
        RECT 128.840 62.440 129.445 64.450 ;
        RECT 130.675 64.325 131.265 64.545 ;
        RECT 132.495 64.325 133.085 64.545 ;
        RECT 130.650 62.510 133.085 64.325 ;
        RECT 134.400 64.060 134.960 64.555 ;
        RECT 130.675 62.440 131.265 62.510 ;
        RECT 132.495 62.440 133.085 62.510 ;
        RECT 133.970 62.655 134.960 64.060 ;
        RECT 128.840 62.420 129.385 62.440 ;
        RECT 126.705 62.155 127.020 62.230 ;
        RECT 133.970 61.920 134.430 62.655 ;
        RECT 134.730 62.630 134.960 62.655 ;
        RECT 135.170 64.530 135.400 64.630 ;
        RECT 135.900 64.530 136.275 67.075 ;
        RECT 137.160 67.025 137.750 67.225 ;
        RECT 138.980 67.025 139.570 67.225 ;
        RECT 137.160 65.210 139.570 67.025 ;
        RECT 137.160 65.120 137.750 65.210 ;
        RECT 138.980 65.120 139.570 65.210 ;
        RECT 140.800 65.230 141.450 67.225 ;
        RECT 142.665 67.085 143.325 72.000 ;
        RECT 143.095 67.015 143.325 67.085 ;
        RECT 143.535 72.995 143.765 73.015 ;
        RECT 143.535 70.410 144.320 72.995 ;
        RECT 145.460 71.215 147.870 73.030 ;
        RECT 145.460 71.110 146.050 71.215 ;
        RECT 147.280 71.110 147.870 71.215 ;
        RECT 145.460 70.410 146.050 70.530 ;
        RECT 143.535 68.595 146.050 70.410 ;
        RECT 147.280 70.290 147.870 70.530 ;
        RECT 143.535 67.830 144.320 68.595 ;
        RECT 145.460 68.425 146.050 68.595 ;
        RECT 147.215 68.425 147.870 70.290 ;
        RECT 143.535 67.095 144.360 67.830 ;
        RECT 143.535 67.015 143.765 67.095 ;
        RECT 143.285 66.755 143.575 66.810 ;
        RECT 143.285 66.745 143.800 66.755 ;
        RECT 143.255 66.310 143.800 66.745 ;
        RECT 144.030 66.515 144.360 67.095 ;
        RECT 145.280 66.945 146.280 67.945 ;
        RECT 147.215 67.235 147.840 68.425 ;
        RECT 142.805 65.310 143.805 66.310 ;
        RECT 144.100 65.515 144.360 66.515 ;
        RECT 140.800 65.120 141.390 65.230 ;
        RECT 143.255 64.845 143.800 65.310 ;
        RECT 144.075 65.220 144.360 65.515 ;
        RECT 145.390 65.260 146.105 66.945 ;
        RECT 147.215 65.270 147.870 67.235 ;
        RECT 143.255 64.835 143.730 64.845 ;
        RECT 143.285 64.820 143.730 64.835 ;
        RECT 143.285 64.790 143.575 64.820 ;
        RECT 143.095 64.585 143.325 64.630 ;
        RECT 135.170 62.840 136.275 64.530 ;
        RECT 137.160 64.430 137.750 64.540 ;
        RECT 135.170 62.710 136.235 62.840 ;
        RECT 135.170 62.630 135.400 62.710 ;
        RECT 134.980 62.470 135.295 62.480 ;
        RECT 134.920 62.240 135.295 62.470 ;
        RECT 137.145 62.435 137.750 64.430 ;
        RECT 138.980 64.385 139.570 64.540 ;
        RECT 140.800 64.385 141.390 64.540 ;
        RECT 138.980 62.570 141.390 64.385 ;
        RECT 142.745 64.150 143.325 64.585 ;
        RECT 138.980 62.435 139.570 62.570 ;
        RECT 137.145 62.410 137.690 62.435 ;
        RECT 139.915 62.420 140.460 62.570 ;
        RECT 140.800 62.435 141.390 62.570 ;
        RECT 142.325 62.685 143.325 64.150 ;
        RECT 134.980 62.190 135.295 62.240 ;
        RECT 142.325 61.920 142.785 62.685 ;
        RECT 143.095 62.630 143.325 62.685 ;
        RECT 143.535 64.570 143.765 64.630 ;
        RECT 144.030 64.570 144.360 65.220 ;
        RECT 145.460 65.225 146.065 65.260 ;
        RECT 145.460 65.130 146.050 65.225 ;
        RECT 147.280 65.130 147.870 65.270 ;
        RECT 143.535 63.075 144.360 64.570 ;
        RECT 145.460 64.365 146.050 64.550 ;
        RECT 147.280 64.365 147.870 64.550 ;
        RECT 143.535 62.690 144.135 63.075 ;
        RECT 143.535 62.630 143.765 62.690 ;
        RECT 145.460 62.550 147.870 64.365 ;
        RECT 143.260 62.180 143.575 62.470 ;
        RECT 145.460 62.445 146.050 62.550 ;
        RECT 147.280 62.445 147.870 62.550 ;
        RECT 79.960 61.440 148.575 61.920 ;
        RECT 79.950 60.860 148.580 61.440 ;
        RECT 11.390 57.310 14.350 57.410 ;
        RECT 2.570 57.280 4.675 57.310 ;
        RECT 2.510 56.720 4.675 57.280 ;
        RECT 5.255 57.280 7.360 57.310 ;
        RECT 8.550 57.280 10.655 57.310 ;
        RECT 5.255 56.720 10.655 57.280 ;
        RECT 11.235 56.720 14.350 57.310 ;
        RECT 2.510 55.490 4.410 56.720 ;
        RECT 5.310 56.680 10.610 56.720 ;
        RECT 11.390 56.630 14.350 56.720 ;
        RECT 2.510 54.900 4.675 55.490 ;
        RECT 5.255 55.480 7.360 55.490 ;
        RECT 8.550 55.480 10.655 55.490 ;
        RECT 5.255 54.900 10.655 55.480 ;
        RECT 11.235 54.900 13.340 55.490 ;
        RECT 2.510 54.880 4.410 54.900 ;
        RECT 5.310 54.880 10.610 54.900 ;
        RECT 2.710 53.670 4.610 53.680 ;
        RECT 5.310 53.670 10.610 53.680 ;
        RECT 11.310 53.670 13.210 54.900 ;
        RECT 2.570 53.080 4.675 53.670 ;
        RECT 5.255 53.080 10.655 53.670 ;
        RECT 11.235 53.080 13.340 53.670 ;
        RECT 2.710 51.850 4.610 53.080 ;
        RECT 61.840 52.540 62.050 52.570 ;
        RECT 61.840 52.090 68.090 52.540 ;
        RECT 61.840 52.060 62.050 52.090 ;
        RECT 11.310 51.875 13.635 51.880 ;
        RECT 11.310 51.850 16.600 51.875 ;
        RECT 26.165 51.850 26.540 51.945 ;
        RECT 41.485 51.875 46.610 51.880 ;
        RECT 29.240 51.850 46.610 51.875 ;
        RECT 47.310 51.850 52.610 51.980 ;
        RECT 53.310 51.850 58.610 51.880 ;
        RECT 59.310 51.850 70.710 51.880 ;
        RECT 71.310 51.850 76.610 51.880 ;
        RECT 77.310 51.850 82.610 51.880 ;
        RECT 2.570 51.260 4.675 51.850 ;
        RECT 5.255 51.780 7.360 51.850 ;
        RECT 8.550 51.780 10.655 51.850 ;
        RECT 5.255 51.260 10.655 51.780 ;
        RECT 11.235 51.260 16.635 51.850 ;
        RECT 17.215 51.260 22.615 51.850 ;
        RECT 23.195 51.810 25.300 51.850 ;
        RECT 26.165 51.810 28.595 51.850 ;
        RECT 23.195 51.260 28.595 51.810 ;
        RECT 29.175 51.270 46.695 51.850 ;
        RECT 29.175 51.260 31.280 51.270 ;
        RECT 41.485 51.260 46.695 51.270 ;
        RECT 47.275 51.280 52.675 51.850 ;
        RECT 47.275 51.260 49.380 51.280 ;
        RECT 50.570 51.260 52.675 51.280 ;
        RECT 53.255 51.260 58.655 51.850 ;
        RECT 59.235 51.260 70.710 51.850 ;
        RECT 71.275 51.260 76.675 51.850 ;
        RECT 77.255 51.280 82.655 51.850 ;
        RECT 77.255 51.260 79.360 51.280 ;
        RECT 80.550 51.260 82.655 51.280 ;
        RECT 83.235 51.260 85.340 51.850 ;
        RECT 5.310 51.180 10.610 51.260 ;
        RECT 11.310 51.180 16.600 51.260 ;
        RECT 17.260 51.255 22.580 51.260 ;
        RECT 13.140 51.170 16.600 51.180 ;
        RECT 1.980 50.360 10.405 50.855 ;
        RECT 10.940 50.500 11.445 50.595 ;
        RECT 17.450 50.500 17.705 51.255 ;
        RECT 23.230 51.215 28.550 51.260 ;
        RECT 29.275 50.575 29.680 51.260 ;
        RECT 41.485 51.180 46.610 51.260 ;
        RECT 47.555 50.630 47.930 51.260 ;
        RECT 53.310 51.180 58.610 51.260 ;
        RECT 59.310 51.180 70.710 51.260 ;
        RECT 71.310 51.180 76.610 51.260 ;
        RECT 59.485 50.680 59.890 51.180 ;
        RECT 10.940 50.245 17.705 50.500 ;
        RECT 10.940 50.150 11.445 50.245 ;
        RECT 26.985 50.170 29.680 50.575 ;
        RECT 38.975 50.255 47.930 50.630 ;
        RECT 55.085 50.275 59.890 50.680 ;
        RECT 71.435 50.655 71.785 51.180 ;
        RECT 82.200 50.735 82.540 51.260 ;
        RECT 83.390 51.160 85.330 51.260 ;
        RECT 83.550 50.755 83.945 51.160 ;
        RECT 66.985 50.305 71.785 50.655 ;
        RECT 78.210 50.170 80.780 50.690 ;
        RECT 82.170 50.395 82.570 50.735 ;
        RECT 83.130 50.360 83.945 50.755 ;
        RECT 84.890 51.100 85.330 51.160 ;
        RECT 144.610 51.100 146.610 51.180 ;
        RECT 84.890 50.660 146.610 51.100 ;
        RECT 27.910 49.960 30.610 49.980 ;
        RECT 55.810 49.960 58.510 49.980 ;
        RECT 83.910 49.960 86.210 49.980 ;
        RECT 112.010 49.960 114.310 49.980 ;
        RECT 1.870 49.280 140.345 49.960 ;
        RECT 144.610 49.310 146.610 50.660 ;
        RECT 1.870 49.260 28.345 49.280 ;
        RECT 29.870 49.260 56.345 49.280 ;
        RECT 57.870 49.260 84.345 49.280 ;
        RECT 85.870 49.260 112.345 49.280 ;
        RECT 113.870 49.260 140.345 49.280 ;
        RECT 2.840 48.635 4.750 49.260 ;
        RECT 6.840 48.925 8.725 48.930 ;
        RECT 10.285 48.925 12.170 48.930 ;
        RECT 6.830 48.695 8.790 48.925 ;
        RECT 10.260 48.695 12.220 48.925 ;
        RECT 2.805 48.405 4.805 48.635 ;
        RECT 6.550 48.410 6.780 48.490 ;
        RECT 2.010 48.355 2.505 48.375 ;
        RECT 2.010 45.060 2.600 48.355 ;
        RECT 5.010 48.275 5.240 48.355 ;
        RECT 4.980 45.060 5.240 48.275 ;
        RECT 2.010 43.245 5.240 45.060 ;
        RECT 2.010 40.395 2.600 43.245 ;
        RECT 3.495 40.640 3.755 40.960 ;
        RECT 4.980 40.645 5.240 43.245 ;
        RECT 6.310 40.990 6.780 48.410 ;
        RECT 7.270 41.775 8.160 48.695 ;
        RECT 8.840 48.390 9.070 48.490 ;
        RECT 8.840 48.380 9.195 48.390 ;
        RECT 9.980 48.380 10.210 48.490 ;
        RECT 3.550 40.480 3.700 40.640 ;
        RECT 2.010 35.255 2.505 40.395 ;
        RECT 3.525 40.345 3.730 40.480 ;
        RECT 5.010 40.395 5.240 40.645 ;
        RECT 6.030 40.550 6.780 40.990 ;
        RECT 7.200 40.775 8.215 41.775 ;
        RECT 2.805 40.115 4.805 40.345 ;
        RECT 6.030 38.355 6.400 40.550 ;
        RECT 6.550 40.490 6.780 40.550 ;
        RECT 7.270 40.285 8.160 40.775 ;
        RECT 8.840 40.580 10.210 48.380 ;
        RECT 10.745 43.635 11.635 48.695 ;
        RECT 12.270 48.410 12.500 48.490 ;
        RECT 10.740 42.015 11.640 43.635 ;
        RECT 10.745 41.605 11.635 42.015 ;
        RECT 10.670 40.605 11.700 41.605 ;
        RECT 12.270 40.625 12.645 48.410 ;
        RECT 12.920 48.025 14.600 49.260 ;
        RECT 15.435 48.025 20.360 48.035 ;
        RECT 12.920 47.545 20.360 48.025 ;
        RECT 12.920 45.285 14.600 47.545 ;
        RECT 15.435 47.125 20.360 47.545 ;
        RECT 14.940 46.935 15.195 46.960 ;
        RECT 14.940 46.920 15.215 46.935 ;
        RECT 14.910 46.645 15.245 46.920 ;
        RECT 15.420 46.895 20.420 47.125 ;
        RECT 20.630 46.935 20.885 46.960 ;
        RECT 14.940 46.630 15.195 46.645 ;
        RECT 15.420 46.455 20.420 46.685 ;
        RECT 20.625 46.645 20.885 46.935 ;
        RECT 20.630 46.630 20.885 46.645 ;
        RECT 15.465 46.445 20.320 46.455 ;
        RECT 15.465 44.920 18.110 44.925 ;
        RECT 14.140 44.720 18.110 44.920 ;
        RECT 14.140 44.690 18.100 44.720 ;
        RECT 12.980 44.335 13.315 44.610 ;
        RECT 13.860 44.440 14.090 44.485 ;
        RECT 8.840 40.560 9.195 40.580 ;
        RECT 8.840 40.490 9.070 40.560 ;
        RECT 9.980 40.490 10.210 40.580 ;
        RECT 10.740 40.465 11.650 40.605 ;
        RECT 12.270 40.490 12.660 40.625 ;
        RECT 10.730 40.285 11.740 40.465 ;
        RECT 6.830 40.055 8.790 40.285 ;
        RECT 10.260 40.055 12.220 40.285 ;
        RECT 7.555 39.065 7.885 40.055 ;
        RECT 10.285 40.050 12.170 40.055 ;
        RECT 12.465 38.355 12.660 40.490 ;
        RECT 13.050 38.830 13.240 44.335 ;
        RECT 13.670 43.105 14.090 44.440 ;
        RECT 15.395 43.105 16.740 44.690 ;
        RECT 13.670 41.720 16.740 43.105 ;
        RECT 13.670 40.990 14.090 41.720 ;
        RECT 13.665 40.485 14.090 40.990 ;
        RECT 13.050 38.640 13.365 38.830 ;
        RECT 3.370 38.125 7.330 38.355 ;
        RECT 8.800 38.125 12.760 38.355 ;
        RECT 13.175 38.130 13.365 38.640 ;
        RECT 3.090 37.515 3.320 37.965 ;
        RECT 4.570 37.515 5.360 38.125 ;
        RECT 3.090 37.210 5.360 37.515 ;
        RECT 3.035 37.195 5.360 37.210 ;
        RECT 2.950 36.350 5.360 37.195 ;
        RECT 2.950 35.975 3.320 36.350 ;
        RECT 3.090 35.965 3.320 35.975 ;
        RECT 4.570 35.805 5.360 36.350 ;
        RECT 7.380 37.880 7.610 37.965 ;
        RECT 8.520 37.880 8.750 37.965 ;
        RECT 7.380 36.055 8.750 37.880 ;
        RECT 7.380 35.965 7.610 36.055 ;
        RECT 3.370 35.575 7.330 35.805 ;
        RECT 2.950 35.255 3.175 35.265 ;
        RECT 7.850 35.255 8.340 36.055 ;
        RECT 8.520 35.965 8.750 36.055 ;
        RECT 10.235 37.745 11.575 38.125 ;
        RECT 12.810 37.745 13.040 37.965 ;
        RECT 10.235 36.150 13.040 37.745 ;
        RECT 10.235 35.805 11.575 36.150 ;
        RECT 12.810 35.965 13.040 36.150 ;
        RECT 8.800 35.575 12.760 35.805 ;
        RECT 13.190 35.785 13.365 38.130 ;
        RECT 13.665 37.965 13.960 40.485 ;
        RECT 15.395 40.280 16.740 41.720 ;
        RECT 18.150 44.390 18.380 44.485 ;
        RECT 18.625 44.390 19.115 46.445 ;
        RECT 19.685 44.920 20.320 44.925 ;
        RECT 19.570 44.690 23.530 44.920 ;
        RECT 19.290 44.390 19.520 44.485 ;
        RECT 18.150 40.565 19.520 44.390 ;
        RECT 18.150 40.485 18.380 40.565 ;
        RECT 19.290 40.485 19.520 40.565 ;
        RECT 20.945 40.280 22.290 44.690 ;
        RECT 23.580 44.420 23.810 44.485 ;
        RECT 24.465 44.425 24.940 49.260 ;
        RECT 26.265 48.455 26.945 49.260 ;
        RECT 27.365 48.735 27.700 48.985 ;
        RECT 27.380 48.710 27.670 48.735 ;
        RECT 30.840 48.635 32.750 49.260 ;
        RECT 34.840 48.925 36.725 48.930 ;
        RECT 38.285 48.925 40.170 48.930 ;
        RECT 34.830 48.695 36.790 48.925 ;
        RECT 38.260 48.695 40.220 48.925 ;
        RECT 27.190 48.455 27.420 48.505 ;
        RECT 26.265 47.955 27.420 48.455 ;
        RECT 25.335 44.735 25.670 44.985 ;
        RECT 25.355 44.705 25.645 44.735 ;
        RECT 25.165 44.425 25.395 44.500 ;
        RECT 23.580 40.485 24.035 44.420 ;
        RECT 24.465 43.680 25.395 44.425 ;
        RECT 24.800 40.565 25.395 43.680 ;
        RECT 25.165 40.500 25.395 40.565 ;
        RECT 25.605 44.475 25.835 44.500 ;
        RECT 25.605 40.920 26.115 44.475 ;
        RECT 25.605 40.550 26.300 40.920 ;
        RECT 26.800 40.600 27.420 47.955 ;
        RECT 25.605 40.500 25.835 40.550 ;
        RECT 14.140 40.250 18.100 40.280 ;
        RECT 19.570 40.250 23.530 40.280 ;
        RECT 14.140 40.090 23.530 40.250 ;
        RECT 14.140 40.050 18.100 40.090 ;
        RECT 19.570 40.050 23.530 40.090 ;
        RECT 23.695 38.660 24.035 40.485 ;
        RECT 25.345 38.660 25.765 40.305 ;
        RECT 23.695 38.505 25.765 38.660 ;
        RECT 23.770 38.390 25.765 38.505 ;
        RECT 14.230 38.125 18.190 38.355 ;
        RECT 19.660 38.125 23.620 38.355 ;
        RECT 13.665 37.205 14.180 37.965 ;
        RECT 13.735 36.025 14.180 37.205 ;
        RECT 13.950 35.965 14.180 36.025 ;
        RECT 15.610 35.805 16.565 38.125 ;
        RECT 18.240 37.900 18.470 37.965 ;
        RECT 19.380 37.900 19.610 37.965 ;
        RECT 18.240 36.030 19.610 37.900 ;
        RECT 18.240 35.965 18.470 36.030 ;
        RECT 13.175 35.255 13.365 35.785 ;
        RECT 14.230 35.575 18.190 35.805 ;
        RECT 18.645 35.255 19.200 36.030 ;
        RECT 19.380 35.965 19.610 36.030 ;
        RECT 21.055 35.805 22.010 38.125 ;
        RECT 23.770 37.970 24.035 38.390 ;
        RECT 25.345 38.115 25.765 38.390 ;
        RECT 26.000 39.355 26.300 40.550 ;
        RECT 27.190 40.505 27.420 40.600 ;
        RECT 27.630 48.430 27.860 48.505 ;
        RECT 27.630 41.110 28.405 48.430 ;
        RECT 30.805 48.405 32.805 48.635 ;
        RECT 34.550 48.410 34.780 48.490 ;
        RECT 30.370 45.060 30.600 48.355 ;
        RECT 33.010 48.275 33.240 48.355 ;
        RECT 32.980 45.060 33.240 48.275 ;
        RECT 30.370 43.245 33.240 45.060 ;
        RECT 27.630 40.580 28.480 41.110 ;
        RECT 30.370 40.825 30.600 43.245 ;
        RECT 27.630 40.505 27.860 40.580 ;
        RECT 27.295 39.825 27.810 40.315 ;
        RECT 28.110 39.825 28.480 40.580 ;
        RECT 30.010 40.395 30.600 40.825 ;
        RECT 31.495 40.640 31.755 40.960 ;
        RECT 32.980 40.645 33.240 43.245 ;
        RECT 34.310 40.990 34.780 48.410 ;
        RECT 35.270 41.775 36.160 48.695 ;
        RECT 36.840 48.390 37.070 48.490 ;
        RECT 36.840 48.380 37.195 48.390 ;
        RECT 37.980 48.380 38.210 48.490 ;
        RECT 31.550 40.480 31.700 40.640 ;
        RECT 27.295 39.360 27.805 39.825 ;
        RECT 26.930 39.355 27.805 39.360 ;
        RECT 26.000 38.950 27.805 39.355 ;
        RECT 26.000 38.110 26.300 38.950 ;
        RECT 26.930 38.935 27.805 38.950 ;
        RECT 27.295 38.825 27.805 38.935 ;
        RECT 27.295 38.125 27.810 38.825 ;
        RECT 28.035 38.795 29.035 39.825 ;
        RECT 23.695 37.965 24.035 37.970 ;
        RECT 23.670 36.020 24.035 37.965 ;
        RECT 25.250 37.900 25.480 37.970 ;
        RECT 24.755 37.230 25.480 37.900 ;
        RECT 24.745 37.040 25.480 37.230 ;
        RECT 24.745 36.240 25.100 37.040 ;
        RECT 25.250 36.970 25.480 37.040 ;
        RECT 25.690 37.925 25.920 37.970 ;
        RECT 26.060 37.925 26.300 38.110 ;
        RECT 25.690 37.595 26.300 37.925 ;
        RECT 27.275 37.870 27.505 37.975 ;
        RECT 25.690 37.040 26.185 37.595 ;
        RECT 25.690 36.970 25.920 37.040 ;
        RECT 25.440 36.785 25.730 36.810 ;
        RECT 25.425 36.535 25.760 36.785 ;
        RECT 27.045 36.765 27.505 37.870 ;
        RECT 26.725 36.240 27.505 36.765 ;
        RECT 24.305 36.060 27.505 36.240 ;
        RECT 23.670 35.965 23.900 36.020 ;
        RECT 19.660 35.575 23.620 35.805 ;
        RECT 24.305 35.620 27.110 36.060 ;
        RECT 27.275 35.975 27.505 36.060 ;
        RECT 27.715 37.910 27.945 37.975 ;
        RECT 28.110 37.910 28.480 38.795 ;
        RECT 27.715 37.585 28.480 37.910 ;
        RECT 27.715 36.045 28.475 37.585 ;
        RECT 27.715 35.975 27.945 36.045 ;
        RECT 27.465 35.795 27.755 35.815 ;
        RECT 24.305 35.255 26.770 35.620 ;
        RECT 27.440 35.545 27.775 35.795 ;
        RECT 30.010 35.280 30.505 40.395 ;
        RECT 31.525 40.345 31.730 40.480 ;
        RECT 33.010 40.395 33.240 40.645 ;
        RECT 34.030 40.550 34.780 40.990 ;
        RECT 35.200 40.775 36.215 41.775 ;
        RECT 30.805 40.115 32.805 40.345 ;
        RECT 34.030 38.355 34.400 40.550 ;
        RECT 34.550 40.490 34.780 40.550 ;
        RECT 35.270 40.285 36.160 40.775 ;
        RECT 36.840 40.580 38.210 48.380 ;
        RECT 38.745 43.635 39.635 48.695 ;
        RECT 40.270 48.410 40.500 48.490 ;
        RECT 38.740 42.015 39.640 43.635 ;
        RECT 38.745 41.605 39.635 42.015 ;
        RECT 38.670 40.605 39.700 41.605 ;
        RECT 40.270 40.625 40.645 48.410 ;
        RECT 40.920 48.025 42.600 49.260 ;
        RECT 43.435 48.025 48.360 48.035 ;
        RECT 40.920 47.545 48.360 48.025 ;
        RECT 40.920 45.285 42.600 47.545 ;
        RECT 43.435 47.125 48.360 47.545 ;
        RECT 42.940 46.935 43.195 46.960 ;
        RECT 42.940 46.920 43.215 46.935 ;
        RECT 42.910 46.645 43.245 46.920 ;
        RECT 43.420 46.895 48.420 47.125 ;
        RECT 48.630 46.935 48.885 46.960 ;
        RECT 42.940 46.630 43.195 46.645 ;
        RECT 43.420 46.455 48.420 46.685 ;
        RECT 48.625 46.645 48.885 46.935 ;
        RECT 48.630 46.630 48.885 46.645 ;
        RECT 43.465 46.445 48.320 46.455 ;
        RECT 43.465 44.920 46.110 44.925 ;
        RECT 42.140 44.720 46.110 44.920 ;
        RECT 42.140 44.690 46.100 44.720 ;
        RECT 40.980 44.335 41.315 44.610 ;
        RECT 41.860 44.440 42.090 44.485 ;
        RECT 36.840 40.560 37.195 40.580 ;
        RECT 36.840 40.490 37.070 40.560 ;
        RECT 37.980 40.490 38.210 40.580 ;
        RECT 38.740 40.465 39.650 40.605 ;
        RECT 40.270 40.490 40.660 40.625 ;
        RECT 38.730 40.285 39.740 40.465 ;
        RECT 34.830 40.055 36.790 40.285 ;
        RECT 38.260 40.055 40.220 40.285 ;
        RECT 35.540 39.340 35.890 40.055 ;
        RECT 38.285 40.050 40.170 40.055 ;
        RECT 40.465 38.355 40.660 40.490 ;
        RECT 41.050 38.830 41.240 44.335 ;
        RECT 41.670 43.105 42.090 44.440 ;
        RECT 43.395 43.105 44.740 44.690 ;
        RECT 41.670 41.720 44.740 43.105 ;
        RECT 41.670 40.990 42.090 41.720 ;
        RECT 41.665 40.485 42.090 40.990 ;
        RECT 41.050 38.640 41.365 38.830 ;
        RECT 31.370 38.125 35.330 38.355 ;
        RECT 36.800 38.125 40.760 38.355 ;
        RECT 41.175 38.130 41.365 38.640 ;
        RECT 31.090 37.515 31.320 37.965 ;
        RECT 32.570 37.515 33.360 38.125 ;
        RECT 31.090 37.210 33.360 37.515 ;
        RECT 31.035 37.195 33.360 37.210 ;
        RECT 30.950 36.350 33.360 37.195 ;
        RECT 30.950 35.975 31.320 36.350 ;
        RECT 31.090 35.965 31.320 35.975 ;
        RECT 32.570 35.805 33.360 36.350 ;
        RECT 35.380 37.880 35.610 37.965 ;
        RECT 36.520 37.880 36.750 37.965 ;
        RECT 35.380 36.055 36.750 37.880 ;
        RECT 35.380 35.965 35.610 36.055 ;
        RECT 31.370 35.575 35.330 35.805 ;
        RECT 28.410 35.255 30.505 35.280 ;
        RECT 30.950 35.255 31.175 35.265 ;
        RECT 35.850 35.255 36.340 36.055 ;
        RECT 36.520 35.965 36.750 36.055 ;
        RECT 38.235 37.745 39.575 38.125 ;
        RECT 40.810 37.745 41.040 37.965 ;
        RECT 38.235 36.150 41.040 37.745 ;
        RECT 38.235 35.805 39.575 36.150 ;
        RECT 40.810 35.965 41.040 36.150 ;
        RECT 36.800 35.575 40.760 35.805 ;
        RECT 41.190 35.785 41.365 38.130 ;
        RECT 41.665 37.965 41.960 40.485 ;
        RECT 43.395 40.280 44.740 41.720 ;
        RECT 46.150 44.390 46.380 44.485 ;
        RECT 46.625 44.390 47.115 46.445 ;
        RECT 47.685 44.920 48.320 44.925 ;
        RECT 47.570 44.690 51.530 44.920 ;
        RECT 47.290 44.390 47.520 44.485 ;
        RECT 46.150 40.565 47.520 44.390 ;
        RECT 46.150 40.485 46.380 40.565 ;
        RECT 47.290 40.485 47.520 40.565 ;
        RECT 48.945 40.280 50.290 44.690 ;
        RECT 51.580 44.420 51.810 44.485 ;
        RECT 52.465 44.425 52.940 49.260 ;
        RECT 54.265 48.455 54.945 49.260 ;
        RECT 55.365 48.735 55.700 48.985 ;
        RECT 55.380 48.710 55.670 48.735 ;
        RECT 58.840 48.635 60.750 49.260 ;
        RECT 62.840 48.925 64.725 48.930 ;
        RECT 66.285 48.925 68.170 48.930 ;
        RECT 62.830 48.695 64.790 48.925 ;
        RECT 66.260 48.695 68.220 48.925 ;
        RECT 55.190 48.455 55.420 48.505 ;
        RECT 54.265 47.955 55.420 48.455 ;
        RECT 53.335 44.735 53.670 44.985 ;
        RECT 53.355 44.705 53.645 44.735 ;
        RECT 53.165 44.425 53.395 44.500 ;
        RECT 51.580 40.485 52.035 44.420 ;
        RECT 52.465 43.680 53.395 44.425 ;
        RECT 52.800 40.565 53.395 43.680 ;
        RECT 53.165 40.500 53.395 40.565 ;
        RECT 53.605 44.475 53.835 44.500 ;
        RECT 53.605 40.920 54.115 44.475 ;
        RECT 53.605 40.550 54.300 40.920 ;
        RECT 54.800 40.600 55.420 47.955 ;
        RECT 53.605 40.500 53.835 40.550 ;
        RECT 42.140 40.250 46.100 40.280 ;
        RECT 47.570 40.250 51.530 40.280 ;
        RECT 42.140 40.090 51.530 40.250 ;
        RECT 42.140 40.050 46.100 40.090 ;
        RECT 47.570 40.050 51.530 40.090 ;
        RECT 51.695 38.660 52.035 40.485 ;
        RECT 53.345 38.660 53.765 40.305 ;
        RECT 51.695 38.505 53.765 38.660 ;
        RECT 51.770 38.390 53.765 38.505 ;
        RECT 42.230 38.125 46.190 38.355 ;
        RECT 47.660 38.125 51.620 38.355 ;
        RECT 41.665 37.205 42.180 37.965 ;
        RECT 41.735 36.025 42.180 37.205 ;
        RECT 41.950 35.965 42.180 36.025 ;
        RECT 43.610 35.805 44.565 38.125 ;
        RECT 46.240 37.900 46.470 37.965 ;
        RECT 47.380 37.900 47.610 37.965 ;
        RECT 46.240 36.030 47.610 37.900 ;
        RECT 46.240 35.965 46.470 36.030 ;
        RECT 41.175 35.255 41.365 35.785 ;
        RECT 42.230 35.575 46.190 35.805 ;
        RECT 46.645 35.255 47.200 36.030 ;
        RECT 47.380 35.965 47.610 36.030 ;
        RECT 49.055 35.805 50.010 38.125 ;
        RECT 51.770 37.970 52.035 38.390 ;
        RECT 53.345 38.115 53.765 38.390 ;
        RECT 54.000 39.355 54.300 40.550 ;
        RECT 55.190 40.505 55.420 40.600 ;
        RECT 55.630 48.430 55.860 48.505 ;
        RECT 55.630 41.110 56.405 48.430 ;
        RECT 58.805 48.405 60.805 48.635 ;
        RECT 62.550 48.410 62.780 48.490 ;
        RECT 58.370 45.060 58.600 48.355 ;
        RECT 61.010 48.275 61.240 48.355 ;
        RECT 60.980 45.060 61.240 48.275 ;
        RECT 58.370 43.245 61.240 45.060 ;
        RECT 55.630 40.580 56.480 41.110 ;
        RECT 58.370 40.825 58.600 43.245 ;
        RECT 55.630 40.505 55.860 40.580 ;
        RECT 55.295 39.825 55.810 40.315 ;
        RECT 55.295 39.360 55.805 39.825 ;
        RECT 56.110 39.795 56.480 40.580 ;
        RECT 58.010 40.395 58.600 40.825 ;
        RECT 59.495 40.640 59.755 40.960 ;
        RECT 60.980 40.645 61.240 43.245 ;
        RECT 62.310 40.990 62.780 48.410 ;
        RECT 63.270 41.775 64.160 48.695 ;
        RECT 64.840 48.390 65.070 48.490 ;
        RECT 64.840 48.380 65.195 48.390 ;
        RECT 65.980 48.380 66.210 48.490 ;
        RECT 59.550 40.480 59.700 40.640 ;
        RECT 54.930 39.355 55.805 39.360 ;
        RECT 54.000 38.950 55.805 39.355 ;
        RECT 54.000 38.110 54.300 38.950 ;
        RECT 54.930 38.935 55.805 38.950 ;
        RECT 55.295 38.825 55.805 38.935 ;
        RECT 55.295 38.125 55.810 38.825 ;
        RECT 56.005 38.795 57.035 39.795 ;
        RECT 51.695 37.965 52.035 37.970 ;
        RECT 51.670 36.020 52.035 37.965 ;
        RECT 53.250 37.900 53.480 37.970 ;
        RECT 52.755 37.230 53.480 37.900 ;
        RECT 52.745 37.040 53.480 37.230 ;
        RECT 52.745 36.240 53.100 37.040 ;
        RECT 53.250 36.970 53.480 37.040 ;
        RECT 53.690 37.925 53.920 37.970 ;
        RECT 54.060 37.925 54.300 38.110 ;
        RECT 53.690 37.595 54.300 37.925 ;
        RECT 55.275 37.870 55.505 37.975 ;
        RECT 53.690 37.040 54.185 37.595 ;
        RECT 53.690 36.970 53.920 37.040 ;
        RECT 53.440 36.785 53.730 36.810 ;
        RECT 53.425 36.535 53.760 36.785 ;
        RECT 55.045 36.765 55.505 37.870 ;
        RECT 54.725 36.240 55.505 36.765 ;
        RECT 52.305 36.060 55.505 36.240 ;
        RECT 51.670 35.965 51.900 36.020 ;
        RECT 47.660 35.575 51.620 35.805 ;
        RECT 52.305 35.620 55.110 36.060 ;
        RECT 55.275 35.975 55.505 36.060 ;
        RECT 55.715 37.910 55.945 37.975 ;
        RECT 56.110 37.910 56.480 38.795 ;
        RECT 55.715 37.585 56.480 37.910 ;
        RECT 55.715 36.045 56.475 37.585 ;
        RECT 55.715 35.975 55.945 36.045 ;
        RECT 55.465 35.795 55.755 35.815 ;
        RECT 52.305 35.255 54.770 35.620 ;
        RECT 55.440 35.545 55.775 35.795 ;
        RECT 58.010 35.280 58.505 40.395 ;
        RECT 59.525 40.345 59.730 40.480 ;
        RECT 61.010 40.395 61.240 40.645 ;
        RECT 62.030 40.550 62.780 40.990 ;
        RECT 63.200 40.775 64.215 41.775 ;
        RECT 58.805 40.115 60.805 40.345 ;
        RECT 62.030 38.355 62.400 40.550 ;
        RECT 62.550 40.490 62.780 40.550 ;
        RECT 63.270 40.285 64.160 40.775 ;
        RECT 64.840 40.580 66.210 48.380 ;
        RECT 66.745 43.635 67.635 48.695 ;
        RECT 68.270 48.410 68.500 48.490 ;
        RECT 66.740 42.015 67.640 43.635 ;
        RECT 66.745 41.605 67.635 42.015 ;
        RECT 66.670 40.605 67.700 41.605 ;
        RECT 68.270 40.625 68.645 48.410 ;
        RECT 68.920 48.025 70.600 49.260 ;
        RECT 71.435 48.025 76.360 48.035 ;
        RECT 68.920 47.545 76.360 48.025 ;
        RECT 68.920 45.285 70.600 47.545 ;
        RECT 71.435 47.125 76.360 47.545 ;
        RECT 70.940 46.935 71.195 46.960 ;
        RECT 70.940 46.920 71.215 46.935 ;
        RECT 70.910 46.645 71.245 46.920 ;
        RECT 71.420 46.895 76.420 47.125 ;
        RECT 76.630 46.935 76.885 46.960 ;
        RECT 70.940 46.630 71.195 46.645 ;
        RECT 71.420 46.455 76.420 46.685 ;
        RECT 76.625 46.645 76.885 46.935 ;
        RECT 76.630 46.630 76.885 46.645 ;
        RECT 71.465 46.445 76.320 46.455 ;
        RECT 71.465 44.920 74.110 44.925 ;
        RECT 70.140 44.720 74.110 44.920 ;
        RECT 70.140 44.690 74.100 44.720 ;
        RECT 68.980 44.335 69.315 44.610 ;
        RECT 69.860 44.440 70.090 44.485 ;
        RECT 64.840 40.560 65.195 40.580 ;
        RECT 64.840 40.490 65.070 40.560 ;
        RECT 65.980 40.490 66.210 40.580 ;
        RECT 66.740 40.465 67.650 40.605 ;
        RECT 68.270 40.490 68.660 40.625 ;
        RECT 66.730 40.285 67.740 40.465 ;
        RECT 62.830 40.055 64.790 40.285 ;
        RECT 66.260 40.055 68.220 40.285 ;
        RECT 63.535 39.230 63.880 40.055 ;
        RECT 66.285 40.050 68.170 40.055 ;
        RECT 68.465 38.355 68.660 40.490 ;
        RECT 69.050 38.830 69.240 44.335 ;
        RECT 69.670 43.105 70.090 44.440 ;
        RECT 71.395 43.105 72.740 44.690 ;
        RECT 69.670 41.720 72.740 43.105 ;
        RECT 69.670 40.990 70.090 41.720 ;
        RECT 69.665 40.485 70.090 40.990 ;
        RECT 69.050 38.640 69.365 38.830 ;
        RECT 59.370 38.125 63.330 38.355 ;
        RECT 64.800 38.125 68.760 38.355 ;
        RECT 69.175 38.130 69.365 38.640 ;
        RECT 59.090 37.515 59.320 37.965 ;
        RECT 60.570 37.515 61.360 38.125 ;
        RECT 59.090 37.210 61.360 37.515 ;
        RECT 59.035 37.195 61.360 37.210 ;
        RECT 58.950 36.350 61.360 37.195 ;
        RECT 58.950 35.975 59.320 36.350 ;
        RECT 59.090 35.965 59.320 35.975 ;
        RECT 60.570 35.805 61.360 36.350 ;
        RECT 63.380 37.880 63.610 37.965 ;
        RECT 64.520 37.880 64.750 37.965 ;
        RECT 63.380 36.055 64.750 37.880 ;
        RECT 63.380 35.965 63.610 36.055 ;
        RECT 59.370 35.575 63.330 35.805 ;
        RECT 56.010 35.255 58.505 35.280 ;
        RECT 58.950 35.255 59.175 35.265 ;
        RECT 63.850 35.255 64.340 36.055 ;
        RECT 64.520 35.965 64.750 36.055 ;
        RECT 66.235 37.745 67.575 38.125 ;
        RECT 68.810 37.745 69.040 37.965 ;
        RECT 66.235 36.150 69.040 37.745 ;
        RECT 66.235 35.805 67.575 36.150 ;
        RECT 68.810 35.965 69.040 36.150 ;
        RECT 64.800 35.575 68.760 35.805 ;
        RECT 69.190 35.785 69.365 38.130 ;
        RECT 69.665 37.965 69.960 40.485 ;
        RECT 71.395 40.280 72.740 41.720 ;
        RECT 74.150 44.390 74.380 44.485 ;
        RECT 74.625 44.390 75.115 46.445 ;
        RECT 75.685 44.920 76.320 44.925 ;
        RECT 75.570 44.690 79.530 44.920 ;
        RECT 75.290 44.390 75.520 44.485 ;
        RECT 74.150 40.565 75.520 44.390 ;
        RECT 74.150 40.485 74.380 40.565 ;
        RECT 75.290 40.485 75.520 40.565 ;
        RECT 76.945 40.280 78.290 44.690 ;
        RECT 79.580 44.420 79.810 44.485 ;
        RECT 80.465 44.425 80.940 49.260 ;
        RECT 82.265 48.455 82.945 49.260 ;
        RECT 83.365 48.735 83.700 48.985 ;
        RECT 83.380 48.710 83.670 48.735 ;
        RECT 86.840 48.635 88.750 49.260 ;
        RECT 90.840 48.925 92.725 48.930 ;
        RECT 94.285 48.925 96.170 48.930 ;
        RECT 90.830 48.695 92.790 48.925 ;
        RECT 94.260 48.695 96.220 48.925 ;
        RECT 83.190 48.455 83.420 48.505 ;
        RECT 82.265 47.955 83.420 48.455 ;
        RECT 81.335 44.735 81.670 44.985 ;
        RECT 81.355 44.705 81.645 44.735 ;
        RECT 81.165 44.425 81.395 44.500 ;
        RECT 79.580 40.485 80.035 44.420 ;
        RECT 80.465 43.680 81.395 44.425 ;
        RECT 80.800 40.565 81.395 43.680 ;
        RECT 81.165 40.500 81.395 40.565 ;
        RECT 81.605 44.475 81.835 44.500 ;
        RECT 81.605 40.920 82.115 44.475 ;
        RECT 81.605 40.550 82.300 40.920 ;
        RECT 82.800 40.600 83.420 47.955 ;
        RECT 81.605 40.500 81.835 40.550 ;
        RECT 70.140 40.250 74.100 40.280 ;
        RECT 75.570 40.250 79.530 40.280 ;
        RECT 70.140 40.090 79.530 40.250 ;
        RECT 70.140 40.050 74.100 40.090 ;
        RECT 75.570 40.050 79.530 40.090 ;
        RECT 79.695 38.660 80.035 40.485 ;
        RECT 81.345 38.660 81.765 40.305 ;
        RECT 79.695 38.505 81.765 38.660 ;
        RECT 79.770 38.390 81.765 38.505 ;
        RECT 70.230 38.125 74.190 38.355 ;
        RECT 75.660 38.125 79.620 38.355 ;
        RECT 69.665 37.205 70.180 37.965 ;
        RECT 69.735 36.025 70.180 37.205 ;
        RECT 69.950 35.965 70.180 36.025 ;
        RECT 71.610 35.805 72.565 38.125 ;
        RECT 74.240 37.900 74.470 37.965 ;
        RECT 75.380 37.900 75.610 37.965 ;
        RECT 74.240 36.030 75.610 37.900 ;
        RECT 74.240 35.965 74.470 36.030 ;
        RECT 69.175 35.255 69.365 35.785 ;
        RECT 70.230 35.575 74.190 35.805 ;
        RECT 74.645 35.255 75.200 36.030 ;
        RECT 75.380 35.965 75.610 36.030 ;
        RECT 77.055 35.805 78.010 38.125 ;
        RECT 79.770 37.970 80.035 38.390 ;
        RECT 81.345 38.115 81.765 38.390 ;
        RECT 82.000 39.355 82.300 40.550 ;
        RECT 83.190 40.505 83.420 40.600 ;
        RECT 83.630 48.430 83.860 48.505 ;
        RECT 83.630 41.110 84.405 48.430 ;
        RECT 86.805 48.405 88.805 48.635 ;
        RECT 90.550 48.410 90.780 48.490 ;
        RECT 86.370 45.060 86.600 48.355 ;
        RECT 89.010 48.275 89.240 48.355 ;
        RECT 88.980 45.060 89.240 48.275 ;
        RECT 86.370 43.245 89.240 45.060 ;
        RECT 83.630 40.580 84.480 41.110 ;
        RECT 86.370 40.825 86.600 43.245 ;
        RECT 83.630 40.505 83.860 40.580 ;
        RECT 83.295 39.825 83.810 40.315 ;
        RECT 83.295 39.360 83.805 39.825 ;
        RECT 84.110 39.795 84.480 40.580 ;
        RECT 86.010 40.395 86.600 40.825 ;
        RECT 87.495 40.640 87.755 40.960 ;
        RECT 88.980 40.645 89.240 43.245 ;
        RECT 90.310 40.990 90.780 48.410 ;
        RECT 91.270 41.775 92.160 48.695 ;
        RECT 92.840 48.390 93.070 48.490 ;
        RECT 92.840 48.380 93.195 48.390 ;
        RECT 93.980 48.380 94.210 48.490 ;
        RECT 87.550 40.480 87.700 40.640 ;
        RECT 82.930 39.355 83.805 39.360 ;
        RECT 82.000 38.950 83.805 39.355 ;
        RECT 82.000 38.110 82.300 38.950 ;
        RECT 82.930 38.935 83.805 38.950 ;
        RECT 83.295 38.825 83.805 38.935 ;
        RECT 83.295 38.125 83.810 38.825 ;
        RECT 84.005 38.795 85.035 39.795 ;
        RECT 79.695 37.965 80.035 37.970 ;
        RECT 79.670 36.020 80.035 37.965 ;
        RECT 81.250 37.900 81.480 37.970 ;
        RECT 80.755 37.230 81.480 37.900 ;
        RECT 80.745 37.040 81.480 37.230 ;
        RECT 80.745 36.240 81.100 37.040 ;
        RECT 81.250 36.970 81.480 37.040 ;
        RECT 81.690 37.925 81.920 37.970 ;
        RECT 82.060 37.925 82.300 38.110 ;
        RECT 81.690 37.595 82.300 37.925 ;
        RECT 83.275 37.870 83.505 37.975 ;
        RECT 81.690 37.040 82.185 37.595 ;
        RECT 81.690 36.970 81.920 37.040 ;
        RECT 81.440 36.785 81.730 36.810 ;
        RECT 81.425 36.535 81.760 36.785 ;
        RECT 83.045 36.765 83.505 37.870 ;
        RECT 82.725 36.240 83.505 36.765 ;
        RECT 80.305 36.060 83.505 36.240 ;
        RECT 79.670 35.965 79.900 36.020 ;
        RECT 80.305 35.960 83.110 36.060 ;
        RECT 83.275 35.975 83.505 36.060 ;
        RECT 83.715 37.910 83.945 37.975 ;
        RECT 84.110 37.910 84.480 38.795 ;
        RECT 83.715 37.585 84.480 37.910 ;
        RECT 83.715 36.045 84.475 37.585 ;
        RECT 83.715 35.975 83.945 36.045 ;
        RECT 75.660 35.575 79.620 35.805 ;
        RECT 80.250 35.785 83.110 35.960 ;
        RECT 83.465 35.795 83.755 35.815 ;
        RECT 80.290 35.620 83.110 35.785 ;
        RECT 80.290 35.255 82.770 35.620 ;
        RECT 83.440 35.545 83.775 35.795 ;
        RECT 86.010 35.280 86.505 40.395 ;
        RECT 87.525 40.345 87.730 40.480 ;
        RECT 89.010 40.395 89.240 40.645 ;
        RECT 90.030 40.550 90.780 40.990 ;
        RECT 91.200 40.775 92.215 41.775 ;
        RECT 86.805 40.115 88.805 40.345 ;
        RECT 90.030 38.355 90.400 40.550 ;
        RECT 90.550 40.490 90.780 40.550 ;
        RECT 91.270 40.285 92.160 40.775 ;
        RECT 92.840 40.580 94.210 48.380 ;
        RECT 94.745 43.635 95.635 48.695 ;
        RECT 96.270 48.410 96.500 48.490 ;
        RECT 94.740 42.015 95.640 43.635 ;
        RECT 94.745 41.605 95.635 42.015 ;
        RECT 94.670 40.605 95.700 41.605 ;
        RECT 96.270 40.625 96.645 48.410 ;
        RECT 96.920 48.025 98.600 49.260 ;
        RECT 99.435 48.025 104.360 48.035 ;
        RECT 96.920 47.545 104.360 48.025 ;
        RECT 96.920 45.285 98.600 47.545 ;
        RECT 99.435 47.125 104.360 47.545 ;
        RECT 98.940 46.935 99.195 46.960 ;
        RECT 98.940 46.920 99.215 46.935 ;
        RECT 98.910 46.645 99.245 46.920 ;
        RECT 99.420 46.895 104.420 47.125 ;
        RECT 104.630 46.935 104.885 46.960 ;
        RECT 98.940 46.630 99.195 46.645 ;
        RECT 99.420 46.455 104.420 46.685 ;
        RECT 104.625 46.645 104.885 46.935 ;
        RECT 104.630 46.630 104.885 46.645 ;
        RECT 99.465 46.445 104.320 46.455 ;
        RECT 99.465 44.920 102.110 44.925 ;
        RECT 98.140 44.720 102.110 44.920 ;
        RECT 98.140 44.690 102.100 44.720 ;
        RECT 96.980 44.335 97.315 44.610 ;
        RECT 97.860 44.440 98.090 44.485 ;
        RECT 92.840 40.560 93.195 40.580 ;
        RECT 92.840 40.490 93.070 40.560 ;
        RECT 93.980 40.490 94.210 40.580 ;
        RECT 94.740 40.465 95.650 40.605 ;
        RECT 96.270 40.490 96.660 40.625 ;
        RECT 94.730 40.285 95.740 40.465 ;
        RECT 90.830 40.055 92.790 40.285 ;
        RECT 94.260 40.055 96.220 40.285 ;
        RECT 91.515 39.170 91.915 40.055 ;
        RECT 94.285 40.050 96.170 40.055 ;
        RECT 96.465 38.355 96.660 40.490 ;
        RECT 97.050 38.830 97.240 44.335 ;
        RECT 97.670 43.105 98.090 44.440 ;
        RECT 99.395 43.105 100.740 44.690 ;
        RECT 97.670 41.720 100.740 43.105 ;
        RECT 97.670 40.990 98.090 41.720 ;
        RECT 97.665 40.485 98.090 40.990 ;
        RECT 97.050 38.640 97.365 38.830 ;
        RECT 87.370 38.125 91.330 38.355 ;
        RECT 92.800 38.125 96.760 38.355 ;
        RECT 97.175 38.130 97.365 38.640 ;
        RECT 87.090 37.515 87.320 37.965 ;
        RECT 88.570 37.515 89.360 38.125 ;
        RECT 87.090 37.210 89.360 37.515 ;
        RECT 87.035 37.195 89.360 37.210 ;
        RECT 86.950 36.350 89.360 37.195 ;
        RECT 86.950 35.975 87.320 36.350 ;
        RECT 87.090 35.965 87.320 35.975 ;
        RECT 88.570 35.805 89.360 36.350 ;
        RECT 91.380 37.880 91.610 37.965 ;
        RECT 92.520 37.880 92.750 37.965 ;
        RECT 91.380 36.055 92.750 37.880 ;
        RECT 91.380 35.965 91.610 36.055 ;
        RECT 87.370 35.575 91.330 35.805 ;
        RECT 84.010 35.255 86.505 35.280 ;
        RECT 86.950 35.255 87.175 35.265 ;
        RECT 91.850 35.255 92.340 36.055 ;
        RECT 92.520 35.965 92.750 36.055 ;
        RECT 94.235 37.745 95.575 38.125 ;
        RECT 96.810 37.745 97.040 37.965 ;
        RECT 94.235 36.150 97.040 37.745 ;
        RECT 94.235 35.805 95.575 36.150 ;
        RECT 96.810 35.965 97.040 36.150 ;
        RECT 92.800 35.575 96.760 35.805 ;
        RECT 97.190 35.785 97.365 38.130 ;
        RECT 97.665 37.965 97.960 40.485 ;
        RECT 99.395 40.280 100.740 41.720 ;
        RECT 102.150 44.390 102.380 44.485 ;
        RECT 102.625 44.390 103.115 46.445 ;
        RECT 103.685 44.920 104.320 44.925 ;
        RECT 103.570 44.690 107.530 44.920 ;
        RECT 103.290 44.390 103.520 44.485 ;
        RECT 102.150 40.565 103.520 44.390 ;
        RECT 102.150 40.485 102.380 40.565 ;
        RECT 103.290 40.485 103.520 40.565 ;
        RECT 104.945 40.280 106.290 44.690 ;
        RECT 107.580 44.420 107.810 44.485 ;
        RECT 108.465 44.425 108.940 49.260 ;
        RECT 110.265 48.455 110.945 49.260 ;
        RECT 111.365 48.735 111.700 48.985 ;
        RECT 111.380 48.710 111.670 48.735 ;
        RECT 114.840 48.635 116.750 49.260 ;
        RECT 118.840 48.925 120.725 48.930 ;
        RECT 122.285 48.925 124.170 48.930 ;
        RECT 118.830 48.695 120.790 48.925 ;
        RECT 122.260 48.695 124.220 48.925 ;
        RECT 111.190 48.455 111.420 48.505 ;
        RECT 110.265 47.955 111.420 48.455 ;
        RECT 109.335 44.735 109.670 44.985 ;
        RECT 109.355 44.705 109.645 44.735 ;
        RECT 109.165 44.425 109.395 44.500 ;
        RECT 107.580 40.485 108.035 44.420 ;
        RECT 108.465 43.680 109.395 44.425 ;
        RECT 108.800 40.565 109.395 43.680 ;
        RECT 109.165 40.500 109.395 40.565 ;
        RECT 109.605 44.475 109.835 44.500 ;
        RECT 109.605 40.920 110.115 44.475 ;
        RECT 109.605 40.550 110.300 40.920 ;
        RECT 110.800 40.600 111.420 47.955 ;
        RECT 109.605 40.500 109.835 40.550 ;
        RECT 98.140 40.250 102.100 40.280 ;
        RECT 103.570 40.250 107.530 40.280 ;
        RECT 98.140 40.090 107.530 40.250 ;
        RECT 98.140 40.050 102.100 40.090 ;
        RECT 103.570 40.050 107.530 40.090 ;
        RECT 107.695 38.660 108.035 40.485 ;
        RECT 109.345 38.660 109.765 40.305 ;
        RECT 107.695 38.505 109.765 38.660 ;
        RECT 107.770 38.390 109.765 38.505 ;
        RECT 98.230 38.125 102.190 38.355 ;
        RECT 103.660 38.125 107.620 38.355 ;
        RECT 97.665 37.205 98.180 37.965 ;
        RECT 97.735 36.025 98.180 37.205 ;
        RECT 97.950 35.965 98.180 36.025 ;
        RECT 99.610 35.805 100.565 38.125 ;
        RECT 102.240 37.900 102.470 37.965 ;
        RECT 103.380 37.900 103.610 37.965 ;
        RECT 102.240 36.030 103.610 37.900 ;
        RECT 102.240 35.965 102.470 36.030 ;
        RECT 97.175 35.255 97.365 35.785 ;
        RECT 98.230 35.575 102.190 35.805 ;
        RECT 102.645 35.255 103.200 36.030 ;
        RECT 103.380 35.965 103.610 36.030 ;
        RECT 105.055 35.805 106.010 38.125 ;
        RECT 107.770 37.970 108.035 38.390 ;
        RECT 109.345 38.115 109.765 38.390 ;
        RECT 110.000 39.355 110.300 40.550 ;
        RECT 111.190 40.505 111.420 40.600 ;
        RECT 111.630 48.430 111.860 48.505 ;
        RECT 111.630 41.110 112.405 48.430 ;
        RECT 114.805 48.405 116.805 48.635 ;
        RECT 118.550 48.410 118.780 48.490 ;
        RECT 114.370 45.060 114.600 48.355 ;
        RECT 117.010 48.275 117.240 48.355 ;
        RECT 116.980 45.060 117.240 48.275 ;
        RECT 114.370 43.245 117.240 45.060 ;
        RECT 111.630 40.580 112.480 41.110 ;
        RECT 114.370 40.825 114.600 43.245 ;
        RECT 111.630 40.505 111.860 40.580 ;
        RECT 111.295 39.825 111.810 40.315 ;
        RECT 111.295 39.360 111.805 39.825 ;
        RECT 112.110 39.795 112.480 40.580 ;
        RECT 114.010 40.395 114.600 40.825 ;
        RECT 115.495 40.640 115.755 40.960 ;
        RECT 116.980 40.645 117.240 43.245 ;
        RECT 118.310 40.990 118.780 48.410 ;
        RECT 119.270 41.775 120.160 48.695 ;
        RECT 120.840 48.390 121.070 48.490 ;
        RECT 120.840 48.380 121.195 48.390 ;
        RECT 121.980 48.380 122.210 48.490 ;
        RECT 115.550 40.480 115.700 40.640 ;
        RECT 110.930 39.355 111.805 39.360 ;
        RECT 110.000 38.950 111.805 39.355 ;
        RECT 110.000 38.110 110.300 38.950 ;
        RECT 110.930 38.935 111.805 38.950 ;
        RECT 111.295 38.825 111.805 38.935 ;
        RECT 111.295 38.125 111.810 38.825 ;
        RECT 112.005 38.795 113.035 39.795 ;
        RECT 107.695 37.965 108.035 37.970 ;
        RECT 107.670 36.020 108.035 37.965 ;
        RECT 109.250 37.900 109.480 37.970 ;
        RECT 108.755 37.230 109.480 37.900 ;
        RECT 108.745 37.040 109.480 37.230 ;
        RECT 108.745 36.240 109.100 37.040 ;
        RECT 109.250 36.970 109.480 37.040 ;
        RECT 109.690 37.925 109.920 37.970 ;
        RECT 110.060 37.925 110.300 38.110 ;
        RECT 109.690 37.595 110.300 37.925 ;
        RECT 111.275 37.870 111.505 37.975 ;
        RECT 109.690 37.040 110.185 37.595 ;
        RECT 109.690 36.970 109.920 37.040 ;
        RECT 109.440 36.785 109.730 36.810 ;
        RECT 109.425 36.535 109.760 36.785 ;
        RECT 111.045 36.765 111.505 37.870 ;
        RECT 110.725 36.240 111.505 36.765 ;
        RECT 108.305 36.060 111.505 36.240 ;
        RECT 107.670 35.965 107.900 36.020 ;
        RECT 103.660 35.575 107.620 35.805 ;
        RECT 108.305 35.620 111.110 36.060 ;
        RECT 111.275 35.975 111.505 36.060 ;
        RECT 111.715 37.910 111.945 37.975 ;
        RECT 112.110 37.910 112.480 38.795 ;
        RECT 111.715 37.585 112.480 37.910 ;
        RECT 111.715 36.045 112.475 37.585 ;
        RECT 111.715 35.975 111.945 36.045 ;
        RECT 111.465 35.795 111.755 35.815 ;
        RECT 108.305 35.255 110.770 35.620 ;
        RECT 111.440 35.545 111.775 35.795 ;
        RECT 114.010 35.280 114.505 40.395 ;
        RECT 115.525 40.345 115.730 40.480 ;
        RECT 117.010 40.395 117.240 40.645 ;
        RECT 118.030 40.550 118.780 40.990 ;
        RECT 119.200 40.775 120.215 41.775 ;
        RECT 114.805 40.115 116.805 40.345 ;
        RECT 118.030 38.355 118.400 40.550 ;
        RECT 118.550 40.490 118.780 40.550 ;
        RECT 119.270 40.285 120.160 40.775 ;
        RECT 120.840 40.580 122.210 48.380 ;
        RECT 122.745 43.635 123.635 48.695 ;
        RECT 124.270 48.410 124.500 48.490 ;
        RECT 122.740 42.015 123.640 43.635 ;
        RECT 122.745 41.605 123.635 42.015 ;
        RECT 122.670 40.605 123.700 41.605 ;
        RECT 124.270 40.625 124.645 48.410 ;
        RECT 124.920 48.025 126.600 49.260 ;
        RECT 127.435 48.025 132.360 48.035 ;
        RECT 124.920 47.545 132.360 48.025 ;
        RECT 124.920 45.285 126.600 47.545 ;
        RECT 127.435 47.125 132.360 47.545 ;
        RECT 126.940 46.935 127.195 46.960 ;
        RECT 126.940 46.920 127.215 46.935 ;
        RECT 126.910 46.645 127.245 46.920 ;
        RECT 127.420 46.895 132.420 47.125 ;
        RECT 132.630 46.935 132.885 46.960 ;
        RECT 126.940 46.630 127.195 46.645 ;
        RECT 127.420 46.455 132.420 46.685 ;
        RECT 132.625 46.645 132.885 46.935 ;
        RECT 132.630 46.630 132.885 46.645 ;
        RECT 127.465 46.445 132.320 46.455 ;
        RECT 127.465 44.920 130.110 44.925 ;
        RECT 126.140 44.720 130.110 44.920 ;
        RECT 126.140 44.690 130.100 44.720 ;
        RECT 124.980 44.335 125.315 44.610 ;
        RECT 125.860 44.440 126.090 44.485 ;
        RECT 120.840 40.560 121.195 40.580 ;
        RECT 120.840 40.490 121.070 40.560 ;
        RECT 121.980 40.490 122.210 40.580 ;
        RECT 122.740 40.465 123.650 40.605 ;
        RECT 124.270 40.490 124.660 40.625 ;
        RECT 122.730 40.285 123.740 40.465 ;
        RECT 118.830 40.055 120.790 40.285 ;
        RECT 122.260 40.055 124.220 40.285 ;
        RECT 119.565 39.135 119.850 40.055 ;
        RECT 122.285 40.050 124.170 40.055 ;
        RECT 124.465 38.355 124.660 40.490 ;
        RECT 125.050 38.830 125.240 44.335 ;
        RECT 125.670 43.105 126.090 44.440 ;
        RECT 127.395 43.105 128.740 44.690 ;
        RECT 125.670 41.720 128.740 43.105 ;
        RECT 125.670 40.990 126.090 41.720 ;
        RECT 125.665 40.485 126.090 40.990 ;
        RECT 125.050 38.640 125.365 38.830 ;
        RECT 115.370 38.125 119.330 38.355 ;
        RECT 120.800 38.125 124.760 38.355 ;
        RECT 125.175 38.130 125.365 38.640 ;
        RECT 115.090 37.515 115.320 37.965 ;
        RECT 116.570 37.515 117.360 38.125 ;
        RECT 115.090 37.210 117.360 37.515 ;
        RECT 115.035 37.195 117.360 37.210 ;
        RECT 114.950 36.350 117.360 37.195 ;
        RECT 114.950 35.975 115.320 36.350 ;
        RECT 115.090 35.965 115.320 35.975 ;
        RECT 116.570 35.805 117.360 36.350 ;
        RECT 119.380 37.880 119.610 37.965 ;
        RECT 120.520 37.880 120.750 37.965 ;
        RECT 119.380 36.055 120.750 37.880 ;
        RECT 119.380 35.965 119.610 36.055 ;
        RECT 115.370 35.575 119.330 35.805 ;
        RECT 111.910 35.255 114.610 35.280 ;
        RECT 114.950 35.255 115.175 35.265 ;
        RECT 119.850 35.255 120.340 36.055 ;
        RECT 120.520 35.965 120.750 36.055 ;
        RECT 122.235 37.745 123.575 38.125 ;
        RECT 124.810 37.745 125.040 37.965 ;
        RECT 122.235 36.150 125.040 37.745 ;
        RECT 122.235 35.805 123.575 36.150 ;
        RECT 124.810 35.965 125.040 36.150 ;
        RECT 120.800 35.575 124.760 35.805 ;
        RECT 125.190 35.785 125.365 38.130 ;
        RECT 125.665 37.965 125.960 40.485 ;
        RECT 127.395 40.280 128.740 41.720 ;
        RECT 130.150 44.390 130.380 44.485 ;
        RECT 130.625 44.390 131.115 46.445 ;
        RECT 131.685 44.920 132.320 44.925 ;
        RECT 131.570 44.690 135.530 44.920 ;
        RECT 131.290 44.390 131.520 44.485 ;
        RECT 130.150 40.565 131.520 44.390 ;
        RECT 130.150 40.485 130.380 40.565 ;
        RECT 131.290 40.485 131.520 40.565 ;
        RECT 132.945 40.280 134.290 44.690 ;
        RECT 135.580 44.420 135.810 44.485 ;
        RECT 136.465 44.425 136.940 49.260 ;
        RECT 138.265 48.455 138.945 49.260 ;
        RECT 139.365 48.735 139.700 48.985 ;
        RECT 139.380 48.710 139.670 48.735 ;
        RECT 144.570 48.720 146.675 49.310 ;
        RECT 147.255 48.720 149.360 49.310 ;
        RECT 139.190 48.455 139.420 48.505 ;
        RECT 138.265 47.955 139.420 48.455 ;
        RECT 137.335 44.735 137.670 44.985 ;
        RECT 137.355 44.705 137.645 44.735 ;
        RECT 137.165 44.425 137.395 44.500 ;
        RECT 135.580 40.485 136.035 44.420 ;
        RECT 136.465 43.680 137.395 44.425 ;
        RECT 136.800 40.565 137.395 43.680 ;
        RECT 137.165 40.500 137.395 40.565 ;
        RECT 137.605 44.475 137.835 44.500 ;
        RECT 137.605 40.920 138.115 44.475 ;
        RECT 137.605 40.550 138.300 40.920 ;
        RECT 138.800 40.600 139.420 47.955 ;
        RECT 137.605 40.500 137.835 40.550 ;
        RECT 126.140 40.250 130.100 40.280 ;
        RECT 131.570 40.250 135.530 40.280 ;
        RECT 126.140 40.090 135.530 40.250 ;
        RECT 126.140 40.050 130.100 40.090 ;
        RECT 131.570 40.050 135.530 40.090 ;
        RECT 135.695 38.660 136.035 40.485 ;
        RECT 137.345 38.660 137.765 40.305 ;
        RECT 135.695 38.505 137.765 38.660 ;
        RECT 135.770 38.390 137.765 38.505 ;
        RECT 126.230 38.125 130.190 38.355 ;
        RECT 131.660 38.125 135.620 38.355 ;
        RECT 125.665 37.205 126.180 37.965 ;
        RECT 125.735 36.025 126.180 37.205 ;
        RECT 125.950 35.965 126.180 36.025 ;
        RECT 127.610 35.805 128.565 38.125 ;
        RECT 130.240 37.900 130.470 37.965 ;
        RECT 131.380 37.900 131.610 37.965 ;
        RECT 130.240 36.030 131.610 37.900 ;
        RECT 130.240 35.965 130.470 36.030 ;
        RECT 125.175 35.255 125.365 35.785 ;
        RECT 126.230 35.575 130.190 35.805 ;
        RECT 130.645 35.255 131.200 36.030 ;
        RECT 131.380 35.965 131.610 36.030 ;
        RECT 133.055 35.805 134.010 38.125 ;
        RECT 135.770 37.970 136.035 38.390 ;
        RECT 137.345 38.115 137.765 38.390 ;
        RECT 138.000 39.355 138.300 40.550 ;
        RECT 139.190 40.505 139.420 40.600 ;
        RECT 139.630 48.430 139.860 48.505 ;
        RECT 139.630 41.110 140.405 48.430 ;
        RECT 147.280 47.490 149.310 48.720 ;
        RECT 144.570 46.900 146.675 47.490 ;
        RECT 147.255 46.900 149.360 47.490 ;
        RECT 144.580 45.670 146.610 46.900 ;
        RECT 147.310 46.880 149.310 46.900 ;
        RECT 147.310 45.670 155.310 45.680 ;
        RECT 144.570 45.080 146.675 45.670 ;
        RECT 147.255 45.180 155.310 45.670 ;
        RECT 147.255 45.080 149.360 45.180 ;
        RECT 144.610 43.850 146.610 43.880 ;
        RECT 144.570 43.260 146.675 43.850 ;
        RECT 147.255 43.780 149.360 43.850 ;
        RECT 149.845 43.780 150.345 44.125 ;
        RECT 153.310 43.850 155.310 45.180 ;
        RECT 150.550 43.780 152.655 43.850 ;
        RECT 147.255 43.280 152.655 43.780 ;
        RECT 147.255 43.260 149.360 43.280 ;
        RECT 150.550 43.260 152.655 43.280 ;
        RECT 153.235 43.260 155.340 43.850 ;
        RECT 144.610 42.945 146.610 43.260 ;
        RECT 142.210 42.505 146.610 42.945 ;
        RECT 144.610 42.030 146.610 42.505 ;
        RECT 144.570 41.440 146.675 42.030 ;
        RECT 147.255 41.980 149.360 42.030 ;
        RECT 150.550 41.980 152.655 42.030 ;
        RECT 147.255 41.480 152.655 41.980 ;
        RECT 147.255 41.440 149.360 41.480 ;
        RECT 149.950 41.440 152.655 41.480 ;
        RECT 153.235 41.440 155.340 42.030 ;
        RECT 149.950 41.240 150.730 41.440 ;
        RECT 139.630 40.580 140.480 41.110 ;
        RECT 149.950 41.035 150.450 41.240 ;
        RECT 139.630 40.505 139.860 40.580 ;
        RECT 139.295 39.825 139.810 40.315 ;
        RECT 139.295 39.360 139.805 39.825 ;
        RECT 140.110 39.795 140.480 40.580 ;
        RECT 142.770 40.535 150.450 41.035 ;
        RECT 153.985 40.995 154.775 41.440 ;
        RECT 151.205 40.205 154.775 40.995 ;
        RECT 151.205 40.055 151.995 40.205 ;
        RECT 138.930 39.355 139.805 39.360 ;
        RECT 138.000 38.950 139.805 39.355 ;
        RECT 138.000 38.110 138.300 38.950 ;
        RECT 138.930 38.935 139.805 38.950 ;
        RECT 139.295 38.825 139.805 38.935 ;
        RECT 139.295 38.125 139.810 38.825 ;
        RECT 140.005 38.795 141.035 39.795 ;
        RECT 141.525 39.265 151.995 40.055 ;
        RECT 135.695 37.965 136.035 37.970 ;
        RECT 135.670 36.020 136.035 37.965 ;
        RECT 137.250 37.900 137.480 37.970 ;
        RECT 136.755 37.230 137.480 37.900 ;
        RECT 136.745 37.040 137.480 37.230 ;
        RECT 136.745 36.240 137.100 37.040 ;
        RECT 137.250 36.970 137.480 37.040 ;
        RECT 137.690 37.925 137.920 37.970 ;
        RECT 138.060 37.925 138.300 38.110 ;
        RECT 137.690 37.595 138.300 37.925 ;
        RECT 139.275 37.870 139.505 37.975 ;
        RECT 137.690 37.040 138.185 37.595 ;
        RECT 137.690 36.970 137.920 37.040 ;
        RECT 137.440 36.785 137.730 36.810 ;
        RECT 137.425 36.535 137.760 36.785 ;
        RECT 139.045 36.765 139.505 37.870 ;
        RECT 138.725 36.240 139.505 36.765 ;
        RECT 136.305 36.060 139.505 36.240 ;
        RECT 135.670 35.965 135.900 36.020 ;
        RECT 131.660 35.575 135.620 35.805 ;
        RECT 136.305 35.620 139.110 36.060 ;
        RECT 139.275 35.975 139.505 36.060 ;
        RECT 139.715 37.910 139.945 37.975 ;
        RECT 140.110 37.910 140.480 38.795 ;
        RECT 139.715 37.585 140.480 37.910 ;
        RECT 139.715 36.045 140.475 37.585 ;
        RECT 139.715 35.975 139.945 36.045 ;
        RECT 139.465 35.795 139.755 35.815 ;
        RECT 136.305 35.335 138.770 35.620 ;
        RECT 139.440 35.545 139.775 35.795 ;
        RECT 141.525 35.335 142.315 39.265 ;
        RECT 136.305 35.255 142.315 35.335 ;
        RECT 1.895 34.545 142.315 35.255 ;
        RECT 1.895 34.380 140.500 34.545 ;
        RECT 28.210 33.960 30.910 33.980 ;
        RECT 55.810 33.960 58.410 33.980 ;
        RECT 83.810 33.960 86.710 33.980 ;
        RECT 111.610 33.960 114.610 33.980 ;
        RECT 1.870 33.280 140.345 33.960 ;
        RECT 1.870 33.260 28.345 33.280 ;
        RECT 29.870 33.260 84.345 33.280 ;
        RECT 85.870 33.260 112.345 33.280 ;
        RECT 113.870 33.260 140.345 33.280 ;
        RECT 2.840 32.635 4.750 33.260 ;
        RECT 6.840 32.925 8.725 32.930 ;
        RECT 10.285 32.925 12.170 32.930 ;
        RECT 6.830 32.695 8.790 32.925 ;
        RECT 10.260 32.695 12.220 32.925 ;
        RECT 2.805 32.405 4.805 32.635 ;
        RECT 6.550 32.410 6.780 32.490 ;
        RECT 2.370 29.060 2.600 32.355 ;
        RECT 5.010 32.275 5.240 32.355 ;
        RECT 4.980 29.060 5.240 32.275 ;
        RECT 2.370 27.245 5.240 29.060 ;
        RECT 2.370 24.825 2.600 27.245 ;
        RECT 2.010 24.395 2.600 24.825 ;
        RECT 3.495 24.640 3.755 24.960 ;
        RECT 4.980 24.645 5.240 27.245 ;
        RECT 6.310 24.990 6.780 32.410 ;
        RECT 7.270 25.775 8.160 32.695 ;
        RECT 8.840 32.390 9.070 32.490 ;
        RECT 8.840 32.380 9.195 32.390 ;
        RECT 9.980 32.380 10.210 32.490 ;
        RECT 3.550 24.480 3.700 24.640 ;
        RECT 2.010 19.255 2.505 24.395 ;
        RECT 3.525 24.345 3.730 24.480 ;
        RECT 5.010 24.395 5.240 24.645 ;
        RECT 6.030 24.550 6.780 24.990 ;
        RECT 7.200 24.775 8.215 25.775 ;
        RECT 2.805 24.115 4.805 24.345 ;
        RECT 6.030 22.355 6.400 24.550 ;
        RECT 6.550 24.490 6.780 24.550 ;
        RECT 7.270 24.285 8.160 24.775 ;
        RECT 8.840 24.580 10.210 32.380 ;
        RECT 10.745 27.635 11.635 32.695 ;
        RECT 12.270 32.410 12.500 32.490 ;
        RECT 10.740 26.015 11.640 27.635 ;
        RECT 10.745 25.605 11.635 26.015 ;
        RECT 10.670 24.605 11.700 25.605 ;
        RECT 12.270 24.625 12.645 32.410 ;
        RECT 12.920 32.025 14.600 33.260 ;
        RECT 15.435 32.025 20.360 32.035 ;
        RECT 12.920 31.545 20.360 32.025 ;
        RECT 12.920 29.285 14.600 31.545 ;
        RECT 15.435 31.125 20.360 31.545 ;
        RECT 14.940 30.935 15.195 30.960 ;
        RECT 14.940 30.920 15.215 30.935 ;
        RECT 14.910 30.645 15.245 30.920 ;
        RECT 15.420 30.895 20.420 31.125 ;
        RECT 20.630 30.935 20.885 30.960 ;
        RECT 14.940 30.630 15.195 30.645 ;
        RECT 15.420 30.455 20.420 30.685 ;
        RECT 20.625 30.645 20.885 30.935 ;
        RECT 20.630 30.630 20.885 30.645 ;
        RECT 15.465 30.445 20.320 30.455 ;
        RECT 15.465 28.920 18.110 28.925 ;
        RECT 14.140 28.720 18.110 28.920 ;
        RECT 14.140 28.690 18.100 28.720 ;
        RECT 12.980 28.335 13.315 28.610 ;
        RECT 13.860 28.440 14.090 28.485 ;
        RECT 8.840 24.560 9.195 24.580 ;
        RECT 8.840 24.490 9.070 24.560 ;
        RECT 9.980 24.490 10.210 24.580 ;
        RECT 10.740 24.465 11.650 24.605 ;
        RECT 12.270 24.490 12.660 24.625 ;
        RECT 10.730 24.285 11.740 24.465 ;
        RECT 6.830 24.055 8.790 24.285 ;
        RECT 10.260 24.055 12.220 24.285 ;
        RECT 7.585 23.035 7.915 24.055 ;
        RECT 10.285 24.050 12.170 24.055 ;
        RECT 12.465 22.355 12.660 24.490 ;
        RECT 13.050 22.830 13.240 28.335 ;
        RECT 13.670 27.105 14.090 28.440 ;
        RECT 15.395 27.105 16.740 28.690 ;
        RECT 13.670 25.720 16.740 27.105 ;
        RECT 13.670 24.990 14.090 25.720 ;
        RECT 13.665 24.485 14.090 24.990 ;
        RECT 13.050 22.640 13.365 22.830 ;
        RECT 3.370 22.125 7.330 22.355 ;
        RECT 8.800 22.125 12.760 22.355 ;
        RECT 13.175 22.130 13.365 22.640 ;
        RECT 3.090 21.515 3.320 21.965 ;
        RECT 4.570 21.515 5.360 22.125 ;
        RECT 3.090 21.210 5.360 21.515 ;
        RECT 3.035 21.195 5.360 21.210 ;
        RECT 2.950 20.350 5.360 21.195 ;
        RECT 2.950 19.975 3.320 20.350 ;
        RECT 3.090 19.965 3.320 19.975 ;
        RECT 4.570 19.805 5.360 20.350 ;
        RECT 7.380 21.880 7.610 21.965 ;
        RECT 8.520 21.880 8.750 21.965 ;
        RECT 7.380 20.055 8.750 21.880 ;
        RECT 7.380 19.965 7.610 20.055 ;
        RECT 3.370 19.575 7.330 19.805 ;
        RECT 2.950 19.255 3.175 19.265 ;
        RECT 7.850 19.255 8.340 20.055 ;
        RECT 8.520 19.965 8.750 20.055 ;
        RECT 10.235 21.745 11.575 22.125 ;
        RECT 12.810 21.745 13.040 21.965 ;
        RECT 10.235 20.150 13.040 21.745 ;
        RECT 10.235 19.805 11.575 20.150 ;
        RECT 12.810 19.965 13.040 20.150 ;
        RECT 8.800 19.575 12.760 19.805 ;
        RECT 13.190 19.785 13.365 22.130 ;
        RECT 13.665 21.965 13.960 24.485 ;
        RECT 15.395 24.280 16.740 25.720 ;
        RECT 18.150 28.390 18.380 28.485 ;
        RECT 18.625 28.390 19.115 30.445 ;
        RECT 19.685 28.920 20.320 28.925 ;
        RECT 19.570 28.690 23.530 28.920 ;
        RECT 19.290 28.390 19.520 28.485 ;
        RECT 18.150 24.565 19.520 28.390 ;
        RECT 18.150 24.485 18.380 24.565 ;
        RECT 19.290 24.485 19.520 24.565 ;
        RECT 20.945 24.280 22.290 28.690 ;
        RECT 23.580 28.420 23.810 28.485 ;
        RECT 24.465 28.425 24.940 33.260 ;
        RECT 26.265 32.455 26.945 33.260 ;
        RECT 27.365 32.735 27.700 32.985 ;
        RECT 27.380 32.710 27.670 32.735 ;
        RECT 30.840 32.635 32.750 33.260 ;
        RECT 34.840 32.925 36.725 32.930 ;
        RECT 38.285 32.925 40.170 32.930 ;
        RECT 34.830 32.695 36.790 32.925 ;
        RECT 38.260 32.695 40.220 32.925 ;
        RECT 27.190 32.455 27.420 32.505 ;
        RECT 26.265 31.955 27.420 32.455 ;
        RECT 25.335 28.735 25.670 28.985 ;
        RECT 25.355 28.705 25.645 28.735 ;
        RECT 25.165 28.425 25.395 28.500 ;
        RECT 23.580 24.485 24.035 28.420 ;
        RECT 24.465 27.680 25.395 28.425 ;
        RECT 24.800 24.565 25.395 27.680 ;
        RECT 25.165 24.500 25.395 24.565 ;
        RECT 25.605 28.475 25.835 28.500 ;
        RECT 25.605 24.920 26.115 28.475 ;
        RECT 25.605 24.550 26.300 24.920 ;
        RECT 26.800 24.600 27.420 31.955 ;
        RECT 25.605 24.500 25.835 24.550 ;
        RECT 14.140 24.250 18.100 24.280 ;
        RECT 19.570 24.250 23.530 24.280 ;
        RECT 14.140 24.090 23.530 24.250 ;
        RECT 14.140 24.050 18.100 24.090 ;
        RECT 19.570 24.050 23.530 24.090 ;
        RECT 23.695 22.660 24.035 24.485 ;
        RECT 25.345 22.660 25.765 24.305 ;
        RECT 23.695 22.505 25.765 22.660 ;
        RECT 23.770 22.390 25.765 22.505 ;
        RECT 14.230 22.125 18.190 22.355 ;
        RECT 19.660 22.125 23.620 22.355 ;
        RECT 13.665 21.205 14.180 21.965 ;
        RECT 13.735 20.025 14.180 21.205 ;
        RECT 13.950 19.965 14.180 20.025 ;
        RECT 15.610 19.805 16.565 22.125 ;
        RECT 18.240 21.900 18.470 21.965 ;
        RECT 19.380 21.900 19.610 21.965 ;
        RECT 18.240 20.030 19.610 21.900 ;
        RECT 18.240 19.965 18.470 20.030 ;
        RECT 13.175 19.255 13.365 19.785 ;
        RECT 14.230 19.575 18.190 19.805 ;
        RECT 18.645 19.255 19.200 20.030 ;
        RECT 19.380 19.965 19.610 20.030 ;
        RECT 21.055 19.805 22.010 22.125 ;
        RECT 23.770 21.970 24.035 22.390 ;
        RECT 25.345 22.115 25.765 22.390 ;
        RECT 26.000 23.355 26.300 24.550 ;
        RECT 27.190 24.505 27.420 24.600 ;
        RECT 27.630 32.430 27.860 32.505 ;
        RECT 27.630 25.110 28.405 32.430 ;
        RECT 30.805 32.405 32.805 32.635 ;
        RECT 34.550 32.410 34.780 32.490 ;
        RECT 30.370 29.060 30.600 32.355 ;
        RECT 33.010 32.275 33.240 32.355 ;
        RECT 32.980 29.060 33.240 32.275 ;
        RECT 30.370 27.245 33.240 29.060 ;
        RECT 27.630 24.580 28.480 25.110 ;
        RECT 30.370 24.825 30.600 27.245 ;
        RECT 27.630 24.505 27.860 24.580 ;
        RECT 27.295 23.825 27.810 24.315 ;
        RECT 28.110 23.825 28.480 24.580 ;
        RECT 30.010 24.395 30.600 24.825 ;
        RECT 31.495 24.640 31.755 24.960 ;
        RECT 32.980 24.645 33.240 27.245 ;
        RECT 34.310 24.990 34.780 32.410 ;
        RECT 35.270 25.775 36.160 32.695 ;
        RECT 36.840 32.390 37.070 32.490 ;
        RECT 36.840 32.380 37.195 32.390 ;
        RECT 37.980 32.380 38.210 32.490 ;
        RECT 31.550 24.480 31.700 24.640 ;
        RECT 27.295 23.360 27.805 23.825 ;
        RECT 26.930 23.355 27.805 23.360 ;
        RECT 26.000 22.950 27.805 23.355 ;
        RECT 26.000 22.110 26.300 22.950 ;
        RECT 26.930 22.935 27.805 22.950 ;
        RECT 27.295 22.825 27.805 22.935 ;
        RECT 27.295 22.125 27.810 22.825 ;
        RECT 28.035 22.795 29.035 23.825 ;
        RECT 23.695 21.965 24.035 21.970 ;
        RECT 23.670 20.020 24.035 21.965 ;
        RECT 25.250 21.900 25.480 21.970 ;
        RECT 24.755 21.230 25.480 21.900 ;
        RECT 24.745 21.040 25.480 21.230 ;
        RECT 24.745 20.240 25.100 21.040 ;
        RECT 25.250 20.970 25.480 21.040 ;
        RECT 25.690 21.925 25.920 21.970 ;
        RECT 26.060 21.925 26.300 22.110 ;
        RECT 25.690 21.595 26.300 21.925 ;
        RECT 27.275 21.870 27.505 21.975 ;
        RECT 25.690 21.040 26.185 21.595 ;
        RECT 25.690 20.970 25.920 21.040 ;
        RECT 25.440 20.785 25.730 20.810 ;
        RECT 25.425 20.535 25.760 20.785 ;
        RECT 27.045 20.765 27.505 21.870 ;
        RECT 26.725 20.240 27.505 20.765 ;
        RECT 24.305 20.060 27.505 20.240 ;
        RECT 23.670 19.965 23.900 20.020 ;
        RECT 19.660 19.575 23.620 19.805 ;
        RECT 24.305 19.620 27.110 20.060 ;
        RECT 27.275 19.975 27.505 20.060 ;
        RECT 27.715 21.910 27.945 21.975 ;
        RECT 28.110 21.910 28.480 22.795 ;
        RECT 27.715 21.585 28.480 21.910 ;
        RECT 27.715 20.045 28.475 21.585 ;
        RECT 27.715 19.975 27.945 20.045 ;
        RECT 27.465 19.795 27.755 19.815 ;
        RECT 24.305 19.255 26.770 19.620 ;
        RECT 27.440 19.545 27.775 19.795 ;
        RECT 30.010 19.280 30.505 24.395 ;
        RECT 31.525 24.345 31.730 24.480 ;
        RECT 33.010 24.395 33.240 24.645 ;
        RECT 34.030 24.550 34.780 24.990 ;
        RECT 35.200 24.775 36.215 25.775 ;
        RECT 30.805 24.115 32.805 24.345 ;
        RECT 34.030 22.355 34.400 24.550 ;
        RECT 34.550 24.490 34.780 24.550 ;
        RECT 35.270 24.285 36.160 24.775 ;
        RECT 36.840 24.580 38.210 32.380 ;
        RECT 38.745 27.635 39.635 32.695 ;
        RECT 40.270 32.410 40.500 32.490 ;
        RECT 38.740 26.015 39.640 27.635 ;
        RECT 38.745 25.605 39.635 26.015 ;
        RECT 38.670 24.605 39.700 25.605 ;
        RECT 40.270 24.625 40.645 32.410 ;
        RECT 40.920 32.025 42.600 33.260 ;
        RECT 43.435 32.025 48.360 32.035 ;
        RECT 40.920 31.545 48.360 32.025 ;
        RECT 40.920 29.285 42.600 31.545 ;
        RECT 43.435 31.125 48.360 31.545 ;
        RECT 42.940 30.935 43.195 30.960 ;
        RECT 42.940 30.920 43.215 30.935 ;
        RECT 42.910 30.645 43.245 30.920 ;
        RECT 43.420 30.895 48.420 31.125 ;
        RECT 48.630 30.935 48.885 30.960 ;
        RECT 42.940 30.630 43.195 30.645 ;
        RECT 43.420 30.455 48.420 30.685 ;
        RECT 48.625 30.645 48.885 30.935 ;
        RECT 48.630 30.630 48.885 30.645 ;
        RECT 43.465 30.445 48.320 30.455 ;
        RECT 43.465 28.920 46.110 28.925 ;
        RECT 42.140 28.720 46.110 28.920 ;
        RECT 42.140 28.690 46.100 28.720 ;
        RECT 40.980 28.335 41.315 28.610 ;
        RECT 41.860 28.440 42.090 28.485 ;
        RECT 36.840 24.560 37.195 24.580 ;
        RECT 36.840 24.490 37.070 24.560 ;
        RECT 37.980 24.490 38.210 24.580 ;
        RECT 38.740 24.465 39.650 24.605 ;
        RECT 40.270 24.490 40.660 24.625 ;
        RECT 38.730 24.285 39.740 24.465 ;
        RECT 34.830 24.055 36.790 24.285 ;
        RECT 38.260 24.055 40.220 24.285 ;
        RECT 35.535 23.005 35.885 24.055 ;
        RECT 38.285 24.050 40.170 24.055 ;
        RECT 40.465 22.355 40.660 24.490 ;
        RECT 41.050 22.830 41.240 28.335 ;
        RECT 41.670 27.105 42.090 28.440 ;
        RECT 43.395 27.105 44.740 28.690 ;
        RECT 41.670 25.720 44.740 27.105 ;
        RECT 41.670 24.990 42.090 25.720 ;
        RECT 41.665 24.485 42.090 24.990 ;
        RECT 41.050 22.640 41.365 22.830 ;
        RECT 31.370 22.125 35.330 22.355 ;
        RECT 36.800 22.125 40.760 22.355 ;
        RECT 41.175 22.130 41.365 22.640 ;
        RECT 31.090 21.515 31.320 21.965 ;
        RECT 32.570 21.515 33.360 22.125 ;
        RECT 31.090 21.210 33.360 21.515 ;
        RECT 31.035 21.195 33.360 21.210 ;
        RECT 30.950 20.350 33.360 21.195 ;
        RECT 30.950 19.975 31.320 20.350 ;
        RECT 31.090 19.965 31.320 19.975 ;
        RECT 32.570 19.805 33.360 20.350 ;
        RECT 35.380 21.880 35.610 21.965 ;
        RECT 36.520 21.880 36.750 21.965 ;
        RECT 35.380 20.055 36.750 21.880 ;
        RECT 35.380 19.965 35.610 20.055 ;
        RECT 31.370 19.575 35.330 19.805 ;
        RECT 28.310 19.255 30.505 19.280 ;
        RECT 30.950 19.255 31.175 19.265 ;
        RECT 35.850 19.255 36.340 20.055 ;
        RECT 36.520 19.965 36.750 20.055 ;
        RECT 38.235 21.745 39.575 22.125 ;
        RECT 40.810 21.745 41.040 21.965 ;
        RECT 38.235 20.150 41.040 21.745 ;
        RECT 38.235 19.805 39.575 20.150 ;
        RECT 40.810 19.965 41.040 20.150 ;
        RECT 36.800 19.575 40.760 19.805 ;
        RECT 41.190 19.785 41.365 22.130 ;
        RECT 41.665 21.965 41.960 24.485 ;
        RECT 43.395 24.280 44.740 25.720 ;
        RECT 46.150 28.390 46.380 28.485 ;
        RECT 46.625 28.390 47.115 30.445 ;
        RECT 47.685 28.920 48.320 28.925 ;
        RECT 47.570 28.690 51.530 28.920 ;
        RECT 47.290 28.390 47.520 28.485 ;
        RECT 46.150 24.565 47.520 28.390 ;
        RECT 46.150 24.485 46.380 24.565 ;
        RECT 47.290 24.485 47.520 24.565 ;
        RECT 48.945 24.280 50.290 28.690 ;
        RECT 51.580 28.420 51.810 28.485 ;
        RECT 52.465 28.425 52.940 33.260 ;
        RECT 54.265 32.455 54.945 33.260 ;
        RECT 55.810 33.180 58.410 33.260 ;
        RECT 55.365 32.735 55.700 32.985 ;
        RECT 55.380 32.710 55.670 32.735 ;
        RECT 58.840 32.635 60.750 33.260 ;
        RECT 62.840 32.925 64.725 32.930 ;
        RECT 66.285 32.925 68.170 32.930 ;
        RECT 62.830 32.695 64.790 32.925 ;
        RECT 66.260 32.695 68.220 32.925 ;
        RECT 55.190 32.455 55.420 32.505 ;
        RECT 54.265 31.955 55.420 32.455 ;
        RECT 53.335 28.735 53.670 28.985 ;
        RECT 53.355 28.705 53.645 28.735 ;
        RECT 53.165 28.425 53.395 28.500 ;
        RECT 51.580 24.485 52.035 28.420 ;
        RECT 52.465 27.680 53.395 28.425 ;
        RECT 52.800 24.565 53.395 27.680 ;
        RECT 53.165 24.500 53.395 24.565 ;
        RECT 53.605 28.475 53.835 28.500 ;
        RECT 53.605 24.920 54.115 28.475 ;
        RECT 53.605 24.550 54.300 24.920 ;
        RECT 54.800 24.600 55.420 31.955 ;
        RECT 53.605 24.500 53.835 24.550 ;
        RECT 42.140 24.250 46.100 24.280 ;
        RECT 47.570 24.250 51.530 24.280 ;
        RECT 42.140 24.090 51.530 24.250 ;
        RECT 42.140 24.050 46.100 24.090 ;
        RECT 47.570 24.050 51.530 24.090 ;
        RECT 51.695 22.660 52.035 24.485 ;
        RECT 53.345 22.660 53.765 24.305 ;
        RECT 51.695 22.505 53.765 22.660 ;
        RECT 51.770 22.390 53.765 22.505 ;
        RECT 42.230 22.125 46.190 22.355 ;
        RECT 47.660 22.125 51.620 22.355 ;
        RECT 41.665 21.205 42.180 21.965 ;
        RECT 41.735 20.025 42.180 21.205 ;
        RECT 41.950 19.965 42.180 20.025 ;
        RECT 43.610 19.805 44.565 22.125 ;
        RECT 46.240 21.900 46.470 21.965 ;
        RECT 47.380 21.900 47.610 21.965 ;
        RECT 46.240 20.030 47.610 21.900 ;
        RECT 46.240 19.965 46.470 20.030 ;
        RECT 41.175 19.255 41.365 19.785 ;
        RECT 42.230 19.575 46.190 19.805 ;
        RECT 46.645 19.255 47.200 20.030 ;
        RECT 47.380 19.965 47.610 20.030 ;
        RECT 49.055 19.805 50.010 22.125 ;
        RECT 51.770 21.970 52.035 22.390 ;
        RECT 53.345 22.115 53.765 22.390 ;
        RECT 54.000 23.355 54.300 24.550 ;
        RECT 55.190 24.505 55.420 24.600 ;
        RECT 55.630 32.430 55.860 32.505 ;
        RECT 55.630 25.110 56.405 32.430 ;
        RECT 58.805 32.405 60.805 32.635 ;
        RECT 62.550 32.410 62.780 32.490 ;
        RECT 58.370 29.060 58.600 32.355 ;
        RECT 61.010 32.275 61.240 32.355 ;
        RECT 60.980 29.060 61.240 32.275 ;
        RECT 58.370 27.245 61.240 29.060 ;
        RECT 55.630 24.580 56.480 25.110 ;
        RECT 58.370 24.825 58.600 27.245 ;
        RECT 55.630 24.505 55.860 24.580 ;
        RECT 55.295 23.825 55.810 24.315 ;
        RECT 55.295 23.360 55.805 23.825 ;
        RECT 56.110 23.795 56.480 24.580 ;
        RECT 58.010 24.395 58.600 24.825 ;
        RECT 59.495 24.640 59.755 24.960 ;
        RECT 60.980 24.645 61.240 27.245 ;
        RECT 62.310 24.990 62.780 32.410 ;
        RECT 63.270 25.775 64.160 32.695 ;
        RECT 64.840 32.390 65.070 32.490 ;
        RECT 64.840 32.380 65.195 32.390 ;
        RECT 65.980 32.380 66.210 32.490 ;
        RECT 59.550 24.480 59.700 24.640 ;
        RECT 54.930 23.355 55.805 23.360 ;
        RECT 54.000 22.950 55.805 23.355 ;
        RECT 54.000 22.110 54.300 22.950 ;
        RECT 54.930 22.935 55.805 22.950 ;
        RECT 55.295 22.825 55.805 22.935 ;
        RECT 55.295 22.125 55.810 22.825 ;
        RECT 56.005 22.795 57.035 23.795 ;
        RECT 51.695 21.965 52.035 21.970 ;
        RECT 51.670 20.020 52.035 21.965 ;
        RECT 53.250 21.900 53.480 21.970 ;
        RECT 52.755 21.230 53.480 21.900 ;
        RECT 52.745 21.040 53.480 21.230 ;
        RECT 52.745 20.240 53.100 21.040 ;
        RECT 53.250 20.970 53.480 21.040 ;
        RECT 53.690 21.925 53.920 21.970 ;
        RECT 54.060 21.925 54.300 22.110 ;
        RECT 53.690 21.595 54.300 21.925 ;
        RECT 55.275 21.870 55.505 21.975 ;
        RECT 53.690 21.040 54.185 21.595 ;
        RECT 53.690 20.970 53.920 21.040 ;
        RECT 53.440 20.785 53.730 20.810 ;
        RECT 53.425 20.535 53.760 20.785 ;
        RECT 55.045 20.765 55.505 21.870 ;
        RECT 54.725 20.240 55.505 20.765 ;
        RECT 52.305 20.060 55.505 20.240 ;
        RECT 51.670 19.965 51.900 20.020 ;
        RECT 47.660 19.575 51.620 19.805 ;
        RECT 52.305 19.620 55.110 20.060 ;
        RECT 55.275 19.975 55.505 20.060 ;
        RECT 55.715 21.910 55.945 21.975 ;
        RECT 56.110 21.910 56.480 22.795 ;
        RECT 55.715 21.585 56.480 21.910 ;
        RECT 55.715 20.045 56.475 21.585 ;
        RECT 55.715 19.975 55.945 20.045 ;
        RECT 55.465 19.795 55.755 19.815 ;
        RECT 52.305 19.255 54.770 19.620 ;
        RECT 55.440 19.545 55.775 19.795 ;
        RECT 58.010 19.280 58.505 24.395 ;
        RECT 59.525 24.345 59.730 24.480 ;
        RECT 61.010 24.395 61.240 24.645 ;
        RECT 62.030 24.550 62.780 24.990 ;
        RECT 63.200 24.775 64.215 25.775 ;
        RECT 58.805 24.115 60.805 24.345 ;
        RECT 62.030 22.355 62.400 24.550 ;
        RECT 62.550 24.490 62.780 24.550 ;
        RECT 63.270 24.285 64.160 24.775 ;
        RECT 64.840 24.580 66.210 32.380 ;
        RECT 66.745 27.635 67.635 32.695 ;
        RECT 68.270 32.410 68.500 32.490 ;
        RECT 66.740 26.015 67.640 27.635 ;
        RECT 66.745 25.605 67.635 26.015 ;
        RECT 66.670 24.605 67.700 25.605 ;
        RECT 68.270 24.625 68.645 32.410 ;
        RECT 68.920 32.025 70.600 33.260 ;
        RECT 71.435 32.025 76.360 32.035 ;
        RECT 68.920 31.545 76.360 32.025 ;
        RECT 68.920 29.285 70.600 31.545 ;
        RECT 71.435 31.125 76.360 31.545 ;
        RECT 70.940 30.935 71.195 30.960 ;
        RECT 70.940 30.920 71.215 30.935 ;
        RECT 70.910 30.645 71.245 30.920 ;
        RECT 71.420 30.895 76.420 31.125 ;
        RECT 76.630 30.935 76.885 30.960 ;
        RECT 70.940 30.630 71.195 30.645 ;
        RECT 71.420 30.455 76.420 30.685 ;
        RECT 76.625 30.645 76.885 30.935 ;
        RECT 76.630 30.630 76.885 30.645 ;
        RECT 71.465 30.445 76.320 30.455 ;
        RECT 71.465 28.920 74.110 28.925 ;
        RECT 70.140 28.720 74.110 28.920 ;
        RECT 70.140 28.690 74.100 28.720 ;
        RECT 68.980 28.335 69.315 28.610 ;
        RECT 69.860 28.440 70.090 28.485 ;
        RECT 64.840 24.560 65.195 24.580 ;
        RECT 64.840 24.490 65.070 24.560 ;
        RECT 65.980 24.490 66.210 24.580 ;
        RECT 66.740 24.465 67.650 24.605 ;
        RECT 68.270 24.490 68.660 24.625 ;
        RECT 66.730 24.285 67.740 24.465 ;
        RECT 62.830 24.055 64.790 24.285 ;
        RECT 66.260 24.055 68.220 24.285 ;
        RECT 63.585 23.050 63.930 24.055 ;
        RECT 66.285 24.050 68.170 24.055 ;
        RECT 68.465 22.355 68.660 24.490 ;
        RECT 69.050 22.830 69.240 28.335 ;
        RECT 69.670 27.105 70.090 28.440 ;
        RECT 71.395 27.105 72.740 28.690 ;
        RECT 69.670 25.720 72.740 27.105 ;
        RECT 69.670 24.990 70.090 25.720 ;
        RECT 69.665 24.485 70.090 24.990 ;
        RECT 69.050 22.640 69.365 22.830 ;
        RECT 59.370 22.125 63.330 22.355 ;
        RECT 64.800 22.125 68.760 22.355 ;
        RECT 69.175 22.130 69.365 22.640 ;
        RECT 59.090 21.515 59.320 21.965 ;
        RECT 60.570 21.515 61.360 22.125 ;
        RECT 59.090 21.210 61.360 21.515 ;
        RECT 59.035 21.195 61.360 21.210 ;
        RECT 58.950 20.350 61.360 21.195 ;
        RECT 58.950 19.975 59.320 20.350 ;
        RECT 59.090 19.965 59.320 19.975 ;
        RECT 60.570 19.805 61.360 20.350 ;
        RECT 63.380 21.880 63.610 21.965 ;
        RECT 64.520 21.880 64.750 21.965 ;
        RECT 63.380 20.055 64.750 21.880 ;
        RECT 63.380 19.965 63.610 20.055 ;
        RECT 59.370 19.575 63.330 19.805 ;
        RECT 55.910 19.255 58.505 19.280 ;
        RECT 58.950 19.255 59.175 19.265 ;
        RECT 63.850 19.255 64.340 20.055 ;
        RECT 64.520 19.965 64.750 20.055 ;
        RECT 66.235 21.745 67.575 22.125 ;
        RECT 68.810 21.745 69.040 21.965 ;
        RECT 66.235 20.150 69.040 21.745 ;
        RECT 66.235 19.805 67.575 20.150 ;
        RECT 68.810 19.965 69.040 20.150 ;
        RECT 64.800 19.575 68.760 19.805 ;
        RECT 69.190 19.785 69.365 22.130 ;
        RECT 69.665 21.965 69.960 24.485 ;
        RECT 71.395 24.280 72.740 25.720 ;
        RECT 74.150 28.390 74.380 28.485 ;
        RECT 74.625 28.390 75.115 30.445 ;
        RECT 75.685 28.920 76.320 28.925 ;
        RECT 75.570 28.690 79.530 28.920 ;
        RECT 75.290 28.390 75.520 28.485 ;
        RECT 74.150 24.565 75.520 28.390 ;
        RECT 74.150 24.485 74.380 24.565 ;
        RECT 75.290 24.485 75.520 24.565 ;
        RECT 76.945 24.280 78.290 28.690 ;
        RECT 79.580 28.420 79.810 28.485 ;
        RECT 80.465 28.425 80.940 33.260 ;
        RECT 82.265 32.455 82.945 33.260 ;
        RECT 83.365 32.735 83.700 32.985 ;
        RECT 83.380 32.710 83.670 32.735 ;
        RECT 86.840 32.635 88.750 33.260 ;
        RECT 90.840 32.925 92.725 32.930 ;
        RECT 94.285 32.925 96.170 32.930 ;
        RECT 90.830 32.695 92.790 32.925 ;
        RECT 94.260 32.695 96.220 32.925 ;
        RECT 83.190 32.455 83.420 32.505 ;
        RECT 82.265 31.955 83.420 32.455 ;
        RECT 81.335 28.735 81.670 28.985 ;
        RECT 81.355 28.705 81.645 28.735 ;
        RECT 81.165 28.425 81.395 28.500 ;
        RECT 79.580 24.485 80.035 28.420 ;
        RECT 80.465 27.680 81.395 28.425 ;
        RECT 80.800 24.565 81.395 27.680 ;
        RECT 81.165 24.500 81.395 24.565 ;
        RECT 81.605 28.475 81.835 28.500 ;
        RECT 81.605 24.920 82.115 28.475 ;
        RECT 81.605 24.550 82.300 24.920 ;
        RECT 82.800 24.600 83.420 31.955 ;
        RECT 81.605 24.500 81.835 24.550 ;
        RECT 70.140 24.250 74.100 24.280 ;
        RECT 75.570 24.250 79.530 24.280 ;
        RECT 70.140 24.090 79.530 24.250 ;
        RECT 70.140 24.050 74.100 24.090 ;
        RECT 75.570 24.050 79.530 24.090 ;
        RECT 79.695 22.660 80.035 24.485 ;
        RECT 81.345 22.660 81.765 24.305 ;
        RECT 79.695 22.505 81.765 22.660 ;
        RECT 79.770 22.390 81.765 22.505 ;
        RECT 70.230 22.125 74.190 22.355 ;
        RECT 75.660 22.125 79.620 22.355 ;
        RECT 69.665 21.205 70.180 21.965 ;
        RECT 69.735 20.025 70.180 21.205 ;
        RECT 69.950 19.965 70.180 20.025 ;
        RECT 71.610 19.805 72.565 22.125 ;
        RECT 74.240 21.900 74.470 21.965 ;
        RECT 75.380 21.900 75.610 21.965 ;
        RECT 74.240 20.030 75.610 21.900 ;
        RECT 74.240 19.965 74.470 20.030 ;
        RECT 69.175 19.255 69.365 19.785 ;
        RECT 70.230 19.575 74.190 19.805 ;
        RECT 74.645 19.255 75.200 20.030 ;
        RECT 75.380 19.965 75.610 20.030 ;
        RECT 77.055 19.805 78.010 22.125 ;
        RECT 79.770 21.970 80.035 22.390 ;
        RECT 81.345 22.115 81.765 22.390 ;
        RECT 82.000 23.355 82.300 24.550 ;
        RECT 83.190 24.505 83.420 24.600 ;
        RECT 83.630 32.430 83.860 32.505 ;
        RECT 83.630 25.110 84.405 32.430 ;
        RECT 86.805 32.405 88.805 32.635 ;
        RECT 90.550 32.410 90.780 32.490 ;
        RECT 86.370 29.060 86.600 32.355 ;
        RECT 89.010 32.275 89.240 32.355 ;
        RECT 88.980 29.060 89.240 32.275 ;
        RECT 86.370 27.245 89.240 29.060 ;
        RECT 83.630 24.580 84.480 25.110 ;
        RECT 86.370 24.825 86.600 27.245 ;
        RECT 83.630 24.505 83.860 24.580 ;
        RECT 83.295 23.825 83.810 24.315 ;
        RECT 83.295 23.360 83.805 23.825 ;
        RECT 84.110 23.795 84.480 24.580 ;
        RECT 86.010 24.395 86.600 24.825 ;
        RECT 87.495 24.640 87.755 24.960 ;
        RECT 88.980 24.645 89.240 27.245 ;
        RECT 90.310 24.990 90.780 32.410 ;
        RECT 91.270 25.775 92.160 32.695 ;
        RECT 92.840 32.390 93.070 32.490 ;
        RECT 92.840 32.380 93.195 32.390 ;
        RECT 93.980 32.380 94.210 32.490 ;
        RECT 87.550 24.480 87.700 24.640 ;
        RECT 82.930 23.355 83.805 23.360 ;
        RECT 82.000 22.950 83.805 23.355 ;
        RECT 82.000 22.110 82.300 22.950 ;
        RECT 82.930 22.935 83.805 22.950 ;
        RECT 83.295 22.825 83.805 22.935 ;
        RECT 83.295 22.125 83.810 22.825 ;
        RECT 84.035 22.795 85.065 23.795 ;
        RECT 79.695 21.965 80.035 21.970 ;
        RECT 79.670 20.020 80.035 21.965 ;
        RECT 81.250 21.900 81.480 21.970 ;
        RECT 80.755 21.230 81.480 21.900 ;
        RECT 80.745 21.040 81.480 21.230 ;
        RECT 80.745 20.240 81.100 21.040 ;
        RECT 81.250 20.970 81.480 21.040 ;
        RECT 81.690 21.925 81.920 21.970 ;
        RECT 82.060 21.925 82.300 22.110 ;
        RECT 81.690 21.595 82.300 21.925 ;
        RECT 83.275 21.870 83.505 21.975 ;
        RECT 81.690 21.040 82.185 21.595 ;
        RECT 81.690 20.970 81.920 21.040 ;
        RECT 81.440 20.785 81.730 20.810 ;
        RECT 81.425 20.535 81.760 20.785 ;
        RECT 83.045 20.765 83.505 21.870 ;
        RECT 82.725 20.240 83.505 20.765 ;
        RECT 80.305 20.060 83.505 20.240 ;
        RECT 79.670 19.965 79.900 20.020 ;
        RECT 75.660 19.575 79.620 19.805 ;
        RECT 80.305 19.620 83.110 20.060 ;
        RECT 83.275 19.975 83.505 20.060 ;
        RECT 83.715 21.910 83.945 21.975 ;
        RECT 84.110 21.910 84.480 22.795 ;
        RECT 83.715 21.585 84.480 21.910 ;
        RECT 83.715 20.045 84.475 21.585 ;
        RECT 83.715 19.975 83.945 20.045 ;
        RECT 83.465 19.795 83.755 19.815 ;
        RECT 80.305 19.255 82.770 19.620 ;
        RECT 83.440 19.545 83.775 19.795 ;
        RECT 86.010 19.280 86.505 24.395 ;
        RECT 87.525 24.345 87.730 24.480 ;
        RECT 89.010 24.395 89.240 24.645 ;
        RECT 90.030 24.550 90.780 24.990 ;
        RECT 91.200 24.775 92.215 25.775 ;
        RECT 86.805 24.115 88.805 24.345 ;
        RECT 90.030 22.355 90.400 24.550 ;
        RECT 90.550 24.490 90.780 24.550 ;
        RECT 91.270 24.285 92.160 24.775 ;
        RECT 92.840 24.580 94.210 32.380 ;
        RECT 94.745 27.635 95.635 32.695 ;
        RECT 96.270 32.410 96.500 32.490 ;
        RECT 94.740 26.015 95.640 27.635 ;
        RECT 94.745 25.605 95.635 26.015 ;
        RECT 94.670 24.605 95.700 25.605 ;
        RECT 96.270 24.625 96.645 32.410 ;
        RECT 96.920 32.025 98.600 33.260 ;
        RECT 99.435 32.025 104.360 32.035 ;
        RECT 96.920 31.545 104.360 32.025 ;
        RECT 96.920 29.285 98.600 31.545 ;
        RECT 99.435 31.125 104.360 31.545 ;
        RECT 98.940 30.935 99.195 30.960 ;
        RECT 98.940 30.920 99.215 30.935 ;
        RECT 98.910 30.645 99.245 30.920 ;
        RECT 99.420 30.895 104.420 31.125 ;
        RECT 104.630 30.935 104.885 30.960 ;
        RECT 98.940 30.630 99.195 30.645 ;
        RECT 99.420 30.455 104.420 30.685 ;
        RECT 104.625 30.645 104.885 30.935 ;
        RECT 104.630 30.630 104.885 30.645 ;
        RECT 99.465 30.445 104.320 30.455 ;
        RECT 99.465 28.920 102.110 28.925 ;
        RECT 98.140 28.720 102.110 28.920 ;
        RECT 98.140 28.690 102.100 28.720 ;
        RECT 96.980 28.335 97.315 28.610 ;
        RECT 97.860 28.440 98.090 28.485 ;
        RECT 92.840 24.560 93.195 24.580 ;
        RECT 92.840 24.490 93.070 24.560 ;
        RECT 93.980 24.490 94.210 24.580 ;
        RECT 94.740 24.465 95.650 24.605 ;
        RECT 96.270 24.490 96.660 24.625 ;
        RECT 94.730 24.285 95.740 24.465 ;
        RECT 90.830 24.055 92.790 24.285 ;
        RECT 94.260 24.055 96.220 24.285 ;
        RECT 91.545 22.980 91.945 24.055 ;
        RECT 94.285 24.050 96.170 24.055 ;
        RECT 96.465 22.355 96.660 24.490 ;
        RECT 97.050 22.830 97.240 28.335 ;
        RECT 97.670 27.105 98.090 28.440 ;
        RECT 99.395 27.105 100.740 28.690 ;
        RECT 97.670 25.720 100.740 27.105 ;
        RECT 97.670 24.990 98.090 25.720 ;
        RECT 97.665 24.485 98.090 24.990 ;
        RECT 97.050 22.640 97.365 22.830 ;
        RECT 87.370 22.125 91.330 22.355 ;
        RECT 92.800 22.125 96.760 22.355 ;
        RECT 97.175 22.130 97.365 22.640 ;
        RECT 87.090 21.515 87.320 21.965 ;
        RECT 88.570 21.515 89.360 22.125 ;
        RECT 87.090 21.210 89.360 21.515 ;
        RECT 87.035 21.195 89.360 21.210 ;
        RECT 86.950 20.350 89.360 21.195 ;
        RECT 86.950 19.975 87.320 20.350 ;
        RECT 87.090 19.965 87.320 19.975 ;
        RECT 88.570 19.805 89.360 20.350 ;
        RECT 91.380 21.880 91.610 21.965 ;
        RECT 92.520 21.880 92.750 21.965 ;
        RECT 91.380 20.055 92.750 21.880 ;
        RECT 91.380 19.965 91.610 20.055 ;
        RECT 87.370 19.575 91.330 19.805 ;
        RECT 84.210 19.255 86.505 19.280 ;
        RECT 86.950 19.255 87.175 19.265 ;
        RECT 91.850 19.255 92.340 20.055 ;
        RECT 92.520 19.965 92.750 20.055 ;
        RECT 94.235 21.745 95.575 22.125 ;
        RECT 96.810 21.745 97.040 21.965 ;
        RECT 94.235 20.150 97.040 21.745 ;
        RECT 94.235 19.805 95.575 20.150 ;
        RECT 96.810 19.965 97.040 20.150 ;
        RECT 92.800 19.575 96.760 19.805 ;
        RECT 97.190 19.785 97.365 22.130 ;
        RECT 97.665 21.965 97.960 24.485 ;
        RECT 99.395 24.280 100.740 25.720 ;
        RECT 102.150 28.390 102.380 28.485 ;
        RECT 102.625 28.390 103.115 30.445 ;
        RECT 103.685 28.920 104.320 28.925 ;
        RECT 103.570 28.690 107.530 28.920 ;
        RECT 103.290 28.390 103.520 28.485 ;
        RECT 102.150 24.565 103.520 28.390 ;
        RECT 102.150 24.485 102.380 24.565 ;
        RECT 103.290 24.485 103.520 24.565 ;
        RECT 104.945 24.280 106.290 28.690 ;
        RECT 107.580 28.420 107.810 28.485 ;
        RECT 108.465 28.425 108.940 33.260 ;
        RECT 110.265 32.455 110.945 33.260 ;
        RECT 111.365 32.735 111.700 32.985 ;
        RECT 111.380 32.710 111.670 32.735 ;
        RECT 114.840 32.635 116.750 33.260 ;
        RECT 118.840 32.925 120.725 32.930 ;
        RECT 122.285 32.925 124.170 32.930 ;
        RECT 118.830 32.695 120.790 32.925 ;
        RECT 122.260 32.695 124.220 32.925 ;
        RECT 111.190 32.455 111.420 32.505 ;
        RECT 110.265 31.955 111.420 32.455 ;
        RECT 109.335 28.735 109.670 28.985 ;
        RECT 109.355 28.705 109.645 28.735 ;
        RECT 109.165 28.425 109.395 28.500 ;
        RECT 107.580 24.485 108.035 28.420 ;
        RECT 108.465 27.680 109.395 28.425 ;
        RECT 108.800 24.565 109.395 27.680 ;
        RECT 109.165 24.500 109.395 24.565 ;
        RECT 109.605 28.475 109.835 28.500 ;
        RECT 109.605 24.920 110.115 28.475 ;
        RECT 109.605 24.550 110.300 24.920 ;
        RECT 110.800 24.600 111.420 31.955 ;
        RECT 109.605 24.500 109.835 24.550 ;
        RECT 98.140 24.250 102.100 24.280 ;
        RECT 103.570 24.250 107.530 24.280 ;
        RECT 98.140 24.090 107.530 24.250 ;
        RECT 98.140 24.050 102.100 24.090 ;
        RECT 103.570 24.050 107.530 24.090 ;
        RECT 107.695 22.660 108.035 24.485 ;
        RECT 109.345 22.660 109.765 24.305 ;
        RECT 107.695 22.505 109.765 22.660 ;
        RECT 107.770 22.390 109.765 22.505 ;
        RECT 98.230 22.125 102.190 22.355 ;
        RECT 103.660 22.125 107.620 22.355 ;
        RECT 97.665 21.205 98.180 21.965 ;
        RECT 97.735 20.025 98.180 21.205 ;
        RECT 97.950 19.965 98.180 20.025 ;
        RECT 99.610 19.805 100.565 22.125 ;
        RECT 102.240 21.900 102.470 21.965 ;
        RECT 103.380 21.900 103.610 21.965 ;
        RECT 102.240 20.030 103.610 21.900 ;
        RECT 102.240 19.965 102.470 20.030 ;
        RECT 97.175 19.255 97.365 19.785 ;
        RECT 98.230 19.575 102.190 19.805 ;
        RECT 102.645 19.255 103.200 20.030 ;
        RECT 103.380 19.965 103.610 20.030 ;
        RECT 105.055 19.805 106.010 22.125 ;
        RECT 107.770 21.970 108.035 22.390 ;
        RECT 109.345 22.115 109.765 22.390 ;
        RECT 110.000 23.355 110.300 24.550 ;
        RECT 111.190 24.505 111.420 24.600 ;
        RECT 111.630 32.430 111.860 32.505 ;
        RECT 111.630 25.110 112.405 32.430 ;
        RECT 114.805 32.405 116.805 32.635 ;
        RECT 118.550 32.410 118.780 32.490 ;
        RECT 114.370 29.060 114.600 32.355 ;
        RECT 117.010 32.275 117.240 32.355 ;
        RECT 116.980 29.060 117.240 32.275 ;
        RECT 114.370 27.245 117.240 29.060 ;
        RECT 111.630 24.580 112.480 25.110 ;
        RECT 114.370 24.825 114.600 27.245 ;
        RECT 111.630 24.505 111.860 24.580 ;
        RECT 111.295 23.825 111.810 24.315 ;
        RECT 111.295 23.360 111.805 23.825 ;
        RECT 112.110 23.795 112.480 24.580 ;
        RECT 114.010 24.395 114.600 24.825 ;
        RECT 115.495 24.640 115.755 24.960 ;
        RECT 116.980 24.645 117.240 27.245 ;
        RECT 118.310 24.990 118.780 32.410 ;
        RECT 119.270 25.775 120.160 32.695 ;
        RECT 120.840 32.390 121.070 32.490 ;
        RECT 120.840 32.380 121.195 32.390 ;
        RECT 121.980 32.380 122.210 32.490 ;
        RECT 115.550 24.480 115.700 24.640 ;
        RECT 110.930 23.355 111.805 23.360 ;
        RECT 110.000 22.950 111.805 23.355 ;
        RECT 110.000 22.110 110.300 22.950 ;
        RECT 110.930 22.935 111.805 22.950 ;
        RECT 111.295 22.825 111.805 22.935 ;
        RECT 111.295 22.125 111.810 22.825 ;
        RECT 112.005 22.795 113.035 23.795 ;
        RECT 107.695 21.965 108.035 21.970 ;
        RECT 107.670 20.020 108.035 21.965 ;
        RECT 109.250 21.900 109.480 21.970 ;
        RECT 108.755 21.230 109.480 21.900 ;
        RECT 108.745 21.040 109.480 21.230 ;
        RECT 108.745 20.240 109.100 21.040 ;
        RECT 109.250 20.970 109.480 21.040 ;
        RECT 109.690 21.925 109.920 21.970 ;
        RECT 110.060 21.925 110.300 22.110 ;
        RECT 109.690 21.595 110.300 21.925 ;
        RECT 111.275 21.870 111.505 21.975 ;
        RECT 109.690 21.040 110.185 21.595 ;
        RECT 109.690 20.970 109.920 21.040 ;
        RECT 109.440 20.785 109.730 20.810 ;
        RECT 109.425 20.535 109.760 20.785 ;
        RECT 111.045 20.765 111.505 21.870 ;
        RECT 110.725 20.240 111.505 20.765 ;
        RECT 108.305 20.060 111.505 20.240 ;
        RECT 107.670 19.965 107.900 20.020 ;
        RECT 103.660 19.575 107.620 19.805 ;
        RECT 108.305 19.620 111.110 20.060 ;
        RECT 111.275 19.975 111.505 20.060 ;
        RECT 111.715 21.910 111.945 21.975 ;
        RECT 112.110 21.910 112.480 22.795 ;
        RECT 111.715 21.585 112.480 21.910 ;
        RECT 111.715 20.045 112.475 21.585 ;
        RECT 111.715 19.975 111.945 20.045 ;
        RECT 111.465 19.795 111.755 19.815 ;
        RECT 108.305 19.255 110.770 19.620 ;
        RECT 111.440 19.545 111.775 19.795 ;
        RECT 114.010 19.255 114.505 24.395 ;
        RECT 115.525 24.345 115.730 24.480 ;
        RECT 117.010 24.395 117.240 24.645 ;
        RECT 118.030 24.550 118.780 24.990 ;
        RECT 119.200 24.775 120.215 25.775 ;
        RECT 114.805 24.115 116.805 24.345 ;
        RECT 118.030 22.355 118.400 24.550 ;
        RECT 118.550 24.490 118.780 24.550 ;
        RECT 119.270 24.285 120.160 24.775 ;
        RECT 120.840 24.580 122.210 32.380 ;
        RECT 122.745 27.635 123.635 32.695 ;
        RECT 124.270 32.410 124.500 32.490 ;
        RECT 122.740 26.015 123.640 27.635 ;
        RECT 122.745 25.605 123.635 26.015 ;
        RECT 122.670 24.605 123.700 25.605 ;
        RECT 124.270 24.625 124.645 32.410 ;
        RECT 124.920 32.025 126.600 33.260 ;
        RECT 127.435 32.025 132.360 32.035 ;
        RECT 124.920 31.545 132.360 32.025 ;
        RECT 124.920 29.285 126.600 31.545 ;
        RECT 127.435 31.125 132.360 31.545 ;
        RECT 126.940 30.935 127.195 30.960 ;
        RECT 126.940 30.920 127.215 30.935 ;
        RECT 126.910 30.645 127.245 30.920 ;
        RECT 127.420 30.895 132.420 31.125 ;
        RECT 132.630 30.935 132.885 30.960 ;
        RECT 126.940 30.630 127.195 30.645 ;
        RECT 127.420 30.455 132.420 30.685 ;
        RECT 132.625 30.645 132.885 30.935 ;
        RECT 132.630 30.630 132.885 30.645 ;
        RECT 127.465 30.445 132.320 30.455 ;
        RECT 127.465 28.920 130.110 28.925 ;
        RECT 126.140 28.720 130.110 28.920 ;
        RECT 126.140 28.690 130.100 28.720 ;
        RECT 124.980 28.335 125.315 28.610 ;
        RECT 125.860 28.440 126.090 28.485 ;
        RECT 120.840 24.560 121.195 24.580 ;
        RECT 120.840 24.490 121.070 24.560 ;
        RECT 121.980 24.490 122.210 24.580 ;
        RECT 122.740 24.465 123.650 24.605 ;
        RECT 124.270 24.490 124.660 24.625 ;
        RECT 122.730 24.285 123.740 24.465 ;
        RECT 118.830 24.055 120.790 24.285 ;
        RECT 122.260 24.055 124.220 24.285 ;
        RECT 119.580 23.115 119.865 24.055 ;
        RECT 122.285 24.050 124.170 24.055 ;
        RECT 124.465 22.355 124.660 24.490 ;
        RECT 125.050 22.830 125.240 28.335 ;
        RECT 125.670 27.105 126.090 28.440 ;
        RECT 127.395 27.105 128.740 28.690 ;
        RECT 125.670 25.720 128.740 27.105 ;
        RECT 125.670 24.990 126.090 25.720 ;
        RECT 125.665 24.485 126.090 24.990 ;
        RECT 125.050 22.640 125.365 22.830 ;
        RECT 115.370 22.125 119.330 22.355 ;
        RECT 120.800 22.125 124.760 22.355 ;
        RECT 125.175 22.130 125.365 22.640 ;
        RECT 115.090 21.515 115.320 21.965 ;
        RECT 116.570 21.515 117.360 22.125 ;
        RECT 115.090 21.210 117.360 21.515 ;
        RECT 115.035 21.195 117.360 21.210 ;
        RECT 114.950 20.350 117.360 21.195 ;
        RECT 114.950 19.975 115.320 20.350 ;
        RECT 115.090 19.965 115.320 19.975 ;
        RECT 116.570 19.805 117.360 20.350 ;
        RECT 119.380 21.880 119.610 21.965 ;
        RECT 120.520 21.880 120.750 21.965 ;
        RECT 119.380 20.055 120.750 21.880 ;
        RECT 119.380 19.965 119.610 20.055 ;
        RECT 115.370 19.575 119.330 19.805 ;
        RECT 114.950 19.255 115.175 19.265 ;
        RECT 119.850 19.255 120.340 20.055 ;
        RECT 120.520 19.965 120.750 20.055 ;
        RECT 122.235 21.745 123.575 22.125 ;
        RECT 124.810 21.745 125.040 21.965 ;
        RECT 122.235 20.150 125.040 21.745 ;
        RECT 122.235 19.805 123.575 20.150 ;
        RECT 124.810 19.965 125.040 20.150 ;
        RECT 120.800 19.575 124.760 19.805 ;
        RECT 125.190 19.785 125.365 22.130 ;
        RECT 125.665 21.965 125.960 24.485 ;
        RECT 127.395 24.280 128.740 25.720 ;
        RECT 130.150 28.390 130.380 28.485 ;
        RECT 130.625 28.390 131.115 30.445 ;
        RECT 131.685 28.920 132.320 28.925 ;
        RECT 131.570 28.690 135.530 28.920 ;
        RECT 131.290 28.390 131.520 28.485 ;
        RECT 130.150 24.565 131.520 28.390 ;
        RECT 130.150 24.485 130.380 24.565 ;
        RECT 131.290 24.485 131.520 24.565 ;
        RECT 132.945 24.280 134.290 28.690 ;
        RECT 135.580 28.420 135.810 28.485 ;
        RECT 136.465 28.425 136.940 33.260 ;
        RECT 138.265 32.455 138.945 33.260 ;
        RECT 139.365 32.735 139.700 32.985 ;
        RECT 139.380 32.710 139.670 32.735 ;
        RECT 139.190 32.455 139.420 32.505 ;
        RECT 138.265 31.955 139.420 32.455 ;
        RECT 137.335 28.735 137.670 28.985 ;
        RECT 137.355 28.705 137.645 28.735 ;
        RECT 137.165 28.425 137.395 28.500 ;
        RECT 135.580 24.485 136.035 28.420 ;
        RECT 136.465 27.680 137.395 28.425 ;
        RECT 136.800 24.565 137.395 27.680 ;
        RECT 137.165 24.500 137.395 24.565 ;
        RECT 137.605 28.475 137.835 28.500 ;
        RECT 137.605 24.920 138.115 28.475 ;
        RECT 137.605 24.550 138.300 24.920 ;
        RECT 138.800 24.600 139.420 31.955 ;
        RECT 137.605 24.500 137.835 24.550 ;
        RECT 126.140 24.250 130.100 24.280 ;
        RECT 131.570 24.250 135.530 24.280 ;
        RECT 126.140 24.090 135.530 24.250 ;
        RECT 126.140 24.050 130.100 24.090 ;
        RECT 131.570 24.050 135.530 24.090 ;
        RECT 135.695 22.660 136.035 24.485 ;
        RECT 137.345 22.660 137.765 24.305 ;
        RECT 135.695 22.505 137.765 22.660 ;
        RECT 135.770 22.390 137.765 22.505 ;
        RECT 126.230 22.125 130.190 22.355 ;
        RECT 131.660 22.125 135.620 22.355 ;
        RECT 125.665 21.205 126.180 21.965 ;
        RECT 125.735 20.025 126.180 21.205 ;
        RECT 125.950 19.965 126.180 20.025 ;
        RECT 127.610 19.805 128.565 22.125 ;
        RECT 130.240 21.900 130.470 21.965 ;
        RECT 131.380 21.900 131.610 21.965 ;
        RECT 130.240 20.030 131.610 21.900 ;
        RECT 130.240 19.965 130.470 20.030 ;
        RECT 125.175 19.255 125.365 19.785 ;
        RECT 126.230 19.575 130.190 19.805 ;
        RECT 130.645 19.255 131.200 20.030 ;
        RECT 131.380 19.965 131.610 20.030 ;
        RECT 133.055 19.805 134.010 22.125 ;
        RECT 135.770 21.970 136.035 22.390 ;
        RECT 137.345 22.115 137.765 22.390 ;
        RECT 138.000 23.355 138.300 24.550 ;
        RECT 139.190 24.505 139.420 24.600 ;
        RECT 139.630 32.430 139.860 32.505 ;
        RECT 139.630 25.110 140.405 32.430 ;
        RECT 139.630 24.580 140.480 25.110 ;
        RECT 139.630 24.505 139.860 24.580 ;
        RECT 139.295 23.825 139.810 24.315 ;
        RECT 139.295 23.360 139.805 23.825 ;
        RECT 140.110 23.795 140.480 24.580 ;
        RECT 138.930 23.355 139.805 23.360 ;
        RECT 138.000 22.950 139.805 23.355 ;
        RECT 138.000 22.110 138.300 22.950 ;
        RECT 138.930 22.935 139.805 22.950 ;
        RECT 139.295 22.825 139.805 22.935 ;
        RECT 139.295 22.125 139.810 22.825 ;
        RECT 140.035 22.795 141.065 23.795 ;
        RECT 135.695 21.965 136.035 21.970 ;
        RECT 135.670 20.020 136.035 21.965 ;
        RECT 137.250 21.900 137.480 21.970 ;
        RECT 136.755 21.230 137.480 21.900 ;
        RECT 136.745 21.040 137.480 21.230 ;
        RECT 136.745 20.240 137.100 21.040 ;
        RECT 137.250 20.970 137.480 21.040 ;
        RECT 137.690 21.925 137.920 21.970 ;
        RECT 138.060 21.925 138.300 22.110 ;
        RECT 137.690 21.595 138.300 21.925 ;
        RECT 139.275 21.870 139.505 21.975 ;
        RECT 137.690 21.040 138.185 21.595 ;
        RECT 137.690 20.970 137.920 21.040 ;
        RECT 137.440 20.785 137.730 20.810 ;
        RECT 137.425 20.535 137.760 20.785 ;
        RECT 139.045 20.765 139.505 21.870 ;
        RECT 138.725 20.240 139.505 20.765 ;
        RECT 136.305 20.060 139.505 20.240 ;
        RECT 135.670 19.965 135.900 20.020 ;
        RECT 131.660 19.575 135.620 19.805 ;
        RECT 136.305 19.620 139.110 20.060 ;
        RECT 139.275 19.975 139.505 20.060 ;
        RECT 139.715 21.910 139.945 21.975 ;
        RECT 140.110 21.910 140.480 22.795 ;
        RECT 139.715 21.585 140.480 21.910 ;
        RECT 139.715 20.045 140.475 21.585 ;
        RECT 139.715 19.975 139.945 20.045 ;
        RECT 139.465 19.795 139.755 19.815 ;
        RECT 136.305 19.255 138.770 19.620 ;
        RECT 139.440 19.545 139.775 19.795 ;
        RECT 1.895 18.380 112.500 19.255 ;
        RECT 113.895 18.380 140.500 19.255 ;
        RECT 28.210 17.960 31.110 17.980 ;
        RECT 55.810 17.960 58.310 17.980 ;
        RECT 69.265 17.960 70.205 17.985 ;
        RECT 84.110 17.960 86.610 17.980 ;
        RECT 1.870 17.280 112.345 17.960 ;
        RECT 1.870 17.260 28.345 17.280 ;
        RECT 29.870 17.260 56.345 17.280 ;
        RECT 57.870 17.260 84.345 17.280 ;
        RECT 85.870 17.260 112.345 17.280 ;
        RECT 113.870 17.260 140.345 17.960 ;
        RECT 2.840 16.635 4.750 17.260 ;
        RECT 6.840 16.925 8.725 16.930 ;
        RECT 10.285 16.925 12.170 16.930 ;
        RECT 6.830 16.695 8.790 16.925 ;
        RECT 10.260 16.695 12.220 16.925 ;
        RECT 2.805 16.405 4.805 16.635 ;
        RECT 6.550 16.410 6.780 16.490 ;
        RECT 2.370 13.060 2.600 16.355 ;
        RECT 5.010 16.275 5.240 16.355 ;
        RECT 4.980 13.060 5.240 16.275 ;
        RECT 2.370 11.245 5.240 13.060 ;
        RECT 2.370 8.825 2.600 11.245 ;
        RECT 2.010 8.395 2.600 8.825 ;
        RECT 3.495 8.640 3.755 8.960 ;
        RECT 4.980 8.645 5.240 11.245 ;
        RECT 6.310 8.990 6.780 16.410 ;
        RECT 7.270 9.775 8.160 16.695 ;
        RECT 8.840 16.390 9.070 16.490 ;
        RECT 8.840 16.380 9.195 16.390 ;
        RECT 9.980 16.380 10.210 16.490 ;
        RECT 3.550 8.480 3.700 8.640 ;
        RECT 2.010 3.255 2.505 8.395 ;
        RECT 3.525 8.345 3.730 8.480 ;
        RECT 5.010 8.395 5.240 8.645 ;
        RECT 6.030 8.550 6.780 8.990 ;
        RECT 7.200 8.775 8.215 9.775 ;
        RECT 2.805 8.115 4.805 8.345 ;
        RECT 6.030 6.355 6.400 8.550 ;
        RECT 6.550 8.490 6.780 8.550 ;
        RECT 7.270 8.285 8.160 8.775 ;
        RECT 8.840 8.580 10.210 16.380 ;
        RECT 10.745 11.635 11.635 16.695 ;
        RECT 12.270 16.410 12.500 16.490 ;
        RECT 10.740 10.015 11.640 11.635 ;
        RECT 10.745 9.605 11.635 10.015 ;
        RECT 10.670 8.605 11.700 9.605 ;
        RECT 12.270 8.625 12.645 16.410 ;
        RECT 12.920 16.025 14.600 17.260 ;
        RECT 15.435 16.025 20.360 16.035 ;
        RECT 12.920 15.545 20.360 16.025 ;
        RECT 12.920 13.285 14.600 15.545 ;
        RECT 15.435 15.125 20.360 15.545 ;
        RECT 14.940 14.935 15.195 14.960 ;
        RECT 14.940 14.920 15.215 14.935 ;
        RECT 14.910 14.645 15.245 14.920 ;
        RECT 15.420 14.895 20.420 15.125 ;
        RECT 20.630 14.935 20.885 14.960 ;
        RECT 14.940 14.630 15.195 14.645 ;
        RECT 15.420 14.455 20.420 14.685 ;
        RECT 20.625 14.645 20.885 14.935 ;
        RECT 20.630 14.630 20.885 14.645 ;
        RECT 15.465 14.445 20.320 14.455 ;
        RECT 15.465 12.920 18.110 12.925 ;
        RECT 14.140 12.720 18.110 12.920 ;
        RECT 14.140 12.690 18.100 12.720 ;
        RECT 12.980 12.335 13.315 12.610 ;
        RECT 13.860 12.440 14.090 12.485 ;
        RECT 8.840 8.560 9.195 8.580 ;
        RECT 8.840 8.490 9.070 8.560 ;
        RECT 9.980 8.490 10.210 8.580 ;
        RECT 10.740 8.465 11.650 8.605 ;
        RECT 12.270 8.490 12.660 8.625 ;
        RECT 10.730 8.285 11.740 8.465 ;
        RECT 6.830 8.055 8.790 8.285 ;
        RECT 10.260 8.055 12.220 8.285 ;
        RECT 7.550 7.085 7.880 8.055 ;
        RECT 10.285 8.050 12.170 8.055 ;
        RECT 12.465 6.355 12.660 8.490 ;
        RECT 13.050 6.830 13.240 12.335 ;
        RECT 13.670 11.105 14.090 12.440 ;
        RECT 15.395 11.105 16.740 12.690 ;
        RECT 13.670 9.720 16.740 11.105 ;
        RECT 13.670 8.990 14.090 9.720 ;
        RECT 13.665 8.485 14.090 8.990 ;
        RECT 13.050 6.640 13.365 6.830 ;
        RECT 3.370 6.125 7.330 6.355 ;
        RECT 8.800 6.125 12.760 6.355 ;
        RECT 13.175 6.130 13.365 6.640 ;
        RECT 3.090 5.515 3.320 5.965 ;
        RECT 4.570 5.515 5.360 6.125 ;
        RECT 3.090 5.210 5.360 5.515 ;
        RECT 3.035 5.195 5.360 5.210 ;
        RECT 2.950 4.350 5.360 5.195 ;
        RECT 2.950 3.975 3.320 4.350 ;
        RECT 3.090 3.965 3.320 3.975 ;
        RECT 4.570 3.805 5.360 4.350 ;
        RECT 7.380 5.880 7.610 5.965 ;
        RECT 8.520 5.880 8.750 5.965 ;
        RECT 7.380 4.055 8.750 5.880 ;
        RECT 7.380 3.965 7.610 4.055 ;
        RECT 3.370 3.575 7.330 3.805 ;
        RECT 2.950 3.255 3.175 3.265 ;
        RECT 7.850 3.255 8.340 4.055 ;
        RECT 8.520 3.965 8.750 4.055 ;
        RECT 10.235 5.745 11.575 6.125 ;
        RECT 12.810 5.745 13.040 5.965 ;
        RECT 10.235 4.150 13.040 5.745 ;
        RECT 10.235 3.805 11.575 4.150 ;
        RECT 12.810 3.965 13.040 4.150 ;
        RECT 8.800 3.575 12.760 3.805 ;
        RECT 13.190 3.785 13.365 6.130 ;
        RECT 13.665 5.965 13.960 8.485 ;
        RECT 15.395 8.280 16.740 9.720 ;
        RECT 18.150 12.390 18.380 12.485 ;
        RECT 18.625 12.390 19.115 14.445 ;
        RECT 19.685 12.920 20.320 12.925 ;
        RECT 19.570 12.690 23.530 12.920 ;
        RECT 19.290 12.390 19.520 12.485 ;
        RECT 18.150 8.565 19.520 12.390 ;
        RECT 18.150 8.485 18.380 8.565 ;
        RECT 19.290 8.485 19.520 8.565 ;
        RECT 20.945 8.280 22.290 12.690 ;
        RECT 23.580 12.420 23.810 12.485 ;
        RECT 24.465 12.425 24.940 17.260 ;
        RECT 26.265 16.455 26.945 17.260 ;
        RECT 27.365 16.735 27.700 16.985 ;
        RECT 27.380 16.710 27.670 16.735 ;
        RECT 30.840 16.635 32.750 17.260 ;
        RECT 34.840 16.925 36.725 16.930 ;
        RECT 38.285 16.925 40.170 16.930 ;
        RECT 34.830 16.695 36.790 16.925 ;
        RECT 38.260 16.695 40.220 16.925 ;
        RECT 27.190 16.455 27.420 16.505 ;
        RECT 26.265 15.955 27.420 16.455 ;
        RECT 25.335 12.735 25.670 12.985 ;
        RECT 25.355 12.705 25.645 12.735 ;
        RECT 25.165 12.425 25.395 12.500 ;
        RECT 23.580 8.485 24.035 12.420 ;
        RECT 24.465 11.680 25.395 12.425 ;
        RECT 24.800 8.565 25.395 11.680 ;
        RECT 25.165 8.500 25.395 8.565 ;
        RECT 25.605 12.475 25.835 12.500 ;
        RECT 25.605 8.920 26.115 12.475 ;
        RECT 25.605 8.550 26.300 8.920 ;
        RECT 26.800 8.600 27.420 15.955 ;
        RECT 25.605 8.500 25.835 8.550 ;
        RECT 14.140 8.250 18.100 8.280 ;
        RECT 19.570 8.250 23.530 8.280 ;
        RECT 14.140 8.090 23.530 8.250 ;
        RECT 14.140 8.050 18.100 8.090 ;
        RECT 19.570 8.050 23.530 8.090 ;
        RECT 23.695 6.660 24.035 8.485 ;
        RECT 25.345 6.660 25.765 8.305 ;
        RECT 23.695 6.505 25.765 6.660 ;
        RECT 23.770 6.390 25.765 6.505 ;
        RECT 14.230 6.125 18.190 6.355 ;
        RECT 19.660 6.125 23.620 6.355 ;
        RECT 13.665 5.205 14.180 5.965 ;
        RECT 13.735 4.025 14.180 5.205 ;
        RECT 13.950 3.965 14.180 4.025 ;
        RECT 15.610 3.805 16.565 6.125 ;
        RECT 18.240 5.900 18.470 5.965 ;
        RECT 19.380 5.900 19.610 5.965 ;
        RECT 18.240 4.030 19.610 5.900 ;
        RECT 18.240 3.965 18.470 4.030 ;
        RECT 13.175 3.255 13.365 3.785 ;
        RECT 14.230 3.575 18.190 3.805 ;
        RECT 18.645 3.255 19.200 4.030 ;
        RECT 19.380 3.965 19.610 4.030 ;
        RECT 21.055 3.805 22.010 6.125 ;
        RECT 23.770 5.970 24.035 6.390 ;
        RECT 25.345 6.115 25.765 6.390 ;
        RECT 26.000 7.355 26.300 8.550 ;
        RECT 27.190 8.505 27.420 8.600 ;
        RECT 27.630 16.430 27.860 16.505 ;
        RECT 27.630 9.110 28.405 16.430 ;
        RECT 30.805 16.405 32.805 16.635 ;
        RECT 34.550 16.410 34.780 16.490 ;
        RECT 30.370 13.060 30.600 16.355 ;
        RECT 33.010 16.275 33.240 16.355 ;
        RECT 32.980 13.060 33.240 16.275 ;
        RECT 30.370 11.245 33.240 13.060 ;
        RECT 27.630 8.580 28.480 9.110 ;
        RECT 30.370 8.825 30.600 11.245 ;
        RECT 27.630 8.505 27.860 8.580 ;
        RECT 27.295 7.825 27.810 8.315 ;
        RECT 28.110 7.825 28.480 8.580 ;
        RECT 30.010 8.395 30.600 8.825 ;
        RECT 31.495 8.640 31.755 8.960 ;
        RECT 32.980 8.645 33.240 11.245 ;
        RECT 34.310 8.990 34.780 16.410 ;
        RECT 35.270 9.775 36.160 16.695 ;
        RECT 36.840 16.390 37.070 16.490 ;
        RECT 36.840 16.380 37.195 16.390 ;
        RECT 37.980 16.380 38.210 16.490 ;
        RECT 31.550 8.480 31.700 8.640 ;
        RECT 27.295 7.360 27.805 7.825 ;
        RECT 26.930 7.355 27.805 7.360 ;
        RECT 26.000 6.950 27.805 7.355 ;
        RECT 26.000 6.110 26.300 6.950 ;
        RECT 26.930 6.935 27.805 6.950 ;
        RECT 27.295 6.825 27.805 6.935 ;
        RECT 27.295 6.125 27.810 6.825 ;
        RECT 28.035 6.795 29.035 7.825 ;
        RECT 23.695 5.965 24.035 5.970 ;
        RECT 23.670 4.020 24.035 5.965 ;
        RECT 25.250 5.900 25.480 5.970 ;
        RECT 24.755 5.230 25.480 5.900 ;
        RECT 24.745 5.040 25.480 5.230 ;
        RECT 24.745 4.240 25.100 5.040 ;
        RECT 25.250 4.970 25.480 5.040 ;
        RECT 25.690 5.925 25.920 5.970 ;
        RECT 26.060 5.925 26.300 6.110 ;
        RECT 25.690 5.595 26.300 5.925 ;
        RECT 27.275 5.870 27.505 5.975 ;
        RECT 25.690 5.040 26.185 5.595 ;
        RECT 25.690 4.970 25.920 5.040 ;
        RECT 25.440 4.785 25.730 4.810 ;
        RECT 25.425 4.535 25.760 4.785 ;
        RECT 27.045 4.765 27.505 5.870 ;
        RECT 26.725 4.240 27.505 4.765 ;
        RECT 24.305 4.060 27.505 4.240 ;
        RECT 23.670 3.965 23.900 4.020 ;
        RECT 19.660 3.575 23.620 3.805 ;
        RECT 24.305 3.620 27.110 4.060 ;
        RECT 27.275 3.975 27.505 4.060 ;
        RECT 27.715 5.910 27.945 5.975 ;
        RECT 28.110 5.910 28.480 6.795 ;
        RECT 27.715 5.585 28.480 5.910 ;
        RECT 27.715 4.045 28.475 5.585 ;
        RECT 27.715 3.975 27.945 4.045 ;
        RECT 27.465 3.795 27.755 3.815 ;
        RECT 24.305 3.255 26.770 3.620 ;
        RECT 27.440 3.545 27.775 3.795 ;
        RECT 30.010 3.280 30.505 8.395 ;
        RECT 31.525 8.345 31.730 8.480 ;
        RECT 33.010 8.395 33.240 8.645 ;
        RECT 34.030 8.550 34.780 8.990 ;
        RECT 35.200 8.775 36.215 9.775 ;
        RECT 30.805 8.115 32.805 8.345 ;
        RECT 34.030 6.355 34.400 8.550 ;
        RECT 34.550 8.490 34.780 8.550 ;
        RECT 35.270 8.285 36.160 8.775 ;
        RECT 36.840 8.580 38.210 16.380 ;
        RECT 38.745 11.635 39.635 16.695 ;
        RECT 40.270 16.410 40.500 16.490 ;
        RECT 38.740 10.015 39.640 11.635 ;
        RECT 38.745 9.605 39.635 10.015 ;
        RECT 38.670 8.605 39.700 9.605 ;
        RECT 40.270 8.625 40.645 16.410 ;
        RECT 40.920 16.025 42.600 17.260 ;
        RECT 43.435 16.025 48.360 16.035 ;
        RECT 40.920 15.545 48.360 16.025 ;
        RECT 40.920 13.285 42.600 15.545 ;
        RECT 43.435 15.125 48.360 15.545 ;
        RECT 42.940 14.935 43.195 14.960 ;
        RECT 42.940 14.920 43.215 14.935 ;
        RECT 42.910 14.645 43.245 14.920 ;
        RECT 43.420 14.895 48.420 15.125 ;
        RECT 48.630 14.935 48.885 14.960 ;
        RECT 42.940 14.630 43.195 14.645 ;
        RECT 43.420 14.455 48.420 14.685 ;
        RECT 48.625 14.645 48.885 14.935 ;
        RECT 48.630 14.630 48.885 14.645 ;
        RECT 43.465 14.445 48.320 14.455 ;
        RECT 43.465 12.920 46.110 12.925 ;
        RECT 42.140 12.720 46.110 12.920 ;
        RECT 42.140 12.690 46.100 12.720 ;
        RECT 40.980 12.335 41.315 12.610 ;
        RECT 41.860 12.440 42.090 12.485 ;
        RECT 36.840 8.560 37.195 8.580 ;
        RECT 36.840 8.490 37.070 8.560 ;
        RECT 37.980 8.490 38.210 8.580 ;
        RECT 38.740 8.465 39.650 8.605 ;
        RECT 40.270 8.490 40.660 8.625 ;
        RECT 38.730 8.285 39.740 8.465 ;
        RECT 34.830 8.055 36.790 8.285 ;
        RECT 38.260 8.055 40.220 8.285 ;
        RECT 35.630 7.040 35.980 8.055 ;
        RECT 38.285 8.050 40.170 8.055 ;
        RECT 40.465 6.355 40.660 8.490 ;
        RECT 41.050 6.830 41.240 12.335 ;
        RECT 41.670 11.105 42.090 12.440 ;
        RECT 43.395 11.105 44.740 12.690 ;
        RECT 41.670 9.720 44.740 11.105 ;
        RECT 41.670 8.990 42.090 9.720 ;
        RECT 41.665 8.485 42.090 8.990 ;
        RECT 41.050 6.640 41.365 6.830 ;
        RECT 31.370 6.125 35.330 6.355 ;
        RECT 36.800 6.125 40.760 6.355 ;
        RECT 41.175 6.130 41.365 6.640 ;
        RECT 31.090 5.515 31.320 5.965 ;
        RECT 32.570 5.515 33.360 6.125 ;
        RECT 31.090 5.210 33.360 5.515 ;
        RECT 31.035 5.195 33.360 5.210 ;
        RECT 30.950 4.350 33.360 5.195 ;
        RECT 30.950 3.975 31.320 4.350 ;
        RECT 31.090 3.965 31.320 3.975 ;
        RECT 32.570 3.805 33.360 4.350 ;
        RECT 35.380 5.880 35.610 5.965 ;
        RECT 36.520 5.880 36.750 5.965 ;
        RECT 35.380 4.055 36.750 5.880 ;
        RECT 35.380 3.965 35.610 4.055 ;
        RECT 31.370 3.575 35.330 3.805 ;
        RECT 28.410 3.255 30.510 3.280 ;
        RECT 30.950 3.255 31.175 3.265 ;
        RECT 35.850 3.255 36.340 4.055 ;
        RECT 36.520 3.965 36.750 4.055 ;
        RECT 38.235 5.745 39.575 6.125 ;
        RECT 40.810 5.745 41.040 5.965 ;
        RECT 38.235 4.150 41.040 5.745 ;
        RECT 38.235 3.805 39.575 4.150 ;
        RECT 40.810 3.965 41.040 4.150 ;
        RECT 36.800 3.575 40.760 3.805 ;
        RECT 41.190 3.785 41.365 6.130 ;
        RECT 41.665 5.965 41.960 8.485 ;
        RECT 43.395 8.280 44.740 9.720 ;
        RECT 46.150 12.390 46.380 12.485 ;
        RECT 46.625 12.390 47.115 14.445 ;
        RECT 47.685 12.920 48.320 12.925 ;
        RECT 47.570 12.690 51.530 12.920 ;
        RECT 47.290 12.390 47.520 12.485 ;
        RECT 46.150 8.565 47.520 12.390 ;
        RECT 46.150 8.485 46.380 8.565 ;
        RECT 47.290 8.485 47.520 8.565 ;
        RECT 48.945 8.280 50.290 12.690 ;
        RECT 51.580 12.420 51.810 12.485 ;
        RECT 52.465 12.425 52.940 17.260 ;
        RECT 54.265 16.455 54.945 17.260 ;
        RECT 55.365 16.735 55.700 16.985 ;
        RECT 55.380 16.710 55.670 16.735 ;
        RECT 58.840 16.635 60.750 17.260 ;
        RECT 62.840 16.925 64.725 16.930 ;
        RECT 66.285 16.925 68.170 16.930 ;
        RECT 62.830 16.695 64.790 16.925 ;
        RECT 66.260 16.695 68.220 16.925 ;
        RECT 55.190 16.455 55.420 16.505 ;
        RECT 54.265 15.955 55.420 16.455 ;
        RECT 53.335 12.735 53.670 12.985 ;
        RECT 53.355 12.705 53.645 12.735 ;
        RECT 53.165 12.425 53.395 12.500 ;
        RECT 51.580 8.485 52.035 12.420 ;
        RECT 52.465 11.680 53.395 12.425 ;
        RECT 52.800 8.565 53.395 11.680 ;
        RECT 53.165 8.500 53.395 8.565 ;
        RECT 53.605 12.475 53.835 12.500 ;
        RECT 53.605 8.920 54.115 12.475 ;
        RECT 53.605 8.550 54.300 8.920 ;
        RECT 54.800 8.600 55.420 15.955 ;
        RECT 53.605 8.500 53.835 8.550 ;
        RECT 42.140 8.250 46.100 8.280 ;
        RECT 47.570 8.250 51.530 8.280 ;
        RECT 42.140 8.090 51.530 8.250 ;
        RECT 42.140 8.050 46.100 8.090 ;
        RECT 47.570 8.050 51.530 8.090 ;
        RECT 51.695 6.660 52.035 8.485 ;
        RECT 53.345 6.660 53.765 8.305 ;
        RECT 51.695 6.505 53.765 6.660 ;
        RECT 51.770 6.390 53.765 6.505 ;
        RECT 42.230 6.125 46.190 6.355 ;
        RECT 47.660 6.125 51.620 6.355 ;
        RECT 41.665 5.205 42.180 5.965 ;
        RECT 41.735 4.025 42.180 5.205 ;
        RECT 41.950 3.965 42.180 4.025 ;
        RECT 43.610 3.805 44.565 6.125 ;
        RECT 46.240 5.900 46.470 5.965 ;
        RECT 47.380 5.900 47.610 5.965 ;
        RECT 46.240 4.030 47.610 5.900 ;
        RECT 46.240 3.965 46.470 4.030 ;
        RECT 41.175 3.255 41.365 3.785 ;
        RECT 42.230 3.575 46.190 3.805 ;
        RECT 46.645 3.255 47.200 4.030 ;
        RECT 47.380 3.965 47.610 4.030 ;
        RECT 49.055 3.805 50.010 6.125 ;
        RECT 51.770 5.970 52.035 6.390 ;
        RECT 53.345 6.115 53.765 6.390 ;
        RECT 54.000 7.355 54.300 8.550 ;
        RECT 55.190 8.505 55.420 8.600 ;
        RECT 55.630 16.430 55.860 16.505 ;
        RECT 55.630 9.110 56.405 16.430 ;
        RECT 58.805 16.405 60.805 16.635 ;
        RECT 62.550 16.410 62.780 16.490 ;
        RECT 58.370 13.060 58.600 16.355 ;
        RECT 61.010 16.275 61.240 16.355 ;
        RECT 60.980 13.060 61.240 16.275 ;
        RECT 58.370 11.245 61.240 13.060 ;
        RECT 55.630 8.580 56.480 9.110 ;
        RECT 58.370 8.825 58.600 11.245 ;
        RECT 55.630 8.505 55.860 8.580 ;
        RECT 55.295 7.825 55.810 8.315 ;
        RECT 55.295 7.360 55.805 7.825 ;
        RECT 56.110 7.795 56.480 8.580 ;
        RECT 58.010 8.395 58.600 8.825 ;
        RECT 59.495 8.640 59.755 8.960 ;
        RECT 60.980 8.645 61.240 11.245 ;
        RECT 62.310 8.990 62.780 16.410 ;
        RECT 63.270 9.775 64.160 16.695 ;
        RECT 64.840 16.390 65.070 16.490 ;
        RECT 64.840 16.380 65.195 16.390 ;
        RECT 65.980 16.380 66.210 16.490 ;
        RECT 59.550 8.480 59.700 8.640 ;
        RECT 54.930 7.355 55.805 7.360 ;
        RECT 54.000 6.950 55.805 7.355 ;
        RECT 54.000 6.110 54.300 6.950 ;
        RECT 54.930 6.935 55.805 6.950 ;
        RECT 55.295 6.825 55.805 6.935 ;
        RECT 55.295 6.125 55.810 6.825 ;
        RECT 56.035 6.795 57.065 7.795 ;
        RECT 51.695 5.965 52.035 5.970 ;
        RECT 51.670 4.020 52.035 5.965 ;
        RECT 53.250 5.900 53.480 5.970 ;
        RECT 52.755 5.230 53.480 5.900 ;
        RECT 52.745 5.040 53.480 5.230 ;
        RECT 52.745 4.240 53.100 5.040 ;
        RECT 53.250 4.970 53.480 5.040 ;
        RECT 53.690 5.925 53.920 5.970 ;
        RECT 54.060 5.925 54.300 6.110 ;
        RECT 53.690 5.595 54.300 5.925 ;
        RECT 55.275 5.870 55.505 5.975 ;
        RECT 53.690 5.040 54.185 5.595 ;
        RECT 53.690 4.970 53.920 5.040 ;
        RECT 53.440 4.785 53.730 4.810 ;
        RECT 53.425 4.535 53.760 4.785 ;
        RECT 55.045 4.765 55.505 5.870 ;
        RECT 54.725 4.240 55.505 4.765 ;
        RECT 52.305 4.060 55.505 4.240 ;
        RECT 51.670 3.965 51.900 4.020 ;
        RECT 47.660 3.575 51.620 3.805 ;
        RECT 52.305 3.620 55.110 4.060 ;
        RECT 55.275 3.975 55.505 4.060 ;
        RECT 55.715 5.910 55.945 5.975 ;
        RECT 56.110 5.910 56.480 6.795 ;
        RECT 55.715 5.585 56.480 5.910 ;
        RECT 55.715 4.045 56.475 5.585 ;
        RECT 55.715 3.975 55.945 4.045 ;
        RECT 55.465 3.795 55.755 3.815 ;
        RECT 52.305 3.255 54.770 3.620 ;
        RECT 55.440 3.545 55.775 3.795 ;
        RECT 58.010 3.280 58.505 8.395 ;
        RECT 59.525 8.345 59.730 8.480 ;
        RECT 61.010 8.395 61.240 8.645 ;
        RECT 62.030 8.550 62.780 8.990 ;
        RECT 63.200 8.775 64.215 9.775 ;
        RECT 58.805 8.115 60.805 8.345 ;
        RECT 62.030 6.355 62.400 8.550 ;
        RECT 62.550 8.490 62.780 8.550 ;
        RECT 63.270 8.285 64.160 8.775 ;
        RECT 64.840 8.580 66.210 16.380 ;
        RECT 66.745 11.635 67.635 16.695 ;
        RECT 68.270 16.410 68.500 16.490 ;
        RECT 66.740 10.015 67.640 11.635 ;
        RECT 66.745 9.605 67.635 10.015 ;
        RECT 66.670 8.605 67.700 9.605 ;
        RECT 68.270 8.625 68.645 16.410 ;
        RECT 68.920 16.025 70.600 17.260 ;
        RECT 71.435 16.025 76.360 16.035 ;
        RECT 68.920 15.545 76.360 16.025 ;
        RECT 68.920 13.285 70.600 15.545 ;
        RECT 71.435 15.125 76.360 15.545 ;
        RECT 70.940 14.935 71.195 14.960 ;
        RECT 70.940 14.920 71.215 14.935 ;
        RECT 70.910 14.645 71.245 14.920 ;
        RECT 71.420 14.895 76.420 15.125 ;
        RECT 76.630 14.935 76.885 14.960 ;
        RECT 70.940 14.630 71.195 14.645 ;
        RECT 71.420 14.455 76.420 14.685 ;
        RECT 76.625 14.645 76.885 14.935 ;
        RECT 76.630 14.630 76.885 14.645 ;
        RECT 71.465 14.445 76.320 14.455 ;
        RECT 71.465 12.920 74.110 12.925 ;
        RECT 70.140 12.720 74.110 12.920 ;
        RECT 70.140 12.690 74.100 12.720 ;
        RECT 68.980 12.335 69.315 12.610 ;
        RECT 69.860 12.440 70.090 12.485 ;
        RECT 64.840 8.560 65.195 8.580 ;
        RECT 64.840 8.490 65.070 8.560 ;
        RECT 65.980 8.490 66.210 8.580 ;
        RECT 66.740 8.465 67.650 8.605 ;
        RECT 68.270 8.490 68.660 8.625 ;
        RECT 66.730 8.285 67.740 8.465 ;
        RECT 62.830 8.055 64.790 8.285 ;
        RECT 66.260 8.055 68.220 8.285 ;
        RECT 63.545 7.090 63.890 8.055 ;
        RECT 66.285 8.050 68.170 8.055 ;
        RECT 68.465 6.355 68.660 8.490 ;
        RECT 69.050 6.830 69.240 12.335 ;
        RECT 69.670 11.105 70.090 12.440 ;
        RECT 71.395 11.105 72.740 12.690 ;
        RECT 69.670 9.720 72.740 11.105 ;
        RECT 69.670 8.990 70.090 9.720 ;
        RECT 69.665 8.485 70.090 8.990 ;
        RECT 69.050 6.640 69.365 6.830 ;
        RECT 59.370 6.125 63.330 6.355 ;
        RECT 64.800 6.125 68.760 6.355 ;
        RECT 69.175 6.130 69.365 6.640 ;
        RECT 59.090 5.515 59.320 5.965 ;
        RECT 60.570 5.515 61.360 6.125 ;
        RECT 59.090 5.210 61.360 5.515 ;
        RECT 59.035 5.195 61.360 5.210 ;
        RECT 58.950 4.350 61.360 5.195 ;
        RECT 58.950 3.975 59.320 4.350 ;
        RECT 59.090 3.965 59.320 3.975 ;
        RECT 60.570 3.805 61.360 4.350 ;
        RECT 63.380 5.880 63.610 5.965 ;
        RECT 64.520 5.880 64.750 5.965 ;
        RECT 63.380 4.055 64.750 5.880 ;
        RECT 63.380 3.965 63.610 4.055 ;
        RECT 59.370 3.575 63.330 3.805 ;
        RECT 56.210 3.255 58.505 3.280 ;
        RECT 58.950 3.255 59.175 3.265 ;
        RECT 63.850 3.255 64.340 4.055 ;
        RECT 64.520 3.965 64.750 4.055 ;
        RECT 66.235 5.745 67.575 6.125 ;
        RECT 68.810 5.745 69.040 5.965 ;
        RECT 66.235 4.150 69.040 5.745 ;
        RECT 66.235 3.805 67.575 4.150 ;
        RECT 68.810 3.965 69.040 4.150 ;
        RECT 64.800 3.575 68.760 3.805 ;
        RECT 69.190 3.785 69.365 6.130 ;
        RECT 69.665 5.965 69.960 8.485 ;
        RECT 71.395 8.280 72.740 9.720 ;
        RECT 74.150 12.390 74.380 12.485 ;
        RECT 74.625 12.390 75.115 14.445 ;
        RECT 75.685 12.920 76.320 12.925 ;
        RECT 75.570 12.690 79.530 12.920 ;
        RECT 75.290 12.390 75.520 12.485 ;
        RECT 74.150 8.565 75.520 12.390 ;
        RECT 74.150 8.485 74.380 8.565 ;
        RECT 75.290 8.485 75.520 8.565 ;
        RECT 76.945 8.280 78.290 12.690 ;
        RECT 79.580 12.420 79.810 12.485 ;
        RECT 80.465 12.425 80.940 17.260 ;
        RECT 82.265 16.455 82.945 17.260 ;
        RECT 83.365 16.735 83.700 16.985 ;
        RECT 83.380 16.710 83.670 16.735 ;
        RECT 86.840 16.635 88.750 17.260 ;
        RECT 90.840 16.925 92.725 16.930 ;
        RECT 94.285 16.925 96.170 16.930 ;
        RECT 90.830 16.695 92.790 16.925 ;
        RECT 94.260 16.695 96.220 16.925 ;
        RECT 83.190 16.455 83.420 16.505 ;
        RECT 82.265 15.955 83.420 16.455 ;
        RECT 81.335 12.735 81.670 12.985 ;
        RECT 81.355 12.705 81.645 12.735 ;
        RECT 81.165 12.425 81.395 12.500 ;
        RECT 79.580 8.485 80.035 12.420 ;
        RECT 80.465 11.680 81.395 12.425 ;
        RECT 80.800 8.565 81.395 11.680 ;
        RECT 81.165 8.500 81.395 8.565 ;
        RECT 81.605 12.475 81.835 12.500 ;
        RECT 81.605 8.920 82.115 12.475 ;
        RECT 81.605 8.550 82.300 8.920 ;
        RECT 82.800 8.600 83.420 15.955 ;
        RECT 81.605 8.500 81.835 8.550 ;
        RECT 70.140 8.250 74.100 8.280 ;
        RECT 75.570 8.250 79.530 8.280 ;
        RECT 70.140 8.090 79.530 8.250 ;
        RECT 70.140 8.050 74.100 8.090 ;
        RECT 75.570 8.050 79.530 8.090 ;
        RECT 79.695 6.660 80.035 8.485 ;
        RECT 81.345 6.660 81.765 8.305 ;
        RECT 79.695 6.505 81.765 6.660 ;
        RECT 79.770 6.390 81.765 6.505 ;
        RECT 70.230 6.125 74.190 6.355 ;
        RECT 75.660 6.125 79.620 6.355 ;
        RECT 69.665 5.205 70.180 5.965 ;
        RECT 69.735 4.025 70.180 5.205 ;
        RECT 69.950 3.965 70.180 4.025 ;
        RECT 71.610 3.805 72.565 6.125 ;
        RECT 74.240 5.900 74.470 5.965 ;
        RECT 75.380 5.900 75.610 5.965 ;
        RECT 74.240 4.030 75.610 5.900 ;
        RECT 74.240 3.965 74.470 4.030 ;
        RECT 69.175 3.255 69.365 3.785 ;
        RECT 70.230 3.575 74.190 3.805 ;
        RECT 74.645 3.255 75.200 4.030 ;
        RECT 75.380 3.965 75.610 4.030 ;
        RECT 77.055 3.805 78.010 6.125 ;
        RECT 79.770 5.970 80.035 6.390 ;
        RECT 81.345 6.115 81.765 6.390 ;
        RECT 82.000 7.355 82.300 8.550 ;
        RECT 83.190 8.505 83.420 8.600 ;
        RECT 83.630 16.430 83.860 16.505 ;
        RECT 83.630 9.110 84.405 16.430 ;
        RECT 86.805 16.405 88.805 16.635 ;
        RECT 90.550 16.410 90.780 16.490 ;
        RECT 86.370 13.060 86.600 16.355 ;
        RECT 89.010 16.275 89.240 16.355 ;
        RECT 88.980 13.060 89.240 16.275 ;
        RECT 86.370 11.245 89.240 13.060 ;
        RECT 83.630 8.580 84.480 9.110 ;
        RECT 86.370 8.825 86.600 11.245 ;
        RECT 83.630 8.505 83.860 8.580 ;
        RECT 83.295 7.825 83.810 8.315 ;
        RECT 83.295 7.360 83.805 7.825 ;
        RECT 84.110 7.795 84.480 8.580 ;
        RECT 86.010 8.395 86.600 8.825 ;
        RECT 87.495 8.640 87.755 8.960 ;
        RECT 88.980 8.645 89.240 11.245 ;
        RECT 90.310 8.990 90.780 16.410 ;
        RECT 91.270 9.775 92.160 16.695 ;
        RECT 92.840 16.390 93.070 16.490 ;
        RECT 92.840 16.380 93.195 16.390 ;
        RECT 93.980 16.380 94.210 16.490 ;
        RECT 87.550 8.480 87.700 8.640 ;
        RECT 82.930 7.355 83.805 7.360 ;
        RECT 82.000 6.950 83.805 7.355 ;
        RECT 82.000 6.110 82.300 6.950 ;
        RECT 82.930 6.935 83.805 6.950 ;
        RECT 83.295 6.825 83.805 6.935 ;
        RECT 83.295 6.125 83.810 6.825 ;
        RECT 84.035 6.795 85.065 7.795 ;
        RECT 79.695 5.965 80.035 5.970 ;
        RECT 79.670 4.020 80.035 5.965 ;
        RECT 81.250 5.900 81.480 5.970 ;
        RECT 80.755 5.230 81.480 5.900 ;
        RECT 80.745 5.040 81.480 5.230 ;
        RECT 80.745 4.240 81.100 5.040 ;
        RECT 81.250 4.970 81.480 5.040 ;
        RECT 81.690 5.925 81.920 5.970 ;
        RECT 82.060 5.925 82.300 6.110 ;
        RECT 81.690 5.595 82.300 5.925 ;
        RECT 83.275 5.870 83.505 5.975 ;
        RECT 81.690 5.040 82.185 5.595 ;
        RECT 81.690 4.970 81.920 5.040 ;
        RECT 81.440 4.785 81.730 4.810 ;
        RECT 81.425 4.535 81.760 4.785 ;
        RECT 83.045 4.765 83.505 5.870 ;
        RECT 82.725 4.240 83.505 4.765 ;
        RECT 80.305 4.060 83.505 4.240 ;
        RECT 79.670 3.965 79.900 4.020 ;
        RECT 75.660 3.575 79.620 3.805 ;
        RECT 80.305 3.620 83.110 4.060 ;
        RECT 83.275 3.975 83.505 4.060 ;
        RECT 83.715 5.910 83.945 5.975 ;
        RECT 84.110 5.910 84.480 6.795 ;
        RECT 83.715 5.585 84.480 5.910 ;
        RECT 83.715 4.045 84.475 5.585 ;
        RECT 83.715 3.975 83.945 4.045 ;
        RECT 83.465 3.795 83.755 3.815 ;
        RECT 80.305 3.255 82.770 3.620 ;
        RECT 83.440 3.545 83.775 3.795 ;
        RECT 86.010 3.280 86.505 8.395 ;
        RECT 87.525 8.345 87.730 8.480 ;
        RECT 89.010 8.395 89.240 8.645 ;
        RECT 90.030 8.550 90.780 8.990 ;
        RECT 91.200 8.775 92.215 9.775 ;
        RECT 86.805 8.115 88.805 8.345 ;
        RECT 90.030 6.355 90.400 8.550 ;
        RECT 90.550 8.490 90.780 8.550 ;
        RECT 91.270 8.285 92.160 8.775 ;
        RECT 92.840 8.580 94.210 16.380 ;
        RECT 94.745 11.635 95.635 16.695 ;
        RECT 96.270 16.410 96.500 16.490 ;
        RECT 94.740 10.015 95.640 11.635 ;
        RECT 94.745 9.605 95.635 10.015 ;
        RECT 94.670 8.605 95.700 9.605 ;
        RECT 96.270 8.625 96.645 16.410 ;
        RECT 96.920 16.025 98.600 17.260 ;
        RECT 99.435 16.025 104.360 16.035 ;
        RECT 96.920 15.545 104.360 16.025 ;
        RECT 96.920 13.285 98.600 15.545 ;
        RECT 99.435 15.125 104.360 15.545 ;
        RECT 98.940 14.935 99.195 14.960 ;
        RECT 98.940 14.920 99.215 14.935 ;
        RECT 98.910 14.645 99.245 14.920 ;
        RECT 99.420 14.895 104.420 15.125 ;
        RECT 104.630 14.935 104.885 14.960 ;
        RECT 98.940 14.630 99.195 14.645 ;
        RECT 99.420 14.455 104.420 14.685 ;
        RECT 104.625 14.645 104.885 14.935 ;
        RECT 104.630 14.630 104.885 14.645 ;
        RECT 99.465 14.445 104.320 14.455 ;
        RECT 99.465 12.920 102.110 12.925 ;
        RECT 98.140 12.720 102.110 12.920 ;
        RECT 98.140 12.690 102.100 12.720 ;
        RECT 96.980 12.335 97.315 12.610 ;
        RECT 97.860 12.440 98.090 12.485 ;
        RECT 92.840 8.560 93.195 8.580 ;
        RECT 92.840 8.490 93.070 8.560 ;
        RECT 93.980 8.490 94.210 8.580 ;
        RECT 94.740 8.465 95.650 8.605 ;
        RECT 96.270 8.490 96.660 8.625 ;
        RECT 94.730 8.285 95.740 8.465 ;
        RECT 90.830 8.055 92.790 8.285 ;
        RECT 94.260 8.055 96.220 8.285 ;
        RECT 91.515 6.975 91.915 8.055 ;
        RECT 94.285 8.050 96.170 8.055 ;
        RECT 96.465 6.355 96.660 8.490 ;
        RECT 97.050 6.830 97.240 12.335 ;
        RECT 97.670 11.105 98.090 12.440 ;
        RECT 99.395 11.105 100.740 12.690 ;
        RECT 97.670 9.720 100.740 11.105 ;
        RECT 97.670 8.990 98.090 9.720 ;
        RECT 97.665 8.485 98.090 8.990 ;
        RECT 97.050 6.640 97.365 6.830 ;
        RECT 87.370 6.125 91.330 6.355 ;
        RECT 92.800 6.125 96.760 6.355 ;
        RECT 97.175 6.130 97.365 6.640 ;
        RECT 87.090 5.515 87.320 5.965 ;
        RECT 88.570 5.515 89.360 6.125 ;
        RECT 87.090 5.210 89.360 5.515 ;
        RECT 87.035 5.195 89.360 5.210 ;
        RECT 86.950 4.350 89.360 5.195 ;
        RECT 86.950 3.975 87.320 4.350 ;
        RECT 87.090 3.965 87.320 3.975 ;
        RECT 88.570 3.805 89.360 4.350 ;
        RECT 91.380 5.880 91.610 5.965 ;
        RECT 92.520 5.880 92.750 5.965 ;
        RECT 91.380 4.055 92.750 5.880 ;
        RECT 91.380 3.965 91.610 4.055 ;
        RECT 87.370 3.575 91.330 3.805 ;
        RECT 84.310 3.255 86.505 3.280 ;
        RECT 86.950 3.255 87.175 3.265 ;
        RECT 91.850 3.255 92.340 4.055 ;
        RECT 92.520 3.965 92.750 4.055 ;
        RECT 94.235 5.745 95.575 6.125 ;
        RECT 96.810 5.745 97.040 5.965 ;
        RECT 94.235 4.150 97.040 5.745 ;
        RECT 94.235 3.805 95.575 4.150 ;
        RECT 96.810 3.965 97.040 4.150 ;
        RECT 92.800 3.575 96.760 3.805 ;
        RECT 97.190 3.785 97.365 6.130 ;
        RECT 97.665 5.965 97.960 8.485 ;
        RECT 99.395 8.280 100.740 9.720 ;
        RECT 102.150 12.390 102.380 12.485 ;
        RECT 102.625 12.390 103.115 14.445 ;
        RECT 103.685 12.920 104.320 12.925 ;
        RECT 103.570 12.690 107.530 12.920 ;
        RECT 103.290 12.390 103.520 12.485 ;
        RECT 102.150 8.565 103.520 12.390 ;
        RECT 102.150 8.485 102.380 8.565 ;
        RECT 103.290 8.485 103.520 8.565 ;
        RECT 104.945 8.280 106.290 12.690 ;
        RECT 107.580 12.420 107.810 12.485 ;
        RECT 108.465 12.425 108.940 17.260 ;
        RECT 110.265 16.455 110.945 17.260 ;
        RECT 111.365 16.735 111.700 16.985 ;
        RECT 111.380 16.710 111.670 16.735 ;
        RECT 114.840 16.635 116.750 17.260 ;
        RECT 118.840 16.925 120.725 16.930 ;
        RECT 122.285 16.925 124.170 16.930 ;
        RECT 118.830 16.695 120.790 16.925 ;
        RECT 122.260 16.695 124.220 16.925 ;
        RECT 111.190 16.455 111.420 16.505 ;
        RECT 110.265 15.955 111.420 16.455 ;
        RECT 109.335 12.735 109.670 12.985 ;
        RECT 109.355 12.705 109.645 12.735 ;
        RECT 109.165 12.425 109.395 12.500 ;
        RECT 107.580 8.485 108.035 12.420 ;
        RECT 108.465 11.680 109.395 12.425 ;
        RECT 108.800 8.565 109.395 11.680 ;
        RECT 109.165 8.500 109.395 8.565 ;
        RECT 109.605 12.475 109.835 12.500 ;
        RECT 109.605 8.920 110.115 12.475 ;
        RECT 109.605 8.550 110.300 8.920 ;
        RECT 110.800 8.600 111.420 15.955 ;
        RECT 109.605 8.500 109.835 8.550 ;
        RECT 98.140 8.250 102.100 8.280 ;
        RECT 103.570 8.250 107.530 8.280 ;
        RECT 98.140 8.090 107.530 8.250 ;
        RECT 98.140 8.050 102.100 8.090 ;
        RECT 103.570 8.050 107.530 8.090 ;
        RECT 107.695 6.660 108.035 8.485 ;
        RECT 109.345 6.660 109.765 8.305 ;
        RECT 107.695 6.505 109.765 6.660 ;
        RECT 107.770 6.390 109.765 6.505 ;
        RECT 98.230 6.125 102.190 6.355 ;
        RECT 103.660 6.125 107.620 6.355 ;
        RECT 97.665 5.205 98.180 5.965 ;
        RECT 97.735 4.025 98.180 5.205 ;
        RECT 97.950 3.965 98.180 4.025 ;
        RECT 99.610 3.805 100.565 6.125 ;
        RECT 102.240 5.900 102.470 5.965 ;
        RECT 103.380 5.900 103.610 5.965 ;
        RECT 102.240 4.030 103.610 5.900 ;
        RECT 102.240 3.965 102.470 4.030 ;
        RECT 97.175 3.255 97.365 3.785 ;
        RECT 98.230 3.575 102.190 3.805 ;
        RECT 102.645 3.255 103.200 4.030 ;
        RECT 103.380 3.965 103.610 4.030 ;
        RECT 105.055 3.805 106.010 6.125 ;
        RECT 107.770 5.970 108.035 6.390 ;
        RECT 109.345 6.115 109.765 6.390 ;
        RECT 110.000 7.355 110.300 8.550 ;
        RECT 111.190 8.505 111.420 8.600 ;
        RECT 111.630 16.430 111.860 16.505 ;
        RECT 111.630 9.110 112.405 16.430 ;
        RECT 114.805 16.405 116.805 16.635 ;
        RECT 118.550 16.410 118.780 16.490 ;
        RECT 114.370 13.060 114.600 16.355 ;
        RECT 117.010 16.275 117.240 16.355 ;
        RECT 116.980 13.060 117.240 16.275 ;
        RECT 114.370 11.245 117.240 13.060 ;
        RECT 111.630 8.580 112.480 9.110 ;
        RECT 114.370 8.825 114.600 11.245 ;
        RECT 111.630 8.505 111.860 8.580 ;
        RECT 111.295 7.825 111.810 8.315 ;
        RECT 111.295 7.360 111.805 7.825 ;
        RECT 112.110 7.795 112.480 8.580 ;
        RECT 114.010 8.395 114.600 8.825 ;
        RECT 115.495 8.640 115.755 8.960 ;
        RECT 116.980 8.645 117.240 11.245 ;
        RECT 118.310 8.990 118.780 16.410 ;
        RECT 119.270 9.775 120.160 16.695 ;
        RECT 120.840 16.390 121.070 16.490 ;
        RECT 120.840 16.380 121.195 16.390 ;
        RECT 121.980 16.380 122.210 16.490 ;
        RECT 115.550 8.480 115.700 8.640 ;
        RECT 110.930 7.355 111.805 7.360 ;
        RECT 110.000 6.950 111.805 7.355 ;
        RECT 110.000 6.110 110.300 6.950 ;
        RECT 110.930 6.935 111.805 6.950 ;
        RECT 111.295 6.825 111.805 6.935 ;
        RECT 111.295 6.125 111.810 6.825 ;
        RECT 112.035 6.795 113.065 7.795 ;
        RECT 107.695 5.965 108.035 5.970 ;
        RECT 107.670 4.020 108.035 5.965 ;
        RECT 109.250 5.900 109.480 5.970 ;
        RECT 108.755 5.230 109.480 5.900 ;
        RECT 108.745 5.040 109.480 5.230 ;
        RECT 108.745 4.240 109.100 5.040 ;
        RECT 109.250 4.970 109.480 5.040 ;
        RECT 109.690 5.925 109.920 5.970 ;
        RECT 110.060 5.925 110.300 6.110 ;
        RECT 109.690 5.595 110.300 5.925 ;
        RECT 111.275 5.870 111.505 5.975 ;
        RECT 109.690 5.040 110.185 5.595 ;
        RECT 109.690 4.970 109.920 5.040 ;
        RECT 109.440 4.785 109.730 4.810 ;
        RECT 109.425 4.535 109.760 4.785 ;
        RECT 111.045 4.765 111.505 5.870 ;
        RECT 110.725 4.240 111.505 4.765 ;
        RECT 108.305 4.060 111.505 4.240 ;
        RECT 107.670 3.965 107.900 4.020 ;
        RECT 103.660 3.575 107.620 3.805 ;
        RECT 108.305 3.620 111.110 4.060 ;
        RECT 111.275 3.975 111.505 4.060 ;
        RECT 111.715 5.910 111.945 5.975 ;
        RECT 112.110 5.910 112.480 6.795 ;
        RECT 111.715 5.585 112.480 5.910 ;
        RECT 111.715 4.045 112.475 5.585 ;
        RECT 111.715 3.975 111.945 4.045 ;
        RECT 111.465 3.795 111.755 3.815 ;
        RECT 108.305 3.255 110.770 3.620 ;
        RECT 111.440 3.545 111.775 3.795 ;
        RECT 114.010 3.280 114.505 8.395 ;
        RECT 115.525 8.345 115.730 8.480 ;
        RECT 117.010 8.395 117.240 8.645 ;
        RECT 118.030 8.550 118.780 8.990 ;
        RECT 119.200 8.775 120.215 9.775 ;
        RECT 114.805 8.115 116.805 8.345 ;
        RECT 118.030 6.355 118.400 8.550 ;
        RECT 118.550 8.490 118.780 8.550 ;
        RECT 119.270 8.285 120.160 8.775 ;
        RECT 120.840 8.580 122.210 16.380 ;
        RECT 122.745 11.635 123.635 16.695 ;
        RECT 124.270 16.410 124.500 16.490 ;
        RECT 122.740 10.015 123.640 11.635 ;
        RECT 122.745 9.605 123.635 10.015 ;
        RECT 122.670 8.605 123.700 9.605 ;
        RECT 124.270 8.625 124.645 16.410 ;
        RECT 124.920 16.025 126.600 17.260 ;
        RECT 127.435 16.025 132.360 16.035 ;
        RECT 124.920 15.545 132.360 16.025 ;
        RECT 124.920 13.285 126.600 15.545 ;
        RECT 127.435 15.125 132.360 15.545 ;
        RECT 126.940 14.935 127.195 14.960 ;
        RECT 126.940 14.920 127.215 14.935 ;
        RECT 126.910 14.645 127.245 14.920 ;
        RECT 127.420 14.895 132.420 15.125 ;
        RECT 132.630 14.935 132.885 14.960 ;
        RECT 126.940 14.630 127.195 14.645 ;
        RECT 127.420 14.455 132.420 14.685 ;
        RECT 132.625 14.645 132.885 14.935 ;
        RECT 132.630 14.630 132.885 14.645 ;
        RECT 127.465 14.445 132.320 14.455 ;
        RECT 127.465 12.920 130.110 12.925 ;
        RECT 126.140 12.720 130.110 12.920 ;
        RECT 126.140 12.690 130.100 12.720 ;
        RECT 124.980 12.335 125.315 12.610 ;
        RECT 125.860 12.440 126.090 12.485 ;
        RECT 120.840 8.560 121.195 8.580 ;
        RECT 120.840 8.490 121.070 8.560 ;
        RECT 121.980 8.490 122.210 8.580 ;
        RECT 122.740 8.465 123.650 8.605 ;
        RECT 124.270 8.490 124.660 8.625 ;
        RECT 122.730 8.285 123.740 8.465 ;
        RECT 118.830 8.055 120.790 8.285 ;
        RECT 122.260 8.055 124.220 8.285 ;
        RECT 119.570 7.155 119.855 8.055 ;
        RECT 122.285 8.050 124.170 8.055 ;
        RECT 124.465 6.355 124.660 8.490 ;
        RECT 125.050 6.830 125.240 12.335 ;
        RECT 125.670 11.105 126.090 12.440 ;
        RECT 127.395 11.105 128.740 12.690 ;
        RECT 125.670 9.720 128.740 11.105 ;
        RECT 125.670 8.990 126.090 9.720 ;
        RECT 125.665 8.485 126.090 8.990 ;
        RECT 125.050 6.640 125.365 6.830 ;
        RECT 115.370 6.125 119.330 6.355 ;
        RECT 120.800 6.125 124.760 6.355 ;
        RECT 125.175 6.130 125.365 6.640 ;
        RECT 115.090 5.515 115.320 5.965 ;
        RECT 116.570 5.515 117.360 6.125 ;
        RECT 115.090 5.210 117.360 5.515 ;
        RECT 115.035 5.195 117.360 5.210 ;
        RECT 114.950 4.350 117.360 5.195 ;
        RECT 114.950 3.975 115.320 4.350 ;
        RECT 115.090 3.965 115.320 3.975 ;
        RECT 116.570 3.805 117.360 4.350 ;
        RECT 119.380 5.880 119.610 5.965 ;
        RECT 120.520 5.880 120.750 5.965 ;
        RECT 119.380 4.055 120.750 5.880 ;
        RECT 119.380 3.965 119.610 4.055 ;
        RECT 115.370 3.575 119.330 3.805 ;
        RECT 112.010 3.255 114.505 3.280 ;
        RECT 114.950 3.255 115.175 3.265 ;
        RECT 119.850 3.255 120.340 4.055 ;
        RECT 120.520 3.965 120.750 4.055 ;
        RECT 122.235 5.745 123.575 6.125 ;
        RECT 124.810 5.745 125.040 5.965 ;
        RECT 122.235 4.150 125.040 5.745 ;
        RECT 122.235 3.805 123.575 4.150 ;
        RECT 124.810 3.965 125.040 4.150 ;
        RECT 120.800 3.575 124.760 3.805 ;
        RECT 125.190 3.785 125.365 6.130 ;
        RECT 125.665 5.965 125.960 8.485 ;
        RECT 127.395 8.280 128.740 9.720 ;
        RECT 130.150 12.390 130.380 12.485 ;
        RECT 130.625 12.390 131.115 14.445 ;
        RECT 131.685 12.920 132.320 12.925 ;
        RECT 131.570 12.690 135.530 12.920 ;
        RECT 131.290 12.390 131.520 12.485 ;
        RECT 130.150 8.565 131.520 12.390 ;
        RECT 130.150 8.485 130.380 8.565 ;
        RECT 131.290 8.485 131.520 8.565 ;
        RECT 132.945 8.280 134.290 12.690 ;
        RECT 135.580 12.420 135.810 12.485 ;
        RECT 136.465 12.425 136.940 17.260 ;
        RECT 138.265 16.455 138.945 17.260 ;
        RECT 139.365 16.735 139.700 16.985 ;
        RECT 139.380 16.710 139.670 16.735 ;
        RECT 139.190 16.455 139.420 16.505 ;
        RECT 138.265 15.955 139.420 16.455 ;
        RECT 137.335 12.735 137.670 12.985 ;
        RECT 137.355 12.705 137.645 12.735 ;
        RECT 137.165 12.425 137.395 12.500 ;
        RECT 135.580 8.485 136.035 12.420 ;
        RECT 136.465 11.680 137.395 12.425 ;
        RECT 136.800 8.565 137.395 11.680 ;
        RECT 137.165 8.500 137.395 8.565 ;
        RECT 137.605 12.475 137.835 12.500 ;
        RECT 137.605 8.920 138.115 12.475 ;
        RECT 137.605 8.550 138.300 8.920 ;
        RECT 138.800 8.600 139.420 15.955 ;
        RECT 137.605 8.500 137.835 8.550 ;
        RECT 126.140 8.250 130.100 8.280 ;
        RECT 131.570 8.250 135.530 8.280 ;
        RECT 126.140 8.090 135.530 8.250 ;
        RECT 126.140 8.050 130.100 8.090 ;
        RECT 131.570 8.050 135.530 8.090 ;
        RECT 135.695 6.660 136.035 8.485 ;
        RECT 137.345 6.660 137.765 8.305 ;
        RECT 135.695 6.505 137.765 6.660 ;
        RECT 135.770 6.390 137.765 6.505 ;
        RECT 126.230 6.125 130.190 6.355 ;
        RECT 131.660 6.125 135.620 6.355 ;
        RECT 125.665 5.205 126.180 5.965 ;
        RECT 125.735 4.025 126.180 5.205 ;
        RECT 125.950 3.965 126.180 4.025 ;
        RECT 127.610 3.805 128.565 6.125 ;
        RECT 130.240 5.900 130.470 5.965 ;
        RECT 131.380 5.900 131.610 5.965 ;
        RECT 130.240 4.030 131.610 5.900 ;
        RECT 130.240 3.965 130.470 4.030 ;
        RECT 125.175 3.255 125.365 3.785 ;
        RECT 126.230 3.575 130.190 3.805 ;
        RECT 130.645 3.255 131.200 4.030 ;
        RECT 131.380 3.965 131.610 4.030 ;
        RECT 133.055 3.805 134.010 6.125 ;
        RECT 135.770 5.970 136.035 6.390 ;
        RECT 137.345 6.115 137.765 6.390 ;
        RECT 138.000 7.355 138.300 8.550 ;
        RECT 139.190 8.505 139.420 8.600 ;
        RECT 139.630 16.430 139.860 16.505 ;
        RECT 139.630 9.110 140.405 16.430 ;
        RECT 139.630 8.580 140.480 9.110 ;
        RECT 139.630 8.505 139.860 8.580 ;
        RECT 139.295 7.825 139.810 8.315 ;
        RECT 139.295 7.360 139.805 7.825 ;
        RECT 140.110 7.795 140.480 8.580 ;
        RECT 138.930 7.355 139.805 7.360 ;
        RECT 138.000 6.950 139.805 7.355 ;
        RECT 138.000 6.110 138.300 6.950 ;
        RECT 138.930 6.935 139.805 6.950 ;
        RECT 139.295 6.825 139.805 6.935 ;
        RECT 139.295 6.125 139.810 6.825 ;
        RECT 140.035 6.795 141.065 7.795 ;
        RECT 135.695 5.965 136.035 5.970 ;
        RECT 135.670 4.020 136.035 5.965 ;
        RECT 137.250 5.900 137.480 5.970 ;
        RECT 136.755 5.230 137.480 5.900 ;
        RECT 136.745 5.040 137.480 5.230 ;
        RECT 136.745 4.240 137.100 5.040 ;
        RECT 137.250 4.970 137.480 5.040 ;
        RECT 137.690 5.925 137.920 5.970 ;
        RECT 138.060 5.925 138.300 6.110 ;
        RECT 137.690 5.595 138.300 5.925 ;
        RECT 139.275 5.870 139.505 5.975 ;
        RECT 137.690 5.040 138.185 5.595 ;
        RECT 137.690 4.970 137.920 5.040 ;
        RECT 137.440 4.785 137.730 4.810 ;
        RECT 137.425 4.535 137.760 4.785 ;
        RECT 139.045 4.765 139.505 5.870 ;
        RECT 138.725 4.240 139.505 4.765 ;
        RECT 136.305 4.060 139.505 4.240 ;
        RECT 135.670 3.965 135.900 4.020 ;
        RECT 131.660 3.575 135.620 3.805 ;
        RECT 136.305 3.620 139.110 4.060 ;
        RECT 139.275 3.975 139.505 4.060 ;
        RECT 139.715 5.910 139.945 5.975 ;
        RECT 140.110 5.910 140.480 6.795 ;
        RECT 139.715 5.585 140.480 5.910 ;
        RECT 139.715 4.045 140.475 5.585 ;
        RECT 139.715 3.975 139.945 4.045 ;
        RECT 139.465 3.795 139.755 3.815 ;
        RECT 136.305 3.255 138.770 3.620 ;
        RECT 139.440 3.545 139.775 3.795 ;
        RECT 1.895 2.380 140.500 3.255 ;
      LAYER met2 ;
        RECT 72.390 93.020 78.385 93.655 ;
        RECT 72.390 77.085 73.025 93.020 ;
        RECT 73.775 88.750 74.180 92.565 ;
        RECT 76.180 91.825 76.585 91.855 ;
        RECT 78.860 91.825 79.265 98.800 ;
        RECT 76.180 91.420 79.265 91.825 ;
        RECT 76.180 91.390 76.585 91.420 ;
        RECT 81.175 91.015 82.060 100.300 ;
        RECT 87.390 97.730 92.205 98.995 ;
        RECT 87.390 97.340 92.280 97.730 ;
        RECT 75.700 90.200 82.090 91.015 ;
        RECT 83.490 90.950 83.870 95.595 ;
        RECT 88.375 95.345 92.280 97.340 ;
        RECT 91.965 95.340 92.280 95.345 ;
        RECT 87.400 92.690 87.870 92.720 ;
        RECT 87.400 92.220 100.225 92.690 ;
        RECT 87.400 92.190 87.870 92.220 ;
        RECT 75.670 90.130 82.090 90.200 ;
        RECT 83.095 90.570 83.870 90.950 ;
        RECT 75.670 89.315 76.615 90.130 ;
        RECT 75.285 88.750 75.690 88.780 ;
        RECT 73.775 88.345 75.690 88.750 ;
        RECT 75.285 88.315 75.690 88.345 ;
        RECT 83.095 84.040 83.475 90.570 ;
        RECT 96.340 88.455 96.800 88.485 ;
        RECT 93.535 87.995 96.800 88.455 ;
        RECT 99.755 88.260 100.225 92.220 ;
        RECT 96.340 87.965 96.800 87.995 ;
        RECT 87.425 86.140 88.035 86.210 ;
        RECT 84.070 85.665 88.035 86.140 ;
        RECT 87.425 85.605 88.035 85.665 ;
        RECT 89.360 80.535 94.395 81.595 ;
        RECT 75.715 80.135 94.395 80.535 ;
        RECT 89.360 79.185 94.395 80.135 ;
        RECT 94.580 78.790 94.975 78.890 ;
        RECT 99.190 78.875 99.450 79.115 ;
        RECT 99.045 78.795 99.450 78.875 ;
        RECT 99.045 78.790 99.445 78.795 ;
        RECT 94.580 78.540 99.445 78.790 ;
        RECT 94.580 78.435 94.975 78.540 ;
        RECT 87.095 63.720 98.640 64.310 ;
        RECT 145.520 64.195 146.065 66.195 ;
        RECT 103.685 64.145 104.335 64.165 ;
        RECT 103.685 63.600 115.625 64.145 ;
        RECT 103.685 63.530 104.335 63.600 ;
        RECT 120.545 63.595 132.195 64.140 ;
        RECT 137.115 63.650 146.065 64.195 ;
        RECT 89.765 62.965 90.360 63.405 ;
        RECT 82.445 62.370 90.360 62.965 ;
        RECT 95.425 62.665 106.995 63.255 ;
        RECT 112.165 62.455 123.775 63.045 ;
        RECT 128.810 62.450 140.490 62.995 ;
        RECT 2.010 48.345 2.505 50.885 ;
        RECT 10.970 48.800 11.415 50.625 ;
        RECT 10.715 48.355 11.665 48.800 ;
        RECT 13.540 48.430 14.320 57.440 ;
        RECT 1.980 47.850 2.535 48.345 ;
        RECT 14.940 46.920 15.215 46.950 ;
        RECT 13.010 46.645 15.215 46.920 ;
        RECT 13.010 44.305 13.285 46.645 ;
        RECT 14.940 46.615 15.215 46.645 ;
        RECT 3.465 40.875 3.785 40.930 ;
        RECT 9.345 40.875 9.665 40.930 ;
        RECT 3.465 40.725 9.665 40.875 ;
        RECT 3.465 40.670 3.785 40.725 ;
        RECT 9.345 40.670 9.665 40.725 ;
        RECT 2.310 39.095 7.915 39.425 ;
        RECT 2.310 23.395 2.640 39.095 ;
        RECT 4.260 37.265 4.580 37.290 ;
        RECT 21.380 37.265 21.700 37.290 ;
        RECT 4.260 37.055 21.700 37.265 ;
        RECT 4.260 37.030 4.580 37.055 ;
        RECT 21.380 37.030 21.700 37.055 ;
        RECT 11.715 36.260 16.220 36.555 ;
        RECT 26.165 32.720 26.540 51.710 ;
        RECT 10.715 32.345 26.540 32.720 ;
        RECT 14.940 30.920 15.215 30.950 ;
        RECT 13.010 30.645 15.215 30.920 ;
        RECT 13.010 28.305 13.285 30.645 ;
        RECT 14.940 30.615 15.215 30.645 ;
        RECT 3.465 24.875 3.785 24.930 ;
        RECT 9.345 24.875 9.665 24.930 ;
        RECT 3.465 24.725 9.665 24.875 ;
        RECT 3.465 24.670 3.785 24.725 ;
        RECT 9.345 24.670 9.665 24.725 ;
        RECT 2.310 23.065 7.945 23.395 ;
        RECT 2.320 7.445 2.650 23.065 ;
        RECT 4.260 21.265 4.580 21.290 ;
        RECT 21.380 21.265 21.700 21.290 ;
        RECT 4.260 21.055 21.700 21.265 ;
        RECT 4.260 21.030 4.580 21.055 ;
        RECT 21.380 21.030 21.700 21.055 ;
        RECT 11.715 20.260 16.220 20.555 ;
        RECT 27.015 16.035 27.420 50.605 ;
        RECT 28.410 39.880 28.660 53.505 ;
        RECT 28.410 39.795 28.910 39.880 ;
        RECT 28.005 39.535 28.910 39.795 ;
        RECT 28.610 39.480 28.910 39.535 ;
        RECT 29.135 39.050 29.480 53.450 ;
        RECT 28.365 38.705 29.480 39.050 ;
        RECT 28.365 23.795 28.710 38.705 ;
        RECT 30.070 38.120 30.350 53.420 ;
        RECT 39.005 48.715 39.380 50.660 ;
        RECT 38.715 48.340 39.665 48.715 ;
        RECT 42.940 46.920 43.215 46.950 ;
        RECT 41.010 46.645 43.215 46.920 ;
        RECT 41.010 44.305 41.285 46.645 ;
        RECT 42.940 46.615 43.215 46.645 ;
        RECT 31.465 40.875 31.785 40.930 ;
        RECT 37.345 40.875 37.665 40.930 ;
        RECT 31.465 40.725 37.665 40.875 ;
        RECT 31.465 40.670 31.785 40.725 ;
        RECT 37.345 40.670 37.665 40.725 ;
        RECT 29.270 37.840 30.350 38.120 ;
        RECT 30.810 39.370 35.920 39.720 ;
        RECT 28.005 23.450 29.065 23.795 ;
        RECT 29.270 23.220 29.550 37.840 ;
        RECT 10.715 15.630 27.420 16.035 ;
        RECT 28.395 22.940 29.550 23.220 ;
        RECT 30.810 23.385 31.160 39.370 ;
        RECT 32.260 37.265 32.580 37.290 ;
        RECT 49.380 37.265 49.700 37.290 ;
        RECT 32.260 37.055 49.700 37.265 ;
        RECT 32.260 37.030 32.580 37.055 ;
        RECT 49.380 37.030 49.700 37.055 ;
        RECT 39.715 36.260 44.220 36.555 ;
        RECT 54.230 32.600 54.630 51.745 ;
        RECT 38.715 32.200 54.630 32.600 ;
        RECT 42.940 30.920 43.215 30.950 ;
        RECT 41.010 30.645 43.215 30.920 ;
        RECT 41.010 28.305 41.285 30.645 ;
        RECT 42.940 30.615 43.215 30.645 ;
        RECT 31.465 24.875 31.785 24.930 ;
        RECT 37.345 24.875 37.665 24.930 ;
        RECT 31.465 24.725 37.665 24.875 ;
        RECT 31.465 24.670 31.785 24.725 ;
        RECT 37.345 24.670 37.665 24.725 ;
        RECT 30.810 23.035 35.915 23.385 ;
        RECT 14.940 14.920 15.215 14.950 ;
        RECT 13.010 14.645 15.215 14.920 ;
        RECT 13.010 12.305 13.285 14.645 ;
        RECT 14.940 14.615 15.215 14.645 ;
        RECT 3.465 8.875 3.785 8.930 ;
        RECT 9.345 8.875 9.665 8.930 ;
        RECT 3.465 8.725 9.665 8.875 ;
        RECT 3.465 8.670 3.785 8.725 ;
        RECT 9.345 8.670 9.665 8.725 ;
        RECT 28.395 7.795 28.675 22.940 ;
        RECT 28.005 7.515 29.065 7.795 ;
        RECT 2.320 7.115 8.170 7.445 ;
        RECT 30.810 7.420 31.160 23.035 ;
        RECT 32.260 21.265 32.580 21.290 ;
        RECT 49.380 21.265 49.700 21.290 ;
        RECT 32.260 21.055 49.700 21.265 ;
        RECT 32.260 21.030 32.580 21.055 ;
        RECT 49.380 21.030 49.700 21.055 ;
        RECT 39.715 20.260 44.220 20.555 ;
        RECT 55.115 16.730 55.520 50.710 ;
        RECT 56.035 38.765 56.310 53.615 ;
        RECT 56.785 38.100 57.030 53.600 ;
        RECT 56.045 37.855 57.030 38.100 ;
        RECT 56.045 23.825 56.290 37.855 ;
        RECT 57.445 37.140 57.770 53.540 ;
        RECT 67.015 48.470 67.365 50.685 ;
        RECT 79.900 50.170 80.470 50.690 ;
        RECT 68.985 48.855 70.550 49.935 ;
        RECT 66.715 48.120 67.665 48.470 ;
        RECT 70.940 46.920 71.215 46.950 ;
        RECT 69.010 46.645 71.215 46.920 ;
        RECT 69.010 44.305 69.285 46.645 ;
        RECT 70.940 46.615 71.215 46.645 ;
        RECT 59.465 40.875 59.785 40.930 ;
        RECT 65.345 40.875 65.665 40.930 ;
        RECT 59.465 40.725 65.665 40.875 ;
        RECT 59.465 40.670 59.785 40.725 ;
        RECT 65.345 40.670 65.665 40.725 ;
        RECT 56.710 36.815 57.770 37.140 ;
        RECT 58.025 39.260 63.910 39.605 ;
        RECT 56.035 22.765 56.295 23.825 ;
        RECT 38.715 16.325 55.520 16.730 ;
        RECT 42.940 14.920 43.215 14.950 ;
        RECT 41.010 14.645 43.215 14.920 ;
        RECT 41.010 12.305 41.285 14.645 ;
        RECT 42.940 14.615 43.215 14.645 ;
        RECT 31.465 8.875 31.785 8.930 ;
        RECT 37.345 8.875 37.665 8.930 ;
        RECT 31.465 8.725 37.665 8.875 ;
        RECT 31.465 8.670 31.785 8.725 ;
        RECT 37.345 8.670 37.665 8.725 ;
        RECT 36.100 7.445 36.380 7.465 ;
        RECT 35.625 7.420 36.405 7.445 ;
        RECT 30.810 7.115 36.405 7.420 ;
        RECT 30.810 7.095 36.380 7.115 ;
        RECT 30.810 7.070 36.225 7.095 ;
        RECT 35.785 7.065 36.225 7.070 ;
        RECT 56.710 6.765 57.035 36.815 ;
        RECT 58.025 23.425 58.370 39.260 ;
        RECT 60.260 37.265 60.580 37.290 ;
        RECT 77.380 37.265 77.700 37.290 ;
        RECT 60.260 37.055 77.700 37.265 ;
        RECT 60.260 37.030 60.580 37.055 ;
        RECT 77.380 37.030 77.700 37.055 ;
        RECT 67.715 36.260 72.220 36.555 ;
        RECT 80.225 34.570 81.600 36.025 ;
        RECT 69.065 33.350 70.415 34.205 ;
        RECT 69.110 33.320 70.370 33.350 ;
        RECT 82.200 32.540 82.540 50.765 ;
        RECT 83.160 37.785 83.555 50.785 ;
        RECT 84.055 39.825 84.275 53.395 ;
        RECT 84.035 38.765 84.295 39.825 ;
        RECT 83.160 37.390 84.285 37.785 ;
        RECT 66.715 32.200 82.540 32.540 ;
        RECT 70.940 30.920 71.215 30.950 ;
        RECT 69.010 30.645 71.215 30.920 ;
        RECT 69.010 28.305 69.285 30.645 ;
        RECT 70.940 30.615 71.215 30.645 ;
        RECT 59.465 24.875 59.785 24.930 ;
        RECT 65.345 24.875 65.665 24.930 ;
        RECT 59.465 24.725 65.665 24.875 ;
        RECT 59.465 24.670 59.785 24.725 ;
        RECT 65.345 24.670 65.665 24.725 ;
        RECT 58.025 23.080 63.960 23.425 ;
        RECT 58.045 7.465 58.390 23.080 ;
        RECT 60.260 21.265 60.580 21.290 ;
        RECT 77.380 21.265 77.700 21.290 ;
        RECT 60.260 21.055 77.700 21.265 ;
        RECT 60.260 21.030 60.580 21.055 ;
        RECT 77.380 21.030 77.700 21.055 ;
        RECT 67.715 20.260 72.220 20.555 ;
        RECT 80.880 18.535 82.255 19.990 ;
        RECT 69.165 16.870 70.310 18.105 ;
        RECT 83.890 16.550 84.285 37.390 ;
        RECT 84.735 22.765 85.035 53.320 ;
        RECT 85.535 52.855 85.900 53.355 ;
        RECT 85.530 22.360 85.900 52.855 ;
        RECT 86.315 47.895 86.620 53.345 ;
        RECT 86.955 48.445 87.280 53.330 ;
        RECT 87.630 49.015 87.935 53.345 ;
        RECT 88.280 49.660 88.625 53.340 ;
        RECT 88.985 50.245 89.335 53.325 ;
        RECT 89.740 51.020 90.130 53.215 ;
        RECT 89.740 50.630 141.735 51.020 ;
        RECT 88.985 49.895 141.035 50.245 ;
        RECT 88.280 49.315 140.380 49.660 ;
        RECT 87.630 48.710 113.550 49.015 ;
        RECT 86.955 48.120 112.960 48.445 ;
        RECT 86.315 47.620 112.340 47.895 ;
        RECT 86.315 47.590 108.230 47.620 ;
        RECT 109.280 47.590 112.340 47.620 ;
        RECT 98.940 46.920 99.215 46.950 ;
        RECT 94.895 46.100 95.660 46.800 ;
        RECT 97.010 46.645 99.215 46.920 ;
        RECT 97.010 44.305 97.285 46.645 ;
        RECT 98.940 46.615 99.215 46.645 ;
        RECT 87.465 40.875 87.785 40.930 ;
        RECT 93.345 40.875 93.665 40.930 ;
        RECT 87.465 40.725 93.665 40.875 ;
        RECT 87.465 40.670 87.785 40.725 ;
        RECT 93.345 40.670 93.665 40.725 ;
        RECT 86.400 39.200 91.945 39.600 ;
        RECT 66.715 16.155 84.285 16.550 ;
        RECT 84.665 21.990 85.900 22.360 ;
        RECT 86.430 23.410 86.830 39.200 ;
        RECT 112.035 38.765 112.340 47.590 ;
        RECT 112.635 37.960 112.960 48.120 ;
        RECT 112.035 37.635 112.960 37.960 ;
        RECT 88.260 37.265 88.580 37.290 ;
        RECT 105.380 37.265 105.700 37.290 ;
        RECT 88.260 37.055 105.700 37.265 ;
        RECT 88.260 37.030 88.580 37.055 ;
        RECT 105.380 37.030 105.700 37.055 ;
        RECT 95.715 36.260 100.220 36.555 ;
        RECT 95.025 31.765 95.790 32.465 ;
        RECT 98.940 30.920 99.215 30.950 ;
        RECT 97.010 30.645 99.215 30.920 ;
        RECT 97.010 28.305 97.285 30.645 ;
        RECT 98.940 30.615 99.215 30.645 ;
        RECT 87.465 24.875 87.785 24.930 ;
        RECT 93.345 24.875 93.665 24.930 ;
        RECT 87.465 24.725 93.665 24.875 ;
        RECT 87.465 24.670 87.785 24.725 ;
        RECT 93.345 24.670 93.665 24.725 ;
        RECT 86.430 23.010 91.975 23.410 ;
        RECT 70.940 14.920 71.215 14.950 ;
        RECT 69.010 14.645 71.215 14.920 ;
        RECT 69.010 12.305 69.285 14.645 ;
        RECT 70.940 14.615 71.215 14.645 ;
        RECT 59.465 8.875 59.785 8.930 ;
        RECT 65.345 8.875 65.665 8.930 ;
        RECT 59.465 8.725 65.665 8.875 ;
        RECT 59.465 8.670 59.785 8.725 ;
        RECT 65.345 8.670 65.665 8.725 ;
        RECT 58.045 7.120 63.920 7.465 ;
        RECT 58.925 7.115 59.685 7.120 ;
        RECT 58.950 7.095 59.230 7.115 ;
        RECT 84.665 6.765 85.035 21.990 ;
        RECT 86.430 7.405 86.830 23.010 ;
        RECT 112.035 22.765 112.360 37.635 ;
        RECT 113.245 37.195 113.550 48.710 ;
        RECT 126.940 46.920 127.215 46.950 ;
        RECT 125.010 46.645 127.215 46.920 ;
        RECT 125.010 44.305 125.285 46.645 ;
        RECT 126.940 46.615 127.215 46.645 ;
        RECT 122.840 43.515 123.515 44.300 ;
        RECT 115.465 40.875 115.785 40.930 ;
        RECT 121.345 40.875 121.665 40.930 ;
        RECT 115.465 40.725 121.665 40.875 ;
        RECT 115.465 40.670 115.785 40.725 ;
        RECT 121.345 40.670 121.665 40.725 ;
        RECT 112.675 36.890 113.550 37.195 ;
        RECT 114.525 39.165 119.880 39.450 ;
        RECT 88.260 21.265 88.580 21.290 ;
        RECT 105.380 21.265 105.700 21.290 ;
        RECT 88.260 21.055 105.700 21.265 ;
        RECT 88.260 21.030 88.580 21.055 ;
        RECT 105.380 21.030 105.700 21.055 ;
        RECT 95.715 20.260 100.220 20.555 ;
        RECT 94.795 15.590 95.560 16.290 ;
        RECT 98.940 14.920 99.215 14.950 ;
        RECT 97.010 14.645 99.215 14.920 ;
        RECT 97.010 12.305 97.285 14.645 ;
        RECT 98.940 14.615 99.215 14.645 ;
        RECT 87.465 8.875 87.785 8.930 ;
        RECT 93.345 8.875 93.665 8.930 ;
        RECT 87.465 8.725 93.665 8.875 ;
        RECT 87.465 8.670 87.785 8.725 ;
        RECT 93.345 8.670 93.665 8.725 ;
        RECT 112.675 7.825 112.980 36.890 ;
        RECT 114.525 23.430 114.810 39.165 ;
        RECT 140.035 38.765 140.380 49.315 ;
        RECT 116.260 37.265 116.580 37.290 ;
        RECT 133.380 37.265 133.700 37.290 ;
        RECT 116.260 37.055 133.700 37.265 ;
        RECT 116.260 37.030 116.580 37.055 ;
        RECT 133.380 37.030 133.700 37.055 ;
        RECT 123.715 36.260 128.220 36.555 ;
        RECT 126.940 30.920 127.215 30.950 ;
        RECT 125.010 30.645 127.215 30.920 ;
        RECT 125.010 28.305 125.285 30.645 ;
        RECT 126.940 30.615 127.215 30.645 ;
        RECT 122.925 27.090 123.600 27.875 ;
        RECT 115.465 24.875 115.785 24.930 ;
        RECT 121.345 24.875 121.665 24.930 ;
        RECT 115.465 24.725 121.665 24.875 ;
        RECT 115.465 24.670 115.785 24.725 ;
        RECT 121.345 24.670 121.665 24.725 ;
        RECT 114.525 23.145 119.895 23.430 ;
        RECT 87.285 7.445 87.565 7.465 ;
        RECT 87.260 7.405 88.160 7.445 ;
        RECT 86.430 7.005 91.945 7.405 ;
        RECT 112.620 6.765 113.035 7.825 ;
        RECT 114.525 7.470 114.810 23.145 ;
        RECT 140.685 22.765 141.035 49.895 ;
        RECT 141.345 22.085 141.735 50.630 ;
        RECT 147.310 48.490 147.715 49.315 ;
        RECT 146.910 48.085 147.715 48.490 ;
        RECT 144.610 46.565 145.040 47.380 ;
        RECT 147.310 47.255 147.715 48.085 ;
        RECT 143.985 46.135 145.040 46.565 ;
        RECT 144.610 45.320 145.040 46.135 ;
        RECT 151.190 45.100 151.955 45.800 ;
        RECT 149.360 43.595 150.375 44.095 ;
        RECT 142.240 42.945 142.680 42.975 ;
        RECT 141.945 42.475 142.680 42.945 ;
        RECT 141.945 27.170 142.385 42.475 ;
        RECT 140.645 21.695 141.735 22.085 ;
        RECT 116.260 21.265 116.580 21.290 ;
        RECT 133.380 21.265 133.700 21.290 ;
        RECT 116.260 21.055 133.700 21.265 ;
        RECT 116.260 21.030 116.580 21.055 ;
        RECT 133.380 21.030 133.700 21.055 ;
        RECT 123.715 20.260 128.220 20.555 ;
        RECT 126.940 14.920 127.215 14.950 ;
        RECT 125.010 14.645 127.215 14.920 ;
        RECT 122.885 13.335 123.560 14.120 ;
        RECT 125.010 12.305 125.285 14.645 ;
        RECT 126.940 14.615 127.215 14.645 ;
        RECT 115.465 8.875 115.785 8.930 ;
        RECT 121.345 8.875 121.665 8.930 ;
        RECT 115.465 8.725 121.665 8.875 ;
        RECT 115.465 8.670 115.785 8.725 ;
        RECT 121.345 8.670 121.665 8.725 ;
        RECT 114.525 7.185 119.885 7.470 ;
        RECT 115.220 7.115 116.010 7.185 ;
        RECT 115.245 7.095 115.525 7.115 ;
        RECT 140.645 6.765 141.035 21.695 ;
        RECT 142.800 13.435 143.300 41.065 ;
        RECT 4.260 5.265 4.580 5.290 ;
        RECT 21.380 5.265 21.700 5.290 ;
        RECT 4.260 5.055 21.700 5.265 ;
        RECT 4.260 5.030 4.580 5.055 ;
        RECT 21.380 5.030 21.700 5.055 ;
        RECT 32.260 5.265 32.580 5.290 ;
        RECT 49.380 5.265 49.700 5.290 ;
        RECT 32.260 5.055 49.700 5.265 ;
        RECT 32.260 5.030 32.580 5.055 ;
        RECT 49.380 5.030 49.700 5.055 ;
        RECT 60.260 5.265 60.580 5.290 ;
        RECT 77.380 5.265 77.700 5.290 ;
        RECT 60.260 5.055 77.700 5.265 ;
        RECT 60.260 5.030 60.580 5.055 ;
        RECT 77.380 5.030 77.700 5.055 ;
        RECT 88.260 5.265 88.580 5.290 ;
        RECT 105.380 5.265 105.700 5.290 ;
        RECT 88.260 5.055 105.700 5.265 ;
        RECT 88.260 5.030 88.580 5.055 ;
        RECT 105.380 5.030 105.700 5.055 ;
        RECT 116.260 5.265 116.580 5.290 ;
        RECT 133.380 5.265 133.700 5.290 ;
        RECT 116.260 5.055 133.700 5.265 ;
        RECT 116.260 5.030 116.580 5.055 ;
        RECT 133.380 5.030 133.700 5.055 ;
        RECT 11.715 4.260 16.220 4.555 ;
        RECT 39.715 4.260 44.220 4.555 ;
        RECT 67.715 4.260 72.220 4.555 ;
        RECT 80.835 2.885 82.210 4.340 ;
        RECT 95.715 4.260 100.220 4.555 ;
        RECT 123.715 4.260 128.220 4.555 ;
      LAYER met3 ;
        RECT 79.900 50.170 80.470 50.690 ;
        RECT 69.085 49.870 70.395 49.875 ;
        RECT 69.055 48.950 70.425 49.870 ;
        RECT 69.085 48.945 70.395 48.950 ;
        RECT 146.930 48.490 147.385 48.515 ;
        RECT 95.065 48.085 147.385 48.490 ;
        RECT 95.065 46.215 95.470 48.085 ;
        RECT 146.930 48.060 147.385 48.085 ;
        RECT 144.005 46.565 144.485 46.590 ;
        RECT 95.985 46.470 107.915 46.565 ;
        RECT 109.595 46.470 144.485 46.565 ;
        RECT 95.985 46.135 144.485 46.470 ;
        RECT 80.225 34.570 81.600 36.025 ;
        RECT 69.085 34.225 70.395 34.230 ;
        RECT 69.055 33.330 70.425 34.225 ;
        RECT 69.085 33.325 70.395 33.330 ;
        RECT 95.985 32.295 96.415 46.135 ;
        RECT 144.005 46.110 144.485 46.135 ;
        RECT 151.245 45.680 151.795 45.705 ;
        RECT 95.115 31.865 96.415 32.295 ;
        RECT 97.190 45.180 151.795 45.680 ;
        RECT 80.880 18.535 82.255 19.990 ;
        RECT 69.080 16.800 70.400 18.180 ;
        RECT 97.190 16.190 97.690 45.180 ;
        RECT 151.245 45.155 151.795 45.180 ;
        RECT 149.380 44.095 149.930 44.120 ;
        RECT 122.915 43.595 149.930 44.095 ;
        RECT 149.380 43.570 149.930 43.595 ;
        RECT 141.920 27.655 142.410 27.680 ;
        RECT 123.010 27.215 142.410 27.655 ;
        RECT 141.920 27.190 142.410 27.215 ;
        RECT 94.950 15.690 97.690 16.190 ;
        RECT 142.775 13.980 143.325 14.005 ;
        RECT 122.980 13.480 143.325 13.980 ;
        RECT 142.775 13.455 143.325 13.480 ;
        RECT 7.770 7.445 8.150 7.470 ;
        RECT 7.770 7.115 143.325 7.445 ;
        RECT 7.770 7.090 8.150 7.115 ;
        RECT 80.835 2.885 82.210 4.340 ;
      LAYER met4 ;
        RECT 30.640 224.970 30.670 225.530 ;
        RECT 30.970 224.970 33.430 225.530 ;
        RECT 33.730 224.970 36.190 225.530 ;
        RECT 36.490 224.970 38.950 225.530 ;
        RECT 42.010 224.920 44.470 225.480 ;
        RECT 44.770 224.920 47.230 225.480 ;
        RECT 47.530 224.920 49.990 225.480 ;
        RECT 45.610 224.910 46.170 224.920 ;
        RECT 53.050 224.840 55.510 225.140 ;
        RECT 55.810 224.840 58.270 225.140 ;
        RECT 58.570 224.840 61.030 225.140 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 52.750 224.560 53.050 224.760 ;
        RECT 1.650 220.760 2.210 220.770 ;
        RECT 6.000 220.440 6.020 220.740 ;
        RECT 6.000 212.060 6.010 213.245 ;
        RECT 80.945 50.625 82.125 50.740 ;
        RECT 79.955 50.230 82.125 50.625 ;
        RECT 3.000 19.330 3.010 23.100 ;
        RECT 69.080 18.155 70.400 49.875 ;
        RECT 80.945 35.855 82.125 50.230 ;
        RECT 80.290 34.675 82.125 35.855 ;
        RECT 69.075 16.825 70.405 18.155 ;
        RECT 80.945 4.270 82.125 34.675 ;
        RECT 80.915 3.030 82.155 4.270 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
        RECT 151.490 1.000 152.930 1.740 ;
        RECT 151.490 0.480 151.810 1.000 ;
        RECT 152.710 0.480 152.930 1.000 ;
  END
END tt_um_adc_dac_tern_alu
END LIBRARY

