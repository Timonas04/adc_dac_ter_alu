magic
tech sky130A
magscale 1 2
timestamp 1757921826
<< viali >>
rect 9873 10761 9907 10795
rect 11713 10761 11747 10795
rect 14289 10761 14323 10795
rect 15117 10761 15151 10795
rect 15577 10761 15611 10795
rect 16129 10761 16163 10795
rect 16957 10761 16991 10795
rect 17601 10761 17635 10795
rect 19533 10761 19567 10795
rect 20913 10761 20947 10795
rect 18429 10693 18463 10727
rect 22937 10693 22971 10727
rect 23305 10693 23339 10727
rect 1685 10625 1719 10659
rect 3893 10625 3927 10659
rect 4169 10625 4203 10659
rect 4261 10625 4295 10659
rect 9137 10625 9171 10659
rect 10057 10625 10091 10659
rect 11069 10625 11103 10659
rect 11897 10625 11931 10659
rect 12265 10625 12299 10659
rect 12725 10625 12759 10659
rect 13001 10625 13035 10659
rect 14105 10625 14139 10659
rect 14657 10625 14691 10659
rect 14933 10625 14967 10659
rect 15301 10625 15335 10659
rect 15761 10625 15795 10659
rect 15945 10625 15979 10659
rect 16497 10625 16531 10659
rect 17141 10625 17175 10659
rect 17417 10625 17451 10659
rect 17785 10625 17819 10659
rect 18061 10625 18095 10659
rect 18613 10625 18647 10659
rect 18797 10625 18831 10659
rect 18889 10625 18923 10659
rect 19717 10625 19751 10659
rect 19993 10625 20027 10659
rect 20545 10625 20579 10659
rect 20821 10625 20855 10659
rect 21097 10625 21131 10659
rect 21465 10625 21499 10659
rect 21833 10625 21867 10659
rect 22385 10625 22419 10659
rect 22569 10625 22603 10659
rect 22661 10625 22695 10659
rect 1777 10557 1811 10591
rect 13277 10557 13311 10591
rect 19809 10557 19843 10591
rect 21189 10557 21223 10591
rect 21649 10557 21683 10591
rect 22477 10557 22511 10591
rect 23121 10557 23155 10591
rect 14841 10489 14875 10523
rect 16313 10489 16347 10523
rect 17877 10489 17911 10523
rect 20177 10489 20211 10523
rect 23213 10489 23247 10523
rect 1501 10421 1535 10455
rect 3985 10421 4019 10455
rect 4445 10421 4479 10455
rect 9321 10421 9355 10455
rect 11253 10421 11287 10455
rect 12449 10421 12483 10455
rect 12633 10421 12667 10455
rect 12909 10421 12943 10455
rect 15485 10421 15519 10455
rect 17233 10421 17267 10455
rect 18245 10421 18279 10455
rect 19073 10421 19107 10455
rect 20453 10421 20487 10455
rect 20637 10421 20671 10455
rect 21281 10421 21315 10455
rect 22017 10421 22051 10455
rect 22845 10421 22879 10455
rect 22937 10421 22971 10455
rect 1961 10217 1995 10251
rect 4077 10217 4111 10251
rect 6101 10217 6135 10251
rect 9965 10217 9999 10251
rect 13921 10217 13955 10251
rect 16497 10217 16531 10251
rect 18797 10217 18831 10251
rect 22109 10217 22143 10251
rect 6193 10149 6227 10183
rect 9873 10149 9907 10183
rect 10333 10149 10367 10183
rect 11713 10149 11747 10183
rect 13553 10149 13587 10183
rect 23029 10149 23063 10183
rect 4721 10081 4755 10115
rect 7021 10081 7055 10115
rect 7757 10081 7791 10115
rect 19349 10081 19383 10115
rect 19717 10081 19751 10115
rect 1685 10013 1719 10047
rect 2145 10013 2179 10047
rect 5273 10013 5307 10047
rect 5825 10013 5859 10047
rect 6469 10013 6503 10047
rect 6561 10013 6595 10047
rect 6745 10013 6779 10047
rect 6837 10013 6871 10047
rect 7113 10013 7147 10047
rect 8217 10013 8251 10047
rect 9505 10013 9539 10047
rect 9597 10013 9631 10047
rect 9873 10013 9907 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 10517 10013 10551 10047
rect 11342 10013 11376 10047
rect 11805 10013 11839 10047
rect 12081 10013 12115 10047
rect 12909 10013 12943 10047
rect 13093 10013 13127 10047
rect 13185 10013 13219 10047
rect 13461 10013 13495 10047
rect 13737 10013 13771 10047
rect 14289 10013 14323 10047
rect 14473 10013 14507 10047
rect 14933 10013 14967 10047
rect 15117 10013 15151 10047
rect 15301 10013 15335 10047
rect 15485 10013 15519 10047
rect 15753 10023 15787 10057
rect 16037 10013 16071 10047
rect 16221 10013 16255 10047
rect 16313 10013 16347 10047
rect 16957 10013 16991 10047
rect 17693 10013 17727 10047
rect 17877 10013 17911 10047
rect 18061 10013 18095 10047
rect 18521 10013 18555 10047
rect 18705 10013 18739 10047
rect 18981 10013 19015 10047
rect 19533 10013 19567 10047
rect 21925 10013 21959 10047
rect 22477 10013 22511 10047
rect 22753 10013 22787 10047
rect 22937 10013 22971 10047
rect 23305 10013 23339 10047
rect 4445 9945 4479 9979
rect 5089 9945 5123 9979
rect 6101 9945 6135 9979
rect 6193 9945 6227 9979
rect 8033 9945 8067 9979
rect 10701 9945 10735 9979
rect 12265 9945 12299 9979
rect 14749 9945 14783 9979
rect 15853 9945 15887 9979
rect 18245 9945 18279 9979
rect 18337 9945 18371 9979
rect 19993 9945 20027 9979
rect 23029 9945 23063 9979
rect 1501 9877 1535 9911
rect 4537 9877 4571 9911
rect 4905 9877 4939 9911
rect 5917 9877 5951 9911
rect 6377 9877 6411 9911
rect 7205 9877 7239 9911
rect 7573 9877 7607 9911
rect 7665 9877 7699 9911
rect 9321 9877 9355 9911
rect 9689 9877 9723 9911
rect 11161 9877 11195 9911
rect 11345 9877 11379 9911
rect 11897 9877 11931 9911
rect 14657 9877 14691 9911
rect 15669 9877 15703 9911
rect 16129 9877 16163 9911
rect 21281 9877 21315 9911
rect 22293 9877 22327 9911
rect 23213 9877 23247 9911
rect 1961 9673 1995 9707
rect 4353 9673 4387 9707
rect 5733 9673 5767 9707
rect 8033 9673 8067 9707
rect 8493 9673 8527 9707
rect 12909 9673 12943 9707
rect 7665 9605 7699 9639
rect 9045 9605 9079 9639
rect 10333 9605 10367 9639
rect 13369 9605 13403 9639
rect 14933 9605 14967 9639
rect 15117 9605 15151 9639
rect 15761 9605 15795 9639
rect 17325 9605 17359 9639
rect 17417 9605 17451 9639
rect 2145 9537 2179 9571
rect 4445 9537 4479 9571
rect 5365 9537 5399 9571
rect 5549 9537 5583 9571
rect 5825 9537 5859 9571
rect 6009 9537 6043 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 7067 9537 7101 9571
rect 7573 9537 7607 9571
rect 8401 9537 8435 9571
rect 8953 9537 8987 9571
rect 9137 9537 9171 9571
rect 9413 9537 9447 9571
rect 9505 9537 9539 9571
rect 9689 9537 9723 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 12449 9537 12483 9571
rect 13277 9537 13311 9571
rect 14289 9537 14323 9571
rect 14473 9537 14507 9571
rect 14565 9537 14599 9571
rect 14841 9537 14875 9571
rect 15577 9537 15611 9571
rect 15669 9537 15703 9571
rect 15945 9537 15979 9571
rect 16037 9537 16071 9571
rect 16221 9537 16255 9571
rect 16313 9537 16347 9571
rect 16681 9537 16715 9571
rect 16773 9537 16807 9571
rect 17207 9537 17241 9571
rect 17509 9537 17543 9571
rect 17785 9537 17819 9571
rect 17963 9537 17997 9571
rect 19809 9537 19843 9571
rect 19993 9537 20027 9571
rect 21465 9537 21499 9571
rect 22017 9537 22051 9571
rect 22293 9537 22327 9571
rect 22477 9537 22511 9571
rect 22753 9537 22787 9571
rect 23029 9537 23063 9571
rect 4537 9469 4571 9503
rect 7757 9469 7791 9503
rect 8585 9469 8619 9503
rect 9873 9469 9907 9503
rect 10241 9469 10275 9503
rect 10517 9469 10551 9503
rect 12541 9469 12575 9503
rect 12725 9469 12759 9503
rect 13553 9469 13587 9503
rect 17049 9469 17083 9503
rect 3985 9401 4019 9435
rect 14105 9401 14139 9435
rect 15393 9401 15427 9435
rect 17785 9401 17819 9435
rect 22937 9401 22971 9435
rect 6193 9333 6227 9367
rect 6561 9333 6595 9367
rect 7021 9333 7055 9367
rect 7205 9333 7239 9367
rect 10057 9333 10091 9367
rect 12081 9333 12115 9367
rect 15117 9333 15151 9367
rect 16037 9333 16071 9367
rect 17693 9333 17727 9367
rect 18521 9333 18555 9367
rect 21833 9333 21867 9367
rect 23213 9333 23247 9367
rect 3065 9129 3099 9163
rect 6837 9129 6871 9163
rect 7205 9129 7239 9163
rect 8493 9129 8527 9163
rect 9505 9129 9539 9163
rect 10885 9129 10919 9163
rect 11713 9129 11747 9163
rect 15025 9129 15059 9163
rect 15945 9129 15979 9163
rect 16497 9129 16531 9163
rect 16681 9129 16715 9163
rect 17417 9129 17451 9163
rect 17693 9129 17727 9163
rect 18521 9129 18555 9163
rect 19993 9129 20027 9163
rect 20729 9129 20763 9163
rect 23213 9129 23247 9163
rect 3525 9061 3559 9095
rect 3801 9061 3835 9095
rect 6285 9061 6319 9095
rect 11161 9061 11195 9095
rect 16221 9061 16255 9095
rect 17325 9061 17359 9095
rect 4445 8993 4479 9027
rect 5273 8993 5307 9027
rect 7665 8993 7699 9027
rect 7757 8993 7791 9027
rect 9229 8993 9263 9027
rect 10609 8993 10643 9027
rect 11805 8993 11839 9027
rect 11989 8993 12023 9027
rect 12541 8993 12575 9027
rect 13829 8993 13863 9027
rect 16957 8993 16991 9027
rect 3249 8925 3283 8959
rect 3341 8925 3375 8959
rect 3617 8925 3651 8959
rect 4721 8925 4755 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 5365 8925 5399 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 6009 8925 6043 8959
rect 6101 8925 6135 8959
rect 6377 8925 6411 8959
rect 6653 8925 6687 8959
rect 8401 8925 8435 8959
rect 8585 8925 8619 8959
rect 9045 8925 9079 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 10241 8925 10275 8959
rect 10424 8925 10458 8959
rect 10517 8925 10551 8959
rect 10793 8925 10827 8959
rect 11342 8925 11376 8959
rect 11897 8925 11931 8959
rect 12081 8925 12115 8959
rect 13553 8925 13587 8959
rect 14841 8925 14875 8959
rect 15117 8925 15151 8959
rect 15393 8925 15427 8959
rect 15577 8925 15611 8959
rect 15669 8925 15703 8959
rect 15785 8925 15819 8959
rect 16037 8925 16071 8959
rect 16313 8925 16347 8959
rect 16497 8925 16531 8959
rect 16773 8925 16807 8959
rect 17049 8925 17083 8959
rect 17141 8925 17175 8959
rect 17601 8925 17635 8959
rect 17877 8925 17911 8959
rect 17969 8925 18003 8959
rect 18153 8925 18187 8959
rect 18705 8925 18739 8959
rect 18797 8925 18831 8959
rect 18981 8925 19015 8959
rect 19073 8925 19107 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 19533 8925 19567 8959
rect 19626 8925 19660 8959
rect 20177 8925 20211 8959
rect 22293 8925 22327 8959
rect 22477 8925 22511 8959
rect 22753 8925 22787 8959
rect 23029 8925 23063 8959
rect 4261 8857 4295 8891
rect 6285 8857 6319 8891
rect 19901 8857 19935 8891
rect 22017 8857 22051 8891
rect 4169 8789 4203 8823
rect 4997 8789 5031 8823
rect 5641 8789 5675 8823
rect 6469 8789 6503 8823
rect 7573 8789 7607 8823
rect 11345 8789 11379 8823
rect 12633 8789 12667 8823
rect 12725 8789 12759 8823
rect 13093 8789 13127 8823
rect 13185 8789 13219 8823
rect 13645 8789 13679 8823
rect 14657 8789 14691 8823
rect 18337 8789 18371 8823
rect 22937 8789 22971 8823
rect 3433 8585 3467 8619
rect 3801 8585 3835 8619
rect 3893 8585 3927 8619
rect 4261 8585 4295 8619
rect 4813 8585 4847 8619
rect 9873 8585 9907 8619
rect 11713 8585 11747 8619
rect 12173 8585 12207 8619
rect 14105 8585 14139 8619
rect 15209 8585 15243 8619
rect 16037 8585 16071 8619
rect 17325 8585 17359 8619
rect 18429 8585 18463 8619
rect 19165 8585 19199 8619
rect 21189 8585 21223 8619
rect 21373 8585 21407 8619
rect 23029 8585 23063 8619
rect 9045 8517 9079 8551
rect 14611 8517 14645 8551
rect 16405 8517 16439 8551
rect 17785 8517 17819 8551
rect 18319 8517 18353 8551
rect 20453 8517 20487 8551
rect 20821 8517 20855 8551
rect 20913 8517 20947 8551
rect 4475 8449 4509 8483
rect 4629 8449 4663 8483
rect 4905 8449 4939 8483
rect 5917 8449 5951 8483
rect 6469 8449 6503 8483
rect 6653 8449 6687 8483
rect 9137 8449 9171 8483
rect 9229 8449 9263 8483
rect 9413 8449 9447 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 12633 8449 12667 8483
rect 12817 8449 12851 8483
rect 14289 8449 14323 8483
rect 14381 8449 14415 8483
rect 14473 8449 14507 8483
rect 14749 8449 14783 8483
rect 15025 8449 15059 8483
rect 15301 8449 15335 8483
rect 15485 8449 15519 8483
rect 15577 8449 15611 8483
rect 15853 8449 15887 8483
rect 16313 8449 16347 8483
rect 16497 8449 16531 8483
rect 16681 8449 16715 8483
rect 16957 8449 16991 8483
rect 17141 8449 17175 8483
rect 17233 8449 17267 8483
rect 17417 8449 17451 8483
rect 17509 8449 17543 8483
rect 17693 8449 17727 8483
rect 17877 8449 17911 8483
rect 18153 8449 18187 8483
rect 18521 8449 18555 8483
rect 19165 8449 19199 8483
rect 19533 8449 19567 8483
rect 19625 8449 19659 8483
rect 19947 8449 19981 8483
rect 20545 8449 20579 8483
rect 20638 8449 20672 8483
rect 21010 8449 21044 8483
rect 21557 8449 21591 8483
rect 21833 8449 21867 8483
rect 22017 8449 22051 8483
rect 22293 8449 22327 8483
rect 22477 8449 22511 8483
rect 22753 8449 22787 8483
rect 22937 8449 22971 8483
rect 23213 8449 23247 8483
rect 4077 8381 4111 8415
rect 9781 8381 9815 8415
rect 12173 8381 12207 8415
rect 14933 8381 14967 8415
rect 15669 8381 15703 8415
rect 18705 8381 18739 8415
rect 18797 8381 18831 8415
rect 19349 8381 19383 8415
rect 20085 8381 20119 8415
rect 6009 8313 6043 8347
rect 6561 8313 6595 8347
rect 8861 8313 8895 8347
rect 16865 8313 16899 8347
rect 22109 8313 22143 8347
rect 9597 8245 9631 8279
rect 11989 8245 12023 8279
rect 12725 8245 12759 8279
rect 17049 8245 17083 8279
rect 18061 8245 18095 8279
rect 3525 8041 3559 8075
rect 4353 8041 4387 8075
rect 5457 8041 5491 8075
rect 6101 8041 6135 8075
rect 7757 8041 7791 8075
rect 8953 8041 8987 8075
rect 12081 8041 12115 8075
rect 15209 8041 15243 8075
rect 15393 8041 15427 8075
rect 15577 8041 15611 8075
rect 18981 8041 19015 8075
rect 23029 8041 23063 8075
rect 3433 7973 3467 8007
rect 4261 7973 4295 8007
rect 6377 7973 6411 8007
rect 6929 7973 6963 8007
rect 7849 7973 7883 8007
rect 8769 7973 8803 8007
rect 12541 7973 12575 8007
rect 12633 7973 12667 8007
rect 13277 7973 13311 8007
rect 16037 7973 16071 8007
rect 3617 7905 3651 7939
rect 4445 7905 4479 7939
rect 5917 7905 5951 7939
rect 6009 7905 6043 7939
rect 6561 7905 6595 7939
rect 7941 7905 7975 7939
rect 9597 7905 9631 7939
rect 12173 7905 12207 7939
rect 13645 7905 13679 7939
rect 14749 7905 14783 7939
rect 18429 7905 18463 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 3341 7837 3375 7871
rect 3801 7837 3835 7871
rect 4169 7837 4203 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 6285 7837 6319 7871
rect 6469 7837 6503 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7021 7837 7055 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 7665 7837 7699 7871
rect 8033 7837 8067 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 9137 7837 9171 7871
rect 9459 7837 9493 7871
rect 9868 7837 9902 7871
rect 10240 7837 10274 7871
rect 10326 7837 10360 7871
rect 11897 7837 11931 7871
rect 11989 7837 12023 7871
rect 12449 7837 12483 7871
rect 12725 7837 12759 7871
rect 13093 7837 13127 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 13553 7837 13587 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14473 7837 14507 7871
rect 14611 7837 14645 7871
rect 15025 7837 15059 7871
rect 16221 7837 16255 7871
rect 16313 7837 16347 7871
rect 16681 7837 16715 7871
rect 16957 7837 16991 7871
rect 17141 7837 17175 7871
rect 17601 7837 17635 7871
rect 17785 7837 17819 7871
rect 17969 7837 18003 7871
rect 18153 7837 18187 7871
rect 18705 7837 18739 7871
rect 18797 7837 18831 7871
rect 21097 7837 21131 7871
rect 23213 7837 23247 7871
rect 7205 7769 7239 7803
rect 8217 7769 8251 7803
rect 8401 7769 8435 7803
rect 9229 7769 9263 7803
rect 9322 7769 9356 7803
rect 9965 7769 9999 7803
rect 10057 7769 10091 7803
rect 14381 7769 14415 7803
rect 14933 7769 14967 7803
rect 15945 7769 15979 7803
rect 18061 7769 18095 7803
rect 18613 7769 18647 7803
rect 19349 7769 19383 7803
rect 21005 7769 21039 7803
rect 3985 7701 4019 7735
rect 9689 7701 9723 7735
rect 12265 7701 12299 7735
rect 12909 7701 12943 7735
rect 15568 7701 15602 7735
rect 16865 7701 16899 7735
rect 18337 7701 18371 7735
rect 22385 7701 22419 7735
rect 4353 7497 4387 7531
rect 5549 7497 5583 7531
rect 6193 7497 6227 7531
rect 6837 7497 6871 7531
rect 9045 7497 9079 7531
rect 14933 7497 14967 7531
rect 15577 7497 15611 7531
rect 17601 7497 17635 7531
rect 21925 7497 21959 7531
rect 3985 7429 4019 7463
rect 5181 7429 5215 7463
rect 5365 7429 5399 7463
rect 6377 7429 6411 7463
rect 13093 7429 13127 7463
rect 14841 7429 14875 7463
rect 15945 7429 15979 7463
rect 17693 7429 17727 7463
rect 21281 7429 21315 7463
rect 22201 7429 22235 7463
rect 22293 7429 22327 7463
rect 1685 7361 1719 7395
rect 3617 7361 3651 7395
rect 4261 7361 4295 7395
rect 4445 7361 4479 7395
rect 5089 7361 5123 7395
rect 5457 7361 5491 7395
rect 5733 7361 5767 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 6745 7361 6779 7395
rect 6929 7361 6963 7395
rect 9321 7361 9355 7395
rect 9413 7361 9447 7395
rect 9781 7361 9815 7395
rect 12449 7361 12483 7395
rect 15117 7361 15151 7395
rect 15209 7361 15243 7395
rect 15301 7361 15335 7395
rect 15485 7361 15519 7395
rect 15761 7361 15795 7395
rect 16221 7361 16255 7395
rect 16497 7361 16531 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 17325 7361 17359 7395
rect 17417 7361 17451 7395
rect 19533 7361 19567 7395
rect 19711 7361 19745 7395
rect 20637 7361 20671 7395
rect 20821 7361 20855 7395
rect 20913 7361 20947 7395
rect 22109 7361 22143 7395
rect 22385 7361 22419 7395
rect 22569 7361 22603 7395
rect 22753 7361 22787 7395
rect 22937 7361 22971 7395
rect 23029 7361 23063 7395
rect 8585 7293 8619 7327
rect 9689 7293 9723 7327
rect 12725 7293 12759 7327
rect 12909 7293 12943 7327
rect 19625 7293 19659 7327
rect 23213 7293 23247 7327
rect 4169 7225 4203 7259
rect 5365 7225 5399 7259
rect 5825 7225 5859 7259
rect 8861 7225 8895 7259
rect 12541 7225 12575 7259
rect 22845 7225 22879 7259
rect 1501 7157 1535 7191
rect 3985 7157 4019 7191
rect 5917 7157 5951 7191
rect 6377 7157 6411 7191
rect 9137 7157 9171 7191
rect 16037 7157 16071 7191
rect 16405 7157 16439 7191
rect 17141 7157 17175 7191
rect 19165 7157 19199 7191
rect 20729 7157 20763 7191
rect 21097 7157 21131 7191
rect 10057 6953 10091 6987
rect 10977 6953 11011 6987
rect 13001 6953 13035 6987
rect 2237 6885 2271 6919
rect 2881 6885 2915 6919
rect 6469 6885 6503 6919
rect 9229 6885 9263 6919
rect 9413 6885 9447 6919
rect 18981 6885 19015 6919
rect 1961 6817 1995 6851
rect 4286 6817 4320 6851
rect 5917 6817 5951 6851
rect 9965 6817 9999 6851
rect 10793 6817 10827 6851
rect 11621 6817 11655 6851
rect 12173 6817 12207 6851
rect 18245 6817 18279 6851
rect 18337 6817 18371 6851
rect 18429 6817 18463 6851
rect 18705 6817 18739 6851
rect 1685 6749 1719 6783
rect 2605 6749 2639 6783
rect 3157 6749 3191 6783
rect 3341 6749 3375 6783
rect 3801 6749 3835 6783
rect 5273 6749 5307 6783
rect 5457 6749 5491 6783
rect 5733 6749 5767 6783
rect 6193 6749 6227 6783
rect 6469 6749 6503 6783
rect 7757 6749 7791 6783
rect 8953 6749 8987 6783
rect 9689 6749 9723 6783
rect 10333 6749 10367 6783
rect 10609 6749 10643 6783
rect 10885 6749 10919 6783
rect 11069 6749 11103 6783
rect 11529 6749 11563 6783
rect 11805 6749 11839 6783
rect 11897 6749 11931 6783
rect 12357 6749 12391 6783
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 12726 6749 12760 6783
rect 12909 6749 12943 6783
rect 13185 6749 13219 6783
rect 13277 6749 13311 6783
rect 13737 6749 13771 6783
rect 14289 6749 14323 6783
rect 14473 6749 14507 6783
rect 14749 6749 14783 6783
rect 14933 6749 14967 6783
rect 15117 6749 15151 6783
rect 17049 6749 17083 6783
rect 17233 6749 17267 6783
rect 18061 6749 18095 6783
rect 18521 6749 18555 6783
rect 18889 6749 18923 6783
rect 19073 6749 19107 6783
rect 21097 6749 21131 6783
rect 23029 6749 23063 6783
rect 4077 6681 4111 6715
rect 6285 6681 6319 6715
rect 13001 6681 13035 6715
rect 14841 6681 14875 6715
rect 16957 6681 16991 6715
rect 19257 6681 19291 6715
rect 22661 6681 22695 6715
rect 1777 6613 1811 6647
rect 2421 6613 2455 6647
rect 3065 6613 3099 6647
rect 3525 6613 3559 6647
rect 4169 6613 4203 6647
rect 4445 6613 4479 6647
rect 7849 6613 7883 6647
rect 10241 6613 10275 6647
rect 10425 6613 10459 6647
rect 12081 6613 12115 6647
rect 13645 6613 13679 6647
rect 13921 6613 13955 6647
rect 14381 6613 14415 6647
rect 14565 6613 14599 6647
rect 15669 6613 15703 6647
rect 17141 6613 17175 6647
rect 20545 6613 20579 6647
rect 23213 6613 23247 6647
rect 1593 6409 1627 6443
rect 1961 6409 1995 6443
rect 4077 6409 4111 6443
rect 9597 6409 9631 6443
rect 9781 6409 9815 6443
rect 10609 6409 10643 6443
rect 13645 6409 13679 6443
rect 14565 6409 14599 6443
rect 4537 6341 4571 6375
rect 12725 6341 12759 6375
rect 15025 6341 15059 6375
rect 15301 6341 15335 6375
rect 20085 6341 20119 6375
rect 20637 6341 20671 6375
rect 21833 6341 21867 6375
rect 21925 6341 21959 6375
rect 1501 6273 1535 6307
rect 2145 6273 2179 6307
rect 3433 6273 3467 6307
rect 3985 6273 4019 6307
rect 4169 6273 4203 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 9137 6273 9171 6307
rect 9643 6273 9677 6307
rect 9965 6273 9999 6307
rect 10241 6273 10275 6307
rect 10977 6273 11011 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 11989 6273 12023 6307
rect 12081 6273 12115 6307
rect 12265 6273 12299 6307
rect 12357 6273 12391 6307
rect 12450 6273 12484 6307
rect 13001 6273 13035 6307
rect 13737 6273 13771 6307
rect 14565 6273 14599 6307
rect 14742 6273 14776 6307
rect 14928 6273 14962 6307
rect 15117 6273 15151 6307
rect 15485 6273 15519 6307
rect 15669 6273 15703 6307
rect 16037 6273 16071 6307
rect 16313 6273 16347 6307
rect 16497 6273 16531 6307
rect 16865 6273 16899 6307
rect 16957 6273 16991 6307
rect 17049 6273 17083 6307
rect 19349 6273 19383 6307
rect 20453 6273 20487 6307
rect 20729 6273 20763 6307
rect 21097 6273 21131 6307
rect 21373 6273 21407 6307
rect 22201 6273 22235 6307
rect 22661 6273 22695 6307
rect 22753 6273 22787 6307
rect 22937 6273 22971 6307
rect 23029 6273 23063 6307
rect 3617 6205 3651 6239
rect 10793 6205 10827 6239
rect 10885 6205 10919 6239
rect 11069 6205 11103 6239
rect 13369 6205 13403 6239
rect 13461 6205 13495 6239
rect 14105 6205 14139 6239
rect 14197 6205 14231 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 17233 6205 17267 6239
rect 17417 6205 17451 6239
rect 22313 6205 22347 6239
rect 4353 6137 4387 6171
rect 4905 6137 4939 6171
rect 11989 6137 12023 6171
rect 4537 6069 4571 6103
rect 5365 6069 5399 6103
rect 9229 6069 9263 6103
rect 10333 6069 10367 6103
rect 10517 6069 10551 6103
rect 14381 6069 14415 6103
rect 15301 6069 15335 6103
rect 16221 6069 16255 6103
rect 16497 6069 16531 6103
rect 18061 6069 18095 6103
rect 22477 6069 22511 6103
rect 23213 6069 23247 6103
rect 5365 5865 5399 5899
rect 8033 5865 8067 5899
rect 8401 5865 8435 5899
rect 9597 5865 9631 5899
rect 12357 5865 12391 5899
rect 13553 5865 13587 5899
rect 13921 5865 13955 5899
rect 14565 5865 14599 5899
rect 15301 5865 15335 5899
rect 16405 5865 16439 5899
rect 18981 5865 19015 5899
rect 20545 5865 20579 5899
rect 1961 5797 1995 5831
rect 4997 5797 5031 5831
rect 10425 5797 10459 5831
rect 13093 5797 13127 5831
rect 14657 5797 14691 5831
rect 18521 5797 18555 5831
rect 21373 5797 21407 5831
rect 4169 5729 4203 5763
rect 5089 5729 5123 5763
rect 10517 5729 10551 5763
rect 11345 5729 11379 5763
rect 15485 5729 15519 5763
rect 17417 5729 17451 5763
rect 1685 5661 1719 5695
rect 2145 5661 2179 5695
rect 4353 5661 4387 5695
rect 4813 5661 4847 5695
rect 5181 5661 5215 5695
rect 5549 5661 5583 5695
rect 5733 5661 5767 5695
rect 7665 5661 7699 5695
rect 7941 5661 7975 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 9873 5661 9907 5695
rect 9965 5661 9999 5695
rect 10057 5661 10091 5695
rect 10241 5661 10275 5695
rect 10333 5661 10367 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 10977 5661 11011 5695
rect 12541 5661 12575 5695
rect 12633 5661 12667 5695
rect 12817 5661 12851 5695
rect 13093 5661 13127 5695
rect 13645 5661 13679 5695
rect 13737 5661 13771 5695
rect 14192 5671 14226 5705
rect 14381 5661 14415 5695
rect 14565 5661 14599 5695
rect 14841 5661 14875 5695
rect 14933 5661 14967 5695
rect 15025 5661 15059 5695
rect 15209 5661 15243 5695
rect 15577 5661 15611 5695
rect 15945 5661 15979 5695
rect 16129 5661 16163 5695
rect 16221 5661 16255 5695
rect 16773 5661 16807 5695
rect 16865 5661 16899 5695
rect 16957 5661 16991 5695
rect 17141 5661 17175 5695
rect 17601 5661 17635 5695
rect 18061 5661 18095 5695
rect 18153 5661 18187 5695
rect 18889 5661 18923 5695
rect 21465 5661 21499 5695
rect 21557 5661 21591 5695
rect 23121 5661 23155 5695
rect 11161 5593 11195 5627
rect 12357 5593 12391 5627
rect 12909 5593 12943 5627
rect 13461 5593 13495 5627
rect 14289 5593 14323 5627
rect 15853 5593 15887 5627
rect 16405 5593 16439 5627
rect 19257 5593 19291 5627
rect 1501 5525 1535 5559
rect 4537 5525 4571 5559
rect 4629 5525 4663 5559
rect 5917 5525 5951 5559
rect 10609 5525 10643 5559
rect 13277 5525 13311 5559
rect 16497 5525 16531 5559
rect 3985 5321 4019 5355
rect 4997 5321 5031 5355
rect 7113 5321 7147 5355
rect 7849 5321 7883 5355
rect 8493 5321 8527 5355
rect 11253 5321 11287 5355
rect 15669 5321 15703 5355
rect 16957 5321 16991 5355
rect 17877 5321 17911 5355
rect 23121 5321 23155 5355
rect 4353 5253 4387 5287
rect 6653 5253 6687 5287
rect 6745 5253 6779 5287
rect 6863 5253 6897 5287
rect 12725 5253 12759 5287
rect 15025 5253 15059 5287
rect 15117 5253 15151 5287
rect 17141 5253 17175 5287
rect 20177 5253 20211 5287
rect 1501 5185 1535 5219
rect 3893 5185 3927 5219
rect 4169 5185 4203 5219
rect 4445 5185 4479 5219
rect 4537 5185 4571 5219
rect 4721 5185 4755 5219
rect 4813 5185 4847 5219
rect 5273 5185 5307 5219
rect 5457 5185 5491 5219
rect 5549 5185 5583 5219
rect 5641 5185 5675 5219
rect 5825 5185 5859 5219
rect 6561 5185 6595 5219
rect 7021 5185 7055 5219
rect 7297 5185 7331 5219
rect 7389 5185 7423 5219
rect 7481 5185 7515 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 8401 5185 8435 5219
rect 8585 5185 8619 5219
rect 11161 5185 11195 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 11897 5185 11931 5219
rect 11989 5185 12023 5219
rect 12173 5185 12207 5219
rect 13001 5185 13035 5219
rect 13369 5185 13403 5219
rect 13645 5185 13679 5219
rect 13921 5185 13955 5219
rect 14473 5185 14507 5219
rect 14933 5185 14967 5219
rect 15301 5185 15335 5219
rect 15577 5185 15611 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 16037 5185 16071 5219
rect 16221 5185 16255 5219
rect 16497 5185 16531 5219
rect 17233 5185 17267 5219
rect 17416 5185 17450 5219
rect 17509 5185 17543 5219
rect 17785 5185 17819 5219
rect 18061 5185 18095 5219
rect 18245 5185 18279 5219
rect 18337 5185 18371 5219
rect 21373 5185 21407 5219
rect 21649 5185 21683 5219
rect 21833 5185 21867 5219
rect 22845 5185 22879 5219
rect 23029 5185 23063 5219
rect 23305 5185 23339 5219
rect 17601 5117 17635 5151
rect 18153 5117 18187 5151
rect 21557 5117 21591 5151
rect 22385 5117 22419 5151
rect 1685 5049 1719 5083
rect 7941 5049 7975 5083
rect 14105 5049 14139 5083
rect 14289 5049 14323 5083
rect 14749 5049 14783 5083
rect 21189 5049 21223 5083
rect 22293 5049 22327 5083
rect 6009 4981 6043 5015
rect 6377 4981 6411 5015
rect 12817 4981 12851 5015
rect 13185 4981 13219 5015
rect 13553 4981 13587 5015
rect 13829 4981 13863 5015
rect 14565 4981 14599 5015
rect 16313 4981 16347 5015
rect 16773 4981 16807 5015
rect 16957 4981 16991 5015
rect 19625 4981 19659 5015
rect 21649 4981 21683 5015
rect 22201 4981 22235 5015
rect 22661 4981 22695 5015
rect 4537 4777 4571 4811
rect 6469 4777 6503 4811
rect 8677 4777 8711 4811
rect 9045 4777 9079 4811
rect 13001 4777 13035 4811
rect 16037 4777 16071 4811
rect 21373 4777 21407 4811
rect 4445 4709 4479 4743
rect 5089 4709 5123 4743
rect 11253 4709 11287 4743
rect 11989 4709 12023 4743
rect 13461 4709 13495 4743
rect 17601 4709 17635 4743
rect 20545 4709 20579 4743
rect 5181 4641 5215 4675
rect 7297 4641 7331 4675
rect 5917 4573 5951 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 6285 4573 6319 4607
rect 7205 4573 7239 4607
rect 7389 4573 7423 4607
rect 7481 4573 7515 4607
rect 7635 4573 7669 4607
rect 8033 4573 8067 4607
rect 8125 4573 8159 4607
rect 8309 4573 8343 4607
rect 8493 4573 8527 4607
rect 9229 4573 9263 4607
rect 10885 4573 10919 4607
rect 11161 4573 11195 4607
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 12265 4573 12299 4607
rect 12357 4573 12391 4607
rect 12450 4573 12484 4607
rect 12822 4573 12856 4607
rect 13185 4573 13219 4607
rect 13645 4573 13679 4607
rect 13737 4573 13771 4607
rect 14289 4573 14323 4607
rect 14443 4573 14477 4607
rect 15025 4573 15059 4607
rect 15301 4573 15335 4607
rect 16221 4573 16255 4607
rect 16405 4573 16439 4607
rect 16497 4573 16531 4607
rect 16957 4573 16991 4607
rect 17049 4573 17083 4607
rect 17233 4573 17267 4607
rect 19073 4573 19107 4607
rect 22845 4573 22879 4607
rect 23029 4573 23063 4607
rect 4077 4505 4111 4539
rect 4721 4505 4755 4539
rect 8401 4505 8435 4539
rect 11253 4505 11287 4539
rect 12633 4505 12667 4539
rect 12725 4505 12759 4539
rect 13461 4505 13495 4539
rect 14657 4505 14691 4539
rect 14933 4505 14967 4539
rect 15761 4505 15795 4539
rect 19257 4505 19291 4539
rect 7849 4437 7883 4471
rect 10701 4437 10735 4471
rect 11069 4437 11103 4471
rect 11437 4437 11471 4471
rect 12173 4437 12207 4471
rect 13277 4437 13311 4471
rect 13921 4437 13955 4471
rect 16589 4437 16623 4471
rect 23213 4437 23247 4471
rect 4997 4233 5031 4267
rect 5549 4233 5583 4267
rect 8677 4233 8711 4267
rect 11729 4233 11763 4267
rect 12189 4233 12223 4267
rect 12817 4233 12851 4267
rect 15209 4233 15243 4267
rect 4261 4165 4295 4199
rect 5641 4165 5675 4199
rect 8861 4165 8895 4199
rect 9045 4165 9079 4199
rect 9597 4165 9631 4199
rect 10885 4165 10919 4199
rect 11529 4165 11563 4199
rect 11989 4165 12023 4199
rect 13001 4165 13035 4199
rect 14841 4165 14875 4199
rect 20821 4165 20855 4199
rect 4077 4097 4111 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 8125 4097 8159 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 8493 4097 8527 4131
rect 8585 4097 8619 4131
rect 9137 4097 9171 4131
rect 9321 4097 9355 4131
rect 9413 4097 9447 4131
rect 9505 4097 9539 4131
rect 9689 4097 9723 4131
rect 11069 4097 11103 4131
rect 11161 4097 11195 4131
rect 12725 4097 12759 4131
rect 13277 4097 13311 4131
rect 13369 4097 13403 4131
rect 13553 4097 13587 4131
rect 13645 4097 13679 4131
rect 14013 4097 14047 4131
rect 14657 4097 14691 4131
rect 15853 4097 15887 4131
rect 16129 4097 16163 4131
rect 16497 4097 16531 4131
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 17785 4097 17819 4131
rect 18337 4097 18371 4131
rect 20453 4097 20487 4131
rect 20545 4097 20579 4131
rect 20913 4097 20947 4131
rect 21005 4097 21039 4131
rect 21189 4097 21223 4131
rect 21281 4097 21315 4131
rect 21378 4097 21412 4131
rect 22477 4097 22511 4131
rect 22661 4097 22695 4131
rect 22845 4097 22879 4131
rect 23121 4097 23155 4131
rect 7665 4029 7699 4063
rect 14933 4029 14967 4063
rect 15669 4029 15703 4063
rect 16037 4029 16071 4063
rect 16221 4029 16255 4063
rect 16313 4029 16347 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 18153 4029 18187 4063
rect 20729 4029 20763 4063
rect 23213 4029 23247 4063
rect 7941 3961 7975 3995
rect 9137 3961 9171 3995
rect 11897 3961 11931 3995
rect 13001 3961 13035 3995
rect 14381 3961 14415 3995
rect 15301 3961 15335 3995
rect 19625 3961 19659 3995
rect 21557 3961 21591 3995
rect 22293 3961 22327 3995
rect 10885 3893 10919 3927
rect 11345 3893 11379 3927
rect 11713 3893 11747 3927
rect 12173 3893 12207 3927
rect 12357 3893 12391 3927
rect 13093 3893 13127 3927
rect 14473 3893 14507 3927
rect 20269 3893 20303 3927
rect 7389 3689 7423 3723
rect 8769 3689 8803 3723
rect 10241 3689 10275 3723
rect 10609 3689 10643 3723
rect 11437 3689 11471 3723
rect 11713 3689 11747 3723
rect 11989 3689 12023 3723
rect 12357 3689 12391 3723
rect 13737 3689 13771 3723
rect 20545 3689 20579 3723
rect 7941 3621 7975 3655
rect 10793 3621 10827 3655
rect 11897 3621 11931 3655
rect 14657 3621 14691 3655
rect 15117 3621 15151 3655
rect 17141 3621 17175 3655
rect 22385 3621 22419 3655
rect 8309 3553 8343 3587
rect 9045 3553 9079 3587
rect 9505 3553 9539 3587
rect 10977 3553 11011 3587
rect 13369 3553 13403 3587
rect 13461 3553 13495 3587
rect 14565 3553 14599 3587
rect 17325 3553 17359 3587
rect 7113 3485 7147 3519
rect 7481 3485 7515 3519
rect 7757 3485 7791 3519
rect 8217 3485 8251 3519
rect 8493 3485 8527 3519
rect 8585 3485 8619 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 9321 3485 9355 3519
rect 9597 3485 9631 3519
rect 9873 3485 9907 3519
rect 10149 3485 10183 3519
rect 10885 3485 10919 3519
rect 11161 3485 11195 3519
rect 11253 3485 11287 3519
rect 11989 3485 12023 3519
rect 12081 3485 12115 3519
rect 12449 3485 12483 3519
rect 12633 3485 12667 3519
rect 12909 3485 12943 3519
rect 13277 3485 13311 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 14197 3485 14231 3519
rect 14381 3485 14415 3519
rect 14933 3485 14967 3519
rect 15301 3485 15335 3519
rect 15485 3485 15519 3519
rect 16037 3485 16071 3519
rect 16497 3485 16531 3519
rect 16681 3485 16715 3519
rect 16773 3485 16807 3519
rect 16866 3485 16900 3519
rect 18981 3485 19015 3519
rect 19257 3485 19291 3519
rect 22937 3485 22971 3519
rect 23121 3485 23155 3519
rect 7389 3417 7423 3451
rect 10425 3417 10459 3451
rect 10641 3417 10675 3451
rect 11529 3417 11563 3451
rect 11729 3417 11763 3451
rect 16221 3417 16255 3451
rect 21097 3417 21131 3451
rect 7205 3349 7239 3383
rect 7573 3349 7607 3383
rect 9689 3349 9723 3383
rect 10057 3349 10091 3383
rect 13093 3349 13127 3383
rect 14473 3349 14507 3383
rect 15669 3349 15703 3383
rect 16129 3349 16163 3383
rect 23029 3349 23063 3383
rect 6653 3145 6687 3179
rect 7849 3145 7883 3179
rect 9229 3145 9263 3179
rect 10517 3145 10551 3179
rect 12173 3145 12207 3179
rect 12541 3145 12575 3179
rect 12725 3145 12759 3179
rect 13277 3145 13311 3179
rect 14105 3145 14139 3179
rect 15209 3145 15243 3179
rect 16773 3145 16807 3179
rect 17969 3145 18003 3179
rect 22293 3145 22327 3179
rect 23213 3145 23247 3179
rect 7665 3077 7699 3111
rect 9413 3077 9447 3111
rect 19349 3077 19383 3111
rect 19533 3077 19567 3111
rect 19901 3077 19935 3111
rect 21649 3077 21683 3111
rect 6837 3009 6871 3043
rect 7021 3009 7055 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 8033 3009 8067 3043
rect 8401 3009 8435 3043
rect 8677 3009 8711 3043
rect 9045 3009 9079 3043
rect 9781 3009 9815 3043
rect 9965 3009 9999 3043
rect 10057 3009 10091 3043
rect 10333 3009 10367 3043
rect 10793 3009 10827 3043
rect 10885 3009 10919 3043
rect 11161 3009 11195 3043
rect 11345 3009 11379 3043
rect 11529 3009 11563 3043
rect 11713 3009 11747 3043
rect 11989 3009 12023 3043
rect 12633 3009 12667 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 13461 3009 13495 3043
rect 13645 3009 13679 3043
rect 13829 3009 13863 3043
rect 14013 3009 14047 3043
rect 14381 3009 14415 3043
rect 16497 3009 16531 3043
rect 16681 3009 16715 3043
rect 17049 3009 17083 3043
rect 19257 3009 19291 3043
rect 22017 3009 22051 3043
rect 22385 3009 22419 3043
rect 22569 3009 22603 3043
rect 22753 3009 22787 3043
rect 23029 3009 23063 3043
rect 8585 2941 8619 2975
rect 10701 2941 10735 2975
rect 11253 2941 11287 2975
rect 13737 2941 13771 2975
rect 14197 2941 14231 2975
rect 17141 2941 17175 2975
rect 21833 2941 21867 2975
rect 14289 2873 14323 2907
rect 1409 2805 1443 2839
rect 8217 2805 8251 2839
rect 9045 2805 9079 2839
rect 11069 2805 11103 2839
rect 12909 2805 12943 2839
rect 14565 2805 14599 2839
rect 19533 2805 19567 2839
rect 19717 2805 19751 2839
rect 4169 2601 4203 2635
rect 6101 2601 6135 2635
rect 7297 2601 7331 2635
rect 7481 2601 7515 2635
rect 8125 2601 8159 2635
rect 15209 2601 15243 2635
rect 18889 2601 18923 2635
rect 23305 2601 23339 2635
rect 4813 2533 4847 2567
rect 8769 2533 8803 2567
rect 9321 2533 9355 2567
rect 11897 2533 11931 2567
rect 13093 2533 13127 2567
rect 22937 2533 22971 2567
rect 6837 2465 6871 2499
rect 19901 2465 19935 2499
rect 21833 2465 21867 2499
rect 22109 2465 22143 2499
rect 23029 2465 23063 2499
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 5917 2397 5951 2431
rect 6929 2397 6963 2431
rect 7297 2397 7331 2431
rect 7941 2397 7975 2431
rect 8585 2397 8619 2431
rect 9137 2397 9171 2431
rect 9505 2397 9539 2431
rect 10057 2397 10091 2431
rect 10793 2397 10827 2431
rect 10885 2397 10919 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 12265 2397 12299 2431
rect 12449 2397 12483 2431
rect 12909 2397 12943 2431
rect 13185 2397 13219 2431
rect 13369 2397 13403 2431
rect 13829 2397 13863 2431
rect 14105 2397 14139 2431
rect 14565 2397 14599 2431
rect 16497 2397 16531 2431
rect 18429 2397 18463 2431
rect 18521 2397 18555 2431
rect 18981 2397 19015 2431
rect 19533 2397 19567 2431
rect 22845 2397 22879 2431
rect 23121 2397 23155 2431
rect 7665 2329 7699 2363
rect 7849 2329 7883 2363
rect 10517 2329 10551 2363
rect 14381 2329 14415 2363
rect 16681 2329 16715 2363
rect 19257 2329 19291 2363
rect 19717 2329 19751 2363
rect 21649 2329 21683 2363
rect 5457 2261 5491 2295
rect 8493 2261 8527 2295
rect 9689 2261 9723 2295
rect 9965 2261 9999 2295
rect 10241 2261 10275 2295
rect 11069 2261 11103 2295
rect 11345 2261 11379 2295
rect 12173 2261 12207 2295
rect 12357 2261 12391 2295
rect 12725 2261 12759 2295
rect 19349 2261 19383 2295
<< metal1 >>
rect 16206 13268 16212 13320
rect 16264 13308 16270 13320
rect 23106 13308 23112 13320
rect 16264 13280 23112 13308
rect 16264 13268 16270 13280
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 16942 11024 16948 11076
rect 17000 11064 17006 11076
rect 20622 11064 20628 11076
rect 17000 11036 20628 11064
rect 17000 11024 17006 11036
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 15010 10996 15016 11008
rect 14240 10968 15016 10996
rect 14240 10956 14246 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 21450 10996 21456 11008
rect 16448 10968 21456 10996
rect 16448 10956 16454 10968
rect 21450 10956 21456 10968
rect 21508 10956 21514 11008
rect 21542 10956 21548 11008
rect 21600 10996 21606 11008
rect 22646 10996 22652 11008
rect 21600 10968 22652 10996
rect 21600 10956 21606 10968
rect 22646 10956 22652 10968
rect 22704 10956 22710 11008
rect 1104 10906 23644 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 23644 10906
rect 1104 10832 23644 10854
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 9861 10795 9919 10801
rect 9861 10792 9873 10795
rect 9732 10764 9873 10792
rect 9732 10752 9738 10764
rect 9861 10761 9873 10764
rect 9907 10761 9919 10795
rect 9861 10755 9919 10761
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11664 10764 11713 10792
rect 11664 10752 11670 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 13538 10752 13544 10804
rect 13596 10792 13602 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 13596 10764 14289 10792
rect 13596 10752 13602 10764
rect 14277 10761 14289 10764
rect 14323 10761 14335 10795
rect 14277 10755 14335 10761
rect 14826 10752 14832 10804
rect 14884 10792 14890 10804
rect 15105 10795 15163 10801
rect 15105 10792 15117 10795
rect 14884 10764 15117 10792
rect 14884 10752 14890 10764
rect 15105 10761 15117 10764
rect 15151 10761 15163 10795
rect 15105 10755 15163 10761
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 15565 10795 15623 10801
rect 15565 10792 15577 10795
rect 15528 10764 15577 10792
rect 15528 10752 15534 10764
rect 15565 10761 15577 10764
rect 15611 10761 15623 10795
rect 15565 10755 15623 10761
rect 16114 10752 16120 10804
rect 16172 10752 16178 10804
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 16945 10795 17003 10801
rect 16945 10792 16957 10795
rect 16816 10764 16957 10792
rect 16816 10752 16822 10764
rect 16945 10761 16957 10764
rect 16991 10761 17003 10795
rect 16945 10755 17003 10761
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 17589 10795 17647 10801
rect 17589 10792 17601 10795
rect 17460 10764 17601 10792
rect 17460 10752 17466 10764
rect 17589 10761 17601 10764
rect 17635 10761 17647 10795
rect 17589 10755 17647 10761
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19521 10795 19579 10801
rect 19521 10792 19533 10795
rect 19392 10764 19533 10792
rect 19392 10752 19398 10764
rect 19521 10761 19533 10764
rect 19567 10761 19579 10795
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 19521 10755 19579 10761
rect 20548 10764 20913 10792
rect 15194 10724 15200 10736
rect 11900 10696 15200 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1946 10656 1952 10668
rect 1719 10628 1952 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3384 10628 3893 10656
rect 3384 10616 3390 10628
rect 3881 10625 3893 10628
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4706 10656 4712 10668
rect 4295 10628 4712 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1360 10560 1777 10588
rect 1360 10548 1366 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 4172 10588 4200 10619
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 9088 10628 9137 10656
rect 9088 10616 9094 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 10008 10628 10057 10656
rect 10008 10616 10014 10628
rect 10045 10625 10057 10628
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 10962 10616 10968 10668
rect 11020 10656 11026 10668
rect 11900 10665 11928 10696
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 17862 10724 17868 10736
rect 15948 10696 17868 10724
rect 11057 10659 11115 10665
rect 11057 10656 11069 10659
rect 11020 10628 11069 10656
rect 11020 10616 11026 10628
rect 11057 10625 11069 10628
rect 11103 10625 11115 10659
rect 11057 10619 11115 10625
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 12250 10616 12256 10668
rect 12308 10616 12314 10668
rect 12710 10616 12716 10668
rect 12768 10616 12774 10668
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12952 10628 13001 10656
rect 12952 10616 12958 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13906 10616 13912 10668
rect 13964 10656 13970 10668
rect 14093 10659 14151 10665
rect 14093 10656 14105 10659
rect 13964 10628 14105 10656
rect 13964 10616 13970 10628
rect 14093 10625 14105 10628
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14642 10616 14648 10668
rect 14700 10616 14706 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14844 10628 14933 10656
rect 4798 10588 4804 10600
rect 4172 10560 4804 10588
rect 1765 10551 1823 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 13078 10548 13084 10600
rect 13136 10588 13142 10600
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 13136 10560 13277 10588
rect 13136 10548 13142 10560
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 5442 10480 5448 10532
rect 5500 10520 5506 10532
rect 12066 10520 12072 10532
rect 5500 10492 12072 10520
rect 5500 10480 5506 10492
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 14844 10529 14872 10628
rect 14921 10625 14933 10628
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 15948 10665 15976 10696
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 18417 10727 18475 10733
rect 18417 10693 18429 10727
rect 18463 10724 18475 10727
rect 20548 10724 20576 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 18463 10696 18828 10724
rect 18463 10693 18475 10696
rect 18417 10687 18475 10693
rect 18800 10668 18828 10696
rect 19812 10696 20576 10724
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 15068 10628 15301 10656
rect 15068 10616 15074 10628
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 15764 10588 15792 10619
rect 16482 10616 16488 10668
rect 16540 10616 16546 10668
rect 17126 10616 17132 10668
rect 17184 10616 17190 10668
rect 17405 10659 17463 10665
rect 17405 10625 17417 10659
rect 17451 10656 17463 10659
rect 17678 10656 17684 10668
rect 17451 10628 17684 10656
rect 17451 10625 17463 10628
rect 17405 10619 17463 10625
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 17770 10616 17776 10668
rect 17828 10616 17834 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18095 10628 18613 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18506 10588 18512 10600
rect 15764 10560 18512 10588
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 18616 10532 18644 10619
rect 18782 10616 18788 10668
rect 18840 10616 18846 10668
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 18892 10588 18920 10619
rect 19702 10616 19708 10668
rect 19760 10616 19766 10668
rect 19812 10597 19840 10696
rect 20548 10665 20576 10696
rect 22462 10684 22468 10736
rect 22520 10724 22526 10736
rect 22738 10724 22744 10736
rect 22520 10696 22744 10724
rect 22520 10684 22526 10696
rect 19981 10659 20039 10665
rect 19981 10625 19993 10659
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 20533 10659 20591 10665
rect 20533 10625 20545 10659
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 19797 10591 19855 10597
rect 19797 10588 19809 10591
rect 18892 10560 19809 10588
rect 19797 10557 19809 10560
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 14829 10523 14887 10529
rect 14829 10489 14841 10523
rect 14875 10489 14887 10523
rect 14829 10483 14887 10489
rect 15396 10492 15976 10520
rect 382 10412 388 10464
rect 440 10452 446 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 440 10424 1501 10452
rect 440 10412 446 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 3973 10455 4031 10461
rect 3973 10421 3985 10455
rect 4019 10452 4031 10455
rect 4062 10452 4068 10464
rect 4019 10424 4068 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 5810 10452 5816 10464
rect 4479 10424 5816 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 9306 10412 9312 10464
rect 9364 10412 9370 10464
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11606 10452 11612 10464
rect 11287 10424 11612 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 12621 10455 12679 10461
rect 12621 10421 12633 10455
rect 12667 10452 12679 10455
rect 12710 10452 12716 10464
rect 12667 10424 12716 10452
rect 12667 10421 12679 10424
rect 12621 10415 12679 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 15396 10452 15424 10492
rect 12943 10424 15424 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 15470 10412 15476 10464
rect 15528 10412 15534 10464
rect 15948 10452 15976 10492
rect 16022 10480 16028 10532
rect 16080 10520 16086 10532
rect 16301 10523 16359 10529
rect 16301 10520 16313 10523
rect 16080 10492 16313 10520
rect 16080 10480 16086 10492
rect 16301 10489 16313 10492
rect 16347 10489 16359 10523
rect 16301 10483 16359 10489
rect 16574 10480 16580 10532
rect 16632 10520 16638 10532
rect 16632 10492 16804 10520
rect 16632 10480 16638 10492
rect 16666 10452 16672 10464
rect 15948 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16776 10452 16804 10492
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 17865 10523 17923 10529
rect 17865 10520 17877 10523
rect 17184 10492 17877 10520
rect 17184 10480 17190 10492
rect 17865 10489 17877 10492
rect 17911 10489 17923 10523
rect 17865 10483 17923 10489
rect 18156 10492 18552 10520
rect 17221 10455 17279 10461
rect 17221 10452 17233 10455
rect 16776 10424 17233 10452
rect 17221 10421 17233 10424
rect 17267 10452 17279 10455
rect 18156 10452 18184 10492
rect 17267 10424 18184 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 18230 10412 18236 10464
rect 18288 10412 18294 10464
rect 18524 10452 18552 10492
rect 18598 10480 18604 10532
rect 18656 10520 18662 10532
rect 18656 10492 19380 10520
rect 18656 10480 18662 10492
rect 18874 10452 18880 10464
rect 18524 10424 18880 10452
rect 18874 10412 18880 10424
rect 18932 10412 18938 10464
rect 19061 10455 19119 10461
rect 19061 10421 19073 10455
rect 19107 10452 19119 10455
rect 19242 10452 19248 10464
rect 19107 10424 19248 10452
rect 19107 10421 19119 10424
rect 19061 10415 19119 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 19352 10452 19380 10492
rect 19518 10480 19524 10532
rect 19576 10520 19582 10532
rect 19996 10520 20024 10619
rect 20806 10616 20812 10668
rect 20864 10616 20870 10668
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 21450 10616 21456 10668
rect 21508 10616 21514 10668
rect 21818 10616 21824 10668
rect 21876 10616 21882 10668
rect 22370 10616 22376 10668
rect 22428 10616 22434 10668
rect 22572 10665 22600 10696
rect 22738 10684 22744 10696
rect 22796 10724 22802 10736
rect 22925 10727 22983 10733
rect 22925 10724 22937 10727
rect 22796 10696 22937 10724
rect 22796 10684 22802 10696
rect 22925 10693 22937 10696
rect 22971 10693 22983 10727
rect 22925 10687 22983 10693
rect 23106 10684 23112 10736
rect 23164 10724 23170 10736
rect 23293 10727 23351 10733
rect 23293 10724 23305 10727
rect 23164 10696 23305 10724
rect 23164 10684 23170 10696
rect 23293 10693 23305 10696
rect 23339 10693 23351 10727
rect 23293 10687 23351 10693
rect 22557 10659 22615 10665
rect 22557 10625 22569 10659
rect 22603 10625 22615 10659
rect 22557 10619 22615 10625
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 21174 10548 21180 10600
rect 21232 10548 21238 10600
rect 21637 10591 21695 10597
rect 21637 10557 21649 10591
rect 21683 10588 21695 10591
rect 22465 10591 22523 10597
rect 22465 10588 22477 10591
rect 21683 10560 22477 10588
rect 21683 10557 21695 10560
rect 21637 10551 21695 10557
rect 22465 10557 22477 10560
rect 22511 10557 22523 10591
rect 22664 10588 22692 10619
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22465 10551 22523 10557
rect 22572 10560 23121 10588
rect 19576 10492 20024 10520
rect 20165 10523 20223 10529
rect 19576 10480 19582 10492
rect 20165 10489 20177 10523
rect 20211 10520 20223 10523
rect 22370 10520 22376 10532
rect 20211 10492 22376 10520
rect 20211 10489 20223 10492
rect 20165 10483 20223 10489
rect 22370 10480 22376 10492
rect 22428 10480 22434 10532
rect 20441 10455 20499 10461
rect 20441 10452 20453 10455
rect 19352 10424 20453 10452
rect 20441 10421 20453 10424
rect 20487 10421 20499 10455
rect 20441 10415 20499 10421
rect 20622 10412 20628 10464
rect 20680 10412 20686 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 21450 10412 21456 10464
rect 21508 10452 21514 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21508 10424 22017 10452
rect 21508 10412 21514 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22572 10452 22600 10560
rect 23109 10557 23121 10560
rect 23155 10557 23167 10591
rect 23109 10551 23167 10557
rect 22646 10480 22652 10532
rect 22704 10520 22710 10532
rect 23201 10523 23259 10529
rect 23201 10520 23213 10523
rect 22704 10492 23213 10520
rect 22704 10480 22710 10492
rect 23201 10489 23213 10492
rect 23247 10489 23259 10523
rect 23201 10483 23259 10489
rect 22152 10424 22600 10452
rect 22152 10412 22158 10424
rect 22830 10412 22836 10464
rect 22888 10412 22894 10464
rect 22922 10412 22928 10464
rect 22980 10412 22986 10464
rect 1104 10362 23644 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 23644 10362
rect 1104 10288 23644 10310
rect 1946 10208 1952 10260
rect 2004 10208 2010 10260
rect 4062 10208 4068 10260
rect 4120 10208 4126 10260
rect 6089 10251 6147 10257
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 6546 10248 6552 10260
rect 6135 10220 6552 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12618 10248 12624 10260
rect 12124 10220 12624 10248
rect 12124 10208 12130 10220
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13906 10208 13912 10260
rect 13964 10208 13970 10260
rect 14660 10220 16436 10248
rect 14660 10192 14688 10220
rect 6181 10183 6239 10189
rect 6181 10149 6193 10183
rect 6227 10180 6239 10183
rect 9861 10183 9919 10189
rect 6227 10152 9720 10180
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 5350 10112 5356 10124
rect 4755 10084 5356 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 7006 10072 7012 10124
rect 7064 10072 7070 10124
rect 7742 10072 7748 10124
rect 7800 10072 7806 10124
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10044 2191 10047
rect 3326 10044 3332 10056
rect 2179 10016 3332 10044
rect 2179 10013 2191 10016
rect 2133 10007 2191 10013
rect 3326 10004 3332 10016
rect 3384 10004 3390 10056
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5442 10044 5448 10056
rect 5307 10016 5448 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5810 10004 5816 10056
rect 5868 10004 5874 10056
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10044 6515 10047
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6503 10016 6561 10044
rect 6503 10013 6515 10016
rect 6457 10007 6515 10013
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 4614 9976 4620 9988
rect 4479 9948 4620 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 5077 9979 5135 9985
rect 5077 9945 5089 9979
rect 5123 9976 5135 9979
rect 5166 9976 5172 9988
rect 5123 9948 5172 9976
rect 5123 9945 5135 9948
rect 5077 9939 5135 9945
rect 5166 9936 5172 9948
rect 5224 9936 5230 9988
rect 6089 9979 6147 9985
rect 6089 9945 6101 9979
rect 6135 9976 6147 9979
rect 6178 9976 6184 9988
rect 6135 9948 6184 9976
rect 6135 9945 6147 9948
rect 6089 9939 6147 9945
rect 6178 9936 6184 9948
rect 6236 9936 6242 9988
rect 6748 9976 6776 10007
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 7098 10004 7104 10056
rect 7156 10004 7162 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 9306 10044 9312 10056
rect 8251 10016 9312 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 6914 9976 6920 9988
rect 6748 9948 6920 9976
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 8021 9979 8079 9985
rect 8021 9976 8033 9979
rect 7576 9948 8033 9976
rect 382 9868 388 9920
rect 440 9908 446 9920
rect 1489 9911 1547 9917
rect 1489 9908 1501 9911
rect 440 9880 1501 9908
rect 440 9868 446 9880
rect 1489 9877 1501 9880
rect 1535 9877 1547 9911
rect 1489 9871 1547 9877
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 4893 9911 4951 9917
rect 4893 9908 4905 9911
rect 4580 9880 4905 9908
rect 4580 9868 4586 9880
rect 4893 9877 4905 9880
rect 4939 9877 4951 9911
rect 4893 9871 4951 9877
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 5776 9880 5917 9908
rect 5776 9868 5782 9880
rect 5905 9877 5917 9880
rect 5951 9908 5963 9911
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 5951 9880 6377 9908
rect 5951 9877 5963 9880
rect 5905 9871 5963 9877
rect 6365 9877 6377 9880
rect 6411 9877 6423 9911
rect 6365 9871 6423 9877
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 7193 9911 7251 9917
rect 7193 9908 7205 9911
rect 6788 9880 7205 9908
rect 6788 9868 6794 9880
rect 7193 9877 7205 9880
rect 7239 9877 7251 9911
rect 7193 9871 7251 9877
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 7576 9917 7604 9948
rect 8021 9945 8033 9948
rect 8067 9945 8079 9979
rect 9508 9976 9536 10007
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 9692 10044 9720 10152
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 10321 10183 10379 10189
rect 10321 10180 10333 10183
rect 9907 10152 10333 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 10321 10149 10333 10152
rect 10367 10149 10379 10183
rect 10321 10143 10379 10149
rect 11701 10183 11759 10189
rect 11701 10149 11713 10183
rect 11747 10180 11759 10183
rect 12894 10180 12900 10192
rect 11747 10152 12900 10180
rect 11747 10149 11759 10152
rect 11701 10143 11759 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13541 10183 13599 10189
rect 13541 10149 13553 10183
rect 13587 10180 13599 10183
rect 14642 10180 14648 10192
rect 13587 10152 14648 10180
rect 13587 10149 13599 10152
rect 13541 10143 13599 10149
rect 14642 10140 14648 10152
rect 14700 10140 14706 10192
rect 14936 10152 16068 10180
rect 11606 10112 11612 10124
rect 11164 10084 11612 10112
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9692 10016 9873 10044
rect 9861 10013 9873 10016
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 10134 10004 10140 10056
rect 10192 10004 10198 10056
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10044 10287 10047
rect 10410 10044 10416 10056
rect 10275 10016 10416 10044
rect 10275 10013 10287 10016
rect 10229 10007 10287 10013
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 11164 10044 11192 10084
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11716 10084 12112 10112
rect 10612 10016 11192 10044
rect 11330 10047 11388 10053
rect 10612 9976 10640 10016
rect 11330 10013 11342 10047
rect 11376 10044 11388 10047
rect 11422 10044 11428 10056
rect 11376 10016 11428 10044
rect 11376 10013 11388 10016
rect 11330 10007 11388 10013
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 9508 9948 10640 9976
rect 8021 9939 8079 9945
rect 10686 9936 10692 9988
rect 10744 9936 10750 9988
rect 11716 9976 11744 10084
rect 12084 10056 12112 10084
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 14936 10112 14964 10152
rect 15378 10112 15384 10124
rect 12492 10084 13216 10112
rect 12492 10072 12498 10084
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 11348 9948 11744 9976
rect 11348 9920 11376 9948
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 7524 9880 7573 9908
rect 7524 9868 7530 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 7561 9871 7619 9877
rect 7650 9868 7656 9920
rect 7708 9868 7714 9920
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 9355 9880 9689 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9677 9877 9689 9880
rect 9723 9908 9735 9911
rect 9766 9908 9772 9920
rect 9723 9880 9772 9908
rect 9723 9877 9735 9880
rect 9677 9871 9735 9877
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 10652 9880 11161 9908
rect 10652 9868 10658 9880
rect 11149 9877 11161 9880
rect 11195 9877 11207 9911
rect 11149 9871 11207 9877
rect 11330 9868 11336 9920
rect 11388 9868 11394 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 11808 9908 11836 10007
rect 12066 10004 12072 10056
rect 12124 10004 12130 10056
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12216 10016 12909 10044
rect 12216 10004 12222 10016
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13188 10053 13216 10084
rect 14292 10084 14964 10112
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 13219 10016 13461 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14292 10053 14320 10084
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 14240 10016 14289 10044
rect 14240 10004 14246 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 14826 10044 14832 10056
rect 14507 10016 14832 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 14826 10004 14832 10016
rect 14884 10004 14890 10056
rect 14936 10053 14964 10084
rect 15120 10084 15384 10112
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 12253 9979 12311 9985
rect 12253 9945 12265 9979
rect 12299 9976 12311 9979
rect 12618 9976 12624 9988
rect 12299 9948 12624 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 13740 9976 13768 10004
rect 14737 9979 14795 9985
rect 14737 9976 14749 9979
rect 12860 9948 13768 9976
rect 14292 9948 14749 9976
rect 12860 9936 12866 9948
rect 14292 9920 14320 9948
rect 14737 9945 14749 9948
rect 14783 9945 14795 9979
rect 14936 9976 14964 10007
rect 15010 10004 15016 10056
rect 15068 10044 15074 10056
rect 15120 10053 15148 10084
rect 15378 10072 15384 10084
rect 15436 10112 15442 10124
rect 15436 10084 15700 10112
rect 15436 10072 15442 10084
rect 15672 10054 15700 10084
rect 15741 10057 15799 10063
rect 15741 10054 15753 10057
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 15068 10016 15117 10044
rect 15068 10004 15074 10016
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10013 15531 10047
rect 15672 10026 15753 10054
rect 15741 10023 15753 10026
rect 15787 10023 15799 10057
rect 16040 10053 16068 10152
rect 16408 10112 16436 10220
rect 16482 10208 16488 10260
rect 16540 10208 16546 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 17828 10220 18797 10248
rect 17828 10208 17834 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 18785 10211 18843 10217
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 21542 10248 21548 10260
rect 18932 10220 21548 10248
rect 18932 10208 18938 10220
rect 21542 10208 21548 10220
rect 21600 10208 21606 10260
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22097 10251 22155 10257
rect 22097 10248 22109 10251
rect 21968 10220 22109 10248
rect 21968 10208 21974 10220
rect 22097 10217 22109 10220
rect 22143 10217 22155 10251
rect 22097 10211 22155 10217
rect 17310 10140 17316 10192
rect 17368 10180 17374 10192
rect 23017 10183 23075 10189
rect 17368 10152 17954 10180
rect 17368 10140 17374 10152
rect 17926 10112 17954 10152
rect 23017 10149 23029 10183
rect 23063 10149 23075 10183
rect 23017 10143 23075 10149
rect 16408 10084 17816 10112
rect 17926 10084 18092 10112
rect 17788 10056 17816 10084
rect 18064 10056 18092 10084
rect 18138 10072 18144 10124
rect 18196 10072 18202 10124
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18288 10084 19012 10112
rect 18288 10072 18294 10084
rect 15741 10017 15799 10023
rect 16025 10047 16083 10053
rect 15473 10007 15531 10013
rect 16025 10013 16037 10047
rect 16071 10013 16083 10047
rect 16025 10007 16083 10013
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10044 16267 10047
rect 16301 10047 16359 10053
rect 16301 10044 16313 10047
rect 16255 10016 16313 10044
rect 16255 10013 16267 10016
rect 16209 10007 16267 10013
rect 16301 10013 16313 10016
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 15304 9976 15332 10007
rect 14936 9948 15332 9976
rect 15488 9976 15516 10007
rect 15841 9979 15899 9985
rect 15841 9976 15853 9979
rect 15488 9948 15853 9976
rect 14737 9939 14795 9945
rect 15841 9945 15853 9948
rect 15887 9976 15899 9979
rect 16224 9976 16252 10007
rect 16942 10004 16948 10056
rect 17000 10004 17006 10056
rect 17681 10047 17739 10053
rect 17681 10013 17693 10047
rect 17727 10013 17739 10047
rect 17681 10007 17739 10013
rect 15887 9948 16252 9976
rect 15887 9945 15899 9948
rect 15841 9939 15899 9945
rect 11885 9911 11943 9917
rect 11885 9908 11897 9911
rect 11756 9880 11897 9908
rect 11756 9868 11762 9880
rect 11885 9877 11897 9880
rect 11931 9877 11943 9911
rect 11885 9871 11943 9877
rect 14274 9868 14280 9920
rect 14332 9868 14338 9920
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 14608 9880 14657 9908
rect 14608 9868 14614 9880
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 14645 9871 14703 9877
rect 15562 9868 15568 9920
rect 15620 9908 15626 9920
rect 15657 9911 15715 9917
rect 15657 9908 15669 9911
rect 15620 9880 15669 9908
rect 15620 9868 15626 9880
rect 15657 9877 15669 9880
rect 15703 9877 15715 9911
rect 15657 9871 15715 9877
rect 15746 9868 15752 9920
rect 15804 9908 15810 9920
rect 16117 9911 16175 9917
rect 16117 9908 16129 9911
rect 15804 9880 16129 9908
rect 15804 9868 15810 9880
rect 16117 9877 16129 9880
rect 16163 9877 16175 9911
rect 17696 9908 17724 10007
rect 17770 10004 17776 10056
rect 17828 10044 17834 10056
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17828 10016 17877 10044
rect 17828 10004 17834 10016
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 18046 10004 18052 10056
rect 18104 10004 18110 10056
rect 18156 10044 18184 10072
rect 18509 10047 18567 10053
rect 18156 10016 18276 10044
rect 18248 9985 18276 10016
rect 18509 10013 18521 10047
rect 18555 10044 18567 10047
rect 18598 10044 18604 10056
rect 18555 10016 18604 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 18782 10044 18788 10056
rect 18739 10016 18788 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 18984 10053 19012 10084
rect 19150 10072 19156 10124
rect 19208 10112 19214 10124
rect 19337 10115 19395 10121
rect 19337 10112 19349 10115
rect 19208 10084 19349 10112
rect 19208 10072 19214 10084
rect 19337 10081 19349 10084
rect 19383 10081 19395 10115
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19337 10075 19395 10081
rect 19444 10084 19717 10112
rect 18969 10047 19027 10053
rect 18969 10013 18981 10047
rect 19015 10013 19027 10047
rect 18969 10007 19027 10013
rect 19058 10004 19064 10056
rect 19116 10044 19122 10056
rect 19444 10044 19472 10084
rect 19705 10081 19717 10084
rect 19751 10112 19763 10115
rect 20622 10112 20628 10124
rect 19751 10084 20628 10112
rect 19751 10081 19763 10084
rect 19705 10075 19763 10081
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 23032 10112 23060 10143
rect 22756 10084 23060 10112
rect 19116 10016 19472 10044
rect 19116 10004 19122 10016
rect 19518 10004 19524 10056
rect 19576 10004 19582 10056
rect 21174 10004 21180 10056
rect 21232 10044 21238 10056
rect 21913 10047 21971 10053
rect 21913 10044 21925 10047
rect 21232 10016 21925 10044
rect 21232 10004 21238 10016
rect 21913 10013 21925 10016
rect 21959 10013 21971 10047
rect 21913 10007 21971 10013
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 22646 10044 22652 10056
rect 22511 10016 22652 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 22756 10053 22784 10084
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10013 22799 10047
rect 22741 10007 22799 10013
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10044 22983 10047
rect 23106 10044 23112 10056
rect 22971 10016 23112 10044
rect 22971 10013 22983 10016
rect 22925 10007 22983 10013
rect 23106 10004 23112 10016
rect 23164 10004 23170 10056
rect 23293 10047 23351 10053
rect 23293 10013 23305 10047
rect 23339 10044 23351 10047
rect 23339 10016 23704 10044
rect 23339 10013 23351 10016
rect 23293 10007 23351 10013
rect 18233 9979 18291 9985
rect 18233 9945 18245 9979
rect 18279 9945 18291 9979
rect 18233 9939 18291 9945
rect 18322 9936 18328 9988
rect 18380 9936 18386 9988
rect 19978 9936 19984 9988
rect 20036 9936 20042 9988
rect 21082 9976 21088 9988
rect 20088 9948 21088 9976
rect 20088 9908 20116 9948
rect 21082 9936 21088 9948
rect 21140 9936 21146 9988
rect 21358 9936 21364 9988
rect 21416 9976 21422 9988
rect 23017 9979 23075 9985
rect 23017 9976 23029 9979
rect 21416 9948 23029 9976
rect 21416 9936 21422 9948
rect 23017 9945 23029 9948
rect 23063 9945 23075 9979
rect 23017 9939 23075 9945
rect 17696 9880 20116 9908
rect 16117 9871 16175 9877
rect 20162 9868 20168 9920
rect 20220 9908 20226 9920
rect 21269 9911 21327 9917
rect 21269 9908 21281 9911
rect 20220 9880 21281 9908
rect 20220 9868 20226 9880
rect 21269 9877 21281 9880
rect 21315 9877 21327 9911
rect 21269 9871 21327 9877
rect 22281 9911 22339 9917
rect 22281 9877 22293 9911
rect 22327 9908 22339 9911
rect 22462 9908 22468 9920
rect 22327 9880 22468 9908
rect 22327 9877 22339 9880
rect 22281 9871 22339 9877
rect 22462 9868 22468 9880
rect 22520 9868 22526 9920
rect 23198 9868 23204 9920
rect 23256 9868 23262 9920
rect 1104 9818 23644 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 23644 9818
rect 1104 9744 23644 9766
rect 1670 9664 1676 9716
rect 1728 9704 1734 9716
rect 1949 9707 2007 9713
rect 1949 9704 1961 9707
rect 1728 9676 1961 9704
rect 1728 9664 1734 9676
rect 1949 9673 1961 9676
rect 1995 9673 2007 9707
rect 1949 9667 2007 9673
rect 4341 9707 4399 9713
rect 4341 9673 4353 9707
rect 4387 9704 4399 9707
rect 4522 9704 4528 9716
rect 4387 9676 4528 9704
rect 4387 9673 4399 9676
rect 4341 9667 4399 9673
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 5718 9664 5724 9716
rect 5776 9664 5782 9716
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6822 9704 6828 9716
rect 6052 9676 6828 9704
rect 6052 9664 6058 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 8021 9707 8079 9713
rect 8021 9704 8033 9707
rect 7064 9676 8033 9704
rect 7064 9664 7070 9676
rect 8021 9673 8033 9676
rect 8067 9673 8079 9707
rect 8021 9667 8079 9673
rect 8478 9664 8484 9716
rect 8536 9664 8542 9716
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 12158 9704 12164 9716
rect 11572 9676 12164 9704
rect 11572 9664 11578 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12434 9704 12440 9716
rect 12268 9676 12440 9704
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5132 9608 6960 9636
rect 5132 9596 5138 9608
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 4614 9568 4620 9580
rect 4479 9540 4620 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 2148 9364 2176 9531
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 5350 9528 5356 9580
rect 5408 9528 5414 9580
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 5368 9500 5396 9528
rect 4571 9472 5396 9500
rect 5552 9500 5580 9531
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 5626 9500 5632 9512
rect 5552 9472 5632 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 5626 9460 5632 9472
rect 5684 9500 5690 9512
rect 6012 9500 6040 9531
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 6932 9568 6960 9608
rect 7650 9596 7656 9648
rect 7708 9636 7714 9648
rect 9033 9639 9091 9645
rect 9033 9636 9045 9639
rect 7708 9608 9045 9636
rect 7708 9596 7714 9608
rect 9033 9605 9045 9608
rect 9079 9605 9091 9639
rect 9858 9636 9864 9648
rect 9033 9599 9091 9605
rect 9416 9608 9864 9636
rect 7006 9568 7012 9580
rect 6932 9540 7012 9568
rect 7006 9528 7012 9540
rect 7064 9577 7070 9580
rect 7064 9571 7113 9577
rect 7064 9537 7067 9571
rect 7101 9537 7113 9571
rect 7064 9531 7113 9537
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 8294 9568 8300 9580
rect 7607 9540 8300 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 7064 9528 7070 9531
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9568 8447 9571
rect 8662 9568 8668 9580
rect 8435 9540 8668 9568
rect 8435 9537 8447 9540
rect 8389 9531 8447 9537
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9568 9183 9571
rect 9214 9568 9220 9580
rect 9171 9540 9220 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 9416 9577 9444 9608
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 10321 9639 10379 9645
rect 10321 9636 10333 9639
rect 10284 9608 10333 9636
rect 10284 9596 10290 9608
rect 10321 9605 10333 9608
rect 10367 9605 10379 9639
rect 10321 9599 10379 9605
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 10410 9568 10416 9580
rect 9723 9540 10416 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 5684 9472 6040 9500
rect 6748 9472 7757 9500
rect 5684 9460 5690 9472
rect 3973 9435 4031 9441
rect 3973 9401 3985 9435
rect 4019 9432 4031 9435
rect 4706 9432 4712 9444
rect 4019 9404 4712 9432
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 5810 9392 5816 9444
rect 5868 9432 5874 9444
rect 6748 9432 6776 9472
rect 7745 9469 7757 9472
rect 7791 9500 7803 9503
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 7791 9472 8585 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 5868 9404 6776 9432
rect 5868 9392 5874 9404
rect 6822 9392 6828 9444
rect 6880 9432 6886 9444
rect 9508 9432 9536 9531
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 12268 9568 12296 9676
rect 12434 9664 12440 9676
rect 12492 9704 12498 9716
rect 12802 9704 12808 9716
rect 12492 9676 12808 9704
rect 12492 9664 12498 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 12894 9664 12900 9716
rect 12952 9664 12958 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13136 9676 16574 9704
rect 13136 9664 13142 9676
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 13357 9639 13415 9645
rect 13357 9636 13369 9639
rect 12400 9608 13369 9636
rect 12400 9596 12406 9608
rect 13357 9605 13369 9608
rect 13403 9605 13415 9639
rect 14921 9639 14979 9645
rect 14921 9636 14933 9639
rect 13357 9599 13415 9605
rect 14476 9608 14933 9636
rect 14476 9580 14504 9608
rect 14921 9605 14933 9608
rect 14967 9605 14979 9639
rect 14921 9599 14979 9605
rect 10836 9540 12296 9568
rect 12437 9571 12495 9577
rect 10836 9528 10842 9540
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10229 9503 10287 9509
rect 10229 9500 10241 9503
rect 9907 9472 10241 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 10229 9469 10241 9472
rect 10275 9469 10287 9503
rect 10229 9463 10287 9469
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9500 10563 9503
rect 10686 9500 10692 9512
rect 10551 9472 10692 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 12250 9460 12256 9512
rect 12308 9500 12314 9512
rect 12452 9500 12480 9531
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 12860 9540 13277 9568
rect 12860 9528 12866 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14148 9540 14289 9568
rect 14148 9528 14154 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14458 9528 14464 9580
rect 14516 9528 14522 9580
rect 14553 9571 14611 9577
rect 14553 9537 14565 9571
rect 14599 9568 14611 9571
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 14599 9540 14841 9568
rect 14599 9537 14611 9540
rect 14553 9531 14611 9537
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14936 9568 14964 9599
rect 15102 9596 15108 9648
rect 15160 9596 15166 9648
rect 15746 9596 15752 9648
rect 15804 9596 15810 9648
rect 16546 9636 16574 9676
rect 16666 9664 16672 9716
rect 16724 9704 16730 9716
rect 23676 9704 23704 10016
rect 16724 9676 23704 9704
rect 16724 9664 16730 9676
rect 17310 9636 17316 9648
rect 15856 9608 16436 9636
rect 16546 9608 17316 9636
rect 14936 9540 15424 9568
rect 14829 9531 14887 9537
rect 12308 9472 12480 9500
rect 12308 9460 12314 9472
rect 12526 9460 12532 9512
rect 12584 9460 12590 9512
rect 12713 9503 12771 9509
rect 12713 9469 12725 9503
rect 12759 9500 12771 9503
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 12759 9472 13553 9500
rect 12759 9469 12771 9472
rect 12713 9463 12771 9469
rect 13541 9469 13553 9472
rect 13587 9500 13599 9503
rect 14844 9500 14872 9531
rect 15396 9500 15424 9540
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15528 9540 15577 9568
rect 15528 9528 15534 9540
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 15856 9568 15884 9608
rect 15712 9540 15884 9568
rect 15712 9528 15718 9540
rect 15930 9528 15936 9580
rect 15988 9528 15994 9580
rect 16022 9528 16028 9580
rect 16080 9528 16086 9580
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 16224 9500 16252 9531
rect 16298 9528 16304 9580
rect 16356 9528 16362 9580
rect 16408 9568 16436 9608
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 17405 9639 17463 9645
rect 17405 9605 17417 9639
rect 17451 9636 17463 9639
rect 18046 9636 18052 9648
rect 17451 9608 17632 9636
rect 17451 9605 17463 9608
rect 17405 9599 17463 9605
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16408 9540 16681 9568
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16758 9528 16764 9580
rect 16816 9528 16822 9580
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17195 9571 17253 9577
rect 17195 9568 17207 9571
rect 16908 9566 17162 9568
rect 17190 9566 17207 9568
rect 16908 9540 17207 9566
rect 16908 9528 16914 9540
rect 17134 9538 17207 9540
rect 17195 9537 17207 9538
rect 17241 9537 17253 9571
rect 17195 9531 17253 9537
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9537 17555 9571
rect 17604 9568 17632 9608
rect 17966 9608 18052 9636
rect 17770 9568 17776 9580
rect 17604 9540 17776 9568
rect 17497 9531 17555 9537
rect 13587 9472 14223 9500
rect 14844 9472 15332 9500
rect 15396 9472 15884 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 6880 9404 9536 9432
rect 6880 9392 6886 9404
rect 11422 9392 11428 9444
rect 11480 9432 11486 9444
rect 12894 9432 12900 9444
rect 11480 9404 12900 9432
rect 11480 9392 11486 9404
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 14056 9404 14105 9432
rect 14056 9392 14062 9404
rect 14093 9401 14105 9404
rect 14139 9401 14151 9435
rect 14195 9432 14223 9472
rect 15304 9432 15332 9472
rect 15381 9435 15439 9441
rect 15381 9432 15393 9435
rect 14195 9404 15240 9432
rect 15304 9404 15393 9432
rect 14093 9395 14151 9401
rect 4062 9364 4068 9376
rect 2148 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9364 4126 9376
rect 4982 9364 4988 9376
rect 4120 9336 4988 9364
rect 4120 9324 4126 9336
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 6086 9324 6092 9376
rect 6144 9364 6150 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 6144 9336 6193 9364
rect 6144 9324 6150 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6420 9336 6561 9364
rect 6420 9324 6426 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 7055 9336 7205 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 9950 9364 9956 9376
rect 7340 9336 9956 9364
rect 7340 9324 7346 9336
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10042 9324 10048 9376
rect 10100 9324 10106 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11848 9336 12081 9364
rect 11848 9324 11854 9336
rect 12069 9333 12081 9336
rect 12115 9333 12127 9367
rect 12069 9327 12127 9333
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 13872 9336 15117 9364
rect 13872 9324 13878 9336
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15212 9364 15240 9404
rect 15381 9401 15393 9404
rect 15427 9401 15439 9435
rect 15856 9432 15884 9472
rect 16132 9472 16252 9500
rect 16132 9432 16160 9472
rect 17034 9460 17040 9512
rect 17092 9460 17098 9512
rect 17512 9500 17540 9531
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17966 9577 17994 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 24486 9636 24492 9648
rect 22020 9608 24492 9636
rect 17951 9571 18009 9577
rect 17951 9537 17963 9571
rect 17997 9537 18009 9571
rect 18690 9568 18696 9580
rect 17951 9531 18009 9537
rect 18064 9540 18696 9568
rect 18064 9512 18092 9540
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19797 9571 19855 9577
rect 19797 9568 19809 9571
rect 19392 9540 19809 9568
rect 19392 9528 19398 9540
rect 19797 9537 19809 9540
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 19981 9571 20039 9577
rect 19981 9537 19993 9571
rect 20027 9568 20039 9571
rect 20162 9568 20168 9580
rect 20027 9540 20168 9568
rect 20027 9537 20039 9540
rect 19981 9531 20039 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 22020 9577 22048 9608
rect 24486 9596 24492 9608
rect 24544 9596 24550 9648
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 20772 9540 21465 9568
rect 20772 9528 20778 9540
rect 21453 9537 21465 9540
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 22005 9571 22063 9577
rect 22005 9537 22017 9571
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9537 22339 9571
rect 22281 9531 22339 9537
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 17134 9472 17540 9500
rect 15856 9404 16160 9432
rect 15381 9395 15439 9401
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 17134 9432 17162 9472
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 21266 9500 21272 9512
rect 18196 9472 21272 9500
rect 18196 9460 18202 9472
rect 21266 9460 21272 9472
rect 21324 9460 21330 9512
rect 22296 9500 22324 9531
rect 22066 9472 22324 9500
rect 16816 9404 17162 9432
rect 16816 9392 16822 9404
rect 17494 9392 17500 9444
rect 17552 9432 17558 9444
rect 17773 9435 17831 9441
rect 17773 9432 17785 9435
rect 17552 9404 17785 9432
rect 17552 9392 17558 9404
rect 17773 9401 17785 9404
rect 17819 9401 17831 9435
rect 17773 9395 17831 9401
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 15212 9336 16037 9364
rect 15105 9327 15163 9333
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 16025 9327 16083 9333
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 17402 9364 17408 9376
rect 16632 9336 17408 9364
rect 16632 9324 16638 9336
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17681 9367 17739 9373
rect 17681 9333 17693 9367
rect 17727 9364 17739 9367
rect 17954 9364 17960 9376
rect 17727 9336 17960 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 18414 9324 18420 9376
rect 18472 9364 18478 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18472 9336 18521 9364
rect 18472 9324 18478 9336
rect 18509 9333 18521 9336
rect 18555 9364 18567 9367
rect 21726 9364 21732 9376
rect 18555 9336 21732 9364
rect 18555 9333 18567 9336
rect 18509 9327 18567 9333
rect 21726 9324 21732 9336
rect 21784 9324 21790 9376
rect 21818 9324 21824 9376
rect 21876 9364 21882 9376
rect 22066 9364 22094 9472
rect 22278 9392 22284 9444
rect 22336 9432 22342 9444
rect 22480 9432 22508 9531
rect 22554 9528 22560 9580
rect 22612 9568 22618 9580
rect 22741 9571 22799 9577
rect 22741 9568 22753 9571
rect 22612 9540 22753 9568
rect 22612 9528 22618 9540
rect 22741 9537 22753 9540
rect 22787 9537 22799 9571
rect 22741 9531 22799 9537
rect 23014 9528 23020 9580
rect 23072 9528 23078 9580
rect 22336 9404 22508 9432
rect 22925 9435 22983 9441
rect 22336 9392 22342 9404
rect 22925 9401 22937 9435
rect 22971 9432 22983 9435
rect 23382 9432 23388 9444
rect 22971 9404 23388 9432
rect 22971 9401 22983 9404
rect 22925 9395 22983 9401
rect 23382 9392 23388 9404
rect 23440 9392 23446 9444
rect 21876 9336 22094 9364
rect 21876 9324 21882 9336
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 23201 9367 23259 9373
rect 23201 9364 23213 9367
rect 22704 9336 23213 9364
rect 22704 9324 22710 9336
rect 23201 9333 23213 9336
rect 23247 9333 23259 9367
rect 23201 9327 23259 9333
rect 1104 9274 23644 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 23644 9274
rect 1104 9200 23644 9222
rect 3053 9163 3111 9169
rect 3053 9129 3065 9163
rect 3099 9160 3111 9163
rect 5902 9160 5908 9172
rect 3099 9132 5908 9160
rect 3099 9129 3111 9132
rect 3053 9123 3111 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6822 9120 6828 9172
rect 6880 9120 6886 9172
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 6972 9132 7205 9160
rect 6972 9120 6978 9132
rect 7193 9129 7205 9132
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 8478 9120 8484 9172
rect 8536 9120 8542 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 9582 9160 9588 9172
rect 9539 9132 9588 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10560 9132 10885 9160
rect 10560 9120 10566 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 10873 9123 10931 9129
rect 11698 9120 11704 9172
rect 11756 9120 11762 9172
rect 13538 9160 13544 9172
rect 12406 9132 13544 9160
rect 3513 9095 3571 9101
rect 3513 9061 3525 9095
rect 3559 9092 3571 9095
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 3559 9064 3801 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 3789 9061 3801 9064
rect 3835 9061 3847 9095
rect 5350 9092 5356 9104
rect 3789 9055 3847 9061
rect 4448 9064 5356 9092
rect 4448 9033 4476 9064
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 6270 9052 6276 9104
rect 6328 9052 6334 9104
rect 8496 9092 8524 9120
rect 7668 9064 8524 9092
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 5074 9024 5080 9036
rect 4433 8987 4491 8993
rect 4632 8996 5080 9024
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3326 8916 3332 8968
rect 3384 8916 3390 8968
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 4356 8956 4476 8958
rect 4632 8956 4660 8996
rect 5074 8984 5080 8996
rect 5132 9024 5138 9036
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 5132 8996 5273 9024
rect 5132 8984 5138 8996
rect 5261 8993 5273 8996
rect 5307 8993 5319 9027
rect 7282 9024 7288 9036
rect 5261 8987 5319 8993
rect 5552 8996 7288 9024
rect 5552 8968 5580 8996
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7668 9033 7696 9064
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 9306 9092 9312 9104
rect 8904 9064 9312 9092
rect 8904 9052 8910 9064
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 11149 9095 11207 9101
rect 11149 9092 11161 9095
rect 10612 9064 11161 9092
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 8993 7711 9027
rect 7653 8987 7711 8993
rect 7742 8984 7748 9036
rect 7800 8984 7806 9036
rect 8938 9024 8944 9036
rect 8404 8996 8944 9024
rect 3651 8930 4660 8956
rect 3651 8928 4384 8930
rect 4448 8928 4660 8930
rect 4709 8959 4767 8965
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 4709 8925 4721 8959
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8956 4859 8959
rect 4982 8956 4988 8968
rect 4847 8928 4988 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 3786 8848 3792 8900
rect 3844 8888 3850 8900
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 3844 8860 4261 8888
rect 3844 8848 3850 8860
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 4724 8888 4752 8919
rect 4982 8916 4988 8928
rect 5040 8956 5046 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 5040 8928 5181 8956
rect 5040 8916 5046 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8956 5411 8959
rect 5534 8956 5540 8968
rect 5399 8928 5540 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 5368 8888 5396 8919
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5718 8916 5724 8968
rect 5776 8916 5782 8968
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5960 8928 6009 8956
rect 5960 8916 5966 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 8294 8956 8300 8968
rect 6687 8928 8300 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 4724 8860 5396 8888
rect 4249 8851 4307 8857
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 4985 8823 5043 8829
rect 4985 8820 4997 8823
rect 4856 8792 4997 8820
rect 4856 8780 4862 8792
rect 4985 8789 4997 8792
rect 5031 8789 5043 8823
rect 4985 8783 5043 8789
rect 5626 8780 5632 8832
rect 5684 8780 5690 8832
rect 6104 8820 6132 8916
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 6273 8891 6331 8897
rect 6273 8888 6285 8891
rect 6236 8860 6285 8888
rect 6236 8848 6242 8860
rect 6273 8857 6285 8860
rect 6319 8888 6331 8891
rect 6656 8888 6684 8919
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8404 8965 8432 8996
rect 8938 8984 8944 8996
rect 8996 9024 9002 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8996 8996 9229 9024
rect 8996 8984 9002 8996
rect 9217 8993 9229 8996
rect 9263 9024 9275 9027
rect 9582 9024 9588 9036
rect 9263 8996 9588 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 10612 9033 10640 9064
rect 11149 9061 11161 9064
rect 11195 9061 11207 9095
rect 12406 9092 12434 9132
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 15010 9120 15016 9172
rect 15068 9120 15074 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 15470 9160 15476 9172
rect 15160 9132 15476 9160
rect 15160 9120 15166 9132
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16298 9160 16304 9172
rect 15979 9132 16304 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16448 9132 16497 9160
rect 16448 9120 16454 9132
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 16485 9123 16543 9129
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 17402 9120 17408 9172
rect 17460 9120 17466 9172
rect 17678 9120 17684 9172
rect 17736 9120 17742 9172
rect 18506 9120 18512 9172
rect 18564 9120 18570 9172
rect 18708 9132 19334 9160
rect 12802 9092 12808 9104
rect 11149 9055 11207 9061
rect 11716 9064 12434 9092
rect 12469 9064 12808 9092
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 8993 10655 9027
rect 11514 9024 11520 9036
rect 10597 8987 10655 8993
rect 10704 8996 11520 9024
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 6319 8860 6684 8888
rect 6319 8857 6331 8860
rect 6273 8851 6331 8857
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 8404 8888 8432 8919
rect 8076 8860 8432 8888
rect 8588 8888 8616 8919
rect 9030 8916 9036 8968
rect 9088 8916 9094 8968
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8956 9367 8959
rect 9398 8956 9404 8968
rect 9355 8928 9404 8956
rect 9355 8925 9367 8928
rect 9309 8919 9367 8925
rect 9324 8888 9352 8919
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 10410 8916 10416 8968
rect 10468 8916 10474 8968
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8956 10563 8959
rect 10704 8956 10732 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 10551 8928 10732 8956
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 10778 8916 10784 8968
rect 10836 8916 10842 8968
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 11330 8959 11388 8965
rect 11330 8956 11342 8959
rect 10928 8928 11342 8956
rect 10928 8916 10934 8928
rect 11330 8925 11342 8928
rect 11376 8956 11388 8959
rect 11716 8956 11744 9064
rect 11790 8984 11796 9036
rect 11848 8984 11854 9036
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 9024 12035 9027
rect 12469 9024 12497 9064
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 15194 9052 15200 9104
rect 15252 9092 15258 9104
rect 16022 9092 16028 9104
rect 15252 9064 16028 9092
rect 15252 9052 15258 9064
rect 16022 9052 16028 9064
rect 16080 9052 16086 9104
rect 16206 9052 16212 9104
rect 16264 9052 16270 9104
rect 17034 9092 17040 9104
rect 16546 9064 17040 9092
rect 12023 8996 12497 9024
rect 12529 9027 12587 9033
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 12529 8993 12541 9027
rect 12575 9024 12587 9027
rect 13814 9024 13820 9036
rect 12575 8996 13820 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 16546 9024 16574 9064
rect 17034 9052 17040 9064
rect 17092 9052 17098 9104
rect 17310 9052 17316 9104
rect 17368 9052 17374 9104
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 18322 9092 18328 9104
rect 17828 9064 18328 9092
rect 17828 9052 17834 9064
rect 18322 9052 18328 9064
rect 18380 9052 18386 9104
rect 16316 8996 16574 9024
rect 11376 8928 11744 8956
rect 11376 8925 11388 8928
rect 11330 8919 11388 8925
rect 11882 8916 11888 8968
rect 11940 8916 11946 8968
rect 12066 8916 12072 8968
rect 12124 8916 12130 8968
rect 12250 8916 12256 8968
rect 12308 8956 12314 8968
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 12308 8928 13553 8956
rect 12308 8916 12314 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 14550 8916 14556 8968
rect 14608 8956 14614 8968
rect 14829 8959 14887 8965
rect 14829 8956 14841 8959
rect 14608 8928 14841 8956
rect 14608 8916 14614 8928
rect 14829 8925 14841 8928
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15102 8956 15108 8968
rect 14976 8928 15108 8956
rect 14976 8916 14982 8928
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15252 8928 15393 8956
rect 15252 8916 15258 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 15562 8916 15568 8968
rect 15620 8916 15626 8968
rect 15654 8916 15660 8968
rect 15712 8916 15718 8968
rect 15746 8916 15752 8968
rect 15804 8965 15810 8968
rect 15804 8959 15831 8965
rect 15819 8925 15831 8959
rect 15804 8919 15831 8925
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 16114 8956 16120 8968
rect 16071 8928 16120 8956
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 15804 8916 15810 8919
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16316 8965 16344 8996
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 16724 8996 16957 9024
rect 16724 8984 16730 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 17494 9024 17500 9036
rect 16945 8987 17003 8993
rect 17052 8996 17500 9024
rect 17052 8968 17080 8996
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8925 16359 8959
rect 16301 8919 16359 8925
rect 16482 8916 16488 8968
rect 16540 8916 16546 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 16761 8959 16819 8965
rect 16632 8952 16712 8956
rect 16761 8952 16773 8959
rect 16632 8928 16773 8952
rect 16632 8916 16638 8928
rect 16684 8925 16773 8928
rect 16807 8925 16819 8959
rect 16684 8924 16819 8925
rect 16761 8919 16819 8924
rect 17034 8916 17040 8968
rect 17092 8916 17098 8968
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8956 17187 8959
rect 17175 8928 17540 8956
rect 17175 8925 17187 8928
rect 17129 8919 17187 8925
rect 8588 8860 9352 8888
rect 10244 8888 10272 8916
rect 12986 8888 12992 8900
rect 10244 8860 12992 8888
rect 8076 8848 8082 8860
rect 12986 8848 12992 8860
rect 13044 8848 13050 8900
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 17512 8888 17540 8928
rect 17586 8916 17592 8968
rect 17644 8916 17650 8968
rect 17862 8916 17868 8968
rect 17920 8916 17926 8968
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18046 8956 18052 8968
rect 18003 8928 18052 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 18230 8956 18236 8968
rect 18187 8928 18236 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 18708 8965 18736 9132
rect 18782 9052 18788 9104
rect 18840 9052 18846 9104
rect 19306 9092 19334 9132
rect 19702 9120 19708 9172
rect 19760 9160 19766 9172
rect 19981 9163 20039 9169
rect 19981 9160 19993 9163
rect 19760 9132 19993 9160
rect 19760 9120 19766 9132
rect 19981 9129 19993 9132
rect 20027 9129 20039 9163
rect 19981 9123 20039 9129
rect 20714 9120 20720 9172
rect 20772 9120 20778 9172
rect 23201 9163 23259 9169
rect 23201 9129 23213 9163
rect 23247 9160 23259 9163
rect 23842 9160 23848 9172
rect 23247 9132 23848 9160
rect 23247 9129 23259 9132
rect 23201 9123 23259 9129
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 20990 9092 20996 9104
rect 19306 9064 20996 9092
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 18799 8965 18827 9052
rect 19536 8996 20392 9024
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 18966 8916 18972 8968
rect 19024 8916 19030 8968
rect 19058 8916 19064 8968
rect 19116 8916 19122 8968
rect 19150 8916 19156 8968
rect 19208 8956 19214 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 19208 8928 19257 8956
rect 19208 8916 19214 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19426 8916 19432 8968
rect 19484 8916 19490 8968
rect 19536 8965 19564 8996
rect 19521 8959 19579 8965
rect 19521 8925 19533 8959
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 20165 8959 20223 8965
rect 20165 8956 20177 8959
rect 19668 8928 19713 8956
rect 20088 8928 20177 8956
rect 19668 8916 19674 8928
rect 19794 8888 19800 8900
rect 13320 8860 16574 8888
rect 17512 8860 19800 8888
rect 13320 8848 13326 8860
rect 6457 8823 6515 8829
rect 6457 8820 6469 8823
rect 6104 8792 6469 8820
rect 6457 8789 6469 8792
rect 6503 8789 6515 8823
rect 6457 8783 6515 8789
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 8662 8820 8668 8832
rect 7607 8792 8668 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 11146 8820 11152 8832
rect 9180 8792 11152 8820
rect 9180 8780 9186 8792
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 11330 8780 11336 8832
rect 11388 8780 11394 8832
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 11882 8820 11888 8832
rect 11480 8792 11888 8820
rect 11480 8780 11486 8792
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 12066 8780 12072 8832
rect 12124 8820 12130 8832
rect 12342 8820 12348 8832
rect 12124 8792 12348 8820
rect 12124 8780 12130 8792
rect 12342 8780 12348 8792
rect 12400 8820 12406 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 12400 8792 12633 8820
rect 12400 8780 12406 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 12621 8783 12679 8789
rect 12713 8823 12771 8829
rect 12713 8789 12725 8823
rect 12759 8820 12771 8823
rect 12802 8820 12808 8832
rect 12759 8792 12808 8820
rect 12759 8789 12771 8792
rect 12713 8783 12771 8789
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13078 8780 13084 8832
rect 13136 8780 13142 8832
rect 13170 8780 13176 8832
rect 13228 8780 13234 8832
rect 13630 8780 13636 8832
rect 13688 8780 13694 8832
rect 14642 8780 14648 8832
rect 14700 8780 14706 8832
rect 16546 8820 16574 8860
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 19886 8848 19892 8900
rect 19944 8848 19950 8900
rect 16850 8820 16856 8832
rect 16546 8792 16856 8820
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17954 8820 17960 8832
rect 17368 8792 17960 8820
rect 17368 8780 17374 8792
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 18325 8823 18383 8829
rect 18325 8789 18337 8823
rect 18371 8820 18383 8823
rect 18966 8820 18972 8832
rect 18371 8792 18972 8820
rect 18371 8789 18383 8792
rect 18325 8783 18383 8789
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 20088 8820 20116 8928
rect 20165 8925 20177 8928
rect 20211 8925 20223 8959
rect 20364 8956 20392 8996
rect 22370 8984 22376 9036
rect 22428 9024 22434 9036
rect 22428 8996 23060 9024
rect 22428 8984 22434 8996
rect 21910 8956 21916 8968
rect 20364 8928 21916 8956
rect 20165 8919 20223 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 22094 8916 22100 8968
rect 22152 8956 22158 8968
rect 22281 8959 22339 8965
rect 22281 8956 22293 8959
rect 22152 8928 22293 8956
rect 22152 8916 22158 8928
rect 22281 8925 22293 8928
rect 22327 8925 22339 8959
rect 22281 8919 22339 8925
rect 22462 8916 22468 8968
rect 22520 8916 22526 8968
rect 22738 8916 22744 8968
rect 22796 8916 22802 8968
rect 23032 8965 23060 8996
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8925 23075 8959
rect 23017 8919 23075 8925
rect 22005 8891 22063 8897
rect 22005 8857 22017 8891
rect 22051 8888 22063 8891
rect 22186 8888 22192 8900
rect 22051 8860 22192 8888
rect 22051 8857 22063 8860
rect 22005 8851 22063 8857
rect 22186 8848 22192 8860
rect 22244 8848 22250 8900
rect 19300 8792 20116 8820
rect 19300 8780 19306 8792
rect 20254 8780 20260 8832
rect 20312 8820 20318 8832
rect 21358 8820 21364 8832
rect 20312 8792 21364 8820
rect 20312 8780 20318 8792
rect 21358 8780 21364 8792
rect 21416 8780 21422 8832
rect 22830 8780 22836 8832
rect 22888 8820 22894 8832
rect 22925 8823 22983 8829
rect 22925 8820 22937 8823
rect 22888 8792 22937 8820
rect 22888 8780 22894 8792
rect 22925 8789 22937 8792
rect 22971 8789 22983 8823
rect 22925 8783 22983 8789
rect 1104 8730 23644 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 23644 8730
rect 1104 8656 23644 8678
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 3421 8619 3479 8625
rect 3421 8616 3433 8619
rect 3292 8588 3433 8616
rect 3292 8576 3298 8588
rect 3421 8585 3433 8588
rect 3467 8585 3479 8619
rect 3421 8579 3479 8585
rect 3786 8576 3792 8628
rect 3844 8576 3850 8628
rect 3881 8619 3939 8625
rect 3881 8585 3893 8619
rect 3927 8616 3939 8619
rect 4154 8616 4160 8628
rect 3927 8588 4160 8616
rect 3927 8585 3939 8588
rect 3881 8579 3939 8585
rect 4154 8576 4160 8588
rect 4212 8616 4218 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4212 8588 4261 8616
rect 4212 8576 4218 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4249 8579 4307 8585
rect 4356 8588 4813 8616
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4356 8548 4384 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 7742 8616 7748 8628
rect 5408 8588 7748 8616
rect 5408 8576 5414 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 7852 8588 9674 8616
rect 5442 8548 5448 8560
rect 4120 8520 4384 8548
rect 4632 8520 5448 8548
rect 4120 8508 4126 8520
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 4632 8489 4660 8520
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 7006 8548 7012 8560
rect 5552 8520 7012 8548
rect 4463 8483 4521 8489
rect 4463 8480 4475 8483
rect 3936 8452 4475 8480
rect 3936 8440 3942 8452
rect 4463 8449 4475 8452
rect 4509 8449 4521 8483
rect 4463 8443 4521 8449
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 4798 8480 4804 8492
rect 4663 8452 4804 8480
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 5552 8480 5580 8520
rect 7006 8508 7012 8520
rect 7064 8548 7070 8560
rect 7852 8548 7880 8588
rect 9646 8560 9674 8588
rect 9858 8576 9864 8628
rect 9916 8576 9922 8628
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8585 11759 8619
rect 11701 8579 11759 8585
rect 12161 8619 12219 8625
rect 12161 8585 12173 8619
rect 12207 8616 12219 8619
rect 12526 8616 12532 8628
rect 12207 8588 12532 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 7064 8520 7880 8548
rect 7064 8508 7070 8520
rect 8846 8508 8852 8560
rect 8904 8548 8910 8560
rect 9033 8551 9091 8557
rect 9033 8548 9045 8551
rect 8904 8520 9045 8548
rect 8904 8508 8910 8520
rect 9033 8517 9045 8520
rect 9079 8517 9091 8551
rect 9646 8520 9680 8560
rect 9033 8511 9091 8517
rect 9674 8508 9680 8520
rect 9732 8548 9738 8560
rect 10594 8548 10600 8560
rect 9732 8520 10600 8548
rect 9732 8508 9738 8520
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 11716 8548 11744 8579
rect 12526 8576 12532 8588
rect 12584 8616 12590 8628
rect 13630 8616 13636 8628
rect 12584 8588 13636 8616
rect 12584 8576 12590 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 14090 8576 14096 8628
rect 14148 8576 14154 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 15197 8619 15255 8625
rect 14516 8588 14780 8616
rect 14516 8576 14522 8588
rect 12250 8548 12256 8560
rect 11716 8520 12256 8548
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 14642 8557 14648 8560
rect 14599 8551 14648 8557
rect 14599 8517 14611 8551
rect 14645 8517 14648 8551
rect 14599 8511 14648 8517
rect 14642 8508 14648 8511
rect 14700 8508 14706 8560
rect 5040 8452 5580 8480
rect 5040 8440 5046 8452
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5684 8452 5917 8480
rect 5684 8440 5690 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6454 8440 6460 8492
rect 6512 8440 6518 8492
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9447 8452 9505 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8412 4123 8415
rect 5350 8412 5356 8424
rect 4111 8384 5356 8412
rect 4111 8381 4123 8384
rect 4065 8375 4123 8381
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 8938 8412 8944 8424
rect 6012 8384 8944 8412
rect 5902 8304 5908 8356
rect 5960 8344 5966 8356
rect 6012 8353 6040 8384
rect 8938 8372 8944 8384
rect 8996 8412 9002 8424
rect 9140 8412 9168 8443
rect 8996 8384 9168 8412
rect 9232 8412 9260 8443
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9640 8452 9873 8480
rect 9640 8440 9646 8452
rect 9861 8449 9873 8452
rect 9907 8480 9919 8483
rect 11422 8480 11428 8492
rect 9907 8452 11428 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 11422 8440 11428 8452
rect 11480 8480 11486 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11480 8452 11529 8480
rect 11480 8440 11486 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 9232 8384 9444 8412
rect 8996 8372 9002 8384
rect 9416 8356 9444 8384
rect 9766 8372 9772 8424
rect 9824 8372 9830 8424
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 11716 8412 11744 8443
rect 11204 8384 11744 8412
rect 11204 8372 11210 8384
rect 5997 8347 6055 8353
rect 5997 8344 6009 8347
rect 5960 8316 6009 8344
rect 5960 8304 5966 8316
rect 5997 8313 6009 8316
rect 6043 8313 6055 8347
rect 5997 8307 6055 8313
rect 6086 8304 6092 8356
rect 6144 8344 6150 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6144 8316 6561 8344
rect 6144 8304 6150 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8849 8347 8907 8353
rect 8849 8344 8861 8347
rect 8260 8316 8861 8344
rect 8260 8304 8266 8316
rect 8849 8313 8861 8316
rect 8895 8313 8907 8347
rect 8849 8307 8907 8313
rect 9398 8304 9404 8356
rect 9456 8304 9462 8356
rect 9508 8316 9904 8344
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5442 8276 5448 8288
rect 4948 8248 5448 8276
rect 4948 8236 4954 8248
rect 5442 8236 5448 8248
rect 5500 8276 5506 8288
rect 5626 8276 5632 8288
rect 5500 8248 5632 8276
rect 5500 8236 5506 8248
rect 5626 8236 5632 8248
rect 5684 8276 5690 8288
rect 7742 8276 7748 8288
rect 5684 8248 7748 8276
rect 5684 8236 5690 8248
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 9508 8276 9536 8316
rect 8628 8248 9536 8276
rect 8628 8236 8634 8248
rect 9582 8236 9588 8288
rect 9640 8236 9646 8288
rect 9876 8276 9904 8316
rect 9950 8304 9956 8356
rect 10008 8344 10014 8356
rect 11900 8344 11928 8443
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 12584 8452 12633 8480
rect 12584 8440 12590 8452
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 13262 8480 13268 8492
rect 12851 8452 13268 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 12158 8372 12164 8424
rect 12216 8372 12222 8424
rect 10008 8316 11928 8344
rect 14292 8344 14320 8443
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 14752 8489 14780 8588
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15243 8588 15792 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15654 8548 15660 8560
rect 15488 8520 15660 8548
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 14476 8412 14504 8443
rect 14550 8412 14556 8424
rect 14476 8384 14556 8412
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 15028 8412 15056 8443
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 15488 8489 15516 8520
rect 15654 8508 15660 8520
rect 15712 8508 15718 8560
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15562 8440 15568 8492
rect 15620 8440 15626 8492
rect 14976 8384 15056 8412
rect 15657 8415 15715 8421
rect 14976 8372 14982 8384
rect 15657 8381 15669 8415
rect 15703 8381 15715 8415
rect 15764 8412 15792 8588
rect 15838 8576 15844 8628
rect 15896 8576 15902 8628
rect 16022 8576 16028 8628
rect 16080 8576 16086 8628
rect 17218 8616 17224 8628
rect 16684 8588 17224 8616
rect 15856 8548 15884 8576
rect 16393 8551 16451 8557
rect 16393 8548 16405 8551
rect 15856 8520 16405 8548
rect 16393 8517 16405 8520
rect 16439 8517 16451 8551
rect 16393 8511 16451 8517
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8449 16359 8483
rect 16301 8443 16359 8449
rect 16316 8412 16344 8443
rect 16482 8440 16488 8492
rect 16540 8440 16546 8492
rect 16684 8489 16712 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8616 17371 8619
rect 18417 8619 18475 8625
rect 18417 8616 18429 8619
rect 17359 8588 18429 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 18417 8585 18429 8588
rect 18463 8616 18475 8619
rect 18690 8616 18696 8628
rect 18463 8588 18696 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 19153 8619 19211 8625
rect 19153 8585 19165 8619
rect 19199 8616 19211 8619
rect 19199 8588 20300 8616
rect 19199 8585 19211 8588
rect 19153 8579 19211 8585
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 16908 8520 17540 8548
rect 16908 8508 16914 8520
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16942 8440 16948 8492
rect 17000 8440 17006 8492
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 16574 8412 16580 8424
rect 15764 8384 16580 8412
rect 15657 8375 15715 8381
rect 15286 8344 15292 8356
rect 14292 8316 15292 8344
rect 10008 8304 10014 8316
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 11882 8276 11888 8288
rect 9876 8248 11888 8276
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 11974 8236 11980 8288
rect 12032 8236 12038 8288
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 13354 8276 13360 8288
rect 12759 8248 13360 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 15672 8276 15700 8375
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 17236 8412 17264 8443
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 17512 8489 17540 8520
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 17773 8551 17831 8557
rect 17773 8548 17785 8551
rect 17644 8520 17785 8548
rect 17644 8508 17650 8520
rect 17773 8517 17785 8520
rect 17819 8517 17831 8551
rect 17954 8548 17960 8560
rect 17773 8511 17831 8517
rect 17880 8520 17960 8548
rect 17405 8483 17463 8489
rect 17405 8480 17417 8483
rect 17368 8452 17417 8480
rect 17368 8440 17374 8452
rect 17405 8449 17417 8452
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 17880 8489 17908 8520
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 18322 8557 18328 8560
rect 18307 8551 18328 8557
rect 18307 8517 18319 8551
rect 18307 8511 18328 8517
rect 18322 8508 18328 8511
rect 18380 8508 18386 8560
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18598 8480 18604 8492
rect 18555 8452 18604 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18156 8412 18184 8443
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 18708 8480 18736 8576
rect 18966 8508 18972 8560
rect 19024 8548 19030 8560
rect 19024 8520 19656 8548
rect 19024 8508 19030 8520
rect 19628 8489 19656 8520
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 18708 8452 19165 8480
rect 19153 8449 19165 8452
rect 19199 8449 19211 8483
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19153 8443 19211 8449
rect 19260 8452 19533 8480
rect 18693 8415 18751 8421
rect 17236 8384 17447 8412
rect 18156 8384 18552 8412
rect 17419 8356 17447 8384
rect 18524 8356 18552 8384
rect 18693 8381 18705 8415
rect 18739 8412 18751 8415
rect 18785 8415 18843 8421
rect 18785 8412 18797 8415
rect 18739 8384 18797 8412
rect 18739 8381 18751 8384
rect 18693 8375 18751 8381
rect 18785 8381 18797 8384
rect 18831 8381 18843 8415
rect 19260 8412 19288 8452
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 19702 8480 19708 8492
rect 19659 8452 19708 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 19935 8483 19993 8489
rect 19935 8449 19947 8483
rect 19981 8480 19993 8483
rect 20162 8480 20168 8492
rect 19981 8452 20168 8480
rect 19981 8449 19993 8452
rect 19935 8443 19993 8449
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 18785 8375 18843 8381
rect 18892 8384 19288 8412
rect 19337 8415 19395 8421
rect 16850 8304 16856 8356
rect 16908 8304 16914 8356
rect 17402 8304 17408 8356
rect 17460 8304 17466 8356
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 18138 8344 18144 8356
rect 17644 8316 18144 8344
rect 17644 8304 17650 8316
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 18506 8304 18512 8356
rect 18564 8304 18570 8356
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 18892 8344 18920 8384
rect 19337 8381 19349 8415
rect 19383 8381 19395 8415
rect 19337 8375 19395 8381
rect 18656 8316 18920 8344
rect 19352 8344 19380 8375
rect 19794 8372 19800 8424
rect 19852 8412 19858 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19852 8384 20085 8412
rect 19852 8372 19858 8384
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20272 8412 20300 8588
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 21140 8588 21189 8616
rect 21140 8576 21146 8588
rect 21177 8585 21189 8588
rect 21223 8585 21235 8619
rect 21177 8579 21235 8585
rect 21358 8576 21364 8628
rect 21416 8576 21422 8628
rect 23017 8619 23075 8625
rect 21468 8588 22876 8616
rect 20441 8551 20499 8557
rect 20441 8517 20453 8551
rect 20487 8548 20499 8551
rect 20809 8551 20867 8557
rect 20809 8548 20821 8551
rect 20487 8520 20821 8548
rect 20487 8517 20499 8520
rect 20441 8511 20499 8517
rect 20809 8517 20821 8520
rect 20855 8517 20867 8551
rect 20809 8511 20867 8517
rect 20898 8508 20904 8560
rect 20956 8508 20962 8560
rect 21266 8508 21272 8560
rect 21324 8548 21330 8560
rect 21468 8548 21496 8588
rect 21324 8520 21496 8548
rect 21324 8508 21330 8520
rect 21634 8508 21640 8560
rect 21692 8548 21698 8560
rect 22848 8548 22876 8588
rect 23017 8585 23029 8619
rect 23063 8616 23075 8619
rect 23198 8616 23204 8628
rect 23063 8588 23204 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 21692 8520 22508 8548
rect 22848 8520 22968 8548
rect 21692 8508 21698 8520
rect 20346 8440 20352 8492
rect 20404 8480 20410 8492
rect 20533 8483 20591 8489
rect 20533 8480 20545 8483
rect 20404 8452 20545 8480
rect 20404 8440 20410 8452
rect 20533 8449 20545 8452
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 20626 8483 20684 8489
rect 20626 8449 20638 8483
rect 20672 8449 20684 8483
rect 20626 8443 20684 8449
rect 20641 8412 20669 8443
rect 20990 8440 20996 8492
rect 21048 8489 21054 8492
rect 21048 8480 21056 8489
rect 21048 8452 21093 8480
rect 21048 8443 21056 8452
rect 21048 8440 21054 8443
rect 21542 8440 21548 8492
rect 21600 8440 21606 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21784 8452 21833 8480
rect 21784 8440 21790 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21968 8452 22017 8480
rect 21968 8440 21974 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 22480 8489 22508 8520
rect 22465 8483 22523 8489
rect 22465 8449 22477 8483
rect 22511 8449 22523 8483
rect 22465 8443 22523 8449
rect 22741 8483 22799 8489
rect 22741 8449 22753 8483
rect 22787 8480 22799 8483
rect 22830 8480 22836 8492
rect 22787 8452 22836 8480
rect 22787 8449 22799 8452
rect 22741 8443 22799 8449
rect 22830 8440 22836 8452
rect 22888 8440 22894 8492
rect 22940 8489 22968 8520
rect 22925 8483 22983 8489
rect 22925 8449 22937 8483
rect 22971 8449 22983 8483
rect 22925 8443 22983 8449
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8480 23259 8483
rect 24210 8480 24216 8492
rect 23247 8452 24216 8480
rect 23247 8449 23259 8452
rect 23201 8443 23259 8449
rect 24210 8440 24216 8452
rect 24268 8440 24274 8492
rect 20272 8384 20669 8412
rect 20073 8375 20131 8381
rect 22097 8347 22155 8353
rect 22097 8344 22109 8347
rect 19352 8316 22109 8344
rect 18656 8304 18662 8316
rect 22097 8313 22109 8316
rect 22143 8313 22155 8347
rect 22097 8307 22155 8313
rect 13872 8248 15700 8276
rect 13872 8236 13878 8248
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 16942 8276 16948 8288
rect 16724 8248 16948 8276
rect 16724 8236 16730 8248
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 17037 8279 17095 8285
rect 17037 8245 17049 8279
rect 17083 8276 17095 8279
rect 17954 8276 17960 8288
rect 17083 8248 17960 8276
rect 17083 8245 17095 8248
rect 17037 8239 17095 8245
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 18049 8279 18107 8285
rect 18049 8245 18061 8279
rect 18095 8276 18107 8279
rect 18230 8276 18236 8288
rect 18095 8248 18236 8276
rect 18095 8245 18107 8248
rect 18049 8239 18107 8245
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 1104 8186 23644 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 23644 8186
rect 1104 8112 23644 8134
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3786 8072 3792 8084
rect 3559 8044 3792 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 4614 8072 4620 8084
rect 4387 8044 4620 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5408 8044 5457 8072
rect 5408 8032 5414 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6089 8075 6147 8081
rect 6089 8072 6101 8075
rect 5868 8044 6101 8072
rect 5868 8032 5874 8044
rect 6089 8041 6101 8044
rect 6135 8041 6147 8075
rect 6089 8035 6147 8041
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 7190 8072 7196 8084
rect 6880 8044 7196 8072
rect 6880 8032 6886 8044
rect 7190 8032 7196 8044
rect 7248 8072 7254 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7248 8044 7757 8072
rect 7248 8032 7254 8044
rect 7745 8041 7757 8044
rect 7791 8072 7803 8075
rect 8941 8075 8999 8081
rect 7791 8044 8524 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 3326 7964 3332 8016
rect 3384 8004 3390 8016
rect 3421 8007 3479 8013
rect 3421 8004 3433 8007
rect 3384 7976 3433 8004
rect 3384 7964 3390 7976
rect 3421 7973 3433 7976
rect 3467 8004 3479 8007
rect 4249 8007 4307 8013
rect 4249 8004 4261 8007
rect 3467 7976 4261 8004
rect 3467 7973 3479 7976
rect 3421 7967 3479 7973
rect 4249 7973 4261 7976
rect 4295 7973 4307 8007
rect 5626 8004 5632 8016
rect 4249 7967 4307 7973
rect 4356 7976 5632 8004
rect 3605 7939 3663 7945
rect 3605 7905 3617 7939
rect 3651 7936 3663 7939
rect 4356 7936 4384 7976
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 6365 8007 6423 8013
rect 6365 7973 6377 8007
rect 6411 8004 6423 8007
rect 6454 8004 6460 8016
rect 6411 7976 6460 8004
rect 6411 7973 6423 7976
rect 6365 7967 6423 7973
rect 6454 7964 6460 7976
rect 6512 8004 6518 8016
rect 6917 8007 6975 8013
rect 6917 8004 6929 8007
rect 6512 7976 6929 8004
rect 6512 7964 6518 7976
rect 6917 7973 6929 7976
rect 6963 7973 6975 8007
rect 6917 7967 6975 7973
rect 7837 8007 7895 8013
rect 7837 7973 7849 8007
rect 7883 7973 7895 8007
rect 7837 7967 7895 7973
rect 3651 7908 4384 7936
rect 3651 7905 3663 7908
rect 3605 7899 3663 7905
rect 4430 7896 4436 7948
rect 4488 7896 4494 7948
rect 5350 7896 5356 7948
rect 5408 7936 5414 7948
rect 5905 7939 5963 7945
rect 5905 7936 5917 7939
rect 5408 7908 5917 7936
rect 5408 7896 5414 7908
rect 5905 7905 5917 7908
rect 5951 7905 5963 7939
rect 5905 7899 5963 7905
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7936 6055 7939
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6043 7908 6561 7936
rect 6043 7905 6055 7908
rect 5997 7899 6055 7905
rect 6549 7905 6561 7908
rect 6595 7936 6607 7939
rect 7852 7936 7880 7967
rect 6595 7908 7880 7936
rect 7929 7939 7987 7945
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 7929 7905 7941 7939
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 382 7828 388 7880
rect 440 7868 446 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 440 7840 1409 7868
rect 440 7828 446 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 1946 7868 1952 7880
rect 1719 7840 1952 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3344 7800 3372 7831
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4172 7800 4200 7828
rect 3344 7772 4200 7800
rect 4540 7800 4568 7831
rect 4614 7828 4620 7880
rect 4672 7828 4678 7880
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 6086 7868 6092 7880
rect 5767 7840 6092 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 4706 7800 4712 7812
rect 4540 7772 4712 7800
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 5644 7800 5672 7831
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6178 7800 6184 7812
rect 5644 7772 6184 7800
rect 6178 7760 6184 7772
rect 6236 7800 6242 7812
rect 6288 7800 6316 7831
rect 6236 7772 6316 7800
rect 6472 7800 6500 7831
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7377 7871 7435 7877
rect 7055 7840 7328 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 6638 7800 6644 7812
rect 6472 7772 6644 7800
rect 6236 7760 6242 7772
rect 6638 7760 6644 7772
rect 6696 7800 6702 7812
rect 7193 7803 7251 7809
rect 7193 7800 7205 7803
rect 6696 7772 7205 7800
rect 6696 7760 6702 7772
rect 7193 7769 7205 7772
rect 7239 7769 7251 7803
rect 7193 7763 7251 7769
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3936 7704 3985 7732
rect 3936 7692 3942 7704
rect 3973 7701 3985 7704
rect 4019 7701 4031 7735
rect 7300 7732 7328 7840
rect 7377 7837 7389 7871
rect 7423 7837 7435 7871
rect 7377 7831 7435 7837
rect 7392 7800 7420 7831
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7616 7840 7665 7868
rect 7616 7828 7622 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7944 7868 7972 7899
rect 8018 7868 8024 7880
rect 7944 7840 8024 7868
rect 7653 7831 7711 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8496 7877 8524 8044
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9030 8072 9036 8084
rect 8987 8044 9036 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 10042 8072 10048 8084
rect 9548 8044 10048 8072
rect 9548 8032 9554 8044
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 12066 8032 12072 8084
rect 12124 8032 12130 8084
rect 13170 8072 13176 8084
rect 12636 8044 13176 8072
rect 8757 8007 8815 8013
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 8846 8004 8852 8016
rect 8803 7976 8852 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 10318 8004 10324 8016
rect 9140 7976 10324 8004
rect 9140 7936 9168 7976
rect 10318 7964 10324 7976
rect 10376 7964 10382 8016
rect 12526 7964 12532 8016
rect 12584 7964 12590 8016
rect 12636 8013 12664 8044
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 15194 8032 15200 8084
rect 15252 8032 15258 8084
rect 15378 8032 15384 8084
rect 15436 8032 15442 8084
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 12621 8007 12679 8013
rect 12621 7973 12633 8007
rect 12667 7973 12679 8007
rect 12621 7967 12679 7973
rect 13078 7964 13084 8016
rect 13136 8004 13142 8016
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 13136 7976 13277 8004
rect 13136 7964 13142 7976
rect 13265 7973 13277 7976
rect 13311 7973 13323 8007
rect 13265 7967 13323 7973
rect 14366 7964 14372 8016
rect 14424 8004 14430 8016
rect 15580 8004 15608 8035
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17586 8072 17592 8084
rect 17092 8044 17592 8072
rect 17092 8032 17098 8044
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 17696 8044 17908 8072
rect 16025 8007 16083 8013
rect 16025 8004 16037 8007
rect 14424 7976 16037 8004
rect 14424 7964 14430 7976
rect 16025 7973 16037 7976
rect 16071 7973 16083 8007
rect 16025 7967 16083 7973
rect 8772 7908 9168 7936
rect 8481 7871 8539 7877
rect 8128 7840 8432 7868
rect 7466 7800 7472 7812
rect 7392 7772 7472 7800
rect 7466 7760 7472 7772
rect 7524 7800 7530 7812
rect 8128 7800 8156 7840
rect 8404 7812 8432 7840
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 8772 7877 8800 7908
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9272 7908 9597 7936
rect 9272 7896 9278 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 10594 7936 10600 7948
rect 9585 7899 9643 7905
rect 10244 7908 10600 7936
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 9858 7877 9864 7880
rect 9447 7871 9505 7877
rect 9447 7837 9459 7871
rect 9493 7868 9505 7871
rect 9856 7868 9864 7877
rect 9493 7840 9720 7868
rect 9819 7840 9864 7868
rect 9493 7837 9505 7840
rect 9447 7831 9505 7837
rect 7524 7772 8156 7800
rect 7524 7760 7530 7772
rect 8202 7760 8208 7812
rect 8260 7760 8266 7812
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 9217 7803 9275 7809
rect 9217 7800 9229 7803
rect 8996 7772 9229 7800
rect 8996 7760 9002 7772
rect 9217 7769 9229 7772
rect 9263 7769 9275 7803
rect 9217 7763 9275 7769
rect 9310 7803 9368 7809
rect 9310 7769 9322 7803
rect 9356 7769 9368 7803
rect 9310 7763 9368 7769
rect 8220 7732 8248 7760
rect 7300 7704 8248 7732
rect 9324 7732 9352 7763
rect 9582 7732 9588 7744
rect 9324 7704 9588 7732
rect 3973 7695 4031 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 9692 7741 9720 7840
rect 9856 7831 9864 7840
rect 9858 7828 9864 7831
rect 9916 7828 9922 7880
rect 10244 7877 10272 7908
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 12161 7939 12219 7945
rect 12161 7936 12173 7939
rect 11756 7908 12173 7936
rect 11756 7896 11762 7908
rect 12161 7905 12173 7908
rect 12207 7905 12219 7939
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 12161 7899 12219 7905
rect 12728 7908 13645 7936
rect 10318 7877 10324 7880
rect 10228 7871 10286 7877
rect 10228 7837 10240 7871
rect 10274 7837 10286 7871
rect 10228 7831 10286 7837
rect 10314 7831 10324 7877
rect 10376 7868 10382 7880
rect 10376 7840 10414 7868
rect 10318 7828 10324 7831
rect 10376 7828 10382 7840
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12618 7868 12624 7880
rect 12483 7840 12624 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 12728 7877 12756 7908
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7936 14795 7939
rect 15286 7936 15292 7948
rect 14783 7908 15292 7936
rect 14783 7905 14795 7908
rect 14737 7899 14795 7905
rect 15286 7896 15292 7908
rect 15344 7936 15350 7948
rect 15562 7936 15568 7948
rect 15344 7908 15568 7936
rect 15344 7896 15350 7908
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 17402 7936 17408 7948
rect 15712 7908 17408 7936
rect 15712 7896 15718 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 17696 7936 17724 8044
rect 17880 8004 17908 8044
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18598 8072 18604 8084
rect 18012 8044 18604 8072
rect 18012 8032 18018 8044
rect 18598 8032 18604 8044
rect 18656 8072 18662 8084
rect 18782 8072 18788 8084
rect 18656 8044 18788 8072
rect 18656 8032 18662 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 18969 8075 19027 8081
rect 18969 8041 18981 8075
rect 19015 8072 19027 8075
rect 19058 8072 19064 8084
rect 19015 8044 19064 8072
rect 19015 8041 19027 8044
rect 18969 8035 19027 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19150 8032 19156 8084
rect 19208 8072 19214 8084
rect 22278 8072 22284 8084
rect 19208 8044 22284 8072
rect 19208 8032 19214 8044
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 23014 8032 23020 8084
rect 23072 8032 23078 8084
rect 19242 8004 19248 8016
rect 17880 7976 19248 8004
rect 19242 7964 19248 7976
rect 19300 8004 19306 8016
rect 19518 8004 19524 8016
rect 19300 7976 19524 8004
rect 19300 7964 19306 7976
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 20622 7964 20628 8016
rect 20680 8004 20686 8016
rect 20680 7976 23244 8004
rect 20680 7964 20686 7976
rect 18417 7939 18475 7945
rect 17604 7908 17724 7936
rect 17880 7908 18184 7936
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12860 7840 13093 7868
rect 12860 7828 12866 7840
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 9950 7760 9956 7812
rect 10008 7760 10014 7812
rect 10042 7760 10048 7812
rect 10100 7760 10106 7812
rect 11992 7800 12020 7828
rect 11900 7772 12020 7800
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7701 9735 7735
rect 9968 7732 9996 7760
rect 11900 7732 11928 7772
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13188 7800 13216 7831
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 13538 7828 13544 7880
rect 13596 7828 13602 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13771 7840 14105 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 13740 7800 13768 7831
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 14642 7877 14648 7880
rect 14599 7871 14648 7877
rect 14599 7837 14611 7871
rect 14645 7837 14648 7871
rect 14599 7831 14648 7837
rect 14642 7828 14648 7831
rect 14700 7828 14706 7880
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15059 7840 15093 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 12584 7772 13768 7800
rect 12584 7760 12590 7772
rect 14366 7760 14372 7812
rect 14424 7760 14430 7812
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7800 14979 7803
rect 15028 7800 15056 7831
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 15528 7840 16221 7868
rect 15528 7828 15534 7840
rect 16209 7837 16221 7840
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 16301 7871 16359 7877
rect 16301 7837 16313 7871
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 14967 7772 15884 7800
rect 14967 7769 14979 7772
rect 14921 7763 14979 7769
rect 9968 7704 11928 7732
rect 9677 7695 9735 7701
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 12124 7704 12265 7732
rect 12124 7692 12130 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12860 7704 12909 7732
rect 12860 7692 12866 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 12897 7695 12955 7701
rect 15556 7735 15614 7741
rect 15556 7701 15568 7735
rect 15602 7732 15614 7735
rect 15746 7732 15752 7744
rect 15602 7704 15752 7732
rect 15602 7701 15614 7704
rect 15556 7695 15614 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 15856 7732 15884 7772
rect 15930 7760 15936 7812
rect 15988 7760 15994 7812
rect 16114 7760 16120 7812
rect 16172 7800 16178 7812
rect 16316 7800 16344 7831
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16669 7871 16727 7877
rect 16669 7868 16681 7871
rect 16632 7840 16681 7868
rect 16632 7828 16638 7840
rect 16669 7837 16681 7840
rect 16715 7868 16727 7871
rect 16850 7868 16856 7880
rect 16715 7840 16856 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 16942 7828 16948 7880
rect 17000 7828 17006 7880
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17494 7868 17500 7880
rect 17276 7840 17500 7868
rect 17276 7828 17282 7840
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 17604 7877 17632 7908
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 17758 7828 17764 7880
rect 17816 7877 17822 7880
rect 17816 7871 17831 7877
rect 17819 7837 17831 7871
rect 17816 7831 17831 7837
rect 17816 7828 17822 7831
rect 16172 7772 16344 7800
rect 16172 7760 16178 7772
rect 17310 7760 17316 7812
rect 17368 7800 17374 7812
rect 17880 7800 17908 7908
rect 17954 7828 17960 7880
rect 18012 7828 18018 7880
rect 18156 7877 18184 7908
rect 18417 7905 18429 7939
rect 18463 7936 18475 7939
rect 19058 7936 19064 7948
rect 18463 7908 19064 7936
rect 18463 7905 18475 7908
rect 18417 7899 18475 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 20714 7936 20720 7948
rect 19306 7908 20720 7936
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18506 7868 18512 7880
rect 18187 7840 18512 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 18690 7828 18696 7880
rect 18748 7828 18754 7880
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 19306 7868 19334 7908
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 18976 7840 19334 7868
rect 17368 7772 17908 7800
rect 18049 7803 18107 7809
rect 17368 7760 17374 7772
rect 18049 7769 18061 7803
rect 18095 7769 18107 7803
rect 18049 7763 18107 7769
rect 18601 7803 18659 7809
rect 18601 7769 18613 7803
rect 18647 7800 18659 7803
rect 18976 7800 19004 7840
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 23216 7877 23244 7976
rect 21085 7871 21143 7877
rect 21085 7868 21097 7871
rect 20588 7840 21097 7868
rect 20588 7828 20594 7840
rect 21085 7837 21097 7840
rect 21131 7837 21143 7871
rect 21085 7831 21143 7837
rect 23201 7871 23259 7877
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 18647 7772 19004 7800
rect 18647 7769 18659 7772
rect 18601 7763 18659 7769
rect 16298 7732 16304 7744
rect 15856 7704 16304 7732
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16853 7735 16911 7741
rect 16853 7701 16865 7735
rect 16899 7732 16911 7735
rect 17126 7732 17132 7744
rect 16899 7704 17132 7732
rect 16899 7701 16911 7704
rect 16853 7695 16911 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 18064 7732 18092 7763
rect 19334 7760 19340 7812
rect 19392 7760 19398 7812
rect 20990 7760 20996 7812
rect 21048 7760 21054 7812
rect 18138 7732 18144 7744
rect 18064 7704 18144 7732
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18506 7732 18512 7744
rect 18371 7704 18512 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 22373 7735 22431 7741
rect 22373 7732 22385 7735
rect 21140 7704 22385 7732
rect 21140 7692 21146 7704
rect 22373 7701 22385 7704
rect 22419 7732 22431 7735
rect 22646 7732 22652 7744
rect 22419 7704 22652 7732
rect 22419 7701 22431 7704
rect 22373 7695 22431 7701
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 1104 7642 23644 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 23644 7642
rect 1104 7568 23644 7590
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 4798 7528 4804 7540
rect 4387 7500 4804 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5184 7500 5549 7528
rect 3973 7463 4031 7469
rect 3973 7429 3985 7463
rect 4019 7460 4031 7463
rect 4062 7460 4068 7472
rect 4019 7432 4068 7460
rect 4019 7429 4031 7432
rect 3973 7423 4031 7429
rect 4062 7420 4068 7432
rect 4120 7420 4126 7472
rect 4614 7460 4620 7472
rect 4264 7432 4620 7460
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 4264 7401 4292 7432
rect 4614 7420 4620 7432
rect 4672 7460 4678 7472
rect 5184 7469 5212 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 6178 7488 6184 7540
rect 6236 7488 6242 7540
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6788 7500 6837 7528
rect 6788 7488 6794 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9214 7528 9220 7540
rect 9079 7500 9220 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 9858 7488 9864 7540
rect 9916 7528 9922 7540
rect 14366 7528 14372 7540
rect 9916 7500 14372 7528
rect 9916 7488 9922 7500
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 15194 7528 15200 7540
rect 14967 7500 15200 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 15194 7488 15200 7500
rect 15252 7488 15258 7540
rect 15562 7488 15568 7540
rect 15620 7488 15626 7540
rect 17402 7488 17408 7540
rect 17460 7488 17466 7540
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 18046 7528 18052 7540
rect 17635 7500 18052 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 18046 7488 18052 7500
rect 18104 7528 18110 7540
rect 19702 7528 19708 7540
rect 18104 7500 19708 7528
rect 18104 7488 18110 7500
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 20772 7500 21404 7528
rect 20772 7488 20778 7500
rect 5169 7463 5227 7469
rect 5169 7460 5181 7463
rect 4672 7432 5181 7460
rect 4672 7420 4678 7432
rect 5169 7429 5181 7432
rect 5215 7429 5227 7463
rect 5169 7423 5227 7429
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 5353 7463 5411 7469
rect 5353 7460 5365 7463
rect 5316 7432 5365 7460
rect 5316 7420 5322 7432
rect 5353 7429 5365 7432
rect 5399 7460 5411 7463
rect 5399 7432 5764 7460
rect 5399 7429 5411 7432
rect 5353 7423 5411 7429
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 3651 7364 4261 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 5736 7401 5764 7432
rect 6270 7420 6276 7472
rect 6328 7460 6334 7472
rect 6365 7463 6423 7469
rect 6365 7460 6377 7463
rect 6328 7432 6377 7460
rect 6328 7420 6334 7432
rect 6365 7429 6377 7432
rect 6411 7429 6423 7463
rect 9232 7460 9260 7488
rect 12158 7460 12164 7472
rect 9232 7432 12164 7460
rect 6365 7423 6423 7429
rect 12158 7420 12164 7432
rect 12216 7460 12222 7472
rect 12216 7432 12940 7460
rect 12216 7420 12222 7432
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4396 7364 4445 7392
rect 4396 7352 4402 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 5092 7324 5120 7355
rect 5460 7324 5488 7355
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6512 7364 6561 7392
rect 6512 7352 6518 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 3936 7296 5488 7324
rect 3936 7284 3942 7296
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6932 7324 6960 7355
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 9398 7352 9404 7404
rect 9456 7352 9462 7404
rect 9769 7395 9827 7401
rect 9769 7392 9781 7395
rect 9600 7364 9781 7392
rect 6144 7296 6960 7324
rect 6144 7284 6150 7296
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8202 7324 8208 7336
rect 7984 7296 8208 7324
rect 7984 7284 7990 7296
rect 8202 7284 8208 7296
rect 8260 7324 8266 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8260 7296 8585 7324
rect 8260 7284 8266 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 9600 7324 9628 7364
rect 9769 7361 9781 7364
rect 9815 7361 9827 7395
rect 9769 7355 9827 7361
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 11698 7392 11704 7404
rect 10376 7364 11704 7392
rect 10376 7352 10382 7364
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12437 7395 12495 7401
rect 12437 7392 12449 7395
rect 12084 7364 12449 7392
rect 9180 7296 9628 7324
rect 9180 7284 9186 7296
rect 9674 7284 9680 7336
rect 9732 7284 9738 7336
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 12084 7324 12112 7364
rect 12437 7361 12449 7364
rect 12483 7392 12495 7395
rect 12526 7392 12532 7404
rect 12483 7364 12532 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 12912 7392 12940 7432
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 13081 7463 13139 7469
rect 13081 7460 13093 7463
rect 13044 7432 13093 7460
rect 13044 7420 13050 7432
rect 13081 7429 13093 7432
rect 13127 7429 13139 7463
rect 13081 7423 13139 7429
rect 14829 7463 14887 7469
rect 14829 7429 14841 7463
rect 14875 7460 14887 7463
rect 15654 7460 15660 7472
rect 14875 7432 15660 7460
rect 14875 7429 14887 7432
rect 14829 7423 14887 7429
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 15933 7463 15991 7469
rect 15933 7429 15945 7463
rect 15979 7460 15991 7463
rect 17218 7460 17224 7472
rect 15979 7432 17224 7460
rect 15979 7429 15991 7432
rect 15933 7423 15991 7429
rect 14734 7392 14740 7404
rect 12912 7364 14740 7392
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 10560 7296 12112 7324
rect 10560 7284 10566 7296
rect 12158 7284 12164 7336
rect 12216 7324 12222 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12216 7296 12725 7324
rect 12216 7284 12222 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12894 7284 12900 7336
rect 12952 7284 12958 7336
rect 14752 7324 14780 7352
rect 15212 7324 15240 7355
rect 15286 7352 15292 7404
rect 15344 7352 15350 7404
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7392 15531 7395
rect 15562 7392 15568 7404
rect 15519 7364 15568 7392
rect 15519 7361 15531 7364
rect 15473 7355 15531 7361
rect 15562 7352 15568 7364
rect 15620 7392 15626 7404
rect 15749 7395 15807 7401
rect 15749 7392 15761 7395
rect 15620 7364 15761 7392
rect 15620 7352 15626 7364
rect 15749 7361 15761 7364
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 15378 7324 15384 7336
rect 14752 7296 15384 7324
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 4157 7259 4215 7265
rect 4157 7225 4169 7259
rect 4203 7256 4215 7259
rect 5258 7256 5264 7268
rect 4203 7228 5264 7256
rect 4203 7225 4215 7228
rect 4157 7219 4215 7225
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 5350 7216 5356 7268
rect 5408 7216 5414 7268
rect 5810 7216 5816 7268
rect 5868 7256 5874 7268
rect 6730 7256 6736 7268
rect 5868 7228 6736 7256
rect 5868 7216 5874 7228
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 8386 7216 8392 7268
rect 8444 7256 8450 7268
rect 8846 7256 8852 7268
rect 8444 7228 8852 7256
rect 8444 7216 8450 7228
rect 8846 7216 8852 7228
rect 8904 7216 8910 7268
rect 12529 7259 12587 7265
rect 12529 7256 12541 7259
rect 8956 7228 12541 7256
rect 198 7148 204 7200
rect 256 7188 262 7200
rect 1489 7191 1547 7197
rect 1489 7188 1501 7191
rect 256 7160 1501 7188
rect 256 7148 262 7160
rect 1489 7157 1501 7160
rect 1535 7157 1547 7191
rect 1489 7151 1547 7157
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 4338 7188 4344 7200
rect 4028 7160 4344 7188
rect 4028 7148 4034 7160
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 4798 7188 4804 7200
rect 4488 7160 4804 7188
rect 4488 7148 4494 7160
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 6086 7188 6092 7200
rect 5951 7160 6092 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7188 6423 7191
rect 8956 7188 8984 7228
rect 12529 7225 12541 7228
rect 12575 7225 12587 7259
rect 12529 7219 12587 7225
rect 14090 7216 14096 7268
rect 14148 7256 14154 7268
rect 14148 7228 15056 7256
rect 14148 7216 14154 7228
rect 6411 7160 8984 7188
rect 6411 7157 6423 7160
rect 6365 7151 6423 7157
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 9088 7160 9137 7188
rect 9088 7148 9094 7160
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 15028 7188 15056 7228
rect 15102 7216 15108 7268
rect 15160 7256 15166 7268
rect 15948 7256 15976 7423
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 17420 7460 17448 7488
rect 17681 7463 17739 7469
rect 17681 7460 17693 7463
rect 17420 7432 17693 7460
rect 17681 7429 17693 7432
rect 17727 7429 17739 7463
rect 17681 7423 17739 7429
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 18288 7432 20668 7460
rect 18288 7420 18294 7432
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 16574 7392 16580 7404
rect 16531 7364 16580 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 16224 7324 16252 7355
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16758 7324 16764 7336
rect 16224 7296 16764 7324
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 16868 7324 16896 7355
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 17310 7352 17316 7404
rect 17368 7352 17374 7404
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17494 7352 17500 7404
rect 17552 7392 17558 7404
rect 19702 7401 19708 7404
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 17552 7364 19533 7392
rect 17552 7352 17558 7364
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19699 7355 19708 7401
rect 19702 7352 19708 7355
rect 19760 7352 19766 7404
rect 20640 7401 20668 7432
rect 21082 7420 21088 7472
rect 21140 7460 21146 7472
rect 21269 7463 21327 7469
rect 21269 7460 21281 7463
rect 21140 7432 21281 7460
rect 21140 7420 21146 7432
rect 21269 7429 21281 7432
rect 21315 7429 21327 7463
rect 21376 7460 21404 7500
rect 21542 7488 21548 7540
rect 21600 7528 21606 7540
rect 21913 7531 21971 7537
rect 21913 7528 21925 7531
rect 21600 7500 21925 7528
rect 21600 7488 21606 7500
rect 21913 7497 21925 7500
rect 21959 7497 21971 7531
rect 21913 7491 21971 7497
rect 22189 7463 22247 7469
rect 22189 7460 22201 7463
rect 21376 7432 22201 7460
rect 21269 7423 21327 7429
rect 22189 7429 22201 7432
rect 22235 7429 22247 7463
rect 22189 7423 22247 7429
rect 22278 7420 22284 7472
rect 22336 7420 22342 7472
rect 22830 7420 22836 7472
rect 22888 7460 22894 7472
rect 22888 7432 23060 7460
rect 22888 7420 22894 7432
rect 20625 7395 20683 7401
rect 20625 7361 20637 7395
rect 20671 7361 20683 7395
rect 20625 7355 20683 7361
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20772 7364 20821 7392
rect 20772 7352 20778 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 21450 7392 21456 7404
rect 20956 7364 21456 7392
rect 20956 7352 20962 7364
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 19613 7327 19671 7333
rect 16868 7296 17540 7324
rect 15160 7228 15976 7256
rect 15160 7216 15166 7228
rect 16482 7216 16488 7268
rect 16540 7256 16546 7268
rect 17310 7256 17316 7268
rect 16540 7228 17316 7256
rect 16540 7216 16546 7228
rect 17310 7216 17316 7228
rect 17368 7216 17374 7268
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15028 7160 16037 7188
rect 9125 7151 9183 7157
rect 16025 7157 16037 7160
rect 16071 7188 16083 7191
rect 16206 7188 16212 7200
rect 16071 7160 16212 7188
rect 16071 7157 16083 7160
rect 16025 7151 16083 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16390 7148 16396 7200
rect 16448 7148 16454 7200
rect 17034 7148 17040 7200
rect 17092 7188 17098 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 17092 7160 17141 7188
rect 17092 7148 17098 7160
rect 17129 7157 17141 7160
rect 17175 7157 17187 7191
rect 17512 7188 17540 7296
rect 19613 7293 19625 7327
rect 19659 7324 19671 7327
rect 22572 7324 22600 7355
rect 22646 7352 22652 7404
rect 22704 7392 22710 7404
rect 22741 7395 22799 7401
rect 22741 7392 22753 7395
rect 22704 7364 22753 7392
rect 22704 7352 22710 7364
rect 22741 7361 22753 7364
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 22922 7352 22928 7404
rect 22980 7352 22986 7404
rect 23032 7401 23060 7432
rect 23017 7395 23075 7401
rect 23017 7361 23029 7395
rect 23063 7361 23075 7395
rect 23017 7355 23075 7361
rect 23201 7327 23259 7333
rect 23201 7324 23213 7327
rect 19659 7296 22324 7324
rect 22572 7296 23213 7324
rect 19659 7293 19671 7296
rect 19613 7287 19671 7293
rect 18598 7216 18604 7268
rect 18656 7256 18662 7268
rect 21450 7256 21456 7268
rect 18656 7228 21456 7256
rect 18656 7216 18662 7228
rect 21450 7216 21456 7228
rect 21508 7216 21514 7268
rect 18230 7188 18236 7200
rect 17512 7160 18236 7188
rect 17129 7151 17187 7157
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 19153 7191 19211 7197
rect 19153 7157 19165 7191
rect 19199 7188 19211 7191
rect 19242 7188 19248 7200
rect 19199 7160 19248 7188
rect 19199 7157 19211 7160
rect 19153 7151 19211 7157
rect 19242 7148 19248 7160
rect 19300 7188 19306 7200
rect 20438 7188 20444 7200
rect 19300 7160 20444 7188
rect 19300 7148 19306 7160
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20714 7148 20720 7200
rect 20772 7148 20778 7200
rect 21085 7191 21143 7197
rect 21085 7157 21097 7191
rect 21131 7188 21143 7191
rect 21174 7188 21180 7200
rect 21131 7160 21180 7188
rect 21131 7157 21143 7160
rect 21085 7151 21143 7157
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 22296 7188 22324 7296
rect 23201 7293 23213 7296
rect 23247 7293 23259 7327
rect 23201 7287 23259 7293
rect 22833 7259 22891 7265
rect 22833 7225 22845 7259
rect 22879 7256 22891 7259
rect 23290 7256 23296 7268
rect 22879 7228 23296 7256
rect 22879 7225 22891 7228
rect 22833 7219 22891 7225
rect 23290 7216 23296 7228
rect 23348 7216 23354 7268
rect 22370 7188 22376 7200
rect 22296 7160 22376 7188
rect 22370 7148 22376 7160
rect 22428 7148 22434 7200
rect 1104 7098 23644 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 23644 7098
rect 1104 7024 23644 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2004 6956 2912 6984
rect 2004 6944 2010 6956
rect 2884 6925 2912 6956
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 5718 6984 5724 6996
rect 4304 6956 5724 6984
rect 4304 6944 4310 6956
rect 5718 6944 5724 6956
rect 5776 6984 5782 6996
rect 7374 6984 7380 6996
rect 5776 6956 7380 6984
rect 5776 6944 5782 6956
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 9858 6984 9864 6996
rect 7800 6956 9864 6984
rect 7800 6944 7806 6956
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 10008 6956 10057 6984
rect 10008 6944 10014 6956
rect 10045 6953 10057 6956
rect 10091 6984 10103 6987
rect 10965 6987 11023 6993
rect 10965 6984 10977 6987
rect 10091 6956 10977 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 10965 6953 10977 6956
rect 11011 6953 11023 6987
rect 10965 6947 11023 6953
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13354 6984 13360 6996
rect 13035 6956 13360 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13464 6956 16252 6984
rect 2225 6919 2283 6925
rect 2225 6885 2237 6919
rect 2271 6885 2283 6919
rect 2225 6879 2283 6885
rect 2869 6919 2927 6925
rect 2869 6885 2881 6919
rect 2915 6916 2927 6919
rect 3326 6916 3332 6928
rect 2915 6888 3332 6916
rect 2915 6885 2927 6888
rect 2869 6879 2927 6885
rect 1946 6808 1952 6860
rect 2004 6808 2010 6860
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1636 6752 1685 6780
rect 1636 6740 1642 6752
rect 1673 6749 1685 6752
rect 1719 6780 1731 6783
rect 2240 6780 2268 6879
rect 3326 6876 3332 6888
rect 3384 6876 3390 6928
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 6086 6916 6092 6928
rect 5316 6888 6092 6916
rect 5316 6876 5322 6888
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 6454 6876 6460 6928
rect 6512 6876 6518 6928
rect 7926 6876 7932 6928
rect 7984 6916 7990 6928
rect 9217 6919 9275 6925
rect 9217 6916 9229 6919
rect 7984 6888 9229 6916
rect 7984 6876 7990 6888
rect 9217 6885 9229 6888
rect 9263 6885 9275 6919
rect 9217 6879 9275 6885
rect 9401 6919 9459 6925
rect 9401 6885 9413 6919
rect 9447 6916 9459 6919
rect 10318 6916 10324 6928
rect 9447 6888 10324 6916
rect 9447 6885 9459 6888
rect 9401 6879 9459 6885
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 13464 6916 13492 6956
rect 15102 6916 15108 6928
rect 10612 6888 13492 6916
rect 14936 6888 15108 6916
rect 4154 6848 4160 6860
rect 3160 6820 4160 6848
rect 3160 6789 3188 6820
rect 4154 6808 4160 6820
rect 4212 6848 4218 6860
rect 4274 6851 4332 6857
rect 4274 6848 4286 6851
rect 4212 6820 4286 6848
rect 4212 6808 4218 6820
rect 4274 6817 4286 6820
rect 4320 6817 4332 6851
rect 4274 6811 4332 6817
rect 5905 6851 5963 6857
rect 5905 6817 5917 6851
rect 5951 6848 5963 6851
rect 9953 6851 10011 6857
rect 5951 6820 9720 6848
rect 5951 6817 5963 6820
rect 5905 6811 5963 6817
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 1719 6752 2605 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2593 6749 2605 6752
rect 2639 6780 2651 6783
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 2639 6752 3157 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3384 6752 3801 6780
rect 3384 6740 3390 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 4706 6780 4712 6792
rect 3789 6743 3847 6749
rect 3896 6752 4712 6780
rect 3896 6712 3924 6752
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 2746 6684 3924 6712
rect 4065 6715 4123 6721
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 2130 6644 2136 6656
rect 1811 6616 2136 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2746 6644 2774 6684
rect 4065 6681 4077 6715
rect 4111 6712 4123 6715
rect 4522 6712 4528 6724
rect 4111 6684 4528 6712
rect 4111 6681 4123 6684
rect 4065 6675 4123 6681
rect 4522 6672 4528 6684
rect 4580 6672 4586 6724
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 5166 6712 5172 6724
rect 4672 6684 5172 6712
rect 4672 6672 4678 6684
rect 5166 6672 5172 6684
rect 5224 6712 5230 6724
rect 5460 6712 5488 6743
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6546 6780 6552 6792
rect 6503 6752 6552 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8018 6780 8024 6792
rect 7791 6752 8024 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8904 6752 8953 6780
rect 8904 6740 8910 6752
rect 8941 6749 8953 6752
rect 8987 6780 8999 6783
rect 9582 6780 9588 6792
rect 8987 6752 9588 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9692 6789 9720 6820
rect 9953 6817 9965 6851
rect 9999 6848 10011 6851
rect 10042 6848 10048 6860
rect 9999 6820 10048 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 10042 6808 10048 6820
rect 10100 6848 10106 6860
rect 10612 6848 10640 6888
rect 10100 6820 10640 6848
rect 10100 6808 10106 6820
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10744 6820 10793 6848
rect 10744 6808 10750 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 11606 6808 11612 6860
rect 11664 6808 11670 6860
rect 11716 6820 12112 6848
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 9858 6780 9864 6792
rect 9723 6752 9864 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 11238 6780 11244 6792
rect 11103 6752 11244 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 5224 6684 5488 6712
rect 6273 6715 6331 6721
rect 5224 6672 5230 6684
rect 6273 6681 6285 6715
rect 6319 6712 6331 6715
rect 6362 6712 6368 6724
rect 6319 6684 6368 6712
rect 6319 6681 6331 6684
rect 6273 6675 6331 6681
rect 6362 6672 6368 6684
rect 6420 6712 6426 6724
rect 6420 6684 7972 6712
rect 6420 6672 6426 6684
rect 2455 6616 2774 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 3050 6604 3056 6656
rect 3108 6604 3114 6656
rect 3510 6604 3516 6656
rect 3568 6604 3574 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4157 6647 4215 6653
rect 4157 6644 4169 6647
rect 4028 6616 4169 6644
rect 4028 6604 4034 6616
rect 4157 6613 4169 6616
rect 4203 6644 4215 6647
rect 4338 6644 4344 6656
rect 4203 6616 4344 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 4433 6647 4491 6653
rect 4433 6613 4445 6647
rect 4479 6644 4491 6647
rect 5810 6644 5816 6656
rect 4479 6616 5816 6644
rect 4479 6613 4491 6616
rect 4433 6607 4491 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 5994 6604 6000 6656
rect 6052 6644 6058 6656
rect 7834 6644 7840 6656
rect 6052 6616 7840 6644
rect 6052 6604 6058 6616
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 7944 6644 7972 6684
rect 9030 6672 9036 6724
rect 9088 6712 9094 6724
rect 10336 6712 10364 6743
rect 9088 6684 10364 6712
rect 9088 6672 9094 6684
rect 9766 6644 9772 6656
rect 7944 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10229 6647 10287 6653
rect 10229 6613 10241 6647
rect 10275 6644 10287 6647
rect 10318 6644 10324 6656
rect 10275 6616 10324 6644
rect 10275 6613 10287 6616
rect 10229 6607 10287 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10413 6647 10471 6653
rect 10413 6613 10425 6647
rect 10459 6644 10471 6647
rect 10502 6644 10508 6656
rect 10459 6616 10508 6644
rect 10459 6613 10471 6616
rect 10413 6607 10471 6613
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 10612 6644 10640 6743
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 10888 6712 10916 6743
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 11716 6780 11744 6820
rect 11572 6752 11744 6780
rect 11793 6783 11851 6789
rect 11572 6740 11578 6752
rect 11793 6749 11805 6783
rect 11839 6749 11851 6783
rect 11793 6743 11851 6749
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 11974 6780 11980 6792
rect 11931 6752 11980 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 11330 6712 11336 6724
rect 10744 6684 11336 6712
rect 10744 6672 10750 6684
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 11532 6644 11560 6740
rect 11808 6712 11836 6743
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 12084 6780 12112 6820
rect 12158 6808 12164 6860
rect 12216 6808 12222 6860
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 12308 6820 13216 6848
rect 12308 6808 12314 6820
rect 12342 6780 12348 6792
rect 12084 6752 12348 6780
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12492 6752 12541 6780
rect 12492 6740 12498 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 12714 6783 12772 6789
rect 12714 6749 12726 6783
rect 12760 6780 12772 6783
rect 12802 6780 12808 6792
rect 12760 6752 12808 6780
rect 12760 6749 12772 6752
rect 12714 6743 12772 6749
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 13188 6789 13216 6820
rect 14366 6808 14372 6860
rect 14424 6848 14430 6860
rect 14936 6848 14964 6888
rect 15102 6876 15108 6888
rect 15160 6876 15166 6928
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15838 6916 15844 6928
rect 15436 6888 15844 6916
rect 15436 6876 15442 6888
rect 15838 6876 15844 6888
rect 15896 6876 15902 6928
rect 16224 6916 16252 6956
rect 16298 6944 16304 6996
rect 16356 6984 16362 6996
rect 16356 6956 19334 6984
rect 16356 6944 16362 6956
rect 17678 6916 17684 6928
rect 16224 6888 17684 6916
rect 17678 6876 17684 6888
rect 17736 6916 17742 6928
rect 17954 6916 17960 6928
rect 17736 6888 17960 6916
rect 17736 6876 17742 6888
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 18046 6876 18052 6928
rect 18104 6916 18110 6928
rect 18104 6888 18368 6916
rect 18104 6876 18110 6888
rect 14424 6820 14964 6848
rect 14424 6808 14430 6820
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13630 6780 13636 6792
rect 13311 6752 13636 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 14148 6752 14289 6780
rect 14148 6740 14154 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 12636 6712 12664 6740
rect 11808 6684 12664 6712
rect 12989 6715 13047 6721
rect 12989 6681 13001 6715
rect 13035 6681 13047 6715
rect 12989 6675 13047 6681
rect 10612 6616 11560 6644
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6644 12127 6647
rect 12250 6644 12256 6656
rect 12115 6616 12256 6644
rect 12115 6613 12127 6616
rect 12069 6607 12127 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 13004 6644 13032 6675
rect 13446 6672 13452 6724
rect 13504 6712 13510 6724
rect 14476 6712 14504 6743
rect 14734 6740 14740 6792
rect 14792 6740 14798 6792
rect 14936 6789 14964 6820
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 15988 6820 17264 6848
rect 15988 6808 15994 6820
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6780 15163 6783
rect 15286 6780 15292 6792
rect 15151 6752 15292 6780
rect 15151 6749 15163 6752
rect 15105 6743 15163 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 17236 6789 17264 6820
rect 17402 6808 17408 6860
rect 17460 6848 17466 6860
rect 18138 6848 18144 6860
rect 17460 6820 18144 6848
rect 17460 6808 17466 6820
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 18230 6808 18236 6860
rect 18288 6808 18294 6860
rect 18340 6857 18368 6888
rect 18966 6876 18972 6928
rect 19024 6876 19030 6928
rect 19306 6916 19334 6956
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 22094 6984 22100 6996
rect 19576 6956 22100 6984
rect 19576 6944 19582 6956
rect 22094 6944 22100 6956
rect 22152 6944 22158 6996
rect 24394 6916 24400 6928
rect 19306 6888 24400 6916
rect 24394 6876 24400 6888
rect 24452 6876 24458 6928
rect 18325 6851 18383 6857
rect 18325 6817 18337 6851
rect 18371 6817 18383 6851
rect 18325 6811 18383 6817
rect 18414 6808 18420 6860
rect 18472 6808 18478 6860
rect 18693 6851 18751 6857
rect 18693 6817 18705 6851
rect 18739 6848 18751 6851
rect 19426 6848 19432 6860
rect 18739 6820 19432 6848
rect 18739 6817 18751 6820
rect 18693 6811 18751 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 21013 6820 23060 6848
rect 17037 6783 17095 6789
rect 17037 6780 17049 6783
rect 16632 6752 17049 6780
rect 16632 6740 16638 6752
rect 17037 6749 17049 6752
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 17770 6780 17776 6792
rect 17368 6752 17776 6780
rect 17368 6740 17374 6752
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 18046 6740 18052 6792
rect 18104 6740 18110 6792
rect 18156 6780 18184 6808
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 18156 6752 18521 6780
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 18877 6783 18935 6789
rect 18877 6780 18889 6783
rect 18840 6752 18889 6780
rect 18840 6740 18846 6752
rect 18877 6749 18889 6752
rect 18923 6749 18935 6783
rect 18877 6743 18935 6749
rect 19058 6740 19064 6792
rect 19116 6740 19122 6792
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 21013 6780 21041 6820
rect 19208 6752 21041 6780
rect 19208 6740 19214 6752
rect 21082 6740 21088 6792
rect 21140 6740 21146 6792
rect 23032 6789 23060 6820
rect 23017 6783 23075 6789
rect 23017 6749 23029 6783
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 13504 6684 14504 6712
rect 13504 6672 13510 6684
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 14829 6715 14887 6721
rect 14829 6712 14841 6715
rect 14700 6684 14841 6712
rect 14700 6672 14706 6684
rect 14829 6681 14841 6684
rect 14875 6681 14887 6715
rect 14829 6675 14887 6681
rect 13354 6644 13360 6656
rect 13004 6616 13360 6644
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13633 6647 13691 6653
rect 13633 6613 13645 6647
rect 13679 6644 13691 6647
rect 13722 6644 13728 6656
rect 13679 6616 13728 6644
rect 13679 6613 13691 6616
rect 13633 6607 13691 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 13906 6604 13912 6656
rect 13964 6604 13970 6656
rect 14366 6604 14372 6656
rect 14424 6604 14430 6656
rect 14550 6604 14556 6656
rect 14608 6604 14614 6656
rect 14844 6644 14872 6675
rect 15010 6672 15016 6724
rect 15068 6712 15074 6724
rect 16482 6712 16488 6724
rect 15068 6684 16488 6712
rect 15068 6672 15074 6684
rect 16482 6672 16488 6684
rect 16540 6672 16546 6724
rect 16942 6672 16948 6724
rect 17000 6672 17006 6724
rect 17052 6684 19196 6712
rect 15286 6644 15292 6656
rect 14844 6616 15292 6644
rect 15286 6604 15292 6616
rect 15344 6644 15350 6656
rect 15562 6644 15568 6656
rect 15344 6616 15568 6644
rect 15344 6604 15350 6616
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 15654 6604 15660 6656
rect 15712 6604 15718 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 16666 6644 16672 6656
rect 16264 6616 16672 6644
rect 16264 6604 16270 6616
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 17052 6644 17080 6684
rect 16908 6616 17080 6644
rect 17129 6647 17187 6653
rect 16908 6604 16914 6616
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17494 6644 17500 6656
rect 17175 6616 17500 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 19058 6644 19064 6656
rect 17920 6616 19064 6644
rect 17920 6604 17926 6616
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19168 6644 19196 6684
rect 19242 6672 19248 6724
rect 19300 6672 19306 6724
rect 21174 6672 21180 6724
rect 21232 6712 21238 6724
rect 21232 6684 21956 6712
rect 21232 6672 21238 6684
rect 20533 6647 20591 6653
rect 20533 6644 20545 6647
rect 19168 6616 20545 6644
rect 20533 6613 20545 6616
rect 20579 6613 20591 6647
rect 20533 6607 20591 6613
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 21818 6644 21824 6656
rect 20772 6616 21824 6644
rect 20772 6604 20778 6616
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 21928 6644 21956 6684
rect 22186 6672 22192 6724
rect 22244 6712 22250 6724
rect 22554 6712 22560 6724
rect 22244 6684 22560 6712
rect 22244 6672 22250 6684
rect 22554 6672 22560 6684
rect 22612 6712 22618 6724
rect 22649 6715 22707 6721
rect 22649 6712 22661 6715
rect 22612 6684 22661 6712
rect 22612 6672 22618 6684
rect 22649 6681 22661 6684
rect 22695 6681 22707 6715
rect 22649 6675 22707 6681
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 21928 6616 23213 6644
rect 23201 6613 23213 6616
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 1104 6554 23644 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 23644 6554
rect 1104 6480 23644 6502
rect 1578 6400 1584 6452
rect 1636 6400 1642 6452
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 1949 6443 2007 6449
rect 1949 6440 1961 6443
rect 1728 6412 1961 6440
rect 1728 6400 1734 6412
rect 1949 6409 1961 6412
rect 1995 6409 2007 6443
rect 1949 6403 2007 6409
rect 4062 6400 4068 6452
rect 4120 6400 4126 6452
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 7282 6440 7288 6452
rect 4764 6412 7288 6440
rect 4764 6400 4770 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 8720 6412 9597 6440
rect 8720 6400 8726 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 10410 6440 10416 6452
rect 9815 6412 10416 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 12894 6440 12900 6452
rect 12084 6412 12900 6440
rect 4525 6375 4583 6381
rect 4525 6372 4537 6375
rect 3436 6344 4537 6372
rect 750 6264 756 6316
rect 808 6304 814 6316
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 808 6276 1501 6304
rect 808 6264 814 6276
rect 1489 6273 1501 6276
rect 1535 6273 1547 6307
rect 1489 6267 1547 6273
rect 2130 6264 2136 6316
rect 2188 6264 2194 6316
rect 3326 6264 3332 6316
rect 3384 6304 3390 6316
rect 3436 6313 3464 6344
rect 4525 6341 4537 6344
rect 4571 6341 4583 6375
rect 4525 6335 4583 6341
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 6512 6344 11928 6372
rect 6512 6332 6518 6344
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3384 6276 3433 6304
rect 3384 6264 3390 6276
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3970 6264 3976 6316
rect 4028 6264 4034 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4246 6304 4252 6316
rect 4203 6276 4252 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 4890 6304 4896 6316
rect 4396 6276 4896 6304
rect 4396 6264 4402 6276
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5626 6304 5632 6316
rect 5215 6276 5632 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6236 3663 6239
rect 4062 6236 4068 6248
rect 3651 6208 4068 6236
rect 3651 6205 3663 6208
rect 3605 6199 3663 6205
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 5092 6236 5120 6267
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8352 6276 9137 6304
rect 8352 6264 8358 6276
rect 9125 6273 9137 6276
rect 9171 6304 9183 6307
rect 9490 6304 9496 6316
rect 9171 6276 9496 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 9631 6307 9689 6313
rect 9631 6273 9643 6307
rect 9677 6304 9689 6307
rect 9766 6304 9772 6316
rect 9677 6276 9772 6304
rect 9677 6273 9689 6276
rect 9631 6267 9689 6273
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9916 6276 9965 6304
rect 9916 6264 9922 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10100 6276 10241 6304
rect 10100 6264 10106 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10376 6276 10977 6304
rect 10376 6264 10382 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 11790 6264 11796 6316
rect 11848 6264 11854 6316
rect 5718 6236 5724 6248
rect 4172 6208 5724 6236
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 4172 6168 4200 6208
rect 5718 6196 5724 6208
rect 5776 6236 5782 6248
rect 10134 6236 10140 6248
rect 5776 6208 10140 6236
rect 5776 6196 5782 6208
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10778 6196 10784 6248
rect 10836 6196 10842 6248
rect 10873 6239 10931 6245
rect 10873 6205 10885 6239
rect 10919 6205 10931 6239
rect 10873 6199 10931 6205
rect 3568 6140 4200 6168
rect 4341 6171 4399 6177
rect 3568 6128 3574 6140
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 4614 6168 4620 6180
rect 4387 6140 4620 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 4614 6128 4620 6140
rect 4672 6128 4678 6180
rect 4890 6128 4896 6180
rect 4948 6128 4954 6180
rect 4982 6128 4988 6180
rect 5040 6168 5046 6180
rect 5442 6168 5448 6180
rect 5040 6140 5448 6168
rect 5040 6128 5046 6140
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 7834 6128 7840 6180
rect 7892 6168 7898 6180
rect 10042 6168 10048 6180
rect 7892 6140 10048 6168
rect 7892 6128 7898 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10686 6168 10692 6180
rect 10336 6140 10692 6168
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 4706 6100 4712 6112
rect 4580 6072 4712 6100
rect 4580 6060 4586 6072
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5353 6103 5411 6109
rect 5353 6069 5365 6103
rect 5399 6100 5411 6103
rect 5534 6100 5540 6112
rect 5399 6072 5540 6100
rect 5399 6069 5411 6072
rect 5353 6063 5411 6069
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 9582 6100 9588 6112
rect 9263 6072 9588 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10336 6109 10364 6140
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6069 10379 6103
rect 10321 6063 10379 6069
rect 10502 6060 10508 6112
rect 10560 6060 10566 6112
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 10888 6100 10916 6199
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11330 6236 11336 6248
rect 11112 6208 11336 6236
rect 11112 6196 11118 6208
rect 11330 6196 11336 6208
rect 11388 6196 11394 6248
rect 11900 6236 11928 6344
rect 11974 6264 11980 6316
rect 12032 6264 12038 6316
rect 12084 6313 12112 6412
rect 12894 6400 12900 6412
rect 12952 6400 12958 6452
rect 13630 6400 13636 6452
rect 13688 6400 13694 6452
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 14660 6412 15240 6440
rect 12710 6332 12716 6384
rect 12768 6332 12774 6384
rect 14568 6372 14596 6403
rect 13832 6344 14596 6372
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12250 6264 12256 6316
rect 12308 6264 12314 6316
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 12438 6307 12496 6313
rect 12438 6273 12450 6307
rect 12484 6304 12496 6307
rect 12526 6304 12532 6316
rect 12484 6276 12532 6304
rect 12484 6273 12496 6276
rect 12438 6267 12496 6273
rect 12360 6236 12388 6267
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 13035 6276 13737 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13004 6236 13032 6267
rect 11900 6208 12388 6236
rect 12544 6208 13032 6236
rect 13357 6239 13415 6245
rect 11977 6171 12035 6177
rect 11977 6137 11989 6171
rect 12023 6168 12035 6171
rect 12434 6168 12440 6180
rect 12023 6140 12440 6168
rect 12023 6137 12035 6140
rect 11977 6131 12035 6137
rect 12434 6128 12440 6140
rect 12492 6128 12498 6180
rect 10652 6072 10916 6100
rect 10652 6060 10658 6072
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12544 6100 12572 6208
rect 13357 6205 13369 6239
rect 13403 6205 13415 6239
rect 13357 6199 13415 6205
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6236 13507 6239
rect 13630 6236 13636 6248
rect 13495 6208 13636 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 12802 6128 12808 6180
rect 12860 6168 12866 6180
rect 13372 6168 13400 6199
rect 13630 6196 13636 6208
rect 13688 6196 13694 6248
rect 13832 6168 13860 6344
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6304 14611 6307
rect 14660 6304 14688 6412
rect 15212 6384 15240 6412
rect 15378 6400 15384 6452
rect 15436 6400 15442 6452
rect 16298 6400 16304 6452
rect 16356 6440 16362 6452
rect 16356 6412 22692 6440
rect 16356 6400 16362 6412
rect 15013 6375 15071 6381
rect 15013 6372 15025 6375
rect 14844 6344 15025 6372
rect 14599 6276 14688 6304
rect 14730 6307 14788 6313
rect 14730 6282 14742 6307
rect 14776 6304 14788 6307
rect 14844 6304 14872 6344
rect 15013 6341 15025 6344
rect 15059 6341 15071 6375
rect 15013 6335 15071 6341
rect 15194 6332 15200 6384
rect 15252 6372 15258 6384
rect 15289 6375 15347 6381
rect 15289 6372 15301 6375
rect 15252 6344 15301 6372
rect 15252 6332 15258 6344
rect 15289 6341 15301 6344
rect 15335 6341 15347 6375
rect 15396 6372 15424 6400
rect 15396 6344 16068 6372
rect 15289 6335 15347 6341
rect 14776 6282 14872 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 14730 6267 14740 6282
rect 14792 6276 14872 6282
rect 14916 6307 14974 6313
rect 14090 6196 14096 6248
rect 14148 6196 14154 6248
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6236 14243 6239
rect 14231 6208 14596 6236
rect 14734 6230 14740 6267
rect 14792 6230 14798 6276
rect 14916 6273 14928 6307
rect 14962 6273 14974 6307
rect 14916 6267 14974 6273
rect 14931 6236 14959 6267
rect 15102 6264 15108 6316
rect 15160 6264 15166 6316
rect 15473 6307 15531 6313
rect 15473 6304 15485 6307
rect 15304 6276 15485 6304
rect 15304 6248 15332 6276
rect 15473 6273 15485 6276
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 16040 6313 16068 6344
rect 16390 6332 16396 6384
rect 16448 6372 16454 6384
rect 16448 6344 19748 6372
rect 16448 6332 16454 6344
rect 16025 6307 16083 6313
rect 15712 6276 15976 6304
rect 15712 6264 15718 6276
rect 15194 6236 15200 6248
rect 14931 6208 15200 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 12860 6140 13860 6168
rect 14568 6168 14596 6208
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 15286 6196 15292 6248
rect 15344 6196 15350 6248
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6205 15899 6239
rect 15948 6236 15976 6276
rect 16025 6273 16037 6307
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 16264 6276 16313 6304
rect 16264 6264 16270 6276
rect 16301 6273 16313 6276
rect 16347 6273 16359 6307
rect 16485 6307 16543 6313
rect 16485 6304 16497 6307
rect 16301 6267 16359 6273
rect 16408 6276 16497 6304
rect 16408 6236 16436 6276
rect 16485 6273 16497 6276
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 16850 6264 16856 6316
rect 16908 6264 16914 6316
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 15948 6208 16436 6236
rect 15841 6199 15899 6205
rect 14568 6140 14642 6168
rect 12860 6128 12866 6140
rect 11940 6072 12572 6100
rect 11940 6060 11946 6072
rect 13262 6060 13268 6112
rect 13320 6100 13326 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 13320 6072 14381 6100
rect 13320 6060 13326 6072
rect 14369 6069 14381 6072
rect 14415 6069 14427 6103
rect 14614 6100 14642 6140
rect 15102 6128 15108 6180
rect 15160 6168 15166 6180
rect 15562 6168 15568 6180
rect 15160 6140 15568 6168
rect 15160 6128 15166 6140
rect 15562 6128 15568 6140
rect 15620 6128 15626 6180
rect 15289 6103 15347 6109
rect 15289 6100 15301 6103
rect 14614 6072 15301 6100
rect 14369 6063 14427 6069
rect 15289 6069 15301 6072
rect 15335 6069 15347 6103
rect 15764 6100 15792 6199
rect 15856 6168 15884 6199
rect 16758 6196 16764 6248
rect 16816 6236 16822 6248
rect 16960 6236 16988 6267
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 17678 6304 17684 6316
rect 17092 6276 17684 6304
rect 17092 6264 17098 6276
rect 17678 6264 17684 6276
rect 17736 6264 17742 6316
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 19337 6307 19395 6313
rect 18288 6276 19288 6304
rect 18288 6264 18294 6276
rect 16816 6208 16988 6236
rect 17221 6239 17279 6245
rect 16816 6196 16822 6208
rect 17221 6205 17233 6239
rect 17267 6205 17279 6239
rect 17221 6199 17279 6205
rect 17405 6239 17463 6245
rect 17405 6205 17417 6239
rect 17451 6236 17463 6239
rect 19150 6236 19156 6248
rect 17451 6208 19156 6236
rect 17451 6205 17463 6208
rect 17405 6199 17463 6205
rect 16022 6168 16028 6180
rect 15856 6140 16028 6168
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 17236 6168 17264 6199
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19260 6236 19288 6276
rect 19337 6273 19349 6307
rect 19383 6304 19395 6307
rect 19610 6304 19616 6316
rect 19383 6276 19616 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 19720 6304 19748 6344
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 20073 6375 20131 6381
rect 20073 6372 20085 6375
rect 20036 6344 20085 6372
rect 20036 6332 20042 6344
rect 20073 6341 20085 6344
rect 20119 6341 20131 6375
rect 20073 6335 20131 6341
rect 20162 6332 20168 6384
rect 20220 6372 20226 6384
rect 20625 6375 20683 6381
rect 20625 6372 20637 6375
rect 20220 6344 20637 6372
rect 20220 6332 20226 6344
rect 20625 6341 20637 6344
rect 20671 6372 20683 6375
rect 20671 6344 21496 6372
rect 20671 6341 20683 6344
rect 20625 6335 20683 6341
rect 20441 6307 20499 6313
rect 20441 6304 20453 6307
rect 19720 6276 20453 6304
rect 20441 6273 20453 6276
rect 20487 6273 20499 6307
rect 20441 6267 20499 6273
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 20732 6236 20760 6267
rect 20990 6264 20996 6316
rect 21048 6304 21054 6316
rect 21085 6307 21143 6313
rect 21085 6304 21097 6307
rect 21048 6276 21097 6304
rect 21048 6264 21054 6276
rect 21085 6273 21097 6276
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 21358 6264 21364 6316
rect 21416 6264 21422 6316
rect 21468 6304 21496 6344
rect 21818 6332 21824 6384
rect 21876 6332 21882 6384
rect 21910 6332 21916 6384
rect 21968 6332 21974 6384
rect 21468 6276 22094 6304
rect 21542 6236 21548 6248
rect 19260 6208 21548 6236
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 21634 6196 21640 6248
rect 21692 6236 21698 6248
rect 21910 6236 21916 6248
rect 21692 6208 21916 6236
rect 21692 6196 21698 6208
rect 21910 6196 21916 6208
rect 21968 6196 21974 6248
rect 22066 6236 22094 6276
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 22664 6313 22692 6412
rect 22649 6307 22707 6313
rect 22649 6273 22661 6307
rect 22695 6273 22707 6307
rect 22649 6267 22707 6273
rect 22738 6264 22744 6316
rect 22796 6264 22802 6316
rect 22925 6307 22983 6313
rect 22925 6273 22937 6307
rect 22971 6273 22983 6307
rect 22925 6267 22983 6273
rect 22301 6239 22359 6245
rect 22301 6236 22313 6239
rect 22066 6208 22313 6236
rect 22301 6205 22313 6208
rect 22347 6205 22359 6239
rect 22301 6199 22359 6205
rect 22646 6168 22652 6180
rect 17236 6140 22652 6168
rect 22646 6128 22652 6140
rect 22704 6168 22710 6180
rect 22940 6168 22968 6267
rect 23014 6264 23020 6316
rect 23072 6264 23078 6316
rect 22704 6140 22968 6168
rect 22704 6128 22710 6140
rect 15838 6100 15844 6112
rect 15764 6072 15844 6100
rect 15289 6063 15347 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 16114 6060 16120 6112
rect 16172 6100 16178 6112
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 16172 6072 16221 6100
rect 16172 6060 16178 6072
rect 16209 6069 16221 6072
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 16485 6103 16543 6109
rect 16485 6069 16497 6103
rect 16531 6100 16543 6103
rect 17586 6100 17592 6112
rect 16531 6072 17592 6100
rect 16531 6069 16543 6072
rect 16485 6063 16543 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 18046 6060 18052 6112
rect 18104 6060 18110 6112
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 21634 6100 21640 6112
rect 18840 6072 21640 6100
rect 18840 6060 18846 6072
rect 21634 6060 21640 6072
rect 21692 6060 21698 6112
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 22465 6103 22523 6109
rect 22465 6100 22477 6103
rect 22152 6072 22477 6100
rect 22152 6060 22158 6072
rect 22465 6069 22477 6072
rect 22511 6069 22523 6103
rect 22465 6063 22523 6069
rect 23198 6060 23204 6112
rect 23256 6060 23262 6112
rect 1104 6010 23644 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 23644 6010
rect 1104 5936 23644 5958
rect 5353 5899 5411 5905
rect 5353 5865 5365 5899
rect 5399 5896 5411 5899
rect 5626 5896 5632 5908
rect 5399 5868 5632 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8294 5896 8300 5908
rect 8067 5868 8300 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 9030 5896 9036 5908
rect 8435 5868 9036 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9582 5856 9588 5908
rect 9640 5856 9646 5908
rect 10318 5896 10324 5908
rect 9871 5868 10324 5896
rect 1949 5831 2007 5837
rect 1949 5797 1961 5831
rect 1995 5797 2007 5831
rect 1949 5791 2007 5797
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 1964 5692 1992 5791
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 4028 5800 4200 5828
rect 4028 5788 4034 5800
rect 4172 5769 4200 5800
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 4985 5831 5043 5837
rect 4985 5828 4997 5831
rect 4856 5800 4997 5828
rect 4856 5788 4862 5800
rect 4985 5797 4997 5800
rect 5031 5828 5043 5831
rect 5442 5828 5448 5840
rect 5031 5800 5448 5828
rect 5031 5797 5043 5800
rect 4985 5791 5043 5797
rect 5442 5788 5448 5800
rect 5500 5828 5506 5840
rect 9871 5828 9899 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 10836 5868 11376 5896
rect 10836 5856 10842 5868
rect 5500 5800 9899 5828
rect 5500 5788 5506 5800
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 10413 5831 10471 5837
rect 10413 5828 10425 5831
rect 10192 5800 10425 5828
rect 10192 5788 10198 5800
rect 10413 5797 10425 5800
rect 10459 5828 10471 5831
rect 10459 5800 11008 5828
rect 10459 5797 10471 5800
rect 10413 5791 10471 5797
rect 4157 5763 4215 5769
rect 4157 5729 4169 5763
rect 4203 5760 4215 5763
rect 5077 5763 5135 5769
rect 4203 5732 5028 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 5000 5704 5028 5732
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 5626 5760 5632 5772
rect 5123 5732 5632 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 8846 5760 8852 5772
rect 7668 5732 8852 5760
rect 7668 5704 7696 5732
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 9732 5732 10517 5760
rect 9732 5720 9738 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10870 5760 10876 5772
rect 10505 5723 10563 5729
rect 10704 5732 10876 5760
rect 1719 5664 1992 5692
rect 2133 5695 2191 5701
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 3970 5692 3976 5704
rect 2179 5664 3976 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4614 5692 4620 5704
rect 4387 5664 4620 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4816 5624 4844 5655
rect 4982 5652 4988 5704
rect 5040 5652 5046 5704
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 5258 5692 5264 5704
rect 5215 5664 5264 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 5810 5692 5816 5704
rect 5767 5664 5816 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 9766 5692 9772 5704
rect 8527 5664 9772 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 4212 5596 7972 5624
rect 4212 5584 4218 5596
rect 750 5516 756 5568
rect 808 5556 814 5568
rect 1489 5559 1547 5565
rect 1489 5556 1501 5559
rect 808 5528 1501 5556
rect 808 5516 814 5528
rect 1489 5525 1501 5528
rect 1535 5525 1547 5559
rect 1489 5519 1547 5525
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 4525 5559 4583 5565
rect 4525 5556 4537 5559
rect 4488 5528 4537 5556
rect 4488 5516 4494 5528
rect 4525 5525 4537 5528
rect 4571 5525 4583 5559
rect 4525 5519 4583 5525
rect 4614 5516 4620 5568
rect 4672 5516 4678 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 6730 5556 6736 5568
rect 5951 5528 6736 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7944 5556 7972 5596
rect 8018 5584 8024 5636
rect 8076 5624 8082 5636
rect 9968 5624 9996 5655
rect 10042 5652 10048 5704
rect 10100 5652 10106 5704
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10410 5692 10416 5704
rect 10367 5664 10416 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10134 5624 10140 5636
rect 8076 5596 9904 5624
rect 9968 5596 10140 5624
rect 8076 5584 8082 5596
rect 9674 5556 9680 5568
rect 7944 5528 9680 5556
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 9876 5556 9904 5596
rect 10134 5584 10140 5596
rect 10192 5584 10198 5636
rect 10244 5624 10272 5655
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 10704 5701 10732 5732
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 10778 5652 10784 5704
rect 10836 5652 10842 5704
rect 10980 5701 11008 5800
rect 11348 5769 11376 5868
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 12032 5868 12357 5896
rect 12032 5856 12038 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 13504 5868 13553 5896
rect 13504 5856 13510 5868
rect 13541 5865 13553 5868
rect 13587 5865 13599 5899
rect 13541 5859 13599 5865
rect 11606 5788 11612 5840
rect 11664 5828 11670 5840
rect 13081 5831 13139 5837
rect 13081 5828 13093 5831
rect 11664 5800 13093 5828
rect 11664 5788 11670 5800
rect 13081 5797 13093 5800
rect 13127 5797 13139 5831
rect 13081 5791 13139 5797
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5760 11391 5763
rect 12158 5760 12164 5772
rect 11379 5732 12164 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 13262 5760 13268 5772
rect 12636 5732 13268 5760
rect 12636 5701 12664 5732
rect 13262 5720 13268 5732
rect 13320 5720 13326 5772
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5661 11023 5695
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 10965 5655 11023 5661
rect 11072 5664 12541 5692
rect 10502 5624 10508 5636
rect 10244 5596 10508 5624
rect 10502 5584 10508 5596
rect 10560 5624 10566 5636
rect 11072 5624 11100 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12802 5652 12808 5704
rect 12860 5652 12866 5704
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13170 5692 13176 5704
rect 13127 5664 13176 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13556 5636 13584 5859
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 13909 5899 13967 5905
rect 13909 5896 13921 5899
rect 13780 5868 13921 5896
rect 13780 5856 13786 5868
rect 13909 5865 13921 5868
rect 13955 5865 13967 5899
rect 14553 5899 14611 5905
rect 14553 5896 14565 5899
rect 13909 5859 13967 5865
rect 14298 5868 14565 5896
rect 13630 5788 13636 5840
rect 13688 5828 13694 5840
rect 14298 5828 14326 5868
rect 14553 5865 14565 5868
rect 14599 5865 14611 5899
rect 15194 5896 15200 5908
rect 14553 5859 14611 5865
rect 14844 5868 15200 5896
rect 13688 5800 14326 5828
rect 13688 5788 13694 5800
rect 14642 5788 14648 5840
rect 14700 5788 14706 5840
rect 14844 5760 14872 5868
rect 15194 5856 15200 5868
rect 15252 5896 15258 5908
rect 15289 5899 15347 5905
rect 15289 5896 15301 5899
rect 15252 5868 15301 5896
rect 15252 5856 15258 5868
rect 15289 5865 15301 5868
rect 15335 5865 15347 5899
rect 15289 5859 15347 5865
rect 16390 5856 16396 5908
rect 16448 5856 16454 5908
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 17402 5896 17408 5908
rect 16908 5868 17408 5896
rect 16908 5856 16914 5868
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18322 5856 18328 5908
rect 18380 5896 18386 5908
rect 18969 5899 19027 5905
rect 18380 5868 18644 5896
rect 18380 5856 18386 5868
rect 15378 5788 15384 5840
rect 15436 5828 15442 5840
rect 15436 5800 15516 5828
rect 15436 5788 15442 5800
rect 15488 5769 15516 5800
rect 16482 5788 16488 5840
rect 16540 5828 16546 5840
rect 16758 5828 16764 5840
rect 16540 5800 16764 5828
rect 16540 5788 16546 5800
rect 16758 5788 16764 5800
rect 16816 5828 16822 5840
rect 16816 5800 17724 5828
rect 16816 5788 16822 5800
rect 14291 5732 14872 5760
rect 15473 5763 15531 5769
rect 14291 5712 14319 5732
rect 15473 5729 15485 5763
rect 15519 5729 15531 5763
rect 15473 5723 15531 5729
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 15896 5732 17417 5760
rect 15896 5720 15902 5732
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 17405 5723 17463 5729
rect 14200 5711 14319 5712
rect 14180 5705 14319 5711
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 13998 5692 14004 5704
rect 13771 5664 14004 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 10560 5596 11100 5624
rect 11149 5627 11207 5633
rect 10560 5584 10566 5596
rect 11149 5593 11161 5627
rect 11195 5624 11207 5627
rect 11238 5624 11244 5636
rect 11195 5596 11244 5624
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 12345 5627 12403 5633
rect 12345 5624 12357 5627
rect 11388 5596 12357 5624
rect 11388 5584 11394 5596
rect 12345 5593 12357 5596
rect 12391 5624 12403 5627
rect 12434 5624 12440 5636
rect 12391 5596 12440 5624
rect 12391 5593 12403 5596
rect 12345 5587 12403 5593
rect 12434 5584 12440 5596
rect 12492 5584 12498 5636
rect 12897 5627 12955 5633
rect 12897 5624 12909 5627
rect 12544 5596 12909 5624
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 9876 5528 10609 5556
rect 10597 5525 10609 5528
rect 10643 5556 10655 5559
rect 11054 5556 11060 5568
rect 10643 5528 11060 5556
rect 10643 5525 10655 5528
rect 10597 5519 10655 5525
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12544 5556 12572 5596
rect 12897 5593 12909 5596
rect 12943 5593 12955 5627
rect 12897 5587 12955 5593
rect 12986 5584 12992 5636
rect 13044 5624 13050 5636
rect 13449 5627 13507 5633
rect 13449 5624 13461 5627
rect 13044 5596 13461 5624
rect 13044 5584 13050 5596
rect 13449 5593 13461 5596
rect 13495 5593 13507 5627
rect 13449 5587 13507 5593
rect 13538 5584 13544 5636
rect 13596 5584 13602 5636
rect 13648 5624 13676 5655
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 14180 5671 14192 5705
rect 14226 5684 14319 5705
rect 14369 5695 14427 5701
rect 14226 5671 14238 5684
rect 14180 5665 14238 5671
rect 14369 5661 14381 5695
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 13906 5624 13912 5636
rect 13648 5596 13912 5624
rect 13906 5584 13912 5596
rect 13964 5584 13970 5636
rect 14277 5627 14335 5633
rect 14277 5593 14289 5627
rect 14323 5593 14335 5627
rect 14384 5624 14412 5655
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15010 5652 15016 5704
rect 15068 5652 15074 5704
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5692 15255 5695
rect 15286 5692 15292 5704
rect 15243 5664 15292 5692
rect 15243 5661 15255 5664
rect 15197 5655 15255 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 15396 5664 15577 5692
rect 15396 5636 15424 5664
rect 15565 5661 15577 5664
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 16114 5652 16120 5704
rect 16172 5652 16178 5704
rect 16206 5652 16212 5704
rect 16264 5652 16270 5704
rect 16316 5664 16712 5692
rect 15102 5624 15108 5636
rect 14384 5596 15108 5624
rect 14277 5587 14335 5593
rect 11848 5528 12572 5556
rect 13265 5559 13323 5565
rect 11848 5516 11854 5528
rect 13265 5525 13277 5559
rect 13311 5556 13323 5559
rect 13354 5556 13360 5568
rect 13311 5528 13360 5556
rect 13311 5525 13323 5528
rect 13265 5519 13323 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 14291 5556 14319 5587
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 15378 5584 15384 5636
rect 15436 5584 15442 5636
rect 15841 5627 15899 5633
rect 15841 5593 15853 5627
rect 15887 5593 15899 5627
rect 15948 5624 15976 5652
rect 16316 5624 16344 5664
rect 15948 5596 16344 5624
rect 16393 5627 16451 5633
rect 15841 5587 15899 5593
rect 16393 5593 16405 5627
rect 16439 5593 16451 5627
rect 16684 5624 16712 5664
rect 16758 5652 16764 5704
rect 16816 5652 16822 5704
rect 16850 5652 16856 5704
rect 16908 5652 16914 5704
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5661 17003 5695
rect 16945 5655 17003 5661
rect 16960 5624 16988 5655
rect 17126 5652 17132 5704
rect 17184 5652 17190 5704
rect 17586 5652 17592 5704
rect 17644 5652 17650 5704
rect 17696 5692 17724 5800
rect 18230 5788 18236 5840
rect 18288 5828 18294 5840
rect 18509 5831 18567 5837
rect 18509 5828 18521 5831
rect 18288 5800 18521 5828
rect 18288 5788 18294 5800
rect 18509 5797 18521 5800
rect 18555 5797 18567 5831
rect 18616 5828 18644 5868
rect 18969 5865 18981 5899
rect 19015 5896 19027 5899
rect 19518 5896 19524 5908
rect 19015 5868 19524 5896
rect 19015 5865 19027 5868
rect 18969 5859 19027 5865
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20530 5856 20536 5908
rect 20588 5856 20594 5908
rect 21361 5831 21419 5837
rect 21361 5828 21373 5831
rect 18616 5800 21373 5828
rect 18509 5791 18567 5797
rect 21361 5797 21373 5800
rect 21407 5797 21419 5831
rect 21361 5791 21419 5797
rect 21634 5788 21640 5840
rect 21692 5828 21698 5840
rect 23198 5828 23204 5840
rect 21692 5800 23204 5828
rect 21692 5788 21698 5800
rect 23198 5788 23204 5800
rect 23256 5788 23262 5840
rect 18966 5720 18972 5772
rect 19024 5760 19030 5772
rect 20622 5760 20628 5772
rect 19024 5732 20628 5760
rect 19024 5720 19030 5732
rect 20622 5720 20628 5732
rect 20680 5720 20686 5772
rect 21468 5732 22094 5760
rect 21468 5704 21496 5732
rect 17954 5692 17960 5704
rect 17696 5664 17960 5692
rect 17954 5652 17960 5664
rect 18012 5692 18018 5704
rect 18049 5695 18107 5701
rect 18049 5692 18061 5695
rect 18012 5664 18061 5692
rect 18012 5652 18018 5664
rect 18049 5661 18061 5664
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 18141 5695 18199 5701
rect 18141 5661 18153 5695
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 16684 5596 16988 5624
rect 16393 5587 16451 5593
rect 14366 5556 14372 5568
rect 14291 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 15856 5556 15884 5587
rect 16114 5556 16120 5568
rect 15856 5528 16120 5556
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16408 5556 16436 5587
rect 17218 5584 17224 5636
rect 17276 5624 17282 5636
rect 18156 5624 18184 5655
rect 18874 5652 18880 5704
rect 18932 5652 18938 5704
rect 21450 5652 21456 5704
rect 21508 5652 21514 5704
rect 21542 5652 21548 5704
rect 21600 5652 21606 5704
rect 22066 5692 22094 5732
rect 23109 5695 23167 5701
rect 23109 5692 23121 5695
rect 22066 5664 23121 5692
rect 23109 5661 23121 5664
rect 23155 5661 23167 5695
rect 23109 5655 23167 5661
rect 17276 5596 18184 5624
rect 17276 5584 17282 5596
rect 18230 5584 18236 5636
rect 18288 5624 18294 5636
rect 19245 5627 19303 5633
rect 19245 5624 19257 5627
rect 18288 5596 19257 5624
rect 18288 5584 18294 5596
rect 19245 5593 19257 5596
rect 19291 5593 19303 5627
rect 19245 5587 19303 5593
rect 16485 5559 16543 5565
rect 16485 5556 16497 5559
rect 16408 5528 16497 5556
rect 16485 5525 16497 5528
rect 16531 5525 16543 5559
rect 16485 5519 16543 5525
rect 1104 5466 23644 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 23644 5466
rect 1104 5392 23644 5414
rect 3970 5312 3976 5364
rect 4028 5312 4034 5364
rect 4985 5355 5043 5361
rect 4080 5324 4936 5352
rect 566 5176 572 5228
rect 624 5216 630 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 624 5188 1501 5216
rect 624 5176 630 5188
rect 1489 5185 1501 5188
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4080 5216 4108 5324
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 4908 5284 4936 5324
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 6178 5352 6184 5364
rect 5031 5324 6184 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7006 5352 7012 5364
rect 6604 5324 6684 5352
rect 6604 5312 6610 5324
rect 6656 5293 6684 5324
rect 6748 5324 7012 5352
rect 6748 5293 6776 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 7156 5324 7420 5352
rect 7156 5312 7162 5324
rect 6641 5287 6699 5293
rect 4387 5256 4844 5284
rect 4908 5256 6500 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 3936 5188 4108 5216
rect 3936 5176 3942 5188
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4430 5176 4436 5228
rect 4488 5176 4494 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4614 5216 4620 5228
rect 4571 5188 4620 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4816 5225 4844 5256
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5350 5216 5356 5228
rect 5307 5188 5356 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 4724 5080 4752 5179
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5460 5225 5488 5256
rect 6472 5228 6500 5256
rect 6641 5253 6653 5287
rect 6687 5253 6699 5287
rect 6641 5247 6699 5253
rect 6733 5287 6791 5293
rect 6733 5253 6745 5287
rect 6779 5253 6791 5287
rect 6733 5247 6791 5253
rect 6822 5244 6828 5296
rect 6880 5293 6886 5296
rect 6880 5287 6909 5293
rect 6897 5253 6909 5287
rect 7392 5284 7420 5324
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7524 5324 7849 5352
rect 7524 5312 7530 5324
rect 7837 5321 7849 5324
rect 7883 5352 7895 5355
rect 8018 5352 8024 5364
rect 7883 5324 8024 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8481 5355 8539 5361
rect 8481 5321 8493 5355
rect 8527 5352 8539 5355
rect 8570 5352 8576 5364
rect 8527 5324 8576 5352
rect 8527 5321 8539 5324
rect 8481 5315 8539 5321
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11241 5355 11299 5361
rect 11241 5352 11253 5355
rect 11204 5324 11253 5352
rect 11204 5312 11210 5324
rect 11241 5321 11253 5324
rect 11287 5321 11299 5355
rect 11241 5315 11299 5321
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 15286 5352 15292 5364
rect 13504 5324 15292 5352
rect 13504 5312 13510 5324
rect 11330 5284 11336 5296
rect 7392 5256 11336 5284
rect 6880 5247 6909 5253
rect 6880 5244 6886 5247
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 11606 5244 11612 5296
rect 11664 5284 11670 5296
rect 11664 5256 11836 5284
rect 11664 5244 11670 5256
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5534 5176 5540 5228
rect 5592 5176 5598 5228
rect 5626 5176 5632 5228
rect 5684 5176 5690 5228
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 5776 5188 5825 5216
rect 5776 5176 5782 5188
rect 5813 5185 5825 5188
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5828 5148 5856 5179
rect 6454 5176 6460 5228
rect 6512 5214 6518 5228
rect 6549 5219 6607 5225
rect 6549 5214 6561 5219
rect 6512 5186 6561 5214
rect 6512 5176 6518 5186
rect 6549 5185 6561 5186
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 7374 5176 7380 5228
rect 7432 5176 7438 5228
rect 7466 5176 7472 5228
rect 7524 5176 7530 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 7834 5216 7840 5228
rect 7699 5188 7840 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 7834 5176 7840 5188
rect 7892 5216 7898 5228
rect 7892 5188 8156 5216
rect 7892 5176 7898 5188
rect 6178 5148 6184 5160
rect 5828 5120 6184 5148
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 8128 5148 8156 5188
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8260 5188 8309 5216
rect 8260 5176 8266 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8536 5188 8585 5216
rect 8536 5176 8542 5188
rect 8573 5185 8585 5188
rect 8619 5216 8631 5219
rect 8938 5216 8944 5228
rect 8619 5188 8944 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11422 5216 11428 5228
rect 11195 5188 11428 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 11514 5176 11520 5228
rect 11572 5176 11578 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11808 5216 11836 5256
rect 12434 5244 12440 5296
rect 12492 5284 12498 5296
rect 12713 5287 12771 5293
rect 12713 5284 12725 5287
rect 12492 5256 12725 5284
rect 12492 5244 12498 5256
rect 12713 5253 12725 5256
rect 12759 5253 12771 5287
rect 14090 5284 14096 5296
rect 12713 5247 12771 5253
rect 13004 5256 14096 5284
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11808 5188 11897 5216
rect 11701 5179 11759 5185
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 10778 5148 10784 5160
rect 7638 5120 8064 5148
rect 8128 5120 10784 5148
rect 4798 5080 4804 5092
rect 1719 5052 2774 5080
rect 4724 5052 4804 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 2746 5012 2774 5052
rect 4798 5040 4804 5052
rect 4856 5080 4862 5092
rect 6546 5080 6552 5092
rect 4856 5052 6552 5080
rect 4856 5040 4862 5052
rect 6546 5040 6552 5052
rect 6604 5080 6610 5092
rect 7638 5080 7666 5120
rect 6604 5052 7666 5080
rect 6604 5040 6610 5052
rect 7742 5040 7748 5092
rect 7800 5080 7806 5092
rect 7929 5083 7987 5089
rect 7929 5080 7941 5083
rect 7800 5052 7941 5080
rect 7800 5040 7806 5052
rect 7929 5049 7941 5052
rect 7975 5049 7987 5083
rect 8036 5080 8064 5120
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11716 5148 11744 5179
rect 11974 5176 11980 5228
rect 12032 5176 12038 5228
rect 12158 5176 12164 5228
rect 12216 5176 12222 5228
rect 13004 5225 13032 5256
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 15028 5293 15056 5324
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 15657 5355 15715 5361
rect 15657 5352 15669 5355
rect 15620 5324 15669 5352
rect 15620 5312 15626 5324
rect 15657 5321 15669 5324
rect 15703 5321 15715 5355
rect 15657 5315 15715 5321
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16390 5352 16396 5364
rect 15804 5324 16396 5352
rect 15804 5312 15810 5324
rect 16390 5312 16396 5324
rect 16448 5352 16454 5364
rect 16945 5355 17003 5361
rect 16945 5352 16957 5355
rect 16448 5324 16957 5352
rect 16448 5312 16454 5324
rect 16945 5321 16957 5324
rect 16991 5321 17003 5355
rect 17865 5355 17923 5361
rect 16945 5315 17003 5321
rect 17052 5324 17816 5352
rect 15013 5287 15071 5293
rect 15013 5253 15025 5287
rect 15059 5253 15071 5287
rect 15013 5247 15071 5253
rect 15102 5244 15108 5296
rect 15160 5244 15166 5296
rect 15396 5256 16528 5284
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13354 5176 13360 5228
rect 13412 5176 13418 5228
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5216 13967 5219
rect 13998 5216 14004 5228
rect 13955 5188 14004 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 11112 5120 11744 5148
rect 11112 5108 11118 5120
rect 11790 5108 11796 5160
rect 11848 5148 11854 5160
rect 13648 5148 13676 5179
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 14461 5219 14519 5225
rect 14461 5185 14473 5219
rect 14507 5216 14519 5219
rect 14642 5216 14648 5228
rect 14507 5188 14648 5216
rect 14507 5185 14519 5188
rect 14461 5179 14519 5185
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14884 5188 14933 5216
rect 14884 5176 14890 5188
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 14921 5179 14979 5185
rect 15028 5188 15301 5216
rect 14844 5148 14872 5176
rect 15028 5160 15056 5188
rect 15289 5185 15301 5188
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 11848 5120 13676 5148
rect 14292 5120 14872 5148
rect 11848 5108 11854 5120
rect 12250 5080 12256 5092
rect 8036 5052 12256 5080
rect 7929 5043 7987 5049
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 13906 5080 13912 5092
rect 12360 5052 13912 5080
rect 5902 5012 5908 5024
rect 2746 4984 5908 5012
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 12360 5012 12388 5052
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 14093 5083 14151 5089
rect 14093 5049 14105 5083
rect 14139 5080 14151 5083
rect 14182 5080 14188 5092
rect 14139 5052 14188 5080
rect 14139 5049 14151 5052
rect 14093 5043 14151 5049
rect 14182 5040 14188 5052
rect 14240 5040 14246 5092
rect 14292 5089 14320 5120
rect 15010 5108 15016 5160
rect 15068 5108 15074 5160
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15396 5148 15424 5256
rect 15562 5176 15568 5228
rect 15620 5176 15626 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15672 5188 15853 5216
rect 15672 5160 15700 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15930 5176 15936 5228
rect 15988 5176 15994 5228
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 16500 5225 16528 5256
rect 16666 5244 16672 5296
rect 16724 5284 16730 5296
rect 17052 5284 17080 5324
rect 16724 5256 17080 5284
rect 17129 5287 17187 5293
rect 16724 5244 16730 5256
rect 17129 5253 17141 5287
rect 17175 5284 17187 5287
rect 17586 5284 17592 5296
rect 17175 5256 17592 5284
rect 17175 5253 17187 5256
rect 17129 5247 17187 5253
rect 17586 5244 17592 5256
rect 17644 5244 17650 5296
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5185 16267 5219
rect 16209 5179 16267 5185
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5185 16543 5219
rect 16485 5179 16543 5185
rect 15252 5120 15424 5148
rect 15252 5108 15258 5120
rect 15654 5108 15660 5160
rect 15712 5108 15718 5160
rect 15746 5108 15752 5160
rect 15804 5148 15810 5160
rect 16224 5148 16252 5179
rect 17218 5176 17224 5228
rect 17276 5176 17282 5228
rect 17402 5216 17408 5228
rect 17363 5188 17408 5216
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 17788 5225 17816 5324
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 21082 5352 21088 5364
rect 17911 5324 21088 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 21634 5312 21640 5364
rect 21692 5352 21698 5364
rect 22462 5352 22468 5364
rect 21692 5324 22468 5352
rect 21692 5312 21698 5324
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 23014 5312 23020 5364
rect 23072 5352 23078 5364
rect 23109 5355 23167 5361
rect 23109 5352 23121 5355
rect 23072 5324 23121 5352
rect 23072 5312 23078 5324
rect 23109 5321 23121 5324
rect 23155 5321 23167 5355
rect 23109 5315 23167 5321
rect 17954 5244 17960 5296
rect 18012 5284 18018 5296
rect 18012 5256 18276 5284
rect 18012 5244 18018 5256
rect 18248 5225 18276 5256
rect 20162 5244 20168 5296
rect 20220 5244 20226 5296
rect 20806 5244 20812 5296
rect 20864 5284 20870 5296
rect 20864 5256 21864 5284
rect 20864 5244 20870 5256
rect 21836 5228 21864 5256
rect 17773 5219 17831 5225
rect 17773 5185 17785 5219
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5216 18383 5219
rect 18414 5216 18420 5228
rect 18371 5188 18420 5216
rect 18371 5185 18383 5188
rect 18325 5179 18383 5185
rect 17589 5151 17647 5157
rect 17589 5148 17601 5151
rect 15804 5120 17601 5148
rect 15804 5108 15810 5120
rect 17589 5117 17601 5120
rect 17635 5117 17647 5151
rect 18064 5148 18092 5179
rect 18414 5176 18420 5188
rect 18472 5176 18478 5228
rect 18874 5176 18880 5228
rect 18932 5216 18938 5228
rect 21174 5216 21180 5228
rect 18932 5188 21180 5216
rect 18932 5176 18938 5188
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 21266 5176 21272 5228
rect 21324 5216 21330 5228
rect 21361 5219 21419 5225
rect 21361 5216 21373 5219
rect 21324 5188 21373 5216
rect 21324 5176 21330 5188
rect 21361 5185 21373 5188
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 21634 5176 21640 5228
rect 21692 5176 21698 5228
rect 21818 5176 21824 5228
rect 21876 5176 21882 5228
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 22922 5216 22928 5228
rect 22879 5188 22928 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 22922 5176 22928 5188
rect 22980 5176 22986 5228
rect 23014 5176 23020 5228
rect 23072 5176 23078 5228
rect 23106 5176 23112 5228
rect 23164 5216 23170 5228
rect 23293 5219 23351 5225
rect 23293 5216 23305 5219
rect 23164 5188 23305 5216
rect 23164 5176 23170 5188
rect 23293 5185 23305 5188
rect 23339 5185 23351 5219
rect 23293 5179 23351 5185
rect 17589 5111 17647 5117
rect 17696 5120 18092 5148
rect 14277 5083 14335 5089
rect 14277 5049 14289 5083
rect 14323 5049 14335 5083
rect 14277 5043 14335 5049
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 14737 5083 14795 5089
rect 14737 5080 14749 5083
rect 14424 5052 14749 5080
rect 14424 5040 14430 5052
rect 14737 5049 14749 5052
rect 14783 5080 14795 5083
rect 17696 5080 17724 5120
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 21545 5151 21603 5157
rect 20772 5120 21496 5148
rect 20772 5108 20778 5120
rect 21177 5083 21235 5089
rect 21177 5080 21189 5083
rect 14783 5052 17724 5080
rect 17788 5052 21189 5080
rect 14783 5049 14795 5052
rect 14737 5043 14795 5049
rect 6512 4984 12388 5012
rect 12805 5015 12863 5021
rect 6512 4972 6518 4984
rect 12805 4981 12817 5015
rect 12851 5012 12863 5015
rect 13078 5012 13084 5024
rect 12851 4984 13084 5012
rect 12851 4981 12863 4984
rect 12805 4975 12863 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13170 4972 13176 5024
rect 13228 4972 13234 5024
rect 13538 4972 13544 5024
rect 13596 4972 13602 5024
rect 13814 4972 13820 5024
rect 13872 4972 13878 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14553 5015 14611 5021
rect 14553 5012 14565 5015
rect 14056 4984 14565 5012
rect 14056 4972 14062 4984
rect 14553 4981 14565 4984
rect 14599 4981 14611 5015
rect 14553 4975 14611 4981
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 15194 5012 15200 5024
rect 14700 4984 15200 5012
rect 14700 4972 14706 4984
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 16301 5015 16359 5021
rect 16301 5012 16313 5015
rect 15436 4984 16313 5012
rect 15436 4972 15442 4984
rect 16301 4981 16313 4984
rect 16347 4981 16359 5015
rect 16301 4975 16359 4981
rect 16666 4972 16672 5024
rect 16724 5012 16730 5024
rect 16761 5015 16819 5021
rect 16761 5012 16773 5015
rect 16724 4984 16773 5012
rect 16724 4972 16730 4984
rect 16761 4981 16773 4984
rect 16807 4981 16819 5015
rect 16761 4975 16819 4981
rect 16945 5015 17003 5021
rect 16945 4981 16957 5015
rect 16991 5012 17003 5015
rect 17034 5012 17040 5024
rect 16991 4984 17040 5012
rect 16991 4981 17003 4984
rect 16945 4975 17003 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 17678 4972 17684 5024
rect 17736 5012 17742 5024
rect 17788 5012 17816 5052
rect 21177 5049 21189 5052
rect 21223 5049 21235 5083
rect 21468 5080 21496 5120
rect 21545 5117 21557 5151
rect 21591 5148 21603 5151
rect 21726 5148 21732 5160
rect 21591 5120 21732 5148
rect 21591 5117 21603 5120
rect 21545 5111 21603 5117
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 22373 5151 22431 5157
rect 22373 5148 22385 5151
rect 21836 5120 22385 5148
rect 21836 5080 21864 5120
rect 22373 5117 22385 5120
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 21468 5052 21864 5080
rect 21177 5043 21235 5049
rect 22002 5040 22008 5092
rect 22060 5080 22066 5092
rect 22281 5083 22339 5089
rect 22281 5080 22293 5083
rect 22060 5052 22293 5080
rect 22060 5040 22066 5052
rect 22281 5049 22293 5052
rect 22327 5049 22339 5083
rect 22281 5043 22339 5049
rect 17736 4984 17816 5012
rect 17736 4972 17742 4984
rect 18966 4972 18972 5024
rect 19024 5012 19030 5024
rect 19242 5012 19248 5024
rect 19024 4984 19248 5012
rect 19024 4972 19030 4984
rect 19242 4972 19248 4984
rect 19300 5012 19306 5024
rect 19613 5015 19671 5021
rect 19613 5012 19625 5015
rect 19300 4984 19625 5012
rect 19300 4972 19306 4984
rect 19613 4981 19625 4984
rect 19659 4981 19671 5015
rect 19613 4975 19671 4981
rect 21637 5015 21695 5021
rect 21637 4981 21649 5015
rect 21683 5012 21695 5015
rect 21910 5012 21916 5024
rect 21683 4984 21916 5012
rect 21683 4981 21695 4984
rect 21637 4975 21695 4981
rect 21910 4972 21916 4984
rect 21968 4972 21974 5024
rect 22189 5015 22247 5021
rect 22189 4981 22201 5015
rect 22235 5012 22247 5015
rect 22370 5012 22376 5024
rect 22235 4984 22376 5012
rect 22235 4981 22247 4984
rect 22189 4975 22247 4981
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 22646 4972 22652 5024
rect 22704 4972 22710 5024
rect 1104 4922 23644 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 23644 4922
rect 1104 4848 23644 4870
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 5442 4808 5448 4820
rect 4571 4780 5448 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 6638 4808 6644 4820
rect 6503 4780 6644 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 8110 4808 8116 4820
rect 7800 4780 8116 4808
rect 7800 4768 7806 4780
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 8662 4768 8668 4820
rect 8720 4768 8726 4820
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8812 4780 9045 4808
rect 8812 4768 8818 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 11514 4808 11520 4820
rect 10836 4780 11520 4808
rect 10836 4768 10842 4780
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 12710 4808 12716 4820
rect 11808 4780 12716 4808
rect 4433 4743 4491 4749
rect 4433 4709 4445 4743
rect 4479 4740 4491 4743
rect 4706 4740 4712 4752
rect 4479 4712 4712 4740
rect 4479 4709 4491 4712
rect 4433 4703 4491 4709
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 4890 4700 4896 4752
rect 4948 4740 4954 4752
rect 5077 4743 5135 4749
rect 5077 4740 5089 4743
rect 4948 4712 5089 4740
rect 4948 4700 4954 4712
rect 5077 4709 5089 4712
rect 5123 4740 5135 4743
rect 5258 4740 5264 4752
rect 5123 4712 5264 4740
rect 5123 4709 5135 4712
rect 5077 4703 5135 4709
rect 5258 4700 5264 4712
rect 5316 4700 5322 4752
rect 5902 4700 5908 4752
rect 5960 4740 5966 4752
rect 7466 4740 7472 4752
rect 5960 4712 7472 4740
rect 5960 4700 5966 4712
rect 7466 4700 7472 4712
rect 7524 4740 7530 4752
rect 7926 4740 7932 4752
rect 7524 4712 7932 4740
rect 7524 4700 7530 4712
rect 7926 4700 7932 4712
rect 7984 4740 7990 4752
rect 7984 4712 8340 4740
rect 7984 4700 7990 4712
rect 5166 4632 5172 4684
rect 5224 4632 5230 4684
rect 6362 4672 6368 4684
rect 5920 4644 6368 4672
rect 5920 4613 5948 4644
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 8312 4672 8340 4712
rect 11238 4700 11244 4752
rect 11296 4700 11302 4752
rect 8570 4672 8576 4684
rect 7331 4644 8156 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 5994 4564 6000 4616
rect 6052 4564 6058 4616
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4604 6331 4607
rect 7098 4604 7104 4616
rect 6319 4576 7104 4604
rect 6319 4573 6331 4576
rect 6273 4567 6331 4573
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 7190 4564 7196 4616
rect 7248 4564 7254 4616
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 4062 4496 4068 4548
rect 4120 4496 4126 4548
rect 4706 4496 4712 4548
rect 4764 4496 4770 4548
rect 7392 4536 7420 4567
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 7650 4613 7656 4616
rect 7623 4607 7656 4613
rect 7623 4573 7635 4607
rect 7708 4604 7714 4616
rect 7708 4576 7972 4604
rect 7623 4567 7656 4573
rect 7650 4564 7656 4567
rect 7708 4564 7714 4576
rect 7742 4536 7748 4548
rect 7392 4508 7748 4536
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 7944 4536 7972 4576
rect 8018 4564 8024 4616
rect 8076 4564 8082 4616
rect 8128 4613 8156 4644
rect 8312 4644 8576 4672
rect 8312 4613 8340 4644
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11422 4672 11428 4684
rect 11112 4644 11428 4672
rect 11112 4632 11118 4644
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 9030 4604 9036 4616
rect 8527 4576 9036 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10873 4607 10931 4613
rect 10873 4604 10885 4607
rect 9732 4576 10885 4604
rect 9732 4564 9738 4576
rect 10873 4573 10885 4576
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 8202 4536 8208 4548
rect 7944 4508 8208 4536
rect 8202 4496 8208 4508
rect 8260 4536 8266 4548
rect 8389 4539 8447 4545
rect 8389 4536 8401 4539
rect 8260 4508 8401 4536
rect 8260 4496 8266 4508
rect 8389 4505 8401 4508
rect 8435 4505 8447 4539
rect 10888 4536 10916 4567
rect 11146 4564 11152 4616
rect 11204 4564 11210 4616
rect 11514 4564 11520 4616
rect 11572 4564 11578 4616
rect 11808 4613 11836 4780
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12860 4780 13001 4808
rect 12860 4768 12866 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 14366 4808 14372 4820
rect 12989 4771 13047 4777
rect 13372 4780 14372 4808
rect 11977 4743 12035 4749
rect 11977 4709 11989 4743
rect 12023 4740 12035 4743
rect 13372 4740 13400 4780
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15930 4808 15936 4820
rect 14660 4780 15936 4808
rect 12023 4712 13400 4740
rect 13449 4743 13507 4749
rect 12023 4709 12035 4712
rect 11977 4703 12035 4709
rect 13449 4709 13461 4743
rect 13495 4740 13507 4743
rect 13630 4740 13636 4752
rect 13495 4712 13636 4740
rect 13495 4709 13507 4712
rect 13449 4703 13507 4709
rect 13630 4700 13636 4712
rect 13688 4700 13694 4752
rect 14182 4672 14188 4684
rect 12268 4644 14188 4672
rect 12268 4613 12296 4644
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 11241 4539 11299 4545
rect 11241 4536 11253 4539
rect 10888 4508 11253 4536
rect 8389 4499 8447 4505
rect 11241 4505 11253 4508
rect 11287 4505 11299 4539
rect 11241 4499 11299 4505
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 12066 4536 12072 4548
rect 11388 4508 12072 4536
rect 11388 4496 11394 4508
rect 12066 4496 12072 4508
rect 12124 4496 12130 4548
rect 7834 4428 7840 4480
rect 7892 4428 7898 4480
rect 10689 4471 10747 4477
rect 10689 4437 10701 4471
rect 10735 4468 10747 4471
rect 10870 4468 10876 4480
rect 10735 4440 10876 4468
rect 10735 4437 10747 4440
rect 10689 4431 10747 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 11057 4471 11115 4477
rect 11057 4437 11069 4471
rect 11103 4468 11115 4471
rect 11146 4468 11152 4480
rect 11103 4440 11152 4468
rect 11103 4437 11115 4440
rect 11057 4431 11115 4437
rect 11146 4428 11152 4440
rect 11204 4468 11210 4480
rect 11425 4471 11483 4477
rect 11425 4468 11437 4471
rect 11204 4440 11437 4468
rect 11204 4428 11210 4440
rect 11425 4437 11437 4440
rect 11471 4468 11483 4471
rect 11882 4468 11888 4480
rect 11471 4440 11888 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 12158 4428 12164 4480
rect 12216 4428 12222 4480
rect 12360 4468 12388 4567
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12492 4576 12537 4604
rect 12492 4564 12498 4576
rect 12802 4564 12808 4616
rect 12860 4613 12866 4616
rect 12860 4567 12868 4613
rect 12860 4564 12866 4567
rect 13170 4564 13176 4616
rect 13228 4564 13234 4616
rect 13262 4564 13268 4616
rect 13320 4564 13326 4616
rect 13633 4607 13691 4613
rect 13633 4573 13645 4607
rect 13679 4604 13691 4607
rect 13722 4604 13728 4616
rect 13679 4576 13728 4604
rect 13679 4573 13691 4576
rect 13633 4567 13691 4573
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14458 4613 14464 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13964 4576 14289 4604
rect 13964 4564 13970 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14431 4607 14464 4613
rect 14431 4573 14443 4607
rect 14431 4567 14464 4573
rect 14458 4564 14464 4567
rect 14516 4564 14522 4616
rect 12618 4496 12624 4548
rect 12676 4496 12682 4548
rect 12713 4539 12771 4545
rect 12713 4505 12725 4539
rect 12759 4536 12771 4539
rect 13280 4536 13308 4564
rect 14660 4545 14688 4780
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 16025 4811 16083 4817
rect 16025 4777 16037 4811
rect 16071 4808 16083 4811
rect 16482 4808 16488 4820
rect 16071 4780 16488 4808
rect 16071 4777 16083 4780
rect 16025 4771 16083 4777
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 16942 4768 16948 4820
rect 17000 4808 17006 4820
rect 20714 4808 20720 4820
rect 17000 4780 20720 4808
rect 17000 4768 17006 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 21358 4768 21364 4820
rect 21416 4768 21422 4820
rect 14826 4700 14832 4752
rect 14884 4740 14890 4752
rect 16206 4740 16212 4752
rect 14884 4712 16212 4740
rect 14884 4700 14890 4712
rect 16206 4700 16212 4712
rect 16264 4700 16270 4752
rect 16390 4700 16396 4752
rect 16448 4740 16454 4752
rect 17589 4743 17647 4749
rect 17589 4740 17601 4743
rect 16448 4712 17601 4740
rect 16448 4700 16454 4712
rect 17589 4709 17601 4712
rect 17635 4740 17647 4743
rect 18506 4740 18512 4752
rect 17635 4712 18512 4740
rect 17635 4709 17647 4712
rect 17589 4703 17647 4709
rect 18506 4700 18512 4712
rect 18564 4700 18570 4752
rect 20533 4743 20591 4749
rect 20533 4709 20545 4743
rect 20579 4709 20591 4743
rect 20533 4703 20591 4709
rect 15562 4672 15568 4684
rect 15028 4644 15568 4672
rect 15028 4613 15056 4644
rect 15562 4632 15568 4644
rect 15620 4672 15626 4684
rect 20548 4672 20576 4703
rect 15620 4644 20576 4672
rect 15620 4632 15626 4644
rect 22278 4632 22284 4684
rect 22336 4672 22342 4684
rect 22336 4644 23060 4672
rect 22336 4632 22342 4644
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 16022 4604 16028 4616
rect 15335 4576 16028 4604
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 12759 4508 13308 4536
rect 13449 4539 13507 4545
rect 12759 4505 12771 4508
rect 12713 4499 12771 4505
rect 13449 4505 13461 4539
rect 13495 4536 13507 4539
rect 14645 4539 14703 4545
rect 14645 4536 14657 4539
rect 13495 4508 14657 4536
rect 13495 4505 13507 4508
rect 13449 4499 13507 4505
rect 14645 4505 14657 4508
rect 14691 4505 14703 4539
rect 14645 4499 14703 4505
rect 14918 4496 14924 4548
rect 14976 4496 14982 4548
rect 12986 4468 12992 4480
rect 12360 4440 12992 4468
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 13262 4428 13268 4480
rect 13320 4428 13326 4480
rect 13909 4471 13967 4477
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 14090 4468 14096 4480
rect 13955 4440 14096 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 15304 4468 15332 4567
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16206 4564 16212 4616
rect 16264 4564 16270 4616
rect 16298 4564 16304 4616
rect 16356 4604 16362 4616
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 16356 4576 16405 4604
rect 16356 4564 16362 4576
rect 16393 4573 16405 4576
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 16482 4564 16488 4616
rect 16540 4564 16546 4616
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 16632 4576 16957 4604
rect 16632 4564 16638 4576
rect 16945 4573 16957 4576
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 17034 4564 17040 4616
rect 17092 4564 17098 4616
rect 17218 4564 17224 4616
rect 17276 4564 17282 4616
rect 19061 4607 19119 4613
rect 19061 4573 19073 4607
rect 19107 4604 19119 4607
rect 20530 4604 20536 4616
rect 19107 4576 20536 4604
rect 19107 4573 19119 4576
rect 19061 4567 19119 4573
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 23032 4613 23060 4644
rect 22833 4607 22891 4613
rect 22833 4604 22845 4607
rect 22612 4576 22845 4604
rect 22612 4564 22618 4576
rect 22833 4573 22845 4576
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23106 4604 23112 4616
rect 23063 4576 23112 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 15749 4539 15807 4545
rect 15749 4505 15761 4539
rect 15795 4536 15807 4539
rect 16758 4536 16764 4548
rect 15795 4508 16764 4536
rect 15795 4505 15807 4508
rect 15749 4499 15807 4505
rect 16758 4496 16764 4508
rect 16816 4496 16822 4548
rect 19242 4496 19248 4548
rect 19300 4496 19306 4548
rect 14884 4440 15332 4468
rect 14884 4428 14890 4440
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 16577 4471 16635 4477
rect 16577 4468 16589 4471
rect 16356 4440 16589 4468
rect 16356 4428 16362 4440
rect 16577 4437 16589 4440
rect 16623 4468 16635 4471
rect 17126 4468 17132 4480
rect 16623 4440 17132 4468
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 17126 4428 17132 4440
rect 17184 4468 17190 4480
rect 17494 4468 17500 4480
rect 17184 4440 17500 4468
rect 17184 4428 17190 4440
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 23198 4428 23204 4480
rect 23256 4428 23262 4480
rect 1104 4378 23644 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 23644 4378
rect 1104 4304 23644 4326
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 4985 4267 5043 4273
rect 4985 4264 4997 4267
rect 4856 4236 4997 4264
rect 4856 4224 4862 4236
rect 4985 4233 4997 4236
rect 5031 4233 5043 4267
rect 4985 4227 5043 4233
rect 5537 4267 5595 4273
rect 5537 4233 5549 4267
rect 5583 4264 5595 4267
rect 6454 4264 6460 4276
rect 5583 4236 6460 4264
rect 5583 4233 5595 4236
rect 5537 4227 5595 4233
rect 4249 4199 4307 4205
rect 4249 4165 4261 4199
rect 4295 4196 4307 4199
rect 4614 4196 4620 4208
rect 4295 4168 4620 4196
rect 4295 4165 4307 4168
rect 4249 4159 4307 4165
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 5552 4196 5580 4227
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 8386 4264 8392 4276
rect 7800 4236 8392 4264
rect 7800 4224 7806 4236
rect 8386 4224 8392 4236
rect 8444 4264 8450 4276
rect 8665 4267 8723 4273
rect 8665 4264 8677 4267
rect 8444 4236 8677 4264
rect 8444 4224 8450 4236
rect 8665 4233 8677 4236
rect 8711 4233 8723 4267
rect 11717 4267 11775 4273
rect 11717 4264 11729 4267
rect 8665 4227 8723 4233
rect 10888 4236 11729 4264
rect 10888 4208 10916 4236
rect 11717 4233 11729 4236
rect 11763 4233 11775 4267
rect 11717 4227 11775 4233
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 12177 4267 12235 4273
rect 12177 4264 12189 4267
rect 12124 4236 12189 4264
rect 12124 4224 12130 4236
rect 12177 4233 12189 4236
rect 12223 4233 12235 4267
rect 12805 4267 12863 4273
rect 12805 4264 12817 4267
rect 12177 4227 12235 4233
rect 12469 4236 12817 4264
rect 4764 4168 5580 4196
rect 4764 4156 4770 4168
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4120 4100 5181 4128
rect 4120 4088 4126 4100
rect 5169 4097 5181 4100
rect 5215 4128 5227 4131
rect 5258 4128 5264 4140
rect 5215 4100 5264 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 5368 4137 5396 4168
rect 5626 4156 5632 4208
rect 5684 4156 5690 4208
rect 8849 4199 8907 4205
rect 8849 4196 8861 4199
rect 8128 4168 8861 4196
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 7524 4100 7573 4128
rect 7524 4088 7530 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 8128 4137 8156 4168
rect 8849 4165 8861 4168
rect 8895 4165 8907 4199
rect 8849 4159 8907 4165
rect 9030 4156 9036 4208
rect 9088 4196 9094 4208
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 9088 4168 9597 4196
rect 9088 4156 9094 4168
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 9585 4159 9643 4165
rect 10870 4156 10876 4208
rect 10928 4156 10934 4208
rect 11330 4196 11336 4208
rect 11072 4168 11336 4196
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 5276 3924 5304 4088
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4060 7711 4063
rect 8128 4060 8156 4091
rect 8202 4088 8208 4140
rect 8260 4088 8266 4140
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8343 4100 8432 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 7699 4032 8156 4060
rect 7699 4029 7711 4032
rect 7653 4023 7711 4029
rect 7929 3995 7987 4001
rect 7929 3961 7941 3995
rect 7975 3992 7987 3995
rect 8294 3992 8300 4004
rect 7975 3964 8300 3992
rect 7975 3961 7987 3964
rect 7929 3955 7987 3961
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 8404 3992 8432 4100
rect 8478 4088 8484 4140
rect 8536 4088 8542 4140
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 8588 4060 8616 4091
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8812 4100 9137 4128
rect 8812 4088 8818 4100
rect 9125 4097 9137 4100
rect 9171 4128 9183 4131
rect 9214 4128 9220 4140
rect 9171 4100 9220 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9324 4060 9352 4091
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9456 4100 9505 4128
rect 9456 4088 9462 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 9674 4088 9680 4140
rect 9732 4088 9738 4140
rect 11072 4137 11100 4168
rect 11330 4156 11336 4168
rect 11388 4156 11394 4208
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 11977 4199 12035 4205
rect 11977 4196 11989 4199
rect 11572 4168 11989 4196
rect 11572 4156 11578 4168
rect 11977 4165 11989 4168
rect 12023 4165 12035 4199
rect 11977 4159 12035 4165
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4097 11207 4131
rect 12469 4128 12497 4236
rect 12805 4233 12817 4236
rect 12851 4264 12863 4267
rect 13262 4264 13268 4276
rect 12851 4236 13268 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 15010 4264 15016 4276
rect 14240 4236 15016 4264
rect 14240 4224 14246 4236
rect 15010 4224 15016 4236
rect 15068 4224 15074 4276
rect 15197 4267 15255 4273
rect 15197 4233 15209 4267
rect 15243 4264 15255 4267
rect 15286 4264 15292 4276
rect 15243 4236 15292 4264
rect 15243 4233 15255 4236
rect 15197 4227 15255 4233
rect 15286 4224 15292 4236
rect 15344 4264 15350 4276
rect 17034 4264 17040 4276
rect 15344 4236 17040 4264
rect 15344 4224 15350 4236
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 21358 4264 21364 4276
rect 20824 4236 21364 4264
rect 12989 4199 13047 4205
rect 12989 4165 13001 4199
rect 13035 4196 13047 4199
rect 14829 4199 14887 4205
rect 14829 4196 14841 4199
rect 13035 4168 14841 4196
rect 13035 4165 13047 4168
rect 12989 4159 13047 4165
rect 14829 4165 14841 4168
rect 14875 4196 14887 4199
rect 15654 4196 15660 4208
rect 14875 4168 15660 4196
rect 14875 4165 14887 4168
rect 14829 4159 14887 4165
rect 15654 4156 15660 4168
rect 15712 4196 15718 4208
rect 15712 4168 16160 4196
rect 15712 4156 15718 4168
rect 11149 4091 11207 4097
rect 11732 4100 12497 4128
rect 12713 4131 12771 4137
rect 9692 4060 9720 4088
rect 8588 4032 9168 4060
rect 9324 4032 9720 4060
rect 8570 3992 8576 4004
rect 8404 3964 8576 3992
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 9140 4001 9168 4032
rect 9125 3995 9183 4001
rect 9125 3961 9137 3995
rect 9171 3961 9183 3995
rect 9125 3955 9183 3961
rect 9030 3924 9036 3936
rect 5276 3896 9036 3924
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9140 3924 9168 3955
rect 9306 3952 9312 4004
rect 9364 3992 9370 4004
rect 11164 3992 11192 4091
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 11732 4060 11760 4100
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13446 4128 13452 4140
rect 13403 4100 13452 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 12250 4060 12256 4072
rect 11388 4032 11760 4060
rect 11808 4032 12256 4060
rect 11388 4020 11394 4032
rect 11514 3992 11520 4004
rect 9364 3964 11520 3992
rect 9364 3952 9370 3964
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 11808 3992 11836 4032
rect 12250 4020 12256 4032
rect 12308 4060 12314 4072
rect 12728 4060 12756 4091
rect 13280 4060 13308 4091
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 13630 4088 13636 4140
rect 13688 4088 13694 4140
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13872 4100 14013 4128
rect 13872 4088 13878 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 14458 4128 14464 4140
rect 14240 4100 14464 4128
rect 14240 4088 14246 4100
rect 14458 4088 14464 4100
rect 14516 4128 14522 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14516 4100 14657 4128
rect 14516 4088 14522 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14844 4100 15608 4128
rect 12308 4032 12756 4060
rect 12912 4032 13308 4060
rect 12308 4020 12314 4032
rect 11624 3964 11836 3992
rect 10410 3924 10416 3936
rect 9140 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3924 10474 3936
rect 10873 3927 10931 3933
rect 10873 3924 10885 3927
rect 10468 3896 10885 3924
rect 10468 3884 10474 3896
rect 10873 3893 10885 3896
rect 10919 3893 10931 3927
rect 10873 3887 10931 3893
rect 11330 3884 11336 3936
rect 11388 3884 11394 3936
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11624 3924 11652 3964
rect 11882 3952 11888 4004
rect 11940 3952 11946 4004
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 12912 3992 12940 4032
rect 12676 3964 12940 3992
rect 12676 3952 12682 3964
rect 12986 3952 12992 4004
rect 13044 3952 13050 4004
rect 13170 3952 13176 4004
rect 13228 3992 13234 4004
rect 14369 3995 14427 4001
rect 14369 3992 14381 3995
rect 13228 3964 14381 3992
rect 13228 3952 13234 3964
rect 14369 3961 14381 3964
rect 14415 3992 14427 3995
rect 14844 3992 14872 4100
rect 15580 4072 15608 4100
rect 15838 4088 15844 4140
rect 15896 4088 15902 4140
rect 16132 4137 16160 4168
rect 16206 4156 16212 4208
rect 16264 4196 16270 4208
rect 19702 4196 19708 4208
rect 16264 4168 19708 4196
rect 16264 4156 16270 4168
rect 19702 4156 19708 4168
rect 19760 4156 19766 4208
rect 20824 4205 20852 4236
rect 21358 4224 21364 4236
rect 21416 4224 21422 4276
rect 20809 4199 20867 4205
rect 20809 4165 20821 4199
rect 20855 4165 20867 4199
rect 22278 4196 22284 4208
rect 20809 4159 20867 4165
rect 20916 4168 22284 4196
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4097 16543 4131
rect 16485 4091 16543 4097
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 16758 4128 16764 4140
rect 16715 4100 16764 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4029 14979 4063
rect 15470 4060 15476 4072
rect 14921 4023 14979 4029
rect 15304 4032 15476 4060
rect 14415 3964 14872 3992
rect 14415 3961 14427 3964
rect 14369 3955 14427 3961
rect 11480 3896 11652 3924
rect 11701 3927 11759 3933
rect 11480 3884 11486 3896
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 11974 3924 11980 3936
rect 11747 3896 11980 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 11974 3884 11980 3896
rect 12032 3924 12038 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 12032 3896 12173 3924
rect 12032 3884 12038 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12308 3896 12357 3924
rect 12308 3884 12314 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12584 3896 13093 3924
rect 12584 3884 12590 3896
rect 13081 3893 13093 3896
rect 13127 3893 13139 3927
rect 13081 3887 13139 3893
rect 14458 3884 14464 3936
rect 14516 3884 14522 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 14936 3924 14964 4023
rect 15304 4004 15332 4032
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15620 4032 15669 4060
rect 15620 4020 15626 4032
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 16022 4020 16028 4072
rect 16080 4020 16086 4072
rect 16206 4020 16212 4072
rect 16264 4020 16270 4072
rect 16301 4063 16359 4069
rect 16301 4029 16313 4063
rect 16347 4060 16359 4063
rect 16390 4060 16396 4072
rect 16347 4032 16396 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16500 4060 16528 4091
rect 16758 4088 16764 4100
rect 16816 4128 16822 4140
rect 17218 4128 17224 4140
rect 16816 4100 17224 4128
rect 16816 4088 16822 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17310 4088 17316 4140
rect 17368 4128 17374 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17368 4100 17785 4128
rect 17368 4088 17374 4100
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17773 4091 17831 4097
rect 17880 4100 18337 4128
rect 17126 4060 17132 4072
rect 16500 4032 17132 4060
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17880 4060 17908 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 20916 4137 20944 4168
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 22370 4156 22376 4208
rect 22428 4196 22434 4208
rect 22428 4168 23152 4196
rect 22428 4156 22434 4168
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 19208 4100 20453 4128
rect 19208 4088 19214 4100
rect 20441 4097 20453 4100
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4128 20591 4131
rect 20901 4131 20959 4137
rect 20579 4100 20852 4128
rect 20579 4097 20591 4100
rect 20533 4091 20591 4097
rect 20824 4072 20852 4100
rect 20901 4097 20913 4131
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4097 21051 4131
rect 20993 4091 21051 4097
rect 17451 4032 17908 4060
rect 18049 4063 18107 4069
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18141 4063 18199 4069
rect 18141 4029 18153 4063
rect 18187 4060 18199 4063
rect 18414 4060 18420 4072
rect 18187 4032 18420 4060
rect 18187 4029 18199 4032
rect 18141 4023 18199 4029
rect 15286 3952 15292 4004
rect 15344 3952 15350 4004
rect 15378 3952 15384 4004
rect 15436 3992 15442 4004
rect 18064 3992 18092 4023
rect 18414 4020 18420 4032
rect 18472 4020 18478 4072
rect 18506 4020 18512 4072
rect 18564 4060 18570 4072
rect 18564 4032 20484 4060
rect 18564 4020 18570 4032
rect 15436 3964 18092 3992
rect 15436 3952 15442 3964
rect 19610 3952 19616 4004
rect 19668 3952 19674 4004
rect 15930 3924 15936 3936
rect 14700 3896 15936 3924
rect 14700 3884 14706 3896
rect 15930 3884 15936 3896
rect 15988 3924 15994 3936
rect 16114 3924 16120 3936
rect 15988 3896 16120 3924
rect 15988 3884 15994 3896
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 20254 3884 20260 3936
rect 20312 3884 20318 3936
rect 20456 3924 20484 4032
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 20680 4032 20729 4060
rect 20680 4020 20686 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 20806 4020 20812 4072
rect 20864 4020 20870 4072
rect 21008 4060 21036 4091
rect 21174 4088 21180 4140
rect 21232 4088 21238 4140
rect 21269 4131 21327 4137
rect 21269 4097 21281 4131
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 20916 4032 21036 4060
rect 20530 3952 20536 4004
rect 20588 3992 20594 4004
rect 20916 3992 20944 4032
rect 20588 3964 20944 3992
rect 20588 3952 20594 3964
rect 21284 3924 21312 4091
rect 21358 4088 21364 4140
rect 21416 4137 21422 4140
rect 21416 4128 21424 4137
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 21416 4100 21461 4128
rect 22066 4100 22477 4128
rect 21416 4091 21424 4100
rect 21416 4088 21422 4091
rect 21545 3995 21603 4001
rect 21545 3961 21557 3995
rect 21591 3992 21603 3995
rect 22066 3992 22094 4100
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 22646 4088 22652 4140
rect 22704 4088 22710 4140
rect 22830 4088 22836 4140
rect 22888 4088 22894 4140
rect 23124 4137 23152 4168
rect 23109 4131 23167 4137
rect 23109 4097 23121 4131
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 23201 4063 23259 4069
rect 23201 4060 23213 4063
rect 22244 4032 23213 4060
rect 22244 4020 22250 4032
rect 23201 4029 23213 4032
rect 23247 4029 23259 4063
rect 23201 4023 23259 4029
rect 21591 3964 22094 3992
rect 21591 3961 21603 3964
rect 21545 3955 21603 3961
rect 22278 3952 22284 4004
rect 22336 3952 22342 4004
rect 20456 3896 21312 3924
rect 1104 3834 23644 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 23644 3834
rect 1104 3760 23644 3782
rect 7377 3723 7435 3729
rect 7377 3689 7389 3723
rect 7423 3720 7435 3723
rect 8018 3720 8024 3732
rect 7423 3692 8024 3720
rect 7423 3689 7435 3692
rect 7377 3683 7435 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8757 3723 8815 3729
rect 8757 3689 8769 3723
rect 8803 3720 8815 3723
rect 10042 3720 10048 3732
rect 8803 3692 10048 3720
rect 8803 3689 8815 3692
rect 8757 3683 8815 3689
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10226 3680 10232 3732
rect 10284 3680 10290 3732
rect 10597 3723 10655 3729
rect 10597 3689 10609 3723
rect 10643 3689 10655 3723
rect 10597 3683 10655 3689
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 7929 3655 7987 3661
rect 7248 3624 7880 3652
rect 7248 3612 7254 3624
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 7852 3584 7880 3624
rect 7929 3621 7941 3655
rect 7975 3652 7987 3655
rect 7975 3624 10548 3652
rect 7975 3621 7987 3624
rect 7929 3615 7987 3621
rect 8297 3587 8355 3593
rect 7432 3556 7788 3584
rect 7852 3556 8248 3584
rect 7432 3544 7438 3556
rect 7760 3525 7788 3556
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 7147 3488 7481 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7469 3485 7481 3488
rect 7515 3516 7527 3519
rect 7745 3519 7803 3525
rect 7515 3488 7696 3516
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 7374 3408 7380 3460
rect 7432 3408 7438 3460
rect 7668 3392 7696 3488
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 8110 3516 8116 3528
rect 7791 3488 8116 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8220 3525 8248 3556
rect 8297 3553 8309 3587
rect 8343 3584 8355 3587
rect 9033 3587 9091 3593
rect 9033 3584 9045 3587
rect 8343 3556 9045 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 9033 3553 9045 3556
rect 9079 3584 9091 3587
rect 9493 3587 9551 3593
rect 9079 3556 9444 3584
rect 9079 3553 9091 3556
rect 9033 3547 9091 3553
rect 9416 3528 9444 3556
rect 9493 3553 9505 3587
rect 9539 3584 9551 3587
rect 10318 3584 10324 3596
rect 9539 3556 10324 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8478 3476 8484 3528
rect 8536 3476 8542 3528
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 8588 3448 8616 3479
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8938 3516 8944 3528
rect 8720 3488 8944 3516
rect 8720 3476 8726 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9214 3476 9220 3528
rect 9272 3476 9278 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9324 3448 9352 3479
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9585 3519 9643 3525
rect 9585 3516 9597 3519
rect 9456 3488 9597 3516
rect 9456 3476 9462 3488
rect 9585 3485 9597 3488
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 9858 3476 9864 3528
rect 9916 3476 9922 3528
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 10060 3488 10149 3516
rect 10060 3448 10088 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10520 3516 10548 3624
rect 10612 3584 10640 3683
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11146 3720 11152 3732
rect 10928 3692 11152 3720
rect 10928 3680 10934 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11422 3680 11428 3732
rect 11480 3680 11486 3732
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 11701 3723 11759 3729
rect 11701 3720 11713 3723
rect 11664 3692 11713 3720
rect 11664 3680 11670 3692
rect 11701 3689 11713 3692
rect 11747 3689 11759 3723
rect 11977 3723 12035 3729
rect 11977 3720 11989 3723
rect 11701 3683 11759 3689
rect 11808 3692 11989 3720
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 11808 3652 11836 3692
rect 11977 3689 11989 3692
rect 12023 3689 12035 3723
rect 11977 3683 12035 3689
rect 12345 3723 12403 3729
rect 12345 3689 12357 3723
rect 12391 3720 12403 3723
rect 12618 3720 12624 3732
rect 12391 3692 12624 3720
rect 12391 3689 12403 3692
rect 12345 3683 12403 3689
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 12986 3720 12992 3732
rect 12820 3692 12992 3720
rect 10827 3624 11836 3652
rect 11885 3655 11943 3661
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 11716 3596 11744 3624
rect 11885 3621 11897 3655
rect 11931 3621 11943 3655
rect 12820 3652 12848 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13078 3680 13084 3732
rect 13136 3680 13142 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13596 3692 13737 3720
rect 13596 3680 13602 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 20070 3720 20076 3732
rect 13872 3692 14596 3720
rect 13872 3680 13878 3692
rect 13096 3652 13124 3680
rect 11885 3615 11943 3621
rect 12636 3624 12848 3652
rect 12912 3624 14412 3652
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10612 3556 10977 3584
rect 10965 3553 10977 3556
rect 11011 3584 11023 3587
rect 11606 3584 11612 3596
rect 11011 3556 11612 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11698 3544 11704 3596
rect 11756 3544 11762 3596
rect 11900 3584 11928 3615
rect 12636 3584 12664 3624
rect 11900 3556 12664 3584
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10520 3488 10885 3516
rect 10137 3479 10195 3485
rect 10873 3485 10885 3488
rect 10919 3516 10931 3519
rect 11054 3516 11060 3528
rect 10919 3488 11060 3516
rect 10919 3485 10931 3488
rect 10873 3479 10931 3485
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11146 3476 11152 3528
rect 11204 3476 11210 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11296 3488 11652 3516
rect 11296 3476 11302 3488
rect 8496 3420 9352 3448
rect 9692 3420 10088 3448
rect 7193 3383 7251 3389
rect 7193 3349 7205 3383
rect 7239 3380 7251 3383
rect 7466 3380 7472 3392
rect 7239 3352 7472 3380
rect 7239 3349 7251 3352
rect 7193 3343 7251 3349
rect 7466 3340 7472 3352
rect 7524 3380 7530 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 7524 3352 7573 3380
rect 7524 3340 7530 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 8496 3380 8524 3420
rect 9692 3392 9720 3420
rect 10410 3408 10416 3460
rect 10468 3408 10474 3460
rect 10629 3451 10687 3457
rect 10629 3417 10641 3451
rect 10675 3448 10687 3451
rect 11256 3448 11284 3476
rect 10675 3420 11284 3448
rect 10675 3417 10687 3420
rect 10629 3411 10687 3417
rect 11514 3408 11520 3460
rect 11572 3408 11578 3460
rect 11624 3448 11652 3488
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11940 3488 11989 3516
rect 11940 3476 11946 3488
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3516 12127 3519
rect 12250 3516 12256 3528
rect 12115 3488 12256 3516
rect 12115 3485 12127 3488
rect 12069 3479 12127 3485
rect 12250 3476 12256 3488
rect 12308 3476 12314 3528
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12400 3488 12449 3516
rect 12400 3476 12406 3488
rect 12437 3485 12449 3488
rect 12483 3516 12495 3519
rect 12526 3516 12532 3528
rect 12483 3488 12532 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12636 3525 12664 3556
rect 12912 3525 12940 3624
rect 13078 3544 13084 3596
rect 13136 3584 13142 3596
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 13136 3556 13369 3584
rect 13136 3544 13142 3556
rect 13357 3553 13369 3556
rect 13403 3553 13415 3587
rect 13357 3547 13415 3553
rect 13446 3544 13452 3596
rect 13504 3544 13510 3596
rect 12621 3519 12679 3525
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13044 3488 13277 3516
rect 13044 3476 13050 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14384 3525 14412 3624
rect 14568 3593 14596 3692
rect 14660 3692 20076 3720
rect 14660 3661 14688 3692
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 20533 3723 20591 3729
rect 20533 3720 20545 3723
rect 20220 3692 20545 3720
rect 20220 3680 20226 3692
rect 20533 3689 20545 3692
rect 20579 3689 20591 3723
rect 20533 3683 20591 3689
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 21818 3720 21824 3732
rect 20956 3692 21824 3720
rect 20956 3680 20962 3692
rect 21818 3680 21824 3692
rect 21876 3680 21882 3732
rect 14645 3655 14703 3661
rect 14645 3621 14657 3655
rect 14691 3621 14703 3655
rect 14645 3615 14703 3621
rect 14826 3612 14832 3664
rect 14884 3652 14890 3664
rect 15105 3655 15163 3661
rect 15105 3652 15117 3655
rect 14884 3624 15117 3652
rect 14884 3612 14890 3624
rect 15105 3621 15117 3624
rect 15151 3621 15163 3655
rect 15105 3615 15163 3621
rect 15194 3612 15200 3664
rect 15252 3652 15258 3664
rect 15562 3652 15568 3664
rect 15252 3624 15568 3652
rect 15252 3612 15258 3624
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 16482 3612 16488 3664
rect 16540 3652 16546 3664
rect 17129 3655 17187 3661
rect 17129 3652 17141 3655
rect 16540 3624 17141 3652
rect 16540 3612 16546 3624
rect 17129 3621 17141 3624
rect 17175 3621 17187 3655
rect 17129 3615 17187 3621
rect 17218 3612 17224 3664
rect 17276 3652 17282 3664
rect 22373 3655 22431 3661
rect 22373 3652 22385 3655
rect 17276 3624 22385 3652
rect 17276 3612 17282 3624
rect 22373 3621 22385 3624
rect 22419 3621 22431 3655
rect 22373 3615 22431 3621
rect 14553 3587 14611 3593
rect 14553 3553 14565 3587
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 15068 3556 17325 3584
rect 15068 3544 15074 3556
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13596 3488 14105 3516
rect 13596 3476 13602 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 14185 3519 14243 3525
rect 14185 3485 14197 3519
rect 14231 3485 14243 3519
rect 14185 3479 14243 3485
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 14642 3516 14648 3528
rect 14415 3488 14648 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 11717 3451 11775 3457
rect 11717 3448 11729 3451
rect 11624 3420 11729 3448
rect 11717 3417 11729 3420
rect 11763 3417 11775 3451
rect 11717 3411 11775 3417
rect 12158 3408 12164 3460
rect 12216 3448 12222 3460
rect 14200 3448 14228 3479
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 14921 3519 14979 3525
rect 14921 3485 14933 3519
rect 14967 3516 14979 3519
rect 15194 3516 15200 3528
rect 14967 3488 15200 3516
rect 14967 3485 14979 3488
rect 14921 3479 14979 3485
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15286 3476 15292 3528
rect 15344 3476 15350 3528
rect 15470 3476 15476 3528
rect 15528 3476 15534 3528
rect 16025 3519 16083 3525
rect 16025 3485 16037 3519
rect 16071 3516 16083 3519
rect 16298 3516 16304 3528
rect 16071 3488 16304 3516
rect 16071 3485 16083 3488
rect 16025 3479 16083 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16482 3476 16488 3528
rect 16540 3476 16546 3528
rect 16684 3525 16712 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 17828 3556 20024 3584
rect 17828 3544 17834 3556
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 16758 3476 16764 3528
rect 16816 3476 16822 3528
rect 16854 3519 16912 3525
rect 16854 3485 16866 3519
rect 16900 3516 16912 3519
rect 16942 3516 16948 3528
rect 16900 3488 16948 3516
rect 16900 3485 16912 3488
rect 16854 3479 16912 3485
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 18966 3476 18972 3528
rect 19024 3476 19030 3528
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3516 19303 3519
rect 19334 3516 19340 3528
rect 19291 3488 19340 3516
rect 19291 3485 19303 3488
rect 19245 3479 19303 3485
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19996 3516 20024 3556
rect 20070 3544 20076 3596
rect 20128 3584 20134 3596
rect 21174 3584 21180 3596
rect 20128 3556 21180 3584
rect 20128 3544 20134 3556
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 21358 3516 21364 3528
rect 19996 3488 21364 3516
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 22388 3516 22416 3615
rect 22925 3519 22983 3525
rect 22925 3516 22937 3519
rect 22388 3488 22937 3516
rect 22925 3485 22937 3488
rect 22971 3485 22983 3519
rect 22925 3479 22983 3485
rect 23106 3476 23112 3528
rect 23164 3476 23170 3528
rect 16209 3451 16267 3457
rect 16209 3448 16221 3451
rect 12216 3420 14228 3448
rect 14384 3420 16221 3448
rect 12216 3408 12222 3420
rect 7708 3352 8524 3380
rect 7708 3340 7714 3352
rect 9674 3340 9680 3392
rect 9732 3340 9738 3392
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3380 10103 3383
rect 11146 3380 11152 3392
rect 10091 3352 11152 3380
rect 10091 3349 10103 3352
rect 10045 3343 10103 3349
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 12342 3380 12348 3392
rect 11664 3352 12348 3380
rect 11664 3340 11670 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 12986 3380 12992 3392
rect 12768 3352 12992 3380
rect 12768 3340 12774 3352
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13081 3383 13139 3389
rect 13081 3349 13093 3383
rect 13127 3380 13139 3383
rect 13814 3380 13820 3392
rect 13127 3352 13820 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 14274 3380 14280 3392
rect 13964 3352 14280 3380
rect 13964 3340 13970 3352
rect 14274 3340 14280 3352
rect 14332 3380 14338 3392
rect 14384 3380 14412 3420
rect 16209 3417 16221 3420
rect 16255 3448 16267 3451
rect 17034 3448 17040 3460
rect 16255 3420 17040 3448
rect 16255 3417 16267 3420
rect 16209 3411 16267 3417
rect 17034 3408 17040 3420
rect 17092 3408 17098 3460
rect 19886 3408 19892 3460
rect 19944 3448 19950 3460
rect 21085 3451 21143 3457
rect 21085 3448 21097 3451
rect 19944 3420 21097 3448
rect 19944 3408 19950 3420
rect 21085 3417 21097 3420
rect 21131 3417 21143 3451
rect 21085 3411 21143 3417
rect 14332 3352 14412 3380
rect 14332 3340 14338 3352
rect 14458 3340 14464 3392
rect 14516 3340 14522 3392
rect 14734 3340 14740 3392
rect 14792 3380 14798 3392
rect 15657 3383 15715 3389
rect 15657 3380 15669 3383
rect 14792 3352 15669 3380
rect 14792 3340 14798 3352
rect 15657 3349 15669 3352
rect 15703 3349 15715 3383
rect 15657 3343 15715 3349
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 17586 3380 17592 3392
rect 16172 3352 17592 3380
rect 16172 3340 16178 3352
rect 17586 3340 17592 3352
rect 17644 3380 17650 3392
rect 18966 3380 18972 3392
rect 17644 3352 18972 3380
rect 17644 3340 17650 3352
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 20530 3380 20536 3392
rect 19576 3352 20536 3380
rect 19576 3340 19582 3352
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 23017 3383 23075 3389
rect 23017 3380 23029 3383
rect 20772 3352 23029 3380
rect 20772 3340 20778 3352
rect 23017 3349 23029 3352
rect 23063 3349 23075 3383
rect 23017 3343 23075 3349
rect 1104 3290 23644 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 23644 3290
rect 1104 3216 23644 3238
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 6822 3176 6828 3188
rect 6687 3148 6828 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 6822 3136 6828 3148
rect 6880 3176 6886 3188
rect 7006 3176 7012 3188
rect 6880 3148 7012 3176
rect 6880 3136 6886 3148
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7558 3176 7564 3188
rect 7432 3148 7564 3176
rect 7432 3136 7438 3148
rect 7558 3136 7564 3148
rect 7616 3176 7622 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7616 3148 7849 3176
rect 7616 3136 7622 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 9674 3176 9680 3188
rect 9263 3148 9680 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10042 3176 10048 3188
rect 9784 3148 10048 3176
rect 7650 3068 7656 3120
rect 7708 3068 7714 3120
rect 9398 3068 9404 3120
rect 9456 3068 9462 3120
rect 9784 3108 9812 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10505 3179 10563 3185
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 10686 3176 10692 3188
rect 10551 3148 10692 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 12158 3136 12164 3188
rect 12216 3136 12222 3188
rect 12250 3136 12256 3188
rect 12308 3136 12314 3188
rect 12529 3179 12587 3185
rect 12529 3145 12541 3179
rect 12575 3176 12587 3179
rect 12618 3176 12624 3188
rect 12575 3148 12624 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12713 3179 12771 3185
rect 12713 3145 12725 3179
rect 12759 3176 12771 3179
rect 12802 3176 12808 3188
rect 12759 3148 12808 3176
rect 12759 3145 12771 3148
rect 12713 3139 12771 3145
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 13262 3136 13268 3188
rect 13320 3136 13326 3188
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 14458 3176 14464 3188
rect 14139 3148 14464 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3176 15255 3179
rect 15378 3176 15384 3188
rect 15243 3148 15384 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 10888 3108 10916 3136
rect 9646 3080 9812 3108
rect 9968 3080 10916 3108
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 6840 2972 6868 3003
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7282 3040 7288 3052
rect 7239 3012 7288 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 8018 3000 8024 3052
rect 8076 3000 8082 3052
rect 8386 3000 8392 3052
rect 8444 3000 8450 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8496 3012 8677 3040
rect 8110 2972 8116 2984
rect 6840 2944 8116 2972
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 8496 2972 8524 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8904 3012 9045 3040
rect 8904 3000 8910 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 8260 2944 8524 2972
rect 8260 2932 8266 2944
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 9646 2972 9674 3080
rect 9968 3052 9996 3080
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 12268 3108 12296 3136
rect 13538 3108 13544 3120
rect 11296 3080 11376 3108
rect 11296 3068 11302 3080
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 8628 2944 9674 2972
rect 9784 2972 9812 3003
rect 9950 3000 9956 3052
rect 10008 3000 10014 3052
rect 10042 3000 10048 3052
rect 10100 3000 10106 3052
rect 10318 3000 10324 3052
rect 10376 3000 10382 3052
rect 10778 3000 10784 3052
rect 10836 3000 10842 3052
rect 10870 3000 10876 3052
rect 10928 3000 10934 3052
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11348 3049 11376 3080
rect 11532 3080 12296 3108
rect 12912 3080 13544 3108
rect 11532 3049 11560 3080
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 11112 3012 11161 3040
rect 11112 3000 11118 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3009 11391 3043
rect 11333 3003 11391 3009
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12250 3040 12256 3052
rect 12023 3012 12256 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 10594 2972 10600 2984
rect 9784 2944 10600 2972
rect 8628 2932 8634 2944
rect 7006 2864 7012 2916
rect 7064 2904 7070 2916
rect 9784 2904 9812 2944
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2972 10747 2975
rect 10962 2972 10968 2984
rect 10735 2944 10968 2972
rect 10735 2941 10747 2944
rect 10689 2935 10747 2941
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11882 2972 11888 2984
rect 11287 2944 11888 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 11992 2904 12020 3003
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 12492 3012 12633 3040
rect 12492 3000 12498 3012
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 12621 3003 12679 3009
rect 12710 3000 12716 3052
rect 12768 3040 12774 3052
rect 12912 3049 12940 3080
rect 13538 3068 13544 3080
rect 13596 3068 13602 3120
rect 15212 3108 15240 3139
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 16758 3136 16764 3188
rect 16816 3136 16822 3188
rect 17957 3179 18015 3185
rect 17957 3145 17969 3179
rect 18003 3176 18015 3179
rect 18414 3176 18420 3188
rect 18003 3148 18420 3176
rect 18003 3145 18015 3148
rect 17957 3139 18015 3145
rect 18414 3136 18420 3148
rect 18472 3176 18478 3188
rect 19242 3176 19248 3188
rect 18472 3148 19248 3176
rect 18472 3136 18478 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 22002 3176 22008 3188
rect 21652 3148 22008 3176
rect 13648 3080 15240 3108
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 12768 3012 12909 3040
rect 12768 3000 12774 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13078 3000 13084 3052
rect 13136 3000 13142 3052
rect 13446 3000 13452 3052
rect 13504 3000 13510 3052
rect 13648 3049 13676 3080
rect 15470 3068 15476 3120
rect 15528 3108 15534 3120
rect 15528 3080 16620 3108
rect 15528 3068 15534 3080
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13814 3000 13820 3052
rect 13872 3000 13878 3052
rect 13998 3000 14004 3052
rect 14056 3000 14062 3052
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 16485 3043 16543 3049
rect 16485 3009 16497 3043
rect 16531 3009 16543 3043
rect 16592 3040 16620 3080
rect 18966 3068 18972 3120
rect 19024 3108 19030 3120
rect 19337 3111 19395 3117
rect 19337 3108 19349 3111
rect 19024 3080 19349 3108
rect 19024 3068 19030 3080
rect 19337 3077 19349 3080
rect 19383 3077 19395 3111
rect 19337 3071 19395 3077
rect 19521 3111 19579 3117
rect 19521 3077 19533 3111
rect 19567 3077 19579 3111
rect 19521 3071 19579 3077
rect 19889 3111 19947 3117
rect 19889 3077 19901 3111
rect 19935 3108 19947 3111
rect 19978 3108 19984 3120
rect 19935 3080 19984 3108
rect 19935 3077 19947 3080
rect 19889 3071 19947 3077
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16592 3012 16681 3040
rect 16485 3003 16543 3009
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 12124 2944 13737 2972
rect 12124 2932 12130 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13725 2935 13783 2941
rect 13832 2944 14197 2972
rect 7064 2876 9812 2904
rect 10704 2876 12020 2904
rect 7064 2864 7070 2876
rect 750 2796 756 2848
rect 808 2836 814 2848
rect 1397 2839 1455 2845
rect 1397 2836 1409 2839
rect 808 2808 1409 2836
rect 808 2796 814 2808
rect 1397 2805 1409 2808
rect 1443 2805 1455 2839
rect 1397 2799 1455 2805
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 7340 2808 8217 2836
rect 7340 2796 7346 2808
rect 8205 2805 8217 2808
rect 8251 2836 8263 2839
rect 8846 2836 8852 2848
rect 8251 2808 8852 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 9048 2845 9076 2876
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2805 9091 2839
rect 9033 2799 9091 2805
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 10704 2836 10732 2876
rect 9180 2808 10732 2836
rect 9180 2796 9186 2808
rect 10778 2796 10784 2848
rect 10836 2836 10842 2848
rect 10962 2836 10968 2848
rect 10836 2808 10968 2836
rect 10836 2796 10842 2808
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11057 2839 11115 2845
rect 11057 2805 11069 2839
rect 11103 2836 11115 2839
rect 11238 2836 11244 2848
rect 11103 2808 11244 2836
rect 11103 2805 11115 2808
rect 11057 2799 11115 2805
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 12158 2836 12164 2848
rect 11388 2808 12164 2836
rect 11388 2796 11394 2808
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 12526 2796 12532 2848
rect 12584 2836 12590 2848
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12584 2808 12909 2836
rect 12584 2796 12590 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 12897 2799 12955 2805
rect 12986 2796 12992 2848
rect 13044 2836 13050 2848
rect 13722 2836 13728 2848
rect 13044 2808 13728 2836
rect 13044 2796 13050 2808
rect 13722 2796 13728 2808
rect 13780 2836 13786 2848
rect 13832 2836 13860 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14277 2907 14335 2913
rect 14277 2873 14289 2907
rect 14323 2904 14335 2907
rect 16500 2904 16528 3003
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 19242 3000 19248 3052
rect 19300 3000 19306 3052
rect 17126 2932 17132 2984
rect 17184 2932 17190 2984
rect 18506 2932 18512 2984
rect 18564 2972 18570 2984
rect 19536 2972 19564 3071
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 21652 3117 21680 3148
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22281 3179 22339 3185
rect 22281 3145 22293 3179
rect 22327 3176 22339 3179
rect 22830 3176 22836 3188
rect 22327 3148 22836 3176
rect 22327 3145 22339 3148
rect 22281 3139 22339 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 23014 3136 23020 3188
rect 23072 3176 23078 3188
rect 23201 3179 23259 3185
rect 23201 3176 23213 3179
rect 23072 3148 23213 3176
rect 23072 3136 23078 3148
rect 23201 3145 23213 3148
rect 23247 3145 23259 3179
rect 23201 3139 23259 3145
rect 21637 3111 21695 3117
rect 21637 3077 21649 3111
rect 21683 3077 21695 3111
rect 21637 3071 21695 3077
rect 21818 3068 21824 3120
rect 21876 3108 21882 3120
rect 23382 3108 23388 3120
rect 21876 3080 22600 3108
rect 21876 3068 21882 3080
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 20680 3012 22017 3040
rect 20680 3000 20686 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 22370 3000 22376 3052
rect 22428 3000 22434 3052
rect 22572 3049 22600 3080
rect 22756 3080 23388 3108
rect 22756 3049 22784 3080
rect 23382 3068 23388 3080
rect 23440 3068 23446 3120
rect 22557 3043 22615 3049
rect 22557 3009 22569 3043
rect 22603 3009 22615 3043
rect 22557 3003 22615 3009
rect 22741 3043 22799 3049
rect 22741 3009 22753 3043
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 23017 3043 23075 3049
rect 23017 3009 23029 3043
rect 23063 3009 23075 3043
rect 23017 3003 23075 3009
rect 18564 2944 19564 2972
rect 21821 2975 21879 2981
rect 18564 2932 18570 2944
rect 21821 2941 21833 2975
rect 21867 2972 21879 2975
rect 22094 2972 22100 2984
rect 21867 2944 22100 2972
rect 21867 2941 21879 2944
rect 21821 2935 21879 2941
rect 22094 2932 22100 2944
rect 22152 2932 22158 2984
rect 19334 2904 19340 2916
rect 14323 2876 15148 2904
rect 16500 2876 19340 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 13780 2808 13860 2836
rect 13780 2796 13786 2808
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14553 2839 14611 2845
rect 14553 2836 14565 2839
rect 14240 2808 14565 2836
rect 14240 2796 14246 2808
rect 14553 2805 14565 2808
rect 14599 2805 14611 2839
rect 15120 2836 15148 2876
rect 19334 2864 19340 2876
rect 19392 2864 19398 2916
rect 23032 2904 23060 3003
rect 19444 2876 23060 2904
rect 16574 2836 16580 2848
rect 15120 2808 16580 2836
rect 14553 2799 14611 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 19444 2836 19472 2876
rect 17460 2808 19472 2836
rect 19521 2839 19579 2845
rect 17460 2796 17466 2808
rect 19521 2805 19533 2839
rect 19567 2836 19579 2839
rect 19610 2836 19616 2848
rect 19567 2808 19616 2836
rect 19567 2805 19579 2808
rect 19521 2799 19579 2805
rect 19610 2796 19616 2808
rect 19668 2796 19674 2848
rect 19702 2796 19708 2848
rect 19760 2796 19766 2848
rect 1104 2746 23644 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 23644 2746
rect 1104 2672 23644 2694
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4614 2632 4620 2644
rect 4203 2604 4620 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 6089 2635 6147 2641
rect 6089 2632 6101 2635
rect 5684 2604 6101 2632
rect 5684 2592 5690 2604
rect 6089 2601 6101 2604
rect 6135 2601 6147 2635
rect 6089 2595 6147 2601
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 7374 2632 7380 2644
rect 7331 2604 7380 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 7466 2592 7472 2644
rect 7524 2592 7530 2644
rect 8110 2592 8116 2644
rect 8168 2632 8174 2644
rect 8168 2604 9536 2632
rect 8168 2592 8174 2604
rect 4801 2567 4859 2573
rect 4801 2533 4813 2567
rect 4847 2564 4859 2567
rect 8386 2564 8392 2576
rect 4847 2536 8392 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 8386 2524 8392 2536
rect 8444 2524 8450 2576
rect 8754 2524 8760 2576
rect 8812 2524 8818 2576
rect 9309 2567 9367 2573
rect 9309 2533 9321 2567
rect 9355 2533 9367 2567
rect 9508 2564 9536 2604
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11020 2604 13124 2632
rect 11020 2592 11026 2604
rect 11790 2564 11796 2576
rect 9508 2536 11796 2564
rect 9309 2527 9367 2533
rect 6822 2456 6828 2508
rect 6880 2456 6886 2508
rect 7834 2496 7840 2508
rect 6932 2468 7840 2496
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6932 2437 6960 2468
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8404 2496 8432 2524
rect 9324 2496 9352 2527
rect 11790 2524 11796 2536
rect 11848 2524 11854 2576
rect 11885 2567 11943 2573
rect 11885 2533 11897 2567
rect 11931 2564 11943 2567
rect 12986 2564 12992 2576
rect 11931 2536 12992 2564
rect 11931 2533 11943 2536
rect 11885 2527 11943 2533
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 13096 2573 13124 2604
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 15197 2635 15255 2641
rect 15197 2632 15209 2635
rect 13872 2604 15209 2632
rect 13872 2592 13878 2604
rect 15197 2601 15209 2604
rect 15243 2632 15255 2635
rect 16482 2632 16488 2644
rect 15243 2604 16488 2632
rect 15243 2601 15255 2604
rect 15197 2595 15255 2601
rect 16482 2592 16488 2604
rect 16540 2592 16546 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 17218 2632 17224 2644
rect 16632 2604 17224 2632
rect 16632 2592 16638 2604
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 18877 2635 18935 2641
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 19242 2632 19248 2644
rect 18923 2604 19248 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 23290 2592 23296 2644
rect 23348 2592 23354 2644
rect 13081 2567 13139 2573
rect 13081 2533 13093 2567
rect 13127 2533 13139 2567
rect 13081 2527 13139 2533
rect 17862 2524 17868 2576
rect 17920 2564 17926 2576
rect 19426 2564 19432 2576
rect 17920 2536 19432 2564
rect 17920 2524 17926 2536
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 22922 2524 22928 2576
rect 22980 2524 22986 2576
rect 9950 2496 9956 2508
rect 8404 2468 9168 2496
rect 9324 2468 9956 2496
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 5460 2332 6224 2360
rect 5460 2301 5488 2332
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2261 5503 2295
rect 6196 2292 6224 2332
rect 6932 2292 6960 2391
rect 7282 2388 7288 2440
rect 7340 2388 7346 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 9140 2437 9168 2468
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 10796 2468 19104 2496
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7800 2400 7941 2428
rect 7800 2388 7806 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 7929 2391 7987 2397
rect 8496 2400 8585 2428
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 7653 2363 7711 2369
rect 7653 2360 7665 2363
rect 7156 2332 7665 2360
rect 7156 2320 7162 2332
rect 7653 2329 7665 2332
rect 7699 2329 7711 2363
rect 7653 2323 7711 2329
rect 7837 2363 7895 2369
rect 7837 2329 7849 2363
rect 7883 2360 7895 2363
rect 8018 2360 8024 2372
rect 7883 2332 8024 2360
rect 7883 2329 7895 2332
rect 7837 2323 7895 2329
rect 8018 2320 8024 2332
rect 8076 2320 8082 2372
rect 8496 2304 8524 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9490 2388 9496 2440
rect 9548 2388 9554 2440
rect 10042 2388 10048 2440
rect 10100 2388 10106 2440
rect 10796 2437 10824 2468
rect 10781 2431 10839 2437
rect 10781 2397 10793 2431
rect 10827 2397 10839 2431
rect 10781 2391 10839 2397
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 10962 2428 10968 2440
rect 10919 2400 10968 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11698 2388 11704 2440
rect 11756 2388 11762 2440
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 10502 2320 10508 2372
rect 10560 2320 10566 2372
rect 11992 2360 12020 2391
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 12216 2400 12265 2428
rect 12216 2388 12222 2400
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12400 2400 12449 2428
rect 12400 2388 12406 2400
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 12894 2388 12900 2440
rect 12952 2388 12958 2440
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 13078 2360 13084 2372
rect 11992 2332 13084 2360
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 6196 2264 6960 2292
rect 5445 2255 5503 2261
rect 8478 2252 8484 2304
rect 8536 2252 8542 2304
rect 9674 2252 9680 2304
rect 9732 2252 9738 2304
rect 9950 2252 9956 2304
rect 10008 2252 10014 2304
rect 10226 2252 10232 2304
rect 10284 2252 10290 2304
rect 11054 2252 11060 2304
rect 11112 2252 11118 2304
rect 11330 2252 11336 2304
rect 11388 2252 11394 2304
rect 12158 2252 12164 2304
rect 12216 2252 12222 2304
rect 12345 2295 12403 2301
rect 12345 2261 12357 2295
rect 12391 2292 12403 2295
rect 12618 2292 12624 2304
rect 12391 2264 12624 2292
rect 12391 2261 12403 2264
rect 12345 2255 12403 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 12710 2252 12716 2304
rect 12768 2252 12774 2304
rect 13188 2292 13216 2391
rect 13372 2360 13400 2391
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14090 2388 14096 2440
rect 14148 2388 14154 2440
rect 14274 2388 14280 2440
rect 14332 2428 14338 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14332 2400 14565 2428
rect 14332 2388 14338 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2428 16543 2431
rect 17862 2428 17868 2440
rect 16531 2400 17868 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 18414 2388 18420 2440
rect 18472 2388 18478 2440
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 18966 2388 18972 2440
rect 19024 2388 19030 2440
rect 19076 2428 19104 2468
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19886 2496 19892 2508
rect 19392 2468 19892 2496
rect 19392 2456 19398 2468
rect 19886 2456 19892 2468
rect 19944 2456 19950 2508
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 20036 2468 21833 2496
rect 20036 2456 20042 2468
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 22097 2499 22155 2505
rect 22097 2465 22109 2499
rect 22143 2496 22155 2499
rect 22370 2496 22376 2508
rect 22143 2468 22376 2496
rect 22143 2465 22155 2468
rect 22097 2459 22155 2465
rect 22370 2456 22376 2468
rect 22428 2456 22434 2508
rect 22462 2456 22468 2508
rect 22520 2496 22526 2508
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22520 2468 23029 2496
rect 22520 2456 22526 2468
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 23017 2459 23075 2465
rect 19521 2431 19579 2437
rect 19076 2400 19380 2428
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 13372 2332 14381 2360
rect 14369 2329 14381 2332
rect 14415 2360 14427 2363
rect 15746 2360 15752 2372
rect 14415 2332 15752 2360
rect 14415 2329 14427 2332
rect 14369 2323 14427 2329
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 16669 2363 16727 2369
rect 16669 2329 16681 2363
rect 16715 2360 16727 2363
rect 17126 2360 17132 2372
rect 16715 2332 17132 2360
rect 16715 2329 16727 2332
rect 16669 2323 16727 2329
rect 16684 2292 16712 2323
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 17218 2320 17224 2372
rect 17276 2360 17282 2372
rect 19245 2363 19303 2369
rect 19245 2360 19257 2363
rect 17276 2332 19257 2360
rect 17276 2320 17282 2332
rect 19245 2329 19257 2332
rect 19291 2329 19303 2363
rect 19352 2360 19380 2400
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 20254 2428 20260 2440
rect 19567 2400 20260 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 22830 2388 22836 2440
rect 22888 2388 22894 2440
rect 23109 2431 23167 2437
rect 23109 2397 23121 2431
rect 23155 2397 23167 2431
rect 23109 2391 23167 2397
rect 19352 2332 19656 2360
rect 19245 2323 19303 2329
rect 13188 2264 16712 2292
rect 19337 2295 19395 2301
rect 19337 2261 19349 2295
rect 19383 2292 19395 2295
rect 19518 2292 19524 2304
rect 19383 2264 19524 2292
rect 19383 2261 19395 2264
rect 19337 2255 19395 2261
rect 19518 2252 19524 2264
rect 19576 2252 19582 2304
rect 19628 2292 19656 2332
rect 19702 2320 19708 2372
rect 19760 2320 19766 2372
rect 21634 2320 21640 2372
rect 21692 2320 21698 2372
rect 21726 2320 21732 2372
rect 21784 2360 21790 2372
rect 23124 2360 23152 2391
rect 21784 2332 23152 2360
rect 21784 2320 21790 2332
rect 22278 2292 22284 2304
rect 19628 2264 22284 2292
rect 22278 2252 22284 2264
rect 22336 2252 22342 2304
rect 1104 2202 23644 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 23644 2202
rect 1104 2128 23644 2150
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 16758 2088 16764 2100
rect 11204 2060 16764 2088
rect 11204 2048 11210 2060
rect 16758 2048 16764 2060
rect 16816 2048 16822 2100
rect 11698 1980 11704 2032
rect 11756 2020 11762 2032
rect 14734 2020 14740 2032
rect 11756 1992 14740 2020
rect 11756 1980 11762 1992
rect 14734 1980 14740 1992
rect 14792 1980 14798 2032
rect 10870 1912 10876 1964
rect 10928 1952 10934 1964
rect 19702 1952 19708 1964
rect 10928 1924 19708 1952
rect 10928 1912 10934 1924
rect 19702 1912 19708 1924
rect 19760 1912 19766 1964
rect 10042 1844 10048 1896
rect 10100 1884 10106 1896
rect 14918 1884 14924 1896
rect 10100 1856 14924 1884
rect 10100 1844 10106 1856
rect 14918 1844 14924 1856
rect 14976 1844 14982 1896
rect 9490 1776 9496 1828
rect 9548 1816 9554 1828
rect 16666 1816 16672 1828
rect 9548 1788 16672 1816
rect 9548 1776 9554 1788
rect 16666 1776 16672 1788
rect 16724 1776 16730 1828
rect 13078 1708 13084 1760
rect 13136 1748 13142 1760
rect 19610 1748 19616 1760
rect 13136 1720 19616 1748
rect 13136 1708 13142 1720
rect 19610 1708 19616 1720
rect 19668 1708 19674 1760
rect 8018 1640 8024 1692
rect 8076 1680 8082 1692
rect 8076 1652 12434 1680
rect 8076 1640 8082 1652
rect 12406 1612 12434 1652
rect 12710 1640 12716 1692
rect 12768 1680 12774 1692
rect 14826 1680 14832 1692
rect 12768 1652 14832 1680
rect 12768 1640 12774 1652
rect 14826 1640 14832 1652
rect 14884 1640 14890 1692
rect 14090 1612 14096 1624
rect 12406 1584 14096 1612
rect 14090 1572 14096 1584
rect 14148 1612 14154 1624
rect 15470 1612 15476 1624
rect 14148 1584 15476 1612
rect 14148 1572 14154 1584
rect 15470 1572 15476 1584
rect 15528 1572 15534 1624
rect 11238 1300 11244 1352
rect 11296 1340 11302 1352
rect 18690 1340 18696 1352
rect 11296 1312 18696 1340
rect 11296 1300 11302 1312
rect 18690 1300 18696 1312
rect 18748 1300 18754 1352
rect 11054 1232 11060 1284
rect 11112 1272 11118 1284
rect 17402 1272 17408 1284
rect 11112 1244 17408 1272
rect 11112 1232 11118 1244
rect 17402 1232 17408 1244
rect 17460 1232 17466 1284
rect 12158 1164 12164 1216
rect 12216 1204 12222 1216
rect 16114 1204 16120 1216
rect 12216 1176 16120 1204
rect 12216 1164 12222 1176
rect 16114 1164 16120 1176
rect 16172 1164 16178 1216
rect 10226 1096 10232 1148
rect 10284 1136 10290 1148
rect 18046 1136 18052 1148
rect 10284 1108 18052 1136
rect 10284 1096 10290 1108
rect 18046 1096 18052 1108
rect 18104 1096 18110 1148
rect 11330 1028 11336 1080
rect 11388 1068 11394 1080
rect 16758 1068 16764 1080
rect 11388 1040 16764 1068
rect 11388 1028 11394 1040
rect 16758 1028 16764 1040
rect 16816 1028 16822 1080
rect 12986 960 12992 1012
rect 13044 1000 13050 1012
rect 15470 1000 15476 1012
rect 13044 972 15476 1000
rect 13044 960 13050 972
rect 15470 960 15476 972
rect 15528 960 15534 1012
rect 9950 620 9956 672
rect 10008 660 10014 672
rect 21910 660 21916 672
rect 10008 632 21916 660
rect 10008 620 10014 632
rect 21910 620 21916 632
rect 21968 620 21974 672
rect 10502 76 10508 128
rect 10560 116 10566 128
rect 19334 116 19340 128
rect 10560 88 19340 116
rect 10560 76 10566 88
rect 19334 76 19340 88
rect 19392 76 19398 128
<< via1 >>
rect 16212 13268 16264 13320
rect 23112 13268 23164 13320
rect 16948 11024 17000 11076
rect 20628 11024 20680 11076
rect 14188 10956 14240 11008
rect 15016 10956 15068 11008
rect 16396 10956 16448 11008
rect 21456 10956 21508 11008
rect 21548 10956 21600 11008
rect 22652 10956 22704 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 9680 10752 9732 10804
rect 11612 10752 11664 10804
rect 13544 10752 13596 10804
rect 14832 10752 14884 10804
rect 15476 10752 15528 10804
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 16764 10752 16816 10804
rect 17408 10752 17460 10804
rect 19340 10752 19392 10804
rect 1952 10616 2004 10668
rect 3332 10616 3384 10668
rect 1308 10548 1360 10600
rect 4712 10616 4764 10668
rect 9036 10616 9088 10668
rect 9956 10616 10008 10668
rect 10968 10616 11020 10668
rect 15200 10684 15252 10736
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 12900 10616 12952 10668
rect 13912 10616 13964 10668
rect 14648 10659 14700 10668
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 4804 10548 4856 10600
rect 13084 10548 13136 10600
rect 5448 10480 5500 10532
rect 12072 10480 12124 10532
rect 15016 10616 15068 10668
rect 17868 10684 17920 10736
rect 16488 10659 16540 10668
rect 16488 10625 16497 10659
rect 16497 10625 16531 10659
rect 16531 10625 16540 10659
rect 16488 10616 16540 10625
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 17684 10616 17736 10668
rect 17776 10659 17828 10668
rect 17776 10625 17785 10659
rect 17785 10625 17819 10659
rect 17819 10625 17828 10659
rect 17776 10616 17828 10625
rect 18512 10548 18564 10600
rect 18788 10659 18840 10668
rect 18788 10625 18797 10659
rect 18797 10625 18831 10659
rect 18831 10625 18840 10659
rect 18788 10616 18840 10625
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 22468 10684 22520 10736
rect 388 10412 440 10464
rect 4068 10412 4120 10464
rect 5816 10412 5868 10464
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 11612 10412 11664 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 12716 10412 12768 10464
rect 15476 10455 15528 10464
rect 15476 10421 15485 10455
rect 15485 10421 15519 10455
rect 15519 10421 15528 10455
rect 15476 10412 15528 10421
rect 16028 10480 16080 10532
rect 16580 10480 16632 10532
rect 16672 10412 16724 10464
rect 17132 10480 17184 10532
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 18604 10480 18656 10532
rect 18880 10412 18932 10464
rect 19248 10412 19300 10464
rect 19524 10480 19576 10532
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 22376 10659 22428 10668
rect 22376 10625 22385 10659
rect 22385 10625 22419 10659
rect 22419 10625 22428 10659
rect 22376 10616 22428 10625
rect 22744 10684 22796 10736
rect 23112 10684 23164 10736
rect 21180 10591 21232 10600
rect 21180 10557 21189 10591
rect 21189 10557 21223 10591
rect 21223 10557 21232 10591
rect 21180 10548 21232 10557
rect 22376 10480 22428 10532
rect 20628 10455 20680 10464
rect 20628 10421 20637 10455
rect 20637 10421 20671 10455
rect 20671 10421 20680 10455
rect 20628 10412 20680 10421
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 21456 10412 21508 10464
rect 22100 10412 22152 10464
rect 22652 10480 22704 10532
rect 22836 10455 22888 10464
rect 22836 10421 22845 10455
rect 22845 10421 22879 10455
rect 22879 10421 22888 10455
rect 22836 10412 22888 10421
rect 22928 10455 22980 10464
rect 22928 10421 22937 10455
rect 22937 10421 22971 10455
rect 22971 10421 22980 10455
rect 22928 10412 22980 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 6552 10208 6604 10260
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 12072 10208 12124 10260
rect 12624 10208 12676 10260
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 5356 10072 5408 10124
rect 7012 10115 7064 10124
rect 7012 10081 7021 10115
rect 7021 10081 7055 10115
rect 7055 10081 7064 10115
rect 7012 10072 7064 10081
rect 7748 10115 7800 10124
rect 7748 10081 7757 10115
rect 7757 10081 7791 10115
rect 7791 10081 7800 10115
rect 7748 10072 7800 10081
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 3332 10004 3384 10056
rect 5448 10004 5500 10056
rect 5816 10047 5868 10056
rect 5816 10013 5825 10047
rect 5825 10013 5859 10047
rect 5859 10013 5868 10047
rect 5816 10004 5868 10013
rect 4620 9936 4672 9988
rect 5172 9936 5224 9988
rect 6184 9979 6236 9988
rect 6184 9945 6193 9979
rect 6193 9945 6227 9979
rect 6227 9945 6236 9979
rect 6184 9936 6236 9945
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 9312 10004 9364 10056
rect 6920 9936 6972 9988
rect 388 9868 440 9920
rect 4528 9911 4580 9920
rect 4528 9877 4537 9911
rect 4537 9877 4571 9911
rect 4571 9877 4580 9911
rect 4528 9868 4580 9877
rect 5724 9868 5776 9920
rect 6736 9868 6788 9920
rect 7472 9868 7524 9920
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 12900 10140 12952 10192
rect 14648 10140 14700 10192
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 10416 10004 10468 10056
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 11612 10072 11664 10124
rect 11428 10004 11480 10056
rect 10692 9979 10744 9988
rect 10692 9945 10701 9979
rect 10701 9945 10735 9979
rect 10735 9945 10744 9979
rect 10692 9936 10744 9945
rect 12440 10072 12492 10124
rect 7656 9911 7708 9920
rect 7656 9877 7665 9911
rect 7665 9877 7699 9911
rect 7699 9877 7708 9911
rect 7656 9868 7708 9877
rect 9772 9868 9824 9920
rect 10600 9868 10652 9920
rect 11336 9911 11388 9920
rect 11336 9877 11345 9911
rect 11345 9877 11379 9911
rect 11379 9877 11388 9911
rect 11336 9868 11388 9877
rect 11704 9868 11756 9920
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 12164 10004 12216 10056
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 14188 10004 14240 10056
rect 14832 10004 14884 10056
rect 12624 9936 12676 9988
rect 12808 9936 12860 9988
rect 15016 10004 15068 10056
rect 15384 10072 15436 10124
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 17776 10208 17828 10260
rect 18880 10208 18932 10260
rect 21548 10208 21600 10260
rect 21916 10208 21968 10260
rect 17316 10140 17368 10192
rect 18144 10072 18196 10124
rect 18236 10072 18288 10124
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 14280 9868 14332 9920
rect 14556 9868 14608 9920
rect 15568 9868 15620 9920
rect 15752 9868 15804 9920
rect 17776 10004 17828 10056
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 18604 10004 18656 10056
rect 18788 10004 18840 10056
rect 19156 10072 19208 10124
rect 19064 10004 19116 10056
rect 20628 10072 20680 10124
rect 19524 10047 19576 10056
rect 19524 10013 19533 10047
rect 19533 10013 19567 10047
rect 19567 10013 19576 10047
rect 19524 10004 19576 10013
rect 21180 10004 21232 10056
rect 22652 10004 22704 10056
rect 23112 10004 23164 10056
rect 18328 9979 18380 9988
rect 18328 9945 18337 9979
rect 18337 9945 18371 9979
rect 18371 9945 18380 9979
rect 18328 9936 18380 9945
rect 19984 9979 20036 9988
rect 19984 9945 19993 9979
rect 19993 9945 20027 9979
rect 20027 9945 20036 9979
rect 19984 9936 20036 9945
rect 21088 9936 21140 9988
rect 21364 9936 21416 9988
rect 20168 9868 20220 9920
rect 22468 9868 22520 9920
rect 23204 9911 23256 9920
rect 23204 9877 23213 9911
rect 23213 9877 23247 9911
rect 23247 9877 23256 9911
rect 23204 9868 23256 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1676 9664 1728 9716
rect 4528 9664 4580 9716
rect 5724 9707 5776 9716
rect 5724 9673 5733 9707
rect 5733 9673 5767 9707
rect 5767 9673 5776 9707
rect 5724 9664 5776 9673
rect 6000 9664 6052 9716
rect 6828 9664 6880 9716
rect 7012 9664 7064 9716
rect 8484 9707 8536 9716
rect 8484 9673 8493 9707
rect 8493 9673 8527 9707
rect 8527 9673 8536 9707
rect 8484 9664 8536 9673
rect 11520 9664 11572 9716
rect 12164 9664 12216 9716
rect 5080 9596 5132 9648
rect 4620 9528 4672 9580
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 5632 9460 5684 9512
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 7656 9639 7708 9648
rect 7656 9605 7665 9639
rect 7665 9605 7699 9639
rect 7699 9605 7708 9639
rect 7656 9596 7708 9605
rect 7012 9528 7064 9580
rect 8300 9528 8352 9580
rect 8668 9528 8720 9580
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 9220 9528 9272 9580
rect 9864 9596 9916 9648
rect 10232 9596 10284 9648
rect 4712 9392 4764 9444
rect 5816 9392 5868 9444
rect 6828 9392 6880 9444
rect 10416 9528 10468 9580
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 12440 9664 12492 9716
rect 12808 9664 12860 9716
rect 12900 9707 12952 9716
rect 12900 9673 12909 9707
rect 12909 9673 12943 9707
rect 12943 9673 12952 9707
rect 12900 9664 12952 9673
rect 13084 9664 13136 9716
rect 12348 9596 12400 9648
rect 10784 9528 10836 9537
rect 10692 9460 10744 9512
rect 12256 9460 12308 9512
rect 12808 9528 12860 9580
rect 14096 9528 14148 9580
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 15108 9639 15160 9648
rect 15108 9605 15117 9639
rect 15117 9605 15151 9639
rect 15151 9605 15160 9639
rect 15108 9596 15160 9605
rect 15752 9639 15804 9648
rect 15752 9605 15761 9639
rect 15761 9605 15795 9639
rect 15795 9605 15804 9639
rect 15752 9596 15804 9605
rect 16672 9664 16724 9716
rect 17316 9639 17368 9648
rect 12532 9503 12584 9512
rect 12532 9469 12541 9503
rect 12541 9469 12575 9503
rect 12575 9469 12584 9503
rect 12532 9460 12584 9469
rect 15476 9528 15528 9580
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 16028 9571 16080 9580
rect 16028 9537 16037 9571
rect 16037 9537 16071 9571
rect 16071 9537 16080 9571
rect 16028 9528 16080 9537
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 17316 9605 17325 9639
rect 17325 9605 17359 9639
rect 17359 9605 17368 9639
rect 17316 9596 17368 9605
rect 16764 9571 16816 9580
rect 16764 9537 16773 9571
rect 16773 9537 16807 9571
rect 16807 9537 16816 9571
rect 16764 9528 16816 9537
rect 16856 9528 16908 9580
rect 17776 9571 17828 9580
rect 11428 9392 11480 9444
rect 12900 9392 12952 9444
rect 14004 9392 14056 9444
rect 4068 9324 4120 9376
rect 4988 9324 5040 9376
rect 6092 9324 6144 9376
rect 6368 9324 6420 9376
rect 7288 9324 7340 9376
rect 9956 9324 10008 9376
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 11796 9324 11848 9376
rect 13820 9324 13872 9376
rect 17040 9503 17092 9512
rect 17040 9469 17049 9503
rect 17049 9469 17083 9503
rect 17083 9469 17092 9503
rect 17040 9460 17092 9469
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 18052 9596 18104 9648
rect 18696 9528 18748 9580
rect 19340 9528 19392 9580
rect 20168 9528 20220 9580
rect 20720 9528 20772 9580
rect 24492 9596 24544 9648
rect 16764 9392 16816 9444
rect 18052 9460 18104 9512
rect 18144 9460 18196 9512
rect 21272 9460 21324 9512
rect 17500 9392 17552 9444
rect 16580 9324 16632 9376
rect 17408 9324 17460 9376
rect 17960 9324 18012 9376
rect 18420 9324 18472 9376
rect 21732 9324 21784 9376
rect 21824 9367 21876 9376
rect 21824 9333 21833 9367
rect 21833 9333 21867 9367
rect 21867 9333 21876 9367
rect 22284 9392 22336 9444
rect 22560 9528 22612 9580
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 23388 9392 23440 9444
rect 21824 9324 21876 9333
rect 22652 9324 22704 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 5908 9120 5960 9172
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 6920 9120 6972 9172
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 9588 9120 9640 9172
rect 10508 9120 10560 9172
rect 11704 9163 11756 9172
rect 11704 9129 11713 9163
rect 11713 9129 11747 9163
rect 11747 9129 11756 9163
rect 11704 9120 11756 9129
rect 5356 9052 5408 9104
rect 6276 9095 6328 9104
rect 6276 9061 6285 9095
rect 6285 9061 6319 9095
rect 6319 9061 6328 9095
rect 6276 9052 6328 9061
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3332 8959 3384 8968
rect 3332 8925 3341 8959
rect 3341 8925 3375 8959
rect 3375 8925 3384 8959
rect 3332 8916 3384 8925
rect 5080 8984 5132 9036
rect 7288 8984 7340 9036
rect 8852 9052 8904 9104
rect 9312 9052 9364 9104
rect 7748 9027 7800 9036
rect 7748 8993 7757 9027
rect 7757 8993 7791 9027
rect 7791 8993 7800 9027
rect 7748 8984 7800 8993
rect 3792 8848 3844 8900
rect 4988 8916 5040 8968
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 5908 8916 5960 8968
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 4804 8780 4856 8832
rect 5632 8823 5684 8832
rect 5632 8789 5641 8823
rect 5641 8789 5675 8823
rect 5675 8789 5684 8823
rect 5632 8780 5684 8789
rect 6184 8848 6236 8900
rect 8300 8916 8352 8968
rect 8944 8984 8996 9036
rect 9588 8984 9640 9036
rect 13544 9120 13596 9172
rect 15016 9163 15068 9172
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 15108 9120 15160 9172
rect 15476 9120 15528 9172
rect 16304 9120 16356 9172
rect 16396 9120 16448 9172
rect 16672 9163 16724 9172
rect 16672 9129 16681 9163
rect 16681 9129 16715 9163
rect 16715 9129 16724 9163
rect 16672 9120 16724 9129
rect 17408 9163 17460 9172
rect 17408 9129 17417 9163
rect 17417 9129 17451 9163
rect 17451 9129 17460 9163
rect 17408 9120 17460 9129
rect 17684 9163 17736 9172
rect 17684 9129 17693 9163
rect 17693 9129 17727 9163
rect 17727 9129 17736 9163
rect 17684 9120 17736 9129
rect 18512 9163 18564 9172
rect 18512 9129 18521 9163
rect 18521 9129 18555 9163
rect 18555 9129 18564 9163
rect 18512 9120 18564 9129
rect 8024 8848 8076 8900
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9404 8916 9456 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 10416 8959 10468 8968
rect 10416 8925 10424 8959
rect 10424 8925 10458 8959
rect 10458 8925 10468 8959
rect 10416 8916 10468 8925
rect 11520 8984 11572 9036
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 10876 8916 10928 8968
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 12808 9052 12860 9104
rect 15200 9052 15252 9104
rect 16028 9052 16080 9104
rect 16212 9095 16264 9104
rect 16212 9061 16221 9095
rect 16221 9061 16255 9095
rect 16255 9061 16264 9095
rect 16212 9052 16264 9061
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 13820 8984 13872 8993
rect 17040 9052 17092 9104
rect 17316 9095 17368 9104
rect 17316 9061 17325 9095
rect 17325 9061 17359 9095
rect 17359 9061 17368 9095
rect 17316 9052 17368 9061
rect 17776 9052 17828 9104
rect 18328 9052 18380 9104
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 12256 8916 12308 8968
rect 14556 8916 14608 8968
rect 14924 8916 14976 8968
rect 15108 8959 15160 8968
rect 15108 8925 15117 8959
rect 15117 8925 15151 8959
rect 15151 8925 15160 8959
rect 15108 8916 15160 8925
rect 15200 8916 15252 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 15752 8959 15804 8968
rect 15752 8925 15785 8959
rect 15785 8925 15804 8959
rect 15752 8916 15804 8925
rect 16120 8916 16172 8968
rect 16672 8984 16724 9036
rect 17500 8984 17552 9036
rect 16488 8959 16540 8968
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 16580 8916 16632 8968
rect 17040 8959 17092 8968
rect 17040 8925 17049 8959
rect 17049 8925 17083 8959
rect 17083 8925 17092 8959
rect 17040 8916 17092 8925
rect 12992 8848 13044 8900
rect 13268 8848 13320 8900
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 18052 8916 18104 8968
rect 18236 8916 18288 8968
rect 18788 9052 18840 9104
rect 19708 9120 19760 9172
rect 20720 9163 20772 9172
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 23848 9120 23900 9172
rect 20996 9052 21048 9104
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 19064 8959 19116 8968
rect 19064 8925 19073 8959
rect 19073 8925 19107 8959
rect 19107 8925 19116 8959
rect 19064 8916 19116 8925
rect 19156 8916 19208 8968
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 19616 8959 19668 8968
rect 19616 8925 19626 8959
rect 19626 8925 19660 8959
rect 19660 8925 19668 8959
rect 19616 8916 19668 8925
rect 8668 8780 8720 8832
rect 9128 8780 9180 8832
rect 11152 8780 11204 8832
rect 11336 8823 11388 8832
rect 11336 8789 11345 8823
rect 11345 8789 11379 8823
rect 11379 8789 11388 8823
rect 11336 8780 11388 8789
rect 11428 8780 11480 8832
rect 11888 8780 11940 8832
rect 12072 8780 12124 8832
rect 12348 8780 12400 8832
rect 12808 8780 12860 8832
rect 13084 8823 13136 8832
rect 13084 8789 13093 8823
rect 13093 8789 13127 8823
rect 13127 8789 13136 8823
rect 13084 8780 13136 8789
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 19800 8848 19852 8900
rect 19892 8891 19944 8900
rect 19892 8857 19901 8891
rect 19901 8857 19935 8891
rect 19935 8857 19944 8891
rect 19892 8848 19944 8857
rect 16856 8780 16908 8832
rect 17316 8780 17368 8832
rect 17960 8780 18012 8832
rect 18972 8780 19024 8832
rect 19248 8780 19300 8832
rect 22376 8984 22428 9036
rect 21916 8916 21968 8968
rect 22100 8916 22152 8968
rect 22468 8959 22520 8968
rect 22468 8925 22477 8959
rect 22477 8925 22511 8959
rect 22511 8925 22520 8959
rect 22468 8916 22520 8925
rect 22744 8959 22796 8968
rect 22744 8925 22753 8959
rect 22753 8925 22787 8959
rect 22787 8925 22796 8959
rect 22744 8916 22796 8925
rect 22192 8848 22244 8900
rect 20260 8780 20312 8832
rect 21364 8780 21416 8832
rect 22836 8780 22888 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3240 8576 3292 8628
rect 3792 8619 3844 8628
rect 3792 8585 3801 8619
rect 3801 8585 3835 8619
rect 3835 8585 3844 8619
rect 3792 8576 3844 8585
rect 4160 8576 4212 8628
rect 4068 8508 4120 8560
rect 5356 8576 5408 8628
rect 7748 8576 7800 8628
rect 3884 8440 3936 8492
rect 5448 8508 5500 8560
rect 4804 8440 4856 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 4988 8440 5040 8492
rect 7012 8508 7064 8560
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 8852 8508 8904 8560
rect 9680 8508 9732 8560
rect 10600 8508 10652 8560
rect 12532 8576 12584 8628
rect 13636 8576 13688 8628
rect 14096 8619 14148 8628
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 14464 8576 14516 8628
rect 12256 8508 12308 8560
rect 14648 8508 14700 8560
rect 5632 8440 5684 8492
rect 6460 8483 6512 8492
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6460 8440 6512 8449
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 5356 8372 5408 8424
rect 5908 8304 5960 8356
rect 8944 8372 8996 8424
rect 9588 8440 9640 8492
rect 11428 8440 11480 8492
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 11152 8372 11204 8424
rect 6092 8304 6144 8356
rect 8208 8304 8260 8356
rect 9404 8304 9456 8356
rect 4896 8236 4948 8288
rect 5448 8236 5500 8288
rect 5632 8236 5684 8288
rect 7748 8236 7800 8288
rect 8576 8236 8628 8288
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 9956 8304 10008 8356
rect 12532 8440 12584 8492
rect 13268 8440 13320 8492
rect 12164 8415 12216 8424
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 14556 8372 14608 8424
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 15660 8508 15712 8560
rect 15568 8483 15620 8492
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 14924 8372 14976 8381
rect 15844 8576 15896 8628
rect 16028 8619 16080 8628
rect 16028 8585 16037 8619
rect 16037 8585 16071 8619
rect 16071 8585 16080 8619
rect 16028 8576 16080 8585
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 17224 8576 17276 8628
rect 18696 8576 18748 8628
rect 16856 8508 16908 8560
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 15292 8304 15344 8356
rect 11888 8236 11940 8288
rect 11980 8279 12032 8288
rect 11980 8245 11989 8279
rect 11989 8245 12023 8279
rect 12023 8245 12032 8279
rect 11980 8236 12032 8245
rect 13360 8236 13412 8288
rect 13820 8236 13872 8288
rect 16580 8372 16632 8424
rect 17316 8440 17368 8492
rect 17592 8508 17644 8560
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 17960 8508 18012 8560
rect 18328 8551 18380 8560
rect 18328 8517 18353 8551
rect 18353 8517 18380 8551
rect 18328 8508 18380 8517
rect 18604 8440 18656 8492
rect 18972 8508 19024 8560
rect 19708 8440 19760 8492
rect 20168 8440 20220 8492
rect 16856 8347 16908 8356
rect 16856 8313 16865 8347
rect 16865 8313 16899 8347
rect 16899 8313 16908 8347
rect 16856 8304 16908 8313
rect 17408 8304 17460 8356
rect 17592 8304 17644 8356
rect 18144 8304 18196 8356
rect 18512 8304 18564 8356
rect 18604 8304 18656 8356
rect 19800 8372 19852 8424
rect 21088 8576 21140 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 20904 8551 20956 8560
rect 20904 8517 20913 8551
rect 20913 8517 20947 8551
rect 20947 8517 20956 8551
rect 20904 8508 20956 8517
rect 21272 8508 21324 8560
rect 21640 8508 21692 8560
rect 23204 8576 23256 8628
rect 20352 8440 20404 8492
rect 20996 8483 21048 8492
rect 20996 8449 21010 8483
rect 21010 8449 21044 8483
rect 21044 8449 21048 8483
rect 20996 8440 21048 8449
rect 21548 8483 21600 8492
rect 21548 8449 21557 8483
rect 21557 8449 21591 8483
rect 21591 8449 21600 8483
rect 21548 8440 21600 8449
rect 21732 8440 21784 8492
rect 21916 8440 21968 8492
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22836 8440 22888 8492
rect 24216 8440 24268 8492
rect 16672 8236 16724 8288
rect 16948 8236 17000 8288
rect 17960 8236 18012 8288
rect 18236 8236 18288 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3792 8032 3844 8084
rect 4620 8032 4672 8084
rect 5356 8032 5408 8084
rect 5816 8032 5868 8084
rect 6828 8032 6880 8084
rect 7196 8032 7248 8084
rect 3332 7964 3384 8016
rect 5632 7964 5684 8016
rect 6460 7964 6512 8016
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 5356 7896 5408 7948
rect 388 7828 440 7880
rect 1952 7828 2004 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 4712 7760 4764 7812
rect 6092 7828 6144 7880
rect 6184 7760 6236 7812
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 6644 7760 6696 7812
rect 3884 7692 3936 7744
rect 7564 7871 7616 7880
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 9036 8032 9088 8084
rect 9496 8032 9548 8084
rect 10048 8032 10100 8084
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 8852 7964 8904 8016
rect 10324 7964 10376 8016
rect 12532 8007 12584 8016
rect 12532 7973 12541 8007
rect 12541 7973 12575 8007
rect 12575 7973 12584 8007
rect 12532 7964 12584 7973
rect 13176 8032 13228 8084
rect 15200 8075 15252 8084
rect 15200 8041 15209 8075
rect 15209 8041 15243 8075
rect 15243 8041 15252 8075
rect 15200 8032 15252 8041
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 13084 7964 13136 8016
rect 14372 7964 14424 8016
rect 17040 8032 17092 8084
rect 17592 8032 17644 8084
rect 7472 7760 7524 7812
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 9220 7896 9272 7948
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 9864 7871 9916 7880
rect 8208 7803 8260 7812
rect 8208 7769 8217 7803
rect 8217 7769 8251 7803
rect 8251 7769 8260 7803
rect 8208 7760 8260 7769
rect 8392 7803 8444 7812
rect 8392 7769 8401 7803
rect 8401 7769 8435 7803
rect 8435 7769 8444 7803
rect 8392 7760 8444 7769
rect 8944 7760 8996 7812
rect 9588 7692 9640 7744
rect 9864 7837 9868 7871
rect 9868 7837 9902 7871
rect 9902 7837 9916 7871
rect 9864 7828 9916 7837
rect 10600 7896 10652 7948
rect 11704 7896 11756 7948
rect 10324 7871 10376 7880
rect 10324 7837 10326 7871
rect 10326 7837 10360 7871
rect 10360 7837 10376 7871
rect 10324 7828 10376 7837
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12624 7828 12676 7880
rect 15292 7896 15344 7948
rect 15568 7896 15620 7948
rect 15660 7896 15712 7948
rect 17408 7896 17460 7948
rect 17960 8032 18012 8084
rect 18604 8032 18656 8084
rect 18788 8032 18840 8084
rect 19064 8032 19116 8084
rect 19156 8032 19208 8084
rect 22284 8032 22336 8084
rect 23020 8075 23072 8084
rect 23020 8041 23029 8075
rect 23029 8041 23063 8075
rect 23063 8041 23072 8075
rect 23020 8032 23072 8041
rect 19248 7964 19300 8016
rect 19524 7964 19576 8016
rect 20628 7964 20680 8016
rect 12808 7828 12860 7880
rect 9956 7803 10008 7812
rect 9956 7769 9965 7803
rect 9965 7769 9999 7803
rect 9999 7769 10008 7803
rect 9956 7760 10008 7769
rect 10048 7803 10100 7812
rect 10048 7769 10057 7803
rect 10057 7769 10091 7803
rect 10091 7769 10100 7803
rect 10048 7760 10100 7769
rect 12532 7760 12584 7812
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 14648 7828 14700 7880
rect 14372 7803 14424 7812
rect 14372 7769 14381 7803
rect 14381 7769 14415 7803
rect 14415 7769 14424 7803
rect 14372 7760 14424 7769
rect 15476 7828 15528 7880
rect 12072 7692 12124 7744
rect 12808 7692 12860 7744
rect 15752 7692 15804 7744
rect 15936 7803 15988 7812
rect 15936 7769 15945 7803
rect 15945 7769 15979 7803
rect 15979 7769 15988 7803
rect 15936 7760 15988 7769
rect 16120 7760 16172 7812
rect 16580 7828 16632 7880
rect 16856 7828 16908 7880
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 17224 7828 17276 7880
rect 17500 7828 17552 7880
rect 17764 7871 17816 7880
rect 17764 7837 17785 7871
rect 17785 7837 17816 7871
rect 17764 7828 17816 7837
rect 17316 7760 17368 7812
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 19064 7896 19116 7948
rect 18512 7828 18564 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 20720 7896 20772 7948
rect 20536 7828 20588 7880
rect 16304 7692 16356 7744
rect 17132 7692 17184 7744
rect 19340 7803 19392 7812
rect 19340 7769 19349 7803
rect 19349 7769 19383 7803
rect 19383 7769 19392 7803
rect 19340 7760 19392 7769
rect 20996 7803 21048 7812
rect 20996 7769 21005 7803
rect 21005 7769 21039 7803
rect 21039 7769 21048 7803
rect 20996 7760 21048 7769
rect 18144 7692 18196 7744
rect 18512 7692 18564 7744
rect 21088 7692 21140 7744
rect 22652 7692 22704 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4804 7488 4856 7540
rect 4068 7420 4120 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 4620 7420 4672 7472
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 6736 7488 6788 7540
rect 9220 7488 9272 7540
rect 9864 7488 9916 7540
rect 14372 7488 14424 7540
rect 15200 7488 15252 7540
rect 15568 7531 15620 7540
rect 15568 7497 15577 7531
rect 15577 7497 15611 7531
rect 15611 7497 15620 7531
rect 15568 7488 15620 7497
rect 17408 7488 17460 7540
rect 18052 7488 18104 7540
rect 19708 7488 19760 7540
rect 20720 7488 20772 7540
rect 5264 7420 5316 7472
rect 4344 7352 4396 7404
rect 6276 7420 6328 7472
rect 12164 7420 12216 7472
rect 3884 7284 3936 7336
rect 6460 7352 6512 7404
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 6092 7284 6144 7336
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 7932 7284 7984 7336
rect 8208 7284 8260 7336
rect 9128 7284 9180 7336
rect 10324 7352 10376 7404
rect 11704 7352 11756 7404
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 10508 7284 10560 7336
rect 12532 7352 12584 7404
rect 12992 7420 13044 7472
rect 15660 7420 15712 7472
rect 14740 7352 14792 7404
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 12164 7284 12216 7336
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 15568 7352 15620 7404
rect 15384 7284 15436 7336
rect 5264 7216 5316 7268
rect 5356 7259 5408 7268
rect 5356 7225 5365 7259
rect 5365 7225 5399 7259
rect 5399 7225 5408 7259
rect 5356 7216 5408 7225
rect 5816 7259 5868 7268
rect 5816 7225 5825 7259
rect 5825 7225 5859 7259
rect 5859 7225 5868 7259
rect 5816 7216 5868 7225
rect 6736 7216 6788 7268
rect 8392 7216 8444 7268
rect 8852 7259 8904 7268
rect 8852 7225 8861 7259
rect 8861 7225 8895 7259
rect 8895 7225 8904 7259
rect 8852 7216 8904 7225
rect 204 7148 256 7200
rect 3976 7191 4028 7200
rect 3976 7157 3985 7191
rect 3985 7157 4019 7191
rect 4019 7157 4028 7191
rect 3976 7148 4028 7157
rect 4344 7148 4396 7200
rect 4436 7148 4488 7200
rect 4804 7148 4856 7200
rect 6092 7148 6144 7200
rect 14096 7216 14148 7268
rect 9036 7148 9088 7200
rect 15108 7216 15160 7268
rect 17224 7420 17276 7472
rect 18236 7420 18288 7472
rect 16580 7352 16632 7404
rect 16764 7284 16816 7336
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17316 7395 17368 7404
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 17316 7352 17368 7361
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 17500 7352 17552 7404
rect 19708 7395 19760 7404
rect 19708 7361 19711 7395
rect 19711 7361 19745 7395
rect 19745 7361 19760 7395
rect 19708 7352 19760 7361
rect 21088 7420 21140 7472
rect 21548 7488 21600 7540
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 22284 7420 22336 7429
rect 22836 7420 22888 7472
rect 20720 7352 20772 7404
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 21456 7352 21508 7404
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 16488 7216 16540 7268
rect 17316 7216 17368 7268
rect 16212 7148 16264 7200
rect 16396 7191 16448 7200
rect 16396 7157 16405 7191
rect 16405 7157 16439 7191
rect 16439 7157 16448 7191
rect 16396 7148 16448 7157
rect 17040 7148 17092 7200
rect 22652 7352 22704 7404
rect 22928 7395 22980 7404
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 18604 7216 18656 7268
rect 21456 7216 21508 7268
rect 18236 7148 18288 7200
rect 19248 7148 19300 7200
rect 20444 7148 20496 7200
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 21180 7148 21232 7200
rect 23296 7216 23348 7268
rect 22376 7148 22428 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1952 6944 2004 6996
rect 4252 6944 4304 6996
rect 5724 6944 5776 6996
rect 7380 6944 7432 6996
rect 7748 6944 7800 6996
rect 9864 6944 9916 6996
rect 9956 6944 10008 6996
rect 13360 6944 13412 6996
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 1584 6740 1636 6792
rect 3332 6876 3384 6928
rect 5264 6876 5316 6928
rect 6092 6876 6144 6928
rect 6460 6919 6512 6928
rect 6460 6885 6469 6919
rect 6469 6885 6503 6919
rect 6503 6885 6512 6919
rect 6460 6876 6512 6885
rect 7932 6876 7984 6928
rect 10324 6876 10376 6928
rect 4160 6808 4212 6860
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 4712 6740 4764 6792
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 2136 6604 2188 6656
rect 4528 6672 4580 6724
rect 4620 6672 4672 6724
rect 5172 6672 5224 6724
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6552 6740 6604 6792
rect 8024 6740 8076 6792
rect 8852 6740 8904 6792
rect 9588 6740 9640 6792
rect 10048 6808 10100 6860
rect 10692 6808 10744 6860
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 11612 6808 11664 6817
rect 9864 6740 9916 6792
rect 6368 6672 6420 6724
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 3976 6604 4028 6656
rect 4344 6604 4396 6656
rect 5816 6604 5868 6656
rect 6000 6604 6052 6656
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 9036 6672 9088 6724
rect 9772 6604 9824 6656
rect 10324 6604 10376 6656
rect 10508 6604 10560 6656
rect 10692 6672 10744 6724
rect 11244 6740 11296 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11336 6672 11388 6724
rect 11980 6740 12032 6792
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 12256 6808 12308 6860
rect 12348 6783 12400 6792
rect 12348 6749 12357 6783
rect 12357 6749 12391 6783
rect 12391 6749 12400 6783
rect 12348 6740 12400 6749
rect 12440 6740 12492 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 12808 6740 12860 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 14372 6808 14424 6860
rect 15108 6876 15160 6928
rect 15384 6876 15436 6928
rect 15844 6876 15896 6928
rect 16304 6944 16356 6996
rect 17684 6876 17736 6928
rect 17960 6876 18012 6928
rect 18052 6876 18104 6928
rect 13636 6740 13688 6792
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14096 6740 14148 6792
rect 12256 6604 12308 6656
rect 13452 6672 13504 6724
rect 14740 6783 14792 6792
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 15936 6808 15988 6860
rect 15292 6740 15344 6792
rect 16580 6740 16632 6792
rect 17408 6808 17460 6860
rect 18144 6808 18196 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 18972 6919 19024 6928
rect 18972 6885 18981 6919
rect 18981 6885 19015 6919
rect 19015 6885 19024 6919
rect 18972 6876 19024 6885
rect 19524 6944 19576 6996
rect 22100 6944 22152 6996
rect 24400 6876 24452 6928
rect 18420 6851 18472 6860
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 19432 6808 19484 6860
rect 17316 6740 17368 6792
rect 17776 6740 17828 6792
rect 18052 6783 18104 6792
rect 18052 6749 18061 6783
rect 18061 6749 18095 6783
rect 18095 6749 18104 6783
rect 18052 6740 18104 6749
rect 18788 6740 18840 6792
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 19156 6740 19208 6792
rect 21088 6783 21140 6792
rect 21088 6749 21097 6783
rect 21097 6749 21131 6783
rect 21131 6749 21140 6783
rect 21088 6740 21140 6749
rect 14648 6672 14700 6724
rect 13360 6604 13412 6656
rect 13728 6604 13780 6656
rect 13912 6647 13964 6656
rect 13912 6613 13921 6647
rect 13921 6613 13955 6647
rect 13955 6613 13964 6647
rect 13912 6604 13964 6613
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 15016 6672 15068 6724
rect 16488 6672 16540 6724
rect 16948 6715 17000 6724
rect 16948 6681 16957 6715
rect 16957 6681 16991 6715
rect 16991 6681 17000 6715
rect 16948 6672 17000 6681
rect 15292 6604 15344 6656
rect 15568 6604 15620 6656
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 16212 6604 16264 6656
rect 16672 6604 16724 6656
rect 16856 6604 16908 6656
rect 17500 6604 17552 6656
rect 17868 6604 17920 6656
rect 19064 6604 19116 6656
rect 19248 6715 19300 6724
rect 19248 6681 19257 6715
rect 19257 6681 19291 6715
rect 19291 6681 19300 6715
rect 19248 6672 19300 6681
rect 21180 6672 21232 6724
rect 20720 6604 20772 6656
rect 21824 6604 21876 6656
rect 22192 6672 22244 6724
rect 22560 6672 22612 6724
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 1676 6400 1728 6452
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 4712 6400 4764 6452
rect 7288 6400 7340 6452
rect 8668 6400 8720 6452
rect 10416 6400 10468 6452
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 756 6264 808 6316
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 3332 6264 3384 6316
rect 6460 6332 6512 6384
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4252 6264 4304 6316
rect 4344 6264 4396 6316
rect 4896 6264 4948 6316
rect 4068 6196 4120 6248
rect 5632 6264 5684 6316
rect 8300 6264 8352 6316
rect 9496 6264 9548 6316
rect 9772 6264 9824 6316
rect 9864 6264 9916 6316
rect 10048 6264 10100 6316
rect 10324 6264 10376 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 3516 6128 3568 6180
rect 5724 6196 5776 6248
rect 10140 6196 10192 6248
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 4620 6128 4672 6180
rect 4896 6171 4948 6180
rect 4896 6137 4905 6171
rect 4905 6137 4939 6171
rect 4939 6137 4948 6171
rect 4896 6128 4948 6137
rect 4988 6128 5040 6180
rect 5448 6128 5500 6180
rect 7840 6128 7892 6180
rect 10048 6128 10100 6180
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 4712 6060 4764 6112
rect 5540 6060 5592 6112
rect 9588 6060 9640 6112
rect 10692 6128 10744 6180
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 10600 6060 10652 6112
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 11336 6196 11388 6248
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12900 6400 12952 6452
rect 13636 6443 13688 6452
rect 13636 6409 13645 6443
rect 13645 6409 13679 6443
rect 13679 6409 13688 6443
rect 13636 6400 13688 6409
rect 12716 6375 12768 6384
rect 12716 6341 12725 6375
rect 12725 6341 12759 6375
rect 12759 6341 12768 6375
rect 12716 6332 12768 6341
rect 12256 6307 12308 6316
rect 12256 6273 12265 6307
rect 12265 6273 12299 6307
rect 12299 6273 12308 6307
rect 12256 6264 12308 6273
rect 12532 6264 12584 6316
rect 12440 6128 12492 6180
rect 11888 6060 11940 6112
rect 12808 6128 12860 6180
rect 13636 6196 13688 6248
rect 15384 6400 15436 6452
rect 16304 6400 16356 6452
rect 15200 6332 15252 6384
rect 14740 6273 14742 6282
rect 14742 6273 14776 6282
rect 14776 6273 14792 6282
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 14740 6230 14792 6273
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 16396 6332 16448 6384
rect 15660 6264 15712 6273
rect 15200 6196 15252 6248
rect 15292 6196 15344 6248
rect 16212 6264 16264 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 13268 6060 13320 6112
rect 15108 6128 15160 6180
rect 15568 6128 15620 6180
rect 16764 6196 16816 6248
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 17684 6264 17736 6316
rect 18236 6264 18288 6316
rect 16028 6128 16080 6180
rect 19156 6196 19208 6248
rect 19616 6264 19668 6316
rect 19984 6332 20036 6384
rect 20168 6332 20220 6384
rect 20996 6264 21048 6316
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 21824 6375 21876 6384
rect 21824 6341 21833 6375
rect 21833 6341 21867 6375
rect 21867 6341 21876 6375
rect 21824 6332 21876 6341
rect 21916 6375 21968 6384
rect 21916 6341 21925 6375
rect 21925 6341 21959 6375
rect 21959 6341 21968 6375
rect 21916 6332 21968 6341
rect 21548 6196 21600 6248
rect 21640 6196 21692 6248
rect 21916 6196 21968 6248
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 22744 6307 22796 6316
rect 22744 6273 22753 6307
rect 22753 6273 22787 6307
rect 22787 6273 22796 6307
rect 22744 6264 22796 6273
rect 22652 6128 22704 6180
rect 23020 6307 23072 6316
rect 23020 6273 23029 6307
rect 23029 6273 23063 6307
rect 23063 6273 23072 6307
rect 23020 6264 23072 6273
rect 15844 6060 15896 6112
rect 16120 6060 16172 6112
rect 17592 6060 17644 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 18788 6060 18840 6112
rect 21640 6060 21692 6112
rect 22100 6060 22152 6112
rect 23204 6103 23256 6112
rect 23204 6069 23213 6103
rect 23213 6069 23247 6103
rect 23247 6069 23256 6103
rect 23204 6060 23256 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 5632 5856 5684 5908
rect 8300 5856 8352 5908
rect 9036 5856 9088 5908
rect 9588 5899 9640 5908
rect 9588 5865 9597 5899
rect 9597 5865 9631 5899
rect 9631 5865 9640 5899
rect 9588 5856 9640 5865
rect 3976 5788 4028 5840
rect 4804 5788 4856 5840
rect 5448 5788 5500 5840
rect 10324 5856 10376 5908
rect 10784 5856 10836 5908
rect 10140 5788 10192 5840
rect 5632 5720 5684 5772
rect 8852 5720 8904 5772
rect 9680 5720 9732 5772
rect 3976 5652 4028 5704
rect 4620 5652 4672 5704
rect 4160 5584 4212 5636
rect 4988 5652 5040 5704
rect 5264 5652 5316 5704
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 5816 5652 5868 5704
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 9772 5652 9824 5704
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 756 5516 808 5568
rect 4436 5516 4488 5568
rect 4620 5559 4672 5568
rect 4620 5525 4629 5559
rect 4629 5525 4663 5559
rect 4663 5525 4672 5559
rect 4620 5516 4672 5525
rect 6736 5516 6788 5568
rect 8024 5584 8076 5636
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 9680 5516 9732 5568
rect 10140 5584 10192 5636
rect 10416 5652 10468 5704
rect 10876 5720 10928 5772
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 11980 5856 12032 5908
rect 13452 5856 13504 5908
rect 11612 5788 11664 5840
rect 12164 5720 12216 5772
rect 13268 5720 13320 5772
rect 10508 5584 10560 5636
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 13176 5652 13228 5704
rect 13728 5856 13780 5908
rect 13636 5788 13688 5840
rect 14648 5831 14700 5840
rect 14648 5797 14657 5831
rect 14657 5797 14691 5831
rect 14691 5797 14700 5831
rect 14648 5788 14700 5797
rect 15200 5856 15252 5908
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 16856 5856 16908 5908
rect 17408 5856 17460 5908
rect 18328 5856 18380 5908
rect 15384 5788 15436 5840
rect 16488 5788 16540 5840
rect 16764 5788 16816 5840
rect 15844 5720 15896 5772
rect 11244 5584 11296 5636
rect 11336 5584 11388 5636
rect 12440 5584 12492 5636
rect 11060 5516 11112 5568
rect 11796 5516 11848 5568
rect 12992 5584 13044 5636
rect 13544 5584 13596 5636
rect 14004 5652 14056 5704
rect 13912 5584 13964 5636
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 15292 5652 15344 5704
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 13360 5516 13412 5568
rect 15108 5584 15160 5636
rect 15384 5584 15436 5636
rect 16764 5695 16816 5704
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 18236 5788 18288 5840
rect 19524 5856 19576 5908
rect 20536 5899 20588 5908
rect 20536 5865 20545 5899
rect 20545 5865 20579 5899
rect 20579 5865 20588 5899
rect 20536 5856 20588 5865
rect 21640 5788 21692 5840
rect 23204 5788 23256 5840
rect 18972 5720 19024 5772
rect 20628 5720 20680 5772
rect 17960 5652 18012 5704
rect 14372 5516 14424 5568
rect 16120 5516 16172 5568
rect 17224 5584 17276 5636
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 21548 5695 21600 5704
rect 21548 5661 21557 5695
rect 21557 5661 21591 5695
rect 21591 5661 21600 5695
rect 21548 5652 21600 5661
rect 18236 5584 18288 5636
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 3976 5355 4028 5364
rect 3976 5321 3985 5355
rect 3985 5321 4019 5355
rect 4019 5321 4028 5355
rect 3976 5312 4028 5321
rect 572 5176 624 5228
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 6184 5312 6236 5364
rect 6552 5312 6604 5364
rect 7012 5312 7064 5364
rect 7104 5355 7156 5364
rect 7104 5321 7113 5355
rect 7113 5321 7147 5355
rect 7147 5321 7156 5355
rect 7104 5312 7156 5321
rect 3884 5176 3936 5185
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 4620 5176 4672 5228
rect 5356 5176 5408 5228
rect 6828 5287 6880 5296
rect 6828 5253 6863 5287
rect 6863 5253 6880 5287
rect 7472 5312 7524 5364
rect 8024 5312 8076 5364
rect 8576 5312 8628 5364
rect 11152 5312 11204 5364
rect 13452 5312 13504 5364
rect 6828 5244 6880 5253
rect 11336 5244 11388 5296
rect 11612 5244 11664 5296
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 5724 5176 5776 5228
rect 6460 5176 6512 5228
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 7380 5219 7432 5228
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 7840 5176 7892 5228
rect 6184 5108 6236 5160
rect 8208 5176 8260 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8484 5176 8536 5228
rect 8944 5176 8996 5228
rect 11428 5176 11480 5228
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 12440 5244 12492 5296
rect 4804 5040 4856 5092
rect 6552 5040 6604 5092
rect 7748 5040 7800 5092
rect 10784 5108 10836 5160
rect 11060 5108 11112 5160
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 12164 5219 12216 5228
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 14096 5244 14148 5296
rect 15292 5312 15344 5364
rect 15568 5312 15620 5364
rect 15752 5312 15804 5364
rect 16396 5312 16448 5364
rect 15108 5287 15160 5296
rect 15108 5253 15117 5287
rect 15117 5253 15151 5287
rect 15151 5253 15160 5287
rect 15108 5244 15160 5253
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 11796 5108 11848 5160
rect 14004 5176 14056 5228
rect 14648 5176 14700 5228
rect 14832 5176 14884 5228
rect 12256 5040 12308 5092
rect 5908 4972 5960 5024
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 6460 4972 6512 5024
rect 13912 5040 13964 5092
rect 14188 5040 14240 5092
rect 15016 5108 15068 5160
rect 15200 5108 15252 5160
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 16672 5244 16724 5296
rect 17592 5244 17644 5296
rect 15660 5108 15712 5160
rect 15752 5108 15804 5160
rect 17224 5219 17276 5228
rect 17224 5185 17233 5219
rect 17233 5185 17267 5219
rect 17267 5185 17276 5219
rect 17224 5176 17276 5185
rect 17408 5219 17460 5228
rect 17408 5185 17416 5219
rect 17416 5185 17450 5219
rect 17450 5185 17460 5219
rect 17408 5176 17460 5185
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 21088 5312 21140 5364
rect 21640 5312 21692 5364
rect 22468 5312 22520 5364
rect 23020 5312 23072 5364
rect 17960 5244 18012 5296
rect 20168 5287 20220 5296
rect 20168 5253 20177 5287
rect 20177 5253 20211 5287
rect 20211 5253 20220 5287
rect 20168 5244 20220 5253
rect 20812 5244 20864 5296
rect 18420 5176 18472 5228
rect 18880 5176 18932 5228
rect 21180 5176 21232 5228
rect 21272 5176 21324 5228
rect 21640 5219 21692 5228
rect 21640 5185 21649 5219
rect 21649 5185 21683 5219
rect 21683 5185 21692 5219
rect 21640 5176 21692 5185
rect 21824 5219 21876 5228
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 22928 5176 22980 5228
rect 23020 5219 23072 5228
rect 23020 5185 23029 5219
rect 23029 5185 23063 5219
rect 23063 5185 23072 5219
rect 23020 5176 23072 5185
rect 23112 5176 23164 5228
rect 14372 5040 14424 5092
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 20720 5108 20772 5160
rect 13084 4972 13136 5024
rect 13176 5015 13228 5024
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 13544 5015 13596 5024
rect 13544 4981 13553 5015
rect 13553 4981 13587 5015
rect 13587 4981 13596 5015
rect 13544 4972 13596 4981
rect 13820 5015 13872 5024
rect 13820 4981 13829 5015
rect 13829 4981 13863 5015
rect 13863 4981 13872 5015
rect 13820 4972 13872 4981
rect 14004 4972 14056 5024
rect 14648 4972 14700 5024
rect 15200 4972 15252 5024
rect 15384 4972 15436 5024
rect 16672 4972 16724 5024
rect 17040 4972 17092 5024
rect 17684 4972 17736 5024
rect 21732 5108 21784 5160
rect 22008 5040 22060 5092
rect 18972 4972 19024 5024
rect 19248 4972 19300 5024
rect 21916 4972 21968 5024
rect 22376 4972 22428 5024
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 5448 4768 5500 4820
rect 6644 4768 6696 4820
rect 7748 4768 7800 4820
rect 8116 4768 8168 4820
rect 8668 4811 8720 4820
rect 8668 4777 8677 4811
rect 8677 4777 8711 4811
rect 8711 4777 8720 4811
rect 8668 4768 8720 4777
rect 8760 4768 8812 4820
rect 10784 4768 10836 4820
rect 11520 4768 11572 4820
rect 4712 4700 4764 4752
rect 4896 4700 4948 4752
rect 5264 4700 5316 4752
rect 5908 4700 5960 4752
rect 7472 4700 7524 4752
rect 7932 4700 7984 4752
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 6368 4632 6420 4684
rect 11244 4743 11296 4752
rect 11244 4709 11253 4743
rect 11253 4709 11287 4743
rect 11287 4709 11296 4743
rect 11244 4700 11296 4709
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 7104 4564 7156 4616
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 4068 4539 4120 4548
rect 4068 4505 4077 4539
rect 4077 4505 4111 4539
rect 4111 4505 4120 4539
rect 4068 4496 4120 4505
rect 4712 4539 4764 4548
rect 4712 4505 4721 4539
rect 4721 4505 4755 4539
rect 4755 4505 4764 4539
rect 4712 4496 4764 4505
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 7656 4607 7708 4616
rect 7656 4573 7669 4607
rect 7669 4573 7708 4607
rect 7656 4564 7708 4573
rect 7748 4496 7800 4548
rect 8024 4607 8076 4616
rect 8024 4573 8033 4607
rect 8033 4573 8067 4607
rect 8067 4573 8076 4607
rect 8024 4564 8076 4573
rect 8576 4632 8628 4684
rect 11060 4632 11112 4684
rect 11428 4632 11480 4684
rect 9036 4564 9088 4616
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9680 4564 9732 4616
rect 8208 4496 8260 4548
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 12716 4768 12768 4820
rect 12808 4768 12860 4820
rect 14372 4768 14424 4820
rect 13636 4700 13688 4752
rect 14188 4632 14240 4684
rect 11336 4496 11388 4548
rect 12072 4496 12124 4548
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 10876 4428 10928 4480
rect 11152 4428 11204 4480
rect 11888 4428 11940 4480
rect 12164 4471 12216 4480
rect 12164 4437 12173 4471
rect 12173 4437 12207 4471
rect 12207 4437 12216 4471
rect 12164 4428 12216 4437
rect 12440 4607 12492 4616
rect 12440 4573 12450 4607
rect 12450 4573 12484 4607
rect 12484 4573 12492 4607
rect 12440 4564 12492 4573
rect 12808 4607 12860 4616
rect 12808 4573 12822 4607
rect 12822 4573 12856 4607
rect 12856 4573 12860 4607
rect 12808 4564 12860 4573
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 13268 4564 13320 4616
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 13912 4564 13964 4616
rect 14464 4607 14516 4616
rect 14464 4573 14477 4607
rect 14477 4573 14516 4607
rect 14464 4564 14516 4573
rect 12624 4539 12676 4548
rect 12624 4505 12633 4539
rect 12633 4505 12667 4539
rect 12667 4505 12676 4539
rect 12624 4496 12676 4505
rect 15936 4768 15988 4820
rect 16488 4768 16540 4820
rect 16948 4768 17000 4820
rect 20720 4768 20772 4820
rect 21364 4811 21416 4820
rect 21364 4777 21373 4811
rect 21373 4777 21407 4811
rect 21407 4777 21416 4811
rect 21364 4768 21416 4777
rect 14832 4700 14884 4752
rect 16212 4700 16264 4752
rect 16396 4700 16448 4752
rect 18512 4700 18564 4752
rect 15568 4632 15620 4684
rect 22284 4632 22336 4684
rect 14924 4539 14976 4548
rect 14924 4505 14933 4539
rect 14933 4505 14967 4539
rect 14967 4505 14976 4539
rect 14924 4496 14976 4505
rect 12992 4428 13044 4480
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 13268 4428 13320 4437
rect 14096 4428 14148 4480
rect 14832 4428 14884 4480
rect 16028 4564 16080 4616
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 16304 4564 16356 4616
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 16580 4564 16632 4616
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 20536 4564 20588 4616
rect 22560 4564 22612 4616
rect 23112 4564 23164 4616
rect 16764 4496 16816 4548
rect 19248 4539 19300 4548
rect 19248 4505 19257 4539
rect 19257 4505 19291 4539
rect 19291 4505 19300 4539
rect 19248 4496 19300 4505
rect 16304 4428 16356 4480
rect 17132 4428 17184 4480
rect 17500 4428 17552 4480
rect 23204 4471 23256 4480
rect 23204 4437 23213 4471
rect 23213 4437 23247 4471
rect 23247 4437 23256 4471
rect 23204 4428 23256 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4804 4224 4856 4276
rect 4620 4156 4672 4208
rect 4712 4156 4764 4208
rect 6460 4224 6512 4276
rect 7748 4224 7800 4276
rect 8392 4224 8444 4276
rect 12072 4224 12124 4276
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 5264 4088 5316 4140
rect 5632 4199 5684 4208
rect 5632 4165 5641 4199
rect 5641 4165 5675 4199
rect 5675 4165 5684 4199
rect 5632 4156 5684 4165
rect 7472 4088 7524 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 9036 4199 9088 4208
rect 9036 4165 9045 4199
rect 9045 4165 9079 4199
rect 9079 4165 9088 4199
rect 9036 4156 9088 4165
rect 10876 4199 10928 4208
rect 10876 4165 10885 4199
rect 10885 4165 10919 4199
rect 10919 4165 10928 4199
rect 10876 4156 10928 4165
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 8300 3952 8352 4004
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 8760 4088 8812 4140
rect 9220 4088 9272 4140
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 11336 4156 11388 4208
rect 11520 4199 11572 4208
rect 11520 4165 11529 4199
rect 11529 4165 11563 4199
rect 11563 4165 11572 4199
rect 11520 4156 11572 4165
rect 13268 4224 13320 4276
rect 14188 4224 14240 4276
rect 15016 4224 15068 4276
rect 15292 4224 15344 4276
rect 17040 4224 17092 4276
rect 15660 4156 15712 4208
rect 8576 3952 8628 4004
rect 9036 3884 9088 3936
rect 9312 3952 9364 4004
rect 11336 4020 11388 4072
rect 11520 3952 11572 4004
rect 12256 4020 12308 4072
rect 13452 4088 13504 4140
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 13636 4131 13688 4140
rect 13636 4097 13645 4131
rect 13645 4097 13679 4131
rect 13679 4097 13688 4131
rect 13636 4088 13688 4097
rect 13820 4088 13872 4140
rect 14188 4088 14240 4140
rect 14464 4088 14516 4140
rect 10416 3884 10468 3936
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 11428 3884 11480 3936
rect 11888 3995 11940 4004
rect 11888 3961 11897 3995
rect 11897 3961 11931 3995
rect 11931 3961 11940 3995
rect 11888 3952 11940 3961
rect 12624 3952 12676 4004
rect 12992 3995 13044 4004
rect 12992 3961 13001 3995
rect 13001 3961 13035 3995
rect 13035 3961 13044 3995
rect 12992 3952 13044 3961
rect 13176 3952 13228 4004
rect 15844 4131 15896 4140
rect 15844 4097 15853 4131
rect 15853 4097 15887 4131
rect 15887 4097 15896 4131
rect 15844 4088 15896 4097
rect 16212 4156 16264 4208
rect 19708 4156 19760 4208
rect 21364 4224 21416 4276
rect 11980 3884 12032 3936
rect 12256 3884 12308 3936
rect 12532 3884 12584 3936
rect 14464 3927 14516 3936
rect 14464 3893 14473 3927
rect 14473 3893 14507 3927
rect 14507 3893 14516 3927
rect 14464 3884 14516 3893
rect 14648 3884 14700 3936
rect 15476 4020 15528 4072
rect 15568 4020 15620 4072
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 16212 4063 16264 4072
rect 16212 4029 16221 4063
rect 16221 4029 16255 4063
rect 16255 4029 16264 4063
rect 16212 4020 16264 4029
rect 16396 4020 16448 4072
rect 16764 4088 16816 4140
rect 17224 4088 17276 4140
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 17132 4020 17184 4072
rect 19156 4088 19208 4140
rect 22284 4156 22336 4208
rect 22376 4156 22428 4208
rect 15292 3995 15344 4004
rect 15292 3961 15301 3995
rect 15301 3961 15335 3995
rect 15335 3961 15344 3995
rect 15292 3952 15344 3961
rect 15384 3952 15436 4004
rect 18420 4020 18472 4072
rect 18512 4020 18564 4072
rect 19616 3995 19668 4004
rect 19616 3961 19625 3995
rect 19625 3961 19659 3995
rect 19659 3961 19668 3995
rect 19616 3952 19668 3961
rect 15936 3884 15988 3936
rect 16120 3884 16172 3936
rect 20260 3927 20312 3936
rect 20260 3893 20269 3927
rect 20269 3893 20303 3927
rect 20303 3893 20312 3927
rect 20260 3884 20312 3893
rect 20628 4020 20680 4072
rect 20812 4020 20864 4072
rect 21180 4131 21232 4140
rect 21180 4097 21189 4131
rect 21189 4097 21223 4131
rect 21223 4097 21232 4131
rect 21180 4088 21232 4097
rect 20536 3952 20588 4004
rect 21364 4131 21416 4140
rect 21364 4097 21378 4131
rect 21378 4097 21412 4131
rect 21412 4097 21416 4131
rect 21364 4088 21416 4097
rect 22652 4131 22704 4140
rect 22652 4097 22661 4131
rect 22661 4097 22695 4131
rect 22695 4097 22704 4131
rect 22652 4088 22704 4097
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 22192 4020 22244 4072
rect 22284 3995 22336 4004
rect 22284 3961 22293 3995
rect 22293 3961 22327 3995
rect 22327 3961 22336 3995
rect 22284 3952 22336 3961
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 8024 3680 8076 3732
rect 10048 3680 10100 3732
rect 10232 3723 10284 3732
rect 10232 3689 10241 3723
rect 10241 3689 10275 3723
rect 10275 3689 10284 3723
rect 10232 3680 10284 3689
rect 7196 3612 7248 3664
rect 7380 3544 7432 3596
rect 7380 3451 7432 3460
rect 7380 3417 7389 3451
rect 7389 3417 7423 3451
rect 7423 3417 7432 3451
rect 7380 3408 7432 3417
rect 8116 3476 8168 3528
rect 10324 3544 10376 3596
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 8668 3476 8720 3528
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9404 3476 9456 3528
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 10876 3680 10928 3732
rect 11152 3680 11204 3732
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 11612 3680 11664 3732
rect 12624 3680 12676 3732
rect 12992 3680 13044 3732
rect 13084 3680 13136 3732
rect 13544 3680 13596 3732
rect 13820 3680 13872 3732
rect 11612 3544 11664 3596
rect 11704 3544 11756 3596
rect 11060 3476 11112 3528
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 7472 3340 7524 3392
rect 7656 3340 7708 3392
rect 10416 3451 10468 3460
rect 10416 3417 10425 3451
rect 10425 3417 10459 3451
rect 10459 3417 10468 3451
rect 10416 3408 10468 3417
rect 11520 3451 11572 3460
rect 11520 3417 11529 3451
rect 11529 3417 11563 3451
rect 11563 3417 11572 3451
rect 11520 3408 11572 3417
rect 11888 3476 11940 3528
rect 12256 3476 12308 3528
rect 12348 3476 12400 3528
rect 12532 3476 12584 3528
rect 13084 3544 13136 3596
rect 13452 3587 13504 3596
rect 13452 3553 13461 3587
rect 13461 3553 13495 3587
rect 13495 3553 13504 3587
rect 13452 3544 13504 3553
rect 12992 3476 13044 3528
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 20076 3680 20128 3732
rect 20168 3680 20220 3732
rect 20904 3680 20956 3732
rect 21824 3680 21876 3732
rect 14832 3612 14884 3664
rect 15200 3612 15252 3664
rect 15568 3612 15620 3664
rect 16488 3612 16540 3664
rect 17224 3612 17276 3664
rect 15016 3544 15068 3596
rect 13544 3476 13596 3485
rect 12164 3408 12216 3460
rect 14648 3476 14700 3528
rect 15200 3476 15252 3528
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 15476 3519 15528 3528
rect 15476 3485 15485 3519
rect 15485 3485 15519 3519
rect 15519 3485 15528 3519
rect 15476 3476 15528 3485
rect 16304 3476 16356 3528
rect 16488 3519 16540 3528
rect 16488 3485 16497 3519
rect 16497 3485 16531 3519
rect 16531 3485 16540 3519
rect 16488 3476 16540 3485
rect 17776 3544 17828 3596
rect 16764 3519 16816 3528
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 16948 3476 17000 3528
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 19340 3476 19392 3528
rect 20076 3544 20128 3596
rect 21180 3544 21232 3596
rect 21364 3476 21416 3528
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 9680 3383 9732 3392
rect 9680 3349 9689 3383
rect 9689 3349 9723 3383
rect 9723 3349 9732 3383
rect 9680 3340 9732 3349
rect 11152 3340 11204 3392
rect 11612 3340 11664 3392
rect 12348 3340 12400 3392
rect 12716 3340 12768 3392
rect 12992 3340 13044 3392
rect 13820 3340 13872 3392
rect 13912 3340 13964 3392
rect 14280 3340 14332 3392
rect 17040 3408 17092 3460
rect 19892 3408 19944 3460
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14464 3340 14516 3349
rect 14740 3340 14792 3392
rect 16120 3383 16172 3392
rect 16120 3349 16129 3383
rect 16129 3349 16163 3383
rect 16163 3349 16172 3383
rect 16120 3340 16172 3349
rect 17592 3340 17644 3392
rect 18972 3340 19024 3392
rect 19524 3340 19576 3392
rect 20536 3340 20588 3392
rect 20720 3340 20772 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 6828 3136 6880 3188
rect 7012 3136 7064 3188
rect 7380 3136 7432 3188
rect 7564 3136 7616 3188
rect 9680 3136 9732 3188
rect 7656 3111 7708 3120
rect 7656 3077 7665 3111
rect 7665 3077 7699 3111
rect 7699 3077 7708 3111
rect 7656 3068 7708 3077
rect 9404 3111 9456 3120
rect 9404 3077 9413 3111
rect 9413 3077 9447 3111
rect 9447 3077 9456 3111
rect 9404 3068 9456 3077
rect 10048 3136 10100 3188
rect 10692 3136 10744 3188
rect 10876 3136 10928 3188
rect 12164 3179 12216 3188
rect 12164 3145 12173 3179
rect 12173 3145 12207 3179
rect 12207 3145 12216 3179
rect 12164 3136 12216 3145
rect 12256 3136 12308 3188
rect 12624 3136 12676 3188
rect 12808 3136 12860 3188
rect 13268 3179 13320 3188
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 14464 3136 14516 3188
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 7288 3000 7340 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 8116 2932 8168 2984
rect 8208 2932 8260 2984
rect 8852 3000 8904 3052
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 11244 3068 11296 3120
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 11060 3000 11112 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 8576 2932 8628 2941
rect 7012 2864 7064 2916
rect 10600 2932 10652 2984
rect 10968 2932 11020 2984
rect 11888 2932 11940 2984
rect 12256 3000 12308 3052
rect 12440 3000 12492 3052
rect 12716 3000 12768 3052
rect 13544 3068 13596 3120
rect 15384 3136 15436 3188
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 18420 3136 18472 3188
rect 19248 3136 19300 3188
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 15476 3068 15528 3120
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 18972 3068 19024 3120
rect 12072 2932 12124 2984
rect 756 2796 808 2848
rect 7288 2796 7340 2848
rect 8852 2796 8904 2848
rect 9128 2796 9180 2848
rect 10784 2796 10836 2848
rect 10968 2796 11020 2848
rect 11244 2796 11296 2848
rect 11336 2796 11388 2848
rect 12164 2796 12216 2848
rect 12532 2796 12584 2848
rect 12992 2796 13044 2848
rect 13728 2796 13780 2848
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 19248 3043 19300 3052
rect 19248 3009 19257 3043
rect 19257 3009 19291 3043
rect 19291 3009 19300 3043
rect 19248 3000 19300 3009
rect 17132 2975 17184 2984
rect 17132 2941 17141 2975
rect 17141 2941 17175 2975
rect 17175 2941 17184 2975
rect 17132 2932 17184 2941
rect 18512 2932 18564 2984
rect 19984 3068 20036 3120
rect 22008 3136 22060 3188
rect 22836 3136 22888 3188
rect 23020 3136 23072 3188
rect 21824 3068 21876 3120
rect 20628 3000 20680 3052
rect 22376 3043 22428 3052
rect 22376 3009 22385 3043
rect 22385 3009 22419 3043
rect 22419 3009 22428 3043
rect 22376 3000 22428 3009
rect 23388 3068 23440 3120
rect 22100 2932 22152 2984
rect 14188 2796 14240 2848
rect 19340 2864 19392 2916
rect 16580 2796 16632 2848
rect 17408 2796 17460 2848
rect 19616 2796 19668 2848
rect 19708 2839 19760 2848
rect 19708 2805 19717 2839
rect 19717 2805 19751 2839
rect 19751 2805 19760 2839
rect 19708 2796 19760 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 4620 2592 4672 2644
rect 5632 2592 5684 2644
rect 7380 2592 7432 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 8392 2524 8444 2576
rect 8760 2567 8812 2576
rect 8760 2533 8769 2567
rect 8769 2533 8803 2567
rect 8803 2533 8812 2567
rect 8760 2524 8812 2533
rect 10968 2592 11020 2644
rect 6828 2499 6880 2508
rect 6828 2465 6837 2499
rect 6837 2465 6871 2499
rect 6871 2465 6880 2499
rect 6828 2456 6880 2465
rect 3884 2388 3936 2440
rect 4528 2388 4580 2440
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5816 2388 5868 2440
rect 7840 2456 7892 2508
rect 11796 2524 11848 2576
rect 12992 2524 13044 2576
rect 13820 2592 13872 2644
rect 16488 2592 16540 2644
rect 16580 2592 16632 2644
rect 17224 2592 17276 2644
rect 19248 2592 19300 2644
rect 23296 2635 23348 2644
rect 23296 2601 23305 2635
rect 23305 2601 23339 2635
rect 23339 2601 23348 2635
rect 23296 2592 23348 2601
rect 17868 2524 17920 2576
rect 19432 2524 19484 2576
rect 22928 2567 22980 2576
rect 22928 2533 22937 2567
rect 22937 2533 22971 2567
rect 22971 2533 22980 2567
rect 22928 2524 22980 2533
rect 7288 2431 7340 2440
rect 7288 2397 7297 2431
rect 7297 2397 7331 2431
rect 7331 2397 7340 2431
rect 7288 2388 7340 2397
rect 7748 2388 7800 2440
rect 9956 2456 10008 2508
rect 7104 2320 7156 2372
rect 8024 2320 8076 2372
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 10968 2388 11020 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 10508 2363 10560 2372
rect 10508 2329 10517 2363
rect 10517 2329 10551 2363
rect 10551 2329 10560 2363
rect 10508 2320 10560 2329
rect 12164 2388 12216 2440
rect 12348 2388 12400 2440
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13084 2320 13136 2372
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 11060 2295 11112 2304
rect 11060 2261 11069 2295
rect 11069 2261 11103 2295
rect 11103 2261 11112 2295
rect 11060 2252 11112 2261
rect 11336 2295 11388 2304
rect 11336 2261 11345 2295
rect 11345 2261 11379 2295
rect 11379 2261 11388 2295
rect 11336 2252 11388 2261
rect 12164 2295 12216 2304
rect 12164 2261 12173 2295
rect 12173 2261 12207 2295
rect 12207 2261 12216 2295
rect 12164 2252 12216 2261
rect 12624 2252 12676 2304
rect 12716 2295 12768 2304
rect 12716 2261 12725 2295
rect 12725 2261 12759 2295
rect 12759 2261 12768 2295
rect 12716 2252 12768 2261
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 14280 2388 14332 2440
rect 17868 2388 17920 2440
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 18972 2431 19024 2440
rect 18972 2397 18981 2431
rect 18981 2397 19015 2431
rect 19015 2397 19024 2431
rect 18972 2388 19024 2397
rect 19340 2456 19392 2508
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 19984 2456 20036 2508
rect 22376 2456 22428 2508
rect 22468 2456 22520 2508
rect 15752 2320 15804 2372
rect 17132 2320 17184 2372
rect 17224 2320 17276 2372
rect 20260 2388 20312 2440
rect 22836 2431 22888 2440
rect 22836 2397 22845 2431
rect 22845 2397 22879 2431
rect 22879 2397 22888 2431
rect 22836 2388 22888 2397
rect 19524 2252 19576 2304
rect 19708 2363 19760 2372
rect 19708 2329 19717 2363
rect 19717 2329 19751 2363
rect 19751 2329 19760 2363
rect 19708 2320 19760 2329
rect 21640 2363 21692 2372
rect 21640 2329 21649 2363
rect 21649 2329 21683 2363
rect 21683 2329 21692 2363
rect 21640 2320 21692 2329
rect 21732 2320 21784 2372
rect 22284 2252 22336 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 11152 2048 11204 2100
rect 16764 2048 16816 2100
rect 11704 1980 11756 2032
rect 14740 1980 14792 2032
rect 10876 1912 10928 1964
rect 19708 1912 19760 1964
rect 10048 1844 10100 1896
rect 14924 1844 14976 1896
rect 9496 1776 9548 1828
rect 16672 1776 16724 1828
rect 13084 1708 13136 1760
rect 19616 1708 19668 1760
rect 8024 1640 8076 1692
rect 12716 1640 12768 1692
rect 14832 1640 14884 1692
rect 14096 1572 14148 1624
rect 15476 1572 15528 1624
rect 11244 1300 11296 1352
rect 18696 1300 18748 1352
rect 11060 1232 11112 1284
rect 17408 1232 17460 1284
rect 12164 1164 12216 1216
rect 16120 1164 16172 1216
rect 10232 1096 10284 1148
rect 18052 1096 18104 1148
rect 11336 1028 11388 1080
rect 16764 1028 16816 1080
rect 12992 960 13044 1012
rect 15476 960 15528 1012
rect 9956 620 10008 672
rect 21916 620 21968 672
rect 10508 76 10560 128
rect 19340 76 19392 128
<< metal2 >>
rect 9034 13270 9090 13370
rect 9678 13270 9734 13370
rect 10966 13270 11022 13370
rect 11610 13270 11666 13370
rect 12254 13270 12310 13370
rect 12898 13270 12954 13370
rect 13542 13270 13598 13370
rect 14186 13270 14242 13370
rect 14830 13270 14886 13370
rect 15474 13270 15530 13370
rect 16118 13270 16174 13370
rect 16212 13320 16264 13326
rect 1306 10976 1362 10985
rect 1306 10911 1362 10920
rect 1320 10606 1348 10911
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 9048 10674 9076 13270
rect 9692 10810 9720 13270
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 10980 10674 11008 13270
rect 11624 10810 11652 13270
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 12268 10674 12296 13270
rect 12912 10674 12940 13270
rect 13556 10810 13584 13270
rect 14200 11014 14228 13270
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14844 10810 14872 13270
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15028 10674 15056 10950
rect 15488 10810 15516 13270
rect 16132 11234 16160 13270
rect 16762 13270 16818 13370
rect 17406 13270 17462 13370
rect 18050 13270 18106 13370
rect 18694 13270 18750 13370
rect 19338 13270 19394 13370
rect 19982 13274 20038 13370
rect 20088 13306 20300 13334
rect 20088 13274 20116 13306
rect 19982 13270 20116 13274
rect 16212 13262 16264 13268
rect 16040 11206 16160 11234
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15842 10704 15898 10713
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 388 10464 440 10470
rect 388 10406 440 10412
rect 400 10305 428 10406
rect 386 10296 442 10305
rect 1964 10266 1992 10610
rect 386 10231 442 10240
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 3344 10062 3372 10610
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 10266 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 388 9920 440 9926
rect 388 9862 440 9868
rect 400 9625 428 9862
rect 1688 9722 1716 9998
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 386 9616 442 9625
rect 386 9551 442 9560
rect 3344 8974 3372 9998
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9722 4568 9862
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4632 9586 4660 9930
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3240 8968 3292 8974
rect 3332 8968 3384 8974
rect 3240 8910 3292 8916
rect 3330 8936 3332 8945
rect 3384 8936 3386 8945
rect 3252 8634 3280 8910
rect 3330 8871 3386 8880
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3804 8634 3832 8842
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3804 8090 3832 8570
rect 4080 8566 4108 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8634 4200 8774
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 388 7880 440 7886
rect 388 7822 440 7828
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 400 7585 428 7822
rect 386 7576 442 7585
rect 386 7511 442 7520
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 204 7200 256 7206
rect 204 7142 256 7148
rect 216 6905 244 7142
rect 202 6896 258 6905
rect 202 6831 258 6840
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1596 6458 1624 6734
rect 1688 6458 1716 7346
rect 1964 7002 1992 7822
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1964 6866 1992 6938
rect 3344 6934 3372 7958
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3332 6928 3384 6934
rect 3332 6870 3384 6876
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 3344 6798 3372 6870
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 2148 6322 2176 6598
rect 3068 6361 3096 6598
rect 3054 6352 3110 6361
rect 756 6316 808 6322
rect 756 6258 808 6264
rect 2136 6316 2188 6322
rect 3344 6322 3372 6734
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3054 6287 3110 6296
rect 3332 6316 3384 6322
rect 2136 6258 2188 6264
rect 3332 6258 3384 6264
rect 768 6225 796 6258
rect 754 6216 810 6225
rect 3528 6186 3556 6598
rect 3804 6361 3832 7822
rect 3896 7750 3924 8434
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8090 4660 9522
rect 4724 9450 4752 10610
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4816 9704 4844 10542
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5172 9988 5224 9994
rect 5224 9948 5304 9976
rect 5172 9930 5224 9936
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4816 9676 4936 9704
rect 4908 9674 4936 9676
rect 4908 9654 5120 9674
rect 4908 9648 5132 9654
rect 4908 9646 5080 9648
rect 5080 9590 5132 9596
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 8974 5028 9318
rect 5092 9042 5120 9590
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8616 4844 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4816 8588 5028 8616
rect 5000 8498 5028 8588
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7342 3924 7686
rect 4068 7472 4120 7478
rect 4172 7426 4200 7822
rect 4120 7420 4200 7426
rect 4068 7414 4200 7420
rect 4080 7398 4200 7414
rect 4344 7404 4396 7410
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3790 6352 3846 6361
rect 3790 6287 3846 6296
rect 754 6151 810 6160
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 756 5568 808 5574
rect 754 5536 756 5545
rect 808 5536 810 5545
rect 754 5471 810 5480
rect 3896 5234 3924 7278
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6662 4016 7142
rect 4080 6984 4108 7398
rect 4344 7346 4396 7352
rect 4356 7206 4384 7346
rect 4448 7206 4476 7890
rect 4620 7880 4672 7886
rect 4618 7848 4620 7857
rect 4672 7848 4674 7857
rect 4618 7783 4674 7792
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4252 6996 4304 7002
rect 4080 6956 4200 6984
rect 4172 6866 4200 6956
rect 4252 6938 4304 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4172 6474 4200 6802
rect 4080 6458 4200 6474
rect 4068 6452 4200 6458
rect 4120 6446 4200 6452
rect 4068 6394 4120 6400
rect 4264 6322 4292 6938
rect 4632 6916 4660 7414
rect 4540 6888 4660 6916
rect 4540 6730 4568 6888
rect 4724 6798 4752 7754
rect 4816 7546 4844 8434
rect 4908 8294 4936 8434
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 5276 7857 5304 9948
rect 5368 9586 5396 10066
rect 5460 10062 5488 10474
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 5828 10062 5856 10406
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5368 9110 5396 9522
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5368 8634 5396 9046
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 8430 5396 8570
rect 5460 8566 5488 9998
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9722 5764 9862
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 8090 5396 8366
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5262 7848 5318 7857
rect 5262 7783 5318 7792
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 5264 7472 5316 7478
rect 5184 7432 5264 7460
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6322 4384 6598
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 3988 5846 4016 6258
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4080 5794 4108 6190
rect 4540 6118 4568 6666
rect 4632 6186 4660 6666
rect 4724 6458 4752 6734
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4080 5766 4200 5794
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3988 5370 4016 5646
rect 4172 5642 4200 5766
rect 4632 5710 4660 6122
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3988 5273 4016 5306
rect 3974 5264 4030 5273
rect 572 5228 624 5234
rect 572 5170 624 5176
rect 3884 5228 3936 5234
rect 4172 5234 4200 5578
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4448 5234 4476 5510
rect 4632 5234 4660 5510
rect 3974 5199 4030 5208
rect 4160 5228 4212 5234
rect 3884 5170 3936 5176
rect 4160 5170 4212 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 584 4865 612 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 570 4856 626 4865
rect 4214 4859 4522 4868
rect 570 4791 626 4800
rect 4724 4758 4752 6054
rect 4816 5846 4844 7142
rect 5184 6730 5212 7432
rect 5264 7414 5316 7420
rect 5368 7274 5396 7890
rect 5460 7290 5488 8230
rect 5552 8106 5580 8910
rect 5644 8838 5672 9454
rect 5828 9450 5856 9522
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5644 8498 5672 8774
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5736 8378 5764 8910
rect 5644 8350 5764 8378
rect 5644 8294 5672 8350
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5552 8078 5764 8106
rect 5828 8090 5856 9386
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5920 8974 5948 9114
rect 5908 8968 5960 8974
rect 6012 8945 6040 9658
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6104 8974 6132 9318
rect 6092 8968 6144 8974
rect 5908 8910 5960 8916
rect 5998 8936 6054 8945
rect 6092 8910 6144 8916
rect 6196 8906 6224 9930
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 5998 8871 6054 8880
rect 6184 8900 6236 8906
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5356 7268 5408 7274
rect 5460 7262 5580 7290
rect 5356 7210 5408 7216
rect 5276 6934 5304 7210
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5276 6798 5304 6870
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5552 6644 5580 7262
rect 5460 6616 5580 6644
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 6186 4936 6258
rect 5460 6186 5488 6616
rect 5644 6322 5672 7958
rect 5736 7002 5764 8078
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4908 5692 4936 6122
rect 5000 5710 5028 6122
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 4816 5664 4936 5692
rect 4988 5704 5040 5710
rect 4816 5352 4844 5664
rect 4988 5646 5040 5652
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4816 5324 4936 5352
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4724 4554 4752 4694
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4080 4146 4108 4490
rect 4724 4214 4752 4490
rect 4816 4282 4844 5034
rect 4908 4758 4936 5324
rect 5276 5250 5304 5646
rect 5354 5536 5410 5545
rect 5354 5471 5410 5480
rect 5184 5222 5304 5250
rect 5368 5234 5396 5471
rect 5356 5228 5408 5234
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 5184 4690 5212 5222
rect 5356 5170 5408 5176
rect 5460 5114 5488 5782
rect 5552 5710 5580 6054
rect 5644 5953 5672 6258
rect 5736 6254 5764 6734
rect 5828 6662 5856 7210
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5630 5944 5686 5953
rect 5630 5879 5632 5888
rect 5684 5879 5686 5888
rect 5632 5850 5684 5856
rect 5644 5778 5672 5850
rect 5632 5772 5684 5778
rect 5684 5732 5764 5760
rect 5632 5714 5684 5720
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5234 5580 5646
rect 5736 5234 5764 5732
rect 5828 5710 5856 6598
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5920 5273 5948 8298
rect 6012 6662 6040 8871
rect 6184 8842 6236 8848
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6104 7886 6132 8298
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6196 7546 6224 7754
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7478 6316 9046
rect 6380 8974 6408 9318
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6472 8022 6500 8434
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6460 7404 6512 7410
rect 6380 7364 6460 7392
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 7206 6132 7278
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6934 6132 7142
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6196 5370 6224 6734
rect 6380 6730 6408 7364
rect 6460 7346 6512 7352
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6472 6390 6500 6870
rect 6564 6798 6592 10202
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9586 6776 9862
rect 6840 9722 6868 9998
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6840 9586 6868 9658
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 6840 9178 6868 9386
rect 6932 9178 6960 9930
rect 7024 9722 7052 10066
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7012 9580 7064 9586
rect 7116 9568 7144 9998
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7064 9540 7144 9568
rect 7012 9522 7064 9528
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7300 9042 7328 9318
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6656 7818 6684 8434
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6840 7886 6868 8026
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6748 7546 6776 7822
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6458 5400 6514 5409
rect 6184 5364 6236 5370
rect 6458 5335 6514 5344
rect 6552 5364 6604 5370
rect 6184 5306 6236 5312
rect 5906 5264 5962 5273
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5724 5228 5776 5234
rect 6472 5234 6500 5335
rect 6552 5306 6604 5312
rect 5906 5199 5962 5208
rect 6460 5228 6512 5234
rect 5724 5170 5776 5176
rect 6460 5170 6512 5176
rect 5644 5114 5672 5170
rect 5460 5086 5672 5114
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 5460 4826 5488 5086
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5630 4856 5686 4865
rect 5448 4820 5500 4826
rect 5630 4791 5686 4800
rect 5448 4762 5500 4768
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 4593 5212 4626
rect 5170 4584 5226 4593
rect 5170 4519 5226 4528
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3505 4660 4150
rect 5276 4146 5304 4694
rect 5644 4214 5672 4791
rect 5920 4758 5948 4966
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6012 4622 6040 4966
rect 6196 4622 6224 5102
rect 6564 5098 6592 5306
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6380 4690 6408 4966
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6472 4282 6500 4966
rect 6656 4826 6684 7346
rect 6748 7274 6776 7346
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6736 5568 6788 5574
rect 7024 5545 7052 8502
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 6736 5510 6788 5516
rect 7010 5536 7066 5545
rect 6748 5284 6776 5510
rect 7010 5471 7066 5480
rect 7024 5370 7052 5471
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 6828 5296 6880 5302
rect 6748 5256 6828 5284
rect 6828 5238 6880 5244
rect 7010 5264 7066 5273
rect 7010 5199 7012 5208
rect 7064 5199 7066 5208
rect 7012 5170 7064 5176
rect 7010 5128 7066 5137
rect 7010 5063 7066 5072
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4618 3496 4674 3505
rect 4618 3431 4674 3440
rect 756 2848 808 2854
rect 754 2816 756 2825
rect 808 2816 810 2825
rect 754 2751 810 2760
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 3431
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5644 2650 5672 4150
rect 7024 3194 7052 5063
rect 7116 4622 7144 5306
rect 7208 5137 7236 8026
rect 7484 7818 7512 9862
rect 7668 9654 7696 9862
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7760 9042 7788 10066
rect 9324 10062 9352 10406
rect 9968 10266 9996 10610
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 11624 10130 11652 10406
rect 12084 10266 12112 10474
rect 12728 10470 12756 10610
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12452 10130 12480 10406
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10508 10056 10560 10062
rect 11428 10056 11480 10062
rect 10508 9998 10560 10004
rect 10690 10024 10746 10033
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8312 9058 8340 9522
rect 8496 9178 8524 9658
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 7748 9036 7800 9042
rect 8312 9030 8524 9058
rect 7748 8978 7800 8984
rect 7760 8634 7788 8978
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7300 5681 7328 6394
rect 7286 5672 7342 5681
rect 7286 5607 7342 5616
rect 7300 5234 7328 5607
rect 7392 5273 7420 6938
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7378 5264 7434 5273
rect 7288 5228 7340 5234
rect 7484 5234 7512 5306
rect 7378 5199 7380 5208
rect 7288 5170 7340 5176
rect 7432 5199 7434 5208
rect 7472 5228 7524 5234
rect 7380 5170 7432 5176
rect 7472 5170 7524 5176
rect 7194 5128 7250 5137
rect 7194 5063 7250 5072
rect 7194 4992 7250 5001
rect 7194 4927 7250 4936
rect 7208 4622 7236 4927
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7208 3670 7236 4558
rect 7392 3720 7420 5170
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7484 4622 7512 4694
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7300 3692 7420 3720
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6840 2514 6868 3130
rect 7024 3058 7052 3130
rect 7300 3058 7328 3692
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7392 3466 7420 3538
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7484 3398 7512 4082
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7392 3058 7420 3130
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7024 2922 7052 2994
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7300 2854 7328 2994
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7300 2446 7328 2790
rect 7392 2650 7420 2994
rect 7484 2650 7512 3334
rect 7576 3194 7604 7822
rect 7760 7002 7788 8230
rect 8036 7886 8064 8842
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8220 7818 8248 8298
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8220 7342 8248 7754
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7668 4622 7696 5646
rect 7760 5098 7788 6938
rect 7944 6934 7972 7278
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6186 7880 6598
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7944 5710 7972 6870
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7838 5400 7894 5409
rect 7838 5335 7894 5344
rect 7852 5234 7880 5335
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7760 4826 7788 5034
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7944 4758 7972 5646
rect 8036 5642 8064 6734
rect 8312 6322 8340 8910
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7274 8432 7754
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8496 6089 8524 9030
rect 8680 8838 8708 9522
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8668 8832 8720 8838
rect 8720 8792 8800 8820
rect 8668 8774 8720 8780
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8588 7886 8616 8230
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8482 6080 8538 6089
rect 8482 6015 8538 6024
rect 8496 5930 8524 6015
rect 8312 5914 8524 5930
rect 8300 5908 8524 5914
rect 8352 5902 8524 5908
rect 8300 5850 8352 5856
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8036 5370 8064 5578
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8206 5264 8262 5273
rect 8206 5199 8208 5208
rect 8260 5199 8262 5208
rect 8208 5170 8260 5176
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 7932 4752 7984 4758
rect 7838 4720 7894 4729
rect 7932 4694 7984 4700
rect 7838 4655 7894 4664
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7760 4282 7788 4490
rect 7852 4486 7880 4655
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7656 3392 7708 3398
rect 7760 3380 7788 4082
rect 8036 4049 8064 4558
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 8036 3738 8064 3975
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8128 3618 8156 4762
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8220 4146 8248 4490
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8312 4010 8340 5646
rect 8496 5234 8524 5902
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8404 4282 8432 5170
rect 8588 4842 8616 5306
rect 8496 4814 8616 4842
rect 8680 4826 8708 6394
rect 8772 5001 8800 8792
rect 8864 8566 8892 9046
rect 8956 9042 8984 9522
rect 9232 9217 9260 9522
rect 9218 9208 9274 9217
rect 9218 9143 9274 9152
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8864 7449 8892 7958
rect 8956 7818 8984 8366
rect 9048 8090 9076 8910
rect 9140 8838 9168 8910
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9232 8548 9260 9143
rect 9324 9110 9352 9998
rect 9600 9178 9628 9998
rect 9772 9920 9824 9926
rect 9770 9888 9772 9897
rect 9824 9888 9826 9897
rect 9770 9823 9826 9832
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9140 8520 9260 8548
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9034 7984 9090 7993
rect 9034 7919 9090 7928
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8850 7440 8906 7449
rect 8850 7375 8906 7384
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8864 6798 8892 7210
rect 9048 7206 9076 7919
rect 9140 7886 9168 8520
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7342 9168 7822
rect 9232 7546 9260 7890
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9324 7410 9352 9046
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8362 9444 8910
rect 9600 8498 9628 8978
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9416 8072 9444 8298
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9496 8084 9548 8090
rect 9416 8044 9496 8072
rect 9496 8026 9548 8032
rect 9600 7993 9628 8230
rect 9586 7984 9642 7993
rect 9586 7919 9642 7928
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9402 7440 9458 7449
rect 9312 7404 9364 7410
rect 9402 7375 9404 7384
rect 9312 7346 9364 7352
rect 9456 7375 9458 7384
rect 9404 7346 9456 7352
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9600 6798 9628 7686
rect 9692 7342 9720 8502
rect 9784 8430 9812 9823
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9876 8634 9904 9590
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 8864 5778 8892 6734
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9048 5914 9076 6666
rect 9784 6662 9812 8366
rect 9968 8362 9996 9318
rect 10060 9081 10088 9318
rect 10046 9072 10102 9081
rect 10046 9007 10102 9016
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7546 9904 7822
rect 10060 7818 10088 8026
rect 10152 7993 10180 9998
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10244 8974 10272 9590
rect 10428 9586 10456 9998
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10428 9058 10456 9522
rect 10520 9178 10548 9998
rect 11428 9998 11480 10004
rect 10690 9959 10692 9968
rect 10744 9959 10746 9968
rect 10692 9930 10744 9936
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 10612 9586 10640 9862
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10428 9030 10548 9058
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10324 8016 10376 8022
rect 10138 7984 10194 7993
rect 10324 7958 10376 7964
rect 10138 7919 10194 7928
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9968 7426 9996 7754
rect 10060 7721 10088 7754
rect 10046 7712 10102 7721
rect 10046 7647 10102 7656
rect 9876 7398 9996 7426
rect 9876 7002 9904 7398
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9772 6656 9824 6662
rect 9494 6624 9550 6633
rect 9772 6598 9824 6604
rect 9494 6559 9550 6568
rect 9508 6322 9536 6559
rect 9784 6322 9812 6598
rect 9876 6322 9904 6734
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5914 9628 6054
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9692 5574 9720 5714
rect 9784 5710 9812 6258
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9864 5704 9916 5710
rect 9968 5692 9996 6938
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6322 10088 6802
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10060 6186 10088 6258
rect 10152 6254 10180 7919
rect 10336 7886 10364 7958
rect 10324 7880 10376 7886
rect 10244 7840 10324 7868
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9916 5664 9996 5692
rect 10048 5704 10100 5710
rect 9864 5646 9916 5652
rect 10048 5646 10100 5652
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8758 4992 8814 5001
rect 8758 4927 8814 4936
rect 8772 4826 8800 4927
rect 8668 4820 8720 4826
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8496 4146 8524 4814
rect 8668 4762 8720 4768
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8588 4010 8616 4626
rect 8772 4146 8800 4762
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 7708 3352 7788 3380
rect 8036 3590 8156 3618
rect 7656 3334 7708 3340
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7576 3097 7604 3130
rect 7668 3126 7696 3334
rect 8036 3176 8064 3590
rect 8956 3534 8984 5170
rect 9218 4720 9274 4729
rect 9218 4655 9274 4664
rect 9232 4622 9260 4655
rect 9692 4622 9720 5510
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9048 4214 9076 4558
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8116 3528 8168 3534
rect 8484 3528 8536 3534
rect 8168 3488 8484 3516
rect 8116 3470 8168 3476
rect 8668 3528 8720 3534
rect 8536 3488 8668 3516
rect 8484 3470 8536 3476
rect 8668 3470 8720 3476
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 7852 3148 8248 3176
rect 7656 3120 7708 3126
rect 7562 3088 7618 3097
rect 7656 3062 7708 3068
rect 7562 3023 7618 3032
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7852 2514 7880 3148
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 3896 100 3924 2382
rect 4540 100 4568 2382
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1306 5304 2382
rect 5184 1278 5304 1306
rect 5184 100 5212 1278
rect 5828 100 5856 2382
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7116 100 7144 2314
rect 7760 100 7788 2382
rect 8036 2378 8064 2994
rect 8220 2990 8248 3148
rect 8574 3088 8630 3097
rect 8392 3052 8444 3058
rect 8574 3023 8630 3032
rect 8852 3052 8904 3058
rect 8392 2994 8444 3000
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8128 2650 8156 2926
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8404 2582 8432 2994
rect 8588 2990 8616 3023
rect 8852 2994 8904 3000
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8864 2854 8892 2994
rect 8852 2848 8904 2854
rect 9048 2836 9076 3878
rect 9232 3777 9260 4082
rect 9310 4040 9366 4049
rect 9310 3975 9312 3984
rect 9364 3975 9366 3984
rect 9312 3946 9364 3952
rect 9218 3768 9274 3777
rect 9218 3703 9274 3712
rect 9232 3534 9260 3703
rect 9416 3534 9444 4082
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9416 3126 9444 3470
rect 9692 3398 9720 4082
rect 9862 3768 9918 3777
rect 10060 3738 10088 5646
rect 10152 5642 10180 5782
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10138 5536 10194 5545
rect 10138 5471 10194 5480
rect 9862 3703 9918 3712
rect 10048 3732 10100 3738
rect 9876 3534 9904 3703
rect 10048 3674 10100 3680
rect 10046 3632 10102 3641
rect 10046 3567 10102 3576
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 3194 9720 3334
rect 10060 3194 10088 3567
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 10060 3058 10088 3130
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9128 2848 9180 2854
rect 9048 2808 9128 2836
rect 8852 2790 8904 2796
rect 9128 2790 9180 2796
rect 8758 2680 8814 2689
rect 8758 2615 8814 2624
rect 8772 2582 8800 2615
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 9968 2514 9996 2994
rect 10152 2689 10180 5471
rect 10244 3738 10272 7840
rect 10324 7822 10376 7828
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10336 6934 10364 7346
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6322 10364 6598
rect 10428 6458 10456 8910
rect 10520 7342 10548 9030
rect 10598 8936 10654 8945
rect 10598 8871 10654 8880
rect 10612 8566 10640 8871
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10612 7954 10640 8502
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10704 6866 10732 9454
rect 10796 8974 10824 9522
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10782 8120 10838 8129
rect 10782 8055 10838 8064
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10508 6656 10560 6662
rect 10560 6616 10640 6644
rect 10508 6598 10560 6604
rect 10506 6488 10562 6497
rect 10416 6452 10468 6458
rect 10612 6458 10640 6616
rect 10506 6423 10562 6432
rect 10600 6452 10652 6458
rect 10416 6394 10468 6400
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10520 6202 10548 6423
rect 10600 6394 10652 6400
rect 10428 6174 10548 6202
rect 10704 6186 10732 6666
rect 10796 6338 10824 8055
rect 10888 6497 10916 8910
rect 11348 8838 11376 9862
rect 11440 9450 11468 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11532 9042 11560 9658
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11164 8430 11192 8774
rect 11440 8498 11468 8774
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 10966 7440 11022 7449
rect 10966 7375 11022 7384
rect 10874 6488 10930 6497
rect 10874 6423 10930 6432
rect 10796 6310 10916 6338
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10692 6180 10744 6186
rect 10324 5908 10376 5914
rect 10428 5896 10456 6174
rect 10692 6122 10744 6128
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10376 5868 10456 5896
rect 10324 5850 10376 5856
rect 10428 5710 10456 5868
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10520 5642 10548 6054
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10612 4026 10640 6054
rect 10796 5914 10824 6190
rect 10888 5953 10916 6310
rect 10874 5944 10930 5953
rect 10784 5908 10836 5914
rect 10874 5879 10930 5888
rect 10784 5850 10836 5856
rect 10690 5808 10746 5817
rect 10888 5778 10916 5879
rect 10690 5743 10746 5752
rect 10876 5772 10928 5778
rect 10336 3998 10640 4026
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10336 3602 10364 3998
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10428 3466 10456 3878
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10704 3194 10732 5743
rect 10876 5714 10928 5720
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10796 5166 10824 5646
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10796 4826 10824 5102
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10888 4214 10916 4422
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10888 3194 10916 3674
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10336 2825 10364 2994
rect 10600 2984 10652 2990
rect 10796 2961 10824 2994
rect 10600 2926 10652 2932
rect 10782 2952 10838 2961
rect 10612 2836 10640 2926
rect 10782 2887 10838 2896
rect 10784 2848 10836 2854
rect 10322 2816 10378 2825
rect 10612 2808 10784 2836
rect 10784 2790 10836 2796
rect 10322 2751 10378 2760
rect 10138 2680 10194 2689
rect 10138 2615 10194 2624
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 8036 1698 8064 2314
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 1873 8524 2246
rect 8482 1864 8538 1873
rect 9508 1834 9536 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 8482 1799 8538 1808
rect 9496 1828 9548 1834
rect 9496 1770 9548 1776
rect 8024 1692 8076 1698
rect 8024 1634 8076 1640
rect 9692 105 9720 2246
rect 9968 678 9996 2246
rect 10060 1902 10088 2382
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10048 1896 10100 1902
rect 10048 1838 10100 1844
rect 10244 1154 10272 2246
rect 10232 1148 10284 1154
rect 10232 1090 10284 1096
rect 9956 672 10008 678
rect 9956 614 10008 620
rect 10520 134 10548 2314
rect 10888 1970 10916 2994
rect 10980 2990 11008 7375
rect 11058 6624 11114 6633
rect 11058 6559 11114 6568
rect 11072 6254 11100 6559
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11060 5568 11112 5574
rect 11164 5556 11192 8366
rect 11532 6798 11560 8978
rect 11624 8922 11652 10066
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9178 11744 9862
rect 12084 9489 12112 9998
rect 12176 9722 12204 9998
rect 12636 9994 12664 10202
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12256 9512 12308 9518
rect 12070 9480 12126 9489
rect 12256 9454 12308 9460
rect 12070 9415 12126 9424
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11808 9042 11836 9318
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 12268 8974 12296 9454
rect 11888 8968 11940 8974
rect 11624 8894 11836 8922
rect 12072 8968 12124 8974
rect 11888 8910 11940 8916
rect 12070 8936 12072 8945
rect 12256 8968 12308 8974
rect 12124 8936 12126 8945
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7410 11744 7890
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 7041 11744 7346
rect 11702 7032 11758 7041
rect 11702 6967 11758 6976
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11256 5642 11284 6734
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11348 6497 11376 6666
rect 11334 6488 11390 6497
rect 11334 6423 11390 6432
rect 11426 6352 11482 6361
rect 11426 6287 11482 6296
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 5642 11376 6190
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11112 5528 11192 5556
rect 11060 5510 11112 5516
rect 11072 5166 11100 5510
rect 11256 5409 11284 5578
rect 11242 5400 11298 5409
rect 11152 5364 11204 5370
rect 11242 5335 11298 5344
rect 11152 5306 11204 5312
rect 11164 5273 11192 5306
rect 11336 5296 11388 5302
rect 11150 5264 11206 5273
rect 11336 5238 11388 5244
rect 11150 5199 11206 5208
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11072 3534 11100 4626
rect 11164 4622 11192 5199
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 3738 11192 4422
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11256 3534 11284 4694
rect 11348 4554 11376 5238
rect 11440 5234 11468 6287
rect 11624 5846 11652 6802
rect 11808 6322 11836 8894
rect 11900 8838 11928 8910
rect 12256 8910 12308 8916
rect 12070 8871 12126 8880
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11900 7886 11928 8230
rect 11992 7886 12020 8230
rect 12084 8090 12112 8774
rect 12268 8566 12296 8910
rect 12360 8838 12388 9590
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11532 4826 11560 5170
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 4214 11376 4490
rect 11440 4298 11468 4626
rect 11532 4622 11560 4762
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11440 4270 11560 4298
rect 11532 4214 11560 4270
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11348 3942 11376 4014
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3738 11468 3878
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11072 3058 11100 3470
rect 11164 3398 11192 3470
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 11164 2938 11192 3334
rect 11256 3126 11284 3470
rect 11532 3466 11560 3946
rect 11624 3738 11652 5238
rect 11716 4185 11744 6258
rect 11808 5574 11836 6258
rect 11900 6118 11928 7822
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11980 6792 12032 6798
rect 12084 6780 12112 7686
rect 12176 7478 12204 8366
rect 12452 7698 12480 9658
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 8634 12572 9454
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8022 12572 8434
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12544 7818 12572 7958
rect 12636 7886 12664 9930
rect 12728 9761 12756 10406
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12714 9752 12770 9761
rect 12820 9722 12848 9930
rect 12912 9722 12940 10134
rect 13096 10062 13124 10542
rect 13924 10266 13952 10610
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14660 10198 14688 10610
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14832 10056 14884 10062
rect 15016 10056 15068 10062
rect 14884 10016 15016 10044
rect 14832 9998 14884 10004
rect 15016 9998 15068 10004
rect 13096 9722 13124 9998
rect 12714 9687 12770 9696
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9110 12848 9522
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12820 8838 12848 9046
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12912 8129 12940 9386
rect 13740 9353 13768 9998
rect 14200 9897 14228 9998
rect 14280 9920 14332 9926
rect 14186 9888 14242 9897
rect 14280 9862 14332 9868
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14186 9823 14242 9832
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14002 9480 14058 9489
rect 14002 9415 14004 9424
rect 14056 9415 14058 9424
rect 14004 9386 14056 9392
rect 13820 9376 13872 9382
rect 13726 9344 13782 9353
rect 13820 9318 13872 9324
rect 13726 9279 13782 9288
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 12898 8120 12954 8129
rect 12898 8055 12954 8064
rect 12624 7880 12676 7886
rect 12808 7880 12860 7886
rect 12676 7840 12808 7868
rect 12624 7822 12676 7828
rect 12808 7822 12860 7828
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12808 7744 12860 7750
rect 12452 7670 12664 7698
rect 12808 7686 12860 7692
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12176 6866 12204 7278
rect 12544 7177 12572 7346
rect 12530 7168 12586 7177
rect 12530 7103 12586 7112
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12032 6752 12112 6780
rect 12268 6746 12296 6802
rect 11980 6734 12032 6740
rect 12176 6718 12296 6746
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11900 5216 11928 6054
rect 11992 5914 12020 6258
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12176 5778 12204 6718
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6322 12296 6598
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12162 5672 12218 5681
rect 12162 5607 12218 5616
rect 12176 5234 12204 5607
rect 11980 5228 12032 5234
rect 11900 5188 11980 5216
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11702 4176 11758 4185
rect 11702 4111 11758 4120
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11624 3602 11652 3674
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11624 3398 11652 3538
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11716 3058 11744 3538
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11164 2910 11376 2938
rect 11348 2854 11376 2910
rect 10968 2848 11020 2854
rect 11244 2848 11296 2854
rect 11020 2808 11100 2836
rect 10968 2790 11020 2796
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10980 2446 11008 2586
rect 11072 2553 11100 2808
rect 11244 2790 11296 2796
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11058 2544 11114 2553
rect 11058 2479 11114 2488
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 10876 1964 10928 1970
rect 10876 1906 10928 1912
rect 11072 1290 11100 2246
rect 11164 2106 11192 2382
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11256 1358 11284 2790
rect 11808 2582 11836 5102
rect 11900 4486 11928 5188
rect 11980 5170 12032 5176
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12268 4729 12296 5034
rect 12254 4720 12310 4729
rect 12254 4655 12310 4664
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 12084 4282 12112 4490
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12254 4448 12310 4457
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12176 4049 12204 4422
rect 12254 4383 12310 4392
rect 12268 4078 12296 4383
rect 12360 4128 12388 6734
rect 12452 6186 12480 6734
rect 12544 6322 12572 7103
rect 12636 6798 12664 7670
rect 12714 6896 12770 6905
rect 12714 6831 12770 6840
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12622 6624 12678 6633
rect 12622 6559 12678 6568
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12440 5636 12492 5642
rect 12636 5624 12664 6559
rect 12728 6390 12756 6831
rect 12820 6798 12848 7686
rect 13004 7478 13032 8842
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13096 8022 13124 8774
rect 13188 8090 13216 8774
rect 13280 8498 13308 8842
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12900 7336 12952 7342
rect 12898 7304 12900 7313
rect 12952 7304 12954 7313
rect 12898 7239 12954 7248
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12900 6792 12952 6798
rect 13004 6780 13032 7414
rect 12952 6752 13032 6780
rect 13174 6760 13230 6769
rect 12900 6734 12952 6740
rect 12806 6488 12862 6497
rect 12912 6458 12940 6734
rect 13174 6695 13230 6704
rect 13082 6488 13138 6497
rect 12806 6423 12862 6432
rect 12900 6452 12952 6458
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12820 6186 12848 6423
rect 13082 6423 13138 6432
rect 12900 6394 12952 6400
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12492 5596 12664 5624
rect 12440 5578 12492 5584
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12452 4865 12480 5238
rect 12438 4856 12494 4865
rect 12820 4826 12848 5646
rect 12992 5636 13044 5642
rect 13096 5624 13124 6423
rect 13188 5710 13216 6695
rect 13280 6202 13308 8434
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 7886 13400 8230
rect 13556 7886 13584 9114
rect 13832 9042 13860 9318
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 8634 13676 8774
rect 14108 8634 14136 9522
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14186 8528 14242 8537
rect 14186 8463 14242 8472
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13372 6769 13400 6938
rect 13358 6760 13414 6769
rect 13358 6695 13414 6704
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13360 6656 13412 6662
rect 13358 6624 13360 6633
rect 13412 6624 13414 6633
rect 13358 6559 13414 6568
rect 13280 6174 13400 6202
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13280 5778 13308 6054
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13176 5704 13228 5710
rect 13372 5658 13400 6174
rect 13464 5914 13492 6666
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13556 5760 13584 7822
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13648 6458 13676 6734
rect 13740 6662 13768 6734
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13636 6248 13688 6254
rect 13740 6225 13768 6598
rect 13636 6190 13688 6196
rect 13726 6216 13782 6225
rect 13648 5846 13676 6190
rect 13726 6151 13782 6160
rect 13726 5944 13782 5953
rect 13726 5879 13728 5888
rect 13780 5879 13782 5888
rect 13728 5850 13780 5856
rect 13636 5840 13688 5846
rect 13636 5782 13688 5788
rect 13176 5646 13228 5652
rect 13044 5596 13124 5624
rect 13280 5630 13400 5658
rect 13464 5732 13584 5760
rect 12992 5578 13044 5584
rect 13004 5545 13032 5578
rect 12990 5536 13046 5545
rect 12990 5471 13046 5480
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 12438 4791 12494 4800
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12438 4720 12494 4729
rect 12438 4655 12494 4664
rect 12452 4622 12480 4655
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12452 4321 12480 4558
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12438 4312 12494 4321
rect 12438 4247 12494 4256
rect 12530 4176 12586 4185
rect 12360 4100 12480 4128
rect 12530 4111 12586 4120
rect 12256 4072 12308 4078
rect 12162 4040 12218 4049
rect 11888 4004 11940 4010
rect 12256 4014 12308 4020
rect 12162 3975 12218 3984
rect 11888 3946 11940 3952
rect 11900 3913 11928 3946
rect 11980 3936 12032 3942
rect 11886 3904 11942 3913
rect 11980 3878 12032 3884
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12346 3904 12402 3913
rect 11886 3839 11942 3848
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 2990 11928 3470
rect 11992 3074 12020 3878
rect 12268 3534 12296 3878
rect 12346 3839 12402 3848
rect 12360 3534 12388 3839
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12176 3194 12204 3402
rect 12268 3194 12296 3470
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12254 3088 12310 3097
rect 11992 3046 12204 3074
rect 11888 2984 11940 2990
rect 12072 2984 12124 2990
rect 11940 2944 12072 2972
rect 11888 2926 11940 2932
rect 12072 2926 12124 2932
rect 12176 2854 12204 3046
rect 12254 3023 12256 3032
rect 12308 3023 12310 3032
rect 12256 2994 12308 3000
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 12176 2446 12204 2790
rect 12360 2446 12388 3334
rect 12452 3058 12480 4100
rect 12544 3942 12572 4111
rect 12636 4010 12664 4490
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12636 3738 12664 3946
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12544 2854 12572 3470
rect 12728 3398 12756 4762
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12624 3188 12676 3194
rect 12728 3176 12756 3334
rect 12820 3194 12848 4558
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12898 4312 12954 4321
rect 12898 4247 12954 4256
rect 12912 3516 12940 4247
rect 13004 4010 13032 4422
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 13096 3738 13124 4966
rect 13188 4729 13216 4966
rect 13174 4720 13230 4729
rect 13174 4655 13230 4664
rect 13280 4622 13308 5630
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5234 13400 5510
rect 13464 5370 13492 5732
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13176 4616 13228 4622
rect 13268 4616 13320 4622
rect 13176 4558 13228 4564
rect 13266 4584 13268 4593
rect 13320 4584 13322 4593
rect 13188 4457 13216 4558
rect 13266 4519 13322 4528
rect 13268 4480 13320 4486
rect 13174 4448 13230 4457
rect 13268 4422 13320 4428
rect 13174 4383 13230 4392
rect 13280 4282 13308 4422
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13372 4185 13400 5170
rect 13358 4176 13414 4185
rect 13464 4146 13492 5306
rect 13556 5030 13584 5578
rect 13726 5536 13782 5545
rect 13726 5471 13782 5480
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4457 13584 4966
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13542 4448 13598 4457
rect 13542 4383 13598 4392
rect 13648 4146 13676 4694
rect 13740 4622 13768 5471
rect 13832 5030 13860 8230
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 6798 14136 7210
rect 14096 6792 14148 6798
rect 14016 6752 14096 6780
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13924 5953 13952 6598
rect 13910 5944 13966 5953
rect 13910 5879 13966 5888
rect 13910 5808 13966 5817
rect 13910 5743 13966 5752
rect 13924 5642 13952 5743
rect 14016 5710 14044 6752
rect 14096 6734 14148 6740
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 14108 5409 14136 6190
rect 14094 5400 14150 5409
rect 14094 5335 14150 5344
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13832 4146 13860 4966
rect 13924 4622 13952 5034
rect 14016 5030 14044 5170
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 4865 14044 4966
rect 14002 4856 14058 4865
rect 14002 4791 14058 4800
rect 14108 4808 14136 5238
rect 14200 5098 14228 8463
rect 14292 7886 14320 9862
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14476 8634 14504 9522
rect 14568 8974 14596 9862
rect 15212 9674 15240 10678
rect 15842 10639 15898 10648
rect 15476 10464 15528 10470
rect 15396 10424 15476 10452
rect 15396 10130 15424 10424
rect 15476 10406 15528 10412
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15568 9920 15620 9926
rect 15752 9920 15804 9926
rect 15568 9862 15620 9868
rect 15672 9880 15752 9908
rect 15108 9648 15160 9654
rect 15212 9646 15424 9674
rect 15160 9596 15240 9602
rect 15108 9590 15240 9596
rect 15120 9574 15240 9590
rect 15014 9208 15070 9217
rect 15014 9143 15016 9152
rect 15068 9143 15070 9152
rect 15108 9172 15160 9178
rect 15016 9114 15068 9120
rect 15108 9114 15160 9120
rect 14556 8968 14608 8974
rect 14924 8968 14976 8974
rect 14556 8910 14608 8916
rect 14844 8928 14924 8956
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14384 8022 14412 8434
rect 14372 8016 14424 8022
rect 14476 7993 14504 8570
rect 14568 8430 14596 8910
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14660 8566 14688 8774
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14372 7958 14424 7964
rect 14462 7984 14518 7993
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14384 7818 14412 7958
rect 14462 7919 14518 7928
rect 14476 7886 14504 7919
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14384 7546 14412 7754
rect 14568 7732 14596 8366
rect 14660 7886 14688 8502
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14476 7704 14596 7732
rect 14844 7721 14872 8928
rect 14924 8910 14976 8916
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14830 7712 14886 7721
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14372 6860 14424 6866
rect 14292 6820 14372 6848
rect 14292 5273 14320 6820
rect 14372 6802 14424 6808
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 5681 14412 6598
rect 14370 5672 14426 5681
rect 14370 5607 14426 5616
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14278 5264 14334 5273
rect 14278 5199 14334 5208
rect 14384 5098 14412 5510
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14476 5012 14504 7704
rect 14830 7647 14886 7656
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14752 6798 14780 7346
rect 14740 6792 14792 6798
rect 14646 6760 14702 6769
rect 14740 6734 14792 6740
rect 14646 6695 14648 6704
rect 14700 6695 14702 6704
rect 14648 6666 14700 6672
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 5710 14596 6598
rect 14740 6282 14792 6288
rect 14740 6224 14792 6230
rect 14648 5840 14700 5846
rect 14752 5828 14780 6224
rect 14700 5800 14780 5828
rect 14648 5782 14700 5788
rect 14844 5710 14872 7647
rect 14936 7585 14964 8366
rect 14922 7576 14978 7585
rect 14922 7511 14978 7520
rect 15028 7460 15056 9114
rect 15120 8974 15148 9114
rect 15212 9110 15240 9574
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15212 8401 15240 8910
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15198 8392 15254 8401
rect 15304 8362 15332 8434
rect 15198 8327 15254 8336
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15198 8120 15254 8129
rect 15198 8055 15200 8064
rect 15252 8055 15254 8064
rect 15200 8026 15252 8032
rect 15304 7954 15332 8298
rect 15396 8090 15424 9646
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15488 9178 15516 9522
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15580 8974 15608 9862
rect 15672 9586 15700 9880
rect 15752 9862 15804 9868
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 8974 15700 9522
rect 15764 9489 15792 9590
rect 15750 9480 15806 9489
rect 15750 9415 15806 9424
rect 15764 9217 15792 9415
rect 15750 9208 15806 9217
rect 15750 9143 15806 9152
rect 15764 8974 15792 9143
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15580 8809 15608 8910
rect 15566 8800 15622 8809
rect 15566 8735 15622 8744
rect 15580 8498 15608 8735
rect 15672 8566 15700 8910
rect 15856 8634 15884 10639
rect 16040 10538 16068 11206
rect 16118 11112 16174 11121
rect 16118 11047 16174 11056
rect 16132 10810 16160 11047
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16118 9888 16174 9897
rect 16118 9823 16174 9832
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15948 8809 15976 9522
rect 16040 9110 16068 9522
rect 16028 9104 16080 9110
rect 16028 9046 16080 9052
rect 15934 8800 15990 8809
rect 15934 8735 15990 8744
rect 16040 8634 16068 9046
rect 16132 8974 16160 9823
rect 16224 9110 16252 13262
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 9178 16344 9522
rect 16408 9178 16436 10950
rect 16670 10840 16726 10849
rect 16776 10810 16804 13270
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16670 10775 16726 10784
rect 16764 10804 16816 10810
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16500 10266 16528 10610
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16592 10146 16620 10474
rect 16684 10470 16712 10775
rect 16764 10746 16816 10752
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16762 10432 16818 10441
rect 16762 10367 16818 10376
rect 16500 10118 16620 10146
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16500 8974 16528 10118
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16776 9674 16804 10367
rect 16960 10062 16988 11018
rect 17420 10810 17448 13270
rect 17682 12336 17738 12345
rect 17682 12271 17738 12280
rect 17498 10976 17554 10985
rect 17498 10911 17554 10920
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17144 10538 17172 10610
rect 17406 10568 17462 10577
rect 17132 10532 17184 10538
rect 17406 10503 17462 10512
rect 17132 10474 17184 10480
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8974 16620 9318
rect 16684 9178 16712 9658
rect 16776 9646 16988 9674
rect 17328 9654 17356 10134
rect 16776 9586 16804 9646
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16868 9489 16896 9522
rect 16854 9480 16910 9489
rect 16764 9444 16816 9450
rect 16854 9415 16910 9424
rect 16764 9386 16816 9392
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16120 8968 16172 8974
rect 16488 8968 16540 8974
rect 16120 8910 16172 8916
rect 16394 8936 16450 8945
rect 16488 8910 16540 8916
rect 16580 8968 16632 8974
rect 16684 8945 16712 8978
rect 16580 8910 16632 8916
rect 16670 8936 16726 8945
rect 16394 8871 16450 8880
rect 16670 8871 16726 8880
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 14936 7432 15056 7460
rect 14936 6440 14964 7432
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15120 7274 15148 7346
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15014 7168 15070 7177
rect 15014 7103 15070 7112
rect 15028 6730 15056 7103
rect 15120 6934 15148 7210
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 14936 6412 15056 6440
rect 14922 6352 14978 6361
rect 14922 6287 14978 6296
rect 14936 5710 14964 6287
rect 15028 5710 15056 6412
rect 15212 6390 15240 7482
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15304 7041 15332 7346
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15290 7032 15346 7041
rect 15290 6967 15346 6976
rect 15304 6798 15332 6967
rect 15396 6934 15424 7278
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15292 6792 15344 6798
rect 15344 6752 15424 6780
rect 15292 6734 15344 6740
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15304 6338 15332 6598
rect 15396 6458 15424 6752
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15108 6316 15160 6322
rect 15304 6310 15424 6338
rect 15108 6258 15160 6264
rect 15120 6186 15148 6258
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 14556 5704 14608 5710
rect 14832 5704 14884 5710
rect 14608 5664 14780 5692
rect 14556 5646 14608 5652
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14660 5137 14688 5170
rect 14646 5128 14702 5137
rect 14646 5063 14702 5072
rect 14648 5024 14700 5030
rect 14476 4984 14648 5012
rect 14372 4820 14424 4826
rect 14108 4780 14320 4808
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14094 4584 14150 4593
rect 14094 4519 14150 4528
rect 14108 4486 14136 4519
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14200 4282 14228 4626
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 13358 4111 13414 4120
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13820 4140 13872 4146
rect 14188 4140 14240 4146
rect 13872 4100 13952 4128
rect 13820 4082 13872 4088
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13004 3618 13032 3674
rect 13188 3641 13216 3946
rect 13450 3904 13506 3913
rect 13450 3839 13506 3848
rect 13174 3632 13230 3641
rect 13004 3602 13124 3618
rect 13004 3596 13136 3602
rect 13004 3590 13084 3596
rect 13464 3602 13492 3839
rect 13556 3738 13584 4082
rect 13740 3738 13860 3754
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13740 3732 13872 3738
rect 13740 3726 13820 3732
rect 13174 3567 13230 3576
rect 13452 3596 13504 3602
rect 13084 3538 13136 3544
rect 13452 3538 13504 3544
rect 12992 3528 13044 3534
rect 12912 3488 12992 3516
rect 12992 3470 13044 3476
rect 12992 3392 13044 3398
rect 12898 3360 12954 3369
rect 12992 3334 13044 3340
rect 12898 3295 12954 3304
rect 12676 3148 12756 3176
rect 12808 3188 12860 3194
rect 12624 3130 12676 3136
rect 12808 3130 12860 3136
rect 12716 3052 12768 3058
rect 12636 3012 12716 3040
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11244 1352 11296 1358
rect 11244 1294 11296 1300
rect 11060 1284 11112 1290
rect 11060 1226 11112 1232
rect 11348 1086 11376 2246
rect 11716 2038 11744 2382
rect 12636 2310 12664 3012
rect 12716 2994 12768 3000
rect 12912 2446 12940 3295
rect 13004 2854 13032 3334
rect 13096 3058 13124 3538
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13266 3224 13322 3233
rect 13266 3159 13268 3168
rect 13320 3159 13322 3168
rect 13268 3130 13320 3136
rect 13556 3126 13584 3470
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13464 2961 13492 2994
rect 13450 2952 13506 2961
rect 13450 2887 13506 2896
rect 13740 2854 13768 3726
rect 13820 3674 13872 3680
rect 13924 3398 13952 4100
rect 14188 4082 14240 4088
rect 14002 3496 14058 3505
rect 14002 3431 14058 3440
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13832 3058 13860 3334
rect 14016 3058 14044 3431
rect 14200 3097 14228 4082
rect 14292 3505 14320 4780
rect 14372 4762 14424 4768
rect 14278 3496 14334 3505
rect 14278 3431 14334 3440
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14186 3088 14242 3097
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14004 3052 14056 3058
rect 14186 3023 14242 3032
rect 14004 2994 14056 3000
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 12176 1222 12204 2246
rect 12728 1698 12756 2246
rect 12716 1692 12768 1698
rect 12716 1634 12768 1640
rect 12164 1216 12216 1222
rect 12164 1158 12216 1164
rect 11336 1080 11388 1086
rect 11336 1022 11388 1028
rect 13004 1018 13032 2518
rect 13832 2446 13860 2586
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13096 1766 13124 2314
rect 13084 1760 13136 1766
rect 13084 1702 13136 1708
rect 14108 1630 14136 2382
rect 14096 1624 14148 1630
rect 14096 1566 14148 1572
rect 12992 1012 13044 1018
rect 12992 954 13044 960
rect 10508 128 10560 134
rect 3882 0 3938 100
rect 4526 0 4582 100
rect 5170 0 5226 100
rect 5814 0 5870 100
rect 7102 0 7158 100
rect 7746 0 7802 100
rect 9678 96 9734 105
rect 14200 100 14228 2790
rect 14292 2446 14320 3334
rect 14384 3058 14412 4762
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14476 4146 14504 4558
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14464 3936 14516 3942
rect 14462 3904 14464 3913
rect 14516 3904 14518 3913
rect 14462 3839 14518 3848
rect 14464 3392 14516 3398
rect 14568 3380 14596 4984
rect 14648 4966 14700 4972
rect 14752 4593 14780 5664
rect 14832 5646 14884 5652
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14844 5234 14872 5646
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14844 4758 14872 5170
rect 14936 5148 14964 5646
rect 15028 5284 15056 5646
rect 15120 5642 15148 6122
rect 15212 5914 15240 6190
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15304 5710 15332 6190
rect 15396 5846 15424 6310
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15304 5370 15332 5646
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15108 5296 15160 5302
rect 15028 5256 15108 5284
rect 15396 5273 15424 5578
rect 15108 5238 15160 5244
rect 15382 5264 15438 5273
rect 15016 5160 15068 5166
rect 14936 5120 15016 5148
rect 15016 5102 15068 5108
rect 15120 5001 15148 5238
rect 15382 5199 15438 5208
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15290 5128 15346 5137
rect 15212 5030 15240 5102
rect 15290 5063 15346 5072
rect 15200 5024 15252 5030
rect 15106 4992 15162 5001
rect 15200 4966 15252 4972
rect 15106 4927 15162 4936
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14738 4584 14794 4593
rect 14738 4519 14794 4528
rect 14924 4548 14976 4554
rect 14924 4490 14976 4496
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14660 3534 14688 3878
rect 14844 3670 14872 4422
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14516 3352 14596 3380
rect 14740 3392 14792 3398
rect 14464 3334 14516 3340
rect 14740 3334 14792 3340
rect 14476 3194 14504 3334
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 14752 2038 14780 3334
rect 14740 2032 14792 2038
rect 14740 1974 14792 1980
rect 14936 1902 14964 4490
rect 15304 4282 15332 5063
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15016 4276 15068 4282
rect 15016 4218 15068 4224
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15028 3602 15056 4218
rect 15396 4128 15424 4966
rect 15120 4100 15424 4128
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15120 3369 15148 4100
rect 15488 4078 15516 7822
rect 15580 7546 15608 7890
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15672 7478 15700 7890
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 6662 15608 7346
rect 15672 6662 15700 7414
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15568 6180 15620 6186
rect 15568 6122 15620 6128
rect 15580 5370 15608 6122
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15672 5250 15700 6258
rect 15764 5370 15792 7686
rect 15856 7041 15884 8434
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15948 7721 15976 7754
rect 15934 7712 15990 7721
rect 15934 7647 15990 7656
rect 16026 7168 16082 7177
rect 16026 7103 16082 7112
rect 15842 7032 15898 7041
rect 15842 6967 15898 6976
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15856 6118 15884 6870
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15844 6112 15896 6118
rect 15948 6089 15976 6802
rect 16040 6186 16068 7103
rect 16132 6361 16160 7754
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6769 16252 7142
rect 16316 7002 16344 7686
rect 16408 7290 16436 8871
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16500 8129 16528 8434
rect 16580 8424 16632 8430
rect 16578 8392 16580 8401
rect 16632 8392 16634 8401
rect 16578 8327 16634 8336
rect 16672 8288 16724 8294
rect 16578 8256 16634 8265
rect 16672 8230 16724 8236
rect 16578 8191 16634 8200
rect 16486 8120 16542 8129
rect 16486 8055 16542 8064
rect 16592 7886 16620 8191
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16408 7274 16528 7290
rect 16408 7268 16540 7274
rect 16408 7262 16488 7268
rect 16488 7210 16540 7216
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 7041 16436 7142
rect 16394 7032 16450 7041
rect 16304 6996 16356 7002
rect 16394 6967 16450 6976
rect 16304 6938 16356 6944
rect 16592 6905 16620 7346
rect 16302 6896 16358 6905
rect 16302 6831 16358 6840
rect 16578 6896 16634 6905
rect 16578 6831 16634 6840
rect 16210 6760 16266 6769
rect 16210 6695 16266 6704
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16118 6352 16174 6361
rect 16224 6322 16252 6598
rect 16316 6458 16344 6831
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16118 6287 16174 6296
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15844 6054 15896 6060
rect 15934 6080 15990 6089
rect 15934 6015 15990 6024
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15568 5228 15620 5234
rect 15672 5222 15792 5250
rect 15568 5170 15620 5176
rect 15580 4690 15608 5170
rect 15764 5166 15792 5222
rect 15660 5160 15712 5166
rect 15658 5128 15660 5137
rect 15752 5160 15804 5166
rect 15712 5128 15714 5137
rect 15752 5102 15804 5108
rect 15658 5063 15714 5072
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15566 4312 15622 4321
rect 15566 4247 15622 4256
rect 15580 4078 15608 4247
rect 15672 4214 15700 5063
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15212 3534 15240 3606
rect 15304 3534 15332 3946
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15106 3360 15162 3369
rect 15106 3295 15162 3304
rect 15304 2553 15332 3470
rect 15396 3194 15424 3946
rect 15580 3670 15608 4014
rect 15568 3664 15620 3670
rect 15474 3632 15530 3641
rect 15568 3606 15620 3612
rect 15474 3567 15530 3576
rect 15488 3534 15516 3567
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15488 3126 15516 3470
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15290 2544 15346 2553
rect 15290 2479 15346 2488
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 14832 1692 14884 1698
rect 14832 1634 14884 1640
rect 14844 100 14872 1634
rect 15488 1630 15516 3062
rect 15764 2378 15792 5102
rect 15856 4146 15884 5714
rect 15948 5710 15976 6015
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15934 5264 15990 5273
rect 16040 5234 16068 6122
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5710 16160 6054
rect 16224 5710 16252 6258
rect 16408 5914 16436 6326
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16500 5846 16528 6666
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16486 5672 16542 5681
rect 16486 5607 16542 5616
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15934 5199 15936 5208
rect 15988 5199 15990 5208
rect 16028 5228 16080 5234
rect 15936 5170 15988 5176
rect 16028 5170 16080 5176
rect 15948 4826 15976 5170
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16040 4622 16068 5170
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15934 4312 15990 4321
rect 15934 4247 15990 4256
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15948 3942 15976 4247
rect 16028 4072 16080 4078
rect 16132 4060 16160 5510
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16408 4758 16436 5306
rect 16500 4826 16528 5607
rect 16592 5273 16620 6734
rect 16684 6662 16712 8230
rect 16776 7993 16804 9386
rect 16960 9092 16988 9646
rect 17316 9648 17368 9654
rect 17038 9616 17094 9625
rect 17316 9590 17368 9596
rect 17038 9551 17094 9560
rect 17052 9518 17080 9551
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17420 9382 17448 10503
rect 17512 9568 17540 10911
rect 17696 10674 17724 12271
rect 18064 11937 18092 13270
rect 18708 12073 18736 13270
rect 18694 12064 18750 12073
rect 18694 11999 18750 12008
rect 18050 11928 18106 11937
rect 18050 11863 18106 11872
rect 18694 11656 18750 11665
rect 18694 11591 18750 11600
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17788 10266 17816 10610
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17682 9616 17738 9625
rect 17512 9540 17632 9568
rect 17788 9586 17816 9998
rect 17682 9551 17738 9560
rect 17776 9580 17828 9586
rect 17500 9444 17552 9450
rect 17500 9386 17552 9392
rect 17408 9376 17460 9382
rect 17038 9344 17094 9353
rect 17038 9279 17094 9288
rect 17222 9344 17278 9353
rect 17408 9318 17460 9324
rect 17222 9279 17278 9288
rect 17052 9110 17080 9279
rect 16868 9064 16988 9092
rect 17040 9104 17092 9110
rect 16868 8956 16896 9064
rect 17040 9046 17092 9052
rect 17040 8968 17092 8974
rect 16868 8928 16988 8956
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 8566 16896 8774
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16960 8498 16988 8928
rect 17092 8928 17172 8956
rect 17040 8910 17092 8916
rect 17144 8616 17172 8928
rect 17236 8634 17264 9279
rect 17314 9208 17370 9217
rect 17420 9178 17448 9318
rect 17314 9143 17370 9152
rect 17408 9172 17460 9178
rect 17328 9110 17356 9143
rect 17408 9114 17460 9120
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17512 9042 17540 9386
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17604 8974 17632 9540
rect 17696 9217 17724 9551
rect 17880 9568 17908 10678
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 17958 10160 18014 10169
rect 18248 10130 18276 10406
rect 17958 10095 18014 10104
rect 18144 10124 18196 10130
rect 17972 9568 18000 10095
rect 18144 10066 18196 10072
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 9654 18092 9998
rect 18156 9761 18184 10066
rect 18142 9752 18198 9761
rect 18142 9687 18198 9696
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17880 9540 18000 9568
rect 17776 9522 17828 9528
rect 18052 9512 18104 9518
rect 17880 9472 18052 9500
rect 17682 9208 17738 9217
rect 17682 9143 17684 9152
rect 17736 9143 17738 9152
rect 17684 9114 17736 9120
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17052 8588 17172 8616
rect 17224 8628 17276 8634
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 16868 8265 16896 8298
rect 16948 8288 17000 8294
rect 16854 8256 16910 8265
rect 17052 8276 17080 8588
rect 17224 8570 17276 8576
rect 17328 8498 17356 8774
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17132 8492 17184 8498
rect 17316 8492 17368 8498
rect 17184 8452 17264 8480
rect 17132 8434 17184 8440
rect 17000 8248 17080 8276
rect 17130 8256 17186 8265
rect 16948 8230 17000 8236
rect 16854 8191 16910 8200
rect 17130 8191 17186 8200
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16762 7984 16818 7993
rect 16762 7919 16818 7928
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16776 6905 16804 7278
rect 16762 6896 16818 6905
rect 16762 6831 16818 6840
rect 16868 6746 16896 7822
rect 16960 6848 16988 7822
rect 17052 7410 17080 8026
rect 17144 7886 17172 8191
rect 17236 7993 17264 8452
rect 17316 8434 17368 8440
rect 17222 7984 17278 7993
rect 17222 7919 17278 7928
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 6914 17080 7142
rect 17144 6984 17172 7686
rect 17236 7478 17264 7822
rect 17328 7818 17356 8434
rect 17604 8362 17632 8502
rect 17684 8492 17736 8498
rect 17788 8480 17816 9046
rect 17880 8974 17908 9472
rect 18144 9512 18196 9518
rect 18052 9454 18104 9460
rect 18142 9480 18144 9489
rect 18196 9480 18198 9489
rect 18142 9415 18198 9424
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17972 8838 18000 9318
rect 18248 9092 18276 10066
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18340 9110 18368 9930
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18156 9064 18276 9092
rect 18328 9104 18380 9110
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17960 8560 18012 8566
rect 17736 8452 17816 8480
rect 17684 8434 17736 8440
rect 17408 8356 17460 8362
rect 17592 8356 17644 8362
rect 17460 8316 17540 8344
rect 17408 8298 17460 8304
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17314 7712 17370 7721
rect 17314 7647 17370 7656
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17328 7410 17356 7647
rect 17420 7546 17448 7890
rect 17512 7886 17540 8316
rect 17592 8298 17644 8304
rect 17604 8090 17632 8298
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17788 7970 17816 8452
rect 17604 7942 17816 7970
rect 17880 8520 17960 8548
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17512 7410 17540 7822
rect 17604 7721 17632 7942
rect 17764 7880 17816 7886
rect 17696 7840 17764 7868
rect 17590 7712 17646 7721
rect 17590 7647 17646 7656
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17316 7268 17368 7274
rect 17419 7256 17447 7346
rect 17419 7228 17448 7256
rect 17316 7210 17368 7216
rect 17328 7018 17356 7210
rect 17420 7177 17448 7228
rect 17406 7168 17462 7177
rect 17406 7103 17462 7112
rect 17328 6990 17448 7018
rect 17144 6956 17264 6984
rect 17052 6886 17172 6914
rect 16960 6820 17080 6848
rect 16776 6718 16896 6746
rect 16948 6724 17000 6730
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 5302 16712 6598
rect 16776 6254 16804 6718
rect 16948 6666 17000 6672
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 6322 16896 6598
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16868 5914 16896 6258
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16764 5840 16816 5846
rect 16764 5782 16816 5788
rect 16776 5710 16804 5782
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16672 5296 16724 5302
rect 16578 5264 16634 5273
rect 16672 5238 16724 5244
rect 16578 5199 16634 5208
rect 16776 5114 16804 5646
rect 16868 5273 16896 5646
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 16592 5086 16804 5114
rect 16854 5128 16910 5137
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16224 4622 16252 4694
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16224 4214 16252 4558
rect 16316 4486 16344 4558
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16212 4208 16264 4214
rect 16408 4162 16436 4694
rect 16592 4622 16620 5086
rect 16854 5063 16910 5072
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16212 4150 16264 4156
rect 16316 4134 16436 4162
rect 16080 4032 16160 4060
rect 16212 4072 16264 4078
rect 16210 4040 16212 4049
rect 16264 4040 16266 4049
rect 16028 4014 16080 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 16040 3777 16068 4014
rect 16210 3975 16266 3984
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16026 3768 16082 3777
rect 16026 3703 16082 3712
rect 16132 3398 16160 3878
rect 16316 3534 16344 4134
rect 16396 4072 16448 4078
rect 16394 4040 16396 4049
rect 16448 4040 16450 4049
rect 16394 3975 16450 3984
rect 16500 3670 16528 4558
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16500 2650 16528 3470
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 2650 16620 2790
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 16684 1834 16712 4966
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16776 4146 16804 4490
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16764 3528 16816 3534
rect 16868 3516 16896 5063
rect 16960 4826 16988 6666
rect 17052 6322 17080 6820
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17144 5794 17172 6886
rect 17236 6780 17264 6956
rect 17420 6866 17448 6990
rect 17696 6934 17724 7840
rect 17764 7822 17816 7828
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17316 6792 17368 6798
rect 17236 6752 17316 6780
rect 17316 6734 17368 6740
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17052 5766 17172 5794
rect 17052 5137 17080 5766
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17222 5672 17278 5681
rect 17038 5128 17094 5137
rect 17038 5063 17094 5072
rect 17040 5024 17092 5030
rect 17038 4992 17040 5001
rect 17092 4992 17094 5001
rect 17038 4927 17094 4936
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17040 4616 17092 4622
rect 17144 4604 17172 5646
rect 17222 5607 17224 5616
rect 17276 5607 17278 5616
rect 17224 5578 17276 5584
rect 17420 5234 17448 5850
rect 17512 5234 17540 6598
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17604 5710 17632 6054
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17236 4622 17264 5170
rect 17314 4720 17370 4729
rect 17314 4655 17370 4664
rect 17092 4576 17172 4604
rect 17224 4616 17276 4622
rect 17040 4558 17092 4564
rect 17224 4558 17276 4564
rect 17052 4282 17080 4558
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17144 4078 17172 4422
rect 17328 4146 17356 4655
rect 17512 4486 17540 5170
rect 17500 4480 17552 4486
rect 17406 4448 17462 4457
rect 17500 4422 17552 4428
rect 17406 4383 17462 4392
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 16946 3768 17002 3777
rect 16946 3703 17002 3712
rect 16960 3534 16988 3703
rect 17236 3670 17264 4082
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 16816 3488 16896 3516
rect 16948 3528 17000 3534
rect 16764 3470 16816 3476
rect 16948 3470 17000 3476
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16776 2106 16804 3130
rect 17052 3058 17080 3402
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 17144 2378 17172 2926
rect 17420 2854 17448 4383
rect 17604 3398 17632 5238
rect 17696 5030 17724 6258
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17788 3602 17816 6734
rect 17880 6662 17908 8520
rect 17960 8502 18012 8508
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17972 8090 18000 8230
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17958 7984 18014 7993
rect 17958 7919 18014 7928
rect 17972 7886 18000 7919
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17958 7712 18014 7721
rect 17958 7647 18014 7656
rect 17972 6934 18000 7647
rect 18064 7546 18092 8910
rect 18156 8362 18184 9064
rect 18328 9046 18380 9052
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8809 18276 8910
rect 18234 8800 18290 8809
rect 18234 8735 18290 8744
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18248 7993 18276 8230
rect 18234 7984 18290 7993
rect 18234 7919 18290 7928
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18064 6934 18092 7482
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18156 6866 18184 7686
rect 18248 7478 18276 7919
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 6866 18276 7142
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 18064 6361 18092 6734
rect 18050 6352 18106 6361
rect 18248 6322 18276 6802
rect 18050 6287 18106 6296
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17960 5704 18012 5710
rect 17958 5672 17960 5681
rect 18012 5672 18014 5681
rect 17958 5607 18014 5616
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17972 4593 18000 5238
rect 17958 4584 18014 4593
rect 17958 4519 18014 4528
rect 18064 4049 18092 6054
rect 18248 5846 18276 6258
rect 18340 5914 18368 8502
rect 18432 6866 18460 9318
rect 18524 9178 18552 10542
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18616 10062 18644 10474
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18708 9586 18736 11591
rect 19352 10810 19380 13270
rect 19996 13246 20116 13270
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 18800 10062 18828 10610
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 18892 10266 18920 10406
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 18788 10056 18840 10062
rect 19064 10056 19116 10062
rect 18840 10016 19064 10044
rect 18788 9998 18840 10004
rect 19064 9998 19116 10004
rect 19168 9897 19196 10066
rect 19154 9888 19210 9897
rect 19154 9823 19210 9832
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18788 9104 18840 9110
rect 18708 9064 18788 9092
rect 18708 9058 18736 9064
rect 18524 9030 18736 9058
rect 18788 9046 18840 9052
rect 18970 9072 19026 9081
rect 18524 8537 18552 9030
rect 18970 9007 19026 9016
rect 18984 8974 19012 9007
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 18972 8832 19024 8838
rect 18878 8800 18934 8809
rect 18972 8774 19024 8780
rect 18878 8735 18934 8744
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18510 8528 18566 8537
rect 18510 8463 18566 8472
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 8362 18644 8434
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18524 7993 18552 8298
rect 18616 8090 18644 8298
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18510 7984 18566 7993
rect 18510 7919 18566 7928
rect 18708 7886 18736 8570
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18800 7886 18828 8026
rect 18512 7880 18564 7886
rect 18696 7880 18748 7886
rect 18564 7840 18644 7868
rect 18512 7822 18564 7828
rect 18512 7744 18564 7750
rect 18616 7732 18644 7840
rect 18696 7822 18748 7828
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18616 7704 18828 7732
rect 18512 7686 18564 7692
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18524 6361 18552 7686
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18510 6352 18566 6361
rect 18510 6287 18566 6296
rect 18616 6089 18644 7210
rect 18800 6798 18828 7704
rect 18892 7188 18920 8735
rect 18984 8566 19012 8774
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 19076 8090 19104 8910
rect 19168 8090 19196 8910
rect 19260 8838 19288 10406
rect 19536 10062 19564 10474
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19064 7948 19116 7954
rect 19168 7936 19196 8026
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19116 7908 19196 7936
rect 19064 7890 19116 7896
rect 19076 7449 19104 7890
rect 19062 7440 19118 7449
rect 19062 7375 19118 7384
rect 19260 7206 19288 7958
rect 19352 7818 19380 9522
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19248 7200 19300 7206
rect 18892 7160 19104 7188
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18878 6352 18934 6361
rect 18878 6287 18934 6296
rect 18788 6112 18840 6118
rect 18602 6080 18658 6089
rect 18602 6015 18658 6024
rect 18786 6080 18788 6089
rect 18840 6080 18842 6089
rect 18786 6015 18842 6024
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 18892 5710 18920 6287
rect 18984 5778 19012 6870
rect 19076 6798 19104 7160
rect 19248 7142 19300 7148
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19064 6656 19116 6662
rect 19168 6644 19196 6734
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19116 6616 19196 6644
rect 19064 6598 19116 6604
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18236 5636 18288 5642
rect 18236 5578 18288 5584
rect 18142 5400 18198 5409
rect 18142 5335 18198 5344
rect 18156 5166 18184 5335
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18050 4040 18106 4049
rect 18050 3975 18106 3984
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 18248 3233 18276 5578
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18432 4078 18460 5170
rect 18892 5001 18920 5170
rect 18972 5024 19024 5030
rect 18878 4992 18934 5001
rect 18972 4966 19024 4972
rect 18878 4927 18934 4936
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18524 4078 18552 4694
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18234 3224 18290 3233
rect 18234 3159 18290 3168
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17236 2378 17264 2586
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 17880 2446 17908 2518
rect 18432 2446 18460 3130
rect 18524 2990 18552 4014
rect 18984 3534 19012 4966
rect 19076 3913 19104 6598
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19168 4146 19196 6190
rect 19260 5030 19288 6666
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19062 3904 19118 3913
rect 19062 3839 19118 3848
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18984 3126 19012 3334
rect 19260 3194 19288 4490
rect 19352 3534 19380 7754
rect 19444 6866 19472 8910
rect 19536 8022 19564 9998
rect 19720 9178 19748 10610
rect 19798 10296 19854 10305
rect 19798 10231 19854 10240
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19628 7721 19656 8910
rect 19812 8906 19840 10231
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19706 8528 19762 8537
rect 19706 8463 19708 8472
rect 19760 8463 19762 8472
rect 19708 8434 19760 8440
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19812 7857 19840 8366
rect 19798 7848 19854 7857
rect 19798 7783 19854 7792
rect 19614 7712 19670 7721
rect 19614 7647 19670 7656
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19720 7410 19748 7482
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19536 5914 19564 6938
rect 19904 6361 19932 8842
rect 19996 6390 20024 9930
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9586 20208 9862
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20180 8498 20208 9522
rect 20272 8838 20300 13306
rect 20626 13270 20682 13370
rect 21270 13270 21326 13370
rect 21914 13270 21970 13370
rect 22558 13270 22614 13370
rect 23112 13320 23164 13326
rect 20640 11082 20668 13270
rect 21086 12064 21142 12073
rect 21086 11999 21142 12008
rect 20810 11928 20866 11937
rect 20810 11863 20866 11872
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20824 10674 20852 11863
rect 21100 10674 21128 11999
rect 21284 11121 21312 13270
rect 21270 11112 21326 11121
rect 21270 11047 21326 11056
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21468 10674 21496 10950
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21180 10600 21232 10606
rect 21178 10568 21180 10577
rect 21232 10568 21234 10577
rect 21178 10503 21234 10512
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 20640 10130 20668 10406
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 21180 10056 21232 10062
rect 20350 10024 20406 10033
rect 21180 9998 21232 10004
rect 20350 9959 20406 9968
rect 21088 9988 21140 9994
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20364 8498 20392 9959
rect 21088 9930 21140 9936
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20732 9178 20760 9522
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20536 7880 20588 7886
rect 20640 7857 20668 7958
rect 20732 7954 20760 9114
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20902 8664 20958 8673
rect 20902 8599 20958 8608
rect 20916 8566 20944 8599
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 21008 8498 21036 9046
rect 21100 8634 21128 9930
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20720 7948 20772 7954
rect 21008 7936 21036 8434
rect 21008 7908 21128 7936
rect 20720 7890 20772 7896
rect 20536 7822 20588 7828
rect 20626 7848 20682 7857
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 19984 6384 20036 6390
rect 19890 6352 19946 6361
rect 19616 6316 19668 6322
rect 19984 6326 20036 6332
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 19890 6287 19946 6296
rect 19616 6258 19668 6264
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19628 4010 19656 6258
rect 19708 4208 19760 4214
rect 19708 4150 19760 4156
rect 19616 4004 19668 4010
rect 19444 3964 19616 3992
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18524 2446 18552 2926
rect 18984 2446 19012 3062
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19260 2650 19288 2994
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19352 2514 19380 2858
rect 19444 2582 19472 3964
rect 19616 3946 19668 3952
rect 19720 3890 19748 4150
rect 19628 3862 19748 3890
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17224 2372 17276 2378
rect 17224 2314 17276 2320
rect 19536 2310 19564 3334
rect 19628 2854 19656 3862
rect 19892 3460 19944 3466
rect 19892 3402 19944 3408
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19720 2496 19748 2790
rect 19904 2514 19932 3402
rect 19996 3126 20024 6326
rect 20180 5302 20208 6326
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 20180 3738 20208 5238
rect 20456 3992 20484 7142
rect 20548 5914 20576 7822
rect 20626 7783 20682 7792
rect 20640 7392 20668 7783
rect 20732 7546 20760 7890
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20720 7404 20772 7410
rect 20640 7364 20720 7392
rect 20904 7404 20956 7410
rect 20720 7346 20772 7352
rect 20824 7364 20904 7392
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20732 6662 20760 7142
rect 20720 6656 20772 6662
rect 20824 6633 20852 7364
rect 20904 7346 20956 7352
rect 20902 6760 20958 6769
rect 20902 6695 20958 6704
rect 20720 6598 20772 6604
rect 20810 6624 20866 6633
rect 20810 6559 20866 6568
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20548 4622 20576 5850
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20640 4078 20668 5714
rect 20824 5386 20852 6559
rect 20732 5358 20852 5386
rect 20732 5166 20760 5358
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20536 4004 20588 4010
rect 20456 3964 20536 3992
rect 20536 3946 20588 3952
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20088 3602 20116 3674
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 19628 2468 19748 2496
rect 19892 2508 19944 2514
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 16764 2100 16816 2106
rect 16764 2042 16816 2048
rect 16672 1828 16724 1834
rect 16672 1770 16724 1776
rect 19628 1766 19656 2468
rect 19892 2450 19944 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19708 2372 19760 2378
rect 19708 2314 19760 2320
rect 19720 1970 19748 2314
rect 19708 1964 19760 1970
rect 19708 1906 19760 1912
rect 19616 1760 19668 1766
rect 19616 1702 19668 1708
rect 15476 1624 15528 1630
rect 15476 1566 15528 1572
rect 18696 1352 18748 1358
rect 18696 1294 18748 1300
rect 17408 1284 17460 1290
rect 17408 1226 17460 1232
rect 16120 1216 16172 1222
rect 16120 1158 16172 1164
rect 15476 1012 15528 1018
rect 15476 954 15528 960
rect 15488 100 15516 954
rect 16132 100 16160 1158
rect 16764 1080 16816 1086
rect 16764 1022 16816 1028
rect 16776 100 16804 1022
rect 17420 100 17448 1226
rect 18052 1148 18104 1154
rect 18052 1090 18104 1096
rect 18064 100 18092 1090
rect 18708 100 18736 1294
rect 19340 128 19392 134
rect 10508 70 10560 76
rect 9678 31 9734 40
rect 14186 0 14242 100
rect 14830 0 14886 100
rect 15474 0 15530 100
rect 16118 0 16174 100
rect 16762 0 16818 100
rect 17406 0 17462 100
rect 18050 0 18106 100
rect 18694 0 18750 100
rect 19338 76 19340 100
rect 19996 100 20024 2450
rect 20272 2446 20300 3878
rect 20548 3398 20576 3946
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20640 3058 20668 4014
rect 20732 3398 20760 4762
rect 20824 4078 20852 5238
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20916 3738 20944 6695
rect 21008 6322 21036 7754
rect 21100 7750 21128 7908
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7478 21128 7686
rect 21088 7472 21140 7478
rect 21088 7414 21140 7420
rect 21192 7206 21220 9998
rect 21284 9976 21312 10406
rect 21364 9988 21416 9994
rect 21284 9948 21364 9976
rect 21284 9518 21312 9948
rect 21364 9930 21416 9936
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21376 8634 21404 8774
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21284 8401 21312 8502
rect 21270 8392 21326 8401
rect 21270 8327 21326 8336
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 21100 5370 21128 6734
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 21192 5234 21220 6666
rect 21284 5234 21312 8327
rect 21468 7410 21496 10406
rect 21560 10266 21588 10950
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21836 10441 21864 10610
rect 21822 10432 21878 10441
rect 21822 10367 21878 10376
rect 21928 10266 21956 13270
rect 22466 10840 22522 10849
rect 22466 10775 22522 10784
rect 22480 10742 22508 10775
rect 22468 10736 22520 10742
rect 22374 10704 22430 10713
rect 22468 10678 22520 10684
rect 22374 10639 22376 10648
rect 22428 10639 22430 10648
rect 22376 10610 22428 10616
rect 22376 10532 22428 10538
rect 22376 10474 22428 10480
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21560 7546 21588 8434
rect 21652 8129 21680 8502
rect 21744 8498 21772 9318
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21638 8120 21694 8129
rect 21638 8055 21694 8064
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21376 4826 21404 6258
rect 21468 5710 21496 7210
rect 21652 6254 21680 8055
rect 21836 6746 21864 9318
rect 22112 8974 22140 10406
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 21916 8968 21968 8974
rect 22100 8968 22152 8974
rect 21968 8928 22048 8956
rect 21916 8910 21968 8916
rect 21914 8528 21970 8537
rect 21914 8463 21916 8472
rect 21968 8463 21970 8472
rect 21916 8434 21968 8440
rect 21914 7032 21970 7041
rect 21914 6967 21970 6976
rect 21744 6718 21864 6746
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21560 5710 21588 6190
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21652 5846 21680 6054
rect 21640 5840 21692 5846
rect 21640 5782 21692 5788
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21640 5364 21692 5370
rect 21640 5306 21692 5312
rect 21652 5273 21680 5306
rect 21638 5264 21694 5273
rect 21638 5199 21640 5208
rect 21692 5199 21694 5208
rect 21640 5170 21692 5176
rect 21744 5166 21772 6718
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21836 6390 21864 6598
rect 21928 6390 21956 6967
rect 21824 6384 21876 6390
rect 21824 6326 21876 6332
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 21836 5234 21864 6326
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21376 4282 21404 4762
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 21192 3602 21220 4082
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 21376 3534 21404 4082
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 21744 2378 21772 5102
rect 21928 5030 21956 6190
rect 22020 5098 22048 8928
rect 22098 8936 22100 8945
rect 22152 8936 22154 8945
rect 22098 8871 22154 8880
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22112 7002 22140 7346
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22204 6730 22232 8842
rect 22296 8498 22324 9386
rect 22388 9042 22416 10474
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22480 8974 22508 9862
rect 22572 9674 22600 13270
rect 23202 13274 23258 13370
rect 23164 13270 23258 13274
rect 23846 13270 23902 13370
rect 24490 13270 24546 13370
rect 23164 13268 23244 13270
rect 23112 13262 23244 13268
rect 23124 13246 23244 13262
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22664 10538 22692 10950
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22664 10062 22692 10474
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22572 9646 22692 9674
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22296 7478 22324 8026
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22008 5092 22060 5098
rect 22008 5034 22060 5040
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 21836 3126 21864 3674
rect 22020 3194 22048 5034
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21824 3120 21876 3126
rect 21824 3062 21876 3068
rect 22112 2990 22140 6054
rect 22204 4078 22232 6258
rect 22296 4690 22324 7414
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22388 7313 22416 7346
rect 22374 7304 22430 7313
rect 22374 7239 22430 7248
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22388 5030 22416 7142
rect 22572 6914 22600 9522
rect 22664 9382 22692 9646
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22756 8974 22784 10678
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22848 9761 22876 10406
rect 22834 9752 22890 9761
rect 22834 9687 22890 9696
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 8498 22876 8774
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22940 8401 22968 10406
rect 23124 10062 23152 10678
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 22926 8392 22982 8401
rect 22926 8327 22982 8336
rect 23032 8090 23060 9522
rect 23124 9217 23152 9998
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23110 9208 23166 9217
rect 23110 9143 23166 9152
rect 23216 8634 23244 9862
rect 23388 9444 23440 9450
rect 23388 9386 23440 9392
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7410 22692 7686
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22480 6886 22600 6914
rect 22480 5370 22508 6886
rect 22560 6724 22612 6730
rect 22560 6666 22612 6672
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22296 4214 22324 4626
rect 22388 4214 22416 4966
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 21640 2372 21692 2378
rect 21640 2314 21692 2320
rect 21732 2372 21784 2378
rect 21732 2314 21784 2320
rect 21652 2145 21680 2314
rect 22296 2310 22324 3946
rect 22374 3224 22430 3233
rect 22374 3159 22430 3168
rect 22388 3058 22416 3159
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22388 2514 22416 2994
rect 22480 2514 22508 5306
rect 22572 4622 22600 6666
rect 22664 6186 22692 7346
rect 22848 6780 22876 7414
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22940 6914 22968 7346
rect 23296 7268 23348 7274
rect 23296 7210 23348 7216
rect 22940 6886 23060 6914
rect 22848 6752 22968 6780
rect 22742 6352 22798 6361
rect 22742 6287 22744 6296
rect 22796 6287 22798 6296
rect 22744 6258 22796 6264
rect 22652 6180 22704 6186
rect 22652 6122 22704 6128
rect 22940 5817 22968 6752
rect 23032 6497 23060 6886
rect 23018 6488 23074 6497
rect 23074 6446 23152 6474
rect 23018 6423 23074 6432
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 22926 5808 22982 5817
rect 22926 5743 22982 5752
rect 22940 5234 22968 5743
rect 23032 5370 23060 6258
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23124 5234 23152 6446
rect 23204 6112 23256 6118
rect 23204 6054 23256 6060
rect 23216 5846 23244 6054
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22664 4146 22692 4966
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22848 3194 22876 4082
rect 23032 3194 23060 5170
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23124 3534 23152 4558
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 22834 2680 22890 2689
rect 22834 2615 22890 2624
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22848 2446 22876 2615
rect 22928 2576 22980 2582
rect 22926 2544 22928 2553
rect 22980 2544 22982 2553
rect 22926 2479 22982 2488
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 22284 2304 22336 2310
rect 22284 2246 22336 2252
rect 21638 2136 21694 2145
rect 21638 2071 21694 2080
rect 23216 785 23244 4422
rect 23308 2650 23336 7210
rect 23400 3126 23428 9386
rect 23860 9178 23888 13270
rect 24214 13016 24270 13025
rect 24214 12951 24270 12960
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 24228 8498 24256 12951
rect 24504 9654 24532 13270
rect 24492 9648 24544 9654
rect 24492 9590 24544 9596
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24398 8256 24454 8265
rect 24398 8191 24454 8200
rect 24412 6934 24440 8191
rect 24400 6928 24452 6934
rect 24400 6870 24452 6876
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23202 776 23258 785
rect 23202 711 23258 720
rect 21916 672 21968 678
rect 21916 614 21968 620
rect 21928 100 21956 614
rect 19392 76 19394 100
rect 19338 0 19394 76
rect 19982 0 20038 100
rect 21914 0 21970 100
<< via2 >>
rect 1306 10920 1362 10976
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 386 10240 442 10296
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 386 9560 442 9616
rect 3330 8916 3332 8936
rect 3332 8916 3384 8936
rect 3384 8916 3386 8936
rect 3330 8880 3386 8916
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 386 7520 442 7576
rect 202 6840 258 6896
rect 3054 6296 3110 6352
rect 754 6160 810 6216
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 3790 6296 3846 6352
rect 754 5516 756 5536
rect 756 5516 808 5536
rect 808 5516 810 5536
rect 754 5480 810 5516
rect 4618 7828 4620 7848
rect 4620 7828 4672 7848
rect 4672 7828 4674 7848
rect 4618 7792 4674 7828
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 5262 7792 5318 7848
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3974 5208 4030 5264
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 570 4800 626 4856
rect 5998 8880 6054 8936
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 5354 5480 5410 5536
rect 5630 5908 5686 5944
rect 5630 5888 5632 5908
rect 5632 5888 5684 5908
rect 5684 5888 5686 5908
rect 6458 5344 6514 5400
rect 5906 5208 5962 5264
rect 5630 4800 5686 4856
rect 5170 4528 5226 4584
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 7010 5480 7066 5536
rect 7010 5228 7066 5264
rect 7010 5208 7012 5228
rect 7012 5208 7064 5228
rect 7064 5208 7066 5228
rect 7010 5072 7066 5128
rect 4618 3440 4674 3496
rect 754 2796 756 2816
rect 756 2796 808 2816
rect 808 2796 810 2816
rect 754 2760 810 2796
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 7286 5616 7342 5672
rect 7378 5228 7434 5264
rect 7378 5208 7380 5228
rect 7380 5208 7432 5228
rect 7432 5208 7434 5228
rect 7194 5072 7250 5128
rect 7194 4936 7250 4992
rect 7838 5344 7894 5400
rect 8482 6024 8538 6080
rect 8206 5228 8262 5264
rect 8206 5208 8208 5228
rect 8208 5208 8260 5228
rect 8260 5208 8262 5228
rect 7838 4664 7894 4720
rect 8022 3984 8078 4040
rect 9218 9152 9274 9208
rect 9770 9868 9772 9888
rect 9772 9868 9824 9888
rect 9824 9868 9826 9888
rect 9770 9832 9826 9868
rect 9034 7928 9090 7984
rect 8850 7384 8906 7440
rect 9586 7928 9642 7984
rect 9402 7404 9458 7440
rect 9402 7384 9404 7404
rect 9404 7384 9456 7404
rect 9456 7384 9458 7404
rect 10046 9016 10102 9072
rect 10690 9988 10746 10024
rect 10690 9968 10692 9988
rect 10692 9968 10744 9988
rect 10744 9968 10746 9988
rect 10138 7928 10194 7984
rect 10046 7656 10102 7712
rect 9494 6568 9550 6624
rect 8758 4936 8814 4992
rect 9218 4664 9274 4720
rect 7562 3032 7618 3088
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 8574 3032 8630 3088
rect 9310 4004 9366 4040
rect 9310 3984 9312 4004
rect 9312 3984 9364 4004
rect 9364 3984 9366 4004
rect 9218 3712 9274 3768
rect 9862 3712 9918 3768
rect 10138 5480 10194 5536
rect 10046 3576 10102 3632
rect 8758 2624 8814 2680
rect 10598 8880 10654 8936
rect 10782 8064 10838 8120
rect 10506 6432 10562 6488
rect 10966 7384 11022 7440
rect 10874 6432 10930 6488
rect 10874 5888 10930 5944
rect 10690 5752 10746 5808
rect 10782 2896 10838 2952
rect 10322 2760 10378 2816
rect 10138 2624 10194 2680
rect 8482 1808 8538 1864
rect 11058 6568 11114 6624
rect 12070 9424 12126 9480
rect 12070 8916 12072 8936
rect 12072 8916 12124 8936
rect 12124 8916 12126 8936
rect 11702 6976 11758 7032
rect 11334 6432 11390 6488
rect 11426 6296 11482 6352
rect 11242 5344 11298 5400
rect 11150 5208 11206 5264
rect 12070 8880 12126 8916
rect 12714 9696 12770 9752
rect 14186 9832 14242 9888
rect 14002 9444 14058 9480
rect 14002 9424 14004 9444
rect 14004 9424 14056 9444
rect 14056 9424 14058 9444
rect 13726 9288 13782 9344
rect 12898 8064 12954 8120
rect 12530 7112 12586 7168
rect 12162 5616 12218 5672
rect 11702 4120 11758 4176
rect 11058 2488 11114 2544
rect 12254 4664 12310 4720
rect 12254 4392 12310 4448
rect 12714 6840 12770 6896
rect 12622 6568 12678 6624
rect 12898 7284 12900 7304
rect 12900 7284 12952 7304
rect 12952 7284 12954 7304
rect 12898 7248 12954 7284
rect 12806 6432 12862 6488
rect 13174 6704 13230 6760
rect 13082 6432 13138 6488
rect 12438 4800 12494 4856
rect 14186 8472 14242 8528
rect 13358 6704 13414 6760
rect 13358 6604 13360 6624
rect 13360 6604 13412 6624
rect 13412 6604 13414 6624
rect 13358 6568 13414 6604
rect 13726 6160 13782 6216
rect 13726 5908 13782 5944
rect 13726 5888 13728 5908
rect 13728 5888 13780 5908
rect 13780 5888 13782 5908
rect 12990 5480 13046 5536
rect 12438 4664 12494 4720
rect 12438 4256 12494 4312
rect 12530 4120 12586 4176
rect 12162 3984 12218 4040
rect 11886 3848 11942 3904
rect 12346 3848 12402 3904
rect 12254 3052 12310 3088
rect 12254 3032 12256 3052
rect 12256 3032 12308 3052
rect 12308 3032 12310 3052
rect 12898 4256 12954 4312
rect 13174 4664 13230 4720
rect 13266 4564 13268 4584
rect 13268 4564 13320 4584
rect 13320 4564 13322 4584
rect 13266 4528 13322 4564
rect 13174 4392 13230 4448
rect 13358 4120 13414 4176
rect 13726 5480 13782 5536
rect 13542 4392 13598 4448
rect 13910 5888 13966 5944
rect 13910 5752 13966 5808
rect 14094 5344 14150 5400
rect 14002 4800 14058 4856
rect 15842 10648 15898 10704
rect 15014 9172 15070 9208
rect 15014 9152 15016 9172
rect 15016 9152 15068 9172
rect 15068 9152 15070 9172
rect 14462 7928 14518 7984
rect 14370 5616 14426 5672
rect 14278 5208 14334 5264
rect 14830 7656 14886 7712
rect 14646 6724 14702 6760
rect 14646 6704 14648 6724
rect 14648 6704 14700 6724
rect 14700 6704 14702 6724
rect 14922 7520 14978 7576
rect 15198 8336 15254 8392
rect 15198 8084 15254 8120
rect 15198 8064 15200 8084
rect 15200 8064 15252 8084
rect 15252 8064 15254 8084
rect 15750 9424 15806 9480
rect 15750 9152 15806 9208
rect 15566 8744 15622 8800
rect 16118 11056 16174 11112
rect 16118 9832 16174 9888
rect 15934 8744 15990 8800
rect 16670 10784 16726 10840
rect 16762 10376 16818 10432
rect 17682 12280 17738 12336
rect 17498 10920 17554 10976
rect 17406 10512 17462 10568
rect 16854 9424 16910 9480
rect 16394 8880 16450 8936
rect 16670 8880 16726 8936
rect 15014 7112 15070 7168
rect 14922 6296 14978 6352
rect 15290 6976 15346 7032
rect 14646 5072 14702 5128
rect 14094 4528 14150 4584
rect 13450 3848 13506 3904
rect 13174 3576 13230 3632
rect 12898 3304 12954 3360
rect 13266 3188 13322 3224
rect 13266 3168 13268 3188
rect 13268 3168 13320 3188
rect 13320 3168 13322 3188
rect 13450 2896 13506 2952
rect 14002 3440 14058 3496
rect 14278 3440 14334 3496
rect 14186 3032 14242 3088
rect 9678 40 9734 96
rect 14462 3884 14464 3904
rect 14464 3884 14516 3904
rect 14516 3884 14518 3904
rect 14462 3848 14518 3884
rect 15382 5208 15438 5264
rect 15290 5072 15346 5128
rect 15106 4936 15162 4992
rect 14738 4528 14794 4584
rect 15934 7656 15990 7712
rect 16026 7112 16082 7168
rect 15842 6976 15898 7032
rect 16578 8372 16580 8392
rect 16580 8372 16632 8392
rect 16632 8372 16634 8392
rect 16578 8336 16634 8372
rect 16578 8200 16634 8256
rect 16486 8064 16542 8120
rect 16394 6976 16450 7032
rect 16302 6840 16358 6896
rect 16578 6840 16634 6896
rect 16210 6704 16266 6760
rect 16118 6296 16174 6352
rect 15934 6024 15990 6080
rect 15658 5108 15660 5128
rect 15660 5108 15712 5128
rect 15712 5108 15714 5128
rect 15658 5072 15714 5108
rect 15566 4256 15622 4312
rect 15106 3304 15162 3360
rect 15474 3576 15530 3632
rect 15290 2488 15346 2544
rect 15934 5228 15990 5264
rect 16486 5616 16542 5672
rect 15934 5208 15936 5228
rect 15936 5208 15988 5228
rect 15988 5208 15990 5228
rect 15934 4256 15990 4312
rect 17038 9560 17094 9616
rect 18694 12008 18750 12064
rect 18050 11872 18106 11928
rect 18694 11600 18750 11656
rect 17682 9560 17738 9616
rect 17038 9288 17094 9344
rect 17222 9288 17278 9344
rect 17314 9152 17370 9208
rect 17958 10104 18014 10160
rect 18142 9696 18198 9752
rect 17682 9172 17738 9208
rect 17682 9152 17684 9172
rect 17684 9152 17736 9172
rect 17736 9152 17738 9172
rect 16854 8200 16910 8256
rect 17130 8200 17186 8256
rect 16762 7928 16818 7984
rect 16762 6840 16818 6896
rect 17222 7928 17278 7984
rect 18142 9460 18144 9480
rect 18144 9460 18196 9480
rect 18196 9460 18198 9480
rect 18142 9424 18198 9460
rect 17314 7656 17370 7712
rect 17590 7656 17646 7712
rect 17406 7112 17462 7168
rect 16578 5208 16634 5264
rect 16854 5208 16910 5264
rect 16854 5072 16910 5128
rect 16210 4020 16212 4040
rect 16212 4020 16264 4040
rect 16264 4020 16266 4040
rect 16210 3984 16266 4020
rect 16026 3712 16082 3768
rect 16394 4020 16396 4040
rect 16396 4020 16448 4040
rect 16448 4020 16450 4040
rect 16394 3984 16450 4020
rect 17038 5072 17094 5128
rect 17038 4972 17040 4992
rect 17040 4972 17092 4992
rect 17092 4972 17094 4992
rect 17038 4936 17094 4972
rect 17222 5636 17278 5672
rect 17222 5616 17224 5636
rect 17224 5616 17276 5636
rect 17276 5616 17278 5636
rect 17314 4664 17370 4720
rect 17406 4392 17462 4448
rect 16946 3712 17002 3768
rect 17958 7928 18014 7984
rect 17958 7656 18014 7712
rect 18234 8744 18290 8800
rect 18234 7928 18290 7984
rect 18050 6296 18106 6352
rect 17958 5652 17960 5672
rect 17960 5652 18012 5672
rect 18012 5652 18014 5672
rect 17958 5616 18014 5652
rect 17958 4528 18014 4584
rect 19154 9832 19210 9888
rect 18970 9016 19026 9072
rect 18878 8744 18934 8800
rect 18510 8472 18566 8528
rect 18510 7928 18566 7984
rect 18510 6296 18566 6352
rect 19062 7384 19118 7440
rect 18878 6296 18934 6352
rect 18602 6024 18658 6080
rect 18786 6060 18788 6080
rect 18788 6060 18840 6080
rect 18840 6060 18842 6080
rect 18786 6024 18842 6060
rect 18142 5344 18198 5400
rect 18050 3984 18106 4040
rect 18878 4936 18934 4992
rect 18234 3168 18290 3224
rect 19062 3848 19118 3904
rect 19798 10240 19854 10296
rect 19706 8492 19762 8528
rect 19706 8472 19708 8492
rect 19708 8472 19760 8492
rect 19760 8472 19762 8492
rect 19798 7792 19854 7848
rect 19614 7656 19670 7712
rect 21086 12008 21142 12064
rect 20810 11872 20866 11928
rect 21270 11056 21326 11112
rect 21178 10548 21180 10568
rect 21180 10548 21232 10568
rect 21232 10548 21234 10568
rect 21178 10512 21234 10548
rect 20350 9968 20406 10024
rect 20902 8608 20958 8664
rect 19890 6296 19946 6352
rect 20626 7792 20682 7848
rect 20902 6704 20958 6760
rect 20810 6568 20866 6624
rect 21270 8336 21326 8392
rect 21822 10376 21878 10432
rect 22466 10784 22522 10840
rect 22374 10668 22430 10704
rect 22374 10648 22376 10668
rect 22376 10648 22428 10668
rect 22428 10648 22430 10668
rect 21638 8064 21694 8120
rect 21914 8492 21970 8528
rect 21914 8472 21916 8492
rect 21916 8472 21968 8492
rect 21968 8472 21970 8492
rect 21914 6976 21970 7032
rect 21638 5228 21694 5264
rect 21638 5208 21640 5228
rect 21640 5208 21692 5228
rect 21692 5208 21694 5228
rect 22098 8916 22100 8936
rect 22100 8916 22152 8936
rect 22152 8916 22154 8936
rect 22098 8880 22154 8916
rect 22374 7248 22430 7304
rect 22834 9696 22890 9752
rect 22926 8336 22982 8392
rect 23110 9152 23166 9208
rect 22374 3168 22430 3224
rect 22742 6316 22798 6352
rect 22742 6296 22744 6316
rect 22744 6296 22796 6316
rect 22796 6296 22798 6316
rect 23018 6432 23074 6488
rect 22926 5752 22982 5808
rect 22834 2624 22890 2680
rect 22926 2524 22928 2544
rect 22928 2524 22980 2544
rect 22980 2524 22982 2544
rect 22926 2488 22982 2524
rect 21638 2080 21694 2136
rect 24214 12960 24270 13016
rect 24398 8200 24454 8256
rect 23202 720 23258 776
<< metal3 >>
rect 24209 13018 24275 13021
rect 24652 13018 24752 13048
rect 24209 13016 24752 13018
rect 24209 12960 24214 13016
rect 24270 12960 24752 13016
rect 24209 12958 24752 12960
rect 24209 12955 24275 12958
rect 24652 12928 24752 12958
rect 17677 12338 17743 12341
rect 24652 12338 24752 12368
rect 17677 12336 24752 12338
rect 17677 12280 17682 12336
rect 17738 12280 24752 12336
rect 17677 12278 24752 12280
rect 17677 12275 17743 12278
rect 24652 12248 24752 12278
rect 18689 12066 18755 12069
rect 21081 12066 21147 12069
rect 18689 12064 21147 12066
rect 18689 12008 18694 12064
rect 18750 12008 21086 12064
rect 21142 12008 21147 12064
rect 18689 12006 21147 12008
rect 18689 12003 18755 12006
rect 21081 12003 21147 12006
rect 18045 11930 18111 11933
rect 20805 11930 20871 11933
rect 18045 11928 20871 11930
rect 18045 11872 18050 11928
rect 18106 11872 20810 11928
rect 20866 11872 20871 11928
rect 18045 11870 20871 11872
rect 18045 11867 18111 11870
rect 20805 11867 20871 11870
rect 18689 11658 18755 11661
rect 24652 11658 24752 11688
rect 18689 11656 24752 11658
rect 18689 11600 18694 11656
rect 18750 11600 24752 11656
rect 18689 11598 24752 11600
rect 18689 11595 18755 11598
rect 24652 11568 24752 11598
rect 16113 11114 16179 11117
rect 21265 11114 21331 11117
rect 16113 11112 21331 11114
rect 16113 11056 16118 11112
rect 16174 11056 21270 11112
rect 21326 11056 21331 11112
rect 16113 11054 21331 11056
rect 16113 11051 16179 11054
rect 21265 11051 21331 11054
rect 0 10978 100 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 100 10918
rect 1301 10915 1367 10918
rect 17493 10978 17559 10981
rect 24652 10978 24752 11008
rect 17493 10976 24752 10978
rect 17493 10920 17498 10976
rect 17554 10920 24752 10976
rect 17493 10918 24752 10920
rect 17493 10915 17559 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 24652 10888 24752 10918
rect 4870 10847 5186 10848
rect 16665 10842 16731 10845
rect 22461 10842 22527 10845
rect 16665 10840 22527 10842
rect 16665 10784 16670 10840
rect 16726 10784 22466 10840
rect 22522 10784 22527 10840
rect 16665 10782 22527 10784
rect 16665 10779 16731 10782
rect 22461 10779 22527 10782
rect 15837 10706 15903 10709
rect 22369 10706 22435 10709
rect 15837 10704 22435 10706
rect 15837 10648 15842 10704
rect 15898 10648 22374 10704
rect 22430 10648 22435 10704
rect 15837 10646 22435 10648
rect 15837 10643 15903 10646
rect 22369 10643 22435 10646
rect 17401 10570 17467 10573
rect 21173 10570 21239 10573
rect 17401 10568 21239 10570
rect 17401 10512 17406 10568
rect 17462 10512 21178 10568
rect 21234 10512 21239 10568
rect 17401 10510 21239 10512
rect 17401 10507 17467 10510
rect 21173 10507 21239 10510
rect 16757 10434 16823 10437
rect 21817 10434 21883 10437
rect 16757 10432 21883 10434
rect 16757 10376 16762 10432
rect 16818 10376 21822 10432
rect 21878 10376 21883 10432
rect 16757 10374 21883 10376
rect 16757 10371 16823 10374
rect 21817 10371 21883 10374
rect 4210 10368 4526 10369
rect 0 10298 100 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 381 10298 447 10301
rect 0 10296 447 10298
rect 0 10240 386 10296
rect 442 10240 447 10296
rect 0 10238 447 10240
rect 0 10208 100 10238
rect 381 10235 447 10238
rect 19793 10298 19859 10301
rect 24652 10298 24752 10328
rect 19793 10296 24752 10298
rect 19793 10240 19798 10296
rect 19854 10240 24752 10296
rect 19793 10238 24752 10240
rect 19793 10235 19859 10238
rect 24652 10208 24752 10238
rect 17953 10162 18019 10165
rect 18822 10162 18828 10164
rect 17953 10160 18828 10162
rect 17953 10104 17958 10160
rect 18014 10104 18828 10160
rect 17953 10102 18828 10104
rect 17953 10099 18019 10102
rect 18822 10100 18828 10102
rect 18892 10100 18898 10164
rect 10685 10026 10751 10029
rect 20345 10026 20411 10029
rect 10685 10024 20411 10026
rect 10685 9968 10690 10024
rect 10746 9968 20350 10024
rect 20406 9968 20411 10024
rect 10685 9966 20411 9968
rect 10685 9963 10751 9966
rect 20345 9963 20411 9966
rect 9765 9890 9831 9893
rect 14181 9890 14247 9893
rect 9765 9888 14247 9890
rect 9765 9832 9770 9888
rect 9826 9832 14186 9888
rect 14242 9832 14247 9888
rect 9765 9830 14247 9832
rect 9765 9827 9831 9830
rect 14181 9827 14247 9830
rect 16113 9890 16179 9893
rect 19149 9890 19215 9893
rect 16113 9888 19215 9890
rect 16113 9832 16118 9888
rect 16174 9832 19154 9888
rect 19210 9832 19215 9888
rect 16113 9830 19215 9832
rect 16113 9827 16179 9830
rect 19149 9827 19215 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 12709 9754 12775 9757
rect 18137 9754 18203 9757
rect 18454 9754 18460 9756
rect 12709 9752 17970 9754
rect 12709 9696 12714 9752
rect 12770 9696 17970 9752
rect 12709 9694 17970 9696
rect 12709 9691 12775 9694
rect 0 9618 100 9648
rect 381 9618 447 9621
rect 0 9616 447 9618
rect 0 9560 386 9616
rect 442 9560 447 9616
rect 0 9558 447 9560
rect 0 9528 100 9558
rect 381 9555 447 9558
rect 9254 9556 9260 9620
rect 9324 9618 9330 9620
rect 17033 9618 17099 9621
rect 17677 9618 17743 9621
rect 9324 9616 17099 9618
rect 9324 9560 17038 9616
rect 17094 9560 17099 9616
rect 9324 9558 17099 9560
rect 9324 9556 9330 9558
rect 17033 9555 17099 9558
rect 17174 9616 17743 9618
rect 17174 9560 17682 9616
rect 17738 9560 17743 9616
rect 17174 9558 17743 9560
rect 17910 9618 17970 9694
rect 18137 9752 18460 9754
rect 18137 9696 18142 9752
rect 18198 9696 18460 9752
rect 18137 9694 18460 9696
rect 18137 9691 18203 9694
rect 18454 9692 18460 9694
rect 18524 9692 18530 9756
rect 21950 9692 21956 9756
rect 22020 9754 22026 9756
rect 22829 9754 22895 9757
rect 22020 9752 22895 9754
rect 22020 9696 22834 9752
rect 22890 9696 22895 9752
rect 22020 9694 22895 9696
rect 22020 9692 22026 9694
rect 22829 9691 22895 9694
rect 24652 9618 24752 9648
rect 17910 9558 24752 9618
rect 12065 9482 12131 9485
rect 13997 9482 14063 9485
rect 12065 9480 14063 9482
rect 12065 9424 12070 9480
rect 12126 9424 14002 9480
rect 14058 9424 14063 9480
rect 12065 9422 14063 9424
rect 12065 9419 12131 9422
rect 13997 9419 14063 9422
rect 15745 9482 15811 9485
rect 16849 9482 16915 9485
rect 17174 9482 17234 9558
rect 17677 9555 17743 9558
rect 24652 9528 24752 9558
rect 15745 9480 16915 9482
rect 15745 9424 15750 9480
rect 15806 9424 16854 9480
rect 16910 9424 16915 9480
rect 15745 9422 16915 9424
rect 15745 9419 15811 9422
rect 16849 9419 16915 9422
rect 17036 9422 17234 9482
rect 17036 9349 17096 9422
rect 17350 9420 17356 9484
rect 17420 9482 17426 9484
rect 18137 9482 18203 9485
rect 17420 9480 18203 9482
rect 17420 9424 18142 9480
rect 18198 9424 18203 9480
rect 17420 9422 18203 9424
rect 17420 9420 17426 9422
rect 18137 9419 18203 9422
rect 13721 9346 13787 9349
rect 16614 9346 16620 9348
rect 13721 9344 16620 9346
rect 13721 9288 13726 9344
rect 13782 9288 16620 9344
rect 13721 9286 16620 9288
rect 13721 9283 13787 9286
rect 16614 9284 16620 9286
rect 16684 9284 16690 9348
rect 17033 9344 17099 9349
rect 17033 9288 17038 9344
rect 17094 9288 17099 9344
rect 17033 9283 17099 9288
rect 17217 9346 17283 9349
rect 17217 9344 23490 9346
rect 17217 9288 17222 9344
rect 17278 9288 23490 9344
rect 17217 9286 23490 9288
rect 17217 9283 17283 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 9213 9210 9279 9213
rect 15009 9210 15075 9213
rect 15745 9210 15811 9213
rect 17309 9212 17375 9213
rect 17309 9210 17356 9212
rect 9213 9208 15811 9210
rect 9213 9152 9218 9208
rect 9274 9152 15014 9208
rect 15070 9152 15750 9208
rect 15806 9152 15811 9208
rect 9213 9150 15811 9152
rect 17264 9208 17356 9210
rect 17264 9152 17314 9208
rect 17264 9150 17356 9152
rect 9213 9147 9279 9150
rect 15009 9147 15075 9150
rect 15745 9147 15811 9150
rect 17309 9148 17356 9150
rect 17420 9148 17426 9212
rect 17677 9210 17743 9213
rect 23105 9210 23171 9213
rect 17677 9208 23171 9210
rect 17677 9152 17682 9208
rect 17738 9152 23110 9208
rect 23166 9152 23171 9208
rect 17677 9150 23171 9152
rect 17309 9147 17375 9148
rect 17677 9147 17743 9150
rect 23105 9147 23171 9150
rect 10041 9074 10107 9077
rect 18965 9074 19031 9077
rect 10041 9072 19031 9074
rect 10041 9016 10046 9072
rect 10102 9016 18970 9072
rect 19026 9016 19031 9072
rect 10041 9014 19031 9016
rect 10041 9011 10107 9014
rect 18965 9011 19031 9014
rect 3325 8938 3391 8941
rect 5993 8938 6059 8941
rect 3325 8936 6059 8938
rect 3325 8880 3330 8936
rect 3386 8880 5998 8936
rect 6054 8880 6059 8936
rect 3325 8878 6059 8880
rect 3325 8875 3391 8878
rect 5993 8875 6059 8878
rect 10593 8938 10659 8941
rect 12065 8938 12131 8941
rect 16389 8938 16455 8941
rect 16665 8940 16731 8941
rect 16614 8938 16620 8940
rect 10593 8936 16455 8938
rect 10593 8880 10598 8936
rect 10654 8880 12070 8936
rect 12126 8880 16394 8936
rect 16450 8880 16455 8936
rect 10593 8878 16455 8880
rect 16574 8878 16620 8938
rect 16684 8936 16731 8940
rect 16726 8880 16731 8936
rect 10593 8875 10659 8878
rect 12065 8875 12131 8878
rect 16389 8875 16455 8878
rect 16614 8876 16620 8878
rect 16684 8876 16731 8880
rect 16982 8876 16988 8940
rect 17052 8938 17058 8940
rect 22093 8938 22159 8941
rect 17052 8936 22159 8938
rect 17052 8880 22098 8936
rect 22154 8880 22159 8936
rect 17052 8878 22159 8880
rect 23430 8938 23490 9286
rect 24652 8938 24752 8968
rect 23430 8878 24752 8938
rect 17052 8876 17058 8878
rect 16665 8875 16731 8876
rect 22093 8875 22159 8878
rect 24652 8848 24752 8878
rect 15561 8802 15627 8805
rect 15929 8802 15995 8805
rect 18229 8802 18295 8805
rect 18873 8802 18939 8805
rect 15561 8800 18939 8802
rect 15561 8744 15566 8800
rect 15622 8744 15934 8800
rect 15990 8744 18234 8800
rect 18290 8744 18878 8800
rect 18934 8744 18939 8800
rect 15561 8742 18939 8744
rect 15561 8739 15627 8742
rect 15929 8739 15995 8742
rect 18229 8739 18295 8742
rect 18873 8739 18939 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 14222 8604 14228 8668
rect 14292 8666 14298 8668
rect 20897 8666 20963 8669
rect 14292 8664 20963 8666
rect 14292 8608 20902 8664
rect 20958 8608 20963 8664
rect 14292 8606 20963 8608
rect 14292 8604 14298 8606
rect 20897 8603 20963 8606
rect 14181 8530 14247 8533
rect 18505 8530 18571 8533
rect 14181 8528 18571 8530
rect 14181 8472 14186 8528
rect 14242 8472 18510 8528
rect 18566 8472 18571 8528
rect 14181 8470 18571 8472
rect 14181 8467 14247 8470
rect 18505 8467 18571 8470
rect 19701 8530 19767 8533
rect 21909 8530 21975 8533
rect 19701 8528 21975 8530
rect 19701 8472 19706 8528
rect 19762 8472 21914 8528
rect 21970 8472 21975 8528
rect 19701 8470 21975 8472
rect 19701 8467 19767 8470
rect 21909 8467 21975 8470
rect 14774 8332 14780 8396
rect 14844 8394 14850 8396
rect 15193 8394 15259 8397
rect 14844 8392 15259 8394
rect 14844 8336 15198 8392
rect 15254 8336 15259 8392
rect 14844 8334 15259 8336
rect 14844 8332 14850 8334
rect 15193 8331 15259 8334
rect 16573 8394 16639 8397
rect 21265 8394 21331 8397
rect 22921 8394 22987 8397
rect 16573 8392 21331 8394
rect 16573 8336 16578 8392
rect 16634 8336 21270 8392
rect 21326 8336 21331 8392
rect 16573 8334 21331 8336
rect 16573 8331 16639 8334
rect 21265 8331 21331 8334
rect 22050 8392 22987 8394
rect 22050 8336 22926 8392
rect 22982 8336 22987 8392
rect 22050 8334 22987 8336
rect 13670 8196 13676 8260
rect 13740 8258 13746 8260
rect 16573 8258 16639 8261
rect 13740 8256 16639 8258
rect 13740 8200 16578 8256
rect 16634 8200 16639 8256
rect 13740 8198 16639 8200
rect 13740 8196 13746 8198
rect 16573 8195 16639 8198
rect 16849 8258 16915 8261
rect 16982 8258 16988 8260
rect 16849 8256 16988 8258
rect 16849 8200 16854 8256
rect 16910 8200 16988 8256
rect 16849 8198 16988 8200
rect 16849 8195 16915 8198
rect 16982 8196 16988 8198
rect 17052 8196 17058 8260
rect 17125 8258 17191 8261
rect 22050 8258 22110 8334
rect 22921 8331 22987 8334
rect 17125 8256 22110 8258
rect 17125 8200 17130 8256
rect 17186 8200 22110 8256
rect 17125 8198 22110 8200
rect 24393 8258 24459 8261
rect 24652 8258 24752 8288
rect 24393 8256 24752 8258
rect 24393 8200 24398 8256
rect 24454 8200 24752 8256
rect 24393 8198 24752 8200
rect 17125 8195 17191 8198
rect 24393 8195 24459 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 24652 8168 24752 8198
rect 4210 8127 4526 8128
rect 10777 8122 10843 8125
rect 12893 8122 12959 8125
rect 15193 8122 15259 8125
rect 16481 8122 16547 8125
rect 21633 8122 21699 8125
rect 10777 8120 15026 8122
rect 10777 8064 10782 8120
rect 10838 8064 12898 8120
rect 12954 8064 15026 8120
rect 10777 8062 15026 8064
rect 10777 8059 10843 8062
rect 12893 8059 12959 8062
rect 9029 7986 9095 7989
rect 9581 7986 9647 7989
rect 9029 7984 9647 7986
rect 9029 7928 9034 7984
rect 9090 7928 9586 7984
rect 9642 7928 9647 7984
rect 9029 7926 9647 7928
rect 9029 7923 9095 7926
rect 9581 7923 9647 7926
rect 10133 7986 10199 7989
rect 14457 7986 14523 7989
rect 14966 7988 15026 8062
rect 15193 8120 21699 8122
rect 15193 8064 15198 8120
rect 15254 8064 16486 8120
rect 16542 8064 21638 8120
rect 21694 8064 21699 8120
rect 15193 8062 21699 8064
rect 15193 8059 15259 8062
rect 16481 8059 16547 8062
rect 21633 8059 21699 8062
rect 10133 7984 14523 7986
rect 10133 7928 10138 7984
rect 10194 7928 14462 7984
rect 14518 7928 14523 7984
rect 10133 7926 14523 7928
rect 10133 7923 10199 7926
rect 14457 7923 14523 7926
rect 14958 7924 14964 7988
rect 15028 7986 15034 7988
rect 16757 7986 16823 7989
rect 15028 7984 16823 7986
rect 15028 7928 16762 7984
rect 16818 7928 16823 7984
rect 15028 7926 16823 7928
rect 15028 7924 15034 7926
rect 16757 7923 16823 7926
rect 17217 7986 17283 7989
rect 17953 7986 18019 7989
rect 18229 7986 18295 7989
rect 17217 7984 18295 7986
rect 17217 7928 17222 7984
rect 17278 7928 17958 7984
rect 18014 7928 18234 7984
rect 18290 7928 18295 7984
rect 17217 7926 18295 7928
rect 17217 7923 17283 7926
rect 17953 7923 18019 7926
rect 18229 7923 18295 7926
rect 18505 7986 18571 7989
rect 18638 7986 18644 7988
rect 18505 7984 18644 7986
rect 18505 7928 18510 7984
rect 18566 7928 18644 7984
rect 18505 7926 18644 7928
rect 18505 7923 18571 7926
rect 18638 7924 18644 7926
rect 18708 7924 18714 7988
rect 4613 7850 4679 7853
rect 5257 7850 5323 7853
rect 19793 7850 19859 7853
rect 20621 7850 20687 7853
rect 4613 7848 20687 7850
rect 4613 7792 4618 7848
rect 4674 7792 5262 7848
rect 5318 7792 19798 7848
rect 19854 7792 20626 7848
rect 20682 7792 20687 7848
rect 4613 7790 20687 7792
rect 4613 7787 4679 7790
rect 5257 7787 5323 7790
rect 19793 7787 19859 7790
rect 20621 7787 20687 7790
rect 10041 7714 10107 7717
rect 14825 7714 14891 7717
rect 15929 7716 15995 7717
rect 10041 7712 14891 7714
rect 10041 7656 10046 7712
rect 10102 7656 14830 7712
rect 14886 7656 14891 7712
rect 10041 7654 14891 7656
rect 10041 7651 10107 7654
rect 14825 7651 14891 7654
rect 15878 7652 15884 7716
rect 15948 7714 15995 7716
rect 17309 7714 17375 7717
rect 17585 7714 17651 7717
rect 15948 7712 16040 7714
rect 15990 7656 16040 7712
rect 15948 7654 16040 7656
rect 17309 7712 17651 7714
rect 17309 7656 17314 7712
rect 17370 7656 17590 7712
rect 17646 7656 17651 7712
rect 17309 7654 17651 7656
rect 15948 7652 15995 7654
rect 15929 7651 15995 7652
rect 17309 7651 17375 7654
rect 17585 7651 17651 7654
rect 17953 7714 18019 7717
rect 19609 7714 19675 7717
rect 17953 7712 19675 7714
rect 17953 7656 17958 7712
rect 18014 7656 19614 7712
rect 19670 7656 19675 7712
rect 17953 7654 19675 7656
rect 17953 7651 18019 7654
rect 19609 7651 19675 7654
rect 4870 7648 5186 7649
rect 0 7578 100 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 381 7578 447 7581
rect 0 7576 447 7578
rect 0 7520 386 7576
rect 442 7520 447 7576
rect 0 7518 447 7520
rect 0 7488 100 7518
rect 381 7515 447 7518
rect 14917 7578 14983 7581
rect 24652 7578 24752 7608
rect 14917 7576 24752 7578
rect 14917 7520 14922 7576
rect 14978 7520 24752 7576
rect 14917 7518 24752 7520
rect 14917 7515 14983 7518
rect 24652 7488 24752 7518
rect 8845 7442 8911 7445
rect 9397 7442 9463 7445
rect 8845 7440 9463 7442
rect 8845 7384 8850 7440
rect 8906 7384 9402 7440
rect 9458 7384 9463 7440
rect 8845 7382 9463 7384
rect 8845 7379 8911 7382
rect 9397 7379 9463 7382
rect 10961 7442 11027 7445
rect 19057 7442 19123 7445
rect 10961 7440 19123 7442
rect 10961 7384 10966 7440
rect 11022 7384 19062 7440
rect 19118 7384 19123 7440
rect 10961 7382 19123 7384
rect 10961 7379 11027 7382
rect 19057 7379 19123 7382
rect 12893 7306 12959 7309
rect 22369 7306 22435 7309
rect 12893 7304 22435 7306
rect 12893 7248 12898 7304
rect 12954 7248 22374 7304
rect 22430 7248 22435 7304
rect 12893 7246 22435 7248
rect 12893 7243 12959 7246
rect 22369 7243 22435 7246
rect 12525 7170 12591 7173
rect 15009 7170 15075 7173
rect 12525 7168 15075 7170
rect 12525 7112 12530 7168
rect 12586 7112 15014 7168
rect 15070 7112 15075 7168
rect 12525 7110 15075 7112
rect 12525 7107 12591 7110
rect 15009 7107 15075 7110
rect 16021 7170 16087 7173
rect 17401 7170 17467 7173
rect 16021 7168 17467 7170
rect 16021 7112 16026 7168
rect 16082 7112 17406 7168
rect 17462 7112 17467 7168
rect 16021 7110 17467 7112
rect 16021 7107 16087 7110
rect 17401 7107 17467 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 11697 7034 11763 7037
rect 15285 7034 15351 7037
rect 11697 7032 15351 7034
rect 11697 6976 11702 7032
rect 11758 6976 15290 7032
rect 15346 6976 15351 7032
rect 11697 6974 15351 6976
rect 11697 6971 11763 6974
rect 15285 6971 15351 6974
rect 15510 6972 15516 7036
rect 15580 7034 15586 7036
rect 15837 7034 15903 7037
rect 15580 7032 15903 7034
rect 15580 6976 15842 7032
rect 15898 6976 15903 7032
rect 15580 6974 15903 6976
rect 15580 6972 15586 6974
rect 15837 6971 15903 6974
rect 16389 7034 16455 7037
rect 21909 7034 21975 7037
rect 16389 7032 21975 7034
rect 16389 6976 16394 7032
rect 16450 6976 21914 7032
rect 21970 6976 21975 7032
rect 16389 6974 21975 6976
rect 16389 6971 16455 6974
rect 21909 6971 21975 6974
rect 0 6898 100 6928
rect 197 6898 263 6901
rect 0 6896 263 6898
rect 0 6840 202 6896
rect 258 6840 263 6896
rect 0 6838 263 6840
rect 0 6808 100 6838
rect 197 6835 263 6838
rect 12709 6898 12775 6901
rect 16297 6898 16363 6901
rect 16573 6900 16639 6901
rect 16573 6898 16620 6900
rect 12709 6896 16363 6898
rect 12709 6840 12714 6896
rect 12770 6840 16302 6896
rect 16358 6840 16363 6896
rect 12709 6838 16363 6840
rect 16528 6896 16620 6898
rect 16528 6840 16578 6896
rect 16528 6838 16620 6840
rect 12709 6835 12775 6838
rect 16297 6835 16363 6838
rect 16573 6836 16620 6838
rect 16684 6836 16690 6900
rect 16757 6898 16823 6901
rect 24652 6898 24752 6928
rect 16757 6896 24752 6898
rect 16757 6840 16762 6896
rect 16818 6840 24752 6896
rect 16757 6838 24752 6840
rect 16573 6835 16639 6836
rect 16757 6835 16823 6838
rect 24652 6808 24752 6838
rect 13169 6762 13235 6765
rect 13353 6762 13419 6765
rect 13169 6760 13419 6762
rect 13169 6704 13174 6760
rect 13230 6704 13358 6760
rect 13414 6704 13419 6760
rect 13169 6702 13419 6704
rect 13169 6699 13235 6702
rect 13353 6699 13419 6702
rect 14038 6700 14044 6764
rect 14108 6762 14114 6764
rect 14641 6762 14707 6765
rect 14108 6760 14707 6762
rect 14108 6704 14646 6760
rect 14702 6704 14707 6760
rect 14108 6702 14707 6704
rect 14108 6700 14114 6702
rect 14641 6699 14707 6702
rect 16205 6762 16271 6765
rect 20897 6762 20963 6765
rect 16205 6760 20963 6762
rect 16205 6704 16210 6760
rect 16266 6704 20902 6760
rect 20958 6704 20963 6760
rect 16205 6702 20963 6704
rect 16205 6699 16271 6702
rect 20897 6699 20963 6702
rect 9489 6626 9555 6629
rect 11053 6626 11119 6629
rect 9489 6624 11119 6626
rect 9489 6568 9494 6624
rect 9550 6568 11058 6624
rect 11114 6568 11119 6624
rect 9489 6566 11119 6568
rect 9489 6563 9555 6566
rect 11053 6563 11119 6566
rect 12617 6626 12683 6629
rect 13353 6626 13419 6629
rect 20805 6626 20871 6629
rect 12617 6624 20871 6626
rect 12617 6568 12622 6624
rect 12678 6568 13358 6624
rect 13414 6568 20810 6624
rect 20866 6568 20871 6624
rect 12617 6566 20871 6568
rect 12617 6563 12683 6566
rect 13353 6563 13419 6566
rect 20805 6563 20871 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 10501 6490 10567 6493
rect 10869 6490 10935 6493
rect 10501 6488 10935 6490
rect 10501 6432 10506 6488
rect 10562 6432 10874 6488
rect 10930 6432 10935 6488
rect 10501 6430 10935 6432
rect 10501 6427 10567 6430
rect 10869 6427 10935 6430
rect 11329 6490 11395 6493
rect 12801 6490 12867 6493
rect 11329 6488 12867 6490
rect 11329 6432 11334 6488
rect 11390 6432 12806 6488
rect 12862 6432 12867 6488
rect 11329 6430 12867 6432
rect 11329 6427 11395 6430
rect 12801 6427 12867 6430
rect 13077 6490 13143 6493
rect 23013 6490 23079 6493
rect 13077 6488 23079 6490
rect 13077 6432 13082 6488
rect 13138 6432 23018 6488
rect 23074 6432 23079 6488
rect 13077 6430 23079 6432
rect 13077 6427 13143 6430
rect 23013 6427 23079 6430
rect 3049 6354 3115 6357
rect 3785 6354 3851 6357
rect 11421 6354 11487 6357
rect 14917 6356 14983 6357
rect 14917 6354 14964 6356
rect 3049 6352 11487 6354
rect 3049 6296 3054 6352
rect 3110 6296 3790 6352
rect 3846 6296 11426 6352
rect 11482 6296 11487 6352
rect 3049 6294 11487 6296
rect 14872 6352 14964 6354
rect 14872 6296 14922 6352
rect 14872 6294 14964 6296
rect 3049 6291 3115 6294
rect 3785 6291 3851 6294
rect 11421 6291 11487 6294
rect 14917 6292 14964 6294
rect 15028 6292 15034 6356
rect 15694 6292 15700 6356
rect 15764 6354 15770 6356
rect 16113 6354 16179 6357
rect 15764 6352 16179 6354
rect 15764 6296 16118 6352
rect 16174 6296 16179 6352
rect 15764 6294 16179 6296
rect 15764 6292 15770 6294
rect 14917 6291 14983 6292
rect 16113 6291 16179 6294
rect 18045 6354 18111 6357
rect 18505 6354 18571 6357
rect 18873 6354 18939 6357
rect 18045 6352 18939 6354
rect 18045 6296 18050 6352
rect 18106 6296 18510 6352
rect 18566 6296 18878 6352
rect 18934 6296 18939 6352
rect 18045 6294 18939 6296
rect 18045 6291 18111 6294
rect 18505 6291 18571 6294
rect 18873 6291 18939 6294
rect 19885 6354 19951 6357
rect 22737 6354 22803 6357
rect 19885 6352 22803 6354
rect 19885 6296 19890 6352
rect 19946 6296 22742 6352
rect 22798 6296 22803 6352
rect 19885 6294 22803 6296
rect 19885 6291 19951 6294
rect 22737 6291 22803 6294
rect 0 6218 100 6248
rect 749 6218 815 6221
rect 0 6216 815 6218
rect 0 6160 754 6216
rect 810 6160 815 6216
rect 0 6158 815 6160
rect 0 6128 100 6158
rect 749 6155 815 6158
rect 13721 6218 13787 6221
rect 24652 6218 24752 6248
rect 13721 6216 24752 6218
rect 13721 6160 13726 6216
rect 13782 6160 24752 6216
rect 13721 6158 24752 6160
rect 13721 6155 13787 6158
rect 24652 6128 24752 6158
rect 8477 6082 8543 6085
rect 15929 6082 15995 6085
rect 8477 6080 15995 6082
rect 8477 6024 8482 6080
rect 8538 6024 15934 6080
rect 15990 6024 15995 6080
rect 8477 6022 15995 6024
rect 8477 6019 8543 6022
rect 15929 6019 15995 6022
rect 16614 6020 16620 6084
rect 16684 6082 16690 6084
rect 18597 6082 18663 6085
rect 16684 6080 18663 6082
rect 16684 6024 18602 6080
rect 18658 6024 18663 6080
rect 16684 6022 18663 6024
rect 16684 6020 16690 6022
rect 18597 6019 18663 6022
rect 18781 6084 18847 6085
rect 18781 6080 18828 6084
rect 18892 6082 18898 6084
rect 18781 6024 18786 6080
rect 18781 6020 18828 6024
rect 18892 6022 18938 6082
rect 18892 6020 18898 6022
rect 18781 6019 18847 6020
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 5625 5946 5691 5949
rect 10869 5946 10935 5949
rect 13721 5948 13787 5949
rect 13670 5946 13676 5948
rect 5625 5944 10935 5946
rect 5625 5888 5630 5944
rect 5686 5888 10874 5944
rect 10930 5888 10935 5944
rect 5625 5886 10935 5888
rect 13630 5886 13676 5946
rect 13740 5944 13787 5948
rect 13782 5888 13787 5944
rect 5625 5883 5691 5886
rect 10869 5883 10935 5886
rect 13670 5884 13676 5886
rect 13740 5884 13787 5888
rect 13721 5883 13787 5884
rect 13905 5946 13971 5949
rect 17902 5946 17908 5948
rect 13905 5944 17908 5946
rect 13905 5888 13910 5944
rect 13966 5888 17908 5944
rect 13905 5886 17908 5888
rect 13905 5883 13971 5886
rect 17902 5884 17908 5886
rect 17972 5884 17978 5948
rect 10685 5810 10751 5813
rect 13905 5810 13971 5813
rect 22921 5810 22987 5813
rect 10685 5808 22987 5810
rect 10685 5752 10690 5808
rect 10746 5752 13910 5808
rect 13966 5752 22926 5808
rect 22982 5752 22987 5808
rect 10685 5750 22987 5752
rect 10685 5747 10751 5750
rect 13905 5747 13971 5750
rect 22921 5747 22987 5750
rect 7281 5674 7347 5677
rect 12157 5674 12223 5677
rect 14038 5674 14044 5676
rect 7281 5672 14044 5674
rect 7281 5616 7286 5672
rect 7342 5616 12162 5672
rect 12218 5616 14044 5672
rect 7281 5614 14044 5616
rect 7281 5611 7347 5614
rect 12157 5611 12223 5614
rect 14038 5612 14044 5614
rect 14108 5612 14114 5676
rect 14365 5674 14431 5677
rect 15142 5674 15148 5676
rect 14365 5672 15148 5674
rect 14365 5616 14370 5672
rect 14426 5616 15148 5672
rect 14365 5614 15148 5616
rect 14365 5611 14431 5614
rect 15142 5612 15148 5614
rect 15212 5612 15218 5676
rect 16481 5674 16547 5677
rect 17217 5674 17283 5677
rect 16481 5672 17283 5674
rect 16481 5616 16486 5672
rect 16542 5616 17222 5672
rect 17278 5616 17283 5672
rect 16481 5614 17283 5616
rect 16481 5611 16547 5614
rect 17217 5611 17283 5614
rect 17953 5674 18019 5677
rect 18454 5674 18460 5676
rect 17953 5672 18460 5674
rect 17953 5616 17958 5672
rect 18014 5616 18460 5672
rect 17953 5614 18460 5616
rect 17953 5611 18019 5614
rect 18454 5612 18460 5614
rect 18524 5612 18530 5676
rect 0 5538 100 5568
rect 749 5538 815 5541
rect 0 5536 815 5538
rect 0 5480 754 5536
rect 810 5480 815 5536
rect 0 5478 815 5480
rect 0 5448 100 5478
rect 749 5475 815 5478
rect 5349 5538 5415 5541
rect 7005 5538 7071 5541
rect 5349 5536 7071 5538
rect 5349 5480 5354 5536
rect 5410 5480 7010 5536
rect 7066 5480 7071 5536
rect 5349 5478 7071 5480
rect 5349 5475 5415 5478
rect 7005 5475 7071 5478
rect 10133 5538 10199 5541
rect 12985 5538 13051 5541
rect 10133 5536 13051 5538
rect 10133 5480 10138 5536
rect 10194 5480 12990 5536
rect 13046 5480 13051 5536
rect 10133 5478 13051 5480
rect 10133 5475 10199 5478
rect 12985 5475 13051 5478
rect 13721 5538 13787 5541
rect 24652 5538 24752 5568
rect 13721 5536 24752 5538
rect 13721 5480 13726 5536
rect 13782 5480 24752 5536
rect 13721 5478 24752 5480
rect 13721 5475 13787 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 24652 5448 24752 5478
rect 4870 5407 5186 5408
rect 6453 5402 6519 5405
rect 7833 5402 7899 5405
rect 6453 5400 7899 5402
rect 6453 5344 6458 5400
rect 6514 5344 7838 5400
rect 7894 5344 7899 5400
rect 6453 5342 7899 5344
rect 6453 5339 6519 5342
rect 7833 5339 7899 5342
rect 11237 5402 11303 5405
rect 14089 5402 14155 5405
rect 18137 5402 18203 5405
rect 11237 5400 18203 5402
rect 11237 5344 11242 5400
rect 11298 5344 14094 5400
rect 14150 5344 18142 5400
rect 18198 5344 18203 5400
rect 11237 5342 18203 5344
rect 11237 5339 11303 5342
rect 14089 5339 14155 5342
rect 18137 5339 18203 5342
rect 3969 5266 4035 5269
rect 5901 5266 5967 5269
rect 7005 5266 7071 5269
rect 3969 5264 7071 5266
rect 3969 5208 3974 5264
rect 4030 5208 5906 5264
rect 5962 5208 7010 5264
rect 7066 5208 7071 5264
rect 3969 5206 7071 5208
rect 3969 5203 4035 5206
rect 5901 5203 5967 5206
rect 7005 5203 7071 5206
rect 7373 5266 7439 5269
rect 8201 5266 8267 5269
rect 7373 5264 8267 5266
rect 7373 5208 7378 5264
rect 7434 5208 8206 5264
rect 8262 5208 8267 5264
rect 7373 5206 8267 5208
rect 7373 5203 7439 5206
rect 8201 5203 8267 5206
rect 11145 5266 11211 5269
rect 14273 5266 14339 5269
rect 15377 5266 15443 5269
rect 11145 5264 15443 5266
rect 11145 5208 11150 5264
rect 11206 5208 14278 5264
rect 14334 5208 15382 5264
rect 15438 5208 15443 5264
rect 11145 5206 15443 5208
rect 11145 5203 11211 5206
rect 14273 5203 14339 5206
rect 15377 5203 15443 5206
rect 15929 5266 15995 5269
rect 16573 5266 16639 5269
rect 16849 5266 16915 5269
rect 15929 5264 16915 5266
rect 15929 5208 15934 5264
rect 15990 5208 16578 5264
rect 16634 5208 16854 5264
rect 16910 5208 16915 5264
rect 15929 5206 16915 5208
rect 15929 5203 15995 5206
rect 16573 5203 16639 5206
rect 16849 5203 16915 5206
rect 17902 5204 17908 5268
rect 17972 5266 17978 5268
rect 21633 5266 21699 5269
rect 17972 5264 21699 5266
rect 17972 5208 21638 5264
rect 21694 5208 21699 5264
rect 17972 5206 21699 5208
rect 17972 5204 17978 5206
rect 21633 5203 21699 5206
rect 7005 5130 7071 5133
rect 7189 5130 7255 5133
rect 7005 5128 7255 5130
rect 7005 5072 7010 5128
rect 7066 5072 7194 5128
rect 7250 5072 7255 5128
rect 7005 5070 7255 5072
rect 7005 5067 7071 5070
rect 7189 5067 7255 5070
rect 14641 5130 14707 5133
rect 14774 5130 14780 5132
rect 14641 5128 14780 5130
rect 14641 5072 14646 5128
rect 14702 5072 14780 5128
rect 14641 5070 14780 5072
rect 14641 5067 14707 5070
rect 14774 5068 14780 5070
rect 14844 5130 14850 5132
rect 15285 5130 15351 5133
rect 14844 5128 15351 5130
rect 14844 5072 15290 5128
rect 15346 5072 15351 5128
rect 14844 5070 15351 5072
rect 14844 5068 14850 5070
rect 15285 5067 15351 5070
rect 15653 5130 15719 5133
rect 16849 5130 16915 5133
rect 17033 5130 17099 5133
rect 15653 5128 17099 5130
rect 15653 5072 15658 5128
rect 15714 5072 16854 5128
rect 16910 5072 17038 5128
rect 17094 5072 17099 5128
rect 15653 5070 17099 5072
rect 15653 5067 15719 5070
rect 16849 5067 16915 5070
rect 17033 5067 17099 5070
rect 7189 4994 7255 4997
rect 8753 4994 8819 4997
rect 7189 4992 8819 4994
rect 7189 4936 7194 4992
rect 7250 4936 8758 4992
rect 8814 4936 8819 4992
rect 7189 4934 8819 4936
rect 7189 4931 7255 4934
rect 8753 4931 8819 4934
rect 15101 4994 15167 4997
rect 17033 4994 17099 4997
rect 18873 4994 18939 4997
rect 15101 4992 18939 4994
rect 15101 4936 15106 4992
rect 15162 4936 17038 4992
rect 17094 4936 18878 4992
rect 18934 4936 18939 4992
rect 15101 4934 18939 4936
rect 15101 4931 15167 4934
rect 17033 4931 17099 4934
rect 18873 4931 18939 4934
rect 4210 4928 4526 4929
rect 0 4858 100 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 565 4858 631 4861
rect 0 4856 631 4858
rect 0 4800 570 4856
rect 626 4800 631 4856
rect 0 4798 631 4800
rect 0 4768 100 4798
rect 565 4795 631 4798
rect 5625 4858 5691 4861
rect 12433 4858 12499 4861
rect 5625 4856 12499 4858
rect 5625 4800 5630 4856
rect 5686 4800 12438 4856
rect 12494 4800 12499 4856
rect 5625 4798 12499 4800
rect 5625 4795 5691 4798
rect 12433 4795 12499 4798
rect 13997 4858 14063 4861
rect 24652 4858 24752 4888
rect 13997 4856 24752 4858
rect 13997 4800 14002 4856
rect 14058 4800 24752 4856
rect 13997 4798 24752 4800
rect 13997 4795 14063 4798
rect 24652 4768 24752 4798
rect 7833 4722 7899 4725
rect 9213 4724 9279 4725
rect 9213 4722 9260 4724
rect 7833 4720 9260 4722
rect 7833 4664 7838 4720
rect 7894 4664 9218 4720
rect 7833 4662 9260 4664
rect 7833 4659 7899 4662
rect 9213 4660 9260 4662
rect 9324 4660 9330 4724
rect 12249 4722 12315 4725
rect 12433 4722 12499 4725
rect 12249 4720 12499 4722
rect 12249 4664 12254 4720
rect 12310 4664 12438 4720
rect 12494 4664 12499 4720
rect 12249 4662 12499 4664
rect 9213 4659 9279 4660
rect 12249 4659 12315 4662
rect 12433 4659 12499 4662
rect 13169 4722 13235 4725
rect 17309 4722 17375 4725
rect 13169 4720 17375 4722
rect 13169 4664 13174 4720
rect 13230 4664 17314 4720
rect 17370 4664 17375 4720
rect 13169 4662 17375 4664
rect 13169 4659 13235 4662
rect 17309 4659 17375 4662
rect 5165 4586 5231 4589
rect 13261 4586 13327 4589
rect 5165 4584 13327 4586
rect 5165 4528 5170 4584
rect 5226 4528 13266 4584
rect 13322 4528 13327 4584
rect 5165 4526 13327 4528
rect 5165 4523 5231 4526
rect 13261 4523 13327 4526
rect 14089 4586 14155 4589
rect 14222 4586 14228 4588
rect 14089 4584 14228 4586
rect 14089 4528 14094 4584
rect 14150 4528 14228 4584
rect 14089 4526 14228 4528
rect 14089 4523 14155 4526
rect 14222 4524 14228 4526
rect 14292 4524 14298 4588
rect 14733 4586 14799 4589
rect 17953 4586 18019 4589
rect 14733 4584 18019 4586
rect 14733 4528 14738 4584
rect 14794 4528 17958 4584
rect 18014 4528 18019 4584
rect 14733 4526 18019 4528
rect 14733 4523 14799 4526
rect 17953 4523 18019 4526
rect 12249 4450 12315 4453
rect 13169 4450 13235 4453
rect 12249 4448 13235 4450
rect 12249 4392 12254 4448
rect 12310 4392 13174 4448
rect 13230 4392 13235 4448
rect 12249 4390 13235 4392
rect 12249 4387 12315 4390
rect 13169 4387 13235 4390
rect 13537 4450 13603 4453
rect 17401 4450 17467 4453
rect 13537 4448 17467 4450
rect 13537 4392 13542 4448
rect 13598 4392 17406 4448
rect 17462 4392 17467 4448
rect 13537 4390 17467 4392
rect 13537 4387 13603 4390
rect 17401 4387 17467 4390
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 12433 4314 12499 4317
rect 12893 4314 12959 4317
rect 12433 4312 12959 4314
rect 12433 4256 12438 4312
rect 12494 4256 12898 4312
rect 12954 4256 12959 4312
rect 12433 4254 12959 4256
rect 12433 4251 12499 4254
rect 12893 4251 12959 4254
rect 15561 4314 15627 4317
rect 15929 4316 15995 4317
rect 15694 4314 15700 4316
rect 15561 4312 15700 4314
rect 15561 4256 15566 4312
rect 15622 4256 15700 4312
rect 15561 4254 15700 4256
rect 15561 4251 15627 4254
rect 15694 4252 15700 4254
rect 15764 4252 15770 4316
rect 15878 4252 15884 4316
rect 15948 4314 15995 4316
rect 15948 4312 16040 4314
rect 15990 4256 16040 4312
rect 15948 4254 16040 4256
rect 15948 4252 15995 4254
rect 15929 4251 15995 4252
rect 11697 4178 11763 4181
rect 12525 4178 12591 4181
rect 11697 4176 12591 4178
rect 11697 4120 11702 4176
rect 11758 4120 12530 4176
rect 12586 4120 12591 4176
rect 11697 4118 12591 4120
rect 11697 4115 11763 4118
rect 12525 4115 12591 4118
rect 13353 4178 13419 4181
rect 24652 4178 24752 4208
rect 13353 4176 24752 4178
rect 13353 4120 13358 4176
rect 13414 4120 24752 4176
rect 13353 4118 24752 4120
rect 13353 4115 13419 4118
rect 24652 4088 24752 4118
rect 8017 4042 8083 4045
rect 9305 4042 9371 4045
rect 8017 4040 9371 4042
rect 8017 3984 8022 4040
rect 8078 3984 9310 4040
rect 9366 3984 9371 4040
rect 8017 3982 9371 3984
rect 8017 3979 8083 3982
rect 9305 3979 9371 3982
rect 12157 4042 12223 4045
rect 16205 4042 16271 4045
rect 12157 4040 16271 4042
rect 12157 3984 12162 4040
rect 12218 3984 16210 4040
rect 16266 3984 16271 4040
rect 12157 3982 16271 3984
rect 12157 3979 12223 3982
rect 16205 3979 16271 3982
rect 16389 4042 16455 4045
rect 18045 4042 18111 4045
rect 16389 4040 18111 4042
rect 16389 3984 16394 4040
rect 16450 3984 18050 4040
rect 18106 3984 18111 4040
rect 16389 3982 18111 3984
rect 16389 3979 16455 3982
rect 18045 3979 18111 3982
rect 11881 3906 11947 3909
rect 12341 3906 12407 3909
rect 13445 3906 13511 3909
rect 11881 3904 13511 3906
rect 11881 3848 11886 3904
rect 11942 3848 12346 3904
rect 12402 3848 13450 3904
rect 13506 3848 13511 3904
rect 11881 3846 13511 3848
rect 11881 3843 11947 3846
rect 12341 3843 12407 3846
rect 13445 3843 13511 3846
rect 14457 3906 14523 3909
rect 19057 3906 19123 3909
rect 14457 3904 19123 3906
rect 14457 3848 14462 3904
rect 14518 3848 19062 3904
rect 19118 3848 19123 3904
rect 14457 3846 19123 3848
rect 14457 3843 14523 3846
rect 19057 3843 19123 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 9213 3770 9279 3773
rect 9857 3770 9923 3773
rect 16021 3770 16087 3773
rect 16941 3770 17007 3773
rect 9213 3768 17007 3770
rect 9213 3712 9218 3768
rect 9274 3712 9862 3768
rect 9918 3712 16026 3768
rect 16082 3712 16946 3768
rect 17002 3712 17007 3768
rect 9213 3710 17007 3712
rect 9213 3707 9279 3710
rect 9857 3707 9923 3710
rect 16021 3707 16087 3710
rect 16941 3707 17007 3710
rect 10041 3634 10107 3637
rect 13169 3634 13235 3637
rect 15469 3636 15535 3637
rect 15469 3634 15516 3636
rect 10041 3632 13235 3634
rect 10041 3576 10046 3632
rect 10102 3576 13174 3632
rect 13230 3576 13235 3632
rect 10041 3574 13235 3576
rect 15424 3632 15516 3634
rect 15424 3576 15474 3632
rect 15424 3574 15516 3576
rect 10041 3571 10107 3574
rect 13169 3571 13235 3574
rect 15469 3572 15516 3574
rect 15580 3572 15586 3636
rect 15469 3571 15535 3572
rect 4613 3498 4679 3501
rect 13997 3498 14063 3501
rect 4613 3496 14063 3498
rect 4613 3440 4618 3496
rect 4674 3440 14002 3496
rect 14058 3440 14063 3496
rect 4613 3438 14063 3440
rect 4613 3435 4679 3438
rect 13997 3435 14063 3438
rect 14273 3498 14339 3501
rect 24652 3498 24752 3528
rect 14273 3496 24752 3498
rect 14273 3440 14278 3496
rect 14334 3440 24752 3496
rect 14273 3438 24752 3440
rect 14273 3435 14339 3438
rect 24652 3408 24752 3438
rect 12893 3362 12959 3365
rect 15101 3362 15167 3365
rect 12893 3360 15167 3362
rect 12893 3304 12898 3360
rect 12954 3304 15106 3360
rect 15162 3304 15167 3360
rect 12893 3302 15167 3304
rect 12893 3299 12959 3302
rect 15101 3299 15167 3302
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 13261 3226 13327 3229
rect 18229 3226 18295 3229
rect 22369 3226 22435 3229
rect 13261 3224 18295 3226
rect 13261 3168 13266 3224
rect 13322 3168 18234 3224
rect 18290 3168 18295 3224
rect 13261 3166 18295 3168
rect 13261 3163 13327 3166
rect 18229 3163 18295 3166
rect 22050 3224 22435 3226
rect 22050 3168 22374 3224
rect 22430 3168 22435 3224
rect 22050 3166 22435 3168
rect 7557 3090 7623 3093
rect 8569 3090 8635 3093
rect 7557 3088 8635 3090
rect 7557 3032 7562 3088
rect 7618 3032 8574 3088
rect 8630 3032 8635 3088
rect 7557 3030 8635 3032
rect 7557 3027 7623 3030
rect 8569 3027 8635 3030
rect 12249 3090 12315 3093
rect 14181 3090 14247 3093
rect 12249 3088 14247 3090
rect 12249 3032 12254 3088
rect 12310 3032 14186 3088
rect 14242 3032 14247 3088
rect 12249 3030 14247 3032
rect 12249 3027 12315 3030
rect 14181 3027 14247 3030
rect 10777 2954 10843 2957
rect 13445 2954 13511 2957
rect 18638 2954 18644 2956
rect 10777 2952 18644 2954
rect 10777 2896 10782 2952
rect 10838 2896 13450 2952
rect 13506 2896 18644 2952
rect 10777 2894 18644 2896
rect 10777 2891 10843 2894
rect 13445 2891 13511 2894
rect 18638 2892 18644 2894
rect 18708 2954 18714 2956
rect 22050 2954 22110 3166
rect 22369 3163 22435 3166
rect 18708 2894 22110 2954
rect 18708 2892 18714 2894
rect 0 2818 100 2848
rect 749 2818 815 2821
rect 0 2816 815 2818
rect 0 2760 754 2816
rect 810 2760 815 2816
rect 0 2758 815 2760
rect 0 2728 100 2758
rect 749 2755 815 2758
rect 10317 2818 10383 2821
rect 24652 2818 24752 2848
rect 10317 2816 24752 2818
rect 10317 2760 10322 2816
rect 10378 2760 24752 2816
rect 10317 2758 24752 2760
rect 10317 2755 10383 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 24652 2728 24752 2758
rect 4210 2687 4526 2688
rect 8753 2682 8819 2685
rect 10133 2682 10199 2685
rect 8753 2680 10199 2682
rect 8753 2624 8758 2680
rect 8814 2624 10138 2680
rect 10194 2624 10199 2680
rect 8753 2622 10199 2624
rect 8753 2619 8819 2622
rect 10133 2619 10199 2622
rect 15142 2620 15148 2684
rect 15212 2682 15218 2684
rect 22829 2682 22895 2685
rect 15212 2680 22895 2682
rect 15212 2624 22834 2680
rect 22890 2624 22895 2680
rect 15212 2622 22895 2624
rect 15212 2620 15218 2622
rect 22829 2619 22895 2622
rect 11053 2546 11119 2549
rect 15285 2546 15351 2549
rect 11053 2544 15351 2546
rect 11053 2488 11058 2544
rect 11114 2488 15290 2544
rect 15346 2488 15351 2544
rect 11053 2486 15351 2488
rect 11053 2483 11119 2486
rect 15285 2483 15351 2486
rect 21950 2484 21956 2548
rect 22020 2546 22026 2548
rect 22921 2546 22987 2549
rect 22020 2544 22987 2546
rect 22020 2488 22926 2544
rect 22982 2488 22987 2544
rect 22020 2486 22987 2488
rect 22020 2484 22026 2486
rect 22921 2483 22987 2486
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 21633 2138 21699 2141
rect 24652 2138 24752 2168
rect 21633 2136 24752 2138
rect 21633 2080 21638 2136
rect 21694 2080 24752 2136
rect 21633 2078 24752 2080
rect 21633 2075 21699 2078
rect 24652 2048 24752 2078
rect 8477 1866 8543 1869
rect 8477 1864 22110 1866
rect 8477 1808 8482 1864
rect 8538 1808 22110 1864
rect 8477 1806 22110 1808
rect 8477 1803 8543 1806
rect 22050 1458 22110 1806
rect 24652 1458 24752 1488
rect 22050 1398 24752 1458
rect 24652 1368 24752 1398
rect 23197 778 23263 781
rect 24652 778 24752 808
rect 23197 776 24752 778
rect 23197 720 23202 776
rect 23258 720 24752 776
rect 23197 718 24752 720
rect 23197 715 23263 718
rect 24652 688 24752 718
rect 9673 98 9739 101
rect 24652 98 24752 128
rect 9673 96 24752 98
rect 9673 40 9678 96
rect 9734 40 24752 96
rect 9673 38 24752 40
rect 9673 35 9739 38
rect 24652 8 24752 38
<< via3 >>
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 18828 10100 18892 10164
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 9260 9556 9324 9620
rect 18460 9692 18524 9756
rect 21956 9692 22020 9756
rect 17356 9420 17420 9484
rect 16620 9284 16684 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 17356 9208 17420 9212
rect 17356 9152 17370 9208
rect 17370 9152 17420 9208
rect 17356 9148 17420 9152
rect 16620 8936 16684 8940
rect 16620 8880 16670 8936
rect 16670 8880 16684 8936
rect 16620 8876 16684 8880
rect 16988 8876 17052 8940
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 14228 8604 14292 8668
rect 14780 8332 14844 8396
rect 13676 8196 13740 8260
rect 16988 8196 17052 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 14964 7924 15028 7988
rect 18644 7924 18708 7988
rect 15884 7712 15948 7716
rect 15884 7656 15934 7712
rect 15934 7656 15948 7712
rect 15884 7652 15948 7656
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 15516 6972 15580 7036
rect 16620 6896 16684 6900
rect 16620 6840 16634 6896
rect 16634 6840 16684 6896
rect 16620 6836 16684 6840
rect 14044 6700 14108 6764
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 14964 6352 15028 6356
rect 14964 6296 14978 6352
rect 14978 6296 15028 6352
rect 14964 6292 15028 6296
rect 15700 6292 15764 6356
rect 16620 6020 16684 6084
rect 18828 6080 18892 6084
rect 18828 6024 18842 6080
rect 18842 6024 18892 6080
rect 18828 6020 18892 6024
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 13676 5944 13740 5948
rect 13676 5888 13726 5944
rect 13726 5888 13740 5944
rect 13676 5884 13740 5888
rect 17908 5884 17972 5948
rect 14044 5612 14108 5676
rect 15148 5612 15212 5676
rect 18460 5612 18524 5676
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 17908 5204 17972 5268
rect 14780 5068 14844 5132
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 9260 4720 9324 4724
rect 9260 4664 9274 4720
rect 9274 4664 9324 4720
rect 9260 4660 9324 4664
rect 14228 4524 14292 4588
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 15700 4252 15764 4316
rect 15884 4312 15948 4316
rect 15884 4256 15934 4312
rect 15934 4256 15948 4312
rect 15884 4252 15948 4256
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 15516 3632 15580 3636
rect 15516 3576 15530 3632
rect 15530 3576 15580 3632
rect 15516 3572 15580 3576
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 18644 2892 18708 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 15148 2620 15212 2684
rect 21956 2484 22020 2548
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 10368 4528 10928
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 10912 5188 10928
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 18827 10164 18893 10165
rect 18827 10100 18828 10164
rect 18892 10100 18893 10164
rect 18827 10099 18893 10100
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 18459 9756 18525 9757
rect 18459 9692 18460 9756
rect 18524 9692 18525 9756
rect 18459 9691 18525 9692
rect 9259 9620 9325 9621
rect 9259 9556 9260 9620
rect 9324 9556 9325 9620
rect 9259 9555 9325 9556
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 9262 4725 9322 9555
rect 17355 9484 17421 9485
rect 17355 9420 17356 9484
rect 17420 9420 17421 9484
rect 17355 9419 17421 9420
rect 16619 9348 16685 9349
rect 16619 9284 16620 9348
rect 16684 9284 16685 9348
rect 16619 9283 16685 9284
rect 16622 8941 16682 9283
rect 17358 9213 17418 9419
rect 17355 9212 17421 9213
rect 17355 9148 17356 9212
rect 17420 9148 17421 9212
rect 17355 9147 17421 9148
rect 16619 8940 16685 8941
rect 16619 8876 16620 8940
rect 16684 8876 16685 8940
rect 16619 8875 16685 8876
rect 16987 8940 17053 8941
rect 16987 8876 16988 8940
rect 17052 8876 17053 8940
rect 16987 8875 17053 8876
rect 14227 8668 14293 8669
rect 14227 8604 14228 8668
rect 14292 8604 14293 8668
rect 14227 8603 14293 8604
rect 13675 8260 13741 8261
rect 13675 8196 13676 8260
rect 13740 8196 13741 8260
rect 13675 8195 13741 8196
rect 13678 5949 13738 8195
rect 14043 6764 14109 6765
rect 14043 6700 14044 6764
rect 14108 6700 14109 6764
rect 14043 6699 14109 6700
rect 13675 5948 13741 5949
rect 13675 5884 13676 5948
rect 13740 5884 13741 5948
rect 13675 5883 13741 5884
rect 14046 5677 14106 6699
rect 14043 5676 14109 5677
rect 14043 5612 14044 5676
rect 14108 5612 14109 5676
rect 14043 5611 14109 5612
rect 9259 4724 9325 4725
rect 9259 4660 9260 4724
rect 9324 4660 9325 4724
rect 9259 4659 9325 4660
rect 14230 4589 14290 8603
rect 14779 8396 14845 8397
rect 14779 8332 14780 8396
rect 14844 8332 14845 8396
rect 14779 8331 14845 8332
rect 14782 5133 14842 8331
rect 16990 8261 17050 8875
rect 16987 8260 17053 8261
rect 16987 8196 16988 8260
rect 17052 8196 17053 8260
rect 16987 8195 17053 8196
rect 14963 7988 15029 7989
rect 14963 7924 14964 7988
rect 15028 7924 15029 7988
rect 14963 7923 15029 7924
rect 14966 6357 15026 7923
rect 15883 7716 15949 7717
rect 15883 7652 15884 7716
rect 15948 7652 15949 7716
rect 15883 7651 15949 7652
rect 15515 7036 15581 7037
rect 15515 6972 15516 7036
rect 15580 6972 15581 7036
rect 15515 6971 15581 6972
rect 14963 6356 15029 6357
rect 14963 6292 14964 6356
rect 15028 6292 15029 6356
rect 14963 6291 15029 6292
rect 15147 5676 15213 5677
rect 15147 5612 15148 5676
rect 15212 5612 15213 5676
rect 15147 5611 15213 5612
rect 14779 5132 14845 5133
rect 14779 5068 14780 5132
rect 14844 5068 14845 5132
rect 14779 5067 14845 5068
rect 14227 4588 14293 4589
rect 14227 4524 14228 4588
rect 14292 4524 14293 4588
rect 14227 4523 14293 4524
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 15150 2685 15210 5611
rect 15518 3637 15578 6971
rect 15699 6356 15765 6357
rect 15699 6292 15700 6356
rect 15764 6292 15765 6356
rect 15699 6291 15765 6292
rect 15702 4317 15762 6291
rect 15886 4317 15946 7651
rect 16619 6900 16685 6901
rect 16619 6836 16620 6900
rect 16684 6836 16685 6900
rect 16619 6835 16685 6836
rect 16622 6085 16682 6835
rect 16619 6084 16685 6085
rect 16619 6020 16620 6084
rect 16684 6020 16685 6084
rect 16619 6019 16685 6020
rect 17907 5948 17973 5949
rect 17907 5884 17908 5948
rect 17972 5884 17973 5948
rect 17907 5883 17973 5884
rect 17910 5269 17970 5883
rect 18462 5677 18522 9691
rect 18643 7988 18709 7989
rect 18643 7924 18644 7988
rect 18708 7924 18709 7988
rect 18643 7923 18709 7924
rect 18459 5676 18525 5677
rect 18459 5612 18460 5676
rect 18524 5612 18525 5676
rect 18459 5611 18525 5612
rect 17907 5268 17973 5269
rect 17907 5204 17908 5268
rect 17972 5204 17973 5268
rect 17907 5203 17973 5204
rect 15699 4316 15765 4317
rect 15699 4252 15700 4316
rect 15764 4252 15765 4316
rect 15699 4251 15765 4252
rect 15883 4316 15949 4317
rect 15883 4252 15884 4316
rect 15948 4252 15949 4316
rect 15883 4251 15949 4252
rect 15515 3636 15581 3637
rect 15515 3572 15516 3636
rect 15580 3572 15581 3636
rect 15515 3571 15581 3572
rect 18646 2957 18706 7923
rect 18830 6085 18890 10099
rect 21955 9756 22021 9757
rect 21955 9692 21956 9756
rect 22020 9692 22021 9756
rect 21955 9691 22021 9692
rect 18827 6084 18893 6085
rect 18827 6020 18828 6084
rect 18892 6020 18893 6084
rect 18827 6019 18893 6020
rect 18643 2956 18709 2957
rect 18643 2892 18644 2956
rect 18708 2892 18709 2956
rect 18643 2891 18709 2892
rect 15147 2684 15213 2685
rect 15147 2620 15148 2684
rect 15212 2620 15213 2684
rect 15147 2619 15213 2620
rect 21958 2549 22018 9691
rect 21955 2548 22021 2549
rect 21955 2484 21956 2548
rect 22020 2484 22021 2548
rect 21955 2483 22021 2484
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1704896540
transform -1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1704896540
transform 1 0 15732 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1704896540
transform 1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1704896540
transform -1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1704896540
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1704896540
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1704896540
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _259_
timestamp 1704896540
transform -1 0 8372 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1704896540
transform 1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16284 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _263_
timestamp 1704896540
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1704896540
transform -1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18676 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1704896540
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14260 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13340 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1704896540
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _272_
timestamp 1704896540
transform 1 0 18676 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22908 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _274_
timestamp 1704896540
transform -1 0 19780 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _275_
timestamp 1704896540
transform 1 0 19780 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _276_
timestamp 1704896540
transform 1 0 17848 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _277_
timestamp 1704896540
transform 1 0 4600 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _278_
timestamp 1704896540
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7452 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _283_
timestamp 1704896540
transform 1 0 4692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _284_
timestamp 1704896540
transform 1 0 14260 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _286_
timestamp 1704896540
transform -1 0 5428 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _288_
timestamp 1704896540
transform 1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _289_
timestamp 1704896540
transform 1 0 4048 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _290_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14536 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _291_
timestamp 1704896540
transform -1 0 4968 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _292_
timestamp 1704896540
transform 1 0 2576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _295_
timestamp 1704896540
transform -1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _296_
timestamp 1704896540
transform -1 0 7636 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _297_
timestamp 1704896540
transform -1 0 16468 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _298_
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _299_
timestamp 1704896540
transform 1 0 7544 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _300_
timestamp 1704896540
transform -1 0 15732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _301_
timestamp 1704896540
transform 1 0 14812 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _302_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1704896540
transform -1 0 8648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _304_
timestamp 1704896540
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _305_
timestamp 1704896540
transform -1 0 14720 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _306_
timestamp 1704896540
transform -1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _309_
timestamp 1704896540
transform 1 0 5336 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _310_
timestamp 1704896540
transform 1 0 7176 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _312_
timestamp 1704896540
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_2  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8464 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1704896540
transform 1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _318_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _319_
timestamp 1704896540
transform 1 0 15272 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _320_
timestamp 1704896540
transform -1 0 9936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16008 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _322_
timestamp 1704896540
transform -1 0 16008 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _324_
timestamp 1704896540
transform 1 0 14076 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _325_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14076 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _326_
timestamp 1704896540
transform -1 0 15180 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _327_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15272 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _328_
timestamp 1704896540
transform 1 0 15364 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _329_
timestamp 1704896540
transform 1 0 16008 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _331_
timestamp 1704896540
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1704896540
transform 1 0 12052 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _333_
timestamp 1704896540
transform -1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _334_
timestamp 1704896540
transform -1 0 12328 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11132 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _336_
timestamp 1704896540
transform -1 0 15548 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _337_
timestamp 1704896540
transform -1 0 15272 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _338_
timestamp 1704896540
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _339_
timestamp 1704896540
transform -1 0 15364 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _340_
timestamp 1704896540
transform -1 0 15180 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _341_
timestamp 1704896540
transform -1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _342_
timestamp 1704896540
transform -1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_2  _343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3404 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a32oi_1  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10304 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _345_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10212 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_2  _346_
timestamp 1704896540
transform 1 0 6900 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _347_
timestamp 1704896540
transform -1 0 8832 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _349_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9936 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _351_
timestamp 1704896540
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _352_
timestamp 1704896540
transform 1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _353_
timestamp 1704896540
transform -1 0 9108 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _354_
timestamp 1704896540
transform -1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _355_
timestamp 1704896540
transform -1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _356_
timestamp 1704896540
transform -1 0 8004 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _358_
timestamp 1704896540
transform -1 0 9844 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _360_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10856 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _361_
timestamp 1704896540
transform -1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _362_
timestamp 1704896540
transform -1 0 16560 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _363_
timestamp 1704896540
transform 1 0 17664 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _364__1
timestamp 1704896540
transform -1 0 12328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _365_
timestamp 1704896540
transform -1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _366_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__o32a_2  _367_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15732 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _368_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16468 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _369_
timestamp 1704896540
transform 1 0 15916 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_4  _370_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17388 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _371__2
timestamp 1704896540
transform -1 0 16560 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371__3
timestamp 1704896540
transform -1 0 21528 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16560 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _373_
timestamp 1704896540
transform 1 0 17204 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _374_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21528 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _375_
timestamp 1704896540
transform -1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _376_
timestamp 1704896540
transform -1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _377_
timestamp 1704896540
transform -1 0 18768 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _378_
timestamp 1704896540
transform -1 0 17664 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _379_
timestamp 1704896540
transform 1 0 17940 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _380_
timestamp 1704896540
transform 1 0 21804 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _381_
timestamp 1704896540
transform 1 0 17480 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _382_
timestamp 1704896540
transform -1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18768 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _384_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19412 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _385_
timestamp 1704896540
transform 1 0 16468 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _386_
timestamp 1704896540
transform 1 0 15456 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _387_
timestamp 1704896540
transform -1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _388_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 20700 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_4  _389_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_2  _390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20516 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _391_
timestamp 1704896540
transform -1 0 9200 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1704896540
transform 1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _393_
timestamp 1704896540
transform 1 0 5796 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1704896540
transform 1 0 7176 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _395_
timestamp 1704896540
transform 1 0 6532 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _396_
timestamp 1704896540
transform -1 0 6900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _397_
timestamp 1704896540
transform -1 0 8832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8832 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _401_
timestamp 1704896540
transform -1 0 9936 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _402_
timestamp 1704896540
transform 1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _403_
timestamp 1704896540
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1704896540
transform 1 0 12880 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _405_
timestamp 1704896540
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _406_
timestamp 1704896540
transform 1 0 9660 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _407_
timestamp 1704896540
transform -1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _408_
timestamp 1704896540
transform 1 0 10948 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _409_
timestamp 1704896540
transform 1 0 10580 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _410_
timestamp 1704896540
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _411_
timestamp 1704896540
transform 1 0 9108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _412_
timestamp 1704896540
transform -1 0 10120 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _413_
timestamp 1704896540
transform 1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _414_
timestamp 1704896540
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _415_
timestamp 1704896540
transform -1 0 10856 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_2  _416_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9936 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and4_2  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _418_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _419_
timestamp 1704896540
transform 1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _420_
timestamp 1704896540
transform -1 0 5336 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1704896540
transform 1 0 4048 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp 1704896540
transform 1 0 3956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _423_
timestamp 1704896540
transform -1 0 4508 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _424_
timestamp 1704896540
transform -1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _425_
timestamp 1704896540
transform 1 0 4140 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _426_
timestamp 1704896540
transform -1 0 4416 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _427_
timestamp 1704896540
transform 1 0 4600 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _428_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5060 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _429_
timestamp 1704896540
transform -1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _430_
timestamp 1704896540
transform 1 0 15272 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _431_
timestamp 1704896540
transform -1 0 16284 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _432_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _433_
timestamp 1704896540
transform 1 0 12972 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _434_
timestamp 1704896540
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _436_
timestamp 1704896540
transform -1 0 7728 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _437_
timestamp 1704896540
transform -1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _438_
timestamp 1704896540
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _439_
timestamp 1704896540
transform 1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _440_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _441_
timestamp 1704896540
transform 1 0 11500 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _442_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13156 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _443_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _444_
timestamp 1704896540
transform -1 0 11500 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _445_
timestamp 1704896540
transform -1 0 13064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _446_
timestamp 1704896540
transform 1 0 11960 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _447_
timestamp 1704896540
transform 1 0 10396 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _448_
timestamp 1704896540
transform -1 0 11408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _449_
timestamp 1704896540
transform 1 0 11960 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _450_
timestamp 1704896540
transform 1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _451_
timestamp 1704896540
transform -1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _452_
timestamp 1704896540
transform -1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _453_
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1704896540
transform 1 0 13156 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _455_
timestamp 1704896540
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _456_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12236 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _457_
timestamp 1704896540
transform -1 0 12144 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _458_
timestamp 1704896540
transform 1 0 12052 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _459_
timestamp 1704896540
transform 1 0 17756 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1704896540
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_2  _461_
timestamp 1704896540
transform -1 0 18860 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _462_
timestamp 1704896540
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _463_
timestamp 1704896540
transform 1 0 23000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _464_
timestamp 1704896540
transform 1 0 22264 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _465_
timestamp 1704896540
transform -1 0 23000 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _466_
timestamp 1704896540
transform 1 0 22264 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _467_
timestamp 1704896540
transform -1 0 23000 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _468_
timestamp 1704896540
transform -1 0 23276 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _469_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23368 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _470_
timestamp 1704896540
transform -1 0 23368 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _471_
timestamp 1704896540
transform -1 0 4692 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _472_
timestamp 1704896540
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _474_
timestamp 1704896540
transform 1 0 3404 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _475_
timestamp 1704896540
transform 1 0 3036 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _476_
timestamp 1704896540
transform -1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _477_
timestamp 1704896540
transform 1 0 4968 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _478_
timestamp 1704896540
transform 1 0 5244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _479_
timestamp 1704896540
transform 1 0 5520 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _480_
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _481_
timestamp 1704896540
transform -1 0 6532 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _482_
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _483_
timestamp 1704896540
transform -1 0 15364 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _484_
timestamp 1704896540
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _485_
timestamp 1704896540
transform 1 0 12328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _486_
timestamp 1704896540
transform -1 0 13800 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _487_
timestamp 1704896540
transform -1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _488_
timestamp 1704896540
transform 1 0 13064 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _489_
timestamp 1704896540
transform -1 0 12052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _490_
timestamp 1704896540
transform 1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _491_
timestamp 1704896540
transform -1 0 13156 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _492_
timestamp 1704896540
transform 1 0 12880 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _493_
timestamp 1704896540
transform -1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_2  _494_
timestamp 1704896540
transform -1 0 13064 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _495_
timestamp 1704896540
transform -1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _496_
timestamp 1704896540
transform -1 0 21712 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _497_
timestamp 1704896540
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _498_
timestamp 1704896540
transform -1 0 22908 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _499_
timestamp 1704896540
transform -1 0 14536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _500_
timestamp 1704896540
transform -1 0 23368 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 23368 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_2  _502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21804 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _503_
timestamp 1704896540
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _504_
timestamp 1704896540
transform -1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _505_
timestamp 1704896540
transform 1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _506_
timestamp 1704896540
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_2  _507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 22632 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21804 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__a21oi_2  _509_
timestamp 1704896540
transform 1 0 21804 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _510_
timestamp 1704896540
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 22908 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _512_
timestamp 1704896540
transform -1 0 21712 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _513_
timestamp 1704896540
transform 1 0 16652 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _514_
timestamp 1704896540
transform -1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_1  _515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14720 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _517_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ba_1  _518_
timestamp 1704896540
transform -1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_1  _519_
timestamp 1704896540
transform -1 0 14352 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _520_
timestamp 1704896540
transform -1 0 17572 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_2  _521_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20148 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _522_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 19872 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _523_
timestamp 1704896540
transform -1 0 19136 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_2  _524_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _525_
timestamp 1704896540
transform 1 0 15456 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _526_
timestamp 1704896540
transform -1 0 13432 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _528_
timestamp 1704896540
transform -1 0 15364 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _529_
timestamp 1704896540
transform 1 0 19320 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _535_
timestamp 1704896540
transform 1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _536_
timestamp 1704896540
transform 1 0 23000 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _537_
timestamp 1704896540
transform 1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _538_
timestamp 1704896540
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _539_
timestamp 1704896540
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _540_
timestamp 1704896540
transform -1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _541_
timestamp 1704896540
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1704896540
transform -1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1704896540
transform -1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _544_
timestamp 1704896540
transform -1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _545_
timestamp 1704896540
transform -1 0 13984 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _546_
timestamp 1704896540
transform 1 0 17848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1704896540
transform 1 0 19964 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1704896540
transform 1 0 18768 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1704896540
transform -1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1704896540
transform -1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1704896540
transform -1 0 8556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1704896540
transform -1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1704896540
transform -1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1704896540
transform -1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1704896540
transform -1 0 13708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19228 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__081_
timestamp 1704896540
transform 1 0 18308 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__084_
timestamp 1704896540
transform 1 0 18308 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__091_
timestamp 1704896540
transform 1 0 21068 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__092_
timestamp 1704896540
transform -1 0 21068 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__235_
timestamp 1704896540
transform -1 0 19320 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__243_
timestamp 1704896540
transform -1 0 17020 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1704896540
transform -1 0 21712 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__079_
timestamp 1704896540
transform -1 0 19136 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__081_
timestamp 1704896540
transform -1 0 19044 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__084_
timestamp 1704896540
transform -1 0 16560 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__091_
timestamp 1704896540
transform -1 0 22908 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__092_
timestamp 1704896540
transform 1 0 19228 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__106_
timestamp 1704896540
transform 1 0 19872 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__235_
timestamp 1704896540
transform -1 0 18492 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__243_
timestamp 1704896540
transform -1 0 14904 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 16560 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__079_
timestamp 1704896540
transform 1 0 21068 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__081_
timestamp 1704896540
transform 1 0 19228 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__084_
timestamp 1704896540
transform -1 0 19412 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__088_
timestamp 1704896540
transform 1 0 21528 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__091_
timestamp 1704896540
transform -1 0 22080 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__092_
timestamp 1704896540
transform -1 0 19872 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__106_
timestamp 1704896540
transform 1 0 19964 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__235_
timestamp 1704896540
transform 1 0 19228 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__243_
timestamp 1704896540
transform 1 0 17664 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 21068 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15916 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 1704896540
transform -1 0 13984 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  clkload2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17020 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 20148 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_8  clkload4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 19964 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  clkload5
timestamp 1704896540
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  clkload6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 21528 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  clkload7
timestamp 1704896540
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  clkload8
timestamp 1704896540
transform -1 0 15640 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  clkload9
timestamp 1704896540
transform -1 0 17756 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout67 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp 1704896540
transform 1 0 23000 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 1704896540
transform -1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 1704896540
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp 1704896540
transform 1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 1704896540
transform -1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 1704896540
transform -1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout75 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13616 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1704896540
transform -1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout77
timestamp 1704896540
transform -1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout79
timestamp 1704896540
transform -1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout80
timestamp 1704896540
transform -1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 1704896540
transform -1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 1704896540
transform -1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout83
timestamp 1704896540
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1704896540
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124
timestamp 1704896540
transform 1 0 12512 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6
timestamp 1704896540
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_18
timestamp 1704896540
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_30
timestamp 1704896540
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_42
timestamp 1704896540
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1704896540
transform 1 0 10212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp 1704896540
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp 1704896540
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_232
timestamp 1704896540
transform 1 0 22448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_241
timestamp 1704896540
transform 1 0 23276 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_75
timestamp 1704896540
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1704896540
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_148
timestamp 1704896540
transform 1 0 14720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 1704896540
transform 1 0 16376 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1704896540
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1704896540
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_73
timestamp 1704896540
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_94
timestamp 1704896540
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1704896540
transform 1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp 1704896540
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1704896540
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_45
timestamp 1704896540
transform 1 0 5244 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_51
timestamp 1704896540
transform 1 0 5796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_59
timestamp 1704896540
transform 1 0 6532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1704896540
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_74
timestamp 1704896540
transform 1 0 7912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1704896540
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_89
timestamp 1704896540
transform 1 0 9292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_101
timestamp 1704896540
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 1704896540
transform 1 0 11592 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_130
timestamp 1704896540
transform 1 0 13064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_148
timestamp 1704896540
transform 1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1704896540
transform 1 0 22908 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 1704896540
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1704896540
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_82
timestamp 1704896540
transform 1 0 8648 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_94
timestamp 1704896540
transform 1 0 9752 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_106
timestamp 1704896540
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1704896540
transform 1 0 12420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_132
timestamp 1704896540
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1704896540
transform 1 0 1748 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_12
timestamp 1704896540
transform 1 0 2208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1704896540
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1704896540
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 1704896540
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_69
timestamp 1704896540
transform 1 0 7452 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_77
timestamp 1704896540
transform 1 0 8188 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1704896540
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1704896540
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_112
timestamp 1704896540
transform 1 0 11408 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1704896540
transform 1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1704896540
transform 1 0 12696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_133
timestamp 1704896540
transform 1 0 13340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1704896540
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_175
timestamp 1704896540
transform 1 0 17204 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_217
timestamp 1704896540
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1704896540
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_12
timestamp 1704896540
transform 1 0 2208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp 1704896540
transform 1 0 3312 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1704896540
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_81
timestamp 1704896540
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp 1704896540
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1704896540
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1704896540
transform 1 0 12788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_145
timestamp 1704896540
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_155
timestamp 1704896540
transform 1 0 15364 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_199
timestamp 1704896540
transform 1 0 19412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1704896540
transform 1 0 19964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1704896540
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_37
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_59
timestamp 1704896540
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp 1704896540
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 1704896540
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_91
timestamp 1704896540
transform 1 0 9476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1704896540
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1704896540
transform 1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_176
timestamp 1704896540
transform 1 0 17296 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_237
timestamp 1704896540
transform 1 0 22908 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7
timestamp 1704896540
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_19
timestamp 1704896540
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_37
timestamp 1704896540
transform 1 0 4508 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_64
timestamp 1704896540
transform 1 0 6992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_76
timestamp 1704896540
transform 1 0 8096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1704896540
transform 1 0 8464 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_95
timestamp 1704896540
transform 1 0 9844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1704896540
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_121
timestamp 1704896540
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_203
timestamp 1704896540
transform 1 0 19780 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1704896540
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_13
timestamp 1704896540
transform 1 0 2300 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp 1704896540
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_40
timestamp 1704896540
transform 1 0 4784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1704896540
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_101
timestamp 1704896540
transform 1 0 10396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_113
timestamp 1704896540
transform 1 0 11500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1704896540
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_167
timestamp 1704896540
transform 1 0 16468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_237
timestamp 1704896540
transform 1 0 22908 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_241
timestamp 1704896540
transform 1 0 23276 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1704896540
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_23
timestamp 1704896540
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_42
timestamp 1704896540
transform 1 0 4968 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1704896540
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1704896540
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_61
timestamp 1704896540
transform 1 0 6716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_73
timestamp 1704896540
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_81
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_97
timestamp 1704896540
transform 1 0 10028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1704896540
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_116
timestamp 1704896540
transform 1 0 11776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_121
timestamp 1704896540
transform 1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_128
timestamp 1704896540
transform 1 0 12880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1704896540
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_163
timestamp 1704896540
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1704896540
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_241
timestamp 1704896540
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1704896540
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1704896540
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_51
timestamp 1704896540
transform 1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_63
timestamp 1704896540
transform 1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1704896540
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1704896540
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_92
timestamp 1704896540
transform 1 0 9568 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_98
timestamp 1704896540
transform 1 0 10120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_108
timestamp 1704896540
transform 1 0 11040 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1704896540
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_153
timestamp 1704896540
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1704896540
transform 1 0 22080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_241
timestamp 1704896540
transform 1 0 23276 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_12
timestamp 1704896540
transform 1 0 2208 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_24
timestamp 1704896540
transform 1 0 3312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_30
timestamp 1704896540
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_40
timestamp 1704896540
transform 1 0 4784 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_84
timestamp 1704896540
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1704896540
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1704896540
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1704896540
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1704896540
transform 1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1704896540
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1704896540
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_172
timestamp 1704896540
transform 1 0 16928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_204
timestamp 1704896540
transform 1 0 19872 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1704896540
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1704896540
transform 1 0 22080 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1704896540
transform 1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_12
timestamp 1704896540
transform 1 0 2208 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1704896540
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1704896540
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_50
timestamp 1704896540
transform 1 0 5704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1704896540
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1704896540
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_106
timestamp 1704896540
transform 1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_122
timestamp 1704896540
transform 1 0 12328 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_133
timestamp 1704896540
transform 1 0 13340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_153
timestamp 1704896540
transform 1 0 15180 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1704896540
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1704896540
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1704896540
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_225
timestamp 1704896540
transform 1 0 21804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_10
timestamp 1704896540
transform 1 0 2024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_22
timestamp 1704896540
transform 1 0 3128 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_29
timestamp 1704896540
transform 1 0 3772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_37
timestamp 1704896540
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1704896540
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1704896540
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1704896540
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_81
timestamp 1704896540
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1704896540
transform 1 0 8924 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 1704896540
transform 1 0 9384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_98
timestamp 1704896540
transform 1 0 10120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1704896540
transform 1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1704896540
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_118
timestamp 1704896540
transform 1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_139
timestamp 1704896540
transform 1 0 13892 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1704896540
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_160
timestamp 1704896540
transform 1 0 15824 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1704896540
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1704896540
transform 1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 1704896540
transform 1 0 22172 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1704896540
transform 1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform -1 0 14168 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform -1 0 13984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 23000 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1704896540
transform -1 0 13984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform -1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1704896540
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1704896540
transform -1 0 17664 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1704896540
transform -1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1704896540
transform -1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1704896540
transform -1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1704896540
transform 1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1704896540
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1704896540
transform -1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1704896540
transform -1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21804 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1704896540
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1704896540
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1704896540
transform 1 0 11040 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1704896540
transform 1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1704896540
transform 1 0 12972 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1704896540
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1704896540
transform 1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1704896540
transform -1 0 21160 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1704896540
transform 1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1704896540
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1704896540
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1704896540
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  main_84 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  main_85
timestamp 1704896540
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  main_86
timestamp 1704896540
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output36
timestamp 1704896540
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output37
timestamp 1704896540
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1704896540
transform 1 0 23000 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output39
timestamp 1704896540
transform 1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output40
timestamp 1704896540
transform -1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output41
timestamp 1704896540
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output42
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1704896540
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1704896540
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1704896540
transform 1 0 14076 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1704896540
transform -1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1704896540
transform -1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1704896540
transform -1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1704896540
transform -1 0 10120 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1704896540
transform 1 0 23000 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1704896540
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1704896540
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1704896540
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1704896540
transform -1 0 16560 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1704896540
transform -1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1704896540
transform 1 0 21896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1704896540
transform 1 0 14904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output58
timestamp 1704896540
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output59
timestamp 1704896540
transform 1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output60
timestamp 1704896540
transform 1 0 23000 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  output61 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17848 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  output62
timestamp 1704896540
transform -1 0 15824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output63
timestamp 1704896540
transform 1 0 15916 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output64
timestamp 1704896540
transform -1 0 21620 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  output65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output66
timestamp 1704896540
transform 1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_16
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_17
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_18
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_19
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 23644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_20
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_21
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 23644 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_22
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_23
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 23644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_24
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_25
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 23644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_26
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_27
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 23644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_28
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_29
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 23644 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_30
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 23644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_31
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 23644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp 1704896540
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp 1704896540
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp 1704896540
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_44
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp 1704896540
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_48
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_49
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_50
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_51
timestamp 1704896540
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_52
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_53
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_54
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp 1704896540
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_56
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_57
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_58
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_59
timestamp 1704896540
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_60
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_61
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_62
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_63
timestamp 1704896540
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_64
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_65
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_66
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_67
timestamp 1704896540
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_68
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_69
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_70
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_71
timestamp 1704896540
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_72
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_73
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_74
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_75
timestamp 1704896540
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_76
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_77
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_78
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_79
timestamp 1704896540
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_80
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_81
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_82
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_83
timestamp 1704896540
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_84
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_85
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_86
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_87
timestamp 1704896540
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_88
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_89
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_90
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_91
timestamp 1704896540
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_92
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_94
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_95
timestamp 1704896540
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_96
timestamp 1704896540
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_97
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_98
timestamp 1704896540
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_99
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_100
timestamp 1704896540
transform 1 0 13984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_101
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_102
timestamp 1704896540
transform 1 0 19136 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_103
timestamp 1704896540
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
<< labels >>
flabel metal2 s 15474 0 15530 100 0 FreeSans 448 0 0 0 DAC6_conn
port 0 nsew signal output
flabel metal2 s 16762 0 16818 100 0 FreeSans 448 0 0 0 DAC8_conn
port 1 nsew signal output
flabel metal4 s 4868 2128 5188 10928 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 10928 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal3 s 24652 3408 24752 3528 0 FreeSans 480 0 0 0 a0
port 4 nsew signal input
flabel metal3 s 24652 688 24752 808 0 FreeSans 480 0 0 0 a0_sel
port 5 nsew signal output
flabel metal2 s 16118 0 16174 100 0 FreeSans 448 0 0 0 aux1_conn
port 6 nsew signal output
flabel metal2 s 11610 13270 11666 13370 0 FreeSans 448 0 0 0 aux2_conn
port 7 nsew signal output
flabel metal3 s 24652 8 24752 128 0 FreeSans 480 0 0 0 buffi_conn
port 8 nsew signal output
flabel metal2 s 18050 0 18106 100 0 FreeSans 448 0 0 0 buffo_conn
port 9 nsew signal output
flabel metal3 s 24652 2048 24752 2168 0 FreeSans 480 0 0 0 clk
port 10 nsew signal input
flabel metal3 s 24652 4768 24752 4888 0 FreeSans 480 0 0 0 compr1
port 11 nsew signal input
flabel metal3 s 24652 5448 24752 5568 0 FreeSans 480 0 0 0 compr2
port 12 nsew signal input
flabel metal3 s 24652 12928 24752 13048 0 FreeSans 480 0 0 0 flash_adc_inp[0]
port 13 nsew signal input
flabel metal3 s 24652 6128 24752 6248 0 FreeSans 480 0 0 0 flash_adc_inp[10]
port 14 nsew signal input
flabel metal3 s 24652 6808 24752 6928 0 FreeSans 480 0 0 0 flash_adc_inp[11]
port 15 nsew signal input
flabel metal3 s 24652 4088 24752 4208 0 FreeSans 480 0 0 0 flash_adc_inp[12]
port 16 nsew signal input
flabel metal3 s 24652 2728 24752 2848 0 FreeSans 480 0 0 0 flash_adc_inp[13]
port 17 nsew signal input
flabel metal3 s 24652 1368 24752 1488 0 FreeSans 480 0 0 0 flash_adc_inp[14]
port 18 nsew signal input
flabel metal3 s 24652 10888 24752 11008 0 FreeSans 480 0 0 0 flash_adc_inp[1]
port 19 nsew signal input
flabel metal3 s 24652 10208 24752 10328 0 FreeSans 480 0 0 0 flash_adc_inp[2]
port 20 nsew signal input
flabel metal3 s 24652 11568 24752 11688 0 FreeSans 480 0 0 0 flash_adc_inp[3]
port 21 nsew signal input
flabel metal3 s 24652 12248 24752 12368 0 FreeSans 480 0 0 0 flash_adc_inp[4]
port 22 nsew signal input
flabel metal3 s 24652 8848 24752 8968 0 FreeSans 480 0 0 0 flash_adc_inp[5]
port 23 nsew signal input
flabel metal3 s 24652 9528 24752 9648 0 FreeSans 480 0 0 0 flash_adc_inp[6]
port 24 nsew signal input
flabel metal3 s 24652 7488 24752 7608 0 FreeSans 480 0 0 0 flash_adc_inp[7]
port 25 nsew signal input
flabel metal3 s 24652 8168 24752 8288 0 FreeSans 480 0 0 0 flash_adc_inp[8]
port 26 nsew signal input
flabel metal2 s 24490 13270 24546 13370 0 FreeSans 448 0 0 0 flash_adc_inp[9]
port 27 nsew signal input
flabel metal2 s 19982 0 20038 100 0 FreeSans 448 0 0 0 rst_n
port 28 nsew signal input
flabel metal3 s 0 6808 100 6928 0 FreeSans 480 0 0 0 tern_dac[0]
port 29 nsew signal output
flabel metal2 s 14186 0 14242 100 0 FreeSans 448 0 0 0 tern_dac[10]
port 30 nsew signal output
flabel metal2 s 13542 13270 13598 13370 0 FreeSans 448 0 0 0 tern_dac[11]
port 31 nsew signal output
flabel metal2 s 16762 13270 16818 13370 0 FreeSans 448 0 0 0 tern_dac[12]
port 32 nsew signal output
flabel metal2 s 19338 13270 19394 13370 0 FreeSans 448 0 0 0 tern_dac[13]
port 33 nsew signal output
flabel metal2 s 17406 13270 17462 13370 0 FreeSans 448 0 0 0 tern_dac[14]
port 34 nsew signal output
flabel metal3 s 0 10888 100 11008 0 FreeSans 480 0 0 0 tern_dac[15]
port 35 nsew signal output
flabel metal3 s 0 2728 100 2848 0 FreeSans 480 0 0 0 tern_dac[16]
port 36 nsew signal output
flabel metal2 s 21914 0 21970 100 0 FreeSans 448 0 0 0 tern_dac[17]
port 37 nsew signal output
flabel metal2 s 9678 13270 9734 13370 0 FreeSans 448 0 0 0 tern_dac[1]
port 38 nsew signal output
flabel metal2 s 22558 13270 22614 13370 0 FreeSans 448 0 0 0 tern_dac[2]
port 39 nsew signal output
flabel metal3 s 0 9528 100 9648 0 FreeSans 480 0 0 0 tern_dac[3]
port 40 nsew signal output
flabel metal3 s 0 5448 100 5568 0 FreeSans 480 0 0 0 tern_dac[4]
port 41 nsew signal output
flabel metal3 s 0 10208 100 10328 0 FreeSans 480 0 0 0 tern_dac[5]
port 42 nsew signal output
flabel metal2 s 16118 13270 16174 13370 0 FreeSans 448 0 0 0 tern_dac[6]
port 43 nsew signal output
flabel metal2 s 14830 0 14886 100 0 FreeSans 448 0 0 0 tern_dac[7]
port 44 nsew signal output
flabel metal2 s 21914 13270 21970 13370 0 FreeSans 448 0 0 0 tern_dac[8]
port 45 nsew signal output
flabel metal2 s 14830 13270 14886 13370 0 FreeSans 448 0 0 0 tern_dac[9]
port 46 nsew signal output
flabel metal2 s 17406 0 17462 100 0 FreeSans 448 0 0 0 ternff_conn
port 47 nsew signal output
flabel metal3 s 0 7488 100 7608 0 FreeSans 480 0 0 0 ui_in[0]
port 48 nsew signal input
flabel metal3 s 0 6128 100 6248 0 FreeSans 480 0 0 0 ui_in[1]
port 49 nsew signal input
flabel metal2 s 4526 0 4582 100 0 FreeSans 448 0 0 0 ui_in[2]
port 50 nsew signal input
flabel metal2 s 5170 0 5226 100 0 FreeSans 448 0 0 0 ui_in[3]
port 51 nsew signal input
flabel metal2 s 10966 13270 11022 13370 0 FreeSans 448 0 0 0 ui_in[4]
port 52 nsew signal input
flabel metal2 s 14186 13270 14242 13370 0 FreeSans 448 0 0 0 ui_in[5]
port 53 nsew signal input
flabel metal2 s 12898 13270 12954 13370 0 FreeSans 448 0 0 0 ui_in[6]
port 54 nsew signal input
flabel metal2 s 12254 13270 12310 13370 0 FreeSans 448 0 0 0 ui_in[7]
port 55 nsew signal input
flabel metal2 s 18050 13270 18106 13370 0 FreeSans 448 0 0 0 uio_in[0]
port 56 nsew signal input
flabel metal2 s 18694 13270 18750 13370 0 FreeSans 448 0 0 0 uio_in[1]
port 57 nsew signal input
flabel metal3 s 0 4768 100 4888 0 FreeSans 480 0 0 0 uio_in[2]
port 58 nsew signal input
flabel metal2 s 9034 13270 9090 13370 0 FreeSans 448 0 0 0 uio_in[3]
port 59 nsew signal input
flabel metal2 s 3882 0 3938 100 0 FreeSans 448 0 0 0 uio_in[4]
port 60 nsew signal input
flabel metal2 s 5814 0 5870 100 0 FreeSans 448 0 0 0 uio_in[5]
port 61 nsew signal input
flabel metal2 s 7102 0 7158 100 0 FreeSans 448 0 0 0 uio_in[6]
port 62 nsew signal input
flabel metal2 s 7746 0 7802 100 0 FreeSans 448 0 0 0 uio_in[7]
port 63 nsew signal input
flabel metal2 s 23202 13270 23258 13370 0 FreeSans 448 0 0 0 uo_out[0]
port 64 nsew signal output
flabel metal2 s 23846 13270 23902 13370 0 FreeSans 448 0 0 0 uo_out[1]
port 65 nsew signal output
flabel metal2 s 20626 13270 20682 13370 0 FreeSans 448 0 0 0 uo_out[2]
port 66 nsew signal output
flabel metal2 s 15474 13270 15530 13370 0 FreeSans 448 0 0 0 uo_out[3]
port 67 nsew signal output
flabel metal2 s 21270 13270 21326 13370 0 FreeSans 448 0 0 0 uo_out[4]
port 68 nsew signal output
flabel metal2 s 19982 13270 20038 13370 0 FreeSans 448 0 0 0 uo_out[5]
port 69 nsew signal output
flabel metal2 s 19338 0 19394 100 0 FreeSans 448 0 0 0 uo_out[6]
port 70 nsew signal output
flabel metal2 s 18694 0 18750 100 0 FreeSans 448 0 0 0 uo_out[7]
port 71 nsew signal output
rlabel metal1 12374 10880 12374 10880 0 VGND
rlabel metal1 12374 10336 12374 10336 0 VPWR
rlabel metal2 15502 534 15502 534 0 DAC6_conn
rlabel metal2 11362 1666 11362 1666 0 DAC8_conn
rlabel metal1 7222 7922 7222 7922 0 _000_
rlabel metal1 13064 8466 13064 8466 0 _001_
rlabel metal1 14076 4522 14076 4522 0 _002_
rlabel metal2 5290 7004 5290 7004 0 _003_
rlabel metal1 6670 5304 6670 5304 0 _004_
rlabel metal1 6302 7242 6302 7242 0 _005_
rlabel metal1 6808 7514 6808 7514 0 _006_
rlabel metal2 5658 5151 5658 5151 0 _007_
rlabel metal1 15778 5202 15778 5202 0 _008_
rlabel metal1 4508 6154 4508 6154 0 _009_
rlabel metal2 3082 6477 3082 6477 0 _010_
rlabel metal2 5382 7582 5382 7582 0 _011_
rlabel metal1 6302 7820 6302 7820 0 _012_
rlabel metal1 6670 7990 6670 7990 0 _013_
rlabel metal1 6486 7820 6486 7820 0 _014_
rlabel metal2 14398 7650 14398 7650 0 _015_
rlabel metal1 11960 7922 11960 7922 0 _016_
rlabel metal1 8188 5882 8188 5882 0 _017_
rlabel metal1 14582 5202 14582 5202 0 _018_
rlabel metal1 15870 6188 15870 6188 0 _019_
rlabel metal2 5842 8806 5842 8806 0 _020_
rlabel metal2 8510 9418 8510 9418 0 _021_
rlabel metal3 16790 3876 16790 3876 0 _022_
rlabel metal1 13892 2346 13892 2346 0 _023_
rlabel metal1 5934 7854 5934 7854 0 _024_
rlabel metal2 7774 9554 7774 9554 0 _025_
rlabel metal1 7544 9690 7544 9690 0 _026_
rlabel metal1 6164 9894 6164 9894 0 _027_
rlabel metal1 7084 9146 7084 9146 0 _028_
rlabel metal1 6532 10030 6532 10030 0 _029_
rlabel metal1 9798 10030 9798 10030 0 _030_
rlabel metal2 9706 3264 9706 3264 0 _031_
rlabel via1 10346 7854 10346 7854 0 _032_
rlabel metal1 7544 3366 7544 3366 0 _033_
rlabel metal1 9591 7854 9591 7854 0 _034_
rlabel metal1 9016 8058 9016 8058 0 _035_
rlabel metal1 9568 9146 9568 9146 0 _036_
rlabel metal1 18216 8942 18216 8942 0 _037_
rlabel metal1 10120 10166 10120 10166 0 _038_
rlabel metal1 14858 9520 14858 9520 0 _039_
rlabel metal1 15180 7922 15180 7922 0 _040_
rlabel via1 14651 8534 14651 8534 0 _041_
rlabel metal2 14122 9078 14122 9078 0 _042_
rlabel metal1 12098 10064 12098 10064 0 _043_
rlabel metal2 14306 8874 14306 8874 0 _044_
rlabel via1 16054 9078 16054 9078 0 _045_
rlabel metal1 16146 9146 16146 9146 0 _046_
rlabel metal1 13889 9486 13889 9486 0 _047_
rlabel metal1 12466 9520 12466 9520 0 _048_
rlabel metal2 12558 9044 12558 9044 0 _049_
rlabel metal2 11822 9180 11822 9180 0 _050_
rlabel metal1 12558 7854 12558 7854 0 _051_
rlabel metal1 11822 9894 11822 9894 0 _052_
rlabel metal1 10626 9044 10626 9044 0 _053_
rlabel metal1 15272 6358 15272 6358 0 _054_
rlabel viali 14762 6290 14762 6290 0 _055_
rlabel metal1 13386 6188 13386 6188 0 _056_
rlabel metal1 18078 5168 18078 5168 0 _057_
rlabel metal2 17986 4913 17986 4913 0 _058_
rlabel metal2 14122 5797 14122 5797 0 _059_
rlabel metal1 10534 6970 10534 6970 0 _060_
rlabel metal2 4186 5491 4186 5491 0 _061_
rlabel metal1 10304 5814 10304 5814 0 _062_
rlabel metal1 9522 3502 9522 3502 0 _063_
rlabel metal1 8602 3468 8602 3468 0 _064_
rlabel metal1 9430 3706 9430 3706 0 _065_
rlabel metal1 9706 6800 9706 6800 0 _066_
rlabel metal1 10258 5644 10258 5644 0 _067_
rlabel metal2 9614 5984 9614 5984 0 _068_
rlabel metal1 8142 4080 8142 4080 0 _069_
rlabel metal2 9062 4386 9062 4386 0 _070_
rlabel metal2 8418 4726 8418 4726 0 _071_
rlabel metal1 8142 4624 8142 4624 0 _072_
rlabel metal2 8050 4148 8050 4148 0 _073_
rlabel metal1 10718 3502 10718 3502 0 _074_
rlabel metal2 8694 5610 8694 5610 0 _075_
rlabel metal1 10120 6426 10120 6426 0 _076_
rlabel metal1 10718 9146 10718 9146 0 _077_
rlabel metal2 20378 9231 20378 9231 0 _078_
rlabel via2 13294 3179 13294 3179 0 _079_
rlabel metal2 17618 5882 17618 5882 0 _080_
rlabel metal1 18308 4046 18308 4046 0 _081_
rlabel metal2 17526 5916 17526 5916 0 _083_
rlabel metal1 17664 4046 17664 4046 0 _084_
rlabel metal2 15870 4930 15870 4930 0 _085_
rlabel metal1 16836 3638 16836 3638 0 _086_
rlabel metal1 16284 4794 16284 4794 0 _087_
rlabel metal1 20746 6256 20746 6256 0 _088_
rlabel metal2 17250 4896 17250 4896 0 _090_
rlabel metal2 21114 6052 21114 6052 0 _091_
rlabel metal1 21068 6290 21068 6290 0 _092_
rlabel metal1 18860 6766 18860 6766 0 _093_
rlabel metal1 17894 8602 17894 8602 0 _094_
rlabel metal2 17756 8466 17756 8466 0 _095_
rlabel metal2 19734 7446 19734 7446 0 _096_
rlabel metal2 18998 8670 18998 8670 0 _097_
rlabel metal1 19366 8364 19366 8364 0 _098_
rlabel metal1 18170 8262 18170 8262 0 _099_
rlabel metal1 18584 8466 18584 8466 0 _100_
rlabel metal1 18768 8398 18768 8398 0 _101_
rlabel metal1 20286 8500 20286 8500 0 _102_
rlabel metal1 16422 5576 16422 5576 0 _103_
rlabel metal2 16146 5882 16146 5882 0 _104_
rlabel metal1 20102 6290 20102 6290 0 _105_
rlabel metal1 20056 6358 20056 6358 0 _106_
rlabel metal1 20654 8534 20654 8534 0 _107_
rlabel metal1 8372 9622 8372 9622 0 _108_
rlabel metal1 7130 9350 7130 9350 0 _109_
rlabel metal2 6118 9146 6118 9146 0 _110_
rlabel metal2 6762 9724 6762 9724 0 _111_
rlabel metal2 6394 9146 6394 9146 0 _112_
rlabel metal2 6854 9282 6854 9282 0 _113_
rlabel via2 9430 7395 9430 7395 0 _114_
rlabel metal1 9476 8466 9476 8466 0 _115_
rlabel metal1 9108 7174 9108 7174 0 _116_
rlabel metal1 9430 9588 9430 9588 0 _117_
rlabel metal1 10074 9486 10074 9486 0 _118_
rlabel metal1 12788 8806 12788 8806 0 _119_
rlabel metal2 12098 8432 12098 8432 0 _120_
rlabel metal2 12926 9928 12926 9928 0 _121_
rlabel metal2 10626 9724 10626 9724 0 _122_
rlabel metal1 10672 6290 10672 6290 0 _123_
rlabel metal1 9936 3570 9936 3570 0 _124_
rlabel metal1 11776 5746 11776 5746 0 _125_
rlabel metal2 10626 6528 10626 6528 0 _126_
rlabel metal2 8510 4471 8510 4471 0 _127_
rlabel metal2 10442 3672 10442 3672 0 _128_
rlabel metal1 12236 2414 12236 2414 0 _129_
rlabel metal1 8142 3978 8142 3978 0 _130_
rlabel metal1 8740 5882 8740 5882 0 _131_
rlabel metal1 10764 6834 10764 6834 0 _132_
rlabel metal2 18998 8993 18998 8993 0 _133_
rlabel metal1 19044 8058 19044 8058 0 _134_
rlabel metal1 4554 9554 4554 9554 0 _135_
rlabel metal1 4738 9894 4738 9894 0 _136_
rlabel metal2 4094 10336 4094 10336 0 _137_
rlabel metal1 4370 9418 4370 9418 0 _138_
rlabel metal2 5842 10234 5842 10234 0 _139_
rlabel metal1 6532 6766 6532 6766 0 _140_
rlabel metal2 4462 5372 4462 5372 0 _141_
rlabel metal1 4830 5236 4830 5236 0 _142_
rlabel metal1 4600 5202 4600 5202 0 _143_
rlabel metal1 5612 5338 5612 5338 0 _144_
rlabel metal1 12374 6256 12374 6256 0 _145_
rlabel metal1 15088 5882 15088 5882 0 _146_
rlabel metal2 15134 6222 15134 6222 0 _147_
rlabel metal1 13570 6222 13570 6222 0 _148_
rlabel metal2 13662 6596 13662 6596 0 _149_
rlabel metal1 13156 5678 13156 5678 0 _150_
rlabel metal1 12420 2414 12420 2414 0 _151_
rlabel metal1 11086 4148 11086 4148 0 _152_
rlabel metal1 12512 2278 12512 2278 0 _153_
rlabel metal2 11270 4114 11270 4114 0 _154_
rlabel metal2 10902 4318 10902 4318 0 _155_
rlabel metal1 12420 3502 12420 3502 0 _156_
rlabel metal1 12650 3536 12650 3536 0 _157_
rlabel metal1 12788 3162 12788 3162 0 _158_
rlabel metal1 12658 4250 12658 4250 0 _159_
rlabel metal1 12742 4080 12742 4080 0 _160_
rlabel metal2 13018 4216 13018 4216 0 _161_
rlabel metal1 12190 3502 12190 3502 0 _162_
rlabel metal1 11914 3706 11914 3706 0 _163_
rlabel metal1 11960 3502 11960 3502 0 _164_
rlabel metal2 12650 4114 12650 4114 0 _165_
rlabel metal1 12926 4794 12926 4794 0 _166_
rlabel metal2 11638 6324 11638 6324 0 _167_
rlabel metal2 13846 9180 13846 9180 0 _168_
rlabel metal2 12558 8228 12558 8228 0 _169_
rlabel metal1 12650 8024 12650 8024 0 _170_
rlabel metal1 12742 7888 12742 7888 0 _171_
rlabel metal1 11960 6766 11960 6766 0 _172_
rlabel metal2 12282 6460 12282 6460 0 _173_
rlabel metal1 22678 6358 22678 6358 0 _174_
rlabel metal2 18078 6545 18078 6545 0 _175_
rlabel metal2 22126 7174 22126 7174 0 _176_
rlabel metal2 19458 7888 19458 7888 0 _177_
rlabel via2 22770 6307 22770 6307 0 _178_
rlabel metal1 22770 10064 22770 10064 0 _179_
rlabel metal2 22494 9418 22494 9418 0 _180_
rlabel metal1 22816 8466 22816 8466 0 _181_
rlabel metal2 22310 8942 22310 8942 0 _182_
rlabel metal1 23092 3094 23092 3094 0 _183_
rlabel metal1 23138 3162 23138 3162 0 _184_
rlabel metal1 23092 5338 23092 5338 0 _185_
rlabel metal1 4094 8602 4094 8602 0 _186_
rlabel metal2 3818 8738 3818 8738 0 _187_
rlabel metal1 3680 9078 3680 9078 0 _188_
rlabel metal1 3358 8602 3358 8602 0 _189_
rlabel metal1 5980 8942 5980 8942 0 _190_
rlabel metal1 6348 7446 6348 7446 0 _191_
rlabel metal2 5566 5882 5566 5882 0 _192_
rlabel metal2 6026 4794 6026 4794 0 _193_
rlabel via1 6867 5270 6867 5270 0 _194_
rlabel metal1 5934 4624 5934 4624 0 _195_
rlabel metal1 6578 4794 6578 4794 0 _196_
rlabel metal1 8970 7208 8970 7208 0 _197_
rlabel metal1 14973 6086 14973 6086 0 _198_
rlabel metal1 12650 5712 12650 5712 0 _199_
rlabel metal1 12190 5882 12190 5882 0 _200_
rlabel metal1 13662 3706 13662 3706 0 _201_
rlabel metal2 13662 4420 13662 4420 0 _202_
rlabel metal2 12558 4029 12558 4029 0 _203_
rlabel metal1 12236 6154 12236 6154 0 _204_
rlabel metal2 13386 8058 13386 8058 0 _205_
rlabel metal1 13202 7990 13202 7990 0 _206_
rlabel metal1 12788 6766 12788 6766 0 _207_
rlabel metal2 12190 7072 12190 7072 0 _208_
rlabel metal2 22402 7327 22402 7327 0 _209_
rlabel metal1 16468 9146 16468 9146 0 _210_
rlabel metal1 22080 10574 22080 10574 0 _211_
rlabel via2 22402 10659 22402 10659 0 _212_
rlabel metal2 22862 10081 22862 10081 0 _213_
rlabel metal3 14789 5644 14789 5644 0 _214_
rlabel metal1 23092 7242 23092 7242 0 _215_
rlabel metal1 22586 7344 22586 7344 0 _216_
rlabel metal1 20700 4046 20700 4046 0 _217_
rlabel metal1 22310 4998 22310 4998 0 _218_
rlabel metal1 22724 4046 22724 4046 0 _219_
rlabel metal2 21850 6494 21850 6494 0 _220_
rlabel metal2 22126 4522 22126 4522 0 _221_
rlabel metal2 22678 4556 22678 4556 0 _222_
rlabel metal2 22862 3638 22862 3638 0 _223_
rlabel metal1 16652 7854 16652 7854 0 _224_
rlabel metal2 22954 9401 22954 9401 0 _225_
rlabel metal1 17388 6290 17388 6290 0 _226_
rlabel via1 21392 4114 21392 4114 0 _227_
rlabel metal1 14214 3468 14214 3468 0 _228_
rlabel metal2 20102 3638 20102 3638 0 _229_
rlabel metal1 22287 4114 22287 4114 0 _230_
rlabel metal2 13846 3196 13846 3196 0 _231_
rlabel metal1 16928 2618 16928 2618 0 _232_
rlabel metal1 19826 4114 19826 4114 0 _233_
rlabel metal1 19918 2414 19918 2414 0 _234_
rlabel metal1 19090 2618 19090 2618 0 _235_
rlabel metal1 23690 9860 23690 9860 0 _236_
rlabel metal1 2599 6630 2599 6630 0 _237_
rlabel metal1 7958 5338 7958 5338 0 _238_
rlabel metal1 15962 9894 15962 9894 0 _239_
rlabel metal1 17802 5270 17802 5270 0 _240_
rlabel metal2 5658 8636 5658 8636 0 _241_
rlabel metal2 12466 3570 12466 3570 0 _242_
rlabel metal2 20746 4080 20746 4080 0 _243_
rlabel metal1 10350 10030 10350 10030 0 _244_
rlabel metal1 4922 8806 4922 8806 0 _245_
rlabel metal1 4186 10608 4186 10608 0 _246_
rlabel metal1 15778 6154 15778 6154 0 _247_
rlabel metal2 9246 4641 9246 4641 0 _248_
rlabel metal1 7958 7888 7958 7888 0 _249_
rlabel metal2 14306 4131 14306 4131 0 a0
rlabel metal3 23951 748 23951 748 0 a0_sel
rlabel metal2 12190 1734 12190 1734 0 aux1_conn
rlabel metal1 11684 10778 11684 10778 0 aux2_conn
rlabel metal2 9706 1173 9706 1173 0 buffi_conn
rlabel metal2 10258 1700 10258 1700 0 buffo_conn
rlabel metal2 21666 2227 21666 2227 0 clk
rlabel metal2 20562 6868 20562 6868 0 clknet_0__079_
rlabel metal2 18998 4250 18998 4250 0 clknet_0__081_
rlabel metal2 19642 5134 19642 5134 0 clknet_0__084_
rlabel metal1 22632 6698 22632 6698 0 clknet_0__091_
rlabel metal2 19366 5644 19366 5644 0 clknet_0__092_
rlabel metal1 18630 3162 18630 3162 0 clknet_0__235_
rlabel metal2 15686 7276 15686 7276 0 clknet_0__243_
rlabel metal1 19642 2482 19642 2482 0 clknet_0_clk
rlabel metal1 16376 5338 16376 5338 0 clknet_1_0__leaf__079_
rlabel metal1 16698 3536 16698 3536 0 clknet_1_0__leaf__081_
rlabel metal1 15870 2618 15870 2618 0 clknet_1_0__leaf__084_
rlabel metal2 21390 5542 21390 5542 0 clknet_1_0__leaf__091_
rlabel metal1 22205 6222 22205 6222 0 clknet_1_0__leaf__092_
rlabel metal1 22172 5066 22172 5066 0 clknet_1_0__leaf__106_
rlabel metal1 16698 2312 16698 2312 0 clknet_1_0__leaf__235_
rlabel metal2 10258 9282 10258 9282 0 clknet_1_0__leaf__243_
rlabel metal1 15318 3162 15318 3162 0 clknet_1_0__leaf_clk
rlabel metal1 22954 6222 22954 6222 0 clknet_1_1__leaf__079_
rlabel metal2 16882 6460 16882 6460 0 clknet_1_1__leaf__081_
rlabel metal1 16376 4046 16376 4046 0 clknet_1_1__leaf__084_
rlabel metal1 22609 5678 22609 5678 0 clknet_1_1__leaf__088_
rlabel metal2 20746 8534 20746 8534 0 clknet_1_1__leaf__091_
rlabel metal1 21804 8466 21804 8466 0 clknet_1_1__leaf__092_
rlabel metal1 20102 9554 20102 9554 0 clknet_1_1__leaf__106_
rlabel metal1 20562 4692 20562 4692 0 clknet_1_1__leaf__235_
rlabel metal1 19458 2278 19458 2278 0 clknet_1_1__leaf__243_
rlabel metal1 22678 3502 22678 3502 0 clknet_1_1__leaf_clk
rlabel metal1 14306 4998 14306 4998 0 compr1
rlabel metal2 13754 5049 13754 5049 0 compr2
rlabel metal3 24457 12988 24457 12988 0 flash_adc_inp[0]
rlabel metal1 13708 6630 13708 6630 0 flash_adc_inp[10]
rlabel metal2 16790 7089 16790 7089 0 flash_adc_inp[11]
rlabel metal2 13386 4675 13386 4675 0 flash_adc_inp[12]
rlabel metal2 10350 2907 10350 2907 0 flash_adc_inp[13]
rlabel metal2 8510 2057 8510 2057 0 flash_adc_inp[14]
rlabel metal3 21099 10948 21099 10948 0 flash_adc_inp[1]
rlabel metal3 22249 10268 22249 10268 0 flash_adc_inp[2]
rlabel metal3 21697 11628 21697 11628 0 flash_adc_inp[3]
rlabel metal2 17710 11475 17710 11475 0 flash_adc_inp[4]
rlabel metal2 17250 8959 17250 8959 0 flash_adc_inp[5]
rlabel metal1 12696 10438 12696 10438 0 flash_adc_inp[6]
rlabel metal2 14950 7973 14950 7973 0 flash_adc_inp[7]
rlabel metal3 24549 8228 24549 8228 0 flash_adc_inp[8]
rlabel metal2 24518 11464 24518 11464 0 flash_adc_inp[9]
rlabel metal2 2162 6460 2162 6460 0 n122_o
rlabel metal1 5106 6256 5106 6256 0 n128_o
rlabel metal1 23230 7922 23230 7922 0 n135_o
rlabel metal1 4922 8942 4922 8942 0 n144_o
rlabel metal2 4002 5508 4002 5508 0 n150_o
rlabel metal1 6440 9690 6440 9690 0 n157_o
rlabel metal1 15686 9962 15686 9962 0 n166_o
rlabel metal1 14628 9894 14628 9894 0 n172_o
rlabel metal2 16790 9979 16790 9979 0 n179_o
rlabel metal2 14674 10404 14674 10404 0 n188_o
rlabel metal1 12604 3162 12604 3162 0 n194_o
rlabel metal2 12834 9826 12834 9826 0 n201_o
rlabel metal1 18630 10574 18630 10574 0 n210_o
rlabel metal2 19274 9622 19274 9622 0 n216_o
rlabel metal1 17710 8534 17710 8534 0 n223_o
rlabel metal2 17342 4403 17342 4403 0 net1
rlabel metal2 17434 9843 17434 9843 0 net10
rlabel metal2 21298 9962 21298 9962 0 net11
rlabel metal1 16330 8976 16330 8976 0 net12
rlabel metal1 22586 10030 22586 10030 0 net13
rlabel metal1 22218 8942 22218 8942 0 net14
rlabel metal1 22586 10676 22586 10676 0 net15
rlabel metal1 22954 8500 22954 8500 0 net16
rlabel metal1 22494 8500 22494 8500 0 net17
rlabel metal1 22310 9520 22310 9520 0 net18
rlabel metal2 22402 3111 22402 3111 0 net19
rlabel metal1 14168 5066 14168 5066 0 net2
rlabel metal2 1978 7344 1978 7344 0 net20
rlabel metal1 1656 6766 1656 6766 0 net21
rlabel metal1 9154 2448 9154 2448 0 net22
rlabel metal1 6210 2312 6210 2312 0 net23
rlabel metal1 12558 5576 12558 5576 0 net24
rlabel metal1 15134 10064 15134 10064 0 net25
rlabel metal2 13110 10302 13110 10302 0 net26
rlabel metal1 13202 10064 13202 10064 0 net27
rlabel metal1 20194 10098 20194 10098 0 net28
rlabel metal1 19366 10574 19366 10574 0 net29
rlabel metal1 14030 4454 14030 4454 0 net3
rlabel metal1 2231 5066 2231 5066 0 net30
rlabel metal1 8786 10030 8786 10030 0 net31
rlabel metal1 4416 2618 4416 2618 0 net32
rlabel metal1 5888 2618 5888 2618 0 net33
rlabel metal1 7958 2346 7958 2346 0 net34
rlabel metal1 8832 2618 8832 2618 0 net35
rlabel metal2 11730 2210 11730 2210 0 net36
rlabel metal2 11178 2244 11178 2244 0 net37
rlabel metal1 23046 4624 23046 4624 0 net38
rlabel metal1 12006 2380 12006 2380 0 net39
rlabel metal1 23138 8602 23138 8602 0 net4
rlabel metal1 11914 10676 11914 10676 0 net40
rlabel metal2 9522 2108 9522 2108 0 net41
rlabel metal2 10074 2142 10074 2142 0 net42
rlabel metal1 1840 6426 1840 6426 0 net43
rlabel metal1 13386 4760 13386 4760 0 net44
rlabel metal2 13938 10438 13938 10438 0 net45
rlabel metal2 17158 10574 17158 10574 0 net46
rlabel metal1 19872 9146 19872 9146 0 net47
rlabel metal1 18308 10234 18308 10234 0 net48
rlabel metal2 9982 10438 9982 10438 0 net49
rlabel metal2 22494 6119 22494 6119 0 net5
rlabel metal2 23046 8806 23046 8806 0 net50
rlabel metal1 1840 9690 1840 9690 0 net51
rlabel metal1 1840 5678 1840 5678 0 net52
rlabel metal2 1978 10438 1978 10438 0 net53
rlabel metal2 16514 10438 16514 10438 0 net54
rlabel metal2 12926 2873 12926 2873 0 net55
rlabel metal1 21160 7174 21160 7174 0 net56
rlabel metal1 14904 10642 14904 10642 0 net57
rlabel metal1 10948 2414 10948 2414 0 net58
rlabel metal1 16100 8942 16100 8942 0 net59
rlabel metal1 22586 3060 22586 3060 0 net6
rlabel metal1 23046 8976 23046 8976 0 net60
rlabel metal1 21160 8602 21160 8602 0 net61
rlabel metal2 18538 9860 18538 9860 0 net62
rlabel metal2 23230 5950 23230 5950 0 net63
rlabel metal1 21758 7514 21758 7514 0 net64
rlabel metal1 19366 2380 19366 2380 0 net65
rlabel metal2 19734 2142 19734 2142 0 net66
rlabel metal1 21206 7378 21206 7378 0 net67
rlabel metal2 21206 5950 21206 5950 0 net68
rlabel metal2 19734 4029 19734 4029 0 net69
rlabel metal1 23046 2958 23046 2958 0 net7
rlabel metal2 11546 4896 11546 4896 0 net70
rlabel metal1 11224 5338 11224 5338 0 net71
rlabel metal1 5520 5882 5520 5882 0 net72
rlabel metal1 8556 9554 8556 9554 0 net73
rlabel metal3 13202 2516 13202 2516 0 net74
rlabel metal2 13846 6630 13846 6630 0 net75
rlabel metal1 7636 7854 7636 7854 0 net76
rlabel metal1 6026 4250 6026 4250 0 net77
rlabel metal2 18998 2754 18998 2754 0 net78
rlabel metal1 5244 4114 5244 4114 0 net79
rlabel metal2 22908 6766 22908 6766 0 net8
rlabel metal1 8924 6766 8924 6766 0 net80
rlabel metal1 9729 6290 9729 6290 0 net81
rlabel metal1 5566 8976 5566 8976 0 net82
rlabel metal1 9338 2516 9338 2516 0 net83
rlabel metal1 1564 10574 1564 10574 0 net84
rlabel metal3 431 2788 431 2788 0 net85
rlabel metal2 9982 1462 9982 1462 0 net86
rlabel via2 16238 4029 16238 4029 0 net87
rlabel metal2 21942 6681 21942 6681 0 net88
rlabel metal1 18492 5882 18492 5882 0 net89
rlabel metal1 23230 5202 23230 5202 0 net9
rlabel metal2 20010 1282 20010 1282 0 rst_n
rlabel metal3 155 6868 155 6868 0 tern_dac[0]
rlabel metal1 14398 2822 14398 2822 0 tern_dac[10]
rlabel metal1 13938 10778 13938 10778 0 tern_dac[11]
rlabel metal1 16882 10778 16882 10778 0 tern_dac[12]
rlabel metal1 19458 10778 19458 10778 0 tern_dac[13]
rlabel metal1 17526 10778 17526 10778 0 tern_dac[14]
rlabel metal1 9798 10778 9798 10778 0 tern_dac[1]
rlabel metal1 22954 9350 22954 9350 0 tern_dac[2]
rlabel metal3 247 9588 247 9588 0 tern_dac[3]
rlabel metal3 431 5508 431 5508 0 tern_dac[4]
rlabel metal3 247 10268 247 10268 0 tern_dac[5]
rlabel metal1 16192 10506 16192 10506 0 tern_dac[6]
rlabel metal2 14858 874 14858 874 0 tern_dac[7]
rlabel metal2 21942 11770 21942 11770 0 tern_dac[8]
rlabel metal1 14996 10778 14996 10778 0 tern_dac[9]
rlabel metal2 11086 1768 11086 1768 0 ternff_conn
rlabel metal3 247 7548 247 7548 0 ui_in[0]
rlabel metal3 431 6188 431 6188 0 ui_in[1]
rlabel metal2 4554 1248 4554 1248 0 ui_in[2]
rlabel metal2 5198 687 5198 687 0 ui_in[3]
rlabel metal2 10994 11974 10994 11974 0 ui_in[4]
rlabel metal2 14214 12144 14214 12144 0 ui_in[5]
rlabel metal2 12926 11974 12926 11974 0 ui_in[6]
rlabel metal2 12282 11974 12282 11974 0 ui_in[7]
rlabel metal2 18078 12603 18078 12603 0 uio_in[0]
rlabel metal2 18722 12671 18722 12671 0 uio_in[1]
rlabel metal3 339 4828 339 4828 0 uio_in[2]
rlabel metal2 9062 11974 9062 11974 0 uio_in[3]
rlabel metal2 3910 1248 3910 1248 0 uio_in[4]
rlabel metal2 5842 1248 5842 1248 0 uio_in[5]
rlabel metal2 7130 1214 7130 1214 0 uio_in[6]
rlabel metal2 7774 1248 7774 1248 0 uio_in[7]
rlabel metal2 23230 13283 23230 13283 0 uo_out[0]
rlabel metal1 23552 9146 23552 9146 0 uo_out[1]
rlabel metal2 16974 10540 16974 10540 0 uo_out[2]
rlabel metal1 15548 10778 15548 10778 0 uo_out[3]
rlabel metal2 16146 10931 16146 10931 0 uo_out[4]
rlabel metal2 20194 13320 20194 13320 0 uo_out[5]
rlabel metal2 10534 1224 10534 1224 0 uo_out[6]
rlabel metal2 18722 704 18722 704 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 24752 13370
<< end >>
